module basic_1000_10000_1500_5_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_922,In_985);
nor U1 (N_1,In_839,In_285);
or U2 (N_2,In_717,In_485);
nor U3 (N_3,In_200,In_503);
xor U4 (N_4,In_257,In_518);
or U5 (N_5,In_446,In_670);
nand U6 (N_6,In_626,In_71);
or U7 (N_7,In_133,In_102);
or U8 (N_8,In_426,In_23);
or U9 (N_9,In_107,In_721);
xor U10 (N_10,In_59,In_984);
nand U11 (N_11,In_662,In_873);
nor U12 (N_12,In_676,In_854);
or U13 (N_13,In_522,In_810);
or U14 (N_14,In_265,In_313);
nand U15 (N_15,In_349,In_971);
xor U16 (N_16,In_920,In_496);
nor U17 (N_17,In_204,In_703);
nand U18 (N_18,In_648,In_126);
and U19 (N_19,In_284,In_163);
xor U20 (N_20,In_905,In_565);
nor U21 (N_21,In_665,In_630);
or U22 (N_22,In_547,In_977);
nor U23 (N_23,In_253,In_138);
nor U24 (N_24,In_412,In_712);
or U25 (N_25,In_802,In_444);
or U26 (N_26,In_814,In_668);
nand U27 (N_27,In_554,In_15);
nand U28 (N_28,In_291,In_220);
nor U29 (N_29,In_577,In_540);
nor U30 (N_30,In_956,In_923);
and U31 (N_31,In_781,In_369);
nor U32 (N_32,In_463,In_606);
nor U33 (N_33,In_599,In_884);
or U34 (N_34,In_889,In_797);
nor U35 (N_35,In_5,In_231);
xor U36 (N_36,In_340,In_413);
or U37 (N_37,In_436,In_302);
and U38 (N_38,In_762,In_916);
nand U39 (N_39,In_862,In_196);
xnor U40 (N_40,In_930,In_298);
nand U41 (N_41,In_545,In_729);
xor U42 (N_42,In_989,In_572);
nand U43 (N_43,In_562,In_11);
xor U44 (N_44,In_46,In_538);
nor U45 (N_45,In_707,In_710);
and U46 (N_46,In_590,In_202);
or U47 (N_47,In_568,In_634);
nand U48 (N_48,In_566,In_469);
or U49 (N_49,In_58,In_207);
and U50 (N_50,In_53,In_387);
xnor U51 (N_51,In_700,In_858);
nor U52 (N_52,In_720,In_639);
xnor U53 (N_53,In_143,In_264);
nand U54 (N_54,In_819,In_696);
xor U55 (N_55,In_63,In_788);
nor U56 (N_56,In_199,In_627);
nand U57 (N_57,In_435,In_746);
nor U58 (N_58,In_687,In_609);
or U59 (N_59,In_432,In_769);
nand U60 (N_60,In_942,In_723);
nand U61 (N_61,In_867,In_113);
nor U62 (N_62,In_124,In_287);
xor U63 (N_63,In_756,In_272);
nor U64 (N_64,In_954,In_56);
nor U65 (N_65,In_679,In_919);
or U66 (N_66,In_289,In_515);
nand U67 (N_67,In_316,In_718);
nor U68 (N_68,In_793,In_31);
or U69 (N_69,In_569,In_643);
nor U70 (N_70,In_119,In_787);
nand U71 (N_71,In_18,In_319);
and U72 (N_72,In_575,In_688);
xor U73 (N_73,In_10,In_417);
xnor U74 (N_74,In_421,In_322);
nand U75 (N_75,In_141,In_871);
nand U76 (N_76,In_821,In_449);
and U77 (N_77,In_683,In_130);
or U78 (N_78,In_224,In_753);
and U79 (N_79,In_212,In_669);
nand U80 (N_80,In_276,In_100);
or U81 (N_81,In_99,In_838);
xor U82 (N_82,In_980,In_418);
or U83 (N_83,In_471,In_438);
xor U84 (N_84,In_589,In_36);
and U85 (N_85,In_500,In_3);
nand U86 (N_86,In_238,In_188);
nor U87 (N_87,In_826,In_189);
and U88 (N_88,In_69,In_926);
xor U89 (N_89,In_403,In_524);
nand U90 (N_90,In_658,In_992);
and U91 (N_91,In_415,In_230);
nor U92 (N_92,In_872,In_972);
nor U93 (N_93,In_686,In_836);
nand U94 (N_94,In_362,In_906);
nor U95 (N_95,In_943,In_278);
xnor U96 (N_96,In_474,In_776);
nor U97 (N_97,In_256,In_663);
or U98 (N_98,In_692,In_636);
or U99 (N_99,In_976,In_945);
nand U100 (N_100,In_55,In_595);
nor U101 (N_101,In_935,In_168);
and U102 (N_102,In_527,In_571);
nor U103 (N_103,In_785,In_125);
nor U104 (N_104,In_135,In_335);
xor U105 (N_105,In_249,In_902);
nand U106 (N_106,In_760,In_892);
nor U107 (N_107,In_47,In_254);
or U108 (N_108,In_817,In_442);
nor U109 (N_109,In_334,In_422);
or U110 (N_110,In_437,In_849);
nand U111 (N_111,In_887,In_445);
nand U112 (N_112,In_573,In_528);
nand U113 (N_113,In_352,In_743);
and U114 (N_114,In_65,In_22);
xnor U115 (N_115,In_150,In_666);
xnor U116 (N_116,In_526,In_592);
nor U117 (N_117,In_675,In_644);
and U118 (N_118,In_560,In_782);
nor U119 (N_119,In_931,In_991);
and U120 (N_120,In_965,In_8);
xnor U121 (N_121,In_811,In_890);
xor U122 (N_122,In_812,In_304);
nand U123 (N_123,In_127,In_516);
nor U124 (N_124,In_139,In_542);
nor U125 (N_125,In_879,In_653);
and U126 (N_126,In_103,In_271);
and U127 (N_127,In_731,In_921);
or U128 (N_128,In_384,In_179);
nor U129 (N_129,In_677,In_633);
nand U130 (N_130,In_341,In_117);
and U131 (N_131,In_391,In_146);
xnor U132 (N_132,In_784,In_363);
and U133 (N_133,In_678,In_217);
xnor U134 (N_134,In_318,In_738);
nor U135 (N_135,In_364,In_702);
nand U136 (N_136,In_358,In_73);
xnor U137 (N_137,In_949,In_79);
or U138 (N_138,In_185,In_973);
or U139 (N_139,In_534,In_519);
xor U140 (N_140,In_619,In_244);
xor U141 (N_141,In_451,In_80);
and U142 (N_142,In_396,In_374);
nand U143 (N_143,In_958,In_295);
nand U144 (N_144,In_689,In_19);
nor U145 (N_145,In_7,In_924);
nor U146 (N_146,In_145,In_600);
nand U147 (N_147,In_452,In_90);
nor U148 (N_148,In_536,In_306);
nor U149 (N_149,In_275,In_321);
nor U150 (N_150,In_122,In_880);
or U151 (N_151,In_457,In_529);
and U152 (N_152,In_732,In_98);
xor U153 (N_153,In_680,In_282);
or U154 (N_154,In_95,In_464);
nand U155 (N_155,In_288,In_852);
nor U156 (N_156,In_280,In_398);
nand U157 (N_157,In_118,In_243);
xnor U158 (N_158,In_48,In_114);
and U159 (N_159,In_567,In_739);
nor U160 (N_160,In_928,In_758);
nand U161 (N_161,In_27,In_376);
and U162 (N_162,In_397,In_402);
and U163 (N_163,In_561,In_440);
xor U164 (N_164,In_941,In_624);
and U165 (N_165,In_510,In_62);
xor U166 (N_166,In_994,In_894);
and U167 (N_167,In_234,In_766);
and U168 (N_168,In_29,In_13);
nand U169 (N_169,In_314,In_470);
xnor U170 (N_170,In_44,In_245);
or U171 (N_171,In_214,In_531);
xnor U172 (N_172,In_443,In_730);
and U173 (N_173,In_74,In_162);
xor U174 (N_174,In_78,In_587);
or U175 (N_175,In_39,In_960);
or U176 (N_176,In_764,In_864);
xor U177 (N_177,In_883,In_727);
and U178 (N_178,In_638,In_621);
nand U179 (N_179,In_49,In_995);
and U180 (N_180,In_734,In_975);
nor U181 (N_181,In_290,In_908);
nor U182 (N_182,In_458,In_998);
nand U183 (N_183,In_848,In_336);
nand U184 (N_184,In_171,In_157);
and U185 (N_185,In_917,In_885);
and U186 (N_186,In_165,In_343);
xnor U187 (N_187,In_448,In_629);
nor U188 (N_188,In_667,In_828);
or U189 (N_189,In_128,In_351);
and U190 (N_190,In_181,In_974);
or U191 (N_191,In_94,In_549);
and U192 (N_192,In_136,In_326);
or U193 (N_193,In_14,In_347);
nand U194 (N_194,In_856,In_355);
xnor U195 (N_195,In_281,In_110);
nor U196 (N_196,In_481,In_886);
and U197 (N_197,In_419,In_927);
nand U198 (N_198,In_876,In_969);
nand U199 (N_199,In_307,In_881);
nand U200 (N_200,In_106,In_578);
and U201 (N_201,In_151,In_770);
or U202 (N_202,In_808,In_115);
or U203 (N_203,In_570,In_618);
nor U204 (N_204,In_952,In_87);
xnor U205 (N_205,In_877,In_532);
nand U206 (N_206,In_901,In_88);
and U207 (N_207,In_851,In_725);
xor U208 (N_208,In_392,In_105);
and U209 (N_209,In_192,In_375);
and U210 (N_210,In_434,In_216);
nand U211 (N_211,In_303,In_733);
nor U212 (N_212,In_76,In_695);
xnor U213 (N_213,In_754,In_903);
and U214 (N_214,In_865,In_612);
or U215 (N_215,In_601,In_713);
xnor U216 (N_216,In_193,In_682);
or U217 (N_217,In_85,In_719);
xor U218 (N_218,In_201,In_967);
and U219 (N_219,In_799,In_409);
and U220 (N_220,In_197,In_17);
or U221 (N_221,In_430,In_365);
and U222 (N_222,In_860,In_24);
nor U223 (N_223,In_914,In_671);
nor U224 (N_224,In_804,In_140);
and U225 (N_225,In_716,In_613);
nor U226 (N_226,In_623,In_91);
nor U227 (N_227,In_246,In_299);
nand U228 (N_228,In_2,In_775);
and U229 (N_229,In_955,In_382);
nor U230 (N_230,In_933,In_827);
nor U231 (N_231,In_475,In_323);
and U232 (N_232,In_360,In_656);
and U233 (N_233,In_320,In_455);
nand U234 (N_234,In_897,In_407);
nor U235 (N_235,In_938,In_904);
nor U236 (N_236,In_649,In_581);
or U237 (N_237,In_383,In_112);
nor U238 (N_238,In_891,In_513);
and U239 (N_239,In_997,In_64);
or U240 (N_240,In_43,In_232);
nor U241 (N_241,In_54,In_778);
xnor U242 (N_242,In_946,In_142);
nand U243 (N_243,In_737,In_68);
nor U244 (N_244,In_585,In_332);
xnor U245 (N_245,In_129,In_959);
xnor U246 (N_246,In_0,In_714);
nor U247 (N_247,In_843,In_504);
nand U248 (N_248,In_424,In_594);
xnor U249 (N_249,In_868,In_439);
nor U250 (N_250,In_664,In_72);
or U251 (N_251,In_774,In_96);
and U252 (N_252,In_429,In_479);
and U253 (N_253,In_465,In_537);
nand U254 (N_254,In_741,In_354);
or U255 (N_255,In_704,In_750);
xnor U256 (N_256,In_605,In_411);
nand U257 (N_257,In_310,In_489);
xnor U258 (N_258,In_616,In_493);
xor U259 (N_259,In_484,In_936);
nor U260 (N_260,In_724,In_400);
and U261 (N_261,In_252,In_416);
and U262 (N_262,In_203,In_308);
nor U263 (N_263,In_711,In_986);
xnor U264 (N_264,In_647,In_357);
and U265 (N_265,In_805,In_981);
nor U266 (N_266,In_806,In_361);
xnor U267 (N_267,In_807,In_657);
nand U268 (N_268,In_833,In_556);
and U269 (N_269,In_350,In_175);
or U270 (N_270,In_52,In_213);
xnor U271 (N_271,In_453,In_480);
xnor U272 (N_272,In_237,In_178);
nand U273 (N_273,In_502,In_507);
or U274 (N_274,In_506,In_89);
xor U275 (N_275,In_498,In_459);
nor U276 (N_276,In_296,In_301);
nor U277 (N_277,In_339,In_698);
nor U278 (N_278,In_30,In_292);
nand U279 (N_279,In_222,In_1);
and U280 (N_280,In_511,In_247);
and U281 (N_281,In_359,In_968);
xnor U282 (N_282,In_353,In_261);
xnor U283 (N_283,In_28,In_116);
or U284 (N_284,In_9,In_267);
nor U285 (N_285,In_912,In_370);
or U286 (N_286,In_944,In_765);
xor U287 (N_287,In_962,In_508);
nor U288 (N_288,In_109,In_158);
nor U289 (N_289,In_255,In_584);
xnor U290 (N_290,In_993,In_517);
and U291 (N_291,In_75,In_789);
or U292 (N_292,In_597,In_239);
nand U293 (N_293,In_603,In_837);
and U294 (N_294,In_86,In_32);
xor U295 (N_295,In_790,In_845);
or U296 (N_296,In_552,In_167);
and U297 (N_297,In_937,In_913);
xor U298 (N_298,In_466,In_777);
and U299 (N_299,In_651,In_205);
xor U300 (N_300,In_184,In_131);
nor U301 (N_301,In_690,In_483);
nand U302 (N_302,In_539,In_441);
and U303 (N_303,In_487,In_652);
nand U304 (N_304,In_389,In_641);
or U305 (N_305,In_970,In_368);
nand U306 (N_306,In_899,In_961);
nor U307 (N_307,In_38,In_558);
nand U308 (N_308,In_911,In_154);
and U309 (N_309,In_366,In_691);
xor U310 (N_310,In_433,In_16);
xor U311 (N_311,In_820,In_66);
or U312 (N_312,In_588,In_497);
nor U313 (N_313,In_274,In_478);
nand U314 (N_314,In_697,In_227);
nand U315 (N_315,In_248,In_210);
xnor U316 (N_316,In_344,In_84);
nor U317 (N_317,In_408,In_694);
or U318 (N_318,In_874,In_742);
or U319 (N_319,In_604,In_57);
xor U320 (N_320,In_541,In_715);
and U321 (N_321,In_798,In_215);
nor U322 (N_322,In_509,In_918);
nand U323 (N_323,In_543,In_614);
nor U324 (N_324,In_462,In_579);
or U325 (N_325,In_783,In_219);
nor U326 (N_326,In_685,In_324);
or U327 (N_327,In_505,In_460);
nand U328 (N_328,In_177,In_759);
or U329 (N_329,In_525,In_70);
nand U330 (N_330,In_813,In_187);
xnor U331 (N_331,In_104,In_144);
nor U332 (N_332,In_866,In_544);
nand U333 (N_333,In_198,In_829);
and U334 (N_334,In_794,In_208);
nor U335 (N_335,In_598,In_423);
nand U336 (N_336,In_786,In_632);
xor U337 (N_337,In_377,In_780);
xor U338 (N_338,In_608,In_186);
xnor U339 (N_339,In_841,In_371);
or U340 (N_340,In_659,In_454);
xor U341 (N_341,In_815,In_660);
or U342 (N_342,In_134,In_425);
nor U343 (N_343,In_747,In_45);
nor U344 (N_344,In_473,In_427);
nor U345 (N_345,In_863,In_34);
xor U346 (N_346,In_241,In_939);
and U347 (N_347,In_315,In_378);
nand U348 (N_348,In_111,In_240);
nand U349 (N_349,In_611,In_751);
nor U350 (N_350,In_499,In_393);
and U351 (N_351,In_132,In_932);
nor U352 (N_352,In_35,In_4);
or U353 (N_353,In_490,In_262);
or U354 (N_354,In_831,In_620);
or U355 (N_355,In_631,In_190);
xnor U356 (N_356,In_492,In_591);
or U357 (N_357,In_878,In_850);
and U358 (N_358,In_228,In_191);
xor U359 (N_359,In_842,In_467);
nor U360 (N_360,In_859,In_486);
nand U361 (N_361,In_576,In_385);
xor U362 (N_362,In_550,In_172);
or U363 (N_363,In_895,In_101);
nand U364 (N_364,In_6,In_218);
or U365 (N_365,In_169,In_844);
xor U366 (N_366,In_800,In_159);
or U367 (N_367,In_963,In_259);
nor U368 (N_368,In_900,In_211);
nand U369 (N_369,In_494,In_174);
or U370 (N_370,In_940,In_748);
or U371 (N_371,In_832,In_661);
or U372 (N_372,In_950,In_728);
nand U373 (N_373,In_999,In_996);
nor U374 (N_374,In_37,In_97);
nor U375 (N_375,In_607,In_21);
xnor U376 (N_376,In_297,In_855);
and U377 (N_377,In_555,In_520);
or U378 (N_378,In_580,In_147);
and U379 (N_379,In_840,In_223);
nand U380 (N_380,In_673,In_672);
and U381 (N_381,In_978,In_166);
xnor U382 (N_382,In_206,In_521);
and U383 (N_383,In_152,In_233);
and U384 (N_384,In_269,In_381);
xor U385 (N_385,In_847,In_761);
and U386 (N_386,In_964,In_557);
nor U387 (N_387,In_20,In_564);
or U388 (N_388,In_835,In_273);
xor U389 (N_389,In_771,In_286);
or U390 (N_390,In_684,In_948);
xnor U391 (N_391,In_910,In_226);
xnor U392 (N_392,In_642,In_929);
or U393 (N_393,In_512,In_283);
and U394 (N_394,In_176,In_325);
and U395 (N_395,In_987,In_757);
nor U396 (N_396,In_796,In_801);
and U397 (N_397,In_160,In_722);
or U398 (N_398,In_153,In_242);
or U399 (N_399,In_779,In_268);
or U400 (N_400,In_530,In_752);
nor U401 (N_401,In_818,In_60);
xor U402 (N_402,In_149,In_553);
and U403 (N_403,In_602,In_472);
xor U404 (N_404,In_164,In_610);
nand U405 (N_405,In_461,In_482);
nand U406 (N_406,In_348,In_294);
xnor U407 (N_407,In_450,In_693);
or U408 (N_408,In_559,In_395);
nor U409 (N_409,In_251,In_983);
xor U410 (N_410,In_477,In_533);
nand U411 (N_411,In_650,In_394);
nor U412 (N_412,In_583,In_83);
xnor U413 (N_413,In_26,In_979);
nor U414 (N_414,In_235,In_250);
nor U415 (N_415,In_311,In_346);
nor U416 (N_416,In_50,In_735);
nand U417 (N_417,In_121,In_373);
xnor U418 (N_418,In_655,In_535);
and U419 (N_419,In_12,In_236);
and U420 (N_420,In_951,In_229);
nand U421 (N_421,In_404,In_338);
nor U422 (N_422,In_744,In_414);
nor U423 (N_423,In_92,In_356);
and U424 (N_424,In_947,In_329);
xnor U425 (N_425,In_681,In_825);
and U426 (N_426,In_401,In_934);
nor U427 (N_427,In_342,In_915);
or U428 (N_428,In_82,In_622);
and U429 (N_429,In_263,In_763);
or U430 (N_430,In_309,In_420);
and U431 (N_431,In_898,In_882);
and U432 (N_432,In_857,In_637);
nand U433 (N_433,In_745,In_646);
and U434 (N_434,In_888,In_51);
or U435 (N_435,In_42,In_156);
or U436 (N_436,In_699,In_551);
nor U437 (N_437,In_41,In_654);
nor U438 (N_438,In_279,In_593);
or U439 (N_439,In_574,In_399);
nand U440 (N_440,In_740,In_331);
and U441 (N_441,In_803,In_170);
nor U442 (N_442,In_221,In_792);
and U443 (N_443,In_456,In_925);
or U444 (N_444,In_330,In_406);
xor U445 (N_445,In_182,In_834);
xnor U446 (N_446,In_277,In_982);
xor U447 (N_447,In_755,In_491);
nand U448 (N_448,In_327,In_173);
nor U449 (N_449,In_388,In_488);
and U450 (N_450,In_645,In_108);
and U451 (N_451,In_736,In_615);
xor U452 (N_452,In_768,In_773);
nand U453 (N_453,In_380,In_137);
nand U454 (N_454,In_791,In_345);
and U455 (N_455,In_816,In_120);
xnor U456 (N_456,In_195,In_405);
and U457 (N_457,In_337,In_386);
nor U458 (N_458,In_333,In_596);
nor U459 (N_459,In_225,In_328);
nor U460 (N_460,In_809,In_180);
and U461 (N_461,In_548,In_183);
and U462 (N_462,In_640,In_701);
or U463 (N_463,In_953,In_767);
nor U464 (N_464,In_25,In_266);
and U465 (N_465,In_447,In_390);
or U466 (N_466,In_822,In_312);
nor U467 (N_467,In_869,In_379);
and U468 (N_468,In_617,In_846);
nand U469 (N_469,In_123,In_305);
or U470 (N_470,In_628,In_966);
xor U471 (N_471,In_148,In_957);
and U472 (N_472,In_81,In_270);
and U473 (N_473,In_372,In_909);
and U474 (N_474,In_772,In_33);
nor U475 (N_475,In_61,In_705);
nor U476 (N_476,In_428,In_875);
nor U477 (N_477,In_907,In_431);
xnor U478 (N_478,In_67,In_209);
or U479 (N_479,In_861,In_824);
or U480 (N_480,In_990,In_635);
xor U481 (N_481,In_709,In_830);
xnor U482 (N_482,In_870,In_706);
or U483 (N_483,In_501,In_161);
nor U484 (N_484,In_300,In_523);
nor U485 (N_485,In_40,In_155);
and U486 (N_486,In_410,In_563);
xnor U487 (N_487,In_795,In_674);
or U488 (N_488,In_194,In_586);
nand U489 (N_489,In_988,In_546);
and U490 (N_490,In_77,In_367);
or U491 (N_491,In_582,In_896);
nor U492 (N_492,In_625,In_93);
nor U493 (N_493,In_708,In_495);
xnor U494 (N_494,In_749,In_468);
and U495 (N_495,In_258,In_853);
nor U496 (N_496,In_260,In_514);
or U497 (N_497,In_476,In_293);
or U498 (N_498,In_893,In_823);
nor U499 (N_499,In_726,In_317);
and U500 (N_500,In_718,In_975);
or U501 (N_501,In_535,In_505);
nand U502 (N_502,In_581,In_242);
and U503 (N_503,In_603,In_881);
and U504 (N_504,In_191,In_562);
nand U505 (N_505,In_271,In_967);
and U506 (N_506,In_991,In_947);
nor U507 (N_507,In_97,In_938);
xnor U508 (N_508,In_894,In_657);
or U509 (N_509,In_996,In_442);
xnor U510 (N_510,In_315,In_376);
xor U511 (N_511,In_306,In_734);
and U512 (N_512,In_714,In_648);
xor U513 (N_513,In_954,In_261);
nand U514 (N_514,In_725,In_574);
nand U515 (N_515,In_46,In_686);
or U516 (N_516,In_683,In_793);
or U517 (N_517,In_130,In_517);
nor U518 (N_518,In_830,In_160);
nand U519 (N_519,In_407,In_805);
xnor U520 (N_520,In_622,In_677);
nor U521 (N_521,In_609,In_329);
nand U522 (N_522,In_655,In_252);
or U523 (N_523,In_142,In_747);
xor U524 (N_524,In_826,In_438);
and U525 (N_525,In_416,In_68);
or U526 (N_526,In_183,In_394);
nand U527 (N_527,In_982,In_763);
or U528 (N_528,In_957,In_973);
nand U529 (N_529,In_411,In_295);
and U530 (N_530,In_116,In_791);
or U531 (N_531,In_670,In_877);
nor U532 (N_532,In_759,In_91);
xnor U533 (N_533,In_514,In_26);
xnor U534 (N_534,In_68,In_115);
nand U535 (N_535,In_898,In_980);
nand U536 (N_536,In_170,In_476);
nand U537 (N_537,In_218,In_470);
nand U538 (N_538,In_614,In_522);
and U539 (N_539,In_759,In_757);
or U540 (N_540,In_914,In_120);
and U541 (N_541,In_879,In_698);
nor U542 (N_542,In_782,In_224);
or U543 (N_543,In_847,In_177);
and U544 (N_544,In_0,In_959);
nor U545 (N_545,In_390,In_119);
nand U546 (N_546,In_272,In_336);
nand U547 (N_547,In_639,In_175);
xnor U548 (N_548,In_793,In_603);
or U549 (N_549,In_597,In_47);
xnor U550 (N_550,In_333,In_135);
nand U551 (N_551,In_361,In_157);
or U552 (N_552,In_567,In_611);
and U553 (N_553,In_42,In_350);
xnor U554 (N_554,In_922,In_656);
xor U555 (N_555,In_462,In_215);
or U556 (N_556,In_105,In_296);
or U557 (N_557,In_883,In_873);
nor U558 (N_558,In_164,In_860);
nand U559 (N_559,In_650,In_679);
xor U560 (N_560,In_769,In_765);
xor U561 (N_561,In_650,In_5);
nor U562 (N_562,In_154,In_172);
xnor U563 (N_563,In_414,In_992);
nand U564 (N_564,In_289,In_525);
or U565 (N_565,In_406,In_213);
nand U566 (N_566,In_846,In_121);
and U567 (N_567,In_976,In_274);
or U568 (N_568,In_553,In_648);
nand U569 (N_569,In_939,In_246);
or U570 (N_570,In_492,In_103);
nor U571 (N_571,In_466,In_580);
xnor U572 (N_572,In_728,In_771);
or U573 (N_573,In_809,In_169);
nand U574 (N_574,In_824,In_576);
nor U575 (N_575,In_403,In_734);
nand U576 (N_576,In_907,In_868);
nor U577 (N_577,In_455,In_88);
nor U578 (N_578,In_434,In_994);
nor U579 (N_579,In_25,In_316);
and U580 (N_580,In_865,In_777);
and U581 (N_581,In_324,In_401);
nand U582 (N_582,In_474,In_87);
or U583 (N_583,In_100,In_395);
nor U584 (N_584,In_71,In_370);
and U585 (N_585,In_72,In_369);
xnor U586 (N_586,In_197,In_183);
nand U587 (N_587,In_83,In_745);
xor U588 (N_588,In_360,In_100);
xor U589 (N_589,In_33,In_641);
nand U590 (N_590,In_324,In_926);
nor U591 (N_591,In_789,In_496);
nor U592 (N_592,In_919,In_967);
xnor U593 (N_593,In_517,In_950);
nand U594 (N_594,In_314,In_563);
nor U595 (N_595,In_761,In_450);
nor U596 (N_596,In_304,In_432);
or U597 (N_597,In_930,In_941);
or U598 (N_598,In_558,In_301);
nand U599 (N_599,In_300,In_799);
xor U600 (N_600,In_967,In_202);
xor U601 (N_601,In_515,In_444);
or U602 (N_602,In_996,In_313);
or U603 (N_603,In_107,In_8);
nand U604 (N_604,In_37,In_975);
nand U605 (N_605,In_640,In_399);
xnor U606 (N_606,In_575,In_190);
and U607 (N_607,In_717,In_832);
and U608 (N_608,In_395,In_692);
nand U609 (N_609,In_304,In_392);
xor U610 (N_610,In_51,In_738);
or U611 (N_611,In_660,In_277);
nand U612 (N_612,In_679,In_796);
or U613 (N_613,In_762,In_181);
nor U614 (N_614,In_98,In_347);
and U615 (N_615,In_402,In_594);
and U616 (N_616,In_959,In_579);
nor U617 (N_617,In_502,In_337);
or U618 (N_618,In_668,In_974);
nand U619 (N_619,In_302,In_327);
nand U620 (N_620,In_324,In_175);
nor U621 (N_621,In_336,In_801);
nand U622 (N_622,In_147,In_774);
xnor U623 (N_623,In_340,In_240);
or U624 (N_624,In_78,In_555);
nor U625 (N_625,In_806,In_894);
or U626 (N_626,In_606,In_27);
nor U627 (N_627,In_81,In_767);
nor U628 (N_628,In_195,In_976);
or U629 (N_629,In_527,In_941);
or U630 (N_630,In_986,In_535);
and U631 (N_631,In_926,In_606);
or U632 (N_632,In_266,In_963);
nand U633 (N_633,In_790,In_473);
or U634 (N_634,In_647,In_421);
xor U635 (N_635,In_673,In_14);
nand U636 (N_636,In_678,In_965);
xor U637 (N_637,In_141,In_571);
or U638 (N_638,In_482,In_427);
and U639 (N_639,In_991,In_545);
or U640 (N_640,In_65,In_222);
nand U641 (N_641,In_844,In_469);
or U642 (N_642,In_831,In_431);
and U643 (N_643,In_917,In_181);
nor U644 (N_644,In_241,In_117);
nor U645 (N_645,In_351,In_864);
and U646 (N_646,In_558,In_918);
or U647 (N_647,In_195,In_879);
and U648 (N_648,In_456,In_323);
nand U649 (N_649,In_499,In_256);
nor U650 (N_650,In_406,In_262);
xnor U651 (N_651,In_963,In_923);
or U652 (N_652,In_159,In_336);
or U653 (N_653,In_616,In_22);
and U654 (N_654,In_744,In_122);
nor U655 (N_655,In_775,In_258);
or U656 (N_656,In_658,In_382);
xor U657 (N_657,In_765,In_312);
or U658 (N_658,In_764,In_599);
nor U659 (N_659,In_357,In_801);
nor U660 (N_660,In_685,In_773);
xnor U661 (N_661,In_887,In_812);
nor U662 (N_662,In_600,In_219);
nand U663 (N_663,In_60,In_425);
xnor U664 (N_664,In_157,In_94);
xor U665 (N_665,In_7,In_766);
xnor U666 (N_666,In_473,In_955);
or U667 (N_667,In_376,In_759);
nand U668 (N_668,In_40,In_515);
and U669 (N_669,In_244,In_151);
xnor U670 (N_670,In_483,In_807);
and U671 (N_671,In_542,In_116);
and U672 (N_672,In_371,In_331);
nor U673 (N_673,In_803,In_475);
nand U674 (N_674,In_94,In_402);
nor U675 (N_675,In_553,In_577);
nand U676 (N_676,In_38,In_901);
and U677 (N_677,In_611,In_585);
nand U678 (N_678,In_560,In_888);
nor U679 (N_679,In_988,In_165);
xnor U680 (N_680,In_196,In_315);
or U681 (N_681,In_617,In_969);
or U682 (N_682,In_59,In_3);
and U683 (N_683,In_544,In_600);
nand U684 (N_684,In_685,In_140);
or U685 (N_685,In_617,In_671);
and U686 (N_686,In_540,In_648);
and U687 (N_687,In_602,In_999);
and U688 (N_688,In_674,In_967);
or U689 (N_689,In_78,In_576);
or U690 (N_690,In_466,In_472);
nand U691 (N_691,In_530,In_674);
xnor U692 (N_692,In_910,In_555);
or U693 (N_693,In_688,In_91);
xnor U694 (N_694,In_794,In_230);
xnor U695 (N_695,In_249,In_569);
or U696 (N_696,In_150,In_73);
xor U697 (N_697,In_493,In_302);
xnor U698 (N_698,In_800,In_289);
or U699 (N_699,In_501,In_939);
xnor U700 (N_700,In_555,In_548);
and U701 (N_701,In_769,In_205);
nand U702 (N_702,In_592,In_340);
xnor U703 (N_703,In_790,In_233);
nor U704 (N_704,In_323,In_904);
or U705 (N_705,In_28,In_960);
or U706 (N_706,In_376,In_876);
nand U707 (N_707,In_576,In_600);
and U708 (N_708,In_392,In_890);
and U709 (N_709,In_869,In_355);
nand U710 (N_710,In_278,In_21);
xor U711 (N_711,In_925,In_692);
and U712 (N_712,In_774,In_720);
nand U713 (N_713,In_748,In_921);
or U714 (N_714,In_735,In_702);
nand U715 (N_715,In_576,In_622);
nor U716 (N_716,In_48,In_712);
xor U717 (N_717,In_491,In_722);
or U718 (N_718,In_926,In_726);
nor U719 (N_719,In_796,In_646);
nand U720 (N_720,In_940,In_312);
nor U721 (N_721,In_223,In_138);
and U722 (N_722,In_45,In_382);
nand U723 (N_723,In_205,In_850);
or U724 (N_724,In_748,In_924);
nand U725 (N_725,In_867,In_191);
nor U726 (N_726,In_813,In_985);
nand U727 (N_727,In_970,In_719);
and U728 (N_728,In_363,In_984);
or U729 (N_729,In_19,In_393);
nand U730 (N_730,In_891,In_381);
nor U731 (N_731,In_792,In_846);
nor U732 (N_732,In_763,In_361);
xor U733 (N_733,In_43,In_274);
nor U734 (N_734,In_345,In_517);
and U735 (N_735,In_382,In_785);
xor U736 (N_736,In_540,In_646);
or U737 (N_737,In_459,In_371);
nor U738 (N_738,In_227,In_976);
nor U739 (N_739,In_648,In_201);
nand U740 (N_740,In_83,In_768);
and U741 (N_741,In_64,In_97);
or U742 (N_742,In_172,In_791);
xor U743 (N_743,In_778,In_220);
nand U744 (N_744,In_305,In_361);
or U745 (N_745,In_610,In_863);
xor U746 (N_746,In_720,In_380);
or U747 (N_747,In_280,In_916);
or U748 (N_748,In_710,In_165);
nand U749 (N_749,In_121,In_337);
nand U750 (N_750,In_208,In_822);
nor U751 (N_751,In_493,In_982);
nor U752 (N_752,In_785,In_673);
or U753 (N_753,In_543,In_66);
nand U754 (N_754,In_567,In_371);
nor U755 (N_755,In_709,In_127);
nor U756 (N_756,In_526,In_262);
nor U757 (N_757,In_291,In_12);
xnor U758 (N_758,In_352,In_944);
or U759 (N_759,In_874,In_397);
nor U760 (N_760,In_525,In_885);
nand U761 (N_761,In_460,In_658);
or U762 (N_762,In_350,In_78);
nand U763 (N_763,In_60,In_247);
nor U764 (N_764,In_236,In_45);
and U765 (N_765,In_704,In_264);
xnor U766 (N_766,In_553,In_903);
or U767 (N_767,In_240,In_936);
nor U768 (N_768,In_700,In_328);
or U769 (N_769,In_827,In_792);
nand U770 (N_770,In_69,In_218);
and U771 (N_771,In_199,In_891);
nor U772 (N_772,In_552,In_883);
or U773 (N_773,In_829,In_787);
nand U774 (N_774,In_431,In_30);
or U775 (N_775,In_178,In_174);
or U776 (N_776,In_532,In_28);
nor U777 (N_777,In_377,In_524);
and U778 (N_778,In_669,In_825);
nor U779 (N_779,In_610,In_249);
and U780 (N_780,In_637,In_942);
or U781 (N_781,In_949,In_510);
nand U782 (N_782,In_394,In_47);
or U783 (N_783,In_153,In_975);
or U784 (N_784,In_888,In_234);
and U785 (N_785,In_81,In_2);
or U786 (N_786,In_460,In_498);
xnor U787 (N_787,In_311,In_543);
xnor U788 (N_788,In_543,In_911);
nand U789 (N_789,In_41,In_474);
or U790 (N_790,In_79,In_224);
xor U791 (N_791,In_902,In_959);
xnor U792 (N_792,In_122,In_865);
xnor U793 (N_793,In_830,In_110);
nor U794 (N_794,In_389,In_966);
xnor U795 (N_795,In_887,In_596);
xnor U796 (N_796,In_193,In_277);
and U797 (N_797,In_639,In_967);
nor U798 (N_798,In_926,In_720);
and U799 (N_799,In_320,In_155);
or U800 (N_800,In_884,In_822);
or U801 (N_801,In_159,In_453);
nor U802 (N_802,In_22,In_729);
and U803 (N_803,In_545,In_684);
nor U804 (N_804,In_532,In_881);
xor U805 (N_805,In_120,In_618);
xnor U806 (N_806,In_590,In_719);
nor U807 (N_807,In_591,In_25);
nand U808 (N_808,In_377,In_590);
nand U809 (N_809,In_812,In_367);
xor U810 (N_810,In_881,In_296);
or U811 (N_811,In_697,In_724);
xor U812 (N_812,In_473,In_255);
and U813 (N_813,In_756,In_366);
and U814 (N_814,In_394,In_756);
nor U815 (N_815,In_309,In_808);
xor U816 (N_816,In_498,In_561);
xor U817 (N_817,In_670,In_188);
or U818 (N_818,In_302,In_238);
and U819 (N_819,In_836,In_106);
or U820 (N_820,In_196,In_559);
nand U821 (N_821,In_72,In_402);
and U822 (N_822,In_486,In_268);
nor U823 (N_823,In_465,In_713);
xor U824 (N_824,In_565,In_11);
nand U825 (N_825,In_838,In_230);
or U826 (N_826,In_509,In_570);
xor U827 (N_827,In_151,In_813);
nor U828 (N_828,In_949,In_679);
nand U829 (N_829,In_921,In_147);
and U830 (N_830,In_611,In_360);
nand U831 (N_831,In_608,In_5);
xor U832 (N_832,In_760,In_49);
nor U833 (N_833,In_967,In_821);
xor U834 (N_834,In_747,In_487);
xnor U835 (N_835,In_860,In_531);
nand U836 (N_836,In_663,In_426);
nor U837 (N_837,In_120,In_636);
nand U838 (N_838,In_803,In_783);
or U839 (N_839,In_87,In_733);
or U840 (N_840,In_495,In_834);
nor U841 (N_841,In_96,In_862);
and U842 (N_842,In_913,In_172);
nand U843 (N_843,In_634,In_828);
and U844 (N_844,In_922,In_908);
xnor U845 (N_845,In_927,In_718);
nand U846 (N_846,In_907,In_231);
or U847 (N_847,In_191,In_634);
nand U848 (N_848,In_512,In_562);
and U849 (N_849,In_512,In_847);
nand U850 (N_850,In_10,In_307);
nand U851 (N_851,In_990,In_906);
nor U852 (N_852,In_63,In_64);
nor U853 (N_853,In_36,In_238);
nor U854 (N_854,In_103,In_638);
nand U855 (N_855,In_713,In_468);
nor U856 (N_856,In_971,In_527);
nor U857 (N_857,In_33,In_207);
nand U858 (N_858,In_401,In_80);
xnor U859 (N_859,In_317,In_856);
xor U860 (N_860,In_776,In_181);
and U861 (N_861,In_411,In_400);
nand U862 (N_862,In_165,In_211);
and U863 (N_863,In_893,In_3);
and U864 (N_864,In_840,In_883);
and U865 (N_865,In_931,In_975);
or U866 (N_866,In_818,In_402);
nand U867 (N_867,In_599,In_456);
nor U868 (N_868,In_913,In_884);
xnor U869 (N_869,In_767,In_467);
xor U870 (N_870,In_241,In_490);
and U871 (N_871,In_611,In_702);
and U872 (N_872,In_50,In_471);
nand U873 (N_873,In_291,In_678);
nor U874 (N_874,In_480,In_214);
nand U875 (N_875,In_700,In_599);
nand U876 (N_876,In_661,In_708);
and U877 (N_877,In_704,In_902);
and U878 (N_878,In_618,In_595);
nor U879 (N_879,In_224,In_352);
xnor U880 (N_880,In_765,In_380);
nand U881 (N_881,In_481,In_525);
or U882 (N_882,In_333,In_367);
xnor U883 (N_883,In_92,In_157);
xor U884 (N_884,In_889,In_925);
and U885 (N_885,In_422,In_113);
xnor U886 (N_886,In_214,In_991);
nand U887 (N_887,In_480,In_539);
nand U888 (N_888,In_473,In_705);
nor U889 (N_889,In_154,In_914);
xnor U890 (N_890,In_559,In_882);
and U891 (N_891,In_114,In_819);
or U892 (N_892,In_692,In_65);
and U893 (N_893,In_597,In_366);
nor U894 (N_894,In_578,In_219);
and U895 (N_895,In_73,In_244);
nand U896 (N_896,In_15,In_537);
or U897 (N_897,In_304,In_800);
nor U898 (N_898,In_553,In_270);
nor U899 (N_899,In_373,In_890);
nand U900 (N_900,In_284,In_456);
or U901 (N_901,In_776,In_75);
xnor U902 (N_902,In_532,In_155);
xor U903 (N_903,In_342,In_927);
nand U904 (N_904,In_337,In_282);
xor U905 (N_905,In_639,In_693);
and U906 (N_906,In_83,In_829);
nor U907 (N_907,In_195,In_395);
nor U908 (N_908,In_149,In_788);
nor U909 (N_909,In_716,In_305);
xor U910 (N_910,In_887,In_952);
or U911 (N_911,In_544,In_473);
and U912 (N_912,In_522,In_764);
nor U913 (N_913,In_637,In_216);
xor U914 (N_914,In_62,In_157);
nand U915 (N_915,In_857,In_771);
and U916 (N_916,In_874,In_627);
or U917 (N_917,In_502,In_473);
nor U918 (N_918,In_340,In_606);
or U919 (N_919,In_604,In_41);
nor U920 (N_920,In_405,In_991);
nand U921 (N_921,In_776,In_647);
or U922 (N_922,In_939,In_53);
nand U923 (N_923,In_296,In_333);
xor U924 (N_924,In_11,In_45);
or U925 (N_925,In_516,In_42);
xor U926 (N_926,In_591,In_101);
and U927 (N_927,In_261,In_164);
nand U928 (N_928,In_597,In_819);
nor U929 (N_929,In_143,In_414);
or U930 (N_930,In_964,In_687);
xor U931 (N_931,In_394,In_558);
or U932 (N_932,In_900,In_811);
nor U933 (N_933,In_644,In_603);
nand U934 (N_934,In_786,In_665);
xnor U935 (N_935,In_921,In_942);
or U936 (N_936,In_640,In_243);
or U937 (N_937,In_408,In_969);
nand U938 (N_938,In_141,In_45);
or U939 (N_939,In_102,In_410);
and U940 (N_940,In_708,In_906);
and U941 (N_941,In_901,In_787);
and U942 (N_942,In_509,In_172);
xor U943 (N_943,In_254,In_241);
xnor U944 (N_944,In_654,In_684);
and U945 (N_945,In_314,In_112);
and U946 (N_946,In_457,In_459);
or U947 (N_947,In_143,In_719);
nand U948 (N_948,In_243,In_583);
or U949 (N_949,In_675,In_160);
or U950 (N_950,In_367,In_529);
xor U951 (N_951,In_345,In_265);
nand U952 (N_952,In_572,In_183);
and U953 (N_953,In_586,In_498);
nor U954 (N_954,In_976,In_594);
nor U955 (N_955,In_577,In_667);
xor U956 (N_956,In_831,In_693);
xnor U957 (N_957,In_576,In_750);
xnor U958 (N_958,In_532,In_777);
nand U959 (N_959,In_283,In_159);
xnor U960 (N_960,In_565,In_896);
or U961 (N_961,In_158,In_157);
and U962 (N_962,In_171,In_277);
xor U963 (N_963,In_330,In_902);
or U964 (N_964,In_772,In_969);
nor U965 (N_965,In_455,In_853);
nor U966 (N_966,In_14,In_479);
nand U967 (N_967,In_310,In_624);
xor U968 (N_968,In_65,In_587);
nor U969 (N_969,In_249,In_603);
nor U970 (N_970,In_288,In_889);
and U971 (N_971,In_242,In_295);
and U972 (N_972,In_808,In_288);
or U973 (N_973,In_226,In_863);
and U974 (N_974,In_385,In_505);
nor U975 (N_975,In_730,In_476);
nor U976 (N_976,In_366,In_74);
or U977 (N_977,In_456,In_414);
nor U978 (N_978,In_554,In_841);
nand U979 (N_979,In_156,In_668);
and U980 (N_980,In_882,In_706);
or U981 (N_981,In_792,In_275);
nor U982 (N_982,In_883,In_523);
nor U983 (N_983,In_830,In_843);
xnor U984 (N_984,In_572,In_52);
xnor U985 (N_985,In_523,In_861);
nor U986 (N_986,In_994,In_667);
nor U987 (N_987,In_274,In_127);
nand U988 (N_988,In_439,In_682);
and U989 (N_989,In_74,In_440);
and U990 (N_990,In_25,In_433);
xnor U991 (N_991,In_455,In_867);
nor U992 (N_992,In_342,In_855);
nand U993 (N_993,In_328,In_364);
nand U994 (N_994,In_35,In_918);
xnor U995 (N_995,In_610,In_742);
or U996 (N_996,In_627,In_280);
and U997 (N_997,In_860,In_818);
and U998 (N_998,In_722,In_34);
or U999 (N_999,In_362,In_461);
nand U1000 (N_1000,In_606,In_331);
nor U1001 (N_1001,In_167,In_338);
nor U1002 (N_1002,In_688,In_10);
xor U1003 (N_1003,In_539,In_348);
and U1004 (N_1004,In_854,In_59);
xnor U1005 (N_1005,In_122,In_435);
nand U1006 (N_1006,In_751,In_774);
and U1007 (N_1007,In_246,In_670);
and U1008 (N_1008,In_573,In_979);
xnor U1009 (N_1009,In_809,In_953);
and U1010 (N_1010,In_631,In_491);
nor U1011 (N_1011,In_273,In_706);
and U1012 (N_1012,In_830,In_504);
nor U1013 (N_1013,In_814,In_183);
nor U1014 (N_1014,In_666,In_753);
and U1015 (N_1015,In_795,In_756);
nor U1016 (N_1016,In_63,In_688);
or U1017 (N_1017,In_934,In_22);
and U1018 (N_1018,In_249,In_66);
and U1019 (N_1019,In_673,In_477);
xnor U1020 (N_1020,In_414,In_967);
or U1021 (N_1021,In_55,In_824);
and U1022 (N_1022,In_972,In_200);
and U1023 (N_1023,In_200,In_891);
nor U1024 (N_1024,In_608,In_853);
xnor U1025 (N_1025,In_566,In_269);
or U1026 (N_1026,In_48,In_698);
nor U1027 (N_1027,In_382,In_112);
or U1028 (N_1028,In_819,In_617);
and U1029 (N_1029,In_720,In_75);
and U1030 (N_1030,In_371,In_276);
nand U1031 (N_1031,In_400,In_805);
and U1032 (N_1032,In_437,In_713);
or U1033 (N_1033,In_810,In_122);
nor U1034 (N_1034,In_524,In_410);
nand U1035 (N_1035,In_725,In_317);
nand U1036 (N_1036,In_339,In_86);
xor U1037 (N_1037,In_903,In_939);
or U1038 (N_1038,In_416,In_141);
nand U1039 (N_1039,In_454,In_358);
nor U1040 (N_1040,In_413,In_722);
or U1041 (N_1041,In_154,In_330);
xnor U1042 (N_1042,In_855,In_719);
and U1043 (N_1043,In_459,In_815);
xnor U1044 (N_1044,In_706,In_929);
or U1045 (N_1045,In_715,In_909);
nand U1046 (N_1046,In_796,In_556);
nor U1047 (N_1047,In_608,In_406);
xnor U1048 (N_1048,In_826,In_434);
or U1049 (N_1049,In_332,In_904);
xnor U1050 (N_1050,In_634,In_874);
nand U1051 (N_1051,In_56,In_635);
nand U1052 (N_1052,In_24,In_40);
nand U1053 (N_1053,In_252,In_216);
or U1054 (N_1054,In_613,In_850);
or U1055 (N_1055,In_36,In_246);
xor U1056 (N_1056,In_24,In_633);
nand U1057 (N_1057,In_162,In_183);
or U1058 (N_1058,In_296,In_937);
xnor U1059 (N_1059,In_883,In_162);
nand U1060 (N_1060,In_416,In_921);
nand U1061 (N_1061,In_84,In_42);
and U1062 (N_1062,In_949,In_902);
xnor U1063 (N_1063,In_400,In_386);
or U1064 (N_1064,In_450,In_822);
xor U1065 (N_1065,In_284,In_402);
nor U1066 (N_1066,In_748,In_626);
and U1067 (N_1067,In_211,In_160);
nor U1068 (N_1068,In_224,In_474);
xnor U1069 (N_1069,In_754,In_857);
or U1070 (N_1070,In_720,In_844);
nor U1071 (N_1071,In_337,In_617);
nand U1072 (N_1072,In_196,In_574);
xor U1073 (N_1073,In_122,In_550);
and U1074 (N_1074,In_597,In_481);
nor U1075 (N_1075,In_768,In_24);
or U1076 (N_1076,In_92,In_29);
nor U1077 (N_1077,In_585,In_506);
xor U1078 (N_1078,In_764,In_828);
nor U1079 (N_1079,In_867,In_292);
or U1080 (N_1080,In_79,In_505);
nand U1081 (N_1081,In_8,In_127);
xor U1082 (N_1082,In_861,In_138);
and U1083 (N_1083,In_850,In_739);
or U1084 (N_1084,In_232,In_793);
nor U1085 (N_1085,In_108,In_266);
and U1086 (N_1086,In_599,In_876);
or U1087 (N_1087,In_443,In_587);
or U1088 (N_1088,In_763,In_12);
xnor U1089 (N_1089,In_795,In_912);
and U1090 (N_1090,In_660,In_44);
nand U1091 (N_1091,In_857,In_872);
nand U1092 (N_1092,In_786,In_559);
nand U1093 (N_1093,In_75,In_429);
nor U1094 (N_1094,In_830,In_995);
nor U1095 (N_1095,In_815,In_451);
xor U1096 (N_1096,In_202,In_206);
nand U1097 (N_1097,In_367,In_120);
nor U1098 (N_1098,In_973,In_375);
or U1099 (N_1099,In_178,In_15);
or U1100 (N_1100,In_61,In_252);
and U1101 (N_1101,In_435,In_605);
or U1102 (N_1102,In_279,In_841);
nand U1103 (N_1103,In_885,In_114);
nand U1104 (N_1104,In_922,In_83);
nand U1105 (N_1105,In_920,In_321);
nand U1106 (N_1106,In_510,In_983);
nor U1107 (N_1107,In_519,In_755);
or U1108 (N_1108,In_497,In_361);
and U1109 (N_1109,In_392,In_625);
xnor U1110 (N_1110,In_851,In_859);
and U1111 (N_1111,In_713,In_897);
and U1112 (N_1112,In_417,In_115);
nand U1113 (N_1113,In_943,In_8);
nor U1114 (N_1114,In_257,In_554);
and U1115 (N_1115,In_572,In_307);
xor U1116 (N_1116,In_416,In_968);
and U1117 (N_1117,In_815,In_67);
and U1118 (N_1118,In_860,In_762);
nand U1119 (N_1119,In_697,In_719);
or U1120 (N_1120,In_497,In_215);
and U1121 (N_1121,In_0,In_595);
xor U1122 (N_1122,In_813,In_409);
nor U1123 (N_1123,In_885,In_577);
or U1124 (N_1124,In_975,In_230);
nor U1125 (N_1125,In_196,In_375);
and U1126 (N_1126,In_486,In_497);
and U1127 (N_1127,In_130,In_383);
and U1128 (N_1128,In_376,In_288);
or U1129 (N_1129,In_113,In_532);
xnor U1130 (N_1130,In_176,In_90);
nor U1131 (N_1131,In_239,In_477);
xnor U1132 (N_1132,In_158,In_949);
nand U1133 (N_1133,In_843,In_784);
or U1134 (N_1134,In_674,In_918);
nand U1135 (N_1135,In_936,In_181);
xor U1136 (N_1136,In_881,In_256);
nor U1137 (N_1137,In_973,In_189);
xor U1138 (N_1138,In_557,In_891);
nand U1139 (N_1139,In_912,In_109);
xor U1140 (N_1140,In_671,In_176);
xnor U1141 (N_1141,In_473,In_156);
nor U1142 (N_1142,In_982,In_669);
and U1143 (N_1143,In_820,In_238);
nand U1144 (N_1144,In_319,In_630);
nand U1145 (N_1145,In_458,In_632);
and U1146 (N_1146,In_829,In_518);
nor U1147 (N_1147,In_491,In_579);
xnor U1148 (N_1148,In_907,In_185);
and U1149 (N_1149,In_288,In_873);
xnor U1150 (N_1150,In_237,In_857);
xor U1151 (N_1151,In_718,In_212);
nor U1152 (N_1152,In_449,In_21);
and U1153 (N_1153,In_656,In_591);
nand U1154 (N_1154,In_76,In_175);
or U1155 (N_1155,In_58,In_900);
nand U1156 (N_1156,In_337,In_526);
or U1157 (N_1157,In_901,In_552);
nand U1158 (N_1158,In_191,In_68);
nand U1159 (N_1159,In_601,In_527);
and U1160 (N_1160,In_206,In_713);
xnor U1161 (N_1161,In_611,In_494);
nor U1162 (N_1162,In_645,In_423);
nand U1163 (N_1163,In_902,In_333);
xnor U1164 (N_1164,In_500,In_897);
nand U1165 (N_1165,In_442,In_997);
nor U1166 (N_1166,In_929,In_761);
nor U1167 (N_1167,In_400,In_827);
or U1168 (N_1168,In_355,In_992);
or U1169 (N_1169,In_870,In_448);
xnor U1170 (N_1170,In_541,In_983);
or U1171 (N_1171,In_496,In_101);
or U1172 (N_1172,In_474,In_166);
and U1173 (N_1173,In_987,In_158);
or U1174 (N_1174,In_621,In_184);
and U1175 (N_1175,In_574,In_628);
or U1176 (N_1176,In_120,In_444);
and U1177 (N_1177,In_588,In_504);
xnor U1178 (N_1178,In_682,In_860);
nor U1179 (N_1179,In_484,In_430);
xnor U1180 (N_1180,In_545,In_392);
xor U1181 (N_1181,In_187,In_742);
nor U1182 (N_1182,In_250,In_924);
or U1183 (N_1183,In_549,In_154);
or U1184 (N_1184,In_475,In_82);
nand U1185 (N_1185,In_629,In_79);
nand U1186 (N_1186,In_180,In_649);
and U1187 (N_1187,In_832,In_93);
nand U1188 (N_1188,In_487,In_877);
or U1189 (N_1189,In_902,In_511);
xor U1190 (N_1190,In_877,In_682);
nor U1191 (N_1191,In_299,In_233);
and U1192 (N_1192,In_62,In_389);
and U1193 (N_1193,In_602,In_838);
xnor U1194 (N_1194,In_488,In_808);
or U1195 (N_1195,In_127,In_824);
xor U1196 (N_1196,In_22,In_219);
and U1197 (N_1197,In_231,In_520);
or U1198 (N_1198,In_835,In_947);
or U1199 (N_1199,In_312,In_518);
and U1200 (N_1200,In_363,In_647);
xnor U1201 (N_1201,In_177,In_714);
or U1202 (N_1202,In_894,In_735);
nor U1203 (N_1203,In_832,In_209);
nand U1204 (N_1204,In_519,In_910);
or U1205 (N_1205,In_173,In_989);
nand U1206 (N_1206,In_907,In_324);
or U1207 (N_1207,In_816,In_910);
nand U1208 (N_1208,In_283,In_417);
and U1209 (N_1209,In_380,In_50);
xnor U1210 (N_1210,In_661,In_601);
and U1211 (N_1211,In_261,In_369);
nand U1212 (N_1212,In_802,In_900);
and U1213 (N_1213,In_631,In_172);
nand U1214 (N_1214,In_616,In_648);
xor U1215 (N_1215,In_174,In_157);
xnor U1216 (N_1216,In_143,In_356);
and U1217 (N_1217,In_997,In_490);
xor U1218 (N_1218,In_72,In_960);
and U1219 (N_1219,In_186,In_936);
or U1220 (N_1220,In_696,In_944);
and U1221 (N_1221,In_711,In_632);
nor U1222 (N_1222,In_791,In_471);
and U1223 (N_1223,In_565,In_345);
or U1224 (N_1224,In_399,In_688);
xor U1225 (N_1225,In_981,In_820);
and U1226 (N_1226,In_981,In_113);
nand U1227 (N_1227,In_138,In_199);
xnor U1228 (N_1228,In_450,In_711);
nand U1229 (N_1229,In_837,In_367);
nor U1230 (N_1230,In_34,In_246);
xor U1231 (N_1231,In_844,In_220);
and U1232 (N_1232,In_32,In_38);
or U1233 (N_1233,In_815,In_736);
xnor U1234 (N_1234,In_850,In_88);
nand U1235 (N_1235,In_397,In_777);
nand U1236 (N_1236,In_244,In_739);
nand U1237 (N_1237,In_172,In_785);
nor U1238 (N_1238,In_856,In_980);
nor U1239 (N_1239,In_107,In_274);
xnor U1240 (N_1240,In_750,In_727);
xnor U1241 (N_1241,In_154,In_759);
and U1242 (N_1242,In_85,In_960);
or U1243 (N_1243,In_677,In_209);
xnor U1244 (N_1244,In_89,In_404);
and U1245 (N_1245,In_228,In_896);
or U1246 (N_1246,In_751,In_859);
nand U1247 (N_1247,In_441,In_440);
or U1248 (N_1248,In_369,In_731);
xor U1249 (N_1249,In_403,In_688);
nand U1250 (N_1250,In_162,In_966);
nand U1251 (N_1251,In_532,In_536);
xor U1252 (N_1252,In_96,In_211);
nor U1253 (N_1253,In_223,In_136);
nor U1254 (N_1254,In_69,In_161);
nand U1255 (N_1255,In_728,In_504);
xor U1256 (N_1256,In_486,In_109);
nor U1257 (N_1257,In_306,In_238);
and U1258 (N_1258,In_886,In_589);
or U1259 (N_1259,In_886,In_440);
or U1260 (N_1260,In_773,In_80);
nand U1261 (N_1261,In_220,In_540);
xnor U1262 (N_1262,In_904,In_123);
nor U1263 (N_1263,In_758,In_139);
xor U1264 (N_1264,In_486,In_654);
xnor U1265 (N_1265,In_901,In_129);
xnor U1266 (N_1266,In_249,In_278);
nor U1267 (N_1267,In_196,In_572);
xnor U1268 (N_1268,In_80,In_755);
nand U1269 (N_1269,In_354,In_622);
xnor U1270 (N_1270,In_572,In_442);
xnor U1271 (N_1271,In_368,In_319);
or U1272 (N_1272,In_856,In_283);
and U1273 (N_1273,In_808,In_292);
and U1274 (N_1274,In_403,In_354);
nor U1275 (N_1275,In_916,In_815);
or U1276 (N_1276,In_833,In_17);
xnor U1277 (N_1277,In_791,In_929);
nor U1278 (N_1278,In_609,In_264);
nand U1279 (N_1279,In_901,In_578);
and U1280 (N_1280,In_353,In_191);
nand U1281 (N_1281,In_795,In_33);
and U1282 (N_1282,In_703,In_467);
and U1283 (N_1283,In_107,In_468);
or U1284 (N_1284,In_712,In_640);
nand U1285 (N_1285,In_201,In_555);
nand U1286 (N_1286,In_856,In_216);
nand U1287 (N_1287,In_83,In_137);
nor U1288 (N_1288,In_970,In_427);
nand U1289 (N_1289,In_397,In_810);
nor U1290 (N_1290,In_775,In_920);
and U1291 (N_1291,In_89,In_640);
or U1292 (N_1292,In_630,In_297);
or U1293 (N_1293,In_728,In_446);
xnor U1294 (N_1294,In_352,In_655);
nand U1295 (N_1295,In_64,In_780);
nor U1296 (N_1296,In_764,In_592);
and U1297 (N_1297,In_702,In_245);
or U1298 (N_1298,In_279,In_979);
and U1299 (N_1299,In_66,In_875);
nand U1300 (N_1300,In_758,In_836);
nand U1301 (N_1301,In_160,In_828);
and U1302 (N_1302,In_811,In_298);
xnor U1303 (N_1303,In_695,In_201);
nor U1304 (N_1304,In_277,In_563);
xor U1305 (N_1305,In_594,In_193);
or U1306 (N_1306,In_750,In_0);
nand U1307 (N_1307,In_162,In_364);
and U1308 (N_1308,In_936,In_590);
xor U1309 (N_1309,In_415,In_986);
xor U1310 (N_1310,In_625,In_477);
and U1311 (N_1311,In_704,In_766);
nor U1312 (N_1312,In_307,In_361);
and U1313 (N_1313,In_341,In_730);
and U1314 (N_1314,In_722,In_692);
nand U1315 (N_1315,In_489,In_246);
or U1316 (N_1316,In_415,In_121);
xnor U1317 (N_1317,In_111,In_93);
nand U1318 (N_1318,In_929,In_744);
xor U1319 (N_1319,In_362,In_132);
xnor U1320 (N_1320,In_557,In_878);
and U1321 (N_1321,In_347,In_847);
xnor U1322 (N_1322,In_940,In_730);
nor U1323 (N_1323,In_234,In_203);
or U1324 (N_1324,In_198,In_140);
or U1325 (N_1325,In_170,In_917);
nor U1326 (N_1326,In_783,In_178);
and U1327 (N_1327,In_851,In_953);
nor U1328 (N_1328,In_212,In_520);
and U1329 (N_1329,In_849,In_256);
nand U1330 (N_1330,In_757,In_571);
nor U1331 (N_1331,In_838,In_909);
or U1332 (N_1332,In_654,In_476);
or U1333 (N_1333,In_664,In_181);
and U1334 (N_1334,In_688,In_267);
and U1335 (N_1335,In_708,In_542);
nand U1336 (N_1336,In_447,In_500);
xnor U1337 (N_1337,In_411,In_546);
xnor U1338 (N_1338,In_346,In_549);
and U1339 (N_1339,In_6,In_894);
nor U1340 (N_1340,In_720,In_786);
nor U1341 (N_1341,In_801,In_838);
nor U1342 (N_1342,In_483,In_12);
and U1343 (N_1343,In_445,In_89);
or U1344 (N_1344,In_603,In_136);
and U1345 (N_1345,In_303,In_627);
or U1346 (N_1346,In_427,In_601);
nor U1347 (N_1347,In_214,In_199);
nor U1348 (N_1348,In_642,In_176);
or U1349 (N_1349,In_833,In_988);
nor U1350 (N_1350,In_425,In_296);
or U1351 (N_1351,In_721,In_985);
nor U1352 (N_1352,In_531,In_647);
and U1353 (N_1353,In_284,In_522);
or U1354 (N_1354,In_553,In_206);
and U1355 (N_1355,In_208,In_73);
nand U1356 (N_1356,In_552,In_541);
nand U1357 (N_1357,In_940,In_560);
nor U1358 (N_1358,In_178,In_721);
xnor U1359 (N_1359,In_192,In_469);
nor U1360 (N_1360,In_220,In_688);
xnor U1361 (N_1361,In_112,In_788);
xnor U1362 (N_1362,In_440,In_189);
xor U1363 (N_1363,In_526,In_581);
nand U1364 (N_1364,In_393,In_341);
xnor U1365 (N_1365,In_94,In_930);
nand U1366 (N_1366,In_471,In_195);
nand U1367 (N_1367,In_714,In_291);
nor U1368 (N_1368,In_355,In_147);
or U1369 (N_1369,In_505,In_313);
or U1370 (N_1370,In_163,In_691);
or U1371 (N_1371,In_696,In_669);
nand U1372 (N_1372,In_776,In_798);
xnor U1373 (N_1373,In_644,In_480);
or U1374 (N_1374,In_566,In_829);
nand U1375 (N_1375,In_973,In_632);
and U1376 (N_1376,In_138,In_845);
and U1377 (N_1377,In_159,In_253);
nand U1378 (N_1378,In_325,In_553);
and U1379 (N_1379,In_78,In_839);
nand U1380 (N_1380,In_585,In_894);
and U1381 (N_1381,In_986,In_436);
nor U1382 (N_1382,In_523,In_373);
or U1383 (N_1383,In_25,In_585);
xor U1384 (N_1384,In_850,In_907);
and U1385 (N_1385,In_392,In_820);
nand U1386 (N_1386,In_221,In_996);
xnor U1387 (N_1387,In_68,In_183);
or U1388 (N_1388,In_108,In_155);
nand U1389 (N_1389,In_999,In_375);
or U1390 (N_1390,In_216,In_682);
nor U1391 (N_1391,In_304,In_82);
nor U1392 (N_1392,In_644,In_213);
nor U1393 (N_1393,In_719,In_422);
and U1394 (N_1394,In_176,In_369);
or U1395 (N_1395,In_666,In_98);
or U1396 (N_1396,In_274,In_718);
nor U1397 (N_1397,In_104,In_896);
or U1398 (N_1398,In_216,In_718);
and U1399 (N_1399,In_286,In_423);
or U1400 (N_1400,In_377,In_342);
and U1401 (N_1401,In_801,In_701);
xor U1402 (N_1402,In_330,In_803);
xnor U1403 (N_1403,In_195,In_886);
and U1404 (N_1404,In_791,In_100);
nor U1405 (N_1405,In_626,In_346);
nor U1406 (N_1406,In_217,In_469);
and U1407 (N_1407,In_283,In_199);
nand U1408 (N_1408,In_297,In_836);
and U1409 (N_1409,In_871,In_168);
xor U1410 (N_1410,In_61,In_282);
nand U1411 (N_1411,In_27,In_388);
and U1412 (N_1412,In_731,In_379);
nor U1413 (N_1413,In_923,In_728);
nand U1414 (N_1414,In_513,In_985);
xor U1415 (N_1415,In_336,In_755);
and U1416 (N_1416,In_899,In_309);
and U1417 (N_1417,In_358,In_665);
nor U1418 (N_1418,In_711,In_833);
nor U1419 (N_1419,In_144,In_150);
or U1420 (N_1420,In_485,In_146);
nor U1421 (N_1421,In_653,In_209);
nor U1422 (N_1422,In_3,In_160);
or U1423 (N_1423,In_441,In_249);
or U1424 (N_1424,In_493,In_366);
nand U1425 (N_1425,In_101,In_481);
nand U1426 (N_1426,In_250,In_475);
xnor U1427 (N_1427,In_161,In_798);
nor U1428 (N_1428,In_919,In_409);
nor U1429 (N_1429,In_70,In_222);
nor U1430 (N_1430,In_537,In_455);
or U1431 (N_1431,In_201,In_954);
xor U1432 (N_1432,In_2,In_826);
and U1433 (N_1433,In_225,In_772);
or U1434 (N_1434,In_666,In_533);
nand U1435 (N_1435,In_821,In_793);
or U1436 (N_1436,In_810,In_380);
nand U1437 (N_1437,In_219,In_11);
and U1438 (N_1438,In_802,In_753);
and U1439 (N_1439,In_328,In_253);
nor U1440 (N_1440,In_12,In_400);
or U1441 (N_1441,In_891,In_750);
xor U1442 (N_1442,In_200,In_77);
or U1443 (N_1443,In_36,In_417);
and U1444 (N_1444,In_442,In_827);
nor U1445 (N_1445,In_463,In_495);
nand U1446 (N_1446,In_770,In_286);
or U1447 (N_1447,In_470,In_375);
and U1448 (N_1448,In_846,In_274);
and U1449 (N_1449,In_408,In_627);
and U1450 (N_1450,In_18,In_631);
xnor U1451 (N_1451,In_83,In_782);
and U1452 (N_1452,In_195,In_524);
nor U1453 (N_1453,In_353,In_815);
nand U1454 (N_1454,In_411,In_55);
or U1455 (N_1455,In_949,In_845);
xnor U1456 (N_1456,In_428,In_421);
or U1457 (N_1457,In_297,In_283);
and U1458 (N_1458,In_994,In_879);
xnor U1459 (N_1459,In_820,In_949);
and U1460 (N_1460,In_758,In_542);
or U1461 (N_1461,In_862,In_579);
or U1462 (N_1462,In_182,In_340);
and U1463 (N_1463,In_64,In_741);
and U1464 (N_1464,In_482,In_838);
xor U1465 (N_1465,In_202,In_715);
xnor U1466 (N_1466,In_158,In_995);
xnor U1467 (N_1467,In_391,In_584);
or U1468 (N_1468,In_226,In_933);
nand U1469 (N_1469,In_199,In_738);
nor U1470 (N_1470,In_65,In_664);
xor U1471 (N_1471,In_461,In_14);
nand U1472 (N_1472,In_615,In_888);
nand U1473 (N_1473,In_416,In_326);
and U1474 (N_1474,In_866,In_744);
nor U1475 (N_1475,In_277,In_719);
and U1476 (N_1476,In_192,In_726);
or U1477 (N_1477,In_765,In_646);
and U1478 (N_1478,In_376,In_367);
and U1479 (N_1479,In_786,In_597);
or U1480 (N_1480,In_634,In_602);
xnor U1481 (N_1481,In_880,In_20);
nor U1482 (N_1482,In_381,In_237);
nor U1483 (N_1483,In_909,In_881);
or U1484 (N_1484,In_157,In_536);
xor U1485 (N_1485,In_818,In_707);
xor U1486 (N_1486,In_233,In_878);
or U1487 (N_1487,In_704,In_896);
nand U1488 (N_1488,In_851,In_79);
and U1489 (N_1489,In_491,In_954);
xnor U1490 (N_1490,In_64,In_235);
nand U1491 (N_1491,In_721,In_185);
xor U1492 (N_1492,In_1,In_42);
and U1493 (N_1493,In_17,In_763);
or U1494 (N_1494,In_547,In_365);
and U1495 (N_1495,In_264,In_409);
xor U1496 (N_1496,In_113,In_813);
nand U1497 (N_1497,In_637,In_541);
nand U1498 (N_1498,In_549,In_40);
and U1499 (N_1499,In_984,In_381);
nand U1500 (N_1500,In_834,In_143);
xnor U1501 (N_1501,In_349,In_865);
and U1502 (N_1502,In_133,In_538);
xnor U1503 (N_1503,In_209,In_123);
and U1504 (N_1504,In_220,In_404);
or U1505 (N_1505,In_789,In_242);
and U1506 (N_1506,In_642,In_503);
or U1507 (N_1507,In_222,In_834);
nand U1508 (N_1508,In_728,In_370);
xor U1509 (N_1509,In_67,In_994);
and U1510 (N_1510,In_474,In_483);
nand U1511 (N_1511,In_373,In_634);
or U1512 (N_1512,In_488,In_380);
nand U1513 (N_1513,In_491,In_176);
or U1514 (N_1514,In_451,In_33);
and U1515 (N_1515,In_406,In_288);
nor U1516 (N_1516,In_827,In_267);
nor U1517 (N_1517,In_559,In_451);
xnor U1518 (N_1518,In_84,In_571);
xnor U1519 (N_1519,In_959,In_91);
or U1520 (N_1520,In_144,In_208);
and U1521 (N_1521,In_412,In_876);
xnor U1522 (N_1522,In_270,In_252);
nor U1523 (N_1523,In_252,In_930);
and U1524 (N_1524,In_522,In_722);
xnor U1525 (N_1525,In_422,In_96);
xor U1526 (N_1526,In_512,In_641);
nor U1527 (N_1527,In_692,In_79);
xor U1528 (N_1528,In_623,In_353);
xnor U1529 (N_1529,In_892,In_960);
and U1530 (N_1530,In_73,In_395);
and U1531 (N_1531,In_121,In_385);
xnor U1532 (N_1532,In_992,In_966);
and U1533 (N_1533,In_772,In_546);
and U1534 (N_1534,In_686,In_72);
and U1535 (N_1535,In_796,In_902);
or U1536 (N_1536,In_3,In_171);
xor U1537 (N_1537,In_158,In_289);
nand U1538 (N_1538,In_944,In_609);
or U1539 (N_1539,In_378,In_537);
nand U1540 (N_1540,In_61,In_523);
or U1541 (N_1541,In_136,In_702);
and U1542 (N_1542,In_342,In_243);
and U1543 (N_1543,In_809,In_992);
xnor U1544 (N_1544,In_610,In_87);
nand U1545 (N_1545,In_635,In_41);
and U1546 (N_1546,In_525,In_20);
or U1547 (N_1547,In_926,In_991);
and U1548 (N_1548,In_715,In_61);
and U1549 (N_1549,In_938,In_257);
or U1550 (N_1550,In_18,In_736);
xnor U1551 (N_1551,In_763,In_73);
xor U1552 (N_1552,In_726,In_635);
and U1553 (N_1553,In_356,In_711);
nor U1554 (N_1554,In_565,In_48);
xnor U1555 (N_1555,In_904,In_592);
and U1556 (N_1556,In_870,In_230);
xnor U1557 (N_1557,In_874,In_818);
and U1558 (N_1558,In_183,In_472);
and U1559 (N_1559,In_602,In_796);
nand U1560 (N_1560,In_561,In_949);
nand U1561 (N_1561,In_825,In_987);
nor U1562 (N_1562,In_8,In_746);
nor U1563 (N_1563,In_808,In_644);
nand U1564 (N_1564,In_566,In_754);
xnor U1565 (N_1565,In_609,In_533);
nand U1566 (N_1566,In_311,In_792);
nand U1567 (N_1567,In_736,In_199);
nand U1568 (N_1568,In_943,In_567);
and U1569 (N_1569,In_444,In_37);
nand U1570 (N_1570,In_697,In_807);
xnor U1571 (N_1571,In_495,In_41);
and U1572 (N_1572,In_205,In_263);
and U1573 (N_1573,In_969,In_982);
or U1574 (N_1574,In_752,In_799);
xor U1575 (N_1575,In_957,In_991);
nor U1576 (N_1576,In_416,In_586);
and U1577 (N_1577,In_549,In_539);
nor U1578 (N_1578,In_884,In_820);
xor U1579 (N_1579,In_964,In_610);
and U1580 (N_1580,In_797,In_446);
nor U1581 (N_1581,In_933,In_572);
and U1582 (N_1582,In_50,In_973);
and U1583 (N_1583,In_102,In_573);
or U1584 (N_1584,In_673,In_272);
or U1585 (N_1585,In_340,In_939);
xnor U1586 (N_1586,In_716,In_819);
nand U1587 (N_1587,In_22,In_223);
or U1588 (N_1588,In_741,In_693);
and U1589 (N_1589,In_646,In_400);
nor U1590 (N_1590,In_629,In_633);
or U1591 (N_1591,In_239,In_159);
xor U1592 (N_1592,In_572,In_339);
or U1593 (N_1593,In_960,In_164);
nand U1594 (N_1594,In_65,In_889);
or U1595 (N_1595,In_662,In_203);
nand U1596 (N_1596,In_367,In_626);
and U1597 (N_1597,In_534,In_161);
or U1598 (N_1598,In_147,In_332);
and U1599 (N_1599,In_899,In_263);
nor U1600 (N_1600,In_974,In_909);
nand U1601 (N_1601,In_589,In_618);
xnor U1602 (N_1602,In_15,In_690);
nor U1603 (N_1603,In_615,In_385);
nor U1604 (N_1604,In_641,In_562);
xor U1605 (N_1605,In_507,In_513);
xor U1606 (N_1606,In_418,In_423);
nand U1607 (N_1607,In_937,In_120);
xnor U1608 (N_1608,In_623,In_521);
xor U1609 (N_1609,In_806,In_314);
or U1610 (N_1610,In_279,In_107);
or U1611 (N_1611,In_716,In_853);
nand U1612 (N_1612,In_961,In_548);
nand U1613 (N_1613,In_634,In_72);
and U1614 (N_1614,In_745,In_947);
or U1615 (N_1615,In_512,In_733);
nor U1616 (N_1616,In_99,In_852);
or U1617 (N_1617,In_740,In_951);
nand U1618 (N_1618,In_865,In_532);
nor U1619 (N_1619,In_225,In_995);
or U1620 (N_1620,In_977,In_228);
nand U1621 (N_1621,In_108,In_562);
and U1622 (N_1622,In_749,In_414);
xnor U1623 (N_1623,In_886,In_532);
or U1624 (N_1624,In_493,In_253);
nand U1625 (N_1625,In_330,In_479);
or U1626 (N_1626,In_931,In_304);
xnor U1627 (N_1627,In_590,In_433);
nand U1628 (N_1628,In_911,In_813);
and U1629 (N_1629,In_572,In_684);
xnor U1630 (N_1630,In_272,In_311);
and U1631 (N_1631,In_84,In_990);
or U1632 (N_1632,In_764,In_798);
xnor U1633 (N_1633,In_765,In_51);
or U1634 (N_1634,In_455,In_670);
nand U1635 (N_1635,In_455,In_595);
xor U1636 (N_1636,In_964,In_852);
nand U1637 (N_1637,In_454,In_625);
xnor U1638 (N_1638,In_390,In_511);
xnor U1639 (N_1639,In_341,In_685);
xnor U1640 (N_1640,In_117,In_738);
nand U1641 (N_1641,In_775,In_24);
xnor U1642 (N_1642,In_287,In_554);
nand U1643 (N_1643,In_599,In_696);
or U1644 (N_1644,In_56,In_160);
nand U1645 (N_1645,In_234,In_919);
xor U1646 (N_1646,In_594,In_522);
or U1647 (N_1647,In_802,In_55);
or U1648 (N_1648,In_843,In_89);
nor U1649 (N_1649,In_52,In_165);
and U1650 (N_1650,In_706,In_277);
nand U1651 (N_1651,In_393,In_305);
nand U1652 (N_1652,In_326,In_940);
nand U1653 (N_1653,In_520,In_970);
and U1654 (N_1654,In_461,In_373);
nor U1655 (N_1655,In_675,In_906);
and U1656 (N_1656,In_85,In_113);
or U1657 (N_1657,In_479,In_47);
nand U1658 (N_1658,In_329,In_187);
nor U1659 (N_1659,In_877,In_996);
and U1660 (N_1660,In_822,In_861);
or U1661 (N_1661,In_916,In_582);
or U1662 (N_1662,In_868,In_418);
nand U1663 (N_1663,In_207,In_891);
or U1664 (N_1664,In_558,In_881);
or U1665 (N_1665,In_845,In_324);
and U1666 (N_1666,In_66,In_204);
xnor U1667 (N_1667,In_741,In_543);
nand U1668 (N_1668,In_1,In_373);
or U1669 (N_1669,In_425,In_48);
nor U1670 (N_1670,In_871,In_220);
nor U1671 (N_1671,In_938,In_497);
or U1672 (N_1672,In_742,In_521);
nand U1673 (N_1673,In_444,In_334);
xor U1674 (N_1674,In_860,In_616);
nor U1675 (N_1675,In_353,In_46);
and U1676 (N_1676,In_921,In_998);
or U1677 (N_1677,In_881,In_375);
and U1678 (N_1678,In_315,In_936);
or U1679 (N_1679,In_956,In_696);
xnor U1680 (N_1680,In_6,In_850);
nand U1681 (N_1681,In_546,In_803);
and U1682 (N_1682,In_152,In_503);
or U1683 (N_1683,In_144,In_854);
nand U1684 (N_1684,In_695,In_696);
nand U1685 (N_1685,In_4,In_426);
nor U1686 (N_1686,In_580,In_753);
xnor U1687 (N_1687,In_42,In_62);
nor U1688 (N_1688,In_795,In_221);
xor U1689 (N_1689,In_405,In_989);
or U1690 (N_1690,In_860,In_689);
or U1691 (N_1691,In_576,In_923);
xor U1692 (N_1692,In_160,In_81);
or U1693 (N_1693,In_719,In_622);
or U1694 (N_1694,In_907,In_556);
and U1695 (N_1695,In_636,In_643);
or U1696 (N_1696,In_514,In_119);
and U1697 (N_1697,In_953,In_198);
nor U1698 (N_1698,In_314,In_752);
xnor U1699 (N_1699,In_599,In_382);
and U1700 (N_1700,In_215,In_945);
nor U1701 (N_1701,In_42,In_538);
nand U1702 (N_1702,In_794,In_899);
xor U1703 (N_1703,In_640,In_886);
nor U1704 (N_1704,In_393,In_982);
xnor U1705 (N_1705,In_575,In_827);
nor U1706 (N_1706,In_822,In_196);
xor U1707 (N_1707,In_109,In_567);
and U1708 (N_1708,In_38,In_597);
or U1709 (N_1709,In_173,In_667);
and U1710 (N_1710,In_571,In_865);
or U1711 (N_1711,In_100,In_729);
nor U1712 (N_1712,In_167,In_554);
xor U1713 (N_1713,In_257,In_524);
or U1714 (N_1714,In_667,In_229);
nand U1715 (N_1715,In_945,In_201);
xnor U1716 (N_1716,In_439,In_923);
xor U1717 (N_1717,In_716,In_466);
nand U1718 (N_1718,In_695,In_565);
xnor U1719 (N_1719,In_619,In_195);
or U1720 (N_1720,In_752,In_883);
xnor U1721 (N_1721,In_325,In_113);
nand U1722 (N_1722,In_126,In_887);
xor U1723 (N_1723,In_349,In_104);
nor U1724 (N_1724,In_392,In_898);
nand U1725 (N_1725,In_839,In_761);
and U1726 (N_1726,In_179,In_627);
xnor U1727 (N_1727,In_788,In_424);
xnor U1728 (N_1728,In_409,In_978);
and U1729 (N_1729,In_394,In_876);
xor U1730 (N_1730,In_493,In_492);
nor U1731 (N_1731,In_715,In_70);
xor U1732 (N_1732,In_513,In_326);
and U1733 (N_1733,In_903,In_8);
xnor U1734 (N_1734,In_575,In_184);
nor U1735 (N_1735,In_533,In_988);
or U1736 (N_1736,In_763,In_948);
nand U1737 (N_1737,In_11,In_943);
nand U1738 (N_1738,In_236,In_536);
nor U1739 (N_1739,In_647,In_970);
nand U1740 (N_1740,In_81,In_909);
nor U1741 (N_1741,In_679,In_415);
or U1742 (N_1742,In_838,In_721);
nor U1743 (N_1743,In_505,In_698);
xnor U1744 (N_1744,In_520,In_455);
nand U1745 (N_1745,In_699,In_485);
nor U1746 (N_1746,In_503,In_197);
xor U1747 (N_1747,In_565,In_463);
nor U1748 (N_1748,In_866,In_284);
nor U1749 (N_1749,In_825,In_869);
nor U1750 (N_1750,In_737,In_709);
nand U1751 (N_1751,In_887,In_302);
nor U1752 (N_1752,In_540,In_667);
or U1753 (N_1753,In_539,In_725);
nor U1754 (N_1754,In_13,In_936);
nand U1755 (N_1755,In_817,In_161);
or U1756 (N_1756,In_228,In_213);
xor U1757 (N_1757,In_137,In_68);
nand U1758 (N_1758,In_961,In_535);
nor U1759 (N_1759,In_817,In_952);
nor U1760 (N_1760,In_264,In_142);
and U1761 (N_1761,In_51,In_815);
or U1762 (N_1762,In_812,In_61);
xnor U1763 (N_1763,In_86,In_700);
or U1764 (N_1764,In_461,In_320);
nand U1765 (N_1765,In_366,In_266);
nand U1766 (N_1766,In_512,In_364);
nor U1767 (N_1767,In_51,In_160);
or U1768 (N_1768,In_163,In_214);
nand U1769 (N_1769,In_106,In_524);
or U1770 (N_1770,In_749,In_196);
xnor U1771 (N_1771,In_61,In_556);
nor U1772 (N_1772,In_969,In_416);
and U1773 (N_1773,In_499,In_331);
and U1774 (N_1774,In_178,In_537);
and U1775 (N_1775,In_137,In_596);
xor U1776 (N_1776,In_542,In_377);
and U1777 (N_1777,In_206,In_742);
and U1778 (N_1778,In_514,In_431);
nor U1779 (N_1779,In_166,In_500);
or U1780 (N_1780,In_186,In_722);
nand U1781 (N_1781,In_806,In_246);
nand U1782 (N_1782,In_436,In_816);
and U1783 (N_1783,In_201,In_609);
or U1784 (N_1784,In_323,In_197);
xnor U1785 (N_1785,In_854,In_976);
and U1786 (N_1786,In_515,In_273);
nand U1787 (N_1787,In_367,In_153);
and U1788 (N_1788,In_595,In_766);
or U1789 (N_1789,In_314,In_879);
nand U1790 (N_1790,In_175,In_65);
and U1791 (N_1791,In_715,In_351);
or U1792 (N_1792,In_412,In_850);
and U1793 (N_1793,In_325,In_563);
nand U1794 (N_1794,In_670,In_456);
nand U1795 (N_1795,In_623,In_696);
and U1796 (N_1796,In_57,In_634);
xnor U1797 (N_1797,In_639,In_785);
and U1798 (N_1798,In_890,In_670);
nor U1799 (N_1799,In_280,In_516);
nor U1800 (N_1800,In_698,In_957);
xor U1801 (N_1801,In_81,In_620);
or U1802 (N_1802,In_431,In_742);
and U1803 (N_1803,In_414,In_976);
nand U1804 (N_1804,In_203,In_892);
nor U1805 (N_1805,In_10,In_705);
xnor U1806 (N_1806,In_532,In_537);
nor U1807 (N_1807,In_116,In_489);
xnor U1808 (N_1808,In_873,In_893);
nor U1809 (N_1809,In_951,In_40);
and U1810 (N_1810,In_396,In_298);
or U1811 (N_1811,In_892,In_749);
nand U1812 (N_1812,In_737,In_39);
xor U1813 (N_1813,In_621,In_243);
and U1814 (N_1814,In_40,In_626);
xor U1815 (N_1815,In_187,In_497);
xnor U1816 (N_1816,In_760,In_201);
or U1817 (N_1817,In_195,In_256);
xor U1818 (N_1818,In_420,In_742);
nand U1819 (N_1819,In_114,In_638);
nor U1820 (N_1820,In_114,In_824);
nor U1821 (N_1821,In_910,In_233);
or U1822 (N_1822,In_273,In_135);
and U1823 (N_1823,In_489,In_981);
nor U1824 (N_1824,In_731,In_695);
or U1825 (N_1825,In_683,In_148);
and U1826 (N_1826,In_642,In_219);
xnor U1827 (N_1827,In_274,In_116);
and U1828 (N_1828,In_857,In_271);
nand U1829 (N_1829,In_967,In_785);
and U1830 (N_1830,In_153,In_410);
and U1831 (N_1831,In_886,In_305);
or U1832 (N_1832,In_915,In_773);
or U1833 (N_1833,In_968,In_959);
xor U1834 (N_1834,In_422,In_995);
nor U1835 (N_1835,In_224,In_114);
nand U1836 (N_1836,In_469,In_528);
nor U1837 (N_1837,In_573,In_902);
nor U1838 (N_1838,In_630,In_225);
nor U1839 (N_1839,In_391,In_73);
nor U1840 (N_1840,In_749,In_146);
nand U1841 (N_1841,In_90,In_673);
and U1842 (N_1842,In_569,In_959);
nand U1843 (N_1843,In_863,In_163);
and U1844 (N_1844,In_896,In_889);
or U1845 (N_1845,In_77,In_500);
nor U1846 (N_1846,In_50,In_418);
or U1847 (N_1847,In_829,In_975);
xnor U1848 (N_1848,In_764,In_647);
nor U1849 (N_1849,In_203,In_856);
nand U1850 (N_1850,In_512,In_215);
and U1851 (N_1851,In_739,In_60);
xor U1852 (N_1852,In_60,In_66);
nand U1853 (N_1853,In_884,In_79);
and U1854 (N_1854,In_455,In_285);
and U1855 (N_1855,In_481,In_662);
or U1856 (N_1856,In_886,In_454);
nand U1857 (N_1857,In_900,In_577);
xor U1858 (N_1858,In_257,In_251);
or U1859 (N_1859,In_690,In_512);
xnor U1860 (N_1860,In_328,In_871);
xor U1861 (N_1861,In_535,In_876);
xnor U1862 (N_1862,In_460,In_784);
nor U1863 (N_1863,In_724,In_647);
nor U1864 (N_1864,In_196,In_368);
and U1865 (N_1865,In_465,In_840);
nand U1866 (N_1866,In_863,In_135);
and U1867 (N_1867,In_881,In_341);
nand U1868 (N_1868,In_813,In_685);
nand U1869 (N_1869,In_105,In_303);
nor U1870 (N_1870,In_547,In_966);
and U1871 (N_1871,In_16,In_546);
nand U1872 (N_1872,In_784,In_820);
or U1873 (N_1873,In_569,In_677);
nand U1874 (N_1874,In_639,In_973);
xor U1875 (N_1875,In_212,In_111);
xor U1876 (N_1876,In_561,In_436);
or U1877 (N_1877,In_704,In_774);
and U1878 (N_1878,In_893,In_478);
nand U1879 (N_1879,In_249,In_476);
and U1880 (N_1880,In_961,In_509);
xor U1881 (N_1881,In_513,In_545);
nor U1882 (N_1882,In_917,In_345);
nand U1883 (N_1883,In_743,In_621);
xnor U1884 (N_1884,In_518,In_415);
and U1885 (N_1885,In_247,In_162);
nand U1886 (N_1886,In_370,In_491);
nand U1887 (N_1887,In_351,In_417);
nor U1888 (N_1888,In_555,In_799);
nand U1889 (N_1889,In_588,In_160);
xnor U1890 (N_1890,In_147,In_421);
xnor U1891 (N_1891,In_111,In_129);
xor U1892 (N_1892,In_713,In_329);
nand U1893 (N_1893,In_505,In_672);
nand U1894 (N_1894,In_82,In_283);
and U1895 (N_1895,In_48,In_584);
or U1896 (N_1896,In_607,In_841);
nor U1897 (N_1897,In_607,In_590);
or U1898 (N_1898,In_416,In_695);
xor U1899 (N_1899,In_983,In_539);
or U1900 (N_1900,In_626,In_756);
or U1901 (N_1901,In_240,In_529);
nor U1902 (N_1902,In_640,In_625);
nor U1903 (N_1903,In_799,In_507);
nand U1904 (N_1904,In_662,In_151);
or U1905 (N_1905,In_620,In_460);
or U1906 (N_1906,In_80,In_794);
and U1907 (N_1907,In_622,In_477);
nand U1908 (N_1908,In_715,In_731);
and U1909 (N_1909,In_984,In_553);
and U1910 (N_1910,In_527,In_958);
nand U1911 (N_1911,In_649,In_809);
xor U1912 (N_1912,In_404,In_410);
and U1913 (N_1913,In_194,In_12);
nand U1914 (N_1914,In_889,In_178);
nand U1915 (N_1915,In_66,In_941);
or U1916 (N_1916,In_117,In_606);
nor U1917 (N_1917,In_386,In_331);
or U1918 (N_1918,In_647,In_319);
or U1919 (N_1919,In_493,In_56);
and U1920 (N_1920,In_344,In_576);
nand U1921 (N_1921,In_634,In_353);
nand U1922 (N_1922,In_655,In_409);
or U1923 (N_1923,In_432,In_764);
nor U1924 (N_1924,In_181,In_282);
xnor U1925 (N_1925,In_919,In_803);
and U1926 (N_1926,In_127,In_904);
nor U1927 (N_1927,In_334,In_225);
and U1928 (N_1928,In_30,In_338);
nor U1929 (N_1929,In_407,In_508);
or U1930 (N_1930,In_347,In_749);
and U1931 (N_1931,In_497,In_291);
or U1932 (N_1932,In_806,In_415);
xnor U1933 (N_1933,In_842,In_179);
and U1934 (N_1934,In_321,In_249);
nor U1935 (N_1935,In_36,In_460);
xnor U1936 (N_1936,In_322,In_260);
nor U1937 (N_1937,In_728,In_443);
nor U1938 (N_1938,In_206,In_31);
and U1939 (N_1939,In_94,In_365);
and U1940 (N_1940,In_391,In_361);
or U1941 (N_1941,In_320,In_497);
or U1942 (N_1942,In_42,In_87);
or U1943 (N_1943,In_23,In_517);
and U1944 (N_1944,In_510,In_66);
nand U1945 (N_1945,In_408,In_787);
xnor U1946 (N_1946,In_563,In_880);
and U1947 (N_1947,In_616,In_108);
nand U1948 (N_1948,In_350,In_823);
xor U1949 (N_1949,In_117,In_770);
and U1950 (N_1950,In_447,In_231);
nor U1951 (N_1951,In_706,In_948);
nand U1952 (N_1952,In_404,In_186);
xnor U1953 (N_1953,In_14,In_250);
xor U1954 (N_1954,In_853,In_13);
nand U1955 (N_1955,In_390,In_610);
and U1956 (N_1956,In_154,In_48);
nand U1957 (N_1957,In_598,In_286);
nand U1958 (N_1958,In_116,In_724);
nand U1959 (N_1959,In_101,In_602);
or U1960 (N_1960,In_347,In_619);
and U1961 (N_1961,In_768,In_153);
xor U1962 (N_1962,In_190,In_211);
nor U1963 (N_1963,In_128,In_261);
nor U1964 (N_1964,In_945,In_105);
nand U1965 (N_1965,In_329,In_97);
or U1966 (N_1966,In_675,In_403);
nand U1967 (N_1967,In_769,In_100);
and U1968 (N_1968,In_248,In_40);
and U1969 (N_1969,In_203,In_575);
and U1970 (N_1970,In_302,In_85);
nor U1971 (N_1971,In_530,In_850);
nand U1972 (N_1972,In_763,In_326);
xor U1973 (N_1973,In_780,In_93);
nor U1974 (N_1974,In_35,In_319);
or U1975 (N_1975,In_720,In_312);
xor U1976 (N_1976,In_859,In_110);
nor U1977 (N_1977,In_34,In_498);
xnor U1978 (N_1978,In_924,In_731);
nor U1979 (N_1979,In_986,In_428);
nand U1980 (N_1980,In_458,In_85);
nor U1981 (N_1981,In_837,In_985);
or U1982 (N_1982,In_983,In_810);
or U1983 (N_1983,In_866,In_475);
nor U1984 (N_1984,In_612,In_853);
xor U1985 (N_1985,In_118,In_225);
nor U1986 (N_1986,In_885,In_162);
and U1987 (N_1987,In_858,In_658);
nor U1988 (N_1988,In_984,In_207);
or U1989 (N_1989,In_702,In_572);
or U1990 (N_1990,In_559,In_716);
nand U1991 (N_1991,In_199,In_718);
xor U1992 (N_1992,In_189,In_593);
xor U1993 (N_1993,In_649,In_319);
or U1994 (N_1994,In_152,In_429);
nand U1995 (N_1995,In_243,In_443);
nand U1996 (N_1996,In_285,In_174);
or U1997 (N_1997,In_351,In_588);
xor U1998 (N_1998,In_734,In_891);
or U1999 (N_1999,In_165,In_725);
nand U2000 (N_2000,N_868,N_416);
xnor U2001 (N_2001,N_1086,N_166);
nor U2002 (N_2002,N_1356,N_1863);
nor U2003 (N_2003,N_1481,N_184);
or U2004 (N_2004,N_226,N_1606);
xor U2005 (N_2005,N_1212,N_1243);
nand U2006 (N_2006,N_242,N_453);
nor U2007 (N_2007,N_472,N_1470);
or U2008 (N_2008,N_1079,N_1991);
and U2009 (N_2009,N_115,N_96);
nand U2010 (N_2010,N_373,N_1432);
nand U2011 (N_2011,N_488,N_255);
nand U2012 (N_2012,N_1067,N_2);
or U2013 (N_2013,N_1018,N_1281);
and U2014 (N_2014,N_1050,N_341);
nand U2015 (N_2015,N_1479,N_1228);
or U2016 (N_2016,N_414,N_1602);
and U2017 (N_2017,N_1822,N_511);
or U2018 (N_2018,N_1007,N_1534);
xnor U2019 (N_2019,N_710,N_958);
xor U2020 (N_2020,N_1156,N_429);
nor U2021 (N_2021,N_314,N_1418);
nor U2022 (N_2022,N_1807,N_1659);
nor U2023 (N_2023,N_933,N_763);
nand U2024 (N_2024,N_1823,N_970);
xor U2025 (N_2025,N_1236,N_366);
xor U2026 (N_2026,N_1248,N_1084);
and U2027 (N_2027,N_1633,N_848);
xnor U2028 (N_2028,N_1502,N_1876);
and U2029 (N_2029,N_380,N_574);
xor U2030 (N_2030,N_1810,N_239);
nand U2031 (N_2031,N_798,N_623);
nor U2032 (N_2032,N_789,N_1589);
nand U2033 (N_2033,N_509,N_1610);
nor U2034 (N_2034,N_1585,N_1398);
and U2035 (N_2035,N_864,N_1170);
or U2036 (N_2036,N_1842,N_362);
nand U2037 (N_2037,N_762,N_375);
and U2038 (N_2038,N_1200,N_1676);
and U2039 (N_2039,N_1045,N_562);
or U2040 (N_2040,N_1406,N_1819);
nand U2041 (N_2041,N_823,N_408);
and U2042 (N_2042,N_838,N_61);
or U2043 (N_2043,N_529,N_1956);
or U2044 (N_2044,N_718,N_135);
and U2045 (N_2045,N_444,N_1485);
and U2046 (N_2046,N_997,N_101);
xnor U2047 (N_2047,N_1094,N_302);
nor U2048 (N_2048,N_1010,N_1405);
nand U2049 (N_2049,N_942,N_849);
or U2050 (N_2050,N_836,N_11);
xnor U2051 (N_2051,N_133,N_833);
and U2052 (N_2052,N_171,N_690);
and U2053 (N_2053,N_622,N_458);
nand U2054 (N_2054,N_1499,N_1533);
xor U2055 (N_2055,N_413,N_1706);
or U2056 (N_2056,N_1446,N_1614);
and U2057 (N_2057,N_1239,N_411);
and U2058 (N_2058,N_437,N_555);
xor U2059 (N_2059,N_1570,N_581);
and U2060 (N_2060,N_670,N_527);
nor U2061 (N_2061,N_1208,N_1076);
nand U2062 (N_2062,N_1512,N_43);
nor U2063 (N_2063,N_1152,N_1039);
nor U2064 (N_2064,N_870,N_1783);
and U2065 (N_2065,N_1015,N_1558);
nor U2066 (N_2066,N_777,N_318);
nand U2067 (N_2067,N_455,N_1594);
nor U2068 (N_2068,N_647,N_1328);
nand U2069 (N_2069,N_493,N_273);
nand U2070 (N_2070,N_1722,N_1518);
nor U2071 (N_2071,N_1225,N_1017);
and U2072 (N_2072,N_258,N_1409);
and U2073 (N_2073,N_1312,N_1429);
nor U2074 (N_2074,N_1548,N_83);
or U2075 (N_2075,N_682,N_816);
or U2076 (N_2076,N_1455,N_1923);
nor U2077 (N_2077,N_1527,N_1615);
and U2078 (N_2078,N_1787,N_1349);
xnor U2079 (N_2079,N_1258,N_1342);
and U2080 (N_2080,N_1472,N_1983);
nor U2081 (N_2081,N_501,N_1544);
or U2082 (N_2082,N_826,N_1126);
and U2083 (N_2083,N_521,N_340);
xnor U2084 (N_2084,N_712,N_272);
and U2085 (N_2085,N_1816,N_1922);
or U2086 (N_2086,N_185,N_1346);
xor U2087 (N_2087,N_391,N_1549);
xnor U2088 (N_2088,N_1153,N_445);
xnor U2089 (N_2089,N_1068,N_1394);
and U2090 (N_2090,N_1888,N_1833);
nand U2091 (N_2091,N_580,N_671);
nand U2092 (N_2092,N_382,N_1764);
nor U2093 (N_2093,N_1901,N_680);
nand U2094 (N_2094,N_1775,N_1114);
or U2095 (N_2095,N_787,N_552);
nand U2096 (N_2096,N_1973,N_528);
and U2097 (N_2097,N_1367,N_1052);
or U2098 (N_2098,N_363,N_1663);
and U2099 (N_2099,N_1118,N_1586);
nand U2100 (N_2100,N_919,N_585);
and U2101 (N_2101,N_434,N_234);
xor U2102 (N_2102,N_74,N_518);
nand U2103 (N_2103,N_1791,N_1392);
and U2104 (N_2104,N_1858,N_791);
nand U2105 (N_2105,N_750,N_1369);
nor U2106 (N_2106,N_1428,N_1458);
nor U2107 (N_2107,N_141,N_1213);
xor U2108 (N_2108,N_945,N_407);
nor U2109 (N_2109,N_1577,N_361);
or U2110 (N_2110,N_1848,N_157);
nor U2111 (N_2111,N_1964,N_1628);
or U2112 (N_2112,N_550,N_223);
and U2113 (N_2113,N_1242,N_1830);
xor U2114 (N_2114,N_47,N_1725);
and U2115 (N_2115,N_312,N_50);
and U2116 (N_2116,N_551,N_315);
nor U2117 (N_2117,N_1305,N_485);
or U2118 (N_2118,N_1645,N_146);
or U2119 (N_2119,N_1662,N_244);
xor U2120 (N_2120,N_820,N_1436);
nor U2121 (N_2121,N_590,N_539);
and U2122 (N_2122,N_1073,N_1237);
or U2123 (N_2123,N_704,N_91);
and U2124 (N_2124,N_1908,N_65);
nor U2125 (N_2125,N_1648,N_1302);
or U2126 (N_2126,N_861,N_1203);
and U2127 (N_2127,N_1252,N_525);
and U2128 (N_2128,N_1077,N_1047);
nand U2129 (N_2129,N_1777,N_1289);
nor U2130 (N_2130,N_1561,N_1853);
nor U2131 (N_2131,N_1595,N_5);
nor U2132 (N_2132,N_3,N_1605);
nor U2133 (N_2133,N_1354,N_1188);
nand U2134 (N_2134,N_337,N_1668);
nand U2135 (N_2135,N_1573,N_9);
and U2136 (N_2136,N_784,N_1206);
xor U2137 (N_2137,N_1732,N_503);
and U2138 (N_2138,N_1849,N_1408);
and U2139 (N_2139,N_1875,N_41);
or U2140 (N_2140,N_751,N_125);
and U2141 (N_2141,N_656,N_1059);
and U2142 (N_2142,N_1509,N_1332);
nor U2143 (N_2143,N_326,N_1139);
or U2144 (N_2144,N_1234,N_1729);
nand U2145 (N_2145,N_1159,N_1207);
xnor U2146 (N_2146,N_107,N_224);
nand U2147 (N_2147,N_37,N_1905);
or U2148 (N_2148,N_1501,N_499);
nand U2149 (N_2149,N_1838,N_1507);
or U2150 (N_2150,N_1099,N_822);
and U2151 (N_2151,N_533,N_1675);
nor U2152 (N_2152,N_918,N_1657);
or U2153 (N_2153,N_876,N_1646);
nand U2154 (N_2154,N_516,N_999);
or U2155 (N_2155,N_1442,N_1269);
nand U2156 (N_2156,N_691,N_253);
and U2157 (N_2157,N_839,N_1181);
or U2158 (N_2158,N_1740,N_433);
or U2159 (N_2159,N_985,N_741);
nor U2160 (N_2160,N_351,N_87);
nand U2161 (N_2161,N_1866,N_1574);
nor U2162 (N_2162,N_1301,N_360);
and U2163 (N_2163,N_759,N_1230);
nand U2164 (N_2164,N_1075,N_967);
nor U2165 (N_2165,N_10,N_1660);
xnor U2166 (N_2166,N_1300,N_1487);
nand U2167 (N_2167,N_1226,N_924);
or U2168 (N_2168,N_1880,N_290);
or U2169 (N_2169,N_1782,N_277);
nor U2170 (N_2170,N_473,N_4);
or U2171 (N_2171,N_486,N_1705);
xnor U2172 (N_2172,N_847,N_752);
or U2173 (N_2173,N_131,N_1115);
xor U2174 (N_2174,N_556,N_769);
or U2175 (N_2175,N_944,N_1467);
xor U2176 (N_2176,N_811,N_929);
nor U2177 (N_2177,N_1388,N_218);
xnor U2178 (N_2178,N_213,N_720);
nand U2179 (N_2179,N_801,N_1380);
nor U2180 (N_2180,N_842,N_229);
nor U2181 (N_2181,N_1927,N_116);
or U2182 (N_2182,N_1308,N_1789);
and U2183 (N_2183,N_1963,N_524);
and U2184 (N_2184,N_597,N_459);
xnor U2185 (N_2185,N_1439,N_1461);
nand U2186 (N_2186,N_678,N_547);
nor U2187 (N_2187,N_236,N_237);
nand U2188 (N_2188,N_1781,N_1263);
nand U2189 (N_2189,N_292,N_320);
xnor U2190 (N_2190,N_1412,N_739);
xnor U2191 (N_2191,N_1343,N_1627);
or U2192 (N_2192,N_1914,N_295);
nor U2193 (N_2193,N_1713,N_1896);
or U2194 (N_2194,N_1065,N_821);
nor U2195 (N_2195,N_860,N_768);
nor U2196 (N_2196,N_20,N_1587);
or U2197 (N_2197,N_1199,N_69);
and U2198 (N_2198,N_1852,N_476);
xnor U2199 (N_2199,N_1172,N_662);
nor U2200 (N_2200,N_1085,N_1641);
xnor U2201 (N_2201,N_711,N_1053);
nand U2202 (N_2202,N_1119,N_467);
nand U2203 (N_2203,N_1674,N_103);
or U2204 (N_2204,N_1588,N_201);
nand U2205 (N_2205,N_1029,N_1462);
nand U2206 (N_2206,N_1478,N_703);
nand U2207 (N_2207,N_1399,N_281);
and U2208 (N_2208,N_183,N_508);
and U2209 (N_2209,N_222,N_1160);
nor U2210 (N_2210,N_832,N_640);
or U2211 (N_2211,N_1489,N_1082);
or U2212 (N_2212,N_1904,N_80);
xnor U2213 (N_2213,N_1035,N_1033);
xor U2214 (N_2214,N_941,N_1293);
nand U2215 (N_2215,N_969,N_770);
and U2216 (N_2216,N_1041,N_173);
xnor U2217 (N_2217,N_460,N_900);
or U2218 (N_2218,N_914,N_491);
nor U2219 (N_2219,N_1621,N_34);
nor U2220 (N_2220,N_1636,N_863);
nand U2221 (N_2221,N_1022,N_1259);
nand U2222 (N_2222,N_692,N_956);
and U2223 (N_2223,N_1210,N_1813);
and U2224 (N_2224,N_1749,N_1750);
nand U2225 (N_2225,N_1966,N_1136);
or U2226 (N_2226,N_254,N_1919);
nor U2227 (N_2227,N_1980,N_1768);
xor U2228 (N_2228,N_464,N_1113);
nor U2229 (N_2229,N_1284,N_1251);
or U2230 (N_2230,N_512,N_305);
or U2231 (N_2231,N_913,N_1530);
nand U2232 (N_2232,N_772,N_383);
and U2233 (N_2233,N_1736,N_1498);
or U2234 (N_2234,N_643,N_162);
nand U2235 (N_2235,N_371,N_1034);
nor U2236 (N_2236,N_1268,N_1821);
or U2237 (N_2237,N_1445,N_188);
xnor U2238 (N_2238,N_134,N_980);
or U2239 (N_2239,N_86,N_1511);
xnor U2240 (N_2240,N_687,N_727);
nor U2241 (N_2241,N_1401,N_1557);
nor U2242 (N_2242,N_728,N_572);
or U2243 (N_2243,N_1555,N_940);
or U2244 (N_2244,N_1786,N_327);
and U2245 (N_2245,N_1395,N_1801);
nand U2246 (N_2246,N_831,N_1358);
xor U2247 (N_2247,N_1471,N_953);
and U2248 (N_2248,N_880,N_1024);
and U2249 (N_2249,N_1138,N_774);
and U2250 (N_2250,N_717,N_565);
nand U2251 (N_2251,N_851,N_1465);
nor U2252 (N_2252,N_1805,N_1744);
or U2253 (N_2253,N_22,N_423);
and U2254 (N_2254,N_1452,N_1148);
nor U2255 (N_2255,N_1196,N_1649);
xnor U2256 (N_2256,N_384,N_653);
nor U2257 (N_2257,N_1917,N_1760);
or U2258 (N_2258,N_1943,N_1309);
or U2259 (N_2259,N_1460,N_660);
nand U2260 (N_2260,N_1667,N_571);
or U2261 (N_2261,N_422,N_335);
nor U2262 (N_2262,N_353,N_28);
nand U2263 (N_2263,N_1746,N_754);
or U2264 (N_2264,N_1889,N_845);
xor U2265 (N_2265,N_420,N_504);
nor U2266 (N_2266,N_377,N_153);
nor U2267 (N_2267,N_1257,N_1482);
and U2268 (N_2268,N_1117,N_136);
nor U2269 (N_2269,N_1921,N_1897);
or U2270 (N_2270,N_1701,N_1049);
nor U2271 (N_2271,N_247,N_256);
or U2272 (N_2272,N_1038,N_99);
nor U2273 (N_2273,N_1036,N_859);
and U2274 (N_2274,N_1984,N_1023);
nand U2275 (N_2275,N_156,N_901);
xor U2276 (N_2276,N_781,N_1270);
or U2277 (N_2277,N_1486,N_1988);
nor U2278 (N_2278,N_0,N_606);
or U2279 (N_2279,N_1870,N_1143);
nand U2280 (N_2280,N_514,N_964);
nand U2281 (N_2281,N_477,N_1319);
nor U2282 (N_2282,N_1865,N_1902);
nand U2283 (N_2283,N_1885,N_1710);
nand U2284 (N_2284,N_357,N_1995);
and U2285 (N_2285,N_303,N_1836);
nor U2286 (N_2286,N_1273,N_252);
nor U2287 (N_2287,N_228,N_1450);
xor U2288 (N_2288,N_825,N_140);
and U2289 (N_2289,N_1638,N_1122);
nand U2290 (N_2290,N_1769,N_1500);
xor U2291 (N_2291,N_144,N_1359);
xnor U2292 (N_2292,N_1491,N_642);
xor U2293 (N_2293,N_1144,N_1697);
nor U2294 (N_2294,N_1435,N_1484);
nand U2295 (N_2295,N_1110,N_1987);
nor U2296 (N_2296,N_1762,N_722);
xnor U2297 (N_2297,N_593,N_1583);
or U2298 (N_2298,N_1330,N_978);
or U2299 (N_2299,N_1282,N_1441);
or U2300 (N_2300,N_1158,N_1569);
nor U2301 (N_2301,N_44,N_744);
and U2302 (N_2302,N_1546,N_1171);
xnor U2303 (N_2303,N_200,N_1021);
and U2304 (N_2304,N_1413,N_345);
nand U2305 (N_2305,N_526,N_646);
and U2306 (N_2306,N_399,N_1808);
xor U2307 (N_2307,N_248,N_1425);
and U2308 (N_2308,N_1344,N_376);
nor U2309 (N_2309,N_672,N_1751);
xor U2310 (N_2310,N_386,N_932);
and U2311 (N_2311,N_1624,N_674);
and U2312 (N_2312,N_1338,N_979);
xnor U2313 (N_2313,N_867,N_1528);
nand U2314 (N_2314,N_534,N_1967);
xnor U2315 (N_2315,N_1072,N_57);
or U2316 (N_2316,N_396,N_996);
nor U2317 (N_2317,N_403,N_1945);
nand U2318 (N_2318,N_348,N_1107);
or U2319 (N_2319,N_1503,N_559);
nand U2320 (N_2320,N_879,N_112);
and U2321 (N_2321,N_782,N_435);
nand U2322 (N_2322,N_1592,N_853);
or U2323 (N_2323,N_190,N_1492);
and U2324 (N_2324,N_1238,N_1521);
nor U2325 (N_2325,N_1757,N_877);
xor U2326 (N_2326,N_517,N_267);
or U2327 (N_2327,N_53,N_1058);
xnor U2328 (N_2328,N_535,N_240);
and U2329 (N_2329,N_1679,N_592);
and U2330 (N_2330,N_1272,N_1316);
nand U2331 (N_2331,N_767,N_994);
xnor U2332 (N_2332,N_790,N_609);
nor U2333 (N_2333,N_1020,N_1133);
nor U2334 (N_2334,N_425,N_158);
nand U2335 (N_2335,N_603,N_1447);
and U2336 (N_2336,N_950,N_614);
and U2337 (N_2337,N_733,N_694);
xnor U2338 (N_2338,N_1579,N_708);
nor U2339 (N_2339,N_344,N_1505);
and U2340 (N_2340,N_1325,N_1796);
or U2341 (N_2341,N_567,N_1102);
and U2342 (N_2342,N_797,N_1229);
xnor U2343 (N_2343,N_1563,N_328);
nand U2344 (N_2344,N_1101,N_888);
or U2345 (N_2345,N_724,N_1256);
nor U2346 (N_2346,N_1797,N_400);
and U2347 (N_2347,N_181,N_1982);
and U2348 (N_2348,N_1504,N_1385);
nand U2349 (N_2349,N_1572,N_289);
nor U2350 (N_2350,N_1913,N_1514);
and U2351 (N_2351,N_1285,N_651);
nor U2352 (N_2352,N_1318,N_788);
or U2353 (N_2353,N_1738,N_1832);
and U2354 (N_2354,N_649,N_756);
nor U2355 (N_2355,N_1989,N_1202);
and U2356 (N_2356,N_427,N_1968);
nor U2357 (N_2357,N_783,N_1981);
and U2358 (N_2358,N_1619,N_579);
xnor U2359 (N_2359,N_147,N_1720);
and U2360 (N_2360,N_1420,N_874);
or U2361 (N_2361,N_1724,N_109);
and U2362 (N_2362,N_1314,N_1522);
xor U2363 (N_2363,N_1222,N_1);
xnor U2364 (N_2364,N_1999,N_1427);
nand U2365 (N_2365,N_1567,N_1828);
or U2366 (N_2366,N_1375,N_887);
and U2367 (N_2367,N_1218,N_192);
or U2368 (N_2368,N_1368,N_1004);
and U2369 (N_2369,N_1307,N_1864);
nand U2370 (N_2370,N_850,N_891);
nor U2371 (N_2371,N_483,N_82);
nand U2372 (N_2372,N_628,N_1673);
or U2373 (N_2373,N_1379,N_178);
nand U2374 (N_2374,N_1878,N_446);
and U2375 (N_2375,N_1915,N_1062);
nand U2376 (N_2376,N_182,N_58);
xor U2377 (N_2377,N_548,N_287);
nand U2378 (N_2378,N_64,N_927);
xnor U2379 (N_2379,N_1407,N_276);
nand U2380 (N_2380,N_990,N_250);
and U2381 (N_2381,N_1524,N_1666);
or U2382 (N_2382,N_417,N_1198);
nor U2383 (N_2383,N_1430,N_1271);
nand U2384 (N_2384,N_755,N_1597);
or U2385 (N_2385,N_988,N_669);
xor U2386 (N_2386,N_232,N_753);
or U2387 (N_2387,N_916,N_1378);
and U2388 (N_2388,N_1942,N_747);
nor U2389 (N_2389,N_1664,N_1827);
nor U2390 (N_2390,N_1096,N_299);
or U2391 (N_2391,N_1591,N_608);
nand U2392 (N_2392,N_1173,N_1695);
nor U2393 (N_2393,N_1814,N_676);
nor U2394 (N_2394,N_1495,N_1979);
or U2395 (N_2395,N_749,N_1778);
xnor U2396 (N_2396,N_1108,N_957);
nor U2397 (N_2397,N_902,N_1217);
nor U2398 (N_2398,N_1684,N_657);
xor U2399 (N_2399,N_1182,N_776);
or U2400 (N_2400,N_626,N_142);
and U2401 (N_2401,N_905,N_428);
nand U2402 (N_2402,N_1806,N_654);
xor U2403 (N_2403,N_1647,N_33);
nor U2404 (N_2404,N_760,N_666);
xor U2405 (N_2405,N_1261,N_36);
nand U2406 (N_2406,N_1468,N_1881);
or U2407 (N_2407,N_1012,N_1879);
or U2408 (N_2408,N_32,N_1179);
and U2409 (N_2409,N_707,N_187);
or U2410 (N_2410,N_1454,N_1262);
xnor U2411 (N_2411,N_1650,N_92);
xnor U2412 (N_2412,N_737,N_589);
nand U2413 (N_2413,N_1765,N_1960);
and U2414 (N_2414,N_679,N_1859);
or U2415 (N_2415,N_284,N_892);
xnor U2416 (N_2416,N_1737,N_196);
nand U2417 (N_2417,N_1011,N_1911);
xor U2418 (N_2418,N_260,N_730);
or U2419 (N_2419,N_1106,N_1166);
xor U2420 (N_2420,N_1895,N_1955);
and U2421 (N_2421,N_280,N_1809);
nand U2422 (N_2422,N_1326,N_309);
nor U2423 (N_2423,N_194,N_426);
and U2424 (N_2424,N_1267,N_634);
nand U2425 (N_2425,N_94,N_1890);
xnor U2426 (N_2426,N_1123,N_81);
and U2427 (N_2427,N_1752,N_904);
nand U2428 (N_2428,N_910,N_1655);
nor U2429 (N_2429,N_1060,N_684);
and U2430 (N_2430,N_1907,N_430);
or U2431 (N_2431,N_1643,N_243);
and U2432 (N_2432,N_169,N_210);
or U2433 (N_2433,N_937,N_577);
nor U2434 (N_2434,N_713,N_949);
nor U2435 (N_2435,N_658,N_55);
nor U2436 (N_2436,N_356,N_137);
nand U2437 (N_2437,N_394,N_1756);
and U2438 (N_2438,N_765,N_1130);
nor U2439 (N_2439,N_492,N_1873);
nor U2440 (N_2440,N_191,N_898);
nor U2441 (N_2441,N_424,N_1735);
xnor U2442 (N_2442,N_946,N_19);
xor U2443 (N_2443,N_1371,N_1554);
xor U2444 (N_2444,N_993,N_110);
and U2445 (N_2445,N_1812,N_1120);
nor U2446 (N_2446,N_163,N_324);
xnor U2447 (N_2447,N_1978,N_1893);
or U2448 (N_2448,N_698,N_1869);
or U2449 (N_2449,N_685,N_66);
and U2450 (N_2450,N_740,N_76);
nand U2451 (N_2451,N_1315,N_1541);
nand U2452 (N_2452,N_1731,N_1165);
nor U2453 (N_2453,N_18,N_1651);
nor U2454 (N_2454,N_1347,N_149);
and U2455 (N_2455,N_764,N_1043);
or U2456 (N_2456,N_1320,N_830);
nand U2457 (N_2457,N_1480,N_1431);
xor U2458 (N_2458,N_489,N_595);
or U2459 (N_2459,N_793,N_804);
xor U2460 (N_2460,N_1950,N_225);
nand U2461 (N_2461,N_1008,N_1088);
and U2462 (N_2462,N_732,N_1721);
nor U2463 (N_2463,N_596,N_561);
and U2464 (N_2464,N_347,N_1404);
nand U2465 (N_2465,N_1613,N_468);
nand U2466 (N_2466,N_1658,N_1032);
or U2467 (N_2467,N_792,N_278);
xor U2468 (N_2468,N_869,N_629);
nor U2469 (N_2469,N_331,N_545);
nand U2470 (N_2470,N_1416,N_878);
nand U2471 (N_2471,N_298,N_145);
nand U2472 (N_2472,N_1124,N_1277);
nor U2473 (N_2473,N_955,N_1834);
nor U2474 (N_2474,N_1582,N_1715);
xnor U2475 (N_2475,N_1656,N_198);
xnor U2476 (N_2476,N_1965,N_117);
or U2477 (N_2477,N_1899,N_1520);
xnor U2478 (N_2478,N_700,N_1607);
and U2479 (N_2479,N_818,N_706);
or U2480 (N_2480,N_922,N_1104);
and U2481 (N_2481,N_1748,N_285);
nor U2482 (N_2482,N_440,N_1985);
xor U2483 (N_2483,N_1103,N_68);
nor U2484 (N_2484,N_97,N_7);
nand U2485 (N_2485,N_965,N_1081);
xor U2486 (N_2486,N_1526,N_1135);
xnor U2487 (N_2487,N_1788,N_321);
nor U2488 (N_2488,N_1176,N_450);
or U2489 (N_2489,N_151,N_715);
or U2490 (N_2490,N_1055,N_406);
xor U2491 (N_2491,N_1547,N_991);
and U2492 (N_2492,N_1411,N_1220);
xor U2493 (N_2493,N_174,N_931);
or U2494 (N_2494,N_936,N_124);
or U2495 (N_2495,N_800,N_1974);
xnor U2496 (N_2496,N_16,N_1028);
nor U2497 (N_2497,N_1704,N_475);
nor U2498 (N_2498,N_478,N_38);
nand U2499 (N_2499,N_743,N_392);
and U2500 (N_2500,N_1860,N_207);
and U2501 (N_2501,N_1449,N_1071);
and U2502 (N_2502,N_443,N_257);
nor U2503 (N_2503,N_1150,N_1850);
and U2504 (N_2504,N_52,N_1977);
xor U2505 (N_2505,N_1383,N_405);
and U2506 (N_2506,N_310,N_917);
nor U2507 (N_2507,N_735,N_1543);
nor U2508 (N_2508,N_336,N_1438);
nand U2509 (N_2509,N_1603,N_573);
nor U2510 (N_2510,N_393,N_1617);
nand U2511 (N_2511,N_1191,N_1565);
and U2512 (N_2512,N_1337,N_461);
nand U2513 (N_2513,N_1244,N_155);
or U2514 (N_2514,N_106,N_1538);
xnor U2515 (N_2515,N_1197,N_387);
nand U2516 (N_2516,N_330,N_264);
nand U2517 (N_2517,N_1799,N_1506);
xor U2518 (N_2518,N_1027,N_249);
nand U2519 (N_2519,N_1488,N_209);
or U2520 (N_2520,N_262,N_165);
nand U2521 (N_2521,N_1831,N_113);
nand U2522 (N_2522,N_1717,N_1232);
and U2523 (N_2523,N_532,N_925);
xnor U2524 (N_2524,N_1903,N_1249);
or U2525 (N_2525,N_359,N_746);
and U2526 (N_2526,N_1469,N_709);
nor U2527 (N_2527,N_1698,N_854);
xnor U2528 (N_2528,N_365,N_494);
and U2529 (N_2529,N_817,N_261);
nand U2530 (N_2530,N_496,N_60);
or U2531 (N_2531,N_1804,N_1064);
or U2532 (N_2532,N_906,N_1374);
xnor U2533 (N_2533,N_293,N_1761);
xnor U2534 (N_2534,N_306,N_1856);
nor U2535 (N_2535,N_1910,N_203);
nor U2536 (N_2536,N_1025,N_1940);
xor U2537 (N_2537,N_419,N_221);
nor U2538 (N_2538,N_570,N_928);
xor U2539 (N_2539,N_814,N_389);
nor U2540 (N_2540,N_1623,N_856);
nor U2541 (N_2541,N_857,N_1304);
and U2542 (N_2542,N_15,N_67);
and U2543 (N_2543,N_1677,N_766);
and U2544 (N_2544,N_824,N_1298);
or U2545 (N_2545,N_502,N_1187);
and U2546 (N_2546,N_1930,N_1996);
or U2547 (N_2547,N_409,N_1525);
nor U2548 (N_2548,N_1798,N_308);
or U2549 (N_2549,N_1440,N_1054);
or U2550 (N_2550,N_1002,N_575);
or U2551 (N_2551,N_600,N_447);
xnor U2552 (N_2552,N_1365,N_63);
nand U2553 (N_2553,N_1685,N_1938);
nand U2554 (N_2554,N_1214,N_1009);
or U2555 (N_2555,N_1351,N_610);
nor U2556 (N_2556,N_1353,N_1993);
or U2557 (N_2557,N_40,N_98);
xnor U2558 (N_2558,N_358,N_1711);
nand U2559 (N_2559,N_1341,N_947);
nor U2560 (N_2560,N_1800,N_693);
and U2561 (N_2561,N_1992,N_259);
xnor U2562 (N_2562,N_1014,N_1311);
nor U2563 (N_2563,N_795,N_961);
xnor U2564 (N_2564,N_481,N_667);
or U2565 (N_2565,N_908,N_1665);
or U2566 (N_2566,N_334,N_1253);
and U2567 (N_2567,N_1894,N_926);
or U2568 (N_2568,N_1393,N_1954);
and U2569 (N_2569,N_1097,N_214);
nor U2570 (N_2570,N_1847,N_1283);
nand U2571 (N_2571,N_1163,N_1006);
nand U2572 (N_2572,N_523,N_1770);
nor U2573 (N_2573,N_355,N_13);
nand U2574 (N_2574,N_815,N_1692);
nor U2575 (N_2575,N_479,N_688);
and U2576 (N_2576,N_1709,N_631);
or U2577 (N_2577,N_959,N_1397);
nand U2578 (N_2578,N_1959,N_1340);
nand U2579 (N_2579,N_1844,N_26);
and U2580 (N_2580,N_1803,N_1483);
nand U2581 (N_2581,N_325,N_42);
nor U2582 (N_2582,N_886,N_1622);
or U2583 (N_2583,N_1475,N_1231);
xnor U2584 (N_2584,N_1609,N_1877);
nor U2585 (N_2585,N_88,N_1635);
nand U2586 (N_2586,N_170,N_1063);
nor U2587 (N_2587,N_75,N_954);
or U2588 (N_2588,N_661,N_1693);
and U2589 (N_2589,N_1519,N_1951);
nand U2590 (N_2590,N_881,N_1157);
xor U2591 (N_2591,N_1703,N_1215);
xor U2592 (N_2592,N_449,N_1183);
nor U2593 (N_2593,N_463,N_1042);
and U2594 (N_2594,N_1019,N_569);
and U2595 (N_2595,N_1590,N_227);
nand U2596 (N_2596,N_530,N_1306);
and U2597 (N_2597,N_161,N_591);
nor U2598 (N_2598,N_268,N_1345);
nor U2599 (N_2599,N_1593,N_418);
or U2600 (N_2600,N_568,N_1802);
nor U2601 (N_2601,N_317,N_862);
nand U2602 (N_2602,N_627,N_490);
and U2603 (N_2603,N_1886,N_808);
or U2604 (N_2604,N_1280,N_177);
nor U2605 (N_2605,N_484,N_655);
nand U2606 (N_2606,N_1400,N_1147);
or U2607 (N_2607,N_59,N_1287);
nand U2608 (N_2608,N_1947,N_962);
xor U2609 (N_2609,N_1083,N_1884);
nor U2610 (N_2610,N_1975,N_1177);
or U2611 (N_2611,N_1194,N_30);
and U2612 (N_2612,N_1370,N_85);
or U2613 (N_2613,N_1560,N_49);
nor U2614 (N_2614,N_454,N_601);
or U2615 (N_2615,N_1240,N_1376);
xnor U2616 (N_2616,N_1542,N_771);
nor U2617 (N_2617,N_1329,N_1125);
nor U2618 (N_2618,N_1186,N_1516);
xnor U2619 (N_2619,N_78,N_866);
or U2620 (N_2620,N_1840,N_1654);
nor U2621 (N_2621,N_683,N_564);
and U2622 (N_2622,N_1246,N_1755);
or U2623 (N_2623,N_675,N_283);
or U2624 (N_2624,N_723,N_588);
and U2625 (N_2625,N_963,N_31);
nor U2626 (N_2626,N_1678,N_404);
xor U2627 (N_2627,N_442,N_673);
or U2628 (N_2628,N_1105,N_25);
xor U2629 (N_2629,N_633,N_1235);
xnor U2630 (N_2630,N_1523,N_976);
nand U2631 (N_2631,N_1719,N_582);
nor U2632 (N_2632,N_193,N_884);
nor U2633 (N_2633,N_1962,N_1513);
nor U2634 (N_2634,N_179,N_865);
and U2635 (N_2635,N_1016,N_677);
nand U2636 (N_2636,N_1219,N_127);
nand U2637 (N_2637,N_1689,N_995);
nand U2638 (N_2638,N_1137,N_1891);
xor U2639 (N_2639,N_1699,N_734);
or U2640 (N_2640,N_1608,N_1618);
xnor U2641 (N_2641,N_1939,N_721);
or U2642 (N_2642,N_981,N_1324);
nand U2643 (N_2643,N_805,N_1255);
nor U2644 (N_2644,N_1779,N_1949);
or U2645 (N_2645,N_1233,N_1151);
nor U2646 (N_2646,N_1294,N_1846);
and U2647 (N_2647,N_681,N_497);
and U2648 (N_2648,N_1372,N_120);
and U2649 (N_2649,N_1423,N_1793);
xor U2650 (N_2650,N_39,N_230);
or U2651 (N_2651,N_1854,N_819);
and U2652 (N_2652,N_54,N_132);
or U2653 (N_2653,N_1681,N_897);
nand U2654 (N_2654,N_500,N_1189);
nor U2655 (N_2655,N_319,N_332);
xor U2656 (N_2656,N_1216,N_742);
xnor U2657 (N_2657,N_1867,N_220);
xnor U2658 (N_2658,N_1087,N_1835);
or U2659 (N_2659,N_1254,N_1364);
nand U2660 (N_2660,N_542,N_507);
and U2661 (N_2661,N_1625,N_1691);
or U2662 (N_2662,N_311,N_566);
nand U2663 (N_2663,N_624,N_1174);
xnor U2664 (N_2664,N_827,N_1490);
and U2665 (N_2665,N_630,N_920);
nor U2666 (N_2666,N_505,N_1976);
and U2667 (N_2667,N_1453,N_45);
nor U2668 (N_2668,N_1630,N_1707);
nor U2669 (N_2669,N_701,N_686);
and U2670 (N_2670,N_664,N_352);
and U2671 (N_2671,N_17,N_1448);
or U2672 (N_2672,N_369,N_316);
and U2673 (N_2673,N_390,N_304);
nand U2674 (N_2674,N_875,N_1149);
or U2675 (N_2675,N_1550,N_1109);
and U2676 (N_2676,N_930,N_172);
xor U2677 (N_2677,N_716,N_24);
xor U2678 (N_2678,N_282,N_1161);
or U2679 (N_2679,N_451,N_1403);
xor U2680 (N_2680,N_8,N_637);
or U2681 (N_2681,N_948,N_90);
xnor U2682 (N_2682,N_1155,N_1291);
or U2683 (N_2683,N_1352,N_620);
xor U2684 (N_2684,N_648,N_645);
or U2685 (N_2685,N_1824,N_531);
nor U2686 (N_2686,N_618,N_1920);
nor U2687 (N_2687,N_1753,N_1227);
xor U2688 (N_2688,N_202,N_1747);
nor U2689 (N_2689,N_1417,N_786);
or U2690 (N_2690,N_275,N_1092);
and U2691 (N_2691,N_1616,N_1632);
and U2692 (N_2692,N_1837,N_1001);
xnor U2693 (N_2693,N_812,N_1473);
xnor U2694 (N_2694,N_1862,N_1741);
or U2695 (N_2695,N_1510,N_1129);
nand U2696 (N_2696,N_1303,N_1296);
xor U2697 (N_2697,N_154,N_1000);
nand U2698 (N_2698,N_705,N_1494);
xor U2699 (N_2699,N_1264,N_123);
xor U2700 (N_2700,N_93,N_1389);
xnor U2701 (N_2701,N_1424,N_130);
nor U2702 (N_2702,N_180,N_388);
and U2703 (N_2703,N_748,N_725);
xnor U2704 (N_2704,N_1696,N_1121);
nor U2705 (N_2705,N_1201,N_432);
nand U2706 (N_2706,N_975,N_1815);
nand U2707 (N_2707,N_1313,N_300);
nor U2708 (N_2708,N_1931,N_960);
nand U2709 (N_2709,N_294,N_520);
or U2710 (N_2710,N_702,N_241);
and U2711 (N_2711,N_1493,N_1459);
or U2712 (N_2712,N_1653,N_894);
and U2713 (N_2713,N_1575,N_939);
xor U2714 (N_2714,N_56,N_95);
nor U2715 (N_2715,N_176,N_1829);
xnor U2716 (N_2716,N_322,N_584);
nor U2717 (N_2717,N_644,N_1851);
nand U2718 (N_2718,N_899,N_1463);
xor U2719 (N_2719,N_1517,N_1327);
or U2720 (N_2720,N_586,N_379);
xnor U2721 (N_2721,N_605,N_843);
or U2722 (N_2722,N_1971,N_160);
and U2723 (N_2723,N_540,N_1826);
and U2724 (N_2724,N_1209,N_1754);
xor U2725 (N_2725,N_114,N_1357);
nand U2726 (N_2726,N_1339,N_368);
nor U2727 (N_2727,N_1952,N_1290);
nand U2728 (N_2728,N_558,N_541);
nand U2729 (N_2729,N_719,N_138);
or U2730 (N_2730,N_714,N_1111);
nor U2731 (N_2731,N_1868,N_778);
nand U2732 (N_2732,N_625,N_1918);
and U2733 (N_2733,N_982,N_1265);
and U2734 (N_2734,N_912,N_1929);
nor U2735 (N_2735,N_35,N_952);
or U2736 (N_2736,N_1180,N_998);
xor U2737 (N_2737,N_1169,N_84);
nand U2738 (N_2738,N_301,N_401);
nor U2739 (N_2739,N_639,N_1336);
and U2740 (N_2740,N_1003,N_1355);
nand U2741 (N_2741,N_1739,N_297);
and U2742 (N_2742,N_374,N_536);
nand U2743 (N_2743,N_1443,N_594);
and U2744 (N_2744,N_538,N_204);
or U2745 (N_2745,N_1811,N_438);
xnor U2746 (N_2746,N_668,N_342);
nand U2747 (N_2747,N_1508,N_1672);
nor U2748 (N_2748,N_522,N_1539);
and U2749 (N_2749,N_1773,N_62);
and U2750 (N_2750,N_1785,N_1335);
and U2751 (N_2751,N_1391,N_1997);
or U2752 (N_2752,N_1131,N_1882);
and U2753 (N_2753,N_1204,N_563);
or U2754 (N_2754,N_343,N_1780);
and U2755 (N_2755,N_121,N_1758);
nand U2756 (N_2756,N_402,N_611);
nand U2757 (N_2757,N_452,N_852);
and U2758 (N_2758,N_1841,N_543);
xnor U2759 (N_2759,N_1185,N_1600);
nand U2760 (N_2760,N_118,N_1223);
and U2761 (N_2761,N_1195,N_1433);
xor U2762 (N_2762,N_108,N_613);
xor U2763 (N_2763,N_844,N_1245);
nor U2764 (N_2764,N_1898,N_1818);
and U2765 (N_2765,N_48,N_271);
and U2766 (N_2766,N_1146,N_1402);
or U2767 (N_2767,N_1192,N_858);
and U2768 (N_2768,N_217,N_105);
xor U2769 (N_2769,N_89,N_1168);
xor U2770 (N_2770,N_29,N_1928);
nor U2771 (N_2771,N_810,N_1132);
xnor U2772 (N_2772,N_829,N_1286);
or U2773 (N_2773,N_951,N_346);
nor U2774 (N_2774,N_1496,N_395);
nand U2775 (N_2775,N_1377,N_1178);
or U2776 (N_2776,N_456,N_738);
nor U2777 (N_2777,N_1924,N_1093);
xnor U2778 (N_2778,N_143,N_1776);
or U2779 (N_2779,N_1566,N_893);
or U2780 (N_2780,N_1141,N_498);
nand U2781 (N_2781,N_546,N_1250);
nand U2782 (N_2782,N_219,N_1193);
or U2783 (N_2783,N_1934,N_974);
nor U2784 (N_2784,N_1790,N_1718);
nand U2785 (N_2785,N_415,N_128);
nand U2786 (N_2786,N_354,N_689);
xnor U2787 (N_2787,N_1089,N_807);
nor U2788 (N_2788,N_779,N_1944);
or U2789 (N_2789,N_1708,N_1184);
nor U2790 (N_2790,N_663,N_635);
and U2791 (N_2791,N_846,N_1299);
xor U2792 (N_2792,N_1912,N_1275);
and U2793 (N_2793,N_1763,N_1317);
nor U2794 (N_2794,N_506,N_871);
and U2795 (N_2795,N_381,N_1759);
nor U2796 (N_2796,N_736,N_1396);
nand U2797 (N_2797,N_216,N_233);
and U2798 (N_2798,N_465,N_1909);
nor U2799 (N_2799,N_1127,N_1070);
nand U2800 (N_2800,N_1410,N_598);
nand U2801 (N_2801,N_1366,N_699);
nand U2802 (N_2802,N_167,N_1743);
xnor U2803 (N_2803,N_1820,N_208);
nand U2804 (N_2804,N_245,N_367);
and U2805 (N_2805,N_872,N_1686);
xor U2806 (N_2806,N_385,N_1205);
nand U2807 (N_2807,N_265,N_1066);
and U2808 (N_2808,N_338,N_1381);
xnor U2809 (N_2809,N_6,N_1167);
nand U2810 (N_2810,N_1297,N_215);
or U2811 (N_2811,N_890,N_796);
nor U2812 (N_2812,N_1774,N_1687);
or U2813 (N_2813,N_1642,N_578);
xnor U2814 (N_2814,N_696,N_935);
or U2815 (N_2815,N_616,N_513);
or U2816 (N_2816,N_641,N_1497);
or U2817 (N_2817,N_1322,N_1545);
or U2818 (N_2818,N_1553,N_1421);
xnor U2819 (N_2819,N_246,N_333);
xor U2820 (N_2820,N_1386,N_1360);
and U2821 (N_2821,N_697,N_837);
and U2822 (N_2822,N_855,N_803);
nand U2823 (N_2823,N_1839,N_1766);
and U2824 (N_2824,N_1661,N_1046);
nand U2825 (N_2825,N_1095,N_71);
nand U2826 (N_2826,N_1584,N_1986);
and U2827 (N_2827,N_269,N_323);
nor U2828 (N_2828,N_896,N_1723);
or U2829 (N_2829,N_195,N_119);
nor U2830 (N_2830,N_1323,N_175);
nor U2831 (N_2831,N_448,N_104);
nand U2832 (N_2832,N_231,N_785);
xor U2833 (N_2833,N_148,N_1334);
xor U2834 (N_2834,N_1190,N_1057);
or U2835 (N_2835,N_636,N_1288);
nand U2836 (N_2836,N_152,N_1321);
nor U2837 (N_2837,N_895,N_1552);
nand U2838 (N_2838,N_1387,N_126);
nand U2839 (N_2839,N_1331,N_1532);
and U2840 (N_2840,N_1266,N_544);
xor U2841 (N_2841,N_1529,N_553);
nor U2842 (N_2842,N_1926,N_695);
xor U2843 (N_2843,N_1578,N_480);
nor U2844 (N_2844,N_1444,N_410);
xnor U2845 (N_2845,N_1434,N_1044);
nand U2846 (N_2846,N_211,N_987);
xor U2847 (N_2847,N_1279,N_665);
and U2848 (N_2848,N_168,N_726);
nand U2849 (N_2849,N_1906,N_159);
and U2850 (N_2850,N_652,N_270);
nand U2851 (N_2851,N_915,N_1857);
and U2852 (N_2852,N_1671,N_378);
nor U2853 (N_2853,N_487,N_1456);
xnor U2854 (N_2854,N_1437,N_1535);
or U2855 (N_2855,N_291,N_1540);
and U2856 (N_2856,N_1652,N_1464);
nor U2857 (N_2857,N_1276,N_607);
xnor U2858 (N_2858,N_1080,N_1714);
nor U2859 (N_2859,N_1680,N_1634);
nand U2860 (N_2860,N_938,N_466);
nand U2861 (N_2861,N_1937,N_1078);
or U2862 (N_2862,N_1670,N_1361);
nand U2863 (N_2863,N_1013,N_903);
and U2864 (N_2864,N_992,N_612);
nor U2865 (N_2865,N_934,N_150);
and U2866 (N_2866,N_1292,N_1745);
xnor U2867 (N_2867,N_809,N_972);
or U2868 (N_2868,N_1090,N_638);
nand U2869 (N_2869,N_457,N_802);
or U2870 (N_2870,N_1612,N_1030);
xnor U2871 (N_2871,N_1916,N_583);
and U2872 (N_2872,N_1363,N_279);
nor U2873 (N_2873,N_1211,N_307);
and U2874 (N_2874,N_470,N_799);
or U2875 (N_2875,N_1700,N_1556);
nor U2876 (N_2876,N_238,N_1476);
nor U2877 (N_2877,N_100,N_1247);
nor U2878 (N_2878,N_1419,N_604);
or U2879 (N_2879,N_1694,N_615);
nand U2880 (N_2880,N_1941,N_14);
nor U2881 (N_2881,N_1100,N_1373);
nor U2882 (N_2882,N_989,N_1175);
nor U2883 (N_2883,N_813,N_780);
nor U2884 (N_2884,N_1477,N_441);
nand U2885 (N_2885,N_1564,N_296);
nand U2886 (N_2886,N_909,N_1026);
xnor U2887 (N_2887,N_1874,N_973);
and U2888 (N_2888,N_794,N_731);
nand U2889 (N_2889,N_1382,N_1415);
nor U2890 (N_2890,N_885,N_1883);
or U2891 (N_2891,N_1639,N_370);
xnor U2892 (N_2892,N_235,N_1784);
or U2893 (N_2893,N_834,N_729);
xor U2894 (N_2894,N_1515,N_835);
and U2895 (N_2895,N_1990,N_70);
nor U2896 (N_2896,N_350,N_1581);
and U2897 (N_2897,N_971,N_632);
nand U2898 (N_2898,N_599,N_1571);
or U2899 (N_2899,N_840,N_1559);
or U2900 (N_2900,N_1742,N_828);
or U2901 (N_2901,N_1726,N_77);
and U2902 (N_2902,N_1074,N_1958);
or U2903 (N_2903,N_164,N_1274);
and U2904 (N_2904,N_1562,N_495);
nor U2905 (N_2905,N_1887,N_1825);
xnor U2906 (N_2906,N_617,N_197);
or U2907 (N_2907,N_1221,N_921);
and U2908 (N_2908,N_1145,N_515);
nor U2909 (N_2909,N_102,N_806);
xnor U2910 (N_2910,N_510,N_1241);
and U2911 (N_2911,N_537,N_1457);
and U2912 (N_2912,N_274,N_251);
xor U2913 (N_2913,N_1932,N_1925);
nor U2914 (N_2914,N_1390,N_1771);
nor U2915 (N_2915,N_1620,N_436);
or U2916 (N_2916,N_1128,N_1611);
or U2917 (N_2917,N_1596,N_1278);
nor U2918 (N_2918,N_1348,N_1601);
or U2919 (N_2919,N_189,N_1892);
or U2920 (N_2920,N_983,N_1466);
and U2921 (N_2921,N_775,N_554);
nand U2922 (N_2922,N_1843,N_1422);
and U2923 (N_2923,N_1712,N_79);
xor U2924 (N_2924,N_1414,N_1224);
and U2925 (N_2925,N_412,N_1957);
nor U2926 (N_2926,N_1795,N_1037);
nand U2927 (N_2927,N_977,N_549);
nand U2928 (N_2928,N_199,N_1994);
nor U2929 (N_2929,N_421,N_1140);
nor U2930 (N_2930,N_1688,N_72);
or U2931 (N_2931,N_1669,N_1961);
nor U2932 (N_2932,N_1637,N_1972);
or U2933 (N_2933,N_1451,N_1900);
xor U2934 (N_2934,N_462,N_1845);
nand U2935 (N_2935,N_23,N_1644);
nor U2936 (N_2936,N_51,N_1295);
or U2937 (N_2937,N_907,N_439);
xnor U2938 (N_2938,N_1626,N_21);
xnor U2939 (N_2939,N_773,N_889);
nand U2940 (N_2940,N_1040,N_1716);
nor U2941 (N_2941,N_761,N_1998);
or U2942 (N_2942,N_1767,N_1604);
and U2943 (N_2943,N_1568,N_1772);
xor U2944 (N_2944,N_288,N_1730);
or U2945 (N_2945,N_1792,N_650);
and U2946 (N_2946,N_1333,N_1260);
and U2947 (N_2947,N_882,N_1056);
xor U2948 (N_2948,N_1576,N_1733);
xor U2949 (N_2949,N_212,N_1682);
and U2950 (N_2950,N_1933,N_474);
and U2951 (N_2951,N_12,N_1474);
or U2952 (N_2952,N_46,N_1855);
nand U2953 (N_2953,N_129,N_757);
and U2954 (N_2954,N_469,N_186);
xor U2955 (N_2955,N_372,N_1599);
xnor U2956 (N_2956,N_984,N_1946);
nand U2957 (N_2957,N_576,N_1702);
xnor U2958 (N_2958,N_397,N_1069);
xnor U2959 (N_2959,N_313,N_27);
or U2960 (N_2960,N_923,N_1164);
and U2961 (N_2961,N_286,N_1362);
xor U2962 (N_2962,N_1969,N_1631);
or U2963 (N_2963,N_873,N_1384);
xor U2964 (N_2964,N_431,N_1728);
and U2965 (N_2965,N_73,N_1551);
xnor U2966 (N_2966,N_1142,N_1727);
nand U2967 (N_2967,N_1048,N_1794);
and U2968 (N_2968,N_339,N_1817);
or U2969 (N_2969,N_1734,N_266);
or U2970 (N_2970,N_1091,N_986);
nor U2971 (N_2971,N_263,N_398);
nand U2972 (N_2972,N_968,N_1598);
nor U2973 (N_2973,N_1948,N_205);
and U2974 (N_2974,N_1116,N_1350);
xnor U2975 (N_2975,N_619,N_943);
and U2976 (N_2976,N_1970,N_1861);
or U2977 (N_2977,N_1640,N_1310);
nand U2978 (N_2978,N_1629,N_911);
xor U2979 (N_2979,N_139,N_1134);
and U2980 (N_2980,N_1537,N_1580);
xor U2981 (N_2981,N_841,N_482);
xnor U2982 (N_2982,N_966,N_122);
or U2983 (N_2983,N_1098,N_471);
nor U2984 (N_2984,N_1051,N_519);
and U2985 (N_2985,N_1536,N_206);
or U2986 (N_2986,N_587,N_1154);
nand U2987 (N_2987,N_111,N_602);
nor U2988 (N_2988,N_1953,N_1005);
and U2989 (N_2989,N_1935,N_758);
nand U2990 (N_2990,N_349,N_1031);
nor U2991 (N_2991,N_1061,N_883);
nor U2992 (N_2992,N_1871,N_745);
nor U2993 (N_2993,N_364,N_557);
and U2994 (N_2994,N_1683,N_1112);
nor U2995 (N_2995,N_1872,N_659);
nand U2996 (N_2996,N_329,N_1162);
nand U2997 (N_2997,N_1936,N_560);
nor U2998 (N_2998,N_1426,N_1690);
nor U2999 (N_2999,N_1531,N_621);
and U3000 (N_3000,N_529,N_1089);
or U3001 (N_3001,N_1198,N_1016);
xnor U3002 (N_3002,N_1838,N_447);
nor U3003 (N_3003,N_697,N_345);
nor U3004 (N_3004,N_1186,N_1095);
xnor U3005 (N_3005,N_507,N_602);
xnor U3006 (N_3006,N_258,N_820);
and U3007 (N_3007,N_46,N_1691);
xnor U3008 (N_3008,N_1494,N_590);
nor U3009 (N_3009,N_810,N_1489);
or U3010 (N_3010,N_376,N_651);
or U3011 (N_3011,N_1188,N_1753);
nor U3012 (N_3012,N_1376,N_775);
nor U3013 (N_3013,N_402,N_1597);
and U3014 (N_3014,N_1936,N_122);
and U3015 (N_3015,N_1702,N_1877);
nor U3016 (N_3016,N_1586,N_1549);
xor U3017 (N_3017,N_826,N_1861);
nand U3018 (N_3018,N_1538,N_1336);
nor U3019 (N_3019,N_1110,N_159);
nand U3020 (N_3020,N_938,N_1965);
or U3021 (N_3021,N_143,N_892);
and U3022 (N_3022,N_339,N_728);
and U3023 (N_3023,N_932,N_393);
nand U3024 (N_3024,N_1597,N_389);
nor U3025 (N_3025,N_1,N_1056);
or U3026 (N_3026,N_719,N_1463);
and U3027 (N_3027,N_1707,N_268);
xnor U3028 (N_3028,N_1250,N_597);
xnor U3029 (N_3029,N_1628,N_531);
or U3030 (N_3030,N_488,N_575);
xnor U3031 (N_3031,N_1488,N_419);
xor U3032 (N_3032,N_786,N_203);
and U3033 (N_3033,N_969,N_598);
nor U3034 (N_3034,N_1221,N_1241);
nand U3035 (N_3035,N_1841,N_1213);
nand U3036 (N_3036,N_1705,N_1710);
nor U3037 (N_3037,N_460,N_1390);
or U3038 (N_3038,N_1788,N_1781);
nor U3039 (N_3039,N_158,N_919);
or U3040 (N_3040,N_684,N_1483);
and U3041 (N_3041,N_341,N_389);
xnor U3042 (N_3042,N_347,N_507);
xor U3043 (N_3043,N_1030,N_518);
xor U3044 (N_3044,N_107,N_781);
nor U3045 (N_3045,N_1724,N_1200);
or U3046 (N_3046,N_1406,N_563);
nand U3047 (N_3047,N_368,N_378);
or U3048 (N_3048,N_453,N_954);
nor U3049 (N_3049,N_1610,N_1711);
or U3050 (N_3050,N_1290,N_1479);
and U3051 (N_3051,N_1160,N_1472);
or U3052 (N_3052,N_1628,N_41);
or U3053 (N_3053,N_1770,N_93);
or U3054 (N_3054,N_1425,N_42);
xor U3055 (N_3055,N_1086,N_1974);
xnor U3056 (N_3056,N_408,N_139);
xor U3057 (N_3057,N_556,N_886);
nor U3058 (N_3058,N_1928,N_1739);
nand U3059 (N_3059,N_128,N_1943);
xor U3060 (N_3060,N_973,N_99);
nand U3061 (N_3061,N_597,N_177);
and U3062 (N_3062,N_1554,N_1029);
or U3063 (N_3063,N_154,N_708);
and U3064 (N_3064,N_1991,N_1044);
or U3065 (N_3065,N_1720,N_1843);
xor U3066 (N_3066,N_1180,N_1269);
nand U3067 (N_3067,N_1622,N_907);
xor U3068 (N_3068,N_598,N_1360);
nand U3069 (N_3069,N_874,N_400);
xor U3070 (N_3070,N_954,N_1859);
nor U3071 (N_3071,N_1898,N_1051);
or U3072 (N_3072,N_1203,N_1116);
or U3073 (N_3073,N_1036,N_53);
and U3074 (N_3074,N_77,N_319);
nand U3075 (N_3075,N_31,N_189);
nor U3076 (N_3076,N_1375,N_918);
or U3077 (N_3077,N_318,N_951);
nor U3078 (N_3078,N_352,N_631);
xnor U3079 (N_3079,N_462,N_138);
or U3080 (N_3080,N_161,N_1047);
nand U3081 (N_3081,N_1897,N_95);
nor U3082 (N_3082,N_361,N_189);
nand U3083 (N_3083,N_1612,N_1302);
and U3084 (N_3084,N_491,N_1267);
xnor U3085 (N_3085,N_1023,N_1908);
xnor U3086 (N_3086,N_576,N_991);
nor U3087 (N_3087,N_489,N_1478);
and U3088 (N_3088,N_776,N_528);
nand U3089 (N_3089,N_1208,N_1897);
xnor U3090 (N_3090,N_1835,N_1110);
and U3091 (N_3091,N_1182,N_1309);
nand U3092 (N_3092,N_801,N_1442);
xor U3093 (N_3093,N_1228,N_1916);
nand U3094 (N_3094,N_469,N_965);
xor U3095 (N_3095,N_1624,N_1448);
nor U3096 (N_3096,N_1249,N_1098);
or U3097 (N_3097,N_1843,N_1121);
nand U3098 (N_3098,N_1257,N_1261);
nor U3099 (N_3099,N_525,N_1790);
nor U3100 (N_3100,N_1964,N_1229);
nand U3101 (N_3101,N_639,N_577);
nand U3102 (N_3102,N_1477,N_1562);
and U3103 (N_3103,N_769,N_1300);
xnor U3104 (N_3104,N_10,N_1871);
or U3105 (N_3105,N_262,N_750);
or U3106 (N_3106,N_1172,N_774);
nand U3107 (N_3107,N_36,N_277);
nand U3108 (N_3108,N_791,N_1703);
nand U3109 (N_3109,N_1218,N_1432);
or U3110 (N_3110,N_1836,N_1061);
or U3111 (N_3111,N_512,N_1608);
nor U3112 (N_3112,N_1260,N_1746);
and U3113 (N_3113,N_1092,N_366);
and U3114 (N_3114,N_1056,N_1803);
and U3115 (N_3115,N_808,N_1386);
nand U3116 (N_3116,N_939,N_77);
or U3117 (N_3117,N_24,N_1678);
xnor U3118 (N_3118,N_927,N_948);
or U3119 (N_3119,N_425,N_1069);
or U3120 (N_3120,N_5,N_222);
nand U3121 (N_3121,N_1290,N_1573);
or U3122 (N_3122,N_548,N_977);
nor U3123 (N_3123,N_1208,N_383);
nor U3124 (N_3124,N_1454,N_1458);
and U3125 (N_3125,N_444,N_1424);
xor U3126 (N_3126,N_1548,N_796);
nand U3127 (N_3127,N_497,N_209);
xor U3128 (N_3128,N_1513,N_104);
and U3129 (N_3129,N_963,N_1227);
xnor U3130 (N_3130,N_1163,N_1900);
nor U3131 (N_3131,N_1529,N_89);
nand U3132 (N_3132,N_1059,N_276);
and U3133 (N_3133,N_898,N_1008);
xor U3134 (N_3134,N_769,N_1161);
and U3135 (N_3135,N_294,N_643);
nor U3136 (N_3136,N_709,N_230);
nor U3137 (N_3137,N_184,N_389);
nand U3138 (N_3138,N_310,N_323);
or U3139 (N_3139,N_1931,N_235);
nor U3140 (N_3140,N_112,N_597);
or U3141 (N_3141,N_7,N_1167);
nor U3142 (N_3142,N_326,N_1160);
nand U3143 (N_3143,N_1093,N_355);
nand U3144 (N_3144,N_1396,N_402);
and U3145 (N_3145,N_1151,N_147);
nand U3146 (N_3146,N_374,N_1341);
xor U3147 (N_3147,N_627,N_1723);
and U3148 (N_3148,N_242,N_1011);
xor U3149 (N_3149,N_1525,N_11);
nor U3150 (N_3150,N_823,N_1563);
nand U3151 (N_3151,N_1551,N_500);
xor U3152 (N_3152,N_1741,N_1982);
xnor U3153 (N_3153,N_376,N_1946);
or U3154 (N_3154,N_1912,N_1553);
nand U3155 (N_3155,N_250,N_1678);
xor U3156 (N_3156,N_1015,N_1537);
and U3157 (N_3157,N_806,N_1987);
nor U3158 (N_3158,N_741,N_1037);
nor U3159 (N_3159,N_1156,N_904);
and U3160 (N_3160,N_1664,N_734);
or U3161 (N_3161,N_574,N_1197);
nand U3162 (N_3162,N_1243,N_1758);
and U3163 (N_3163,N_1547,N_1149);
nor U3164 (N_3164,N_1670,N_1381);
nand U3165 (N_3165,N_1211,N_1039);
nor U3166 (N_3166,N_641,N_1516);
or U3167 (N_3167,N_444,N_753);
nand U3168 (N_3168,N_1135,N_602);
and U3169 (N_3169,N_1374,N_90);
and U3170 (N_3170,N_1064,N_1347);
or U3171 (N_3171,N_514,N_1309);
or U3172 (N_3172,N_1185,N_1997);
nand U3173 (N_3173,N_1064,N_789);
nand U3174 (N_3174,N_1865,N_127);
and U3175 (N_3175,N_1496,N_14);
nor U3176 (N_3176,N_574,N_1161);
xor U3177 (N_3177,N_370,N_143);
nor U3178 (N_3178,N_818,N_134);
nand U3179 (N_3179,N_995,N_327);
xor U3180 (N_3180,N_1283,N_1979);
or U3181 (N_3181,N_583,N_568);
nand U3182 (N_3182,N_825,N_1259);
xor U3183 (N_3183,N_1118,N_655);
nand U3184 (N_3184,N_1373,N_1684);
nor U3185 (N_3185,N_240,N_1999);
and U3186 (N_3186,N_772,N_246);
nor U3187 (N_3187,N_1657,N_932);
nand U3188 (N_3188,N_636,N_608);
and U3189 (N_3189,N_1196,N_131);
xnor U3190 (N_3190,N_187,N_1088);
or U3191 (N_3191,N_1632,N_1575);
and U3192 (N_3192,N_484,N_563);
or U3193 (N_3193,N_172,N_893);
nand U3194 (N_3194,N_608,N_1742);
xnor U3195 (N_3195,N_299,N_1823);
and U3196 (N_3196,N_1612,N_1346);
or U3197 (N_3197,N_633,N_1779);
nor U3198 (N_3198,N_1392,N_649);
or U3199 (N_3199,N_683,N_887);
nor U3200 (N_3200,N_1158,N_1950);
and U3201 (N_3201,N_1704,N_66);
nand U3202 (N_3202,N_1300,N_181);
and U3203 (N_3203,N_1209,N_1469);
and U3204 (N_3204,N_734,N_1012);
or U3205 (N_3205,N_628,N_1784);
nand U3206 (N_3206,N_1073,N_1255);
nand U3207 (N_3207,N_1273,N_1659);
and U3208 (N_3208,N_885,N_1557);
xor U3209 (N_3209,N_601,N_309);
nand U3210 (N_3210,N_82,N_732);
nand U3211 (N_3211,N_141,N_796);
and U3212 (N_3212,N_1485,N_249);
xor U3213 (N_3213,N_163,N_488);
and U3214 (N_3214,N_1844,N_906);
nor U3215 (N_3215,N_1697,N_1598);
xor U3216 (N_3216,N_255,N_1923);
or U3217 (N_3217,N_1724,N_163);
and U3218 (N_3218,N_1870,N_1077);
nor U3219 (N_3219,N_1806,N_1096);
nor U3220 (N_3220,N_664,N_1058);
nand U3221 (N_3221,N_1541,N_326);
and U3222 (N_3222,N_1142,N_1399);
nand U3223 (N_3223,N_1960,N_1495);
xnor U3224 (N_3224,N_1891,N_32);
nand U3225 (N_3225,N_252,N_1124);
nor U3226 (N_3226,N_1088,N_1771);
nand U3227 (N_3227,N_24,N_983);
nor U3228 (N_3228,N_887,N_1078);
nand U3229 (N_3229,N_963,N_1949);
or U3230 (N_3230,N_1632,N_1882);
xnor U3231 (N_3231,N_929,N_59);
nand U3232 (N_3232,N_765,N_1291);
xor U3233 (N_3233,N_1804,N_1753);
nor U3234 (N_3234,N_393,N_384);
and U3235 (N_3235,N_112,N_1574);
xor U3236 (N_3236,N_622,N_1982);
nand U3237 (N_3237,N_1666,N_941);
and U3238 (N_3238,N_1590,N_599);
and U3239 (N_3239,N_785,N_150);
or U3240 (N_3240,N_252,N_401);
nor U3241 (N_3241,N_1275,N_958);
nor U3242 (N_3242,N_697,N_1031);
and U3243 (N_3243,N_730,N_206);
xor U3244 (N_3244,N_951,N_1171);
nand U3245 (N_3245,N_29,N_658);
and U3246 (N_3246,N_1283,N_1977);
nand U3247 (N_3247,N_221,N_915);
or U3248 (N_3248,N_1412,N_1577);
xnor U3249 (N_3249,N_495,N_1225);
nor U3250 (N_3250,N_282,N_1905);
or U3251 (N_3251,N_424,N_1200);
and U3252 (N_3252,N_1105,N_615);
and U3253 (N_3253,N_428,N_602);
or U3254 (N_3254,N_1824,N_191);
or U3255 (N_3255,N_1417,N_1241);
or U3256 (N_3256,N_1855,N_117);
or U3257 (N_3257,N_95,N_1549);
nor U3258 (N_3258,N_1974,N_425);
and U3259 (N_3259,N_238,N_788);
or U3260 (N_3260,N_72,N_536);
xnor U3261 (N_3261,N_1669,N_129);
and U3262 (N_3262,N_460,N_399);
xnor U3263 (N_3263,N_1542,N_1350);
nand U3264 (N_3264,N_1233,N_1767);
or U3265 (N_3265,N_1511,N_1022);
xnor U3266 (N_3266,N_1079,N_1467);
and U3267 (N_3267,N_1151,N_739);
and U3268 (N_3268,N_26,N_800);
nand U3269 (N_3269,N_1060,N_120);
nand U3270 (N_3270,N_232,N_1368);
or U3271 (N_3271,N_1324,N_1584);
nand U3272 (N_3272,N_1566,N_969);
or U3273 (N_3273,N_1865,N_1006);
nor U3274 (N_3274,N_1063,N_201);
xor U3275 (N_3275,N_78,N_1580);
and U3276 (N_3276,N_1787,N_967);
and U3277 (N_3277,N_404,N_1859);
xor U3278 (N_3278,N_1601,N_1290);
xnor U3279 (N_3279,N_1491,N_364);
xnor U3280 (N_3280,N_1889,N_1433);
xnor U3281 (N_3281,N_1611,N_884);
or U3282 (N_3282,N_147,N_89);
nand U3283 (N_3283,N_1271,N_1890);
nand U3284 (N_3284,N_257,N_11);
nand U3285 (N_3285,N_598,N_724);
xor U3286 (N_3286,N_999,N_97);
nor U3287 (N_3287,N_1973,N_372);
or U3288 (N_3288,N_417,N_832);
or U3289 (N_3289,N_1537,N_806);
and U3290 (N_3290,N_243,N_549);
and U3291 (N_3291,N_1474,N_1550);
nor U3292 (N_3292,N_194,N_729);
and U3293 (N_3293,N_799,N_1358);
xor U3294 (N_3294,N_750,N_324);
nand U3295 (N_3295,N_1559,N_1730);
nor U3296 (N_3296,N_612,N_323);
nor U3297 (N_3297,N_91,N_449);
and U3298 (N_3298,N_132,N_1284);
and U3299 (N_3299,N_1674,N_259);
or U3300 (N_3300,N_659,N_1790);
nand U3301 (N_3301,N_339,N_1528);
xor U3302 (N_3302,N_857,N_1311);
or U3303 (N_3303,N_515,N_1249);
and U3304 (N_3304,N_1539,N_811);
nor U3305 (N_3305,N_1927,N_1020);
nor U3306 (N_3306,N_1189,N_1789);
and U3307 (N_3307,N_28,N_596);
and U3308 (N_3308,N_265,N_1384);
nand U3309 (N_3309,N_496,N_1437);
or U3310 (N_3310,N_636,N_1306);
nand U3311 (N_3311,N_1590,N_1117);
xnor U3312 (N_3312,N_1069,N_938);
nand U3313 (N_3313,N_368,N_1162);
nand U3314 (N_3314,N_1260,N_1370);
nor U3315 (N_3315,N_765,N_611);
xnor U3316 (N_3316,N_111,N_645);
xor U3317 (N_3317,N_960,N_1978);
xor U3318 (N_3318,N_1423,N_752);
and U3319 (N_3319,N_1809,N_1028);
and U3320 (N_3320,N_1344,N_1922);
or U3321 (N_3321,N_1627,N_571);
or U3322 (N_3322,N_1625,N_1850);
nand U3323 (N_3323,N_1147,N_1710);
nor U3324 (N_3324,N_897,N_421);
and U3325 (N_3325,N_1217,N_1247);
and U3326 (N_3326,N_1986,N_1597);
and U3327 (N_3327,N_444,N_1953);
or U3328 (N_3328,N_863,N_946);
nand U3329 (N_3329,N_1434,N_1215);
xnor U3330 (N_3330,N_606,N_112);
nand U3331 (N_3331,N_1694,N_703);
or U3332 (N_3332,N_855,N_1321);
or U3333 (N_3333,N_320,N_33);
nor U3334 (N_3334,N_1488,N_1474);
xor U3335 (N_3335,N_1168,N_1461);
xor U3336 (N_3336,N_506,N_1258);
and U3337 (N_3337,N_1113,N_297);
and U3338 (N_3338,N_1574,N_1154);
or U3339 (N_3339,N_1430,N_670);
nand U3340 (N_3340,N_1388,N_1082);
and U3341 (N_3341,N_819,N_658);
nor U3342 (N_3342,N_1925,N_137);
nor U3343 (N_3343,N_1405,N_1021);
and U3344 (N_3344,N_1056,N_818);
nand U3345 (N_3345,N_558,N_759);
nand U3346 (N_3346,N_828,N_1341);
or U3347 (N_3347,N_697,N_465);
and U3348 (N_3348,N_1365,N_1040);
nor U3349 (N_3349,N_1385,N_676);
nor U3350 (N_3350,N_36,N_965);
or U3351 (N_3351,N_94,N_484);
nand U3352 (N_3352,N_1554,N_1076);
and U3353 (N_3353,N_1111,N_1123);
xnor U3354 (N_3354,N_763,N_1905);
xor U3355 (N_3355,N_1631,N_302);
or U3356 (N_3356,N_1351,N_657);
or U3357 (N_3357,N_580,N_200);
and U3358 (N_3358,N_1290,N_175);
xnor U3359 (N_3359,N_1435,N_1316);
and U3360 (N_3360,N_513,N_460);
and U3361 (N_3361,N_1422,N_203);
and U3362 (N_3362,N_424,N_13);
and U3363 (N_3363,N_1415,N_910);
nor U3364 (N_3364,N_481,N_609);
xor U3365 (N_3365,N_1407,N_997);
or U3366 (N_3366,N_1366,N_1766);
nand U3367 (N_3367,N_189,N_1948);
nor U3368 (N_3368,N_696,N_130);
or U3369 (N_3369,N_1069,N_401);
nand U3370 (N_3370,N_1836,N_1419);
xor U3371 (N_3371,N_1923,N_1115);
and U3372 (N_3372,N_1176,N_1934);
nor U3373 (N_3373,N_39,N_21);
or U3374 (N_3374,N_680,N_399);
xor U3375 (N_3375,N_671,N_1554);
nor U3376 (N_3376,N_1988,N_390);
xnor U3377 (N_3377,N_437,N_979);
or U3378 (N_3378,N_1447,N_934);
xnor U3379 (N_3379,N_546,N_543);
xnor U3380 (N_3380,N_793,N_711);
or U3381 (N_3381,N_1500,N_999);
nor U3382 (N_3382,N_808,N_1883);
nand U3383 (N_3383,N_290,N_1468);
nand U3384 (N_3384,N_729,N_879);
nor U3385 (N_3385,N_249,N_1798);
xnor U3386 (N_3386,N_492,N_871);
nor U3387 (N_3387,N_313,N_1549);
and U3388 (N_3388,N_1341,N_707);
and U3389 (N_3389,N_110,N_1658);
or U3390 (N_3390,N_1632,N_673);
or U3391 (N_3391,N_1205,N_1874);
or U3392 (N_3392,N_1497,N_1424);
or U3393 (N_3393,N_1176,N_886);
xor U3394 (N_3394,N_1709,N_1345);
nor U3395 (N_3395,N_323,N_434);
or U3396 (N_3396,N_1484,N_82);
or U3397 (N_3397,N_507,N_644);
or U3398 (N_3398,N_388,N_662);
nand U3399 (N_3399,N_1386,N_1971);
nand U3400 (N_3400,N_185,N_1972);
xnor U3401 (N_3401,N_1468,N_1918);
nor U3402 (N_3402,N_1086,N_1929);
nand U3403 (N_3403,N_844,N_1975);
nor U3404 (N_3404,N_709,N_208);
nand U3405 (N_3405,N_122,N_332);
and U3406 (N_3406,N_1546,N_1944);
nand U3407 (N_3407,N_940,N_643);
xor U3408 (N_3408,N_437,N_1400);
nor U3409 (N_3409,N_1558,N_476);
or U3410 (N_3410,N_514,N_17);
xnor U3411 (N_3411,N_1506,N_1734);
nor U3412 (N_3412,N_1974,N_1710);
and U3413 (N_3413,N_152,N_1624);
nand U3414 (N_3414,N_810,N_1246);
or U3415 (N_3415,N_1151,N_1970);
nand U3416 (N_3416,N_1337,N_712);
xnor U3417 (N_3417,N_1347,N_1986);
xnor U3418 (N_3418,N_1662,N_1618);
or U3419 (N_3419,N_677,N_946);
and U3420 (N_3420,N_1275,N_1874);
nor U3421 (N_3421,N_1552,N_299);
xor U3422 (N_3422,N_537,N_430);
or U3423 (N_3423,N_239,N_398);
nand U3424 (N_3424,N_801,N_39);
xnor U3425 (N_3425,N_1820,N_130);
and U3426 (N_3426,N_1974,N_330);
or U3427 (N_3427,N_1265,N_695);
nand U3428 (N_3428,N_370,N_1317);
or U3429 (N_3429,N_867,N_575);
nand U3430 (N_3430,N_1557,N_1715);
or U3431 (N_3431,N_721,N_280);
nand U3432 (N_3432,N_1399,N_1049);
xor U3433 (N_3433,N_791,N_1196);
nor U3434 (N_3434,N_391,N_812);
nor U3435 (N_3435,N_1676,N_950);
or U3436 (N_3436,N_1637,N_444);
nand U3437 (N_3437,N_12,N_1336);
xnor U3438 (N_3438,N_1366,N_1409);
or U3439 (N_3439,N_430,N_1060);
nand U3440 (N_3440,N_519,N_35);
xor U3441 (N_3441,N_1010,N_1823);
nand U3442 (N_3442,N_715,N_787);
nand U3443 (N_3443,N_291,N_1443);
and U3444 (N_3444,N_1721,N_58);
and U3445 (N_3445,N_429,N_1946);
or U3446 (N_3446,N_1490,N_1180);
and U3447 (N_3447,N_1216,N_510);
or U3448 (N_3448,N_1864,N_674);
nor U3449 (N_3449,N_522,N_478);
or U3450 (N_3450,N_347,N_1723);
nand U3451 (N_3451,N_1610,N_1659);
nand U3452 (N_3452,N_499,N_72);
or U3453 (N_3453,N_198,N_922);
nand U3454 (N_3454,N_1522,N_1581);
nand U3455 (N_3455,N_1237,N_59);
xnor U3456 (N_3456,N_278,N_466);
and U3457 (N_3457,N_844,N_1597);
nor U3458 (N_3458,N_1793,N_909);
and U3459 (N_3459,N_615,N_768);
or U3460 (N_3460,N_1773,N_222);
nand U3461 (N_3461,N_942,N_1843);
nand U3462 (N_3462,N_515,N_728);
and U3463 (N_3463,N_303,N_45);
or U3464 (N_3464,N_1109,N_1699);
nand U3465 (N_3465,N_1571,N_1987);
or U3466 (N_3466,N_1032,N_1724);
or U3467 (N_3467,N_1129,N_702);
xor U3468 (N_3468,N_1861,N_1392);
nor U3469 (N_3469,N_345,N_1419);
nor U3470 (N_3470,N_890,N_1387);
xnor U3471 (N_3471,N_1456,N_204);
and U3472 (N_3472,N_1492,N_1317);
nor U3473 (N_3473,N_911,N_740);
xnor U3474 (N_3474,N_966,N_1299);
or U3475 (N_3475,N_1027,N_822);
xor U3476 (N_3476,N_1970,N_147);
and U3477 (N_3477,N_1623,N_1883);
and U3478 (N_3478,N_1730,N_1463);
xor U3479 (N_3479,N_1142,N_1541);
nor U3480 (N_3480,N_1074,N_790);
nor U3481 (N_3481,N_1217,N_1805);
nand U3482 (N_3482,N_1712,N_293);
or U3483 (N_3483,N_981,N_1416);
or U3484 (N_3484,N_1975,N_647);
nand U3485 (N_3485,N_593,N_1051);
or U3486 (N_3486,N_1673,N_1548);
and U3487 (N_3487,N_110,N_179);
xor U3488 (N_3488,N_1463,N_850);
nor U3489 (N_3489,N_1809,N_322);
xnor U3490 (N_3490,N_214,N_245);
nor U3491 (N_3491,N_1878,N_1242);
and U3492 (N_3492,N_46,N_180);
and U3493 (N_3493,N_1255,N_864);
or U3494 (N_3494,N_186,N_485);
xnor U3495 (N_3495,N_26,N_1063);
or U3496 (N_3496,N_1205,N_274);
nand U3497 (N_3497,N_1428,N_1425);
xor U3498 (N_3498,N_1754,N_106);
nor U3499 (N_3499,N_1662,N_1442);
or U3500 (N_3500,N_920,N_1938);
and U3501 (N_3501,N_1173,N_1506);
or U3502 (N_3502,N_1934,N_1135);
nor U3503 (N_3503,N_1097,N_1621);
nand U3504 (N_3504,N_1204,N_23);
or U3505 (N_3505,N_1342,N_1778);
or U3506 (N_3506,N_326,N_652);
xor U3507 (N_3507,N_1631,N_1724);
nor U3508 (N_3508,N_1954,N_1467);
and U3509 (N_3509,N_426,N_1415);
and U3510 (N_3510,N_1041,N_221);
or U3511 (N_3511,N_448,N_494);
nand U3512 (N_3512,N_459,N_1750);
xnor U3513 (N_3513,N_1187,N_1876);
and U3514 (N_3514,N_228,N_1332);
nor U3515 (N_3515,N_1360,N_1720);
nor U3516 (N_3516,N_41,N_777);
or U3517 (N_3517,N_1264,N_362);
xor U3518 (N_3518,N_722,N_901);
nand U3519 (N_3519,N_45,N_1754);
nand U3520 (N_3520,N_212,N_562);
nor U3521 (N_3521,N_545,N_407);
nand U3522 (N_3522,N_1792,N_717);
xor U3523 (N_3523,N_1183,N_1060);
xnor U3524 (N_3524,N_198,N_1942);
nor U3525 (N_3525,N_1425,N_487);
xor U3526 (N_3526,N_1491,N_698);
or U3527 (N_3527,N_1900,N_1128);
and U3528 (N_3528,N_1666,N_762);
nand U3529 (N_3529,N_1734,N_1872);
nor U3530 (N_3530,N_1066,N_1057);
xnor U3531 (N_3531,N_812,N_913);
and U3532 (N_3532,N_1241,N_678);
nand U3533 (N_3533,N_1432,N_356);
nor U3534 (N_3534,N_1197,N_274);
xnor U3535 (N_3535,N_326,N_52);
and U3536 (N_3536,N_605,N_1641);
and U3537 (N_3537,N_745,N_1149);
or U3538 (N_3538,N_1681,N_1158);
xnor U3539 (N_3539,N_1396,N_1596);
nand U3540 (N_3540,N_1299,N_979);
nor U3541 (N_3541,N_1812,N_44);
or U3542 (N_3542,N_1793,N_334);
xor U3543 (N_3543,N_858,N_125);
and U3544 (N_3544,N_428,N_588);
nand U3545 (N_3545,N_1351,N_1410);
or U3546 (N_3546,N_1410,N_1833);
nor U3547 (N_3547,N_1180,N_205);
nand U3548 (N_3548,N_1405,N_823);
xor U3549 (N_3549,N_637,N_521);
xnor U3550 (N_3550,N_1549,N_992);
and U3551 (N_3551,N_1512,N_1067);
nor U3552 (N_3552,N_1002,N_1996);
nand U3553 (N_3553,N_175,N_1934);
nor U3554 (N_3554,N_1486,N_1002);
or U3555 (N_3555,N_623,N_107);
and U3556 (N_3556,N_7,N_609);
nor U3557 (N_3557,N_1483,N_283);
or U3558 (N_3558,N_629,N_1128);
xor U3559 (N_3559,N_1619,N_1500);
nand U3560 (N_3560,N_1437,N_743);
and U3561 (N_3561,N_1553,N_1100);
xnor U3562 (N_3562,N_787,N_1902);
xor U3563 (N_3563,N_1800,N_1723);
or U3564 (N_3564,N_104,N_1222);
nand U3565 (N_3565,N_597,N_1077);
and U3566 (N_3566,N_1074,N_1226);
xnor U3567 (N_3567,N_1491,N_457);
nand U3568 (N_3568,N_995,N_1669);
nor U3569 (N_3569,N_776,N_1329);
nand U3570 (N_3570,N_141,N_1393);
or U3571 (N_3571,N_852,N_1367);
nand U3572 (N_3572,N_1433,N_868);
nand U3573 (N_3573,N_1057,N_878);
nand U3574 (N_3574,N_803,N_1488);
nor U3575 (N_3575,N_1309,N_877);
or U3576 (N_3576,N_1734,N_1839);
nand U3577 (N_3577,N_1552,N_1969);
nand U3578 (N_3578,N_512,N_142);
nor U3579 (N_3579,N_1686,N_1143);
xor U3580 (N_3580,N_391,N_313);
or U3581 (N_3581,N_422,N_672);
xor U3582 (N_3582,N_1826,N_1266);
nand U3583 (N_3583,N_1296,N_1788);
and U3584 (N_3584,N_1148,N_687);
and U3585 (N_3585,N_1715,N_1940);
or U3586 (N_3586,N_651,N_1497);
xor U3587 (N_3587,N_340,N_567);
xor U3588 (N_3588,N_1957,N_1522);
or U3589 (N_3589,N_1775,N_1196);
xor U3590 (N_3590,N_749,N_1858);
nor U3591 (N_3591,N_1351,N_1526);
or U3592 (N_3592,N_480,N_254);
nor U3593 (N_3593,N_1581,N_1305);
xnor U3594 (N_3594,N_1568,N_840);
and U3595 (N_3595,N_1702,N_240);
or U3596 (N_3596,N_317,N_1045);
or U3597 (N_3597,N_61,N_389);
and U3598 (N_3598,N_94,N_1856);
or U3599 (N_3599,N_744,N_1512);
and U3600 (N_3600,N_735,N_1509);
and U3601 (N_3601,N_1000,N_1939);
xnor U3602 (N_3602,N_1593,N_212);
and U3603 (N_3603,N_800,N_757);
nor U3604 (N_3604,N_280,N_919);
nor U3605 (N_3605,N_995,N_1488);
and U3606 (N_3606,N_1357,N_1435);
nor U3607 (N_3607,N_332,N_455);
or U3608 (N_3608,N_1520,N_1439);
nand U3609 (N_3609,N_1565,N_4);
nand U3610 (N_3610,N_190,N_1704);
and U3611 (N_3611,N_633,N_933);
nor U3612 (N_3612,N_475,N_1147);
nor U3613 (N_3613,N_133,N_1050);
or U3614 (N_3614,N_307,N_1773);
xnor U3615 (N_3615,N_531,N_752);
and U3616 (N_3616,N_1546,N_524);
nor U3617 (N_3617,N_426,N_485);
or U3618 (N_3618,N_1862,N_1574);
xnor U3619 (N_3619,N_1708,N_779);
xor U3620 (N_3620,N_477,N_302);
xor U3621 (N_3621,N_507,N_1566);
or U3622 (N_3622,N_189,N_969);
and U3623 (N_3623,N_682,N_409);
or U3624 (N_3624,N_1,N_1428);
xnor U3625 (N_3625,N_1826,N_1401);
and U3626 (N_3626,N_1507,N_415);
or U3627 (N_3627,N_428,N_527);
xor U3628 (N_3628,N_1084,N_786);
nor U3629 (N_3629,N_1548,N_380);
nand U3630 (N_3630,N_763,N_1718);
and U3631 (N_3631,N_1410,N_1825);
or U3632 (N_3632,N_1808,N_1285);
nand U3633 (N_3633,N_1987,N_1114);
nor U3634 (N_3634,N_711,N_1168);
nor U3635 (N_3635,N_824,N_1706);
and U3636 (N_3636,N_1640,N_547);
nand U3637 (N_3637,N_94,N_1460);
nand U3638 (N_3638,N_698,N_1544);
xnor U3639 (N_3639,N_941,N_1911);
xor U3640 (N_3640,N_459,N_1436);
or U3641 (N_3641,N_1555,N_1424);
nor U3642 (N_3642,N_840,N_954);
nor U3643 (N_3643,N_411,N_1422);
nand U3644 (N_3644,N_400,N_347);
and U3645 (N_3645,N_1803,N_741);
and U3646 (N_3646,N_1948,N_1508);
and U3647 (N_3647,N_218,N_925);
xnor U3648 (N_3648,N_977,N_1180);
xor U3649 (N_3649,N_95,N_1933);
xnor U3650 (N_3650,N_1525,N_561);
nor U3651 (N_3651,N_1866,N_1791);
xnor U3652 (N_3652,N_233,N_46);
nor U3653 (N_3653,N_71,N_518);
nand U3654 (N_3654,N_63,N_441);
and U3655 (N_3655,N_819,N_1150);
nor U3656 (N_3656,N_1210,N_441);
and U3657 (N_3657,N_1143,N_1937);
or U3658 (N_3658,N_1716,N_1851);
nand U3659 (N_3659,N_1757,N_575);
or U3660 (N_3660,N_1115,N_1157);
nand U3661 (N_3661,N_1136,N_1955);
or U3662 (N_3662,N_154,N_1050);
or U3663 (N_3663,N_1752,N_1770);
nor U3664 (N_3664,N_1133,N_1719);
nand U3665 (N_3665,N_1588,N_1263);
nor U3666 (N_3666,N_701,N_925);
xor U3667 (N_3667,N_1436,N_961);
and U3668 (N_3668,N_459,N_1468);
nand U3669 (N_3669,N_374,N_441);
nor U3670 (N_3670,N_209,N_317);
and U3671 (N_3671,N_1876,N_726);
nand U3672 (N_3672,N_1212,N_1485);
or U3673 (N_3673,N_1028,N_724);
nor U3674 (N_3674,N_1523,N_1507);
nor U3675 (N_3675,N_504,N_1934);
nand U3676 (N_3676,N_1234,N_1918);
and U3677 (N_3677,N_657,N_731);
nor U3678 (N_3678,N_1061,N_1206);
and U3679 (N_3679,N_1951,N_1733);
and U3680 (N_3680,N_809,N_540);
nand U3681 (N_3681,N_1336,N_1279);
nand U3682 (N_3682,N_1751,N_1974);
xor U3683 (N_3683,N_139,N_613);
xnor U3684 (N_3684,N_771,N_498);
or U3685 (N_3685,N_448,N_488);
nand U3686 (N_3686,N_628,N_1007);
nor U3687 (N_3687,N_1286,N_1054);
nand U3688 (N_3688,N_749,N_1323);
and U3689 (N_3689,N_488,N_14);
nand U3690 (N_3690,N_1284,N_1435);
xnor U3691 (N_3691,N_188,N_1274);
and U3692 (N_3692,N_740,N_1220);
nor U3693 (N_3693,N_1159,N_526);
xor U3694 (N_3694,N_760,N_426);
and U3695 (N_3695,N_1636,N_670);
nand U3696 (N_3696,N_662,N_137);
nor U3697 (N_3697,N_1417,N_1524);
xor U3698 (N_3698,N_519,N_97);
nand U3699 (N_3699,N_112,N_1004);
nor U3700 (N_3700,N_1454,N_1337);
or U3701 (N_3701,N_411,N_1047);
nor U3702 (N_3702,N_1796,N_1033);
nor U3703 (N_3703,N_1161,N_1304);
nand U3704 (N_3704,N_840,N_656);
or U3705 (N_3705,N_1519,N_1204);
nor U3706 (N_3706,N_8,N_660);
xor U3707 (N_3707,N_1070,N_1291);
nor U3708 (N_3708,N_281,N_736);
xor U3709 (N_3709,N_738,N_1697);
and U3710 (N_3710,N_754,N_866);
nand U3711 (N_3711,N_1974,N_574);
and U3712 (N_3712,N_1350,N_281);
and U3713 (N_3713,N_1014,N_1277);
nand U3714 (N_3714,N_1246,N_244);
or U3715 (N_3715,N_1975,N_1070);
or U3716 (N_3716,N_1011,N_244);
xor U3717 (N_3717,N_1811,N_1673);
xnor U3718 (N_3718,N_863,N_302);
xor U3719 (N_3719,N_1224,N_979);
nand U3720 (N_3720,N_1126,N_388);
xnor U3721 (N_3721,N_1487,N_894);
nor U3722 (N_3722,N_186,N_1408);
and U3723 (N_3723,N_1783,N_330);
nand U3724 (N_3724,N_279,N_1344);
nand U3725 (N_3725,N_103,N_820);
and U3726 (N_3726,N_504,N_814);
nor U3727 (N_3727,N_374,N_769);
or U3728 (N_3728,N_1134,N_1323);
nor U3729 (N_3729,N_712,N_1950);
and U3730 (N_3730,N_737,N_1094);
xor U3731 (N_3731,N_110,N_435);
nor U3732 (N_3732,N_149,N_377);
nor U3733 (N_3733,N_851,N_882);
and U3734 (N_3734,N_501,N_1576);
or U3735 (N_3735,N_923,N_995);
nor U3736 (N_3736,N_524,N_139);
and U3737 (N_3737,N_1301,N_1958);
and U3738 (N_3738,N_1404,N_1421);
or U3739 (N_3739,N_1722,N_243);
and U3740 (N_3740,N_1171,N_677);
nand U3741 (N_3741,N_1560,N_1505);
or U3742 (N_3742,N_1635,N_1054);
nor U3743 (N_3743,N_800,N_16);
nor U3744 (N_3744,N_77,N_1909);
xor U3745 (N_3745,N_1108,N_24);
nand U3746 (N_3746,N_93,N_56);
nor U3747 (N_3747,N_1852,N_564);
nor U3748 (N_3748,N_927,N_1925);
or U3749 (N_3749,N_1709,N_1618);
nand U3750 (N_3750,N_489,N_436);
xnor U3751 (N_3751,N_1397,N_652);
nand U3752 (N_3752,N_1240,N_670);
and U3753 (N_3753,N_97,N_1307);
nand U3754 (N_3754,N_532,N_601);
and U3755 (N_3755,N_983,N_1019);
nand U3756 (N_3756,N_999,N_1176);
nor U3757 (N_3757,N_768,N_40);
nor U3758 (N_3758,N_649,N_407);
and U3759 (N_3759,N_1441,N_682);
xnor U3760 (N_3760,N_1820,N_1274);
and U3761 (N_3761,N_266,N_382);
nand U3762 (N_3762,N_1424,N_1627);
and U3763 (N_3763,N_1987,N_1391);
nor U3764 (N_3764,N_149,N_1151);
or U3765 (N_3765,N_4,N_1716);
and U3766 (N_3766,N_868,N_1378);
xor U3767 (N_3767,N_1244,N_669);
xnor U3768 (N_3768,N_642,N_1775);
or U3769 (N_3769,N_747,N_1312);
nor U3770 (N_3770,N_1098,N_1317);
xnor U3771 (N_3771,N_1877,N_1306);
xor U3772 (N_3772,N_1180,N_269);
nand U3773 (N_3773,N_373,N_458);
and U3774 (N_3774,N_180,N_1294);
or U3775 (N_3775,N_753,N_361);
nand U3776 (N_3776,N_290,N_278);
xor U3777 (N_3777,N_54,N_370);
nand U3778 (N_3778,N_1022,N_1104);
or U3779 (N_3779,N_1047,N_127);
or U3780 (N_3780,N_141,N_1781);
or U3781 (N_3781,N_1155,N_1372);
or U3782 (N_3782,N_1646,N_1856);
nand U3783 (N_3783,N_395,N_367);
nand U3784 (N_3784,N_1085,N_1021);
nor U3785 (N_3785,N_1546,N_673);
and U3786 (N_3786,N_1587,N_1012);
nor U3787 (N_3787,N_924,N_1303);
or U3788 (N_3788,N_325,N_1158);
or U3789 (N_3789,N_1343,N_1360);
and U3790 (N_3790,N_797,N_1237);
nor U3791 (N_3791,N_745,N_1603);
xnor U3792 (N_3792,N_1194,N_837);
xnor U3793 (N_3793,N_52,N_1338);
nor U3794 (N_3794,N_1175,N_1631);
and U3795 (N_3795,N_1542,N_856);
nand U3796 (N_3796,N_1393,N_64);
xnor U3797 (N_3797,N_202,N_1282);
and U3798 (N_3798,N_182,N_1256);
nor U3799 (N_3799,N_1638,N_1470);
nand U3800 (N_3800,N_989,N_1356);
nor U3801 (N_3801,N_1387,N_425);
nand U3802 (N_3802,N_1553,N_1777);
nand U3803 (N_3803,N_1337,N_742);
xor U3804 (N_3804,N_1584,N_912);
xor U3805 (N_3805,N_1633,N_1804);
and U3806 (N_3806,N_783,N_1415);
or U3807 (N_3807,N_1906,N_1856);
xor U3808 (N_3808,N_572,N_1305);
xnor U3809 (N_3809,N_60,N_153);
nor U3810 (N_3810,N_423,N_1784);
and U3811 (N_3811,N_110,N_50);
and U3812 (N_3812,N_1665,N_514);
and U3813 (N_3813,N_30,N_1754);
nand U3814 (N_3814,N_1450,N_456);
xor U3815 (N_3815,N_1209,N_1690);
and U3816 (N_3816,N_1245,N_1894);
or U3817 (N_3817,N_368,N_1821);
xor U3818 (N_3818,N_666,N_1246);
and U3819 (N_3819,N_137,N_1583);
and U3820 (N_3820,N_850,N_1587);
nand U3821 (N_3821,N_737,N_1233);
nor U3822 (N_3822,N_1073,N_412);
nand U3823 (N_3823,N_1323,N_1646);
xor U3824 (N_3824,N_583,N_210);
and U3825 (N_3825,N_982,N_830);
nor U3826 (N_3826,N_1667,N_177);
nor U3827 (N_3827,N_1194,N_235);
nor U3828 (N_3828,N_1176,N_1703);
nand U3829 (N_3829,N_1445,N_678);
nor U3830 (N_3830,N_4,N_665);
or U3831 (N_3831,N_1304,N_814);
or U3832 (N_3832,N_153,N_1347);
and U3833 (N_3833,N_206,N_962);
nor U3834 (N_3834,N_42,N_1070);
nor U3835 (N_3835,N_1597,N_1177);
nor U3836 (N_3836,N_304,N_518);
nand U3837 (N_3837,N_1316,N_1887);
nand U3838 (N_3838,N_1500,N_168);
xor U3839 (N_3839,N_1568,N_617);
or U3840 (N_3840,N_1307,N_614);
nor U3841 (N_3841,N_783,N_868);
nor U3842 (N_3842,N_710,N_217);
and U3843 (N_3843,N_1577,N_1132);
or U3844 (N_3844,N_1283,N_1778);
and U3845 (N_3845,N_1279,N_1870);
nand U3846 (N_3846,N_1571,N_907);
xor U3847 (N_3847,N_994,N_112);
nor U3848 (N_3848,N_335,N_156);
xor U3849 (N_3849,N_1087,N_1795);
nand U3850 (N_3850,N_234,N_614);
nor U3851 (N_3851,N_777,N_1297);
nand U3852 (N_3852,N_860,N_1402);
or U3853 (N_3853,N_832,N_1581);
xnor U3854 (N_3854,N_1409,N_560);
nand U3855 (N_3855,N_1993,N_742);
nand U3856 (N_3856,N_4,N_751);
nand U3857 (N_3857,N_564,N_1833);
nor U3858 (N_3858,N_1729,N_1302);
or U3859 (N_3859,N_1196,N_552);
nand U3860 (N_3860,N_1217,N_594);
nor U3861 (N_3861,N_540,N_1259);
xor U3862 (N_3862,N_1584,N_1681);
xor U3863 (N_3863,N_863,N_1501);
nand U3864 (N_3864,N_1458,N_1796);
nand U3865 (N_3865,N_21,N_1881);
nor U3866 (N_3866,N_293,N_859);
nand U3867 (N_3867,N_1198,N_569);
xnor U3868 (N_3868,N_890,N_944);
xor U3869 (N_3869,N_754,N_409);
and U3870 (N_3870,N_1599,N_1580);
or U3871 (N_3871,N_188,N_1909);
or U3872 (N_3872,N_56,N_273);
nor U3873 (N_3873,N_1545,N_1124);
and U3874 (N_3874,N_1880,N_1305);
xnor U3875 (N_3875,N_454,N_1413);
and U3876 (N_3876,N_185,N_638);
xor U3877 (N_3877,N_1773,N_754);
and U3878 (N_3878,N_921,N_413);
nand U3879 (N_3879,N_1179,N_1541);
nand U3880 (N_3880,N_1464,N_457);
xor U3881 (N_3881,N_1649,N_1797);
and U3882 (N_3882,N_683,N_277);
or U3883 (N_3883,N_880,N_1263);
and U3884 (N_3884,N_451,N_683);
or U3885 (N_3885,N_492,N_494);
or U3886 (N_3886,N_911,N_1621);
xor U3887 (N_3887,N_824,N_304);
nand U3888 (N_3888,N_401,N_1209);
nand U3889 (N_3889,N_1704,N_786);
nor U3890 (N_3890,N_494,N_1346);
xor U3891 (N_3891,N_1424,N_199);
and U3892 (N_3892,N_1002,N_1613);
nand U3893 (N_3893,N_627,N_1985);
xor U3894 (N_3894,N_501,N_809);
nor U3895 (N_3895,N_450,N_1338);
nor U3896 (N_3896,N_1882,N_586);
nor U3897 (N_3897,N_1773,N_1078);
or U3898 (N_3898,N_747,N_1506);
nand U3899 (N_3899,N_824,N_1448);
or U3900 (N_3900,N_853,N_152);
xnor U3901 (N_3901,N_1455,N_600);
and U3902 (N_3902,N_1051,N_420);
or U3903 (N_3903,N_851,N_1975);
xor U3904 (N_3904,N_1181,N_1362);
nor U3905 (N_3905,N_1398,N_960);
nand U3906 (N_3906,N_1350,N_251);
nand U3907 (N_3907,N_1709,N_50);
and U3908 (N_3908,N_81,N_528);
or U3909 (N_3909,N_239,N_624);
nand U3910 (N_3910,N_684,N_1706);
and U3911 (N_3911,N_1192,N_1715);
xor U3912 (N_3912,N_1037,N_1430);
nand U3913 (N_3913,N_947,N_1752);
nand U3914 (N_3914,N_1469,N_1479);
or U3915 (N_3915,N_1224,N_888);
nor U3916 (N_3916,N_201,N_1591);
nor U3917 (N_3917,N_909,N_735);
nand U3918 (N_3918,N_548,N_257);
nand U3919 (N_3919,N_496,N_534);
xor U3920 (N_3920,N_416,N_412);
nor U3921 (N_3921,N_1056,N_837);
and U3922 (N_3922,N_1253,N_1112);
nand U3923 (N_3923,N_1699,N_467);
xnor U3924 (N_3924,N_36,N_229);
xor U3925 (N_3925,N_1894,N_477);
nor U3926 (N_3926,N_65,N_1300);
nor U3927 (N_3927,N_847,N_1564);
or U3928 (N_3928,N_1908,N_452);
nand U3929 (N_3929,N_888,N_446);
and U3930 (N_3930,N_1044,N_247);
nor U3931 (N_3931,N_1409,N_118);
or U3932 (N_3932,N_678,N_965);
or U3933 (N_3933,N_1531,N_1989);
xnor U3934 (N_3934,N_200,N_1978);
or U3935 (N_3935,N_1258,N_152);
xor U3936 (N_3936,N_1850,N_693);
xor U3937 (N_3937,N_1572,N_1143);
and U3938 (N_3938,N_1396,N_352);
xnor U3939 (N_3939,N_1036,N_1730);
nand U3940 (N_3940,N_1123,N_1786);
xnor U3941 (N_3941,N_359,N_1246);
xor U3942 (N_3942,N_119,N_1105);
nand U3943 (N_3943,N_762,N_281);
or U3944 (N_3944,N_403,N_1623);
nand U3945 (N_3945,N_703,N_272);
nor U3946 (N_3946,N_1077,N_1496);
nor U3947 (N_3947,N_1996,N_1018);
xor U3948 (N_3948,N_334,N_1904);
and U3949 (N_3949,N_115,N_1799);
or U3950 (N_3950,N_835,N_1190);
or U3951 (N_3951,N_1073,N_1833);
nor U3952 (N_3952,N_558,N_1690);
or U3953 (N_3953,N_47,N_1964);
and U3954 (N_3954,N_703,N_1030);
xnor U3955 (N_3955,N_406,N_1180);
and U3956 (N_3956,N_603,N_1794);
or U3957 (N_3957,N_469,N_884);
and U3958 (N_3958,N_253,N_1052);
xor U3959 (N_3959,N_1507,N_226);
xnor U3960 (N_3960,N_1856,N_668);
or U3961 (N_3961,N_1510,N_285);
nor U3962 (N_3962,N_93,N_1086);
nor U3963 (N_3963,N_1074,N_274);
or U3964 (N_3964,N_1110,N_148);
xnor U3965 (N_3965,N_1052,N_413);
or U3966 (N_3966,N_78,N_61);
nor U3967 (N_3967,N_833,N_1449);
or U3968 (N_3968,N_898,N_456);
or U3969 (N_3969,N_1597,N_548);
and U3970 (N_3970,N_1581,N_654);
or U3971 (N_3971,N_1516,N_3);
or U3972 (N_3972,N_394,N_1597);
xnor U3973 (N_3973,N_276,N_1747);
nand U3974 (N_3974,N_857,N_1837);
xor U3975 (N_3975,N_202,N_1527);
nor U3976 (N_3976,N_621,N_1664);
nor U3977 (N_3977,N_210,N_266);
and U3978 (N_3978,N_1624,N_1633);
xnor U3979 (N_3979,N_140,N_549);
nor U3980 (N_3980,N_707,N_1468);
nor U3981 (N_3981,N_1288,N_2);
nor U3982 (N_3982,N_644,N_846);
nor U3983 (N_3983,N_1867,N_959);
xor U3984 (N_3984,N_1411,N_546);
nor U3985 (N_3985,N_1081,N_1092);
or U3986 (N_3986,N_1035,N_1270);
nor U3987 (N_3987,N_1574,N_1390);
nand U3988 (N_3988,N_1379,N_1691);
or U3989 (N_3989,N_599,N_1272);
nor U3990 (N_3990,N_524,N_1486);
nand U3991 (N_3991,N_1584,N_0);
or U3992 (N_3992,N_750,N_342);
and U3993 (N_3993,N_854,N_939);
nor U3994 (N_3994,N_1349,N_88);
and U3995 (N_3995,N_1474,N_805);
or U3996 (N_3996,N_1434,N_167);
nand U3997 (N_3997,N_825,N_79);
nor U3998 (N_3998,N_1567,N_1565);
nand U3999 (N_3999,N_923,N_753);
or U4000 (N_4000,N_3964,N_3809);
nor U4001 (N_4001,N_2800,N_2880);
nor U4002 (N_4002,N_3887,N_3422);
nor U4003 (N_4003,N_2543,N_2284);
xor U4004 (N_4004,N_2468,N_3638);
nand U4005 (N_4005,N_2405,N_3859);
nand U4006 (N_4006,N_3173,N_3883);
nor U4007 (N_4007,N_3433,N_3895);
xnor U4008 (N_4008,N_2045,N_2644);
nand U4009 (N_4009,N_3866,N_3586);
nor U4010 (N_4010,N_2229,N_3450);
nand U4011 (N_4011,N_2752,N_3099);
nand U4012 (N_4012,N_3588,N_3216);
or U4013 (N_4013,N_2399,N_2690);
nand U4014 (N_4014,N_3855,N_3485);
nand U4015 (N_4015,N_2595,N_3940);
or U4016 (N_4016,N_3750,N_2280);
and U4017 (N_4017,N_3868,N_3147);
xnor U4018 (N_4018,N_2908,N_3221);
xnor U4019 (N_4019,N_3058,N_3315);
nor U4020 (N_4020,N_3772,N_3881);
or U4021 (N_4021,N_2387,N_2286);
nand U4022 (N_4022,N_2683,N_2178);
xnor U4023 (N_4023,N_3299,N_3959);
xor U4024 (N_4024,N_3548,N_3040);
nor U4025 (N_4025,N_2710,N_3573);
or U4026 (N_4026,N_3563,N_2645);
nor U4027 (N_4027,N_2240,N_2343);
nor U4028 (N_4028,N_3191,N_2790);
or U4029 (N_4029,N_2635,N_3897);
and U4030 (N_4030,N_3672,N_2599);
nand U4031 (N_4031,N_3472,N_3441);
xor U4032 (N_4032,N_2364,N_2504);
xor U4033 (N_4033,N_3415,N_3296);
xnor U4034 (N_4034,N_3062,N_2545);
or U4035 (N_4035,N_3832,N_2228);
nand U4036 (N_4036,N_3131,N_2214);
nor U4037 (N_4037,N_3574,N_2632);
and U4038 (N_4038,N_2384,N_2059);
and U4039 (N_4039,N_3107,N_2922);
and U4040 (N_4040,N_2893,N_2902);
or U4041 (N_4041,N_3014,N_3564);
and U4042 (N_4042,N_3187,N_3265);
nand U4043 (N_4043,N_3506,N_3053);
or U4044 (N_4044,N_2702,N_2986);
nand U4045 (N_4045,N_3807,N_3322);
or U4046 (N_4046,N_3406,N_3145);
xor U4047 (N_4047,N_3434,N_2762);
or U4048 (N_4048,N_3353,N_2032);
nand U4049 (N_4049,N_3876,N_3211);
xnor U4050 (N_4050,N_3411,N_2082);
or U4051 (N_4051,N_2777,N_2782);
nor U4052 (N_4052,N_3421,N_3346);
or U4053 (N_4053,N_3646,N_3015);
nand U4054 (N_4054,N_3439,N_2989);
or U4055 (N_4055,N_3596,N_2218);
nand U4056 (N_4056,N_2542,N_2518);
and U4057 (N_4057,N_3337,N_3529);
and U4058 (N_4058,N_2708,N_3267);
nand U4059 (N_4059,N_3047,N_3643);
or U4060 (N_4060,N_3510,N_2401);
or U4061 (N_4061,N_2612,N_3177);
or U4062 (N_4062,N_2493,N_3320);
xor U4063 (N_4063,N_3373,N_3290);
nor U4064 (N_4064,N_2431,N_3579);
xnor U4065 (N_4065,N_3598,N_2927);
nor U4066 (N_4066,N_2968,N_3377);
nand U4067 (N_4067,N_2135,N_3929);
nand U4068 (N_4068,N_2763,N_2066);
nor U4069 (N_4069,N_2418,N_3117);
or U4070 (N_4070,N_2014,N_2039);
nor U4071 (N_4071,N_3936,N_3307);
nand U4072 (N_4072,N_3224,N_2962);
xnor U4073 (N_4073,N_2126,N_2550);
nand U4074 (N_4074,N_2540,N_2507);
nand U4075 (N_4075,N_2909,N_3631);
nand U4076 (N_4076,N_3995,N_2144);
xor U4077 (N_4077,N_3871,N_2532);
nand U4078 (N_4078,N_2636,N_3258);
and U4079 (N_4079,N_2743,N_2512);
or U4080 (N_4080,N_3851,N_2237);
nor U4081 (N_4081,N_3557,N_2815);
nor U4082 (N_4082,N_3097,N_3526);
nand U4083 (N_4083,N_3812,N_3697);
xor U4084 (N_4084,N_2951,N_2696);
nand U4085 (N_4085,N_2328,N_2633);
nor U4086 (N_4086,N_2967,N_2332);
nor U4087 (N_4087,N_2466,N_2460);
nand U4088 (N_4088,N_2094,N_3449);
nor U4089 (N_4089,N_2368,N_3416);
and U4090 (N_4090,N_2206,N_2067);
nand U4091 (N_4091,N_3059,N_3440);
and U4092 (N_4092,N_3533,N_3055);
or U4093 (N_4093,N_3930,N_3487);
xor U4094 (N_4094,N_2324,N_2615);
or U4095 (N_4095,N_2695,N_2792);
nand U4096 (N_4096,N_2073,N_2728);
and U4097 (N_4097,N_2721,N_2692);
nand U4098 (N_4098,N_3298,N_2597);
nand U4099 (N_4099,N_2724,N_2485);
and U4100 (N_4100,N_2143,N_3823);
or U4101 (N_4101,N_3486,N_3051);
xnor U4102 (N_4102,N_3309,N_2783);
or U4103 (N_4103,N_3981,N_3539);
xnor U4104 (N_4104,N_2230,N_3917);
nor U4105 (N_4105,N_3752,N_3410);
nor U4106 (N_4106,N_2440,N_3644);
and U4107 (N_4107,N_3189,N_3854);
and U4108 (N_4108,N_3786,N_3122);
xnor U4109 (N_4109,N_3597,N_3233);
and U4110 (N_4110,N_3822,N_2247);
or U4111 (N_4111,N_2348,N_3350);
or U4112 (N_4112,N_2575,N_2382);
nand U4113 (N_4113,N_2506,N_2513);
nand U4114 (N_4114,N_2347,N_3060);
and U4115 (N_4115,N_3057,N_2491);
xnor U4116 (N_4116,N_2906,N_3042);
nor U4117 (N_4117,N_2374,N_3085);
or U4118 (N_4118,N_2156,N_2040);
nand U4119 (N_4119,N_2765,N_2873);
or U4120 (N_4120,N_3061,N_2445);
nand U4121 (N_4121,N_3242,N_3474);
xor U4122 (N_4122,N_3056,N_2317);
nor U4123 (N_4123,N_2235,N_3630);
nor U4124 (N_4124,N_2806,N_2589);
xor U4125 (N_4125,N_2684,N_3845);
nor U4126 (N_4126,N_2494,N_2961);
nand U4127 (N_4127,N_2823,N_2581);
nor U4128 (N_4128,N_2946,N_3074);
nand U4129 (N_4129,N_3431,N_3448);
nor U4130 (N_4130,N_2409,N_2876);
or U4131 (N_4131,N_3957,N_3517);
nor U4132 (N_4132,N_2365,N_3490);
or U4133 (N_4133,N_3717,N_2312);
or U4134 (N_4134,N_2606,N_3384);
xnor U4135 (N_4135,N_3654,N_3674);
and U4136 (N_4136,N_3266,N_2878);
nand U4137 (N_4137,N_3587,N_2520);
nand U4138 (N_4138,N_2147,N_2809);
and U4139 (N_4139,N_3788,N_3864);
nor U4140 (N_4140,N_2301,N_3158);
nor U4141 (N_4141,N_2691,N_3162);
or U4142 (N_4142,N_3756,N_2252);
or U4143 (N_4143,N_2323,N_3423);
and U4144 (N_4144,N_2386,N_3225);
or U4145 (N_4145,N_3865,N_3974);
and U4146 (N_4146,N_3137,N_3836);
xnor U4147 (N_4147,N_3240,N_3558);
xor U4148 (N_4148,N_2410,N_2510);
or U4149 (N_4149,N_2569,N_3824);
and U4150 (N_4150,N_2734,N_3483);
xor U4151 (N_4151,N_3444,N_2924);
nand U4152 (N_4152,N_2579,N_3797);
and U4153 (N_4153,N_3541,N_2226);
or U4154 (N_4154,N_3043,N_2225);
xnor U4155 (N_4155,N_2331,N_2795);
nor U4156 (N_4156,N_3291,N_3889);
xor U4157 (N_4157,N_2617,N_2356);
nand U4158 (N_4158,N_2803,N_3610);
or U4159 (N_4159,N_2796,N_2694);
nand U4160 (N_4160,N_3721,N_3341);
xor U4161 (N_4161,N_2498,N_3363);
or U4162 (N_4162,N_3723,N_3479);
nor U4163 (N_4163,N_3451,N_3905);
xor U4164 (N_4164,N_3808,N_3627);
and U4165 (N_4165,N_2448,N_3700);
and U4166 (N_4166,N_2013,N_3943);
and U4167 (N_4167,N_3725,N_2716);
and U4168 (N_4168,N_3910,N_2840);
nand U4169 (N_4169,N_3869,N_2404);
xor U4170 (N_4170,N_3716,N_2231);
nand U4171 (N_4171,N_3387,N_2462);
and U4172 (N_4172,N_3289,N_3821);
xnor U4173 (N_4173,N_2490,N_2105);
xor U4174 (N_4174,N_2098,N_3877);
or U4175 (N_4175,N_3727,N_3075);
nand U4176 (N_4176,N_3664,N_3844);
or U4177 (N_4177,N_3209,N_3914);
xnor U4178 (N_4178,N_2239,N_2487);
nand U4179 (N_4179,N_2836,N_2799);
and U4180 (N_4180,N_3963,N_3382);
and U4181 (N_4181,N_3626,N_2559);
nand U4182 (N_4182,N_3934,N_2903);
or U4183 (N_4183,N_2434,N_3773);
or U4184 (N_4184,N_2288,N_3501);
xnor U4185 (N_4185,N_2877,N_3293);
or U4186 (N_4186,N_3436,N_2667);
nand U4187 (N_4187,N_2580,N_3571);
nand U4188 (N_4188,N_3554,N_3068);
nor U4189 (N_4189,N_3566,N_2276);
xnor U4190 (N_4190,N_2134,N_2771);
xor U4191 (N_4191,N_3530,N_2154);
nor U4192 (N_4192,N_2890,N_3915);
or U4193 (N_4193,N_3193,N_3560);
and U4194 (N_4194,N_2707,N_3657);
nand U4195 (N_4195,N_2954,N_3755);
or U4196 (N_4196,N_2748,N_3276);
nor U4197 (N_4197,N_2307,N_2124);
nand U4198 (N_4198,N_2330,N_2205);
xnor U4199 (N_4199,N_3249,N_2200);
nand U4200 (N_4200,N_2037,N_3527);
xor U4201 (N_4201,N_2339,N_2030);
nor U4202 (N_4202,N_3295,N_2333);
xor U4203 (N_4203,N_3710,N_2236);
nor U4204 (N_4204,N_2981,N_2793);
and U4205 (N_4205,N_2839,N_2122);
or U4206 (N_4206,N_2592,N_3323);
nor U4207 (N_4207,N_3691,N_3453);
nor U4208 (N_4208,N_3690,N_2619);
and U4209 (N_4209,N_2607,N_2990);
or U4210 (N_4210,N_2004,N_3803);
xor U4211 (N_4211,N_3509,N_2081);
or U4212 (N_4212,N_2196,N_3665);
or U4213 (N_4213,N_2290,N_3528);
and U4214 (N_4214,N_3310,N_3802);
nor U4215 (N_4215,N_2647,N_2515);
nor U4216 (N_4216,N_3104,N_2233);
or U4217 (N_4217,N_3467,N_3352);
nor U4218 (N_4218,N_2892,N_3857);
or U4219 (N_4219,N_3362,N_2417);
nand U4220 (N_4220,N_3684,N_2860);
or U4221 (N_4221,N_3961,N_3994);
nand U4222 (N_4222,N_3706,N_2602);
and U4223 (N_4223,N_3123,N_2623);
xnor U4224 (N_4224,N_3159,N_2801);
or U4225 (N_4225,N_3072,N_2408);
nand U4226 (N_4226,N_2258,N_3282);
xnor U4227 (N_4227,N_2705,N_2208);
and U4228 (N_4228,N_3306,N_2488);
xnor U4229 (N_4229,N_3985,N_2654);
or U4230 (N_4230,N_2704,N_3944);
nand U4231 (N_4231,N_2565,N_3863);
or U4232 (N_4232,N_2215,N_2243);
or U4233 (N_4233,N_3918,N_3157);
nor U4234 (N_4234,N_3988,N_3408);
nand U4235 (N_4235,N_3738,N_3703);
nand U4236 (N_4236,N_3124,N_2452);
xor U4237 (N_4237,N_3962,N_2107);
and U4238 (N_4238,N_2574,N_3789);
nand U4239 (N_4239,N_2216,N_3760);
nand U4240 (N_4240,N_2874,N_2531);
xnor U4241 (N_4241,N_3933,N_2920);
or U4242 (N_4242,N_2601,N_3022);
nand U4243 (N_4243,N_3555,N_3997);
and U4244 (N_4244,N_2241,N_2202);
and U4245 (N_4245,N_2807,N_3188);
xnor U4246 (N_4246,N_2572,N_3183);
nor U4247 (N_4247,N_2198,N_3935);
nand U4248 (N_4248,N_2779,N_3196);
and U4249 (N_4249,N_2457,N_2455);
or U4250 (N_4250,N_2766,N_2184);
nand U4251 (N_4251,N_2665,N_2311);
nand U4252 (N_4252,N_3696,N_3271);
or U4253 (N_4253,N_3184,N_2213);
xnor U4254 (N_4254,N_3503,N_2744);
nor U4255 (N_4255,N_3326,N_2825);
xnor U4256 (N_4256,N_3305,N_3941);
nand U4257 (N_4257,N_3837,N_3493);
nand U4258 (N_4258,N_3420,N_2308);
and U4259 (N_4259,N_2188,N_3340);
nor U4260 (N_4260,N_2473,N_2091);
nor U4261 (N_4261,N_3185,N_2291);
nor U4262 (N_4262,N_3312,N_2313);
xnor U4263 (N_4263,N_3460,N_3227);
or U4264 (N_4264,N_2933,N_2772);
or U4265 (N_4265,N_2223,N_2958);
nand U4266 (N_4266,N_3149,N_2011);
nor U4267 (N_4267,N_3237,N_3795);
nor U4268 (N_4268,N_3693,N_2381);
xnor U4269 (N_4269,N_3039,N_3512);
nor U4270 (N_4270,N_2594,N_3300);
or U4271 (N_4271,N_2677,N_2372);
or U4272 (N_4272,N_2857,N_2084);
and U4273 (N_4273,N_3426,N_3902);
nor U4274 (N_4274,N_3076,N_2537);
xnor U4275 (N_4275,N_2598,N_3459);
xnor U4276 (N_4276,N_2912,N_3798);
nand U4277 (N_4277,N_2578,N_3391);
nand U4278 (N_4278,N_2412,N_2556);
or U4279 (N_4279,N_2177,N_2337);
or U4280 (N_4280,N_3470,N_2376);
and U4281 (N_4281,N_3109,N_2056);
and U4282 (N_4282,N_2370,N_2345);
or U4283 (N_4283,N_3916,N_3089);
and U4284 (N_4284,N_3656,N_3390);
nor U4285 (N_4285,N_2207,N_2027);
nand U4286 (N_4286,N_3017,N_2309);
nor U4287 (N_4287,N_3165,N_2971);
nand U4288 (N_4288,N_2630,N_2437);
nor U4289 (N_4289,N_3427,N_2586);
or U4290 (N_4290,N_3600,N_2593);
xnor U4291 (N_4291,N_2625,N_2979);
nand U4292 (N_4292,N_2145,N_3395);
nand U4293 (N_4293,N_2141,N_3906);
nand U4294 (N_4294,N_3903,N_2670);
nand U4295 (N_4295,N_3519,N_3218);
or U4296 (N_4296,N_2173,N_2052);
and U4297 (N_4297,N_3617,N_3719);
nand U4298 (N_4298,N_3791,N_2300);
nand U4299 (N_4299,N_3658,N_3378);
nand U4300 (N_4300,N_2170,N_2031);
nor U4301 (N_4301,N_3160,N_3524);
nor U4302 (N_4302,N_3088,N_2770);
xnor U4303 (N_4303,N_3394,N_3778);
or U4304 (N_4304,N_2957,N_2151);
nor U4305 (N_4305,N_2541,N_2273);
nor U4306 (N_4306,N_2747,N_2183);
nor U4307 (N_4307,N_2383,N_3200);
nor U4308 (N_4308,N_2042,N_2904);
or U4309 (N_4309,N_3376,N_3686);
and U4310 (N_4310,N_2109,N_3615);
xnor U4311 (N_4311,N_3250,N_2563);
and U4312 (N_4312,N_3967,N_2193);
and U4313 (N_4313,N_3311,N_3278);
nand U4314 (N_4314,N_2994,N_3284);
xnor U4315 (N_4315,N_2767,N_3956);
xor U4316 (N_4316,N_3682,N_2919);
or U4317 (N_4317,N_2731,N_2378);
xor U4318 (N_4318,N_2316,N_3446);
or U4319 (N_4319,N_3833,N_2433);
and U4320 (N_4320,N_2834,N_3199);
nor U4321 (N_4321,N_3660,N_3318);
or U4322 (N_4322,N_3590,N_2069);
and U4323 (N_4323,N_2521,N_2864);
nor U4324 (N_4324,N_2481,N_3429);
or U4325 (N_4325,N_2289,N_3077);
xnor U4326 (N_4326,N_3201,N_3398);
nor U4327 (N_4327,N_2931,N_3100);
nor U4328 (N_4328,N_3513,N_2415);
xnor U4329 (N_4329,N_3603,N_3673);
and U4330 (N_4330,N_3167,N_2501);
or U4331 (N_4331,N_3946,N_3839);
xnor U4332 (N_4332,N_3210,N_2053);
or U4333 (N_4333,N_2190,N_3645);
nand U4334 (N_4334,N_3993,N_3805);
nand U4335 (N_4335,N_2071,N_2883);
and U4336 (N_4336,N_3958,N_2470);
or U4337 (N_4337,N_2192,N_2687);
xor U4338 (N_4338,N_2600,N_2535);
nor U4339 (N_4339,N_3980,N_3480);
nor U4340 (N_4340,N_2375,N_2717);
and U4341 (N_4341,N_2789,N_2090);
xor U4342 (N_4342,N_3843,N_2295);
xor U4343 (N_4343,N_3890,N_2078);
and U4344 (N_4344,N_2963,N_2640);
and U4345 (N_4345,N_2087,N_2675);
or U4346 (N_4346,N_3151,N_2167);
nand U4347 (N_4347,N_3360,N_3737);
or U4348 (N_4348,N_2005,N_3662);
nor U4349 (N_4349,N_2830,N_2355);
nand U4350 (N_4350,N_3749,N_3709);
nand U4351 (N_4351,N_2780,N_2499);
or U4352 (N_4352,N_2304,N_2018);
nand U4353 (N_4353,N_3784,N_2282);
or U4354 (N_4354,N_2422,N_2703);
nor U4355 (N_4355,N_3297,N_2523);
or U4356 (N_4356,N_2881,N_2660);
nand U4357 (N_4357,N_3019,N_3259);
nand U4358 (N_4358,N_2776,N_2576);
nand U4359 (N_4359,N_3983,N_2831);
nor U4360 (N_4360,N_3283,N_3425);
nand U4361 (N_4361,N_3150,N_3288);
xnor U4362 (N_4362,N_2588,N_3522);
nand U4363 (N_4363,N_3796,N_2441);
nor U4364 (N_4364,N_3153,N_3009);
nand U4365 (N_4365,N_3438,N_2753);
and U4366 (N_4366,N_2773,N_3888);
or U4367 (N_4367,N_3146,N_3948);
nand U4368 (N_4368,N_3071,N_2058);
nor U4369 (N_4369,N_3601,N_3751);
or U4370 (N_4370,N_2211,N_2938);
and U4371 (N_4371,N_2242,N_3951);
nor U4372 (N_4372,N_3713,N_2165);
nor U4373 (N_4373,N_3507,N_3163);
nand U4374 (N_4374,N_3239,N_2006);
nor U4375 (N_4375,N_3385,N_3031);
or U4376 (N_4376,N_2043,N_2508);
xor U4377 (N_4377,N_2658,N_3286);
nand U4378 (N_4378,N_2294,N_3867);
or U4379 (N_4379,N_3591,N_2794);
xnor U4380 (N_4380,N_2022,N_3356);
nor U4381 (N_4381,N_2676,N_3576);
or U4382 (N_4382,N_2737,N_2464);
and U4383 (N_4383,N_3804,N_2629);
and U4384 (N_4384,N_2643,N_2463);
nor U4385 (N_4385,N_2804,N_3106);
nand U4386 (N_4386,N_2117,N_2935);
or U4387 (N_4387,N_2250,N_3989);
and U4388 (N_4388,N_3593,N_2725);
nand U4389 (N_4389,N_2131,N_3328);
nor U4390 (N_4390,N_3121,N_2814);
or U4391 (N_4391,N_3144,N_2123);
and U4392 (N_4392,N_2723,N_2895);
and U4393 (N_4393,N_3091,N_3336);
or U4394 (N_4394,N_2817,N_2397);
nor U4395 (N_4395,N_3344,N_3858);
nand U4396 (N_4396,N_3893,N_2502);
nand U4397 (N_4397,N_2941,N_3909);
nor U4398 (N_4398,N_3004,N_3032);
or U4399 (N_4399,N_2699,N_3698);
or U4400 (N_4400,N_2844,N_3736);
or U4401 (N_4401,N_3976,N_2302);
xor U4402 (N_4402,N_3820,N_3430);
nand U4403 (N_4403,N_3138,N_2175);
nand U4404 (N_4404,N_3166,N_2162);
xor U4405 (N_4405,N_2764,N_3226);
and U4406 (N_4406,N_2360,N_3081);
nand U4407 (N_4407,N_2972,N_2608);
nor U4408 (N_4408,N_2362,N_3763);
nor U4409 (N_4409,N_3465,N_3886);
xnor U4410 (N_4410,N_3746,N_3634);
or U4411 (N_4411,N_3532,N_3048);
nor U4412 (N_4412,N_2148,N_3852);
xor U4413 (N_4413,N_2451,N_3142);
xnor U4414 (N_4414,N_2742,N_3611);
and U4415 (N_4415,N_2210,N_2065);
xnor U4416 (N_4416,N_2733,N_3370);
nor U4417 (N_4417,N_2274,N_2012);
nand U4418 (N_4418,N_2121,N_2983);
and U4419 (N_4419,N_3632,N_2096);
xnor U4420 (N_4420,N_3937,N_2872);
nand U4421 (N_4421,N_2413,N_3911);
nor U4422 (N_4422,N_2828,N_2756);
nand U4423 (N_4423,N_2662,N_3960);
nor U4424 (N_4424,N_2320,N_3371);
or U4425 (N_4425,N_3670,N_3392);
nand U4426 (N_4426,N_2293,N_2051);
or U4427 (N_4427,N_2325,N_3849);
and U4428 (N_4428,N_3705,N_3388);
or U4429 (N_4429,N_3141,N_2552);
nand U4430 (N_4430,N_3066,N_2757);
or U4431 (N_4431,N_3955,N_3619);
nand U4432 (N_4432,N_3790,N_2685);
nor U4433 (N_4433,N_2719,N_3549);
or U4434 (N_4434,N_3987,N_3484);
and U4435 (N_4435,N_3799,N_2033);
or U4436 (N_4436,N_3650,N_3984);
nor U4437 (N_4437,N_2163,N_2160);
xnor U4438 (N_4438,N_3182,N_3494);
xor U4439 (N_4439,N_2050,N_3575);
and U4440 (N_4440,N_2089,N_2818);
xor U4441 (N_4441,N_3825,N_2582);
or U4442 (N_4442,N_2438,N_2894);
xnor U4443 (N_4443,N_3647,N_3508);
xor U4444 (N_4444,N_2886,N_2641);
or U4445 (N_4445,N_3878,N_3488);
and U4446 (N_4446,N_3179,N_2888);
or U4447 (N_4447,N_2921,N_2843);
xor U4448 (N_4448,N_2259,N_3442);
or U4449 (N_4449,N_3817,N_2750);
nand U4450 (N_4450,N_2539,N_2166);
nor U4451 (N_4451,N_2021,N_2525);
or U4452 (N_4452,N_3248,N_2319);
nand U4453 (N_4453,N_2652,N_3204);
xor U4454 (N_4454,N_3217,N_2560);
and U4455 (N_4455,N_3414,N_3728);
nand U4456 (N_4456,N_2558,N_2260);
xnor U4457 (N_4457,N_2432,N_2453);
or U4458 (N_4458,N_3464,N_2759);
or U4459 (N_4459,N_2187,N_2621);
or U4460 (N_4460,N_3998,N_2140);
xnor U4461 (N_4461,N_2974,N_2544);
and U4462 (N_4462,N_2275,N_3052);
xnor U4463 (N_4463,N_2969,N_3625);
or U4464 (N_4464,N_2930,N_3463);
xnor U4465 (N_4465,N_3111,N_3819);
xnor U4466 (N_4466,N_2516,N_3238);
or U4467 (N_4467,N_2007,N_3007);
xnor U4468 (N_4468,N_2732,N_3722);
or U4469 (N_4469,N_3927,N_3885);
xor U4470 (N_4470,N_2561,N_2256);
xor U4471 (N_4471,N_3792,N_2786);
xnor U4472 (N_4472,N_2847,N_2267);
nor U4473 (N_4473,N_2186,N_2936);
xor U4474 (N_4474,N_2867,N_2570);
or U4475 (N_4475,N_2952,N_3220);
nand U4476 (N_4476,N_2842,N_3604);
nand U4477 (N_4477,N_3112,N_2526);
and U4478 (N_4478,N_3629,N_3578);
xnor U4479 (N_4479,N_3110,N_2845);
and U4480 (N_4480,N_3779,N_2125);
and U4481 (N_4481,N_3403,N_3035);
nor U4482 (N_4482,N_2964,N_3262);
xnor U4483 (N_4483,N_2283,N_3478);
and U4484 (N_4484,N_3481,N_2157);
and U4485 (N_4485,N_2305,N_2863);
and U4486 (N_4486,N_3349,N_2741);
xnor U4487 (N_4487,N_3840,N_2388);
xor U4488 (N_4488,N_3999,N_2975);
nand U4489 (N_4489,N_3417,N_3924);
xnor U4490 (N_4490,N_3456,N_3623);
or U4491 (N_4491,N_2663,N_2503);
nor U4492 (N_4492,N_2149,N_3771);
or U4493 (N_4493,N_3708,N_3928);
and U4494 (N_4494,N_3367,N_2885);
nor U4495 (N_4495,N_3585,N_2064);
and U4496 (N_4496,N_2443,N_3538);
and U4497 (N_4497,N_3701,N_2666);
or U4498 (N_4498,N_2978,N_2195);
or U4499 (N_4499,N_2785,N_2590);
nand U4500 (N_4500,N_3669,N_3569);
or U4501 (N_4501,N_2336,N_3846);
and U4502 (N_4502,N_2875,N_3304);
or U4503 (N_4503,N_2315,N_2261);
nor U4504 (N_4504,N_2899,N_3424);
nand U4505 (N_4505,N_2791,N_2768);
and U4506 (N_4506,N_2054,N_2180);
and U4507 (N_4507,N_2835,N_2740);
xor U4508 (N_4508,N_3641,N_2150);
xnor U4509 (N_4509,N_2379,N_3938);
nor U4510 (N_4510,N_3155,N_2810);
or U4511 (N_4511,N_2634,N_3520);
and U4512 (N_4512,N_2527,N_3202);
nand U4513 (N_4513,N_3256,N_2047);
nand U4514 (N_4514,N_3971,N_3652);
or U4515 (N_4515,N_3681,N_2735);
nand U4516 (N_4516,N_3715,N_3169);
nand U4517 (N_4517,N_3178,N_3949);
nor U4518 (N_4518,N_2517,N_3577);
nor U4519 (N_4519,N_3086,N_2435);
nand U4520 (N_4520,N_2626,N_2650);
nor U4521 (N_4521,N_2070,N_3720);
nand U4522 (N_4522,N_3366,N_3942);
and U4523 (N_4523,N_2573,N_2529);
nor U4524 (N_4524,N_3255,N_3176);
or U4525 (N_4525,N_3996,N_2467);
and U4526 (N_4526,N_3285,N_2271);
nor U4527 (N_4527,N_3194,N_2985);
nand U4528 (N_4528,N_2547,N_3616);
nor U4529 (N_4529,N_3678,N_3477);
nand U4530 (N_4530,N_3800,N_2965);
nand U4531 (N_4531,N_3228,N_2567);
or U4532 (N_4532,N_2158,N_3853);
xor U4533 (N_4533,N_2788,N_2120);
and U4534 (N_4534,N_3908,N_2191);
and U4535 (N_4535,N_3028,N_2862);
nor U4536 (N_4536,N_2450,N_2787);
xor U4537 (N_4537,N_3559,N_3080);
nor U4538 (N_4538,N_3023,N_3572);
and U4539 (N_4539,N_2538,N_2203);
xnor U4540 (N_4540,N_3092,N_3841);
nor U4541 (N_4541,N_3500,N_2861);
nand U4542 (N_4542,N_3033,N_3546);
or U4543 (N_4543,N_2554,N_2928);
and U4544 (N_4544,N_2999,N_3748);
and U4545 (N_4545,N_3354,N_2937);
or U4546 (N_4546,N_3731,N_2342);
and U4547 (N_4547,N_2049,N_2869);
or U4548 (N_4548,N_2357,N_3966);
nor U4549 (N_4549,N_2306,N_3592);
or U4550 (N_4550,N_3287,N_3325);
or U4551 (N_4551,N_2129,N_3335);
nor U4552 (N_4552,N_2628,N_3544);
and U4553 (N_4553,N_3475,N_3770);
nand U4554 (N_4554,N_2546,N_2749);
or U4555 (N_4555,N_3319,N_2371);
and U4556 (N_4556,N_3338,N_2854);
and U4557 (N_4557,N_2292,N_2416);
and U4558 (N_4558,N_3551,N_3098);
or U4559 (N_4559,N_3342,N_3561);
nand U4560 (N_4560,N_2061,N_2940);
or U4561 (N_4561,N_2769,N_3677);
xnor U4562 (N_4562,N_2826,N_3514);
nand U4563 (N_4563,N_2395,N_2103);
and U4564 (N_4564,N_2077,N_2953);
xnor U4565 (N_4565,N_3348,N_3381);
nand U4566 (N_4566,N_3462,N_2279);
and U4567 (N_4567,N_2113,N_3898);
and U4568 (N_4568,N_3389,N_2549);
and U4569 (N_4569,N_3661,N_2426);
nand U4570 (N_4570,N_2603,N_3516);
or U4571 (N_4571,N_2713,N_2829);
nor U4572 (N_4572,N_3518,N_3125);
xor U4573 (N_4573,N_3041,N_3317);
and U4574 (N_4574,N_2651,N_2358);
nor U4575 (N_4575,N_2060,N_2238);
or U4576 (N_4576,N_2697,N_3445);
nand U4577 (N_4577,N_3101,N_3171);
nand U4578 (N_4578,N_2010,N_2528);
and U4579 (N_4579,N_2827,N_3847);
nand U4580 (N_4580,N_2639,N_3119);
and U4581 (N_4581,N_3190,N_2700);
nor U4582 (N_4582,N_2314,N_3329);
nor U4583 (N_4583,N_2681,N_2648);
and U4584 (N_4584,N_2425,N_3829);
xnor U4585 (N_4585,N_3030,N_2185);
and U4586 (N_4586,N_3135,N_2671);
nor U4587 (N_4587,N_2812,N_3765);
xor U4588 (N_4588,N_2993,N_2614);
and U4589 (N_4589,N_3115,N_2522);
or U4590 (N_4590,N_2945,N_2819);
or U4591 (N_4591,N_2201,N_2015);
xnor U4592 (N_4592,N_3679,N_2152);
or U4593 (N_4593,N_3036,N_3618);
nor U4594 (N_4594,N_3810,N_3912);
or U4595 (N_4595,N_3589,N_3787);
nor U4596 (N_4596,N_3082,N_3979);
nor U4597 (N_4597,N_3164,N_2029);
and U4598 (N_4598,N_2976,N_3499);
and U4599 (N_4599,N_2492,N_2001);
and U4600 (N_4600,N_2656,N_3419);
and U4601 (N_4601,N_2264,N_3008);
or U4602 (N_4602,N_2361,N_3743);
and U4603 (N_4603,N_3065,N_3461);
xnor U4604 (N_4604,N_2255,N_3550);
nand U4605 (N_4605,N_3073,N_2778);
xnor U4606 (N_4606,N_2476,N_2139);
and U4607 (N_4607,N_2480,N_2534);
xnor U4608 (N_4608,N_3862,N_3268);
or U4609 (N_4609,N_3212,N_2568);
xor U4610 (N_4610,N_2244,N_3545);
or U4611 (N_4611,N_2913,N_3275);
or U4612 (N_4612,N_3038,N_2016);
xnor U4613 (N_4613,N_2363,N_3161);
nand U4614 (N_4614,N_3970,N_3875);
and U4615 (N_4615,N_3232,N_2914);
nand U4616 (N_4616,N_2484,N_3343);
xnor U4617 (N_4617,N_2551,N_3213);
and U4618 (N_4618,N_2402,N_3969);
nand U4619 (N_4619,N_2400,N_2533);
nand U4620 (N_4620,N_2571,N_2472);
nor U4621 (N_4621,N_2285,N_2596);
nor U4622 (N_4622,N_3502,N_2168);
or U4623 (N_4623,N_2298,N_2500);
xnor U4624 (N_4624,N_2459,N_3396);
xnor U4625 (N_4625,N_3769,N_2068);
or U4626 (N_4626,N_3327,N_2072);
xor U4627 (N_4627,N_3861,N_3511);
nand U4628 (N_4628,N_2424,N_3880);
and U4629 (N_4629,N_2698,N_2988);
or U4630 (N_4630,N_3090,N_2220);
and U4631 (N_4631,N_3521,N_3024);
xor U4632 (N_4632,N_2296,N_2934);
and U4633 (N_4633,N_2898,N_3148);
nor U4634 (N_4634,N_3379,N_2341);
and U4635 (N_4635,N_2948,N_2270);
or U4636 (N_4636,N_2726,N_3607);
nor U4637 (N_4637,N_2161,N_3026);
xnor U4638 (N_4638,N_2808,N_3000);
xnor U4639 (N_4639,N_2136,N_3482);
or U4640 (N_4640,N_2855,N_3872);
nand U4641 (N_4641,N_2973,N_2661);
or U4642 (N_4642,N_2659,N_2367);
nor U4643 (N_4643,N_3537,N_2618);
and U4644 (N_4644,N_3064,N_3899);
or U4645 (N_4645,N_3599,N_2631);
xor U4646 (N_4646,N_2760,N_2101);
and U4647 (N_4647,N_3707,N_2832);
and U4648 (N_4648,N_2841,N_2980);
or U4649 (N_4649,N_2530,N_2146);
or U4650 (N_4650,N_2674,N_3547);
and U4651 (N_4651,N_3473,N_2303);
or U4652 (N_4652,N_3402,N_3206);
nand U4653 (N_4653,N_3496,N_2224);
xnor U4654 (N_4654,N_2585,N_2019);
xor U4655 (N_4655,N_2605,N_2171);
xnor U4656 (N_4656,N_3236,N_3814);
xnor U4657 (N_4657,N_2781,N_2837);
xor U4658 (N_4658,N_3314,N_3628);
xnor U4659 (N_4659,N_2456,N_3540);
and U4660 (N_4660,N_2222,N_2020);
or U4661 (N_4661,N_3324,N_2172);
nand U4662 (N_4662,N_3609,N_2727);
nand U4663 (N_4663,N_3413,N_3815);
nand U4664 (N_4664,N_3001,N_3016);
nand U4665 (N_4665,N_2882,N_2653);
and U4666 (N_4666,N_3754,N_2100);
xnor U4667 (N_4667,N_2212,N_2272);
xnor U4668 (N_4668,N_3045,N_3214);
and U4669 (N_4669,N_3952,N_2245);
xnor U4670 (N_4670,N_3636,N_2859);
nor U4671 (N_4671,N_3025,N_2326);
or U4672 (N_4672,N_3418,N_2754);
xor U4673 (N_4673,N_3010,N_2430);
or U4674 (N_4674,N_3132,N_3767);
nand U4675 (N_4675,N_2209,N_3140);
and U4676 (N_4676,N_2406,N_3034);
or U4677 (N_4677,N_2672,N_3274);
nor U4678 (N_4678,N_2044,N_3531);
xor U4679 (N_4679,N_2564,N_3222);
or U4680 (N_4680,N_2821,N_3269);
nor U4681 (N_4681,N_2471,N_3231);
xor U4682 (N_4682,N_2891,N_3699);
xor U4683 (N_4683,N_2394,N_2108);
nor U4684 (N_4684,N_3801,N_3096);
and U4685 (N_4685,N_2429,N_3926);
and U4686 (N_4686,N_3830,N_3339);
nand U4687 (N_4687,N_2048,N_2414);
xor U4688 (N_4688,N_3768,N_2900);
or U4689 (N_4689,N_2926,N_3671);
nand U4690 (N_4690,N_2411,N_2299);
and U4691 (N_4691,N_3012,N_3945);
or U4692 (N_4692,N_3435,N_3046);
or U4693 (N_4693,N_2884,N_2729);
nor U4694 (N_4694,N_3580,N_2838);
or U4695 (N_4695,N_3246,N_2246);
xor U4696 (N_4696,N_2346,N_2234);
or U4697 (N_4697,N_2093,N_3892);
xnor U4698 (N_4698,N_3264,N_3741);
nor U4699 (N_4699,N_3740,N_3870);
nor U4700 (N_4700,N_2712,N_2249);
xor U4701 (N_4701,N_2128,N_2181);
nand U4702 (N_4702,N_3856,N_3139);
and U4703 (N_4703,N_2620,N_3261);
and U4704 (N_4704,N_2159,N_2392);
xor U4705 (N_4705,N_3105,N_3543);
and U4706 (N_4706,N_2813,N_2390);
nor U4707 (N_4707,N_2000,N_2127);
and U4708 (N_4708,N_2023,N_3393);
nor U4709 (N_4709,N_3633,N_2866);
xor U4710 (N_4710,N_2495,N_2439);
and U4711 (N_4711,N_3978,N_3816);
or U4712 (N_4712,N_3659,N_3458);
nand U4713 (N_4713,N_2701,N_2689);
and U4714 (N_4714,N_3357,N_3118);
and U4715 (N_4715,N_2446,N_2718);
nand U4716 (N_4716,N_3303,N_2269);
nor U4717 (N_4717,N_3515,N_3977);
xnor U4718 (N_4718,N_3714,N_3582);
nor U4719 (N_4719,N_3605,N_2396);
or U4720 (N_4720,N_2678,N_2436);
or U4721 (N_4721,N_2668,N_2865);
and U4722 (N_4722,N_3497,N_3992);
nor U4723 (N_4723,N_3680,N_3333);
and U4724 (N_4724,N_2918,N_3891);
nor U4725 (N_4725,N_3230,N_2354);
nor U4726 (N_4726,N_3842,N_2997);
or U4727 (N_4727,N_2688,N_2915);
or U4728 (N_4728,N_3457,N_2562);
nor U4729 (N_4729,N_2176,N_3873);
and U4730 (N_4730,N_2095,N_2679);
xnor U4731 (N_4731,N_2509,N_3277);
xnor U4732 (N_4732,N_3079,N_2038);
and U4733 (N_4733,N_3950,N_3584);
nand U4734 (N_4734,N_3386,N_2715);
xnor U4735 (N_4735,N_3130,N_3688);
xor U4736 (N_4736,N_3443,N_3542);
and U4737 (N_4737,N_2344,N_3534);
or U4738 (N_4738,N_2947,N_3361);
and U4739 (N_4739,N_2613,N_2849);
and U4740 (N_4740,N_2174,N_2179);
xnor U4741 (N_4741,N_3400,N_2106);
nand U4742 (N_4742,N_2074,N_2197);
xnor U4743 (N_4743,N_2287,N_3021);
nand U4744 (N_4744,N_3018,N_3838);
nor U4745 (N_4745,N_3102,N_2277);
or U4746 (N_4746,N_2075,N_3712);
nor U4747 (N_4747,N_3405,N_2232);
and U4748 (N_4748,N_2901,N_2483);
or U4749 (N_4749,N_3702,N_3774);
and U4750 (N_4750,N_3982,N_2003);
xor U4751 (N_4751,N_2334,N_2998);
and U4752 (N_4752,N_3006,N_3793);
xor U4753 (N_4753,N_3466,N_3203);
nand U4754 (N_4754,N_2929,N_3718);
or U4755 (N_4755,N_2711,N_3620);
and U4756 (N_4756,N_3762,N_2505);
and U4757 (N_4757,N_2846,N_2942);
or U4758 (N_4758,N_2086,N_2248);
nor U4759 (N_4759,N_2669,N_3606);
nand U4760 (N_4760,N_2910,N_3174);
xor U4761 (N_4761,N_3850,N_2118);
nand U4762 (N_4762,N_2092,N_3655);
nor U4763 (N_4763,N_2366,N_2489);
nand U4764 (N_4764,N_3181,N_3711);
nor U4765 (N_4765,N_3848,N_3301);
nand U4766 (N_4766,N_2745,N_3621);
and U4767 (N_4767,N_2002,N_2649);
and U4768 (N_4768,N_2469,N_2465);
nand U4769 (N_4769,N_3308,N_2811);
nor U4770 (N_4770,N_3761,N_2905);
nand U4771 (N_4771,N_3733,N_3726);
nand U4772 (N_4772,N_2577,N_3794);
and U4773 (N_4773,N_3498,N_2943);
nand U4774 (N_4774,N_3067,N_3811);
or U4775 (N_4775,N_2116,N_3922);
and U4776 (N_4776,N_3991,N_2693);
nor U4777 (N_4777,N_3412,N_2925);
nor U4778 (N_4778,N_3608,N_2474);
xnor U4779 (N_4779,N_3947,N_3973);
and U4780 (N_4780,N_3835,N_3622);
or U4781 (N_4781,N_2755,N_2199);
or U4782 (N_4782,N_2646,N_2257);
nand U4783 (N_4783,N_2097,N_2984);
or U4784 (N_4784,N_2153,N_3745);
nand U4785 (N_4785,N_3372,N_2034);
or U4786 (N_4786,N_2377,N_3932);
xnor U4787 (N_4787,N_3027,N_3676);
and U4788 (N_4788,N_3087,N_3975);
xor U4789 (N_4789,N_2420,N_3595);
nand U4790 (N_4790,N_2373,N_3003);
nand U4791 (N_4791,N_3894,N_2816);
nand U4792 (N_4792,N_2407,N_3666);
nand U4793 (N_4793,N_3781,N_3114);
xor U4794 (N_4794,N_3152,N_2110);
nand U4795 (N_4795,N_3907,N_2897);
nor U4796 (N_4796,N_2138,N_2738);
or U4797 (N_4797,N_2461,N_2680);
nand U4798 (N_4798,N_2982,N_3968);
and U4799 (N_4799,N_2254,N_3834);
nand U4800 (N_4800,N_3965,N_3351);
and U4801 (N_4801,N_3247,N_3321);
xnor U4802 (N_4802,N_3775,N_3197);
and U4803 (N_4803,N_3063,N_3925);
nor U4804 (N_4804,N_3828,N_2221);
or U4805 (N_4805,N_3536,N_3613);
nand U4806 (N_4806,N_3552,N_2916);
nor U4807 (N_4807,N_2421,N_2966);
or U4808 (N_4808,N_3113,N_2393);
or U4809 (N_4809,N_3103,N_2642);
nor U4810 (N_4810,N_2477,N_3245);
xnor U4811 (N_4811,N_3785,N_3668);
nand U4812 (N_4812,N_2486,N_3375);
nand U4813 (N_4813,N_3156,N_2889);
nor U4814 (N_4814,N_2566,N_2950);
nor U4815 (N_4815,N_2327,N_3205);
nand U4816 (N_4816,N_3280,N_2583);
or U4817 (N_4817,N_3263,N_3653);
nor U4818 (N_4818,N_3612,N_3272);
nand U4819 (N_4819,N_2114,N_2132);
and U4820 (N_4820,N_2604,N_2458);
nor U4821 (N_4821,N_2281,N_2036);
and U4822 (N_4822,N_3782,N_2079);
or U4823 (N_4823,N_3913,N_3921);
nor U4824 (N_4824,N_2949,N_2995);
xor U4825 (N_4825,N_2591,N_2479);
nor U4826 (N_4826,N_2062,N_3747);
and U4827 (N_4827,N_3695,N_3428);
nand U4828 (N_4828,N_2142,N_2041);
nand U4829 (N_4829,N_2217,N_3602);
xnor U4830 (N_4830,N_2115,N_2335);
nor U4831 (N_4831,N_3535,N_2008);
or U4832 (N_4832,N_2511,N_3583);
nor U4833 (N_4833,N_2722,N_2353);
nor U4834 (N_4834,N_2624,N_2076);
or U4835 (N_4835,N_2322,N_3753);
xor U4836 (N_4836,N_3648,N_3900);
and U4837 (N_4837,N_2352,N_3005);
and U4838 (N_4838,N_3523,N_2959);
nor U4839 (N_4839,N_2736,N_2398);
and U4840 (N_4840,N_3316,N_2482);
nand U4841 (N_4841,N_3777,N_3207);
or U4842 (N_4842,N_3143,N_2887);
or U4843 (N_4843,N_3116,N_2932);
xnor U4844 (N_4844,N_3168,N_3084);
nor U4845 (N_4845,N_3757,N_3491);
and U4846 (N_4846,N_3380,N_3954);
nand U4847 (N_4847,N_3594,N_3134);
xnor U4848 (N_4848,N_3879,N_3223);
or U4849 (N_4849,N_2686,N_2025);
nor U4850 (N_4850,N_3154,N_2784);
nor U4851 (N_4851,N_3108,N_2080);
xnor U4852 (N_4852,N_3685,N_3127);
nor U4853 (N_4853,N_3195,N_2035);
and U4854 (N_4854,N_2359,N_2278);
xor U4855 (N_4855,N_2204,N_2253);
or U4856 (N_4856,N_2870,N_2673);
xor U4857 (N_4857,N_3692,N_3172);
nor U4858 (N_4858,N_2099,N_3783);
nor U4859 (N_4859,N_2321,N_3083);
nor U4860 (N_4860,N_3469,N_3504);
or U4861 (N_4861,N_2944,N_3492);
xnor U4862 (N_4862,N_2389,N_2774);
or U4863 (N_4863,N_3468,N_3489);
xnor U4864 (N_4864,N_3694,N_3923);
and U4865 (N_4865,N_3565,N_2024);
nor U4866 (N_4866,N_3330,N_2751);
or U4867 (N_4867,N_3175,N_3675);
or U4868 (N_4868,N_3637,N_2444);
nand U4869 (N_4869,N_3129,N_3374);
nor U4870 (N_4870,N_2655,N_3614);
or U4871 (N_4871,N_3397,N_3667);
or U4872 (N_4872,N_3931,N_2557);
xor U4873 (N_4873,N_2380,N_2553);
or U4874 (N_4874,N_2497,N_2104);
and U4875 (N_4875,N_3505,N_2318);
or U4876 (N_4876,N_2868,N_3049);
nand U4877 (N_4877,N_3732,N_2063);
nor U4878 (N_4878,N_3050,N_3260);
nand U4879 (N_4879,N_3687,N_2478);
nor U4880 (N_4880,N_2519,N_3759);
xor U4881 (N_4881,N_3095,N_2610);
xnor U4882 (N_4882,N_3904,N_3234);
or U4883 (N_4883,N_3355,N_2419);
nor U4884 (N_4884,N_2102,N_2447);
and U4885 (N_4885,N_2977,N_2351);
nor U4886 (N_4886,N_2046,N_2992);
and U4887 (N_4887,N_2739,N_2297);
nor U4888 (N_4888,N_2761,N_3766);
xnor U4889 (N_4889,N_3281,N_3365);
or U4890 (N_4890,N_2164,N_3383);
and U4891 (N_4891,N_2189,N_2085);
nor U4892 (N_4892,N_2970,N_3689);
and U4893 (N_4893,N_3219,N_3744);
nor U4894 (N_4894,N_2391,N_3581);
nor U4895 (N_4895,N_3002,N_3273);
nor U4896 (N_4896,N_2028,N_2657);
and U4897 (N_4897,N_3128,N_2730);
and U4898 (N_4898,N_3044,N_2709);
nor U4899 (N_4899,N_3525,N_2454);
or U4900 (N_4900,N_2833,N_2853);
xor U4901 (N_4901,N_2385,N_3070);
nor U4902 (N_4902,N_2428,N_2112);
and U4903 (N_4903,N_2923,N_2917);
or U4904 (N_4904,N_3939,N_3972);
or U4905 (N_4905,N_3831,N_2169);
and U4906 (N_4906,N_2851,N_3136);
nand U4907 (N_4907,N_3640,N_3896);
nor U4908 (N_4908,N_2057,N_2227);
or U4909 (N_4909,N_2664,N_3093);
or U4910 (N_4910,N_3120,N_2496);
xnor U4911 (N_4911,N_2805,N_3029);
nand U4912 (N_4912,N_3020,N_3198);
nand U4913 (N_4913,N_3742,N_2960);
or U4914 (N_4914,N_2009,N_2824);
nor U4915 (N_4915,N_2627,N_2587);
xnor U4916 (N_4916,N_2219,N_2955);
or U4917 (N_4917,N_2369,N_3663);
or U4918 (N_4918,N_3635,N_3078);
nand U4919 (N_4919,N_3186,N_2055);
nor U4920 (N_4920,N_3730,N_3332);
and U4921 (N_4921,N_3568,N_3037);
nor U4922 (N_4922,N_3447,N_3215);
xor U4923 (N_4923,N_3229,N_2338);
and U4924 (N_4924,N_2265,N_2802);
and U4925 (N_4925,N_2850,N_3069);
or U4926 (N_4926,N_2797,N_2349);
nand U4927 (N_4927,N_2820,N_3437);
nor U4928 (N_4928,N_2871,N_3170);
nor U4929 (N_4929,N_2858,N_2111);
nor U4930 (N_4930,N_3454,N_3243);
xnor U4931 (N_4931,N_2896,N_2775);
xnor U4932 (N_4932,N_2682,N_2822);
nand U4933 (N_4933,N_3827,N_3764);
and U4934 (N_4934,N_3624,N_3476);
or U4935 (N_4935,N_3432,N_2263);
xnor U4936 (N_4936,N_2536,N_2798);
and U4937 (N_4937,N_3986,N_3874);
nand U4938 (N_4938,N_2423,N_2637);
xor U4939 (N_4939,N_3651,N_2611);
and U4940 (N_4940,N_3639,N_3776);
nand U4941 (N_4941,N_2848,N_3860);
or U4942 (N_4942,N_3208,N_2514);
and U4943 (N_4943,N_2555,N_3013);
and U4944 (N_4944,N_3920,N_3244);
or U4945 (N_4945,N_3399,N_3729);
or U4946 (N_4946,N_2310,N_2340);
xnor U4947 (N_4947,N_3358,N_3495);
nor U4948 (N_4948,N_2133,N_3359);
nand U4949 (N_4949,N_3567,N_3334);
nor U4950 (N_4950,N_3953,N_3826);
xor U4951 (N_4951,N_3133,N_3252);
nor U4952 (N_4952,N_3758,N_3780);
and U4953 (N_4953,N_3368,N_3553);
or U4954 (N_4954,N_3254,N_3401);
nand U4955 (N_4955,N_2475,N_2119);
nand U4956 (N_4956,N_3556,N_2638);
nand U4957 (N_4957,N_3253,N_3806);
nor U4958 (N_4958,N_2609,N_2262);
and U4959 (N_4959,N_3331,N_3369);
nand U4960 (N_4960,N_2622,N_3452);
nor U4961 (N_4961,N_3404,N_2746);
nand U4962 (N_4962,N_2403,N_3570);
xnor U4963 (N_4963,N_3270,N_2130);
nand U4964 (N_4964,N_2616,N_3642);
nor U4965 (N_4965,N_3471,N_3407);
xor U4966 (N_4966,N_2268,N_3257);
and U4967 (N_4967,N_3704,N_3302);
nand U4968 (N_4968,N_3241,N_3235);
and U4969 (N_4969,N_3094,N_2182);
xnor U4970 (N_4970,N_3455,N_3649);
or U4971 (N_4971,N_2907,N_2026);
and U4972 (N_4972,N_3409,N_2442);
or U4973 (N_4973,N_3990,N_3180);
nand U4974 (N_4974,N_3192,N_3292);
and U4975 (N_4975,N_2155,N_2083);
nand U4976 (N_4976,N_3011,N_2758);
xor U4977 (N_4977,N_2856,N_2939);
and U4978 (N_4978,N_2017,N_3901);
or U4979 (N_4979,N_2706,N_2251);
and U4980 (N_4980,N_3279,N_2329);
nand U4981 (N_4981,N_3313,N_3724);
xor U4982 (N_4982,N_2524,N_3294);
or U4983 (N_4983,N_3884,N_2548);
or U4984 (N_4984,N_2991,N_3813);
nand U4985 (N_4985,N_2720,N_3347);
nand U4986 (N_4986,N_2350,N_3562);
and U4987 (N_4987,N_3126,N_3734);
or U4988 (N_4988,N_3683,N_2088);
nor U4989 (N_4989,N_2137,N_3882);
nor U4990 (N_4990,N_2987,N_2852);
or U4991 (N_4991,N_2427,N_2879);
nand U4992 (N_4992,N_2714,N_2266);
or U4993 (N_4993,N_3054,N_3739);
nand U4994 (N_4994,N_2194,N_3818);
and U4995 (N_4995,N_3735,N_2996);
xnor U4996 (N_4996,N_2956,N_2911);
and U4997 (N_4997,N_2449,N_3251);
nor U4998 (N_4998,N_3345,N_2584);
and U4999 (N_4999,N_3919,N_3364);
nor U5000 (N_5000,N_3232,N_3245);
or U5001 (N_5001,N_3222,N_3401);
nand U5002 (N_5002,N_3943,N_3993);
xor U5003 (N_5003,N_2883,N_3549);
nand U5004 (N_5004,N_3601,N_3124);
or U5005 (N_5005,N_2150,N_3185);
xnor U5006 (N_5006,N_2403,N_3314);
and U5007 (N_5007,N_2303,N_2585);
or U5008 (N_5008,N_2681,N_2441);
xnor U5009 (N_5009,N_3445,N_2637);
nor U5010 (N_5010,N_2952,N_2203);
nand U5011 (N_5011,N_3456,N_3696);
nand U5012 (N_5012,N_3117,N_2940);
nand U5013 (N_5013,N_3269,N_2471);
and U5014 (N_5014,N_3990,N_3054);
or U5015 (N_5015,N_3175,N_2628);
or U5016 (N_5016,N_3583,N_2056);
xnor U5017 (N_5017,N_2546,N_3795);
and U5018 (N_5018,N_3337,N_2263);
xnor U5019 (N_5019,N_2525,N_2281);
and U5020 (N_5020,N_2837,N_2808);
nand U5021 (N_5021,N_2364,N_3873);
nand U5022 (N_5022,N_3004,N_2692);
xor U5023 (N_5023,N_3951,N_3740);
nor U5024 (N_5024,N_2117,N_3583);
or U5025 (N_5025,N_2541,N_2879);
and U5026 (N_5026,N_2511,N_2924);
xor U5027 (N_5027,N_2584,N_3121);
or U5028 (N_5028,N_2624,N_3675);
nor U5029 (N_5029,N_2993,N_2306);
nor U5030 (N_5030,N_3430,N_3793);
nand U5031 (N_5031,N_2426,N_3057);
or U5032 (N_5032,N_3501,N_3858);
nor U5033 (N_5033,N_3557,N_2590);
nor U5034 (N_5034,N_2513,N_3535);
xor U5035 (N_5035,N_3987,N_2509);
nor U5036 (N_5036,N_2445,N_2516);
nor U5037 (N_5037,N_3216,N_3627);
and U5038 (N_5038,N_3755,N_2159);
and U5039 (N_5039,N_3333,N_3866);
nand U5040 (N_5040,N_3015,N_3878);
nand U5041 (N_5041,N_2303,N_2607);
or U5042 (N_5042,N_3092,N_2237);
nand U5043 (N_5043,N_3487,N_3520);
or U5044 (N_5044,N_2672,N_2512);
or U5045 (N_5045,N_3453,N_2383);
nor U5046 (N_5046,N_3979,N_3315);
nor U5047 (N_5047,N_3431,N_2915);
and U5048 (N_5048,N_3519,N_2811);
nor U5049 (N_5049,N_2839,N_2126);
nand U5050 (N_5050,N_2086,N_3037);
and U5051 (N_5051,N_3279,N_3461);
or U5052 (N_5052,N_3426,N_3468);
nand U5053 (N_5053,N_3118,N_3880);
or U5054 (N_5054,N_2879,N_3549);
and U5055 (N_5055,N_3251,N_2047);
and U5056 (N_5056,N_2588,N_2342);
xnor U5057 (N_5057,N_3342,N_3190);
or U5058 (N_5058,N_2635,N_2322);
nor U5059 (N_5059,N_2238,N_3389);
or U5060 (N_5060,N_3018,N_3323);
or U5061 (N_5061,N_3325,N_3539);
nor U5062 (N_5062,N_2880,N_3447);
xnor U5063 (N_5063,N_3064,N_2833);
or U5064 (N_5064,N_2352,N_2854);
or U5065 (N_5065,N_2992,N_3466);
xnor U5066 (N_5066,N_3018,N_2811);
nor U5067 (N_5067,N_3362,N_3844);
or U5068 (N_5068,N_2091,N_2552);
nand U5069 (N_5069,N_2181,N_3858);
nand U5070 (N_5070,N_2848,N_2405);
nand U5071 (N_5071,N_2001,N_2698);
nor U5072 (N_5072,N_2107,N_2010);
nor U5073 (N_5073,N_3846,N_2141);
nor U5074 (N_5074,N_2110,N_2267);
xor U5075 (N_5075,N_3996,N_2280);
or U5076 (N_5076,N_3094,N_2991);
xnor U5077 (N_5077,N_2475,N_2718);
xnor U5078 (N_5078,N_3059,N_2268);
nand U5079 (N_5079,N_2370,N_2340);
nor U5080 (N_5080,N_2132,N_3815);
xnor U5081 (N_5081,N_2041,N_3090);
and U5082 (N_5082,N_3514,N_3112);
xor U5083 (N_5083,N_2152,N_2537);
nor U5084 (N_5084,N_3295,N_3990);
nand U5085 (N_5085,N_3103,N_2761);
nor U5086 (N_5086,N_2504,N_2076);
or U5087 (N_5087,N_2708,N_2832);
or U5088 (N_5088,N_2741,N_2441);
nand U5089 (N_5089,N_2517,N_2968);
nor U5090 (N_5090,N_3592,N_2694);
or U5091 (N_5091,N_2120,N_3671);
or U5092 (N_5092,N_3725,N_3368);
or U5093 (N_5093,N_3795,N_2160);
and U5094 (N_5094,N_3917,N_2921);
or U5095 (N_5095,N_2111,N_3483);
and U5096 (N_5096,N_2261,N_3494);
xor U5097 (N_5097,N_3014,N_3123);
or U5098 (N_5098,N_3742,N_2293);
and U5099 (N_5099,N_2491,N_2314);
or U5100 (N_5100,N_2185,N_2118);
xnor U5101 (N_5101,N_2207,N_2313);
and U5102 (N_5102,N_3995,N_2927);
nor U5103 (N_5103,N_2232,N_3316);
nand U5104 (N_5104,N_3704,N_2822);
nand U5105 (N_5105,N_3315,N_3513);
or U5106 (N_5106,N_3212,N_2810);
nor U5107 (N_5107,N_2150,N_3610);
nand U5108 (N_5108,N_2186,N_2531);
xor U5109 (N_5109,N_2744,N_3189);
and U5110 (N_5110,N_3153,N_2492);
nor U5111 (N_5111,N_3727,N_3408);
and U5112 (N_5112,N_2394,N_3450);
nor U5113 (N_5113,N_2451,N_3626);
nor U5114 (N_5114,N_2659,N_3501);
and U5115 (N_5115,N_3578,N_3206);
nor U5116 (N_5116,N_3062,N_2084);
or U5117 (N_5117,N_3502,N_3757);
xor U5118 (N_5118,N_2067,N_3921);
xor U5119 (N_5119,N_3607,N_2492);
nor U5120 (N_5120,N_2991,N_2749);
nand U5121 (N_5121,N_2311,N_3421);
and U5122 (N_5122,N_3739,N_2639);
nor U5123 (N_5123,N_2187,N_3717);
xor U5124 (N_5124,N_2341,N_2616);
xnor U5125 (N_5125,N_2414,N_2667);
xnor U5126 (N_5126,N_2965,N_3739);
nand U5127 (N_5127,N_2760,N_3236);
xor U5128 (N_5128,N_2002,N_3894);
or U5129 (N_5129,N_3940,N_3482);
xnor U5130 (N_5130,N_3446,N_3491);
or U5131 (N_5131,N_3188,N_3681);
and U5132 (N_5132,N_2511,N_3816);
or U5133 (N_5133,N_2167,N_2654);
nor U5134 (N_5134,N_2137,N_2163);
nor U5135 (N_5135,N_2052,N_2906);
and U5136 (N_5136,N_3076,N_2273);
xor U5137 (N_5137,N_2624,N_2959);
xnor U5138 (N_5138,N_2303,N_2289);
nor U5139 (N_5139,N_2711,N_2353);
nor U5140 (N_5140,N_3764,N_2502);
and U5141 (N_5141,N_2200,N_3354);
or U5142 (N_5142,N_2154,N_2238);
and U5143 (N_5143,N_2865,N_3368);
xnor U5144 (N_5144,N_3742,N_2211);
or U5145 (N_5145,N_2980,N_3193);
xor U5146 (N_5146,N_3328,N_2253);
nor U5147 (N_5147,N_2445,N_2141);
nand U5148 (N_5148,N_2758,N_3359);
nand U5149 (N_5149,N_3445,N_3362);
nor U5150 (N_5150,N_3812,N_2190);
and U5151 (N_5151,N_3712,N_2413);
xor U5152 (N_5152,N_2414,N_3655);
nand U5153 (N_5153,N_3850,N_3280);
nand U5154 (N_5154,N_2588,N_2717);
xor U5155 (N_5155,N_2487,N_3706);
and U5156 (N_5156,N_2185,N_2231);
nor U5157 (N_5157,N_3903,N_2075);
and U5158 (N_5158,N_2642,N_2860);
or U5159 (N_5159,N_2592,N_3078);
nand U5160 (N_5160,N_3958,N_3941);
or U5161 (N_5161,N_2328,N_2004);
nand U5162 (N_5162,N_3038,N_3835);
or U5163 (N_5163,N_2515,N_2338);
or U5164 (N_5164,N_2221,N_3161);
nor U5165 (N_5165,N_2042,N_2147);
and U5166 (N_5166,N_3695,N_2943);
xnor U5167 (N_5167,N_3759,N_2815);
or U5168 (N_5168,N_3710,N_3963);
nand U5169 (N_5169,N_2827,N_2558);
xor U5170 (N_5170,N_2394,N_2083);
and U5171 (N_5171,N_3082,N_2986);
xor U5172 (N_5172,N_2489,N_2556);
nand U5173 (N_5173,N_2856,N_2897);
xnor U5174 (N_5174,N_2391,N_3430);
nor U5175 (N_5175,N_3946,N_3578);
nand U5176 (N_5176,N_2840,N_3449);
nand U5177 (N_5177,N_2138,N_2670);
xnor U5178 (N_5178,N_3330,N_2552);
and U5179 (N_5179,N_2145,N_3958);
or U5180 (N_5180,N_2726,N_2033);
nor U5181 (N_5181,N_3218,N_3978);
nor U5182 (N_5182,N_2617,N_2644);
and U5183 (N_5183,N_2756,N_2902);
nand U5184 (N_5184,N_2190,N_3567);
and U5185 (N_5185,N_3284,N_2758);
nor U5186 (N_5186,N_3458,N_2617);
nand U5187 (N_5187,N_2805,N_3875);
nor U5188 (N_5188,N_3262,N_2537);
or U5189 (N_5189,N_2786,N_3087);
or U5190 (N_5190,N_3472,N_3836);
or U5191 (N_5191,N_2015,N_2310);
nand U5192 (N_5192,N_3359,N_2347);
or U5193 (N_5193,N_2103,N_2026);
and U5194 (N_5194,N_3828,N_3641);
nor U5195 (N_5195,N_3148,N_2015);
or U5196 (N_5196,N_2348,N_3665);
xnor U5197 (N_5197,N_2410,N_2781);
nor U5198 (N_5198,N_2646,N_2445);
nor U5199 (N_5199,N_3051,N_3521);
or U5200 (N_5200,N_3693,N_2824);
nand U5201 (N_5201,N_2146,N_3441);
or U5202 (N_5202,N_2380,N_2376);
xor U5203 (N_5203,N_2721,N_2302);
nor U5204 (N_5204,N_3302,N_3188);
or U5205 (N_5205,N_3320,N_2851);
nor U5206 (N_5206,N_2453,N_3036);
xor U5207 (N_5207,N_3687,N_3330);
xor U5208 (N_5208,N_2452,N_2209);
nor U5209 (N_5209,N_3022,N_2311);
and U5210 (N_5210,N_3574,N_3561);
or U5211 (N_5211,N_2997,N_2365);
or U5212 (N_5212,N_3919,N_2595);
xor U5213 (N_5213,N_3573,N_2788);
xor U5214 (N_5214,N_3340,N_2107);
nand U5215 (N_5215,N_2332,N_2545);
nor U5216 (N_5216,N_2329,N_2341);
and U5217 (N_5217,N_2503,N_3739);
and U5218 (N_5218,N_2623,N_3792);
or U5219 (N_5219,N_2674,N_3698);
and U5220 (N_5220,N_3550,N_2211);
nand U5221 (N_5221,N_3913,N_3456);
nor U5222 (N_5222,N_3097,N_3485);
nand U5223 (N_5223,N_2547,N_3227);
nand U5224 (N_5224,N_2422,N_3077);
nand U5225 (N_5225,N_3645,N_2452);
and U5226 (N_5226,N_2566,N_3158);
xor U5227 (N_5227,N_2674,N_2023);
nand U5228 (N_5228,N_2113,N_3832);
nor U5229 (N_5229,N_3617,N_3938);
or U5230 (N_5230,N_2193,N_3235);
and U5231 (N_5231,N_3787,N_3997);
nor U5232 (N_5232,N_3149,N_2006);
and U5233 (N_5233,N_3774,N_2298);
xnor U5234 (N_5234,N_2425,N_2551);
nand U5235 (N_5235,N_3270,N_2111);
and U5236 (N_5236,N_2093,N_3885);
and U5237 (N_5237,N_3997,N_3526);
nand U5238 (N_5238,N_3739,N_3032);
xnor U5239 (N_5239,N_2926,N_2271);
or U5240 (N_5240,N_2638,N_2272);
nor U5241 (N_5241,N_2224,N_2281);
xnor U5242 (N_5242,N_2520,N_3402);
xnor U5243 (N_5243,N_3627,N_2258);
nor U5244 (N_5244,N_2670,N_2513);
and U5245 (N_5245,N_3828,N_2807);
xnor U5246 (N_5246,N_3155,N_2104);
nand U5247 (N_5247,N_3050,N_2416);
and U5248 (N_5248,N_3288,N_3451);
and U5249 (N_5249,N_3544,N_2460);
or U5250 (N_5250,N_2605,N_3430);
or U5251 (N_5251,N_3256,N_3419);
nand U5252 (N_5252,N_2276,N_3889);
nor U5253 (N_5253,N_3623,N_2180);
nor U5254 (N_5254,N_2693,N_3707);
nand U5255 (N_5255,N_2629,N_2981);
or U5256 (N_5256,N_2046,N_2999);
nand U5257 (N_5257,N_3389,N_2514);
nor U5258 (N_5258,N_3528,N_3200);
or U5259 (N_5259,N_3857,N_2961);
and U5260 (N_5260,N_3808,N_2197);
and U5261 (N_5261,N_3068,N_2851);
xor U5262 (N_5262,N_3044,N_2022);
xor U5263 (N_5263,N_2111,N_3819);
xor U5264 (N_5264,N_3237,N_2770);
or U5265 (N_5265,N_2405,N_3184);
and U5266 (N_5266,N_3587,N_3848);
xor U5267 (N_5267,N_3481,N_3706);
or U5268 (N_5268,N_3791,N_3862);
xor U5269 (N_5269,N_3599,N_3659);
nor U5270 (N_5270,N_3026,N_3220);
and U5271 (N_5271,N_2079,N_3296);
and U5272 (N_5272,N_2175,N_3310);
nand U5273 (N_5273,N_3107,N_3988);
or U5274 (N_5274,N_3246,N_3726);
or U5275 (N_5275,N_2354,N_2756);
and U5276 (N_5276,N_3006,N_2643);
nor U5277 (N_5277,N_2248,N_3526);
or U5278 (N_5278,N_2511,N_2730);
and U5279 (N_5279,N_2761,N_2890);
or U5280 (N_5280,N_3054,N_2903);
xor U5281 (N_5281,N_2511,N_3981);
nand U5282 (N_5282,N_3860,N_2117);
or U5283 (N_5283,N_2310,N_2288);
xnor U5284 (N_5284,N_3631,N_3395);
and U5285 (N_5285,N_3313,N_3730);
and U5286 (N_5286,N_3736,N_3291);
xor U5287 (N_5287,N_3708,N_3451);
nor U5288 (N_5288,N_3182,N_3417);
and U5289 (N_5289,N_2960,N_2455);
or U5290 (N_5290,N_3980,N_3932);
nand U5291 (N_5291,N_2215,N_2701);
xor U5292 (N_5292,N_3559,N_3082);
xnor U5293 (N_5293,N_2156,N_3861);
and U5294 (N_5294,N_2533,N_3559);
and U5295 (N_5295,N_3112,N_3264);
and U5296 (N_5296,N_2030,N_2154);
nor U5297 (N_5297,N_2871,N_3289);
nand U5298 (N_5298,N_3714,N_3402);
xor U5299 (N_5299,N_2485,N_3817);
nand U5300 (N_5300,N_3473,N_2170);
nand U5301 (N_5301,N_3881,N_3114);
and U5302 (N_5302,N_2451,N_3855);
nand U5303 (N_5303,N_2640,N_3210);
xnor U5304 (N_5304,N_3742,N_2433);
nand U5305 (N_5305,N_2996,N_3456);
nor U5306 (N_5306,N_3208,N_2985);
or U5307 (N_5307,N_2851,N_3945);
xor U5308 (N_5308,N_2421,N_2743);
nand U5309 (N_5309,N_2370,N_2745);
or U5310 (N_5310,N_3221,N_2814);
nor U5311 (N_5311,N_3573,N_3992);
xor U5312 (N_5312,N_3646,N_2988);
xor U5313 (N_5313,N_3132,N_2222);
and U5314 (N_5314,N_3321,N_3824);
and U5315 (N_5315,N_2007,N_2682);
nor U5316 (N_5316,N_2992,N_2292);
xnor U5317 (N_5317,N_2653,N_3530);
nor U5318 (N_5318,N_3953,N_3685);
or U5319 (N_5319,N_3394,N_3215);
nor U5320 (N_5320,N_3936,N_3051);
or U5321 (N_5321,N_2401,N_3288);
xor U5322 (N_5322,N_3225,N_2684);
nor U5323 (N_5323,N_3434,N_2539);
nand U5324 (N_5324,N_3975,N_3980);
xor U5325 (N_5325,N_2901,N_3554);
nand U5326 (N_5326,N_2927,N_3885);
nand U5327 (N_5327,N_2064,N_3035);
or U5328 (N_5328,N_3634,N_3059);
and U5329 (N_5329,N_3233,N_2697);
or U5330 (N_5330,N_3161,N_2591);
nand U5331 (N_5331,N_2160,N_3041);
xor U5332 (N_5332,N_3127,N_3108);
xor U5333 (N_5333,N_3973,N_2821);
and U5334 (N_5334,N_3629,N_3547);
nand U5335 (N_5335,N_2412,N_2232);
xor U5336 (N_5336,N_2851,N_2148);
xnor U5337 (N_5337,N_2665,N_3883);
and U5338 (N_5338,N_3166,N_3144);
and U5339 (N_5339,N_2891,N_3178);
xor U5340 (N_5340,N_3535,N_2864);
nor U5341 (N_5341,N_2082,N_2517);
and U5342 (N_5342,N_3268,N_3502);
and U5343 (N_5343,N_2072,N_3305);
xor U5344 (N_5344,N_3842,N_2429);
or U5345 (N_5345,N_3543,N_3206);
or U5346 (N_5346,N_2494,N_3980);
nor U5347 (N_5347,N_3438,N_2486);
or U5348 (N_5348,N_3821,N_3888);
or U5349 (N_5349,N_2299,N_3394);
nand U5350 (N_5350,N_3921,N_3852);
xnor U5351 (N_5351,N_3818,N_3455);
and U5352 (N_5352,N_2682,N_2392);
nand U5353 (N_5353,N_2766,N_3488);
xor U5354 (N_5354,N_3562,N_3640);
and U5355 (N_5355,N_3416,N_2920);
xor U5356 (N_5356,N_2412,N_3684);
nand U5357 (N_5357,N_3412,N_3671);
or U5358 (N_5358,N_2443,N_3098);
xnor U5359 (N_5359,N_2490,N_2998);
or U5360 (N_5360,N_3658,N_2806);
nor U5361 (N_5361,N_2918,N_2016);
nor U5362 (N_5362,N_2845,N_2685);
or U5363 (N_5363,N_3287,N_3516);
nor U5364 (N_5364,N_2590,N_3079);
nor U5365 (N_5365,N_2460,N_3337);
nand U5366 (N_5366,N_3749,N_3158);
or U5367 (N_5367,N_3450,N_2165);
xnor U5368 (N_5368,N_3759,N_2570);
nor U5369 (N_5369,N_3459,N_3475);
xor U5370 (N_5370,N_2561,N_3917);
and U5371 (N_5371,N_3816,N_2323);
or U5372 (N_5372,N_2684,N_2632);
nor U5373 (N_5373,N_2715,N_3181);
nor U5374 (N_5374,N_2434,N_2829);
nand U5375 (N_5375,N_3600,N_3588);
and U5376 (N_5376,N_3182,N_2032);
or U5377 (N_5377,N_3395,N_3701);
or U5378 (N_5378,N_3335,N_3731);
and U5379 (N_5379,N_3952,N_3739);
nand U5380 (N_5380,N_3097,N_3785);
and U5381 (N_5381,N_2411,N_2934);
or U5382 (N_5382,N_3085,N_2695);
or U5383 (N_5383,N_2261,N_2969);
nand U5384 (N_5384,N_2338,N_2070);
xor U5385 (N_5385,N_2601,N_3879);
xnor U5386 (N_5386,N_2459,N_3258);
and U5387 (N_5387,N_2087,N_3389);
nand U5388 (N_5388,N_2803,N_2189);
nand U5389 (N_5389,N_3748,N_3745);
xnor U5390 (N_5390,N_2693,N_3036);
xnor U5391 (N_5391,N_2282,N_3876);
nor U5392 (N_5392,N_2561,N_2200);
nand U5393 (N_5393,N_3397,N_3633);
nand U5394 (N_5394,N_2809,N_2796);
or U5395 (N_5395,N_2388,N_3674);
nand U5396 (N_5396,N_2611,N_2746);
xnor U5397 (N_5397,N_2208,N_3271);
nand U5398 (N_5398,N_2773,N_2500);
nor U5399 (N_5399,N_3130,N_3856);
nor U5400 (N_5400,N_3711,N_3361);
nand U5401 (N_5401,N_3063,N_2571);
nand U5402 (N_5402,N_2304,N_3079);
xor U5403 (N_5403,N_2805,N_3175);
and U5404 (N_5404,N_2621,N_3315);
nand U5405 (N_5405,N_2299,N_2881);
xor U5406 (N_5406,N_3601,N_2186);
nand U5407 (N_5407,N_3864,N_2313);
xnor U5408 (N_5408,N_3181,N_2566);
nand U5409 (N_5409,N_3102,N_2756);
or U5410 (N_5410,N_2254,N_2433);
and U5411 (N_5411,N_3223,N_3306);
and U5412 (N_5412,N_2360,N_2161);
nand U5413 (N_5413,N_2829,N_2625);
xnor U5414 (N_5414,N_2060,N_2666);
or U5415 (N_5415,N_3483,N_3496);
xor U5416 (N_5416,N_2633,N_2538);
nand U5417 (N_5417,N_2283,N_2207);
and U5418 (N_5418,N_2237,N_2785);
and U5419 (N_5419,N_3642,N_2393);
nor U5420 (N_5420,N_3863,N_3579);
and U5421 (N_5421,N_3911,N_3412);
and U5422 (N_5422,N_3337,N_3768);
or U5423 (N_5423,N_2078,N_3151);
nand U5424 (N_5424,N_2118,N_3153);
xor U5425 (N_5425,N_2136,N_3263);
and U5426 (N_5426,N_3751,N_2889);
xnor U5427 (N_5427,N_2018,N_3301);
nor U5428 (N_5428,N_3636,N_2929);
xor U5429 (N_5429,N_3547,N_2572);
nand U5430 (N_5430,N_3758,N_3774);
nand U5431 (N_5431,N_2774,N_3839);
nor U5432 (N_5432,N_2255,N_2093);
xor U5433 (N_5433,N_3092,N_3343);
or U5434 (N_5434,N_3302,N_3076);
nand U5435 (N_5435,N_2105,N_2575);
nor U5436 (N_5436,N_2527,N_3300);
xnor U5437 (N_5437,N_3665,N_3308);
and U5438 (N_5438,N_3008,N_3082);
nand U5439 (N_5439,N_3281,N_2619);
nand U5440 (N_5440,N_2722,N_2439);
nor U5441 (N_5441,N_3967,N_2405);
and U5442 (N_5442,N_2973,N_3235);
nor U5443 (N_5443,N_3732,N_3159);
xnor U5444 (N_5444,N_3638,N_2395);
nor U5445 (N_5445,N_2162,N_2243);
and U5446 (N_5446,N_2556,N_3508);
xor U5447 (N_5447,N_2754,N_2891);
xnor U5448 (N_5448,N_2983,N_2698);
xnor U5449 (N_5449,N_3382,N_3801);
nand U5450 (N_5450,N_3535,N_2672);
and U5451 (N_5451,N_2895,N_3061);
xor U5452 (N_5452,N_3053,N_2142);
and U5453 (N_5453,N_3649,N_3900);
or U5454 (N_5454,N_2500,N_3840);
nand U5455 (N_5455,N_2685,N_3961);
nor U5456 (N_5456,N_2061,N_3439);
and U5457 (N_5457,N_2799,N_3144);
nor U5458 (N_5458,N_3174,N_3106);
nand U5459 (N_5459,N_3118,N_3317);
nor U5460 (N_5460,N_3771,N_3897);
xnor U5461 (N_5461,N_3984,N_3949);
nand U5462 (N_5462,N_2363,N_2495);
nand U5463 (N_5463,N_2561,N_2851);
or U5464 (N_5464,N_2696,N_2888);
nand U5465 (N_5465,N_2173,N_2024);
nand U5466 (N_5466,N_3410,N_3731);
xnor U5467 (N_5467,N_3537,N_2419);
xnor U5468 (N_5468,N_2582,N_3989);
nand U5469 (N_5469,N_2774,N_3932);
nor U5470 (N_5470,N_2948,N_2132);
nor U5471 (N_5471,N_2618,N_3397);
nor U5472 (N_5472,N_3491,N_2368);
nor U5473 (N_5473,N_2816,N_3233);
or U5474 (N_5474,N_2091,N_3319);
nor U5475 (N_5475,N_2208,N_3715);
and U5476 (N_5476,N_2718,N_2222);
nand U5477 (N_5477,N_3808,N_3150);
nor U5478 (N_5478,N_2874,N_3562);
and U5479 (N_5479,N_2648,N_2988);
nand U5480 (N_5480,N_3019,N_2124);
nor U5481 (N_5481,N_3862,N_3602);
or U5482 (N_5482,N_3990,N_2220);
or U5483 (N_5483,N_3169,N_3805);
or U5484 (N_5484,N_3983,N_2671);
xnor U5485 (N_5485,N_2043,N_3913);
xnor U5486 (N_5486,N_2333,N_3544);
nor U5487 (N_5487,N_3819,N_2662);
nor U5488 (N_5488,N_2859,N_2959);
or U5489 (N_5489,N_3747,N_3645);
and U5490 (N_5490,N_2921,N_3562);
or U5491 (N_5491,N_3739,N_3587);
xor U5492 (N_5492,N_3558,N_2724);
or U5493 (N_5493,N_2485,N_3073);
xor U5494 (N_5494,N_3257,N_3198);
and U5495 (N_5495,N_3722,N_3589);
nor U5496 (N_5496,N_3220,N_2776);
nor U5497 (N_5497,N_3332,N_2207);
nor U5498 (N_5498,N_3847,N_2031);
or U5499 (N_5499,N_2075,N_3405);
nand U5500 (N_5500,N_2924,N_3153);
xnor U5501 (N_5501,N_3761,N_3444);
nor U5502 (N_5502,N_3744,N_2673);
xnor U5503 (N_5503,N_2530,N_3430);
or U5504 (N_5504,N_2642,N_2780);
nor U5505 (N_5505,N_2042,N_2379);
and U5506 (N_5506,N_3841,N_2100);
nor U5507 (N_5507,N_2703,N_3928);
nand U5508 (N_5508,N_3524,N_2897);
nand U5509 (N_5509,N_2309,N_2311);
nand U5510 (N_5510,N_2237,N_2184);
or U5511 (N_5511,N_2750,N_3393);
nor U5512 (N_5512,N_2777,N_2987);
xnor U5513 (N_5513,N_3671,N_2445);
nor U5514 (N_5514,N_2227,N_3589);
nor U5515 (N_5515,N_3609,N_2187);
nand U5516 (N_5516,N_2678,N_3254);
xor U5517 (N_5517,N_2119,N_2882);
or U5518 (N_5518,N_2924,N_3195);
nand U5519 (N_5519,N_2359,N_2040);
xor U5520 (N_5520,N_3589,N_2312);
and U5521 (N_5521,N_2962,N_2604);
nand U5522 (N_5522,N_3659,N_3930);
xor U5523 (N_5523,N_3111,N_3008);
nand U5524 (N_5524,N_3506,N_2813);
nor U5525 (N_5525,N_3740,N_3015);
and U5526 (N_5526,N_2172,N_2165);
and U5527 (N_5527,N_2838,N_3614);
and U5528 (N_5528,N_3556,N_3753);
or U5529 (N_5529,N_3162,N_3654);
or U5530 (N_5530,N_2863,N_2222);
xnor U5531 (N_5531,N_2124,N_3442);
xor U5532 (N_5532,N_2167,N_3760);
and U5533 (N_5533,N_2099,N_2301);
nor U5534 (N_5534,N_2183,N_2162);
or U5535 (N_5535,N_3887,N_2657);
and U5536 (N_5536,N_3644,N_3713);
or U5537 (N_5537,N_3487,N_2209);
nor U5538 (N_5538,N_2681,N_2067);
and U5539 (N_5539,N_2439,N_3346);
nand U5540 (N_5540,N_3912,N_3556);
and U5541 (N_5541,N_2421,N_2941);
or U5542 (N_5542,N_2808,N_2360);
and U5543 (N_5543,N_2390,N_2348);
nor U5544 (N_5544,N_2402,N_3322);
xor U5545 (N_5545,N_3773,N_2475);
xnor U5546 (N_5546,N_3343,N_3893);
and U5547 (N_5547,N_2825,N_2810);
nor U5548 (N_5548,N_3215,N_3502);
nand U5549 (N_5549,N_3545,N_3544);
and U5550 (N_5550,N_2086,N_3145);
nor U5551 (N_5551,N_2643,N_2368);
and U5552 (N_5552,N_3407,N_2214);
nand U5553 (N_5553,N_2574,N_3346);
nand U5554 (N_5554,N_2330,N_3066);
and U5555 (N_5555,N_3451,N_2407);
and U5556 (N_5556,N_3052,N_3214);
xnor U5557 (N_5557,N_2215,N_2282);
nor U5558 (N_5558,N_3901,N_2448);
nand U5559 (N_5559,N_3748,N_2235);
xor U5560 (N_5560,N_3970,N_2741);
xor U5561 (N_5561,N_2492,N_3718);
xnor U5562 (N_5562,N_3735,N_3215);
nand U5563 (N_5563,N_2422,N_2000);
nor U5564 (N_5564,N_2495,N_3734);
nand U5565 (N_5565,N_3387,N_2961);
or U5566 (N_5566,N_3592,N_3847);
nand U5567 (N_5567,N_3773,N_2710);
nor U5568 (N_5568,N_2629,N_2252);
or U5569 (N_5569,N_2225,N_2192);
and U5570 (N_5570,N_2346,N_3183);
xnor U5571 (N_5571,N_2283,N_3116);
nand U5572 (N_5572,N_2928,N_2871);
nor U5573 (N_5573,N_3334,N_2333);
xnor U5574 (N_5574,N_2459,N_3333);
xor U5575 (N_5575,N_2520,N_3595);
or U5576 (N_5576,N_2386,N_3894);
or U5577 (N_5577,N_3551,N_2959);
or U5578 (N_5578,N_2408,N_3240);
xnor U5579 (N_5579,N_3601,N_3829);
and U5580 (N_5580,N_3132,N_2177);
nor U5581 (N_5581,N_2675,N_3323);
xor U5582 (N_5582,N_3019,N_2805);
xor U5583 (N_5583,N_3476,N_3452);
or U5584 (N_5584,N_3252,N_3260);
nor U5585 (N_5585,N_3900,N_3020);
xnor U5586 (N_5586,N_2641,N_3208);
and U5587 (N_5587,N_3205,N_3111);
or U5588 (N_5588,N_3292,N_2785);
and U5589 (N_5589,N_3372,N_2270);
nor U5590 (N_5590,N_2196,N_3653);
nand U5591 (N_5591,N_3050,N_3489);
nand U5592 (N_5592,N_2468,N_2307);
and U5593 (N_5593,N_2539,N_2631);
nand U5594 (N_5594,N_2572,N_2733);
xnor U5595 (N_5595,N_3407,N_2804);
or U5596 (N_5596,N_2325,N_3661);
nor U5597 (N_5597,N_3697,N_2844);
xor U5598 (N_5598,N_3710,N_2858);
or U5599 (N_5599,N_2135,N_2871);
xnor U5600 (N_5600,N_3022,N_2788);
and U5601 (N_5601,N_3859,N_3696);
and U5602 (N_5602,N_2737,N_2377);
xnor U5603 (N_5603,N_2475,N_2158);
and U5604 (N_5604,N_2245,N_3649);
xnor U5605 (N_5605,N_3591,N_2129);
or U5606 (N_5606,N_2624,N_2330);
xor U5607 (N_5607,N_3890,N_2136);
nor U5608 (N_5608,N_2930,N_2412);
or U5609 (N_5609,N_2140,N_2580);
or U5610 (N_5610,N_3998,N_2055);
and U5611 (N_5611,N_2546,N_2450);
nor U5612 (N_5612,N_3633,N_3387);
nand U5613 (N_5613,N_3856,N_2462);
xnor U5614 (N_5614,N_3053,N_2776);
nor U5615 (N_5615,N_2726,N_2905);
nand U5616 (N_5616,N_2127,N_2596);
xnor U5617 (N_5617,N_3682,N_3936);
nor U5618 (N_5618,N_3734,N_2443);
nand U5619 (N_5619,N_3890,N_2123);
xnor U5620 (N_5620,N_3402,N_2028);
xnor U5621 (N_5621,N_2752,N_3037);
nand U5622 (N_5622,N_3606,N_3387);
and U5623 (N_5623,N_3622,N_3491);
nand U5624 (N_5624,N_2337,N_2483);
nor U5625 (N_5625,N_3822,N_2645);
xnor U5626 (N_5626,N_2491,N_3285);
and U5627 (N_5627,N_2196,N_2954);
nor U5628 (N_5628,N_2391,N_3639);
xnor U5629 (N_5629,N_3076,N_3696);
xnor U5630 (N_5630,N_2742,N_3937);
and U5631 (N_5631,N_2485,N_3803);
or U5632 (N_5632,N_2761,N_2450);
nor U5633 (N_5633,N_2409,N_2670);
or U5634 (N_5634,N_3518,N_2281);
or U5635 (N_5635,N_2069,N_2875);
or U5636 (N_5636,N_2885,N_3587);
xnor U5637 (N_5637,N_2704,N_3812);
or U5638 (N_5638,N_3584,N_3888);
nand U5639 (N_5639,N_2342,N_2650);
xnor U5640 (N_5640,N_2426,N_3093);
and U5641 (N_5641,N_3402,N_2230);
nand U5642 (N_5642,N_2929,N_3337);
nor U5643 (N_5643,N_2980,N_3052);
nand U5644 (N_5644,N_3754,N_2953);
xor U5645 (N_5645,N_3342,N_2420);
or U5646 (N_5646,N_2555,N_3124);
or U5647 (N_5647,N_2308,N_3566);
and U5648 (N_5648,N_3263,N_2203);
or U5649 (N_5649,N_3657,N_2889);
nand U5650 (N_5650,N_2550,N_3315);
or U5651 (N_5651,N_2870,N_3692);
or U5652 (N_5652,N_2129,N_2597);
nand U5653 (N_5653,N_3533,N_2888);
or U5654 (N_5654,N_2369,N_3259);
xor U5655 (N_5655,N_3773,N_3318);
xor U5656 (N_5656,N_2531,N_3748);
nor U5657 (N_5657,N_3972,N_2855);
and U5658 (N_5658,N_3200,N_2278);
and U5659 (N_5659,N_3852,N_2860);
and U5660 (N_5660,N_2806,N_2699);
and U5661 (N_5661,N_2898,N_3603);
or U5662 (N_5662,N_3788,N_2315);
nor U5663 (N_5663,N_3019,N_3955);
xnor U5664 (N_5664,N_2420,N_3425);
and U5665 (N_5665,N_3175,N_2872);
nor U5666 (N_5666,N_2714,N_2767);
or U5667 (N_5667,N_2542,N_2848);
nand U5668 (N_5668,N_2184,N_3297);
or U5669 (N_5669,N_2856,N_2397);
or U5670 (N_5670,N_3374,N_3221);
nor U5671 (N_5671,N_2807,N_3835);
nor U5672 (N_5672,N_3436,N_3437);
nand U5673 (N_5673,N_3329,N_3079);
or U5674 (N_5674,N_2467,N_3786);
nor U5675 (N_5675,N_2882,N_2082);
nor U5676 (N_5676,N_3004,N_2338);
or U5677 (N_5677,N_2344,N_3784);
or U5678 (N_5678,N_2957,N_3463);
or U5679 (N_5679,N_2348,N_2150);
or U5680 (N_5680,N_3482,N_3606);
and U5681 (N_5681,N_2119,N_3699);
or U5682 (N_5682,N_2301,N_3958);
or U5683 (N_5683,N_2725,N_2866);
xor U5684 (N_5684,N_2247,N_3837);
nor U5685 (N_5685,N_2705,N_3569);
xnor U5686 (N_5686,N_3682,N_2533);
nand U5687 (N_5687,N_2793,N_2788);
and U5688 (N_5688,N_3811,N_3178);
or U5689 (N_5689,N_2627,N_2047);
and U5690 (N_5690,N_2988,N_3331);
nor U5691 (N_5691,N_3475,N_3537);
xnor U5692 (N_5692,N_2253,N_2846);
or U5693 (N_5693,N_2337,N_2685);
nand U5694 (N_5694,N_3069,N_2970);
xor U5695 (N_5695,N_3651,N_2865);
or U5696 (N_5696,N_3647,N_2372);
xor U5697 (N_5697,N_2107,N_3469);
xor U5698 (N_5698,N_3544,N_2988);
and U5699 (N_5699,N_2647,N_2822);
xor U5700 (N_5700,N_2932,N_2710);
xnor U5701 (N_5701,N_2327,N_2379);
and U5702 (N_5702,N_3221,N_3810);
nand U5703 (N_5703,N_3497,N_3745);
nand U5704 (N_5704,N_2656,N_3643);
nor U5705 (N_5705,N_3892,N_2880);
and U5706 (N_5706,N_2505,N_3282);
nand U5707 (N_5707,N_2692,N_2364);
xnor U5708 (N_5708,N_2211,N_3740);
xor U5709 (N_5709,N_3262,N_3062);
or U5710 (N_5710,N_2449,N_3885);
xor U5711 (N_5711,N_3274,N_3087);
and U5712 (N_5712,N_3489,N_2030);
nand U5713 (N_5713,N_3703,N_2599);
xor U5714 (N_5714,N_2897,N_2869);
nor U5715 (N_5715,N_2644,N_3979);
and U5716 (N_5716,N_3303,N_3296);
or U5717 (N_5717,N_3072,N_3259);
nor U5718 (N_5718,N_2678,N_2521);
nand U5719 (N_5719,N_3844,N_2559);
xnor U5720 (N_5720,N_3051,N_3614);
xor U5721 (N_5721,N_2009,N_2710);
and U5722 (N_5722,N_3801,N_3501);
xor U5723 (N_5723,N_2660,N_2684);
nand U5724 (N_5724,N_3746,N_3553);
xnor U5725 (N_5725,N_2966,N_2231);
nor U5726 (N_5726,N_3673,N_3680);
xor U5727 (N_5727,N_3263,N_2592);
nand U5728 (N_5728,N_3824,N_3433);
and U5729 (N_5729,N_2039,N_2242);
nor U5730 (N_5730,N_2680,N_3113);
or U5731 (N_5731,N_3490,N_2578);
and U5732 (N_5732,N_2648,N_3559);
nand U5733 (N_5733,N_3747,N_3138);
nand U5734 (N_5734,N_3508,N_3587);
and U5735 (N_5735,N_3310,N_3021);
nor U5736 (N_5736,N_2137,N_2787);
xnor U5737 (N_5737,N_2024,N_2117);
xor U5738 (N_5738,N_3619,N_3175);
nor U5739 (N_5739,N_3728,N_2724);
nor U5740 (N_5740,N_2873,N_3712);
xnor U5741 (N_5741,N_3895,N_3931);
and U5742 (N_5742,N_3487,N_2168);
nor U5743 (N_5743,N_3069,N_2714);
and U5744 (N_5744,N_2277,N_2581);
nand U5745 (N_5745,N_3443,N_3789);
and U5746 (N_5746,N_2973,N_3854);
and U5747 (N_5747,N_2131,N_3958);
nand U5748 (N_5748,N_3466,N_2640);
xor U5749 (N_5749,N_3616,N_3639);
or U5750 (N_5750,N_2464,N_3481);
and U5751 (N_5751,N_2282,N_2513);
or U5752 (N_5752,N_3946,N_2722);
nor U5753 (N_5753,N_2396,N_2511);
and U5754 (N_5754,N_3114,N_2306);
and U5755 (N_5755,N_3331,N_2191);
nand U5756 (N_5756,N_3371,N_3287);
or U5757 (N_5757,N_3912,N_2779);
or U5758 (N_5758,N_3038,N_3469);
nand U5759 (N_5759,N_3228,N_3462);
and U5760 (N_5760,N_3560,N_2793);
and U5761 (N_5761,N_3613,N_2751);
and U5762 (N_5762,N_3225,N_2247);
nor U5763 (N_5763,N_3331,N_2162);
nand U5764 (N_5764,N_2455,N_3106);
nand U5765 (N_5765,N_2911,N_3415);
and U5766 (N_5766,N_3670,N_2667);
nor U5767 (N_5767,N_3810,N_3831);
or U5768 (N_5768,N_2308,N_2890);
or U5769 (N_5769,N_3335,N_3278);
or U5770 (N_5770,N_3954,N_3668);
or U5771 (N_5771,N_3749,N_3342);
and U5772 (N_5772,N_2962,N_2138);
and U5773 (N_5773,N_2737,N_2338);
nor U5774 (N_5774,N_3847,N_2311);
nand U5775 (N_5775,N_3021,N_3897);
nor U5776 (N_5776,N_2281,N_2713);
or U5777 (N_5777,N_2739,N_2713);
nor U5778 (N_5778,N_2976,N_2269);
or U5779 (N_5779,N_3815,N_3492);
nand U5780 (N_5780,N_3000,N_3183);
xor U5781 (N_5781,N_3081,N_3720);
nand U5782 (N_5782,N_2610,N_3098);
xor U5783 (N_5783,N_2286,N_3518);
nand U5784 (N_5784,N_3654,N_3703);
nand U5785 (N_5785,N_3475,N_2064);
nand U5786 (N_5786,N_3716,N_2217);
and U5787 (N_5787,N_3858,N_2550);
nand U5788 (N_5788,N_3794,N_3807);
nand U5789 (N_5789,N_2381,N_2661);
or U5790 (N_5790,N_3130,N_3612);
or U5791 (N_5791,N_3940,N_2581);
nand U5792 (N_5792,N_3758,N_2291);
and U5793 (N_5793,N_2920,N_2554);
nand U5794 (N_5794,N_2246,N_3457);
and U5795 (N_5795,N_2361,N_3164);
xor U5796 (N_5796,N_2852,N_3317);
or U5797 (N_5797,N_2006,N_3899);
nor U5798 (N_5798,N_3088,N_3721);
nor U5799 (N_5799,N_2365,N_2015);
nor U5800 (N_5800,N_3128,N_3297);
or U5801 (N_5801,N_2478,N_2745);
xor U5802 (N_5802,N_3355,N_3438);
nand U5803 (N_5803,N_2465,N_2081);
nand U5804 (N_5804,N_3046,N_2221);
xor U5805 (N_5805,N_3437,N_2393);
nand U5806 (N_5806,N_3089,N_2101);
or U5807 (N_5807,N_3240,N_3575);
xnor U5808 (N_5808,N_3136,N_2411);
xor U5809 (N_5809,N_2909,N_3754);
nand U5810 (N_5810,N_3022,N_3003);
or U5811 (N_5811,N_3967,N_2149);
or U5812 (N_5812,N_2076,N_3494);
and U5813 (N_5813,N_3663,N_3991);
nand U5814 (N_5814,N_3162,N_3257);
nand U5815 (N_5815,N_3901,N_3303);
nor U5816 (N_5816,N_3675,N_3069);
nor U5817 (N_5817,N_2585,N_3388);
xnor U5818 (N_5818,N_2640,N_2303);
and U5819 (N_5819,N_2918,N_2294);
xor U5820 (N_5820,N_2273,N_2475);
and U5821 (N_5821,N_3525,N_2249);
nor U5822 (N_5822,N_2015,N_2124);
xnor U5823 (N_5823,N_3318,N_3515);
nor U5824 (N_5824,N_3081,N_3521);
or U5825 (N_5825,N_3958,N_2582);
and U5826 (N_5826,N_3328,N_2028);
and U5827 (N_5827,N_3217,N_3315);
and U5828 (N_5828,N_2277,N_2023);
and U5829 (N_5829,N_2297,N_2617);
or U5830 (N_5830,N_2082,N_3611);
nand U5831 (N_5831,N_2004,N_3032);
nand U5832 (N_5832,N_2524,N_3560);
and U5833 (N_5833,N_3925,N_2626);
or U5834 (N_5834,N_2312,N_3185);
nor U5835 (N_5835,N_3950,N_2334);
xnor U5836 (N_5836,N_2613,N_3212);
nand U5837 (N_5837,N_2279,N_3992);
nand U5838 (N_5838,N_3382,N_2760);
nand U5839 (N_5839,N_3338,N_2320);
nor U5840 (N_5840,N_2065,N_2300);
nand U5841 (N_5841,N_3431,N_3810);
nor U5842 (N_5842,N_3528,N_3216);
and U5843 (N_5843,N_3985,N_3378);
or U5844 (N_5844,N_3627,N_2435);
and U5845 (N_5845,N_3076,N_3167);
or U5846 (N_5846,N_2771,N_2783);
xor U5847 (N_5847,N_3574,N_2153);
or U5848 (N_5848,N_2768,N_3987);
nor U5849 (N_5849,N_2753,N_3288);
nand U5850 (N_5850,N_2912,N_3241);
nand U5851 (N_5851,N_3716,N_2487);
xnor U5852 (N_5852,N_2531,N_3140);
or U5853 (N_5853,N_3154,N_3377);
nor U5854 (N_5854,N_2911,N_3919);
or U5855 (N_5855,N_2323,N_3226);
nand U5856 (N_5856,N_3826,N_3876);
or U5857 (N_5857,N_2872,N_2692);
or U5858 (N_5858,N_2327,N_2947);
nor U5859 (N_5859,N_3526,N_2934);
and U5860 (N_5860,N_2434,N_2073);
and U5861 (N_5861,N_2847,N_2683);
nor U5862 (N_5862,N_3114,N_3856);
or U5863 (N_5863,N_2512,N_3278);
or U5864 (N_5864,N_2759,N_2559);
nand U5865 (N_5865,N_2542,N_2114);
and U5866 (N_5866,N_3644,N_3832);
nand U5867 (N_5867,N_2348,N_3217);
nand U5868 (N_5868,N_2145,N_2673);
nand U5869 (N_5869,N_3760,N_3183);
and U5870 (N_5870,N_3947,N_3991);
and U5871 (N_5871,N_2195,N_3086);
or U5872 (N_5872,N_2012,N_3308);
nor U5873 (N_5873,N_3977,N_2753);
xor U5874 (N_5874,N_2968,N_3472);
or U5875 (N_5875,N_3675,N_2575);
or U5876 (N_5876,N_2810,N_3618);
or U5877 (N_5877,N_2313,N_3697);
nor U5878 (N_5878,N_3374,N_3680);
nor U5879 (N_5879,N_3612,N_3359);
and U5880 (N_5880,N_3170,N_3538);
nand U5881 (N_5881,N_2589,N_2361);
nand U5882 (N_5882,N_3916,N_3895);
xnor U5883 (N_5883,N_3613,N_2523);
nor U5884 (N_5884,N_2119,N_3408);
and U5885 (N_5885,N_2810,N_2016);
or U5886 (N_5886,N_2236,N_2919);
and U5887 (N_5887,N_3757,N_2587);
nor U5888 (N_5888,N_3479,N_3802);
nand U5889 (N_5889,N_2166,N_2213);
or U5890 (N_5890,N_2747,N_2085);
nand U5891 (N_5891,N_2170,N_3220);
or U5892 (N_5892,N_2752,N_3378);
nor U5893 (N_5893,N_2047,N_2163);
nand U5894 (N_5894,N_3518,N_2767);
or U5895 (N_5895,N_3363,N_2637);
xor U5896 (N_5896,N_3941,N_3225);
xor U5897 (N_5897,N_3081,N_3280);
nand U5898 (N_5898,N_2011,N_3122);
nand U5899 (N_5899,N_3514,N_2563);
nor U5900 (N_5900,N_3925,N_3229);
and U5901 (N_5901,N_2452,N_3727);
or U5902 (N_5902,N_2465,N_2262);
and U5903 (N_5903,N_3627,N_2287);
and U5904 (N_5904,N_3198,N_3909);
xnor U5905 (N_5905,N_3062,N_3375);
nand U5906 (N_5906,N_2684,N_3340);
xor U5907 (N_5907,N_3733,N_3022);
xor U5908 (N_5908,N_3746,N_2359);
xnor U5909 (N_5909,N_3995,N_3270);
and U5910 (N_5910,N_3074,N_3487);
or U5911 (N_5911,N_2998,N_3007);
nor U5912 (N_5912,N_2686,N_2141);
and U5913 (N_5913,N_2905,N_3293);
and U5914 (N_5914,N_2992,N_3323);
or U5915 (N_5915,N_2878,N_3265);
nand U5916 (N_5916,N_3348,N_2243);
xnor U5917 (N_5917,N_2912,N_3453);
nor U5918 (N_5918,N_2796,N_2308);
xor U5919 (N_5919,N_3120,N_3352);
or U5920 (N_5920,N_2668,N_2285);
or U5921 (N_5921,N_2636,N_3797);
and U5922 (N_5922,N_2812,N_2741);
nor U5923 (N_5923,N_2313,N_2711);
xnor U5924 (N_5924,N_3730,N_3370);
nand U5925 (N_5925,N_2916,N_2913);
or U5926 (N_5926,N_3671,N_2156);
nand U5927 (N_5927,N_2378,N_2879);
nand U5928 (N_5928,N_3772,N_3034);
nor U5929 (N_5929,N_3452,N_3970);
nor U5930 (N_5930,N_2836,N_2155);
nor U5931 (N_5931,N_3090,N_3137);
xor U5932 (N_5932,N_3758,N_2473);
and U5933 (N_5933,N_3336,N_2245);
xnor U5934 (N_5934,N_3203,N_2191);
nand U5935 (N_5935,N_2769,N_2456);
nor U5936 (N_5936,N_2974,N_2752);
xnor U5937 (N_5937,N_2788,N_2449);
or U5938 (N_5938,N_2754,N_2796);
nor U5939 (N_5939,N_2106,N_3220);
nor U5940 (N_5940,N_3350,N_2454);
and U5941 (N_5941,N_2405,N_2448);
and U5942 (N_5942,N_3623,N_2290);
nand U5943 (N_5943,N_2515,N_2977);
nor U5944 (N_5944,N_3736,N_3922);
nand U5945 (N_5945,N_3645,N_3249);
and U5946 (N_5946,N_3830,N_3922);
and U5947 (N_5947,N_2876,N_3166);
and U5948 (N_5948,N_3853,N_3551);
nand U5949 (N_5949,N_3804,N_3254);
nand U5950 (N_5950,N_2393,N_3707);
nand U5951 (N_5951,N_2588,N_3983);
and U5952 (N_5952,N_2368,N_2755);
or U5953 (N_5953,N_3208,N_3176);
and U5954 (N_5954,N_2791,N_3058);
and U5955 (N_5955,N_2003,N_2554);
nor U5956 (N_5956,N_3161,N_2488);
nor U5957 (N_5957,N_2454,N_3161);
nor U5958 (N_5958,N_2869,N_2032);
xnor U5959 (N_5959,N_3042,N_2265);
and U5960 (N_5960,N_2937,N_3483);
xor U5961 (N_5961,N_2389,N_3867);
xnor U5962 (N_5962,N_3319,N_3378);
or U5963 (N_5963,N_2693,N_3243);
nand U5964 (N_5964,N_2272,N_3478);
nand U5965 (N_5965,N_2572,N_2151);
or U5966 (N_5966,N_3936,N_2890);
nand U5967 (N_5967,N_2207,N_2272);
and U5968 (N_5968,N_2180,N_3228);
and U5969 (N_5969,N_3390,N_2344);
and U5970 (N_5970,N_2413,N_3455);
or U5971 (N_5971,N_2714,N_2916);
and U5972 (N_5972,N_3205,N_3481);
nand U5973 (N_5973,N_2116,N_2886);
and U5974 (N_5974,N_2918,N_3984);
or U5975 (N_5975,N_2902,N_3835);
nand U5976 (N_5976,N_2401,N_3165);
nand U5977 (N_5977,N_3407,N_3074);
nand U5978 (N_5978,N_2317,N_2374);
nor U5979 (N_5979,N_3752,N_2874);
xor U5980 (N_5980,N_3484,N_3456);
nand U5981 (N_5981,N_3665,N_3377);
or U5982 (N_5982,N_3468,N_2728);
or U5983 (N_5983,N_2624,N_3655);
xor U5984 (N_5984,N_2129,N_2486);
and U5985 (N_5985,N_3984,N_2015);
and U5986 (N_5986,N_2075,N_3247);
xnor U5987 (N_5987,N_3340,N_3297);
xnor U5988 (N_5988,N_3047,N_2243);
xnor U5989 (N_5989,N_2804,N_3645);
and U5990 (N_5990,N_3173,N_2868);
nand U5991 (N_5991,N_2740,N_3626);
and U5992 (N_5992,N_3515,N_3714);
nand U5993 (N_5993,N_3883,N_2723);
nand U5994 (N_5994,N_3981,N_3006);
xnor U5995 (N_5995,N_3849,N_2876);
xnor U5996 (N_5996,N_3554,N_3427);
nor U5997 (N_5997,N_3581,N_3273);
xor U5998 (N_5998,N_2396,N_3533);
or U5999 (N_5999,N_2507,N_2425);
and U6000 (N_6000,N_4685,N_5630);
or U6001 (N_6001,N_4547,N_4833);
nand U6002 (N_6002,N_5840,N_4933);
xnor U6003 (N_6003,N_4487,N_5400);
nor U6004 (N_6004,N_5151,N_4964);
nand U6005 (N_6005,N_5900,N_4045);
xnor U6006 (N_6006,N_5827,N_4407);
xor U6007 (N_6007,N_5516,N_4371);
nand U6008 (N_6008,N_4198,N_4086);
or U6009 (N_6009,N_5156,N_4908);
xnor U6010 (N_6010,N_4264,N_4281);
and U6011 (N_6011,N_5095,N_5925);
or U6012 (N_6012,N_4926,N_4605);
or U6013 (N_6013,N_5573,N_4728);
xor U6014 (N_6014,N_5668,N_4260);
nor U6015 (N_6015,N_4778,N_5339);
nor U6016 (N_6016,N_5950,N_5518);
nand U6017 (N_6017,N_4246,N_5568);
nand U6018 (N_6018,N_4994,N_4769);
xnor U6019 (N_6019,N_5493,N_5442);
nor U6020 (N_6020,N_5542,N_4135);
or U6021 (N_6021,N_4190,N_4340);
or U6022 (N_6022,N_4104,N_5012);
xor U6023 (N_6023,N_4739,N_4784);
and U6024 (N_6024,N_5055,N_4974);
and U6025 (N_6025,N_4834,N_5297);
or U6026 (N_6026,N_4044,N_5933);
nand U6027 (N_6027,N_5797,N_5579);
nand U6028 (N_6028,N_5533,N_4528);
nand U6029 (N_6029,N_4392,N_5713);
xor U6030 (N_6030,N_5642,N_4529);
and U6031 (N_6031,N_4727,N_5105);
and U6032 (N_6032,N_4654,N_4592);
nand U6033 (N_6033,N_5999,N_5547);
and U6034 (N_6034,N_4439,N_4201);
or U6035 (N_6035,N_5209,N_5629);
nor U6036 (N_6036,N_4178,N_5044);
and U6037 (N_6037,N_5779,N_5529);
xnor U6038 (N_6038,N_5766,N_5583);
and U6039 (N_6039,N_5238,N_5927);
and U6040 (N_6040,N_4912,N_4915);
xor U6041 (N_6041,N_5143,N_5316);
nand U6042 (N_6042,N_5009,N_5163);
nor U6043 (N_6043,N_5741,N_5490);
or U6044 (N_6044,N_4786,N_4851);
xnor U6045 (N_6045,N_4173,N_5689);
or U6046 (N_6046,N_4884,N_4875);
xnor U6047 (N_6047,N_5114,N_4212);
or U6048 (N_6048,N_5546,N_4127);
and U6049 (N_6049,N_5962,N_4537);
nand U6050 (N_6050,N_4386,N_4882);
nand U6051 (N_6051,N_4334,N_5102);
nand U6052 (N_6052,N_4269,N_4193);
nor U6053 (N_6053,N_4106,N_4085);
nor U6054 (N_6054,N_5708,N_4907);
xor U6055 (N_6055,N_4189,N_5716);
nand U6056 (N_6056,N_4686,N_4272);
or U6057 (N_6057,N_4634,N_5401);
or U6058 (N_6058,N_5116,N_4922);
nand U6059 (N_6059,N_4877,N_4549);
nand U6060 (N_6060,N_4606,N_5025);
xnor U6061 (N_6061,N_5157,N_4458);
or U6062 (N_6062,N_4620,N_5359);
or U6063 (N_6063,N_5463,N_5075);
and U6064 (N_6064,N_4467,N_5448);
nand U6065 (N_6065,N_4854,N_4338);
and U6066 (N_6066,N_4626,N_5455);
or U6067 (N_6067,N_5698,N_5755);
nand U6068 (N_6068,N_4098,N_5967);
and U6069 (N_6069,N_5084,N_5059);
nor U6070 (N_6070,N_4515,N_4586);
or U6071 (N_6071,N_5210,N_4496);
or U6072 (N_6072,N_5094,N_5253);
nor U6073 (N_6073,N_5386,N_5252);
and U6074 (N_6074,N_5117,N_4510);
xnor U6075 (N_6075,N_5406,N_5745);
and U6076 (N_6076,N_4229,N_4137);
nand U6077 (N_6077,N_4230,N_5544);
or U6078 (N_6078,N_4719,N_5736);
nor U6079 (N_6079,N_4871,N_4435);
nand U6080 (N_6080,N_5505,N_5483);
xor U6081 (N_6081,N_4545,N_4791);
or U6082 (N_6082,N_4289,N_5433);
xnor U6083 (N_6083,N_5378,N_5223);
nand U6084 (N_6084,N_5665,N_5219);
or U6085 (N_6085,N_5908,N_4103);
nand U6086 (N_6086,N_5902,N_4176);
nor U6087 (N_6087,N_5740,N_5302);
nor U6088 (N_6088,N_4368,N_4463);
nor U6089 (N_6089,N_5160,N_5144);
nand U6090 (N_6090,N_5130,N_4244);
or U6091 (N_6091,N_5977,N_5345);
xnor U6092 (N_6092,N_5416,N_4570);
or U6093 (N_6093,N_4992,N_4418);
xnor U6094 (N_6094,N_4355,N_5035);
or U6095 (N_6095,N_4763,N_5266);
and U6096 (N_6096,N_4188,N_5155);
nor U6097 (N_6097,N_5497,N_4629);
nand U6098 (N_6098,N_5732,N_4568);
or U6099 (N_6099,N_4777,N_5299);
nor U6100 (N_6100,N_5435,N_5487);
xor U6101 (N_6101,N_4931,N_4139);
or U6102 (N_6102,N_5717,N_4955);
xnor U6103 (N_6103,N_4141,N_4425);
nand U6104 (N_6104,N_5504,N_4682);
or U6105 (N_6105,N_4431,N_5301);
or U6106 (N_6106,N_4007,N_5992);
and U6107 (N_6107,N_4208,N_5470);
and U6108 (N_6108,N_5702,N_5964);
nand U6109 (N_6109,N_4358,N_4318);
and U6110 (N_6110,N_4258,N_4485);
or U6111 (N_6111,N_5306,N_4783);
or U6112 (N_6112,N_5567,N_5832);
nor U6113 (N_6113,N_5955,N_5620);
or U6114 (N_6114,N_5612,N_4548);
xnor U6115 (N_6115,N_4405,N_5054);
or U6116 (N_6116,N_5310,N_4416);
xor U6117 (N_6117,N_5888,N_4377);
xnor U6118 (N_6118,N_4718,N_4713);
nand U6119 (N_6119,N_5377,N_5217);
or U6120 (N_6120,N_5335,N_4319);
nand U6121 (N_6121,N_4857,N_4107);
or U6122 (N_6122,N_5672,N_5182);
nor U6123 (N_6123,N_4853,N_4025);
or U6124 (N_6124,N_4711,N_5936);
nand U6125 (N_6125,N_5246,N_4301);
and U6126 (N_6126,N_5051,N_5763);
and U6127 (N_6127,N_5334,N_5848);
nand U6128 (N_6128,N_4231,N_4238);
nor U6129 (N_6129,N_4813,N_5778);
nand U6130 (N_6130,N_4027,N_4034);
nor U6131 (N_6131,N_5821,N_4067);
nor U6132 (N_6132,N_5203,N_4333);
and U6133 (N_6133,N_5993,N_5753);
or U6134 (N_6134,N_5859,N_5861);
xor U6135 (N_6135,N_4696,N_5171);
nor U6136 (N_6136,N_4889,N_4112);
or U6137 (N_6137,N_4669,N_4914);
and U6138 (N_6138,N_4291,N_4140);
or U6139 (N_6139,N_5453,N_4966);
and U6140 (N_6140,N_5914,N_4437);
xnor U6141 (N_6141,N_5882,N_4949);
nor U6142 (N_6142,N_4636,N_5935);
nor U6143 (N_6143,N_4276,N_4113);
xnor U6144 (N_6144,N_4445,N_5756);
or U6145 (N_6145,N_5492,N_5699);
nand U6146 (N_6146,N_4808,N_5963);
nand U6147 (N_6147,N_4001,N_4670);
or U6148 (N_6148,N_4794,N_4109);
nor U6149 (N_6149,N_5752,N_4185);
xnor U6150 (N_6150,N_5920,N_5269);
and U6151 (N_6151,N_5363,N_5589);
and U6152 (N_6152,N_5013,N_5304);
or U6153 (N_6153,N_5618,N_4647);
or U6154 (N_6154,N_5479,N_5189);
or U6155 (N_6155,N_4998,N_4972);
or U6156 (N_6156,N_5053,N_4477);
nor U6157 (N_6157,N_5839,N_5564);
nor U6158 (N_6158,N_5198,N_4422);
and U6159 (N_6159,N_5196,N_5838);
xor U6160 (N_6160,N_4052,N_4401);
and U6161 (N_6161,N_4204,N_5293);
nor U6162 (N_6162,N_4183,N_4759);
or U6163 (N_6163,N_4115,N_5358);
and U6164 (N_6164,N_5481,N_5686);
or U6165 (N_6165,N_5909,N_4245);
and U6166 (N_6166,N_5016,N_4604);
nor U6167 (N_6167,N_4500,N_4699);
nand U6168 (N_6168,N_4345,N_5195);
xor U6169 (N_6169,N_4646,N_5785);
nand U6170 (N_6170,N_5636,N_4928);
and U6171 (N_6171,N_5405,N_5186);
and U6172 (N_6172,N_5343,N_4206);
and U6173 (N_6173,N_4664,N_4257);
and U6174 (N_6174,N_5083,N_4362);
or U6175 (N_6175,N_5853,N_5086);
and U6176 (N_6176,N_5657,N_5506);
nor U6177 (N_6177,N_5411,N_5362);
xor U6178 (N_6178,N_4677,N_4169);
nand U6179 (N_6179,N_4698,N_4285);
and U6180 (N_6180,N_4056,N_4880);
nand U6181 (N_6181,N_5872,N_5034);
nor U6182 (N_6182,N_4090,N_5747);
nand U6183 (N_6183,N_4476,N_5422);
or U6184 (N_6184,N_5805,N_4716);
xor U6185 (N_6185,N_4446,N_4822);
and U6186 (N_6186,N_5896,N_5691);
xnor U6187 (N_6187,N_5214,N_5558);
or U6188 (N_6188,N_4066,N_4038);
and U6189 (N_6189,N_4923,N_5773);
nand U6190 (N_6190,N_4232,N_4838);
and U6191 (N_6191,N_4388,N_4743);
nor U6192 (N_6192,N_5141,N_4436);
and U6193 (N_6193,N_4663,N_4890);
or U6194 (N_6194,N_4295,N_4217);
or U6195 (N_6195,N_4396,N_4280);
xnor U6196 (N_6196,N_4505,N_4290);
and U6197 (N_6197,N_5537,N_4651);
and U6198 (N_6198,N_5107,N_4251);
and U6199 (N_6199,N_5849,N_4965);
or U6200 (N_6200,N_4943,N_4200);
nor U6201 (N_6201,N_4424,N_4249);
xor U6202 (N_6202,N_4088,N_5011);
nor U6203 (N_6203,N_5330,N_5918);
and U6204 (N_6204,N_4748,N_5485);
or U6205 (N_6205,N_5289,N_5602);
nor U6206 (N_6206,N_5355,N_4132);
nand U6207 (N_6207,N_4765,N_4754);
and U6208 (N_6208,N_4643,N_5336);
or U6209 (N_6209,N_5447,N_5218);
xor U6210 (N_6210,N_5662,N_5065);
nand U6211 (N_6211,N_5477,N_4900);
and U6212 (N_6212,N_4999,N_4542);
or U6213 (N_6213,N_4835,N_5850);
nor U6214 (N_6214,N_5393,N_4414);
nor U6215 (N_6215,N_4638,N_5561);
and U6216 (N_6216,N_4665,N_5344);
nor U6217 (N_6217,N_4731,N_5278);
nor U6218 (N_6218,N_5553,N_4393);
xnor U6219 (N_6219,N_4522,N_4474);
nor U6220 (N_6220,N_5725,N_4509);
or U6221 (N_6221,N_5879,N_5890);
or U6222 (N_6222,N_4015,N_5600);
or U6223 (N_6223,N_5973,N_5525);
or U6224 (N_6224,N_5031,N_4785);
nand U6225 (N_6225,N_5284,N_5762);
nor U6226 (N_6226,N_4239,N_4552);
nor U6227 (N_6227,N_4453,N_4374);
or U6228 (N_6228,N_4741,N_4196);
xnor U6229 (N_6229,N_5231,N_4224);
nand U6230 (N_6230,N_5645,N_4325);
nand U6231 (N_6231,N_4062,N_4187);
or U6232 (N_6232,N_5027,N_5560);
xor U6233 (N_6233,N_4207,N_5443);
or U6234 (N_6234,N_5757,N_5260);
nand U6235 (N_6235,N_5010,N_4814);
xnor U6236 (N_6236,N_4541,N_5771);
xor U6237 (N_6237,N_4556,N_4473);
and U6238 (N_6238,N_5110,N_5775);
and U6239 (N_6239,N_5634,N_4611);
nor U6240 (N_6240,N_4951,N_5478);
and U6241 (N_6241,N_4790,N_5494);
and U6242 (N_6242,N_5193,N_4110);
nor U6243 (N_6243,N_5996,N_5658);
nor U6244 (N_6244,N_4901,N_5826);
or U6245 (N_6245,N_5421,N_4101);
and U6246 (N_6246,N_4945,N_4977);
and U6247 (N_6247,N_5710,N_4432);
nand U6248 (N_6248,N_4519,N_5104);
nand U6249 (N_6249,N_4958,N_5288);
nor U6250 (N_6250,N_4715,N_5413);
and U6251 (N_6251,N_5078,N_5818);
nor U6252 (N_6252,N_4693,N_4557);
nand U6253 (N_6253,N_4726,N_4956);
nor U6254 (N_6254,N_4560,N_4042);
or U6255 (N_6255,N_4162,N_5235);
and U6256 (N_6256,N_4421,N_4040);
nand U6257 (N_6257,N_5263,N_5910);
xor U6258 (N_6258,N_5975,N_4199);
xnor U6259 (N_6259,N_4271,N_4979);
and U6260 (N_6260,N_4600,N_5664);
xnor U6261 (N_6261,N_5707,N_4466);
nand U6262 (N_6262,N_4982,N_4893);
and U6263 (N_6263,N_5042,N_4029);
xnor U6264 (N_6264,N_5295,N_4740);
and U6265 (N_6265,N_4408,N_5201);
and U6266 (N_6266,N_4623,N_4501);
and U6267 (N_6267,N_4320,N_4910);
xnor U6268 (N_6268,N_5804,N_4582);
nand U6269 (N_6269,N_4511,N_5676);
or U6270 (N_6270,N_5387,N_4525);
xnor U6271 (N_6271,N_5396,N_4041);
nor U6272 (N_6272,N_5291,N_4482);
and U6273 (N_6273,N_4302,N_4216);
nor U6274 (N_6274,N_4717,N_4980);
xor U6275 (N_6275,N_5239,N_4483);
or U6276 (N_6276,N_4729,N_5990);
xor U6277 (N_6277,N_4166,N_4957);
or U6278 (N_6278,N_5709,N_5132);
nor U6279 (N_6279,N_5758,N_4402);
or U6280 (N_6280,N_4091,N_5161);
or U6281 (N_6281,N_5472,N_4228);
nand U6282 (N_6282,N_4761,N_4142);
or U6283 (N_6283,N_5751,N_5704);
or U6284 (N_6284,N_5430,N_4924);
xnor U6285 (N_6285,N_5551,N_4950);
and U6286 (N_6286,N_4802,N_5033);
nor U6287 (N_6287,N_4895,N_5081);
nor U6288 (N_6288,N_5581,N_4220);
nor U6289 (N_6289,N_4642,N_4387);
nor U6290 (N_6290,N_5491,N_5985);
xor U6291 (N_6291,N_4049,N_4680);
or U6292 (N_6292,N_5460,N_5320);
and U6293 (N_6293,N_4546,N_5646);
or U6294 (N_6294,N_5912,N_5966);
and U6295 (N_6295,N_4615,N_5526);
or U6296 (N_6296,N_5450,N_5412);
xnor U6297 (N_6297,N_4565,N_4495);
nor U6298 (N_6298,N_4180,N_5836);
nand U6299 (N_6299,N_5559,N_5326);
and U6300 (N_6300,N_5372,N_5842);
xor U6301 (N_6301,N_5509,N_4913);
xor U6302 (N_6302,N_4593,N_4259);
xor U6303 (N_6303,N_4911,N_4011);
and U6304 (N_6304,N_5532,N_4359);
xnor U6305 (N_6305,N_5347,N_4073);
and U6306 (N_6306,N_4841,N_4048);
xor U6307 (N_6307,N_4095,N_4607);
or U6308 (N_6308,N_5008,N_5585);
xnor U6309 (N_6309,N_5321,N_5425);
xor U6310 (N_6310,N_5591,N_5374);
and U6311 (N_6311,N_4028,N_4734);
and U6312 (N_6312,N_5724,N_5045);
and U6313 (N_6313,N_4478,N_5715);
xnor U6314 (N_6314,N_4266,N_4100);
xnor U6315 (N_6315,N_5830,N_5234);
xor U6316 (N_6316,N_5540,N_5886);
nand U6317 (N_6317,N_4283,N_5873);
nor U6318 (N_6318,N_5735,N_5714);
nand U6319 (N_6319,N_5983,N_5125);
nor U6320 (N_6320,N_4465,N_4869);
xor U6321 (N_6321,N_5122,N_4021);
xnor U6322 (N_6322,N_4591,N_5017);
or U6323 (N_6323,N_4404,N_5582);
xnor U6324 (N_6324,N_4554,N_5337);
xor U6325 (N_6325,N_5557,N_5770);
xor U6326 (N_6326,N_5048,N_4866);
and U6327 (N_6327,N_5801,N_4796);
and U6328 (N_6328,N_4344,N_4969);
nand U6329 (N_6329,N_5168,N_4918);
xnor U6330 (N_6330,N_4016,N_5329);
xor U6331 (N_6331,N_5375,N_4618);
and U6332 (N_6332,N_4504,N_4535);
xor U6333 (N_6333,N_5093,N_4179);
nor U6334 (N_6334,N_4197,N_5145);
and U6335 (N_6335,N_4097,N_5259);
nand U6336 (N_6336,N_4613,N_4614);
or U6337 (N_6337,N_5414,N_5808);
nand U6338 (N_6338,N_5651,N_5028);
nand U6339 (N_6339,N_5989,N_5580);
nand U6340 (N_6340,N_4781,N_4161);
and U6341 (N_6341,N_4250,N_5318);
and U6342 (N_6342,N_4307,N_4701);
or U6343 (N_6343,N_4897,N_5120);
and U6344 (N_6344,N_4017,N_4385);
xnor U6345 (N_6345,N_4703,N_4324);
xnor U6346 (N_6346,N_5594,N_4697);
nor U6347 (N_6347,N_4352,N_4572);
and U6348 (N_6348,N_4879,N_5719);
nand U6349 (N_6349,N_5759,N_4843);
and U6350 (N_6350,N_4215,N_4694);
or U6351 (N_6351,N_4809,N_4798);
xor U6352 (N_6352,N_4026,N_5420);
nor U6353 (N_6353,N_5474,N_4084);
or U6354 (N_6354,N_4375,N_4214);
xor U6355 (N_6355,N_5835,N_5865);
or U6356 (N_6356,N_5466,N_4036);
nand U6357 (N_6357,N_5674,N_5215);
and U6358 (N_6358,N_4054,N_5066);
nor U6359 (N_6359,N_4690,N_4348);
nand U6360 (N_6360,N_4633,N_4752);
xnor U6361 (N_6361,N_5984,N_4002);
nor U6362 (N_6362,N_4948,N_4273);
nand U6363 (N_6363,N_4534,N_4120);
xnor U6364 (N_6364,N_4148,N_4970);
nand U6365 (N_6365,N_4089,N_5515);
or U6366 (N_6366,N_4539,N_5641);
xor U6367 (N_6367,N_5669,N_5097);
xor U6368 (N_6368,N_4906,N_4248);
nand U6369 (N_6369,N_4990,N_5241);
and U6370 (N_6370,N_5074,N_5959);
xnor U6371 (N_6371,N_5325,N_5895);
and U6372 (N_6372,N_4080,N_5911);
nand U6373 (N_6373,N_5593,N_4793);
nand U6374 (N_6374,N_5670,N_5943);
nand U6375 (N_6375,N_5300,N_5368);
or U6376 (N_6376,N_4577,N_5987);
xnor U6377 (N_6377,N_4471,N_4673);
and U6378 (N_6378,N_4865,N_5242);
and U6379 (N_6379,N_5613,N_5124);
and U6380 (N_6380,N_4323,N_5931);
nand U6381 (N_6381,N_5111,N_5191);
and U6382 (N_6382,N_4806,N_4278);
nand U6383 (N_6383,N_5085,N_4288);
and U6384 (N_6384,N_4968,N_4886);
xor U6385 (N_6385,N_5695,N_5883);
and U6386 (N_6386,N_5251,N_4294);
nand U6387 (N_6387,N_5897,N_4013);
or U6388 (N_6388,N_5113,N_4624);
nand U6389 (N_6389,N_4346,N_5574);
xnor U6390 (N_6390,N_5774,N_5350);
xor U6391 (N_6391,N_4531,N_4354);
nand U6392 (N_6392,N_4807,N_4946);
or U6393 (N_6393,N_4448,N_5046);
nor U6394 (N_6394,N_5096,N_4497);
or U6395 (N_6395,N_4464,N_5857);
xnor U6396 (N_6396,N_5623,N_4668);
and U6397 (N_6397,N_4811,N_4508);
or U6398 (N_6398,N_4427,N_5891);
xnor U6399 (N_6399,N_4076,N_4942);
or U6400 (N_6400,N_4125,N_5200);
nand U6401 (N_6401,N_5624,N_4331);
or U6402 (N_6402,N_5528,N_4707);
and U6403 (N_6403,N_4705,N_4170);
xnor U6404 (N_6404,N_5367,N_4175);
or U6405 (N_6405,N_5001,N_5706);
and U6406 (N_6406,N_5489,N_5718);
xor U6407 (N_6407,N_4603,N_5183);
or U6408 (N_6408,N_5584,N_5180);
nor U6409 (N_6409,N_5440,N_5666);
nor U6410 (N_6410,N_4341,N_4064);
or U6411 (N_6411,N_5475,N_5469);
and U6412 (N_6412,N_4299,N_4929);
nor U6413 (N_6413,N_5614,N_5978);
nor U6414 (N_6414,N_5769,N_5795);
nand U6415 (N_6415,N_5852,N_5654);
xnor U6416 (N_6416,N_4369,N_5513);
nand U6417 (N_6417,N_5632,N_4632);
xor U6418 (N_6418,N_5998,N_4996);
nor U6419 (N_6419,N_5134,N_4051);
nor U6420 (N_6420,N_5680,N_5366);
and U6421 (N_6421,N_5471,N_4441);
nor U6422 (N_6422,N_4649,N_5633);
nand U6423 (N_6423,N_5726,N_4061);
or U6424 (N_6424,N_5468,N_5190);
nor U6425 (N_6425,N_4789,N_4389);
nand U6426 (N_6426,N_5968,N_5364);
nand U6427 (N_6427,N_5022,N_4019);
xor U6428 (N_6428,N_5205,N_4909);
nor U6429 (N_6429,N_4960,N_5794);
or U6430 (N_6430,N_4171,N_4057);
or U6431 (N_6431,N_5800,N_4681);
or U6432 (N_6432,N_4517,N_5159);
nand U6433 (N_6433,N_5949,N_4263);
nand U6434 (N_6434,N_4234,N_4018);
nand U6435 (N_6435,N_5225,N_5663);
nor U6436 (N_6436,N_5047,N_4608);
and U6437 (N_6437,N_5408,N_5994);
nor U6438 (N_6438,N_4075,N_5845);
nand U6439 (N_6439,N_4826,N_5701);
nand U6440 (N_6440,N_4033,N_4824);
and U6441 (N_6441,N_4700,N_4156);
and U6442 (N_6442,N_5870,N_5846);
nand U6443 (N_6443,N_4736,N_5554);
and U6444 (N_6444,N_4131,N_5637);
or U6445 (N_6445,N_4595,N_4502);
xor U6446 (N_6446,N_4845,N_5510);
and U6447 (N_6447,N_4203,N_5903);
nand U6448 (N_6448,N_4940,N_4578);
nand U6449 (N_6449,N_4818,N_4308);
nor U6450 (N_6450,N_5748,N_4286);
nor U6451 (N_6451,N_5207,N_4581);
nor U6452 (N_6452,N_5938,N_5913);
nand U6453 (N_6453,N_4653,N_5502);
nand U6454 (N_6454,N_5220,N_5029);
and U6455 (N_6455,N_4621,N_4768);
xnor U6456 (N_6456,N_5222,N_5459);
nand U6457 (N_6457,N_4082,N_5464);
xnor U6458 (N_6458,N_4138,N_4805);
or U6459 (N_6459,N_4395,N_4540);
or U6460 (N_6460,N_5322,N_5142);
nand U6461 (N_6461,N_4306,N_5820);
nor U6462 (N_6462,N_4255,N_4316);
nor U6463 (N_6463,N_4443,N_5930);
xnor U6464 (N_6464,N_5720,N_4390);
and U6465 (N_6465,N_5498,N_4210);
and U6466 (N_6466,N_5817,N_5254);
nor U6467 (N_6467,N_4312,N_5005);
or U6468 (N_6468,N_4714,N_4449);
nor U6469 (N_6469,N_5331,N_5184);
and U6470 (N_6470,N_5446,N_4233);
xor U6471 (N_6471,N_4671,N_5856);
nor U6472 (N_6472,N_4855,N_5939);
or U6473 (N_6473,N_5389,N_5941);
or U6474 (N_6474,N_4072,N_5877);
xnor U6475 (N_6475,N_4532,N_4413);
nor U6476 (N_6476,N_5399,N_4488);
nand U6477 (N_6477,N_5495,N_4297);
nand U6478 (N_6478,N_5893,N_4329);
nor U6479 (N_6479,N_5050,N_5728);
or U6480 (N_6480,N_4724,N_5772);
nand U6481 (N_6481,N_4506,N_4530);
nand U6482 (N_6482,N_5427,N_4708);
nand U6483 (N_6483,N_4394,N_5863);
and U6484 (N_6484,N_4792,N_5862);
nor U6485 (N_6485,N_4936,N_4160);
xor U6486 (N_6486,N_4859,N_5768);
or U6487 (N_6487,N_5965,N_5082);
or U6488 (N_6488,N_5743,N_4426);
nand U6489 (N_6489,N_5415,N_4486);
and U6490 (N_6490,N_5906,N_4253);
xnor U6491 (N_6491,N_4237,N_5373);
or U6492 (N_6492,N_5404,N_4265);
and U6493 (N_6493,N_4952,N_4891);
or U6494 (N_6494,N_4365,N_4887);
and U6495 (N_6495,N_5311,N_4666);
nor U6496 (N_6496,N_5154,N_4378);
and U6497 (N_6497,N_5486,N_5298);
xnor U6498 (N_6498,N_4573,N_4243);
and U6499 (N_6499,N_4235,N_4995);
or U6500 (N_6500,N_5361,N_4744);
nor U6501 (N_6501,N_4874,N_5898);
xor U6502 (N_6502,N_4679,N_4812);
nand U6503 (N_6503,N_5286,N_4118);
and U6504 (N_6504,N_5417,N_5398);
nand U6505 (N_6505,N_5928,N_5070);
xnor U6506 (N_6506,N_5402,N_5004);
nor U6507 (N_6507,N_4195,N_4779);
nor U6508 (N_6508,N_4683,N_5661);
nand U6509 (N_6509,N_5675,N_4020);
xor U6510 (N_6510,N_5851,N_5166);
xnor U6511 (N_6511,N_5652,N_5208);
and U6512 (N_6512,N_4973,N_4507);
and U6513 (N_6513,N_5454,N_5823);
nor U6514 (N_6514,N_4930,N_4584);
nand U6515 (N_6515,N_5960,N_5007);
nand U6516 (N_6516,N_4059,N_4799);
nor U6517 (N_6517,N_5106,N_5014);
nand U6518 (N_6518,N_5333,N_4971);
and U6519 (N_6519,N_5831,N_5940);
nor U6520 (N_6520,N_4356,N_5147);
nor U6521 (N_6521,N_5319,N_5601);
nor U6522 (N_6522,N_4839,N_5410);
xor U6523 (N_6523,N_4810,N_5431);
or U6524 (N_6524,N_4277,N_5426);
and U6525 (N_6525,N_5383,N_5970);
xnor U6526 (N_6526,N_4134,N_5128);
nor U6527 (N_6527,N_5000,N_5812);
or U6528 (N_6528,N_5784,N_4494);
nor U6529 (N_6529,N_5194,N_5566);
nor U6530 (N_6530,N_4347,N_4524);
and U6531 (N_6531,N_4934,N_5162);
xnor U6532 (N_6532,N_5881,N_5855);
or U6533 (N_6533,N_5605,N_5521);
or U6534 (N_6534,N_5227,N_4861);
xnor U6535 (N_6535,N_5265,N_5588);
nand U6536 (N_6536,N_4795,N_4400);
nand U6537 (N_6537,N_5626,N_5232);
or U6538 (N_6538,N_5101,N_4637);
and U6539 (N_6539,N_4984,N_4617);
and U6540 (N_6540,N_5060,N_4157);
and U6541 (N_6541,N_5250,N_4093);
and U6542 (N_6542,N_4339,N_5103);
and U6543 (N_6543,N_4223,N_5257);
xor U6544 (N_6544,N_5049,N_4981);
nand U6545 (N_6545,N_5737,N_4304);
xnor U6546 (N_6546,N_4143,N_4144);
nand U6547 (N_6547,N_5371,N_5866);
nor U6548 (N_6548,N_5780,N_4499);
nand U6549 (N_6549,N_5556,N_4840);
or U6550 (N_6550,N_5276,N_5436);
nand U6551 (N_6551,N_5531,N_5595);
or U6552 (N_6552,N_5204,N_5061);
nor U6553 (N_6553,N_5598,N_5867);
xnor U6554 (N_6554,N_4650,N_5248);
nand U6555 (N_6555,N_4321,N_5569);
xnor U6556 (N_6556,N_5500,N_4292);
and U6557 (N_6557,N_5749,N_5535);
nor U6558 (N_6558,N_5187,N_5874);
nand U6559 (N_6559,N_5380,N_5790);
and U6560 (N_6560,N_5981,N_4240);
nor U6561 (N_6561,N_4450,N_5997);
and U6562 (N_6562,N_4576,N_5236);
and U6563 (N_6563,N_4151,N_4360);
xnor U6564 (N_6564,N_4797,N_5268);
nand U6565 (N_6565,N_5439,N_5843);
and U6566 (N_6566,N_4154,N_4932);
and U6567 (N_6567,N_5575,N_5064);
or U6568 (N_6568,N_5230,N_4518);
or U6569 (N_6569,N_4723,N_5871);
nand U6570 (N_6570,N_4309,N_4514);
nor U6571 (N_6571,N_4764,N_5348);
and U6572 (N_6572,N_4721,N_4848);
nor U6573 (N_6573,N_5980,N_4447);
or U6574 (N_6574,N_5847,N_4167);
nand U6575 (N_6575,N_4594,N_5727);
nand U6576 (N_6576,N_4881,N_5294);
nor U6577 (N_6577,N_4163,N_5381);
and U6578 (N_6578,N_5791,N_4599);
xor U6579 (N_6579,N_5199,N_5555);
and U6580 (N_6580,N_4772,N_4489);
or U6581 (N_6581,N_4397,N_5834);
or U6582 (N_6582,N_4122,N_4124);
or U6583 (N_6583,N_5841,N_5062);
nor U6584 (N_6584,N_5901,N_5764);
and U6585 (N_6585,N_4738,N_4850);
xnor U6586 (N_6586,N_5948,N_5409);
nor U6587 (N_6587,N_5428,N_4702);
nor U6588 (N_6588,N_5653,N_5305);
or U6589 (N_6589,N_5229,N_5255);
nor U6590 (N_6590,N_5961,N_4755);
or U6591 (N_6591,N_4878,N_4872);
nor U6592 (N_6592,N_4762,N_4335);
xor U6593 (N_6593,N_5261,N_4684);
nor U6594 (N_6594,N_4108,N_4361);
nor U6595 (N_6595,N_4712,N_4094);
nor U6596 (N_6596,N_4674,N_4588);
and U6597 (N_6597,N_4876,N_5945);
xor U6598 (N_6598,N_4211,N_4800);
nand U6599 (N_6599,N_4566,N_4380);
xnor U6600 (N_6600,N_5894,N_5150);
or U6601 (N_6601,N_5622,N_5731);
nand U6602 (N_6602,N_5211,N_5810);
or U6603 (N_6603,N_4442,N_5550);
nand U6604 (N_6604,N_5233,N_4083);
xnor U6605 (N_6605,N_4503,N_4689);
xnor U6606 (N_6606,N_5137,N_4481);
xor U6607 (N_6607,N_4986,N_4691);
xor U6608 (N_6608,N_5919,N_4438);
xnor U6609 (N_6609,N_5824,N_4117);
and U6610 (N_6610,N_5971,N_4152);
nor U6611 (N_6611,N_5690,N_5352);
nor U6612 (N_6612,N_4455,N_4720);
or U6613 (N_6613,N_4310,N_4722);
nor U6614 (N_6614,N_4213,N_4863);
nor U6615 (N_6615,N_5677,N_4429);
or U6616 (N_6616,N_5667,N_4904);
or U6617 (N_6617,N_4558,N_5991);
nor U6618 (N_6618,N_5905,N_5792);
nor U6619 (N_6619,N_5828,N_4533);
nand U6620 (N_6620,N_4370,N_5721);
xor U6621 (N_6621,N_5512,N_5173);
xor U6622 (N_6622,N_4096,N_5520);
xor U6623 (N_6623,N_5315,N_5814);
or U6624 (N_6624,N_5733,N_5597);
nor U6625 (N_6625,N_5822,N_4567);
nand U6626 (N_6626,N_5212,N_4959);
nand U6627 (N_6627,N_4937,N_5880);
xnor U6628 (N_6628,N_4336,N_5552);
nor U6629 (N_6629,N_4756,N_4675);
nor U6630 (N_6630,N_5036,N_4384);
and U6631 (N_6631,N_4836,N_5603);
or U6632 (N_6632,N_5392,N_4648);
xnor U6633 (N_6633,N_4284,N_5815);
and U6634 (N_6634,N_5638,N_4074);
nor U6635 (N_6635,N_5287,N_4953);
nand U6636 (N_6636,N_4459,N_5659);
xor U6637 (N_6637,N_5767,N_4658);
nor U6638 (N_6638,N_5307,N_5279);
or U6639 (N_6639,N_5324,N_4619);
or U6640 (N_6640,N_5148,N_4825);
or U6641 (N_6641,N_5712,N_5327);
and U6642 (N_6642,N_4692,N_4351);
xor U6643 (N_6643,N_5807,N_4662);
xor U6644 (N_6644,N_4268,N_4527);
nor U6645 (N_6645,N_4128,N_4031);
or U6646 (N_6646,N_4381,N_5176);
nand U6647 (N_6647,N_5953,N_4043);
or U6648 (N_6648,N_4725,N_5296);
nand U6649 (N_6649,N_5979,N_5969);
nand U6650 (N_6650,N_4564,N_5037);
and U6651 (N_6651,N_4944,N_5876);
and U6652 (N_6652,N_5273,N_4366);
or U6653 (N_6653,N_5649,N_5249);
nor U6654 (N_6654,N_5247,N_4667);
and U6655 (N_6655,N_4186,N_4430);
and U6656 (N_6656,N_5384,N_4296);
nand U6657 (N_6657,N_4829,N_5346);
nand U6658 (N_6658,N_5369,N_4627);
or U6659 (N_6659,N_5100,N_5837);
or U6660 (N_6660,N_4241,N_5711);
or U6661 (N_6661,N_5032,N_4192);
or U6662 (N_6662,N_5015,N_5577);
xnor U6663 (N_6663,N_5467,N_5829);
nor U6664 (N_6664,N_5484,N_5610);
or U6665 (N_6665,N_4423,N_5108);
nor U6666 (N_6666,N_4856,N_5077);
or U6667 (N_6667,N_5332,N_4279);
nor U6668 (N_6668,N_4780,N_5365);
xnor U6669 (N_6669,N_5281,N_4750);
nand U6670 (N_6670,N_5499,N_4287);
nor U6671 (N_6671,N_4939,N_5648);
and U6672 (N_6672,N_5178,N_5738);
and U6673 (N_6673,N_4597,N_5951);
nand U6674 (N_6674,N_4155,N_5854);
or U6675 (N_6675,N_4864,N_5576);
xnor U6676 (N_6676,N_4129,N_5360);
nor U6677 (N_6677,N_4159,N_5693);
and U6678 (N_6678,N_4732,N_4475);
nor U6679 (N_6679,N_5403,N_5274);
nor U6680 (N_6680,N_4610,N_4444);
xor U6681 (N_6681,N_5524,N_5734);
nor U6682 (N_6682,N_4962,N_5615);
or U6683 (N_6683,N_5258,N_5119);
and U6684 (N_6684,N_5860,N_4469);
xor U6685 (N_6685,N_4920,N_5813);
nor U6686 (N_6686,N_4538,N_5179);
nor U6687 (N_6687,N_5974,N_4282);
nor U6688 (N_6688,N_4657,N_5889);
nor U6689 (N_6689,N_5146,N_5213);
nand U6690 (N_6690,N_5181,N_4164);
or U6691 (N_6691,N_4417,N_4218);
nor U6692 (N_6692,N_4559,N_4079);
and U6693 (N_6693,N_5844,N_5946);
or U6694 (N_6694,N_5115,N_5099);
xnor U6695 (N_6695,N_5271,N_5019);
or U6696 (N_6696,N_5744,N_5240);
or U6697 (N_6697,N_4461,N_4219);
or U6698 (N_6698,N_4640,N_5609);
nand U6699 (N_6699,N_4363,N_4008);
xnor U6700 (N_6700,N_5884,N_4069);
nand U6701 (N_6701,N_4571,N_5617);
or U6702 (N_6702,N_5394,N_4536);
xnor U6703 (N_6703,N_4905,N_5165);
and U6704 (N_6704,N_4315,N_5501);
or U6705 (N_6705,N_4804,N_5309);
or U6706 (N_6706,N_4349,N_4523);
nor U6707 (N_6707,N_4006,N_4168);
nand U6708 (N_6708,N_5904,N_5003);
and U6709 (N_6709,N_4938,N_4815);
and U6710 (N_6710,N_4376,N_4782);
nor U6711 (N_6711,N_4883,N_5140);
and U6712 (N_6712,N_4849,N_5158);
or U6713 (N_6713,N_4460,N_5761);
or U6714 (N_6714,N_4326,N_4867);
nor U6715 (N_6715,N_5328,N_5354);
and U6716 (N_6716,N_5314,N_5067);
or U6717 (N_6717,N_4773,N_4520);
nand U6718 (N_6718,N_4561,N_5068);
and U6719 (N_6719,N_5127,N_5292);
xor U6720 (N_6720,N_4660,N_5152);
or U6721 (N_6721,N_4337,N_4526);
and U6722 (N_6722,N_5391,N_4892);
xnor U6723 (N_6723,N_5536,N_4695);
or U6724 (N_6724,N_4622,N_4434);
nor U6725 (N_6725,N_5655,N_4121);
and U6726 (N_6726,N_5892,N_5957);
nand U6727 (N_6727,N_5673,N_5370);
and U6728 (N_6728,N_5833,N_4641);
nor U6729 (N_6729,N_4050,N_4462);
xor U6730 (N_6730,N_5090,N_4925);
nor U6731 (N_6731,N_5072,N_5275);
xnor U6732 (N_6732,N_5563,N_5868);
nand U6733 (N_6733,N_4870,N_5461);
and U6734 (N_6734,N_5424,N_4860);
nand U6735 (N_6735,N_4314,N_4873);
or U6736 (N_6736,N_5202,N_5647);
xnor U6737 (N_6737,N_5917,N_4111);
xor U6738 (N_6738,N_4470,N_5924);
nand U6739 (N_6739,N_5277,N_5538);
xnor U6740 (N_6740,N_5786,N_5080);
and U6741 (N_6741,N_5002,N_5058);
nand U6742 (N_6742,N_5644,N_5480);
or U6743 (N_6743,N_4709,N_5806);
and U6744 (N_6744,N_4226,N_5237);
nor U6745 (N_6745,N_5088,N_5308);
nor U6746 (N_6746,N_5923,N_4024);
xnor U6747 (N_6747,N_5696,N_5226);
nor U6748 (N_6748,N_4544,N_4078);
nand U6749 (N_6749,N_5816,N_5592);
nor U6750 (N_6750,N_5682,N_5341);
nor U6751 (N_6751,N_5071,N_4921);
nand U6752 (N_6752,N_4583,N_4555);
and U6753 (N_6753,N_5548,N_5079);
nor U6754 (N_6754,N_4635,N_4512);
xnor U6755 (N_6755,N_4035,N_4774);
and U6756 (N_6756,N_4379,N_4630);
xnor U6757 (N_6757,N_5507,N_5599);
xnor U6758 (N_6758,N_5452,N_4997);
or U6759 (N_6759,N_4710,N_5723);
xor U6760 (N_6760,N_4428,N_4898);
nand U6761 (N_6761,N_5811,N_5787);
or U6762 (N_6762,N_4105,N_4490);
and U6763 (N_6763,N_5549,N_5730);
and U6764 (N_6764,N_5739,N_5129);
and U6765 (N_6765,N_4830,N_4888);
xnor U6766 (N_6766,N_4551,N_5256);
xor U6767 (N_6767,N_5131,N_4801);
or U6768 (N_6768,N_4454,N_5606);
nand U6769 (N_6769,N_4330,N_4659);
or U6770 (N_6770,N_5089,N_5388);
and U6771 (N_6771,N_5136,N_4274);
xor U6772 (N_6772,N_5476,N_5684);
xnor U6773 (N_6773,N_5026,N_4644);
or U6774 (N_6774,N_4771,N_4313);
nand U6775 (N_6775,N_5519,N_4037);
nand U6776 (N_6776,N_4899,N_5228);
xnor U6777 (N_6777,N_5091,N_4065);
and U6778 (N_6778,N_4569,N_5174);
nand U6779 (N_6779,N_5098,N_5451);
nand U6780 (N_6780,N_5449,N_4403);
nand U6781 (N_6781,N_4327,N_5175);
and U6782 (N_6782,N_5995,N_4989);
xnor U6783 (N_6783,N_4181,N_5508);
xnor U6784 (N_6784,N_5534,N_4409);
nor U6785 (N_6785,N_4753,N_4885);
nor U6786 (N_6786,N_4433,N_4828);
xor U6787 (N_6787,N_4844,N_5541);
xnor U6788 (N_6788,N_5397,N_5224);
nand U6789 (N_6789,N_4553,N_5496);
and U6790 (N_6790,N_5621,N_5465);
xor U6791 (N_6791,N_5562,N_5121);
nor U6792 (N_6792,N_5687,N_5023);
nand U6793 (N_6793,N_4976,N_5216);
or U6794 (N_6794,N_4975,N_4757);
nand U6795 (N_6795,N_5976,N_5869);
xor U6796 (N_6796,N_5809,N_4262);
xnor U6797 (N_6797,N_4656,N_4254);
and U6798 (N_6798,N_5915,N_5958);
and U6799 (N_6799,N_5503,N_4412);
and U6800 (N_6800,N_4823,N_5750);
and U6801 (N_6801,N_5020,N_4935);
xnor U6802 (N_6802,N_5264,N_5429);
nand U6803 (N_6803,N_5376,N_4574);
and U6804 (N_6804,N_4411,N_4256);
or U6805 (N_6805,N_5760,N_4837);
nand U6806 (N_6806,N_4816,N_5407);
nand U6807 (N_6807,N_4221,N_4150);
nand U6808 (N_6808,N_5462,N_4063);
nor U6809 (N_6809,N_5607,N_5522);
or U6810 (N_6810,N_4983,N_5887);
and U6811 (N_6811,N_4172,N_4242);
nor U6812 (N_6812,N_5112,N_5858);
and U6813 (N_6813,N_4009,N_5611);
or U6814 (N_6814,N_5514,N_4492);
nor U6815 (N_6815,N_4587,N_5458);
xor U6816 (N_6816,N_5030,N_4896);
or U6817 (N_6817,N_4060,N_4457);
and U6818 (N_6818,N_5018,N_5656);
nor U6819 (N_6819,N_4222,N_4087);
xor U6820 (N_6820,N_4580,N_4730);
xor U6821 (N_6821,N_5685,N_4760);
and U6822 (N_6822,N_4751,N_5153);
xor U6823 (N_6823,N_4733,N_5631);
xnor U6824 (N_6824,N_5280,N_4770);
or U6825 (N_6825,N_5063,N_5885);
nor U6826 (N_6826,N_5683,N_4126);
xnor U6827 (N_6827,N_5527,N_5342);
nand U6828 (N_6828,N_5937,N_5052);
and U6829 (N_6829,N_4988,N_4133);
and U6830 (N_6830,N_4858,N_4563);
nand U6831 (N_6831,N_5285,N_5705);
or U6832 (N_6832,N_4452,N_5069);
nor U6833 (N_6833,N_4468,N_4382);
xor U6834 (N_6834,N_4842,N_5922);
and U6835 (N_6835,N_4236,N_4961);
nor U6836 (N_6836,N_4406,N_5530);
and U6837 (N_6837,N_4493,N_5473);
or U6838 (N_6838,N_5076,N_4032);
and U6839 (N_6839,N_5572,N_4672);
xor U6840 (N_6840,N_4575,N_5799);
xnor U6841 (N_6841,N_4364,N_5385);
nand U6842 (N_6842,N_4317,N_4655);
and U6843 (N_6843,N_5942,N_4704);
or U6844 (N_6844,N_5056,N_4903);
or U6845 (N_6845,N_5185,N_5282);
nor U6846 (N_6846,N_5627,N_5006);
nand U6847 (N_6847,N_5628,N_5742);
and U6848 (N_6848,N_4202,N_4114);
and U6849 (N_6849,N_5135,N_4985);
and U6850 (N_6850,N_5926,N_4598);
and U6851 (N_6851,N_4941,N_5244);
xor U6852 (N_6852,N_5283,N_4550);
or U6853 (N_6853,N_4012,N_5243);
nor U6854 (N_6854,N_5640,N_4817);
nor U6855 (N_6855,N_5188,N_4332);
nand U6856 (N_6856,N_5206,N_4055);
nand U6857 (N_6857,N_4513,N_4343);
or U6858 (N_6858,N_5565,N_5608);
nor U6859 (N_6859,N_5972,N_4676);
and U6860 (N_6860,N_4182,N_4261);
and U6861 (N_6861,N_5671,N_5349);
nand U6862 (N_6862,N_5746,N_5444);
and U6863 (N_6863,N_4631,N_4123);
nor U6864 (N_6864,N_5793,N_5312);
xor U6865 (N_6865,N_5571,N_5643);
and U6866 (N_6866,N_5092,N_5688);
xnor U6867 (N_6867,N_4967,N_4303);
xnor U6868 (N_6868,N_4005,N_4399);
xor U6869 (N_6869,N_5545,N_4687);
or U6870 (N_6870,N_4645,N_5457);
and U6871 (N_6871,N_5788,N_4585);
or U6872 (N_6872,N_5262,N_4917);
nand U6873 (N_6873,N_4058,N_5038);
and U6874 (N_6874,N_5697,N_4149);
nor U6875 (N_6875,N_5139,N_5678);
nor U6876 (N_6876,N_5650,N_4158);
or U6877 (N_6877,N_4491,N_4119);
or U6878 (N_6878,N_5126,N_4737);
nor U6879 (N_6879,N_4398,N_5351);
nor U6880 (N_6880,N_4827,N_5303);
xor U6881 (N_6881,N_5523,N_4609);
nand U6882 (N_6882,N_5290,N_5781);
and U6883 (N_6883,N_4628,N_4868);
nand U6884 (N_6884,N_4821,N_5982);
xor U6885 (N_6885,N_5177,N_4688);
nor U6886 (N_6886,N_5432,N_4003);
nor U6887 (N_6887,N_4225,N_4472);
nor U6888 (N_6888,N_5353,N_5379);
nand U6889 (N_6889,N_5133,N_4820);
nor U6890 (N_6890,N_4146,N_5907);
nor U6891 (N_6891,N_5798,N_4267);
xnor U6892 (N_6892,N_4978,N_4102);
nand U6893 (N_6893,N_4745,N_5317);
or U6894 (N_6894,N_4293,N_4184);
and U6895 (N_6895,N_4602,N_4596);
xnor U6896 (N_6896,N_4562,N_4022);
or U6897 (N_6897,N_5916,N_4787);
nor U6898 (N_6898,N_5021,N_5356);
and U6899 (N_6899,N_5272,N_5382);
nor U6900 (N_6900,N_4415,N_4070);
nor U6901 (N_6901,N_4322,N_5694);
nor U6902 (N_6902,N_4862,N_5123);
nor U6903 (N_6903,N_4919,N_5517);
nor U6904 (N_6904,N_5073,N_5170);
nor U6905 (N_6905,N_4372,N_4030);
xor U6906 (N_6906,N_4145,N_5952);
and U6907 (N_6907,N_5043,N_4543);
and U6908 (N_6908,N_4579,N_4616);
or U6909 (N_6909,N_4136,N_5419);
nand U6910 (N_6910,N_4735,N_4357);
nand U6911 (N_6911,N_5511,N_4894);
xor U6912 (N_6912,N_4270,N_5221);
and U6913 (N_6913,N_4071,N_4410);
nor U6914 (N_6914,N_4373,N_5878);
or U6915 (N_6915,N_4947,N_5149);
xnor U6916 (N_6916,N_4747,N_5041);
xnor U6917 (N_6917,N_4902,N_4000);
xnor U6918 (N_6918,N_5482,N_5986);
and U6919 (N_6919,N_4010,N_5456);
nand U6920 (N_6920,N_4014,N_4311);
nor U6921 (N_6921,N_5783,N_4068);
nand U6922 (N_6922,N_4153,N_5988);
xor U6923 (N_6923,N_5825,N_4046);
or U6924 (N_6924,N_4832,N_5754);
or U6925 (N_6925,N_4954,N_5899);
xnor U6926 (N_6926,N_5323,N_5722);
and U6927 (N_6927,N_4652,N_4081);
nand U6928 (N_6928,N_4767,N_5057);
nand U6929 (N_6929,N_4803,N_5635);
nand U6930 (N_6930,N_5437,N_4987);
nor U6931 (N_6931,N_4353,N_4004);
nor U6932 (N_6932,N_4479,N_4039);
and U6933 (N_6933,N_4147,N_5438);
nand U6934 (N_6934,N_4788,N_5864);
or U6935 (N_6935,N_4391,N_5167);
or U6936 (N_6936,N_5782,N_4589);
xnor U6937 (N_6937,N_5947,N_5340);
or U6938 (N_6938,N_4639,N_5729);
nand U6939 (N_6939,N_4516,N_4227);
or U6940 (N_6940,N_5418,N_4456);
and U6941 (N_6941,N_4498,N_4746);
nand U6942 (N_6942,N_4749,N_4130);
nor U6943 (N_6943,N_5172,N_5578);
xor U6944 (N_6944,N_4766,N_5586);
nor U6945 (N_6945,N_4847,N_4775);
and U6946 (N_6946,N_4991,N_4484);
or U6947 (N_6947,N_4275,N_5776);
nand U6948 (N_6948,N_4963,N_5875);
and U6949 (N_6949,N_5934,N_5660);
or U6950 (N_6950,N_4350,N_5118);
or U6951 (N_6951,N_4116,N_4993);
and U6952 (N_6952,N_4053,N_4023);
xor U6953 (N_6953,N_4678,N_4047);
nor U6954 (N_6954,N_5039,N_5803);
or U6955 (N_6955,N_4077,N_5789);
or U6956 (N_6956,N_4191,N_5040);
and U6957 (N_6957,N_5164,N_5596);
xnor U6958 (N_6958,N_4383,N_4367);
or U6959 (N_6959,N_4205,N_4092);
or U6960 (N_6960,N_5616,N_5169);
and U6961 (N_6961,N_5639,N_4298);
or U6962 (N_6962,N_5929,N_4420);
nand U6963 (N_6963,N_5932,N_4419);
xor U6964 (N_6964,N_5703,N_4521);
nor U6965 (N_6965,N_4342,N_5700);
nor U6966 (N_6966,N_4209,N_5313);
nand U6967 (N_6967,N_4099,N_5625);
and U6968 (N_6968,N_5087,N_5270);
nand U6969 (N_6969,N_4819,N_5434);
or U6970 (N_6970,N_4758,N_4846);
nand U6971 (N_6971,N_4451,N_4612);
xnor U6972 (N_6972,N_5944,N_4165);
or U6973 (N_6973,N_4300,N_5765);
nor U6974 (N_6974,N_5681,N_5802);
xor U6975 (N_6975,N_4831,N_4927);
xor U6976 (N_6976,N_4177,N_4328);
nand U6977 (N_6977,N_5604,N_5395);
xor U6978 (N_6978,N_4194,N_5587);
xor U6979 (N_6979,N_4174,N_5488);
nand U6980 (N_6980,N_5245,N_5543);
nor U6981 (N_6981,N_5109,N_5796);
nand U6982 (N_6982,N_5777,N_4601);
and U6983 (N_6983,N_5539,N_5619);
or U6984 (N_6984,N_5921,N_4852);
or U6985 (N_6985,N_4590,N_5024);
or U6986 (N_6986,N_5590,N_5423);
and U6987 (N_6987,N_5570,N_5441);
xnor U6988 (N_6988,N_4776,N_4706);
nand U6989 (N_6989,N_5819,N_5679);
nor U6990 (N_6990,N_4661,N_5692);
xnor U6991 (N_6991,N_5197,N_4247);
or U6992 (N_6992,N_4916,N_5445);
nor U6993 (N_6993,N_4305,N_4252);
nor U6994 (N_6994,N_5192,N_4625);
xor U6995 (N_6995,N_5138,N_4742);
xor U6996 (N_6996,N_5267,N_5954);
or U6997 (N_6997,N_5357,N_4440);
nor U6998 (N_6998,N_5390,N_5956);
and U6999 (N_6999,N_5338,N_4480);
and U7000 (N_7000,N_5599,N_5319);
nor U7001 (N_7001,N_5409,N_5102);
nor U7002 (N_7002,N_4112,N_5194);
and U7003 (N_7003,N_5793,N_5813);
nand U7004 (N_7004,N_5054,N_4736);
nor U7005 (N_7005,N_4192,N_4331);
nand U7006 (N_7006,N_5940,N_4290);
xor U7007 (N_7007,N_4837,N_5521);
nand U7008 (N_7008,N_4654,N_5674);
and U7009 (N_7009,N_4384,N_4522);
nand U7010 (N_7010,N_5645,N_4870);
nor U7011 (N_7011,N_4138,N_5756);
nor U7012 (N_7012,N_4604,N_5226);
nand U7013 (N_7013,N_5310,N_4864);
or U7014 (N_7014,N_5410,N_5022);
nor U7015 (N_7015,N_4519,N_4954);
or U7016 (N_7016,N_5857,N_5064);
nand U7017 (N_7017,N_5944,N_5756);
nand U7018 (N_7018,N_5302,N_5915);
xor U7019 (N_7019,N_5197,N_5206);
and U7020 (N_7020,N_5095,N_5815);
xnor U7021 (N_7021,N_5006,N_4488);
xor U7022 (N_7022,N_5115,N_5169);
or U7023 (N_7023,N_4499,N_5179);
nand U7024 (N_7024,N_4733,N_4476);
or U7025 (N_7025,N_5092,N_4545);
and U7026 (N_7026,N_4276,N_4028);
or U7027 (N_7027,N_5452,N_4912);
and U7028 (N_7028,N_5114,N_4236);
nor U7029 (N_7029,N_4012,N_5703);
and U7030 (N_7030,N_4265,N_5668);
nor U7031 (N_7031,N_5229,N_5534);
or U7032 (N_7032,N_4283,N_5086);
nor U7033 (N_7033,N_5627,N_4584);
nor U7034 (N_7034,N_5289,N_4906);
nand U7035 (N_7035,N_4185,N_4112);
and U7036 (N_7036,N_4144,N_5808);
nor U7037 (N_7037,N_4784,N_4086);
and U7038 (N_7038,N_4355,N_5479);
nor U7039 (N_7039,N_5581,N_4354);
nor U7040 (N_7040,N_4715,N_4154);
xor U7041 (N_7041,N_4634,N_4601);
or U7042 (N_7042,N_5696,N_4634);
xor U7043 (N_7043,N_5396,N_4043);
nand U7044 (N_7044,N_4147,N_5163);
or U7045 (N_7045,N_4893,N_5595);
nor U7046 (N_7046,N_5723,N_4952);
nor U7047 (N_7047,N_5476,N_4213);
or U7048 (N_7048,N_4221,N_4015);
or U7049 (N_7049,N_5273,N_4780);
nand U7050 (N_7050,N_5775,N_4030);
and U7051 (N_7051,N_4139,N_5731);
or U7052 (N_7052,N_4889,N_4755);
nand U7053 (N_7053,N_5909,N_4453);
nor U7054 (N_7054,N_5896,N_5883);
nor U7055 (N_7055,N_4378,N_5781);
nand U7056 (N_7056,N_4804,N_4617);
or U7057 (N_7057,N_4658,N_5665);
nand U7058 (N_7058,N_4925,N_5526);
nand U7059 (N_7059,N_4005,N_5560);
nand U7060 (N_7060,N_4205,N_4739);
xor U7061 (N_7061,N_4791,N_4743);
and U7062 (N_7062,N_5796,N_5795);
nor U7063 (N_7063,N_4966,N_5571);
and U7064 (N_7064,N_5780,N_5395);
nor U7065 (N_7065,N_4559,N_5661);
nand U7066 (N_7066,N_4137,N_5747);
nand U7067 (N_7067,N_4417,N_5383);
and U7068 (N_7068,N_4536,N_4640);
nor U7069 (N_7069,N_5822,N_5362);
xnor U7070 (N_7070,N_4674,N_5480);
and U7071 (N_7071,N_4230,N_5741);
nand U7072 (N_7072,N_5566,N_5788);
nor U7073 (N_7073,N_5644,N_5114);
or U7074 (N_7074,N_5008,N_5077);
and U7075 (N_7075,N_4345,N_4361);
nor U7076 (N_7076,N_5607,N_5392);
nand U7077 (N_7077,N_5183,N_5501);
nor U7078 (N_7078,N_5188,N_5330);
or U7079 (N_7079,N_5908,N_4395);
xor U7080 (N_7080,N_5442,N_4975);
xnor U7081 (N_7081,N_4246,N_4850);
nand U7082 (N_7082,N_4207,N_4891);
xor U7083 (N_7083,N_5982,N_4252);
or U7084 (N_7084,N_5782,N_4389);
and U7085 (N_7085,N_4028,N_4134);
nand U7086 (N_7086,N_4457,N_4602);
nor U7087 (N_7087,N_5199,N_4733);
nor U7088 (N_7088,N_5810,N_5411);
xor U7089 (N_7089,N_4603,N_4546);
nand U7090 (N_7090,N_4605,N_5867);
nor U7091 (N_7091,N_5987,N_4640);
or U7092 (N_7092,N_5311,N_4350);
xor U7093 (N_7093,N_4456,N_4460);
xor U7094 (N_7094,N_5697,N_4525);
xor U7095 (N_7095,N_4895,N_5400);
nor U7096 (N_7096,N_5447,N_4510);
nand U7097 (N_7097,N_4753,N_5436);
xnor U7098 (N_7098,N_4753,N_5308);
and U7099 (N_7099,N_4650,N_4801);
nand U7100 (N_7100,N_5978,N_4762);
and U7101 (N_7101,N_5176,N_5369);
and U7102 (N_7102,N_4977,N_4437);
or U7103 (N_7103,N_5011,N_5520);
nor U7104 (N_7104,N_4412,N_4277);
nor U7105 (N_7105,N_4666,N_5155);
nand U7106 (N_7106,N_5446,N_4956);
nor U7107 (N_7107,N_5117,N_5395);
xor U7108 (N_7108,N_5828,N_4384);
xor U7109 (N_7109,N_5455,N_5293);
nand U7110 (N_7110,N_5723,N_5671);
xnor U7111 (N_7111,N_4746,N_4823);
or U7112 (N_7112,N_4818,N_5451);
and U7113 (N_7113,N_4810,N_4546);
nor U7114 (N_7114,N_4623,N_4057);
xnor U7115 (N_7115,N_5350,N_5976);
nor U7116 (N_7116,N_4420,N_4080);
or U7117 (N_7117,N_4140,N_4956);
xnor U7118 (N_7118,N_5995,N_4174);
or U7119 (N_7119,N_4401,N_4081);
or U7120 (N_7120,N_4632,N_4424);
or U7121 (N_7121,N_5077,N_5894);
nand U7122 (N_7122,N_5747,N_4491);
nor U7123 (N_7123,N_5115,N_5861);
nand U7124 (N_7124,N_4326,N_5638);
and U7125 (N_7125,N_5423,N_5594);
xor U7126 (N_7126,N_4622,N_5255);
nand U7127 (N_7127,N_4110,N_4961);
and U7128 (N_7128,N_5021,N_5328);
and U7129 (N_7129,N_5216,N_5759);
nor U7130 (N_7130,N_4087,N_4414);
nand U7131 (N_7131,N_5068,N_5358);
and U7132 (N_7132,N_4321,N_5442);
or U7133 (N_7133,N_5947,N_4625);
nand U7134 (N_7134,N_5086,N_5858);
xnor U7135 (N_7135,N_5811,N_5325);
or U7136 (N_7136,N_4775,N_5294);
nand U7137 (N_7137,N_5264,N_5007);
nor U7138 (N_7138,N_5778,N_5391);
and U7139 (N_7139,N_4835,N_4732);
nor U7140 (N_7140,N_5785,N_4888);
nor U7141 (N_7141,N_4336,N_4463);
xor U7142 (N_7142,N_5263,N_5239);
nor U7143 (N_7143,N_4075,N_5195);
nor U7144 (N_7144,N_4039,N_5716);
nand U7145 (N_7145,N_5254,N_4047);
nor U7146 (N_7146,N_5538,N_4769);
or U7147 (N_7147,N_4356,N_4974);
xnor U7148 (N_7148,N_4754,N_4066);
nor U7149 (N_7149,N_4898,N_5578);
or U7150 (N_7150,N_5218,N_4680);
xor U7151 (N_7151,N_4889,N_5180);
nor U7152 (N_7152,N_4320,N_4811);
or U7153 (N_7153,N_5180,N_5336);
and U7154 (N_7154,N_5168,N_4988);
or U7155 (N_7155,N_4970,N_5321);
or U7156 (N_7156,N_4582,N_4133);
nand U7157 (N_7157,N_5486,N_5814);
xnor U7158 (N_7158,N_4207,N_5761);
or U7159 (N_7159,N_4215,N_5196);
or U7160 (N_7160,N_5953,N_5571);
and U7161 (N_7161,N_4437,N_5260);
nor U7162 (N_7162,N_5627,N_4604);
nor U7163 (N_7163,N_4895,N_4153);
nor U7164 (N_7164,N_5252,N_5816);
xor U7165 (N_7165,N_4715,N_5215);
xnor U7166 (N_7166,N_5882,N_4974);
and U7167 (N_7167,N_4998,N_4801);
nand U7168 (N_7168,N_5504,N_4273);
nor U7169 (N_7169,N_4899,N_5414);
or U7170 (N_7170,N_5076,N_5324);
xnor U7171 (N_7171,N_4444,N_5374);
and U7172 (N_7172,N_5751,N_5732);
and U7173 (N_7173,N_4160,N_4614);
and U7174 (N_7174,N_4659,N_5132);
or U7175 (N_7175,N_4674,N_5225);
or U7176 (N_7176,N_5610,N_5515);
nand U7177 (N_7177,N_4933,N_5786);
nor U7178 (N_7178,N_4063,N_4604);
nand U7179 (N_7179,N_4429,N_4969);
or U7180 (N_7180,N_5762,N_4554);
and U7181 (N_7181,N_5294,N_4898);
nor U7182 (N_7182,N_4183,N_5130);
nor U7183 (N_7183,N_5697,N_5533);
or U7184 (N_7184,N_4395,N_5086);
xnor U7185 (N_7185,N_4937,N_5115);
nor U7186 (N_7186,N_4751,N_4458);
nor U7187 (N_7187,N_5909,N_5399);
nand U7188 (N_7188,N_5077,N_5080);
and U7189 (N_7189,N_5555,N_5872);
nand U7190 (N_7190,N_5956,N_4359);
nor U7191 (N_7191,N_5081,N_5181);
or U7192 (N_7192,N_5020,N_5443);
nor U7193 (N_7193,N_5524,N_5263);
or U7194 (N_7194,N_4217,N_5445);
nor U7195 (N_7195,N_5533,N_4345);
nand U7196 (N_7196,N_5263,N_5750);
or U7197 (N_7197,N_5952,N_5132);
nor U7198 (N_7198,N_5021,N_5396);
and U7199 (N_7199,N_5429,N_4098);
xnor U7200 (N_7200,N_5268,N_5641);
or U7201 (N_7201,N_4531,N_5904);
xor U7202 (N_7202,N_5853,N_5512);
and U7203 (N_7203,N_4322,N_5722);
nand U7204 (N_7204,N_4526,N_5582);
nand U7205 (N_7205,N_5273,N_5375);
nand U7206 (N_7206,N_5010,N_5710);
or U7207 (N_7207,N_4283,N_5170);
or U7208 (N_7208,N_4631,N_5190);
or U7209 (N_7209,N_4349,N_5119);
xnor U7210 (N_7210,N_5937,N_4711);
and U7211 (N_7211,N_4611,N_4232);
nand U7212 (N_7212,N_4665,N_5044);
or U7213 (N_7213,N_4479,N_4812);
xor U7214 (N_7214,N_5902,N_5927);
nand U7215 (N_7215,N_4224,N_5812);
xnor U7216 (N_7216,N_5326,N_5375);
nand U7217 (N_7217,N_5435,N_4784);
nor U7218 (N_7218,N_5650,N_5164);
or U7219 (N_7219,N_5030,N_4377);
and U7220 (N_7220,N_4602,N_5523);
nor U7221 (N_7221,N_5418,N_5587);
or U7222 (N_7222,N_4969,N_5586);
and U7223 (N_7223,N_4730,N_4429);
nor U7224 (N_7224,N_4905,N_5966);
and U7225 (N_7225,N_4851,N_5695);
xnor U7226 (N_7226,N_5753,N_4124);
nor U7227 (N_7227,N_4584,N_5134);
xor U7228 (N_7228,N_4817,N_5883);
and U7229 (N_7229,N_4260,N_4530);
xor U7230 (N_7230,N_5341,N_4568);
nand U7231 (N_7231,N_5232,N_5100);
xor U7232 (N_7232,N_4141,N_4070);
xnor U7233 (N_7233,N_5253,N_4269);
nand U7234 (N_7234,N_4923,N_5428);
nand U7235 (N_7235,N_4034,N_4274);
nand U7236 (N_7236,N_5782,N_5152);
or U7237 (N_7237,N_4657,N_4309);
and U7238 (N_7238,N_4552,N_4127);
and U7239 (N_7239,N_5992,N_4171);
and U7240 (N_7240,N_5017,N_5080);
xnor U7241 (N_7241,N_4408,N_5273);
nor U7242 (N_7242,N_5467,N_4864);
nand U7243 (N_7243,N_4100,N_4057);
or U7244 (N_7244,N_4496,N_5824);
xnor U7245 (N_7245,N_5076,N_5465);
nor U7246 (N_7246,N_4554,N_4672);
or U7247 (N_7247,N_5763,N_4199);
nor U7248 (N_7248,N_5484,N_4762);
nand U7249 (N_7249,N_4111,N_5964);
and U7250 (N_7250,N_4655,N_5369);
and U7251 (N_7251,N_5108,N_5202);
xor U7252 (N_7252,N_5917,N_5004);
nor U7253 (N_7253,N_5236,N_4485);
nand U7254 (N_7254,N_4369,N_4645);
and U7255 (N_7255,N_5857,N_4073);
nand U7256 (N_7256,N_5797,N_5118);
nand U7257 (N_7257,N_5333,N_5389);
nand U7258 (N_7258,N_4741,N_5334);
or U7259 (N_7259,N_4068,N_5053);
or U7260 (N_7260,N_4125,N_5014);
xnor U7261 (N_7261,N_5613,N_4713);
nor U7262 (N_7262,N_5520,N_4372);
nand U7263 (N_7263,N_5609,N_4140);
and U7264 (N_7264,N_4489,N_4275);
xnor U7265 (N_7265,N_4696,N_5136);
nand U7266 (N_7266,N_5981,N_5749);
or U7267 (N_7267,N_4776,N_5203);
nand U7268 (N_7268,N_5565,N_5484);
nand U7269 (N_7269,N_5374,N_4012);
nand U7270 (N_7270,N_4538,N_5817);
nand U7271 (N_7271,N_4912,N_5943);
nand U7272 (N_7272,N_5671,N_4023);
xnor U7273 (N_7273,N_4521,N_5541);
or U7274 (N_7274,N_4109,N_5665);
or U7275 (N_7275,N_5589,N_5155);
xnor U7276 (N_7276,N_4896,N_5689);
or U7277 (N_7277,N_5436,N_5989);
nand U7278 (N_7278,N_5236,N_4935);
nor U7279 (N_7279,N_4139,N_5363);
nor U7280 (N_7280,N_4428,N_5213);
nor U7281 (N_7281,N_5254,N_4936);
or U7282 (N_7282,N_4388,N_4878);
nor U7283 (N_7283,N_5339,N_4170);
nor U7284 (N_7284,N_4525,N_4908);
xnor U7285 (N_7285,N_4914,N_5963);
or U7286 (N_7286,N_4724,N_5211);
xnor U7287 (N_7287,N_4830,N_5351);
xor U7288 (N_7288,N_4230,N_5533);
xor U7289 (N_7289,N_5370,N_4397);
and U7290 (N_7290,N_5748,N_4230);
nor U7291 (N_7291,N_5387,N_4190);
xor U7292 (N_7292,N_4663,N_5772);
nand U7293 (N_7293,N_4698,N_4193);
xnor U7294 (N_7294,N_5745,N_4788);
xor U7295 (N_7295,N_5657,N_4625);
nand U7296 (N_7296,N_5837,N_4758);
xnor U7297 (N_7297,N_4427,N_5072);
and U7298 (N_7298,N_4997,N_4500);
xor U7299 (N_7299,N_5694,N_5793);
nor U7300 (N_7300,N_5389,N_5563);
and U7301 (N_7301,N_4721,N_4853);
xor U7302 (N_7302,N_5330,N_5174);
and U7303 (N_7303,N_5849,N_5299);
and U7304 (N_7304,N_4593,N_4662);
xor U7305 (N_7305,N_4758,N_4973);
xor U7306 (N_7306,N_5304,N_4215);
and U7307 (N_7307,N_4021,N_4894);
nor U7308 (N_7308,N_4900,N_4005);
nand U7309 (N_7309,N_5148,N_5606);
xor U7310 (N_7310,N_4569,N_5099);
nand U7311 (N_7311,N_4180,N_5012);
and U7312 (N_7312,N_5330,N_4945);
or U7313 (N_7313,N_5206,N_4169);
and U7314 (N_7314,N_5034,N_5957);
nor U7315 (N_7315,N_4044,N_4934);
nor U7316 (N_7316,N_5447,N_5554);
xnor U7317 (N_7317,N_4601,N_4002);
xor U7318 (N_7318,N_5960,N_4707);
and U7319 (N_7319,N_5404,N_4392);
nand U7320 (N_7320,N_4063,N_4854);
nor U7321 (N_7321,N_4472,N_5493);
nor U7322 (N_7322,N_4088,N_4765);
and U7323 (N_7323,N_4935,N_4947);
xor U7324 (N_7324,N_5500,N_4238);
nand U7325 (N_7325,N_5457,N_5653);
and U7326 (N_7326,N_4514,N_4444);
and U7327 (N_7327,N_4181,N_4619);
or U7328 (N_7328,N_5006,N_4050);
or U7329 (N_7329,N_4446,N_4358);
and U7330 (N_7330,N_5501,N_5727);
nand U7331 (N_7331,N_4714,N_4128);
or U7332 (N_7332,N_4690,N_5466);
and U7333 (N_7333,N_5517,N_4675);
or U7334 (N_7334,N_4482,N_4899);
or U7335 (N_7335,N_4996,N_5377);
and U7336 (N_7336,N_5792,N_5278);
xnor U7337 (N_7337,N_5649,N_5865);
or U7338 (N_7338,N_4573,N_4719);
nor U7339 (N_7339,N_5110,N_4683);
nor U7340 (N_7340,N_5419,N_5278);
nand U7341 (N_7341,N_5830,N_4720);
or U7342 (N_7342,N_5467,N_5860);
nor U7343 (N_7343,N_5334,N_5003);
nand U7344 (N_7344,N_4835,N_5259);
nand U7345 (N_7345,N_4683,N_4304);
or U7346 (N_7346,N_5032,N_5463);
nor U7347 (N_7347,N_5735,N_5196);
nand U7348 (N_7348,N_4676,N_4080);
nand U7349 (N_7349,N_5512,N_5201);
nand U7350 (N_7350,N_5274,N_5365);
or U7351 (N_7351,N_4227,N_4028);
or U7352 (N_7352,N_4305,N_4733);
or U7353 (N_7353,N_4800,N_5366);
or U7354 (N_7354,N_5016,N_4351);
xor U7355 (N_7355,N_5269,N_5544);
nor U7356 (N_7356,N_4686,N_4702);
xnor U7357 (N_7357,N_4777,N_4608);
nand U7358 (N_7358,N_5313,N_4243);
nand U7359 (N_7359,N_5474,N_5129);
xnor U7360 (N_7360,N_4555,N_5514);
and U7361 (N_7361,N_5328,N_4068);
nand U7362 (N_7362,N_4958,N_4513);
or U7363 (N_7363,N_5720,N_4073);
nor U7364 (N_7364,N_4968,N_4118);
and U7365 (N_7365,N_5924,N_4566);
xor U7366 (N_7366,N_5887,N_4884);
xnor U7367 (N_7367,N_4548,N_4210);
xor U7368 (N_7368,N_4422,N_5260);
nor U7369 (N_7369,N_4112,N_5469);
nand U7370 (N_7370,N_4053,N_4941);
nand U7371 (N_7371,N_4615,N_5248);
nor U7372 (N_7372,N_5181,N_4728);
or U7373 (N_7373,N_4273,N_4503);
nand U7374 (N_7374,N_4459,N_5898);
and U7375 (N_7375,N_4960,N_4163);
nand U7376 (N_7376,N_4412,N_5383);
or U7377 (N_7377,N_4940,N_4672);
nor U7378 (N_7378,N_5965,N_5876);
xor U7379 (N_7379,N_4275,N_5729);
xnor U7380 (N_7380,N_5116,N_5378);
and U7381 (N_7381,N_4485,N_4451);
xnor U7382 (N_7382,N_4235,N_5725);
nor U7383 (N_7383,N_5191,N_5954);
or U7384 (N_7384,N_5828,N_4659);
or U7385 (N_7385,N_4591,N_5590);
nor U7386 (N_7386,N_4497,N_5147);
nand U7387 (N_7387,N_5075,N_4123);
nand U7388 (N_7388,N_4566,N_5353);
and U7389 (N_7389,N_5115,N_4508);
and U7390 (N_7390,N_4830,N_5497);
nor U7391 (N_7391,N_4484,N_4755);
xnor U7392 (N_7392,N_5990,N_4688);
nand U7393 (N_7393,N_5621,N_5461);
xor U7394 (N_7394,N_5849,N_4433);
nand U7395 (N_7395,N_5063,N_5467);
xor U7396 (N_7396,N_4856,N_4497);
or U7397 (N_7397,N_5984,N_5425);
or U7398 (N_7398,N_5864,N_5019);
nor U7399 (N_7399,N_4790,N_4113);
nor U7400 (N_7400,N_4775,N_4516);
nor U7401 (N_7401,N_4452,N_4849);
nor U7402 (N_7402,N_5810,N_5515);
nand U7403 (N_7403,N_5906,N_4120);
and U7404 (N_7404,N_4750,N_5138);
nor U7405 (N_7405,N_5159,N_5165);
nor U7406 (N_7406,N_4107,N_5222);
nand U7407 (N_7407,N_5038,N_4359);
nor U7408 (N_7408,N_4436,N_5353);
or U7409 (N_7409,N_5942,N_4541);
or U7410 (N_7410,N_4615,N_4244);
nand U7411 (N_7411,N_4231,N_4735);
and U7412 (N_7412,N_5047,N_5317);
nor U7413 (N_7413,N_5904,N_4842);
or U7414 (N_7414,N_4158,N_4094);
xor U7415 (N_7415,N_4424,N_4948);
xnor U7416 (N_7416,N_4253,N_5079);
or U7417 (N_7417,N_5461,N_4161);
or U7418 (N_7418,N_5116,N_4278);
xnor U7419 (N_7419,N_4336,N_4762);
or U7420 (N_7420,N_4138,N_4645);
or U7421 (N_7421,N_4930,N_4948);
or U7422 (N_7422,N_4037,N_5360);
nor U7423 (N_7423,N_5543,N_4148);
or U7424 (N_7424,N_5244,N_5995);
and U7425 (N_7425,N_4736,N_5774);
nor U7426 (N_7426,N_5653,N_5765);
or U7427 (N_7427,N_5574,N_5160);
nor U7428 (N_7428,N_4444,N_5861);
and U7429 (N_7429,N_5598,N_5102);
nand U7430 (N_7430,N_5727,N_5611);
nand U7431 (N_7431,N_5357,N_5255);
xor U7432 (N_7432,N_5219,N_4584);
nor U7433 (N_7433,N_4393,N_5126);
or U7434 (N_7434,N_5880,N_5262);
and U7435 (N_7435,N_5216,N_5230);
nand U7436 (N_7436,N_5552,N_5728);
and U7437 (N_7437,N_4036,N_5744);
and U7438 (N_7438,N_4176,N_4522);
nand U7439 (N_7439,N_4599,N_5502);
xor U7440 (N_7440,N_5685,N_5151);
and U7441 (N_7441,N_5811,N_5293);
xor U7442 (N_7442,N_5682,N_5906);
xnor U7443 (N_7443,N_4684,N_5270);
nor U7444 (N_7444,N_4689,N_4023);
nand U7445 (N_7445,N_4772,N_5704);
nand U7446 (N_7446,N_4433,N_4715);
nor U7447 (N_7447,N_5329,N_5814);
and U7448 (N_7448,N_4730,N_4212);
nor U7449 (N_7449,N_4366,N_5693);
xnor U7450 (N_7450,N_4270,N_5261);
and U7451 (N_7451,N_5564,N_5145);
nor U7452 (N_7452,N_5539,N_4112);
or U7453 (N_7453,N_4285,N_4917);
or U7454 (N_7454,N_4253,N_4830);
or U7455 (N_7455,N_4949,N_5755);
nor U7456 (N_7456,N_4664,N_4278);
nor U7457 (N_7457,N_5103,N_5467);
or U7458 (N_7458,N_5979,N_4202);
nor U7459 (N_7459,N_5136,N_4914);
and U7460 (N_7460,N_4062,N_5825);
xnor U7461 (N_7461,N_5224,N_4330);
nand U7462 (N_7462,N_4928,N_5942);
and U7463 (N_7463,N_4116,N_5502);
nand U7464 (N_7464,N_5706,N_4342);
nand U7465 (N_7465,N_5841,N_5709);
nand U7466 (N_7466,N_5119,N_4276);
nor U7467 (N_7467,N_5334,N_4568);
or U7468 (N_7468,N_4439,N_4586);
and U7469 (N_7469,N_5398,N_4354);
and U7470 (N_7470,N_5551,N_5045);
nand U7471 (N_7471,N_4002,N_4552);
xnor U7472 (N_7472,N_4218,N_5442);
nand U7473 (N_7473,N_5927,N_4479);
nor U7474 (N_7474,N_4078,N_4526);
xnor U7475 (N_7475,N_5665,N_4941);
nor U7476 (N_7476,N_4049,N_4215);
nand U7477 (N_7477,N_5434,N_5429);
nor U7478 (N_7478,N_5465,N_5207);
xor U7479 (N_7479,N_4868,N_5132);
nand U7480 (N_7480,N_4724,N_5294);
xor U7481 (N_7481,N_5850,N_4870);
nor U7482 (N_7482,N_4713,N_5366);
xnor U7483 (N_7483,N_4463,N_5904);
or U7484 (N_7484,N_5737,N_5403);
nand U7485 (N_7485,N_4671,N_4258);
nor U7486 (N_7486,N_5491,N_4834);
xnor U7487 (N_7487,N_5960,N_5207);
nand U7488 (N_7488,N_5767,N_5682);
nand U7489 (N_7489,N_4091,N_5554);
and U7490 (N_7490,N_4688,N_4289);
nor U7491 (N_7491,N_5421,N_5012);
and U7492 (N_7492,N_5422,N_4498);
and U7493 (N_7493,N_5351,N_5538);
or U7494 (N_7494,N_4117,N_4434);
and U7495 (N_7495,N_5467,N_5941);
nand U7496 (N_7496,N_4513,N_4743);
or U7497 (N_7497,N_4581,N_5594);
nand U7498 (N_7498,N_5378,N_4962);
nor U7499 (N_7499,N_5299,N_5165);
and U7500 (N_7500,N_5253,N_5549);
nor U7501 (N_7501,N_5997,N_4257);
and U7502 (N_7502,N_4964,N_5755);
nand U7503 (N_7503,N_5275,N_5876);
xnor U7504 (N_7504,N_4268,N_5557);
and U7505 (N_7505,N_5053,N_4482);
xor U7506 (N_7506,N_4440,N_5822);
nor U7507 (N_7507,N_5987,N_4753);
nand U7508 (N_7508,N_4572,N_4423);
xor U7509 (N_7509,N_4617,N_5101);
nor U7510 (N_7510,N_4609,N_5522);
or U7511 (N_7511,N_5454,N_4829);
nand U7512 (N_7512,N_4370,N_5334);
or U7513 (N_7513,N_4766,N_5027);
nor U7514 (N_7514,N_5773,N_5359);
and U7515 (N_7515,N_5997,N_4953);
and U7516 (N_7516,N_5194,N_4298);
and U7517 (N_7517,N_5210,N_5038);
nor U7518 (N_7518,N_4515,N_5065);
nand U7519 (N_7519,N_5469,N_4096);
or U7520 (N_7520,N_5094,N_4495);
and U7521 (N_7521,N_4214,N_4207);
nand U7522 (N_7522,N_4064,N_4538);
nand U7523 (N_7523,N_5491,N_4769);
xnor U7524 (N_7524,N_4851,N_5939);
or U7525 (N_7525,N_5248,N_5302);
xor U7526 (N_7526,N_5952,N_5139);
and U7527 (N_7527,N_5177,N_4897);
nor U7528 (N_7528,N_4704,N_4590);
xor U7529 (N_7529,N_4808,N_4026);
xor U7530 (N_7530,N_4337,N_5772);
and U7531 (N_7531,N_5404,N_4737);
nand U7532 (N_7532,N_4792,N_4898);
nor U7533 (N_7533,N_4299,N_5545);
and U7534 (N_7534,N_4612,N_4338);
nand U7535 (N_7535,N_4869,N_4378);
nand U7536 (N_7536,N_5067,N_4614);
xnor U7537 (N_7537,N_4267,N_4209);
or U7538 (N_7538,N_5651,N_5145);
nor U7539 (N_7539,N_4645,N_5020);
and U7540 (N_7540,N_5306,N_5799);
xor U7541 (N_7541,N_5683,N_5312);
xor U7542 (N_7542,N_5577,N_5549);
or U7543 (N_7543,N_4123,N_5893);
nor U7544 (N_7544,N_5194,N_5482);
nand U7545 (N_7545,N_4363,N_4148);
and U7546 (N_7546,N_4659,N_4718);
and U7547 (N_7547,N_4840,N_4779);
xnor U7548 (N_7548,N_5876,N_4396);
nor U7549 (N_7549,N_4147,N_5038);
nor U7550 (N_7550,N_5034,N_4018);
and U7551 (N_7551,N_4207,N_4535);
or U7552 (N_7552,N_4630,N_5550);
xnor U7553 (N_7553,N_5026,N_5151);
nand U7554 (N_7554,N_4236,N_4470);
nor U7555 (N_7555,N_5324,N_4804);
xnor U7556 (N_7556,N_5916,N_5514);
nand U7557 (N_7557,N_4103,N_5808);
nor U7558 (N_7558,N_4773,N_5016);
and U7559 (N_7559,N_5270,N_5556);
nor U7560 (N_7560,N_5610,N_4282);
nand U7561 (N_7561,N_5980,N_4715);
and U7562 (N_7562,N_5602,N_4941);
and U7563 (N_7563,N_5912,N_4776);
xnor U7564 (N_7564,N_5282,N_5079);
or U7565 (N_7565,N_5674,N_5523);
nand U7566 (N_7566,N_4537,N_4493);
or U7567 (N_7567,N_4469,N_5568);
or U7568 (N_7568,N_4875,N_5555);
xor U7569 (N_7569,N_5483,N_4755);
or U7570 (N_7570,N_4852,N_5746);
xnor U7571 (N_7571,N_5189,N_5738);
nand U7572 (N_7572,N_4587,N_5955);
and U7573 (N_7573,N_5965,N_4416);
nor U7574 (N_7574,N_5539,N_4000);
or U7575 (N_7575,N_5852,N_4879);
or U7576 (N_7576,N_5836,N_4346);
nand U7577 (N_7577,N_4246,N_4992);
and U7578 (N_7578,N_5443,N_5924);
xor U7579 (N_7579,N_4570,N_5417);
or U7580 (N_7580,N_4071,N_5492);
nand U7581 (N_7581,N_5013,N_5119);
xor U7582 (N_7582,N_5129,N_5330);
xor U7583 (N_7583,N_5869,N_4621);
xor U7584 (N_7584,N_4464,N_4835);
nor U7585 (N_7585,N_5593,N_5839);
nand U7586 (N_7586,N_4391,N_5171);
and U7587 (N_7587,N_4734,N_4580);
nor U7588 (N_7588,N_5834,N_5662);
nand U7589 (N_7589,N_4306,N_4659);
and U7590 (N_7590,N_5853,N_4969);
xnor U7591 (N_7591,N_5082,N_4500);
xor U7592 (N_7592,N_5391,N_5927);
or U7593 (N_7593,N_5116,N_5985);
nand U7594 (N_7594,N_4421,N_4626);
xnor U7595 (N_7595,N_4741,N_5850);
nand U7596 (N_7596,N_4909,N_5210);
and U7597 (N_7597,N_5814,N_5312);
nand U7598 (N_7598,N_5280,N_5420);
nand U7599 (N_7599,N_5548,N_4875);
and U7600 (N_7600,N_4908,N_4655);
nor U7601 (N_7601,N_4862,N_5147);
nand U7602 (N_7602,N_4583,N_4551);
and U7603 (N_7603,N_4832,N_4531);
or U7604 (N_7604,N_4794,N_4942);
and U7605 (N_7605,N_5849,N_5640);
nor U7606 (N_7606,N_5635,N_5632);
xor U7607 (N_7607,N_5590,N_5267);
or U7608 (N_7608,N_5004,N_4914);
and U7609 (N_7609,N_4879,N_4617);
nor U7610 (N_7610,N_4926,N_4750);
xnor U7611 (N_7611,N_5095,N_5728);
nor U7612 (N_7612,N_4457,N_5353);
xnor U7613 (N_7613,N_5151,N_4072);
nor U7614 (N_7614,N_4418,N_4310);
and U7615 (N_7615,N_4735,N_5059);
or U7616 (N_7616,N_5812,N_5730);
xnor U7617 (N_7617,N_4794,N_4410);
xor U7618 (N_7618,N_5713,N_5125);
nor U7619 (N_7619,N_4882,N_5214);
nand U7620 (N_7620,N_4218,N_4319);
or U7621 (N_7621,N_5572,N_4984);
nand U7622 (N_7622,N_5555,N_5601);
or U7623 (N_7623,N_5557,N_5644);
and U7624 (N_7624,N_4849,N_4238);
nand U7625 (N_7625,N_5037,N_5036);
xor U7626 (N_7626,N_4634,N_5612);
xor U7627 (N_7627,N_5194,N_5881);
nand U7628 (N_7628,N_4645,N_4852);
nand U7629 (N_7629,N_4503,N_4284);
and U7630 (N_7630,N_5217,N_4471);
and U7631 (N_7631,N_5397,N_5713);
or U7632 (N_7632,N_4471,N_4824);
or U7633 (N_7633,N_4443,N_4178);
nor U7634 (N_7634,N_5311,N_5218);
nor U7635 (N_7635,N_5908,N_4255);
or U7636 (N_7636,N_5709,N_5723);
and U7637 (N_7637,N_4931,N_5291);
nand U7638 (N_7638,N_5114,N_4325);
xor U7639 (N_7639,N_5746,N_5511);
xor U7640 (N_7640,N_4108,N_4685);
and U7641 (N_7641,N_5791,N_5162);
or U7642 (N_7642,N_4889,N_5699);
nand U7643 (N_7643,N_4869,N_5853);
nand U7644 (N_7644,N_4799,N_4516);
xnor U7645 (N_7645,N_4885,N_4211);
nor U7646 (N_7646,N_5106,N_4724);
and U7647 (N_7647,N_5989,N_5910);
xor U7648 (N_7648,N_4371,N_4534);
xor U7649 (N_7649,N_5609,N_5719);
and U7650 (N_7650,N_5344,N_4390);
and U7651 (N_7651,N_5989,N_4599);
and U7652 (N_7652,N_5856,N_4391);
and U7653 (N_7653,N_4923,N_5240);
xnor U7654 (N_7654,N_4487,N_5026);
and U7655 (N_7655,N_4582,N_5811);
xor U7656 (N_7656,N_4660,N_5317);
nand U7657 (N_7657,N_5488,N_4233);
xnor U7658 (N_7658,N_5540,N_4977);
xor U7659 (N_7659,N_4349,N_4680);
nor U7660 (N_7660,N_4433,N_4792);
nand U7661 (N_7661,N_5462,N_5420);
nor U7662 (N_7662,N_5143,N_5333);
nand U7663 (N_7663,N_5844,N_4286);
nor U7664 (N_7664,N_4135,N_4755);
nand U7665 (N_7665,N_5220,N_4948);
or U7666 (N_7666,N_4469,N_4183);
or U7667 (N_7667,N_4886,N_4546);
and U7668 (N_7668,N_5179,N_5086);
nor U7669 (N_7669,N_4801,N_5599);
nor U7670 (N_7670,N_4531,N_4710);
xnor U7671 (N_7671,N_4003,N_4178);
xnor U7672 (N_7672,N_5824,N_4146);
or U7673 (N_7673,N_5281,N_4511);
nand U7674 (N_7674,N_4291,N_4535);
xnor U7675 (N_7675,N_4004,N_5294);
and U7676 (N_7676,N_5474,N_4789);
and U7677 (N_7677,N_4190,N_5170);
nor U7678 (N_7678,N_5108,N_5350);
or U7679 (N_7679,N_4137,N_4312);
xnor U7680 (N_7680,N_5875,N_4837);
nand U7681 (N_7681,N_5168,N_4298);
or U7682 (N_7682,N_4021,N_5490);
and U7683 (N_7683,N_5859,N_4675);
nand U7684 (N_7684,N_4565,N_4509);
xnor U7685 (N_7685,N_4826,N_5454);
nand U7686 (N_7686,N_5368,N_5441);
or U7687 (N_7687,N_4844,N_4491);
nor U7688 (N_7688,N_5925,N_4671);
or U7689 (N_7689,N_4460,N_4808);
nand U7690 (N_7690,N_4631,N_4532);
and U7691 (N_7691,N_5807,N_4468);
nand U7692 (N_7692,N_5612,N_4887);
nand U7693 (N_7693,N_4419,N_5405);
nor U7694 (N_7694,N_5989,N_5074);
and U7695 (N_7695,N_5096,N_5655);
or U7696 (N_7696,N_4379,N_4501);
or U7697 (N_7697,N_4381,N_5063);
nand U7698 (N_7698,N_5043,N_5629);
nor U7699 (N_7699,N_4983,N_5386);
nand U7700 (N_7700,N_5990,N_5745);
nand U7701 (N_7701,N_4337,N_5606);
and U7702 (N_7702,N_4612,N_5822);
nor U7703 (N_7703,N_4163,N_4131);
xnor U7704 (N_7704,N_4902,N_4122);
xor U7705 (N_7705,N_4503,N_5111);
or U7706 (N_7706,N_4937,N_5364);
and U7707 (N_7707,N_5052,N_5780);
or U7708 (N_7708,N_4909,N_5135);
xor U7709 (N_7709,N_4927,N_4445);
xor U7710 (N_7710,N_5599,N_4894);
xnor U7711 (N_7711,N_5818,N_5881);
nand U7712 (N_7712,N_5953,N_4292);
nor U7713 (N_7713,N_4128,N_4732);
nor U7714 (N_7714,N_5346,N_5352);
nand U7715 (N_7715,N_4618,N_5328);
nand U7716 (N_7716,N_5271,N_4926);
or U7717 (N_7717,N_5545,N_4344);
or U7718 (N_7718,N_4603,N_4854);
or U7719 (N_7719,N_4156,N_4666);
or U7720 (N_7720,N_4449,N_5452);
nor U7721 (N_7721,N_5761,N_5243);
nor U7722 (N_7722,N_4746,N_5939);
or U7723 (N_7723,N_4926,N_5414);
and U7724 (N_7724,N_5583,N_4502);
and U7725 (N_7725,N_4347,N_4903);
and U7726 (N_7726,N_5792,N_4133);
or U7727 (N_7727,N_4178,N_5165);
or U7728 (N_7728,N_4787,N_4325);
and U7729 (N_7729,N_5938,N_4212);
nor U7730 (N_7730,N_5632,N_5554);
or U7731 (N_7731,N_5615,N_4680);
and U7732 (N_7732,N_4214,N_5847);
xnor U7733 (N_7733,N_4387,N_4472);
nor U7734 (N_7734,N_5522,N_5154);
or U7735 (N_7735,N_5811,N_4988);
nand U7736 (N_7736,N_5246,N_4735);
nand U7737 (N_7737,N_5000,N_4729);
xnor U7738 (N_7738,N_5062,N_5760);
and U7739 (N_7739,N_4786,N_4463);
nand U7740 (N_7740,N_5235,N_4713);
or U7741 (N_7741,N_5838,N_4894);
nor U7742 (N_7742,N_5609,N_4715);
and U7743 (N_7743,N_5320,N_5269);
xor U7744 (N_7744,N_5210,N_5129);
nor U7745 (N_7745,N_4338,N_5403);
nand U7746 (N_7746,N_5960,N_4381);
or U7747 (N_7747,N_4825,N_4173);
xnor U7748 (N_7748,N_4553,N_4619);
xor U7749 (N_7749,N_4851,N_5639);
xor U7750 (N_7750,N_5463,N_4538);
or U7751 (N_7751,N_5339,N_5979);
nor U7752 (N_7752,N_5785,N_5781);
and U7753 (N_7753,N_5158,N_4773);
or U7754 (N_7754,N_5839,N_5889);
or U7755 (N_7755,N_5907,N_5821);
or U7756 (N_7756,N_4079,N_5869);
and U7757 (N_7757,N_5095,N_5654);
nand U7758 (N_7758,N_4492,N_5410);
nand U7759 (N_7759,N_5274,N_5465);
and U7760 (N_7760,N_5397,N_5672);
and U7761 (N_7761,N_4024,N_4880);
or U7762 (N_7762,N_5716,N_4346);
nor U7763 (N_7763,N_4770,N_4398);
and U7764 (N_7764,N_5667,N_5703);
nor U7765 (N_7765,N_4312,N_5382);
nand U7766 (N_7766,N_4672,N_4193);
and U7767 (N_7767,N_5768,N_4053);
and U7768 (N_7768,N_5510,N_5160);
xor U7769 (N_7769,N_4893,N_5108);
nand U7770 (N_7770,N_5328,N_5408);
or U7771 (N_7771,N_4470,N_4235);
or U7772 (N_7772,N_5950,N_4252);
nand U7773 (N_7773,N_4517,N_5173);
nand U7774 (N_7774,N_4826,N_4753);
or U7775 (N_7775,N_5783,N_4775);
and U7776 (N_7776,N_4611,N_5775);
xor U7777 (N_7777,N_5848,N_5739);
and U7778 (N_7778,N_5623,N_4623);
nand U7779 (N_7779,N_4108,N_5685);
nor U7780 (N_7780,N_4553,N_4596);
xor U7781 (N_7781,N_4734,N_4917);
nor U7782 (N_7782,N_4258,N_5173);
and U7783 (N_7783,N_4643,N_4765);
nand U7784 (N_7784,N_5244,N_4207);
or U7785 (N_7785,N_4475,N_4408);
and U7786 (N_7786,N_5011,N_4598);
and U7787 (N_7787,N_4927,N_5665);
nor U7788 (N_7788,N_5017,N_5028);
xor U7789 (N_7789,N_4337,N_5985);
nand U7790 (N_7790,N_4470,N_4902);
nand U7791 (N_7791,N_5266,N_4747);
and U7792 (N_7792,N_5868,N_4446);
nand U7793 (N_7793,N_5984,N_4449);
nand U7794 (N_7794,N_4517,N_4300);
nand U7795 (N_7795,N_5915,N_4684);
xor U7796 (N_7796,N_4354,N_5157);
or U7797 (N_7797,N_4994,N_4603);
and U7798 (N_7798,N_4926,N_5671);
nand U7799 (N_7799,N_4881,N_4957);
xor U7800 (N_7800,N_5243,N_4090);
and U7801 (N_7801,N_5118,N_4326);
nor U7802 (N_7802,N_5517,N_4183);
or U7803 (N_7803,N_5882,N_5194);
nor U7804 (N_7804,N_4966,N_5357);
and U7805 (N_7805,N_5141,N_5687);
nand U7806 (N_7806,N_5679,N_4410);
or U7807 (N_7807,N_4838,N_4722);
or U7808 (N_7808,N_4843,N_5696);
or U7809 (N_7809,N_4079,N_5634);
or U7810 (N_7810,N_4340,N_4652);
or U7811 (N_7811,N_5671,N_4084);
nand U7812 (N_7812,N_5804,N_4276);
nand U7813 (N_7813,N_5714,N_5326);
and U7814 (N_7814,N_4904,N_4010);
nand U7815 (N_7815,N_4298,N_5697);
xnor U7816 (N_7816,N_5243,N_5297);
nand U7817 (N_7817,N_5560,N_5288);
xor U7818 (N_7818,N_5477,N_4306);
nand U7819 (N_7819,N_4016,N_4663);
nor U7820 (N_7820,N_4672,N_4801);
nor U7821 (N_7821,N_5020,N_5641);
and U7822 (N_7822,N_4018,N_4398);
nor U7823 (N_7823,N_4931,N_4388);
and U7824 (N_7824,N_4538,N_5551);
xor U7825 (N_7825,N_5266,N_5140);
xor U7826 (N_7826,N_4852,N_5843);
nand U7827 (N_7827,N_4193,N_4471);
or U7828 (N_7828,N_5719,N_5893);
and U7829 (N_7829,N_4243,N_5793);
or U7830 (N_7830,N_4795,N_5878);
xor U7831 (N_7831,N_4783,N_5434);
nand U7832 (N_7832,N_4002,N_4079);
xnor U7833 (N_7833,N_5392,N_4989);
nand U7834 (N_7834,N_5824,N_4357);
or U7835 (N_7835,N_4406,N_4327);
and U7836 (N_7836,N_4142,N_5118);
xor U7837 (N_7837,N_4268,N_4395);
nand U7838 (N_7838,N_5232,N_5054);
or U7839 (N_7839,N_5483,N_4864);
nand U7840 (N_7840,N_5388,N_5289);
nand U7841 (N_7841,N_4102,N_5673);
xor U7842 (N_7842,N_5229,N_5292);
or U7843 (N_7843,N_5691,N_4710);
xor U7844 (N_7844,N_4492,N_5423);
nor U7845 (N_7845,N_4506,N_5362);
and U7846 (N_7846,N_4556,N_4995);
nor U7847 (N_7847,N_4667,N_4968);
nand U7848 (N_7848,N_5160,N_4459);
or U7849 (N_7849,N_5084,N_5381);
and U7850 (N_7850,N_4221,N_5095);
and U7851 (N_7851,N_4015,N_4231);
nor U7852 (N_7852,N_5903,N_4757);
or U7853 (N_7853,N_5431,N_5051);
xor U7854 (N_7854,N_5260,N_4943);
xnor U7855 (N_7855,N_4600,N_4020);
xnor U7856 (N_7856,N_4939,N_4879);
or U7857 (N_7857,N_5159,N_5607);
xor U7858 (N_7858,N_4246,N_4677);
xnor U7859 (N_7859,N_5160,N_5485);
or U7860 (N_7860,N_4923,N_5586);
and U7861 (N_7861,N_4413,N_4810);
and U7862 (N_7862,N_5192,N_4043);
nand U7863 (N_7863,N_5405,N_5103);
nor U7864 (N_7864,N_5509,N_4412);
nor U7865 (N_7865,N_5876,N_5078);
nor U7866 (N_7866,N_4426,N_4137);
nand U7867 (N_7867,N_5381,N_4383);
nor U7868 (N_7868,N_4352,N_5459);
or U7869 (N_7869,N_5588,N_5288);
xor U7870 (N_7870,N_5505,N_5173);
or U7871 (N_7871,N_5899,N_5753);
or U7872 (N_7872,N_5026,N_5381);
nand U7873 (N_7873,N_4898,N_5186);
xor U7874 (N_7874,N_5716,N_5077);
nand U7875 (N_7875,N_4876,N_4757);
and U7876 (N_7876,N_4459,N_5350);
or U7877 (N_7877,N_5201,N_4948);
nor U7878 (N_7878,N_4415,N_5222);
or U7879 (N_7879,N_5294,N_4941);
or U7880 (N_7880,N_4958,N_5022);
and U7881 (N_7881,N_5786,N_4371);
nor U7882 (N_7882,N_4459,N_4354);
or U7883 (N_7883,N_4572,N_5899);
nor U7884 (N_7884,N_4215,N_4952);
and U7885 (N_7885,N_5634,N_4052);
nand U7886 (N_7886,N_4802,N_5751);
or U7887 (N_7887,N_4794,N_5208);
or U7888 (N_7888,N_5030,N_5977);
nor U7889 (N_7889,N_5119,N_5012);
and U7890 (N_7890,N_5064,N_5581);
or U7891 (N_7891,N_5193,N_5280);
nand U7892 (N_7892,N_5295,N_5339);
and U7893 (N_7893,N_4174,N_5970);
nor U7894 (N_7894,N_4975,N_5402);
or U7895 (N_7895,N_4308,N_4989);
or U7896 (N_7896,N_5979,N_4575);
nor U7897 (N_7897,N_4250,N_5617);
and U7898 (N_7898,N_5913,N_5777);
or U7899 (N_7899,N_4330,N_5292);
xnor U7900 (N_7900,N_5120,N_5934);
and U7901 (N_7901,N_5390,N_5641);
or U7902 (N_7902,N_5419,N_4442);
or U7903 (N_7903,N_4728,N_4226);
xnor U7904 (N_7904,N_5620,N_4819);
or U7905 (N_7905,N_5609,N_4529);
xor U7906 (N_7906,N_4256,N_4644);
nand U7907 (N_7907,N_5129,N_5421);
xnor U7908 (N_7908,N_4163,N_5266);
or U7909 (N_7909,N_5384,N_4378);
nand U7910 (N_7910,N_5389,N_5543);
and U7911 (N_7911,N_4709,N_5303);
and U7912 (N_7912,N_4495,N_4065);
nand U7913 (N_7913,N_5122,N_5073);
nor U7914 (N_7914,N_5576,N_4868);
and U7915 (N_7915,N_5047,N_4996);
xnor U7916 (N_7916,N_4074,N_5128);
or U7917 (N_7917,N_4343,N_5735);
xnor U7918 (N_7918,N_5062,N_5083);
nor U7919 (N_7919,N_5543,N_4372);
and U7920 (N_7920,N_4561,N_4922);
nand U7921 (N_7921,N_5607,N_4793);
xnor U7922 (N_7922,N_4462,N_5672);
or U7923 (N_7923,N_4065,N_4752);
nor U7924 (N_7924,N_4885,N_5180);
nor U7925 (N_7925,N_4006,N_5557);
or U7926 (N_7926,N_5670,N_4204);
nand U7927 (N_7927,N_5058,N_4808);
nand U7928 (N_7928,N_4383,N_5860);
and U7929 (N_7929,N_4496,N_5615);
and U7930 (N_7930,N_4155,N_5977);
xor U7931 (N_7931,N_5646,N_5960);
xnor U7932 (N_7932,N_5374,N_4945);
nor U7933 (N_7933,N_4177,N_5612);
and U7934 (N_7934,N_5863,N_4004);
or U7935 (N_7935,N_4654,N_5377);
xnor U7936 (N_7936,N_4041,N_4908);
xor U7937 (N_7937,N_5966,N_5146);
or U7938 (N_7938,N_4768,N_5501);
nand U7939 (N_7939,N_5817,N_5066);
and U7940 (N_7940,N_5416,N_5928);
or U7941 (N_7941,N_5238,N_5315);
and U7942 (N_7942,N_4345,N_4593);
xor U7943 (N_7943,N_5110,N_5581);
or U7944 (N_7944,N_4369,N_4161);
nand U7945 (N_7945,N_4871,N_4799);
and U7946 (N_7946,N_5735,N_5738);
xor U7947 (N_7947,N_4994,N_4253);
or U7948 (N_7948,N_5687,N_5011);
nor U7949 (N_7949,N_4104,N_4393);
and U7950 (N_7950,N_4468,N_4770);
xor U7951 (N_7951,N_4261,N_4990);
or U7952 (N_7952,N_4147,N_4807);
nor U7953 (N_7953,N_5924,N_4919);
xnor U7954 (N_7954,N_5071,N_4398);
nand U7955 (N_7955,N_4246,N_5530);
nand U7956 (N_7956,N_5676,N_5624);
nor U7957 (N_7957,N_4311,N_4675);
and U7958 (N_7958,N_5430,N_5505);
and U7959 (N_7959,N_4324,N_5397);
nor U7960 (N_7960,N_5863,N_5034);
or U7961 (N_7961,N_5766,N_4197);
nand U7962 (N_7962,N_4689,N_4756);
and U7963 (N_7963,N_4773,N_4601);
and U7964 (N_7964,N_5611,N_4433);
nor U7965 (N_7965,N_4378,N_5703);
nor U7966 (N_7966,N_5927,N_4173);
nand U7967 (N_7967,N_4314,N_4257);
nor U7968 (N_7968,N_4349,N_4295);
or U7969 (N_7969,N_5351,N_5368);
and U7970 (N_7970,N_4920,N_4117);
or U7971 (N_7971,N_5623,N_5905);
xor U7972 (N_7972,N_5037,N_5511);
nand U7973 (N_7973,N_4020,N_5787);
nand U7974 (N_7974,N_5977,N_5224);
nor U7975 (N_7975,N_5654,N_4475);
nor U7976 (N_7976,N_4520,N_4881);
nand U7977 (N_7977,N_5624,N_4189);
nor U7978 (N_7978,N_5810,N_5607);
or U7979 (N_7979,N_4805,N_5279);
or U7980 (N_7980,N_5153,N_4991);
nor U7981 (N_7981,N_4819,N_4421);
nor U7982 (N_7982,N_4908,N_5394);
or U7983 (N_7983,N_4208,N_4064);
and U7984 (N_7984,N_4880,N_4265);
nand U7985 (N_7985,N_5596,N_5329);
and U7986 (N_7986,N_5363,N_5308);
xor U7987 (N_7987,N_4412,N_4023);
nor U7988 (N_7988,N_5945,N_5605);
and U7989 (N_7989,N_4458,N_4892);
xnor U7990 (N_7990,N_5745,N_4389);
nand U7991 (N_7991,N_5464,N_5936);
or U7992 (N_7992,N_5420,N_4043);
nand U7993 (N_7993,N_5950,N_4341);
and U7994 (N_7994,N_5669,N_5192);
or U7995 (N_7995,N_5759,N_5655);
or U7996 (N_7996,N_5653,N_5569);
xnor U7997 (N_7997,N_4628,N_4677);
nand U7998 (N_7998,N_4829,N_5858);
xor U7999 (N_7999,N_4159,N_4737);
xor U8000 (N_8000,N_7681,N_7085);
nand U8001 (N_8001,N_6281,N_6592);
xor U8002 (N_8002,N_7446,N_7495);
nor U8003 (N_8003,N_6285,N_6909);
and U8004 (N_8004,N_6942,N_7025);
nand U8005 (N_8005,N_6378,N_7518);
and U8006 (N_8006,N_7032,N_6868);
nor U8007 (N_8007,N_6036,N_6741);
nand U8008 (N_8008,N_6043,N_6199);
nand U8009 (N_8009,N_6955,N_7896);
xor U8010 (N_8010,N_7292,N_6913);
nor U8011 (N_8011,N_7321,N_6582);
and U8012 (N_8012,N_7593,N_7147);
nor U8013 (N_8013,N_6792,N_6486);
nand U8014 (N_8014,N_6538,N_7889);
nand U8015 (N_8015,N_6163,N_6459);
xor U8016 (N_8016,N_6771,N_6274);
and U8017 (N_8017,N_6827,N_7206);
or U8018 (N_8018,N_6370,N_7094);
nor U8019 (N_8019,N_7817,N_6034);
nand U8020 (N_8020,N_6910,N_6639);
nor U8021 (N_8021,N_6968,N_6540);
or U8022 (N_8022,N_6371,N_6655);
and U8023 (N_8023,N_7167,N_7275);
or U8024 (N_8024,N_7262,N_6969);
nor U8025 (N_8025,N_7810,N_7306);
nand U8026 (N_8026,N_6665,N_7371);
xnor U8027 (N_8027,N_7764,N_7506);
xnor U8028 (N_8028,N_7178,N_7568);
xor U8029 (N_8029,N_7174,N_6601);
or U8030 (N_8030,N_6580,N_6255);
nand U8031 (N_8031,N_7122,N_7710);
nor U8032 (N_8032,N_6489,N_6682);
nor U8033 (N_8033,N_6651,N_7138);
nand U8034 (N_8034,N_6694,N_7637);
or U8035 (N_8035,N_6401,N_6069);
nand U8036 (N_8036,N_7908,N_7870);
xnor U8037 (N_8037,N_6060,N_7657);
nor U8038 (N_8038,N_6515,N_6751);
xnor U8039 (N_8039,N_6294,N_6480);
and U8040 (N_8040,N_6348,N_6323);
nor U8041 (N_8041,N_6235,N_7440);
and U8042 (N_8042,N_7936,N_6385);
xnor U8043 (N_8043,N_6020,N_7418);
or U8044 (N_8044,N_7691,N_6177);
nor U8045 (N_8045,N_7591,N_6086);
and U8046 (N_8046,N_7117,N_7627);
nor U8047 (N_8047,N_6810,N_7573);
nand U8048 (N_8048,N_7902,N_7348);
nand U8049 (N_8049,N_7245,N_7822);
nand U8050 (N_8050,N_7334,N_7569);
nor U8051 (N_8051,N_7647,N_6689);
nor U8052 (N_8052,N_6330,N_7209);
nand U8053 (N_8053,N_6041,N_7932);
xnor U8054 (N_8054,N_7389,N_6795);
xor U8055 (N_8055,N_7941,N_7677);
xor U8056 (N_8056,N_7879,N_7923);
and U8057 (N_8057,N_7736,N_6088);
and U8058 (N_8058,N_7413,N_7111);
nand U8059 (N_8059,N_6625,N_6193);
xnor U8060 (N_8060,N_6584,N_6539);
and U8061 (N_8061,N_6575,N_6223);
or U8062 (N_8062,N_6988,N_7462);
or U8063 (N_8063,N_7862,N_6596);
or U8064 (N_8064,N_6074,N_6001);
and U8065 (N_8065,N_7678,N_6331);
xor U8066 (N_8066,N_6715,N_6641);
nor U8067 (N_8067,N_6799,N_7126);
and U8068 (N_8068,N_6059,N_6964);
nand U8069 (N_8069,N_6217,N_7071);
nor U8070 (N_8070,N_6202,N_6589);
nor U8071 (N_8071,N_7792,N_6624);
nand U8072 (N_8072,N_6129,N_7247);
or U8073 (N_8073,N_6372,N_7818);
nor U8074 (N_8074,N_6005,N_6408);
nor U8075 (N_8075,N_6593,N_6428);
nand U8076 (N_8076,N_7968,N_7561);
nand U8077 (N_8077,N_7915,N_6500);
and U8078 (N_8078,N_6890,N_6752);
nand U8079 (N_8079,N_6404,N_6626);
nand U8080 (N_8080,N_7123,N_6920);
nor U8081 (N_8081,N_7289,N_6781);
or U8082 (N_8082,N_7700,N_7567);
nor U8083 (N_8083,N_7294,N_6251);
nor U8084 (N_8084,N_6653,N_7885);
nor U8085 (N_8085,N_7027,N_6603);
nand U8086 (N_8086,N_7331,N_7855);
xor U8087 (N_8087,N_6835,N_6176);
xor U8088 (N_8088,N_6513,N_7435);
nand U8089 (N_8089,N_6314,N_7562);
or U8090 (N_8090,N_6338,N_7450);
nand U8091 (N_8091,N_6843,N_7175);
and U8092 (N_8092,N_7938,N_6152);
or U8093 (N_8093,N_7820,N_6073);
nand U8094 (N_8094,N_7979,N_6565);
xor U8095 (N_8095,N_7698,N_7253);
and U8096 (N_8096,N_6687,N_7999);
nand U8097 (N_8097,N_6092,N_6221);
or U8098 (N_8098,N_7617,N_7318);
and U8099 (N_8099,N_7315,N_7866);
nand U8100 (N_8100,N_6878,N_7600);
nor U8101 (N_8101,N_6622,N_6169);
xnor U8102 (N_8102,N_7127,N_6472);
nand U8103 (N_8103,N_6726,N_7758);
or U8104 (N_8104,N_7499,N_6610);
nor U8105 (N_8105,N_6308,N_6057);
nand U8106 (N_8106,N_6007,N_6766);
nor U8107 (N_8107,N_7816,N_6818);
nand U8108 (N_8108,N_6772,N_6194);
nor U8109 (N_8109,N_7464,N_6307);
and U8110 (N_8110,N_6570,N_7179);
nand U8111 (N_8111,N_7091,N_6723);
nand U8112 (N_8112,N_7981,N_7566);
and U8113 (N_8113,N_6290,N_6786);
nor U8114 (N_8114,N_6244,N_6344);
xor U8115 (N_8115,N_7218,N_7695);
xnor U8116 (N_8116,N_6851,N_7633);
or U8117 (N_8117,N_7326,N_6106);
nor U8118 (N_8118,N_7353,N_6932);
or U8119 (N_8119,N_6979,N_6548);
nand U8120 (N_8120,N_7546,N_7096);
and U8121 (N_8121,N_6309,N_6926);
xor U8122 (N_8122,N_6928,N_7782);
nor U8123 (N_8123,N_6735,N_6286);
and U8124 (N_8124,N_7286,N_7631);
xnor U8125 (N_8125,N_6405,N_6514);
or U8126 (N_8126,N_6268,N_6118);
nand U8127 (N_8127,N_7263,N_7121);
nor U8128 (N_8128,N_6329,N_6122);
xor U8129 (N_8129,N_6649,N_6228);
and U8130 (N_8130,N_6559,N_6219);
and U8131 (N_8131,N_6081,N_6119);
xnor U8132 (N_8132,N_6398,N_6383);
xnor U8133 (N_8133,N_6478,N_7594);
and U8134 (N_8134,N_6266,N_6637);
and U8135 (N_8135,N_6809,N_7165);
xnor U8136 (N_8136,N_6275,N_7944);
and U8137 (N_8137,N_6707,N_6600);
xor U8138 (N_8138,N_7552,N_6393);
nand U8139 (N_8139,N_6718,N_6166);
and U8140 (N_8140,N_6941,N_6820);
nor U8141 (N_8141,N_6618,N_6846);
and U8142 (N_8142,N_7125,N_7581);
xnor U8143 (N_8143,N_6499,N_7806);
xnor U8144 (N_8144,N_7737,N_6927);
or U8145 (N_8145,N_6550,N_6120);
nor U8146 (N_8146,N_7007,N_7220);
or U8147 (N_8147,N_6117,N_6949);
or U8148 (N_8148,N_7217,N_7124);
nand U8149 (N_8149,N_6467,N_7844);
nor U8150 (N_8150,N_6922,N_7078);
nor U8151 (N_8151,N_7293,N_7578);
or U8152 (N_8152,N_6136,N_7898);
or U8153 (N_8153,N_6667,N_7668);
or U8154 (N_8154,N_6033,N_7201);
nand U8155 (N_8155,N_7717,N_6834);
nor U8156 (N_8156,N_6142,N_6961);
nand U8157 (N_8157,N_7216,N_6231);
nor U8158 (N_8158,N_6191,N_6278);
xnor U8159 (N_8159,N_6306,N_7531);
nor U8160 (N_8160,N_7441,N_7564);
xor U8161 (N_8161,N_7018,N_6067);
nand U8162 (N_8162,N_7432,N_6644);
and U8163 (N_8163,N_7237,N_6110);
xnor U8164 (N_8164,N_7946,N_6054);
and U8165 (N_8165,N_6506,N_7204);
and U8166 (N_8166,N_6479,N_7359);
nand U8167 (N_8167,N_7757,N_6985);
or U8168 (N_8168,N_6825,N_7159);
nand U8169 (N_8169,N_7040,N_6497);
or U8170 (N_8170,N_6699,N_7059);
nor U8171 (N_8171,N_7261,N_6155);
or U8172 (N_8172,N_7052,N_6319);
nor U8173 (N_8173,N_7832,N_6026);
and U8174 (N_8174,N_6493,N_6945);
xnor U8175 (N_8175,N_7192,N_6183);
xor U8176 (N_8176,N_7228,N_6149);
xnor U8177 (N_8177,N_6396,N_7433);
xnor U8178 (N_8178,N_6635,N_7154);
xor U8179 (N_8179,N_6324,N_6099);
nand U8180 (N_8180,N_6115,N_7360);
and U8181 (N_8181,N_6638,N_6414);
or U8182 (N_8182,N_7718,N_6468);
or U8183 (N_8183,N_7422,N_7576);
nor U8184 (N_8184,N_6018,N_7990);
nor U8185 (N_8185,N_6794,N_6660);
and U8186 (N_8186,N_6808,N_6530);
and U8187 (N_8187,N_6279,N_7749);
nor U8188 (N_8188,N_7417,N_6289);
nand U8189 (N_8189,N_7730,N_6946);
xor U8190 (N_8190,N_7470,N_7434);
nor U8191 (N_8191,N_7533,N_7128);
and U8192 (N_8192,N_7451,N_6688);
and U8193 (N_8193,N_6542,N_7170);
or U8194 (N_8194,N_6146,N_7625);
nand U8195 (N_8195,N_7163,N_7794);
nor U8196 (N_8196,N_7282,N_6953);
or U8197 (N_8197,N_6543,N_6079);
or U8198 (N_8198,N_7504,N_6528);
nor U8199 (N_8199,N_7363,N_6390);
nor U8200 (N_8200,N_7398,N_6705);
and U8201 (N_8201,N_6245,N_7021);
nor U8202 (N_8202,N_7234,N_7519);
nand U8203 (N_8203,N_7966,N_7256);
nor U8204 (N_8204,N_6788,N_6025);
and U8205 (N_8205,N_7692,N_6536);
and U8206 (N_8206,N_7784,N_6813);
and U8207 (N_8207,N_7543,N_7939);
or U8208 (N_8208,N_6270,N_6729);
nor U8209 (N_8209,N_7497,N_7004);
or U8210 (N_8210,N_6661,N_6773);
xnor U8211 (N_8211,N_6426,N_6966);
xor U8212 (N_8212,N_6240,N_6819);
nor U8213 (N_8213,N_6483,N_6925);
nand U8214 (N_8214,N_7424,N_7300);
nor U8215 (N_8215,N_6389,N_7912);
or U8216 (N_8216,N_7488,N_6350);
xnor U8217 (N_8217,N_7368,N_6168);
and U8218 (N_8218,N_6458,N_7055);
and U8219 (N_8219,N_7624,N_7346);
xor U8220 (N_8220,N_7317,N_6755);
nor U8221 (N_8221,N_7804,N_6312);
nor U8222 (N_8222,N_7868,N_6157);
and U8223 (N_8223,N_7861,N_6271);
and U8224 (N_8224,N_6900,N_7354);
xnor U8225 (N_8225,N_6934,N_6828);
or U8226 (N_8226,N_7976,N_7250);
nor U8227 (N_8227,N_6963,N_7874);
or U8228 (N_8228,N_7148,N_7195);
and U8229 (N_8229,N_6779,N_6494);
or U8230 (N_8230,N_7189,N_6887);
or U8231 (N_8231,N_7707,N_6679);
nand U8232 (N_8232,N_6031,N_7310);
or U8233 (N_8233,N_7375,N_7260);
nor U8234 (N_8234,N_7574,N_7232);
or U8235 (N_8235,N_6140,N_6357);
nor U8236 (N_8236,N_7913,N_6447);
and U8237 (N_8237,N_6162,N_7520);
xnor U8238 (N_8238,N_7184,N_7740);
nand U8239 (N_8239,N_7399,N_6989);
nor U8240 (N_8240,N_6195,N_7558);
and U8241 (N_8241,N_7865,N_6429);
or U8242 (N_8242,N_7509,N_7729);
and U8243 (N_8243,N_6366,N_7157);
and U8244 (N_8244,N_6154,N_6583);
xnor U8245 (N_8245,N_7008,N_6365);
nand U8246 (N_8246,N_7928,N_7061);
and U8247 (N_8247,N_6433,N_7425);
xor U8248 (N_8248,N_7809,N_7419);
nand U8249 (N_8249,N_7102,N_7489);
nand U8250 (N_8250,N_6631,N_7609);
nand U8251 (N_8251,N_7408,N_6421);
xnor U8252 (N_8252,N_6091,N_7683);
nor U8253 (N_8253,N_6950,N_7064);
nor U8254 (N_8254,N_7168,N_6427);
and U8255 (N_8255,N_6008,N_7382);
nand U8256 (N_8256,N_6455,N_7927);
xnor U8257 (N_8257,N_6711,N_6521);
nand U8258 (N_8258,N_7442,N_6347);
and U8259 (N_8259,N_7444,N_7301);
or U8260 (N_8260,N_7502,N_6380);
and U8261 (N_8261,N_7200,N_7828);
and U8262 (N_8262,N_7257,N_6367);
and U8263 (N_8263,N_6713,N_6829);
nor U8264 (N_8264,N_7396,N_7841);
or U8265 (N_8265,N_7194,N_6407);
or U8266 (N_8266,N_7635,N_7980);
and U8267 (N_8267,N_7795,N_7051);
nand U8268 (N_8268,N_6643,N_6211);
nor U8269 (N_8269,N_7421,N_6438);
and U8270 (N_8270,N_7093,N_7113);
nor U8271 (N_8271,N_7798,N_7383);
xor U8272 (N_8272,N_6368,N_6084);
or U8273 (N_8273,N_7663,N_7670);
or U8274 (N_8274,N_7611,N_7385);
and U8275 (N_8275,N_6475,N_6340);
nor U8276 (N_8276,N_7974,N_7241);
nand U8277 (N_8277,N_6719,N_7233);
nand U8278 (N_8278,N_7490,N_6229);
nand U8279 (N_8279,N_6800,N_7338);
or U8280 (N_8280,N_7314,N_6097);
or U8281 (N_8281,N_7997,N_7967);
or U8282 (N_8282,N_6919,N_6571);
xor U8283 (N_8283,N_6139,N_7373);
xnor U8284 (N_8284,N_7665,N_6151);
nor U8285 (N_8285,N_7409,N_6743);
xnor U8286 (N_8286,N_6864,N_7231);
and U8287 (N_8287,N_6113,N_6381);
and U8288 (N_8288,N_7541,N_7254);
nand U8289 (N_8289,N_6466,N_6066);
nand U8290 (N_8290,N_7406,N_7544);
and U8291 (N_8291,N_7522,N_7099);
nand U8292 (N_8292,N_6617,N_7297);
or U8293 (N_8293,N_6870,N_6234);
and U8294 (N_8294,N_7449,N_7696);
nand U8295 (N_8295,N_6412,N_7640);
xor U8296 (N_8296,N_6470,N_6696);
nand U8297 (N_8297,N_7176,N_7847);
nor U8298 (N_8298,N_6490,N_7427);
and U8299 (N_8299,N_6673,N_7793);
xor U8300 (N_8300,N_7738,N_6836);
nor U8301 (N_8301,N_6262,N_7395);
nor U8302 (N_8302,N_7347,N_6708);
or U8303 (N_8303,N_6161,N_6220);
nand U8304 (N_8304,N_7416,N_6052);
nor U8305 (N_8305,N_6534,N_7252);
and U8306 (N_8306,N_6701,N_7136);
and U8307 (N_8307,N_6449,N_6205);
nor U8308 (N_8308,N_7158,N_7890);
nor U8309 (N_8309,N_7517,N_6448);
and U8310 (N_8310,N_7343,N_7208);
nand U8311 (N_8311,N_6529,N_7959);
nand U8312 (N_8312,N_7074,N_7788);
xnor U8313 (N_8313,N_6894,N_6675);
or U8314 (N_8314,N_7598,N_7744);
and U8315 (N_8315,N_7903,N_7634);
nand U8316 (N_8316,N_6325,N_6022);
and U8317 (N_8317,N_7177,N_6869);
and U8318 (N_8318,N_7088,N_7856);
and U8319 (N_8319,N_6572,N_6179);
nor U8320 (N_8320,N_6908,N_6297);
nand U8321 (N_8321,N_7769,N_7243);
nand U8322 (N_8322,N_7374,N_7151);
xor U8323 (N_8323,N_6931,N_7777);
nor U8324 (N_8324,N_6442,N_6986);
nand U8325 (N_8325,N_7534,N_6085);
and U8326 (N_8326,N_6105,N_6328);
and U8327 (N_8327,N_6853,N_6840);
and U8328 (N_8328,N_7947,N_6602);
xnor U8329 (N_8329,N_7080,N_6216);
and U8330 (N_8330,N_6629,N_6315);
or U8331 (N_8331,N_6754,N_6634);
or U8332 (N_8332,N_6895,N_7929);
nor U8333 (N_8333,N_6201,N_6188);
nand U8334 (N_8334,N_6874,N_7619);
nand U8335 (N_8335,N_6349,N_6903);
or U8336 (N_8336,N_6024,N_7833);
nor U8337 (N_8337,N_6065,N_7709);
nor U8338 (N_8338,N_6346,N_6141);
xnor U8339 (N_8339,N_7370,N_7863);
and U8340 (N_8340,N_6498,N_6127);
or U8341 (N_8341,N_7762,N_6473);
nor U8342 (N_8342,N_7473,N_7400);
nor U8343 (N_8343,N_7152,N_7791);
nand U8344 (N_8344,N_6068,N_7831);
and U8345 (N_8345,N_7998,N_6303);
nor U8346 (N_8346,N_7423,N_7397);
nor U8347 (N_8347,N_6430,N_6012);
nor U8348 (N_8348,N_7595,N_6173);
nor U8349 (N_8349,N_7101,N_6518);
or U8350 (N_8350,N_7024,N_6558);
xor U8351 (N_8351,N_7039,N_6793);
xor U8352 (N_8352,N_7073,N_6588);
or U8353 (N_8353,N_7662,N_7020);
nand U8354 (N_8354,N_7336,N_7477);
nor U8355 (N_8355,N_7750,N_7349);
nand U8356 (N_8356,N_7770,N_6263);
or U8357 (N_8357,N_7824,N_7867);
or U8358 (N_8358,N_7800,N_6881);
nand U8359 (N_8359,N_6992,N_7642);
or U8360 (N_8360,N_7493,N_6855);
nor U8361 (N_8361,N_7530,N_7249);
nand U8362 (N_8362,N_7725,N_6636);
nor U8363 (N_8363,N_6153,N_7814);
xor U8364 (N_8364,N_7323,N_7259);
xor U8365 (N_8365,N_7853,N_6083);
xnor U8366 (N_8366,N_6444,N_6877);
and U8367 (N_8367,N_6717,N_6889);
nor U8368 (N_8368,N_7081,N_7952);
xnor U8369 (N_8369,N_6627,N_6783);
nor U8370 (N_8370,N_6171,N_7687);
xor U8371 (N_8371,N_6898,N_7162);
xnor U8372 (N_8372,N_7046,N_6050);
and U8373 (N_8373,N_6481,N_6510);
or U8374 (N_8374,N_6545,N_6854);
nor U8375 (N_8375,N_7675,N_6292);
xnor U8376 (N_8376,N_7618,N_6100);
xnor U8377 (N_8377,N_7210,N_7084);
and U8378 (N_8378,N_6677,N_7356);
xor U8379 (N_8379,N_6190,N_6042);
and U8380 (N_8380,N_6023,N_6039);
nor U8381 (N_8381,N_7813,N_7012);
xor U8382 (N_8382,N_7106,N_7789);
xor U8383 (N_8383,N_6769,N_7638);
nor U8384 (N_8384,N_7056,N_6006);
and U8385 (N_8385,N_7143,N_6078);
nor U8386 (N_8386,N_7621,N_6048);
nand U8387 (N_8387,N_7741,N_6958);
or U8388 (N_8388,N_6124,N_7689);
or U8389 (N_8389,N_7671,N_7926);
nor U8390 (N_8390,N_6339,N_7183);
nand U8391 (N_8391,N_6310,N_7654);
and U8392 (N_8392,N_6607,N_7703);
xor U8393 (N_8393,N_6577,N_6464);
or U8394 (N_8394,N_7258,N_7715);
nor U8395 (N_8395,N_6956,N_6880);
or U8396 (N_8396,N_7100,N_7602);
or U8397 (N_8397,N_7511,N_6995);
xor U8398 (N_8398,N_6574,N_6852);
nand U8399 (N_8399,N_6206,N_7065);
nor U8400 (N_8400,N_7212,N_7588);
nand U8401 (N_8401,N_7414,N_7494);
or U8402 (N_8402,N_7554,N_7501);
nor U8403 (N_8403,N_6905,N_7335);
nor U8404 (N_8404,N_6859,N_6112);
or U8405 (N_8405,N_7508,N_7510);
or U8406 (N_8406,N_7897,N_6976);
nor U8407 (N_8407,N_7628,N_6823);
nand U8408 (N_8408,N_7332,N_7022);
and U8409 (N_8409,N_7267,N_6761);
nor U8410 (N_8410,N_7983,N_6247);
xnor U8411 (N_8411,N_6731,N_6361);
nand U8412 (N_8412,N_7134,N_6495);
xor U8413 (N_8413,N_7607,N_6947);
nor U8414 (N_8414,N_7743,N_7222);
and U8415 (N_8415,N_7190,N_7872);
or U8416 (N_8416,N_6971,N_6482);
nand U8417 (N_8417,N_7901,N_7626);
and U8418 (N_8418,N_6114,N_7771);
or U8419 (N_8419,N_7823,N_7783);
nand U8420 (N_8420,N_7010,N_7120);
xnor U8421 (N_8421,N_7072,N_7387);
or U8422 (N_8422,N_6107,N_6998);
nand U8423 (N_8423,N_6875,N_6130);
or U8424 (N_8424,N_7001,N_6628);
and U8425 (N_8425,N_6032,N_6132);
xnor U8426 (N_8426,N_6553,N_7949);
and U8427 (N_8427,N_7112,N_6299);
nand U8428 (N_8428,N_7994,N_6431);
or U8429 (N_8429,N_7644,N_6720);
nand U8430 (N_8430,N_6035,N_6884);
and U8431 (N_8431,N_6222,N_7391);
nand U8432 (N_8432,N_7615,N_6451);
or U8433 (N_8433,N_6460,N_7236);
nor U8434 (N_8434,N_7726,N_6280);
or U8435 (N_8435,N_6453,N_6849);
or U8436 (N_8436,N_7060,N_7679);
xor U8437 (N_8437,N_6561,N_6358);
nand U8438 (N_8438,N_6917,N_6335);
xnor U8439 (N_8439,N_7606,N_7616);
nor U8440 (N_8440,N_7603,N_6203);
nand U8441 (N_8441,N_6496,N_7098);
nor U8442 (N_8442,N_6282,N_7688);
nand U8443 (N_8443,N_7471,N_6776);
nor U8444 (N_8444,N_7169,N_6876);
xnor U8445 (N_8445,N_6170,N_7977);
nand U8446 (N_8446,N_7797,N_6376);
xnor U8447 (N_8447,N_7653,N_7719);
xor U8448 (N_8448,N_7467,N_7888);
nor U8449 (N_8449,N_6445,N_6936);
nor U8450 (N_8450,N_6027,N_6778);
xnor U8451 (N_8451,N_6058,N_6184);
xnor U8452 (N_8452,N_6304,N_6664);
nand U8453 (N_8453,N_7328,N_7532);
and U8454 (N_8454,N_6797,N_6695);
or U8455 (N_8455,N_7116,N_6413);
nand U8456 (N_8456,N_6844,N_6929);
nand U8457 (N_8457,N_6952,N_7951);
xor U8458 (N_8458,N_6526,N_7887);
xor U8459 (N_8459,N_7575,N_6566);
nand U8460 (N_8460,N_7436,N_7956);
or U8461 (N_8461,N_6562,N_7058);
xor U8462 (N_8462,N_7693,N_6509);
and U8463 (N_8463,N_6260,N_7295);
or U8464 (N_8464,N_7720,N_6104);
nand U8465 (N_8465,N_7225,N_6138);
and U8466 (N_8466,N_7587,N_6017);
nor U8467 (N_8467,N_7028,N_7858);
and U8468 (N_8468,N_7655,N_7622);
nand U8469 (N_8469,N_7316,N_7649);
nand U8470 (N_8470,N_7054,N_7840);
and U8471 (N_8471,N_6745,N_7954);
and U8472 (N_8472,N_7579,N_6321);
or U8473 (N_8473,N_6879,N_6135);
and U8474 (N_8474,N_6283,N_7596);
nor U8475 (N_8475,N_7728,N_6614);
nor U8476 (N_8476,N_7911,N_7202);
nand U8477 (N_8477,N_6857,N_6507);
nor U8478 (N_8478,N_6541,N_7992);
nand U8479 (N_8479,N_7131,N_6906);
xor U8480 (N_8480,N_7223,N_6080);
and U8481 (N_8481,N_6108,N_7401);
nand U8482 (N_8482,N_7110,N_7067);
nand U8483 (N_8483,N_7474,N_6739);
nand U8484 (N_8484,N_6567,N_6750);
nand U8485 (N_8485,N_7843,N_7276);
nand U8486 (N_8486,N_6456,N_6450);
nand U8487 (N_8487,N_7246,N_6975);
nand U8488 (N_8488,N_6832,N_7961);
and U8489 (N_8489,N_6210,N_6681);
nor U8490 (N_8490,N_7458,N_7215);
or U8491 (N_8491,N_6016,N_6248);
nor U8492 (N_8492,N_7312,N_7849);
or U8493 (N_8493,N_6186,N_7993);
xor U8494 (N_8494,N_7364,N_6014);
and U8495 (N_8495,N_6666,N_6208);
nor U8496 (N_8496,N_6897,N_7555);
nor U8497 (N_8497,N_7457,N_7407);
xnor U8498 (N_8498,N_7308,N_6838);
or U8499 (N_8499,N_6640,N_7825);
and U8500 (N_8500,N_7014,N_7592);
xor U8501 (N_8501,N_7731,N_6693);
xor U8502 (N_8502,N_6970,N_7732);
nand U8503 (N_8503,N_7448,N_7761);
nor U8504 (N_8504,N_7808,N_7235);
and U8505 (N_8505,N_6753,N_7724);
or U8506 (N_8506,N_7482,N_6264);
and U8507 (N_8507,N_7713,N_7412);
xnor U8508 (N_8508,N_7133,N_6646);
nor U8509 (N_8509,N_7727,N_7006);
or U8510 (N_8510,N_6243,N_7632);
and U8511 (N_8511,N_6273,N_6295);
nand U8512 (N_8512,N_7239,N_6525);
and U8513 (N_8513,N_6609,N_6556);
nor U8514 (N_8514,N_6209,N_6727);
or U8515 (N_8515,N_6990,N_6563);
and U8516 (N_8516,N_6167,N_6446);
xnor U8517 (N_8517,N_6336,N_7563);
nand U8518 (N_8518,N_6103,N_6476);
nand U8519 (N_8519,N_7048,N_6848);
and U8520 (N_8520,N_6569,N_7722);
and U8521 (N_8521,N_6821,N_6356);
and U8522 (N_8522,N_7937,N_7390);
xor U8523 (N_8523,N_7033,N_6246);
and U8524 (N_8524,N_7213,N_7785);
and U8525 (N_8525,N_7404,N_6804);
xor U8526 (N_8526,N_6736,N_7584);
nor U8527 (N_8527,N_7819,N_7229);
xor U8528 (N_8528,N_7381,N_7763);
or U8529 (N_8529,N_6882,N_7641);
xor U8530 (N_8530,N_6301,N_7549);
and U8531 (N_8531,N_6252,N_6757);
or U8532 (N_8532,N_7790,N_7924);
nor U8533 (N_8533,N_7023,N_6488);
nor U8534 (N_8534,N_7747,N_7430);
xnor U8535 (N_8535,N_7883,N_6212);
or U8536 (N_8536,N_7188,N_6733);
xnor U8537 (N_8537,N_6463,N_6796);
nand U8538 (N_8538,N_6242,N_6126);
nor U8539 (N_8539,N_7766,N_6215);
or U8540 (N_8540,N_6517,N_7786);
and U8541 (N_8541,N_7753,N_6109);
xnor U8542 (N_8542,N_6265,N_7917);
and U8543 (N_8543,N_6053,N_6822);
and U8544 (N_8544,N_6999,N_7324);
or U8545 (N_8545,N_6004,N_7812);
or U8546 (N_8546,N_6474,N_7650);
and U8547 (N_8547,N_7108,N_7320);
xor U8548 (N_8548,N_7850,N_7283);
xor U8549 (N_8549,N_6684,N_6269);
and U8550 (N_8550,N_7461,N_6669);
nand U8551 (N_8551,N_6387,N_6734);
xnor U8552 (N_8552,N_6598,N_6038);
and U8553 (N_8553,N_6659,N_7103);
nor U8554 (N_8554,N_7551,N_7015);
and U8555 (N_8555,N_7105,N_6391);
xnor U8556 (N_8556,N_7978,N_6015);
or U8557 (N_8557,N_6354,N_7305);
xor U8558 (N_8558,N_7439,N_7337);
nor U8559 (N_8559,N_7164,N_6411);
and U8560 (N_8560,N_7900,N_6148);
nor U8561 (N_8561,N_6856,N_7034);
xnor U8562 (N_8562,N_6984,N_7884);
or U8563 (N_8563,N_7601,N_6872);
xor U8564 (N_8564,N_6585,N_7107);
or U8565 (N_8565,N_7585,N_6419);
nand U8566 (N_8566,N_6576,N_7571);
or U8567 (N_8567,N_6409,N_6896);
nand U8568 (N_8568,N_6133,N_7226);
xor U8569 (N_8569,N_6613,N_6327);
and U8570 (N_8570,N_6866,N_7772);
and U8571 (N_8571,N_6993,N_6709);
nor U8572 (N_8572,N_7559,N_7660);
and U8573 (N_8573,N_7057,N_6817);
or U8574 (N_8574,N_7708,N_7669);
xor U8575 (N_8575,N_6826,N_7219);
nand U8576 (N_8576,N_7492,N_7921);
and U8577 (N_8577,N_7197,N_7699);
and U8578 (N_8578,N_7153,N_6805);
nor U8579 (N_8579,N_7859,N_6317);
nand U8580 (N_8580,N_7659,N_6440);
nand U8581 (N_8581,N_7077,N_6615);
nand U8582 (N_8582,N_6288,N_7765);
xor U8583 (N_8583,N_7857,N_6604);
nor U8584 (N_8584,N_7620,N_6322);
nand U8585 (N_8585,N_6523,N_6973);
nor U8586 (N_8586,N_7339,N_7577);
nand U8587 (N_8587,N_7542,N_7527);
or U8588 (N_8588,N_6037,N_7330);
nand U8589 (N_8589,N_6061,N_7964);
xor U8590 (N_8590,N_7960,N_6980);
nor U8591 (N_8591,N_6977,N_6663);
and U8592 (N_8592,N_7049,N_7636);
nor U8593 (N_8593,N_7227,N_7666);
and U8594 (N_8594,N_7751,N_7672);
nor U8595 (N_8595,N_6902,N_6400);
and U8596 (N_8596,N_6134,N_7973);
nor U8597 (N_8597,N_7376,N_6316);
or U8598 (N_8598,N_7523,N_6690);
and U8599 (N_8599,N_6801,N_7582);
xnor U8600 (N_8600,N_6076,N_7196);
and U8601 (N_8601,N_7775,N_6180);
nand U8602 (N_8602,N_7876,N_6916);
or U8603 (N_8603,N_7676,N_6862);
xnor U8604 (N_8604,N_7428,N_6768);
xor U8605 (N_8605,N_7714,N_7705);
or U8606 (N_8606,N_7643,N_6258);
or U8607 (N_8607,N_7271,N_7934);
nor U8608 (N_8608,N_7807,N_6143);
nor U8609 (N_8609,N_7274,N_7536);
xnor U8610 (N_8610,N_7919,N_7362);
xnor U8611 (N_8611,N_6597,N_6991);
or U8612 (N_8612,N_6774,N_6386);
and U8613 (N_8613,N_7851,N_6738);
nor U8614 (N_8614,N_6554,N_6164);
or U8615 (N_8615,N_6355,N_7694);
or U8616 (N_8616,N_6044,N_6730);
nor U8617 (N_8617,N_6721,N_7266);
and U8618 (N_8618,N_6824,N_6686);
nand U8619 (N_8619,N_7244,N_6392);
nand U8620 (N_8620,N_6095,N_6533);
or U8621 (N_8621,N_6182,N_7599);
xnor U8622 (N_8622,N_7918,N_6291);
nand U8623 (N_8623,N_7984,N_7514);
and U8624 (N_8624,N_7988,N_6441);
or U8625 (N_8625,N_6865,N_7878);
nand U8626 (N_8626,N_7827,N_7351);
nand U8627 (N_8627,N_7701,N_7557);
nor U8628 (N_8628,N_6842,N_7475);
and U8629 (N_8629,N_7472,N_6485);
nand U8630 (N_8630,N_7799,N_7975);
nand U8631 (N_8631,N_7466,N_6200);
and U8632 (N_8632,N_6363,N_6704);
and U8633 (N_8633,N_7447,N_6384);
nor U8634 (N_8634,N_6535,N_7721);
nand U8635 (N_8635,N_6944,N_7341);
nor U8636 (N_8636,N_7146,N_6587);
xnor U8637 (N_8637,N_6030,N_6402);
or U8638 (N_8638,N_6487,N_7597);
xor U8639 (N_8639,N_6131,N_7986);
xor U8640 (N_8640,N_6951,N_6524);
nor U8641 (N_8641,N_6352,N_7943);
nor U8642 (N_8642,N_6320,N_7240);
and U8643 (N_8643,N_6224,N_7047);
or U8644 (N_8644,N_7042,N_7521);
nand U8645 (N_8645,N_6937,N_6477);
xnor U8646 (N_8646,N_6253,N_7016);
or U8647 (N_8647,N_6207,N_6029);
nor U8648 (N_8648,N_6454,N_6395);
and U8649 (N_8649,N_7656,N_6353);
and U8650 (N_8650,N_7925,N_6332);
nor U8651 (N_8651,N_7759,N_6147);
nand U8652 (N_8652,N_7478,N_6861);
xnor U8653 (N_8653,N_6159,N_7892);
nand U8654 (N_8654,N_7480,N_7465);
nand U8655 (N_8655,N_6983,N_7019);
nor U8656 (N_8656,N_6049,N_6537);
or U8657 (N_8657,N_7269,N_7942);
or U8658 (N_8658,N_7392,N_7242);
nand U8659 (N_8659,N_6833,N_6519);
nor U8660 (N_8660,N_7604,N_7104);
xor U8661 (N_8661,N_7130,N_7166);
xnor U8662 (N_8662,N_6225,N_6187);
xor U8663 (N_8663,N_6551,N_7674);
xnor U8664 (N_8664,N_6863,N_6780);
nor U8665 (N_8665,N_7716,N_6650);
nor U8666 (N_8666,N_7463,N_6296);
nor U8667 (N_8667,N_7614,N_6382);
xnor U8668 (N_8668,N_6318,N_7281);
nand U8669 (N_8669,N_7526,N_6599);
nor U8670 (N_8670,N_6098,N_7528);
nand U8671 (N_8671,N_6375,N_6710);
xnor U8672 (N_8672,N_7752,N_6962);
xnor U8673 (N_8673,N_7648,N_6415);
or U8674 (N_8674,N_7629,N_7503);
and U8675 (N_8675,N_6259,N_7835);
nand U8676 (N_8676,N_7076,N_6045);
xnor U8677 (N_8677,N_7891,N_6237);
and U8678 (N_8678,N_7150,N_6172);
xnor U8679 (N_8679,N_7875,N_7394);
and U8680 (N_8680,N_6656,N_7333);
or U8681 (N_8681,N_6013,N_6775);
nor U8682 (N_8682,N_7583,N_6341);
and U8683 (N_8683,N_6055,N_7156);
nor U8684 (N_8684,N_7685,N_6806);
and U8685 (N_8685,N_6557,N_7483);
xor U8686 (N_8686,N_6439,N_7882);
nor U8687 (N_8687,N_6434,N_6333);
xor U8688 (N_8688,N_6724,N_7288);
nor U8689 (N_8689,N_6002,N_6912);
xor U8690 (N_8690,N_7155,N_7410);
and U8691 (N_8691,N_6612,N_6123);
and U8692 (N_8692,N_6935,N_7075);
nor U8693 (N_8693,N_6648,N_6578);
and U8694 (N_8694,N_7319,N_7299);
nand U8695 (N_8695,N_6605,N_6933);
and U8696 (N_8696,N_6764,N_7755);
or U8697 (N_8697,N_6397,N_7350);
or U8698 (N_8698,N_6740,N_7963);
and U8699 (N_8699,N_6606,N_7895);
nand U8700 (N_8700,N_7781,N_7735);
and U8701 (N_8701,N_7268,N_6505);
nor U8702 (N_8702,N_7070,N_6591);
or U8703 (N_8703,N_6616,N_7612);
and U8704 (N_8704,N_7667,N_6311);
nor U8705 (N_8705,N_6070,N_7608);
nand U8706 (N_8706,N_7512,N_7141);
and U8707 (N_8707,N_7264,N_6581);
or U8708 (N_8708,N_6732,N_6047);
xor U8709 (N_8709,N_6680,N_7011);
or U8710 (N_8710,N_6165,N_7469);
and U8711 (N_8711,N_6749,N_7545);
xnor U8712 (N_8712,N_6185,N_6632);
nor U8713 (N_8713,N_7953,N_6457);
xor U8714 (N_8714,N_6728,N_6373);
or U8715 (N_8715,N_6267,N_7415);
or U8716 (N_8716,N_6249,N_6345);
nor U8717 (N_8717,N_6192,N_7114);
nor U8718 (N_8718,N_6888,N_7090);
nor U8719 (N_8719,N_7205,N_6313);
or U8720 (N_8720,N_6512,N_6918);
nand U8721 (N_8721,N_7965,N_7702);
and U8722 (N_8722,N_6594,N_7658);
or U8723 (N_8723,N_6608,N_7538);
xnor U8724 (N_8724,N_6051,N_6198);
nand U8725 (N_8725,N_7712,N_6342);
nand U8726 (N_8726,N_7684,N_7664);
xor U8727 (N_8727,N_6683,N_6867);
nand U8728 (N_8728,N_6546,N_7043);
xnor U8729 (N_8729,N_7826,N_7661);
and U8730 (N_8730,N_7411,N_7109);
nor U8731 (N_8731,N_7476,N_7767);
xnor U8732 (N_8732,N_6620,N_6484);
nand U8733 (N_8733,N_7255,N_6742);
nand U8734 (N_8734,N_6700,N_6798);
xnor U8735 (N_8735,N_6090,N_6850);
and U8736 (N_8736,N_7864,N_7680);
and U8737 (N_8737,N_6790,N_7733);
and U8738 (N_8738,N_7115,N_7224);
nand U8739 (N_8739,N_7068,N_6676);
or U8740 (N_8740,N_7848,N_7186);
xnor U8741 (N_8741,N_7342,N_6845);
and U8742 (N_8742,N_6337,N_7000);
xor U8743 (N_8743,N_6549,N_6360);
xor U8744 (N_8744,N_7445,N_6914);
xnor U8745 (N_8745,N_6250,N_7854);
or U8746 (N_8746,N_7340,N_7311);
or U8747 (N_8747,N_7906,N_7935);
xor U8748 (N_8748,N_7029,N_6831);
nor U8749 (N_8749,N_7904,N_7087);
and U8750 (N_8750,N_6272,N_7948);
or U8751 (N_8751,N_6560,N_6394);
xnor U8752 (N_8752,N_7193,N_7063);
and U8753 (N_8753,N_7673,N_6452);
or U8754 (N_8754,N_6573,N_7429);
and U8755 (N_8755,N_7086,N_6967);
and U8756 (N_8756,N_6491,N_7172);
nand U8757 (N_8757,N_7605,N_7570);
nor U8758 (N_8758,N_6420,N_6028);
xnor U8759 (N_8759,N_6364,N_6837);
or U8760 (N_8760,N_7378,N_6516);
nor U8761 (N_8761,N_6277,N_6997);
and U8762 (N_8762,N_6101,N_6532);
or U8763 (N_8763,N_6959,N_6416);
nor U8764 (N_8764,N_6232,N_6178);
nand U8765 (N_8765,N_7296,N_6662);
xnor U8766 (N_8766,N_6326,N_7893);
and U8767 (N_8767,N_7357,N_6657);
and U8768 (N_8768,N_6841,N_7610);
or U8769 (N_8769,N_6071,N_7646);
xnor U8770 (N_8770,N_6907,N_7529);
nand U8771 (N_8771,N_6082,N_6144);
nor U8772 (N_8772,N_6697,N_6175);
and U8773 (N_8773,N_6712,N_7369);
nor U8774 (N_8774,N_7871,N_7013);
xnor U8775 (N_8775,N_6714,N_7524);
nand U8776 (N_8776,N_6939,N_6145);
nor U8777 (N_8777,N_6116,N_6672);
nand U8778 (N_8778,N_6586,N_7930);
or U8779 (N_8779,N_6938,N_7214);
nand U8780 (N_8780,N_6077,N_6544);
and U8781 (N_8781,N_7203,N_6789);
or U8782 (N_8782,N_7834,N_7539);
nand U8783 (N_8783,N_6374,N_7639);
and U8784 (N_8784,N_6046,N_7773);
xnor U8785 (N_8785,N_6089,N_7515);
or U8786 (N_8786,N_7460,N_7748);
xor U8787 (N_8787,N_7149,N_7756);
nand U8788 (N_8788,N_6125,N_6424);
or U8789 (N_8789,N_6087,N_6334);
or U8790 (N_8790,N_6150,N_6359);
nand U8791 (N_8791,N_7907,N_6972);
and U8792 (N_8792,N_6633,N_6181);
or U8793 (N_8793,N_7985,N_6765);
nor U8794 (N_8794,N_7438,N_7129);
nor U8795 (N_8795,N_6611,N_7066);
xor U8796 (N_8796,N_7651,N_7774);
and U8797 (N_8797,N_7537,N_6527);
or U8798 (N_8798,N_6362,N_6522);
xor U8799 (N_8799,N_7734,N_6432);
xor U8800 (N_8800,N_7050,N_6093);
nand U8801 (N_8801,N_6568,N_7931);
xnor U8802 (N_8802,N_6784,N_6994);
and U8803 (N_8803,N_6737,N_6064);
nor U8804 (N_8804,N_7181,N_7277);
and U8805 (N_8805,N_7996,N_7344);
or U8806 (N_8806,N_7270,N_6443);
and U8807 (N_8807,N_6137,N_6019);
nand U8808 (N_8808,N_7045,N_7787);
and U8809 (N_8809,N_7837,N_6021);
and U8810 (N_8810,N_7327,N_6957);
or U8811 (N_8811,N_7500,N_6885);
nor U8812 (N_8812,N_6924,N_7279);
nor U8813 (N_8813,N_7182,N_7535);
and U8814 (N_8814,N_7304,N_7026);
nor U8815 (N_8815,N_7437,N_6954);
and U8816 (N_8816,N_7955,N_7365);
xor U8817 (N_8817,N_7491,N_6703);
nor U8818 (N_8818,N_7565,N_6915);
or U8819 (N_8819,N_7982,N_6204);
nand U8820 (N_8820,N_7145,N_6930);
or U8821 (N_8821,N_6227,N_6436);
and U8822 (N_8822,N_7723,N_6128);
nor U8823 (N_8823,N_6785,N_7238);
xnor U8824 (N_8824,N_6003,N_6802);
nand U8825 (N_8825,N_6520,N_6214);
and U8826 (N_8826,N_7265,N_7367);
or U8827 (N_8827,N_7452,N_7754);
nand U8828 (N_8828,N_6901,N_7431);
nand U8829 (N_8829,N_7139,N_7097);
nor U8830 (N_8830,N_7690,N_7525);
and U8831 (N_8831,N_7957,N_7273);
nand U8832 (N_8832,N_7031,N_7135);
or U8833 (N_8833,N_7287,N_6777);
nand U8834 (N_8834,N_6858,N_7796);
or U8835 (N_8835,N_7313,N_6503);
nand U8836 (N_8836,N_6501,N_6619);
and U8837 (N_8837,N_7920,N_6261);
nor U8838 (N_8838,N_7379,N_6595);
and U8839 (N_8839,N_6369,N_7962);
nand U8840 (N_8840,N_7830,N_7187);
xor U8841 (N_8841,N_7132,N_6756);
nand U8842 (N_8842,N_7768,N_6435);
nor U8843 (N_8843,N_6063,N_7484);
nand U8844 (N_8844,N_6236,N_7082);
and U8845 (N_8845,N_6511,N_6763);
and U8846 (N_8846,N_7776,N_7969);
nor U8847 (N_8847,N_7345,N_7971);
and U8848 (N_8848,N_6948,N_7453);
nor U8849 (N_8849,N_7302,N_7355);
or U8850 (N_8850,N_6590,N_7590);
and U8851 (N_8851,N_7479,N_7017);
nand U8852 (N_8852,N_6791,N_6418);
xor U8853 (N_8853,N_6762,N_7940);
or U8854 (N_8854,N_7298,N_6678);
xor U8855 (N_8855,N_6238,N_7284);
nor U8856 (N_8856,N_7586,N_6652);
or U8857 (N_8857,N_6965,N_7910);
nor U8858 (N_8858,N_7697,N_6647);
and U8859 (N_8859,N_7393,N_7366);
and U8860 (N_8860,N_7426,N_7303);
or U8861 (N_8861,N_7325,N_7505);
xnor U8862 (N_8862,N_7950,N_7455);
or U8863 (N_8863,N_7760,N_6094);
xnor U8864 (N_8864,N_7886,N_7894);
nor U8865 (N_8865,N_6377,N_7845);
nand U8866 (N_8866,N_7836,N_6744);
or U8867 (N_8867,N_7062,N_7869);
and U8868 (N_8868,N_7307,N_6241);
nand U8869 (N_8869,N_7548,N_6982);
and U8870 (N_8870,N_7459,N_6812);
or U8871 (N_8871,N_6830,N_7881);
nor U8872 (N_8872,N_6102,N_6630);
nand U8873 (N_8873,N_6847,N_6471);
nor U8874 (N_8874,N_6767,N_7706);
or U8875 (N_8875,N_7852,N_6692);
nand U8876 (N_8876,N_7309,N_6075);
nor U8877 (N_8877,N_7137,N_6978);
nand U8878 (N_8878,N_7118,N_6547);
and U8879 (N_8879,N_6974,N_7251);
nor U8880 (N_8880,N_7191,N_6940);
nand U8881 (N_8881,N_6461,N_6531);
xnor U8882 (N_8882,N_7623,N_6891);
nand U8883 (N_8883,N_7645,N_7486);
or U8884 (N_8884,N_6287,N_6492);
or U8885 (N_8885,N_6706,N_7547);
nor U8886 (N_8886,N_6579,N_7405);
nand U8887 (N_8887,N_7909,N_7198);
nor U8888 (N_8888,N_7873,N_7041);
or U8889 (N_8889,N_7248,N_7207);
nand U8890 (N_8890,N_7221,N_6746);
or U8891 (N_8891,N_7704,N_7860);
and U8892 (N_8892,N_7384,N_7780);
xor U8893 (N_8893,N_6803,N_7380);
or U8894 (N_8894,N_6011,N_7291);
nand U8895 (N_8895,N_6759,N_6621);
nand U8896 (N_8896,N_7550,N_7456);
and U8897 (N_8897,N_6758,N_7377);
xor U8898 (N_8898,N_7388,N_7144);
nor U8899 (N_8899,N_7682,N_7745);
nor U8900 (N_8900,N_7742,N_7746);
xor U8901 (N_8901,N_7513,N_7199);
nor U8902 (N_8902,N_7556,N_6807);
and U8903 (N_8903,N_6871,N_6196);
nor U8904 (N_8904,N_7211,N_6987);
and U8905 (N_8905,N_7002,N_6943);
or U8906 (N_8906,N_6770,N_7230);
xnor U8907 (N_8907,N_6883,N_6465);
nor U8908 (N_8908,N_7811,N_6423);
and U8909 (N_8909,N_6298,N_7285);
nor U8910 (N_8910,N_7386,N_7498);
and U8911 (N_8911,N_6911,N_6860);
nor U8912 (N_8912,N_6725,N_7802);
xnor U8913 (N_8913,N_6437,N_7009);
nor U8914 (N_8914,N_7280,N_7613);
and U8915 (N_8915,N_6658,N_7580);
xor U8916 (N_8916,N_7778,N_6000);
nor U8917 (N_8917,N_6121,N_6156);
nor U8918 (N_8918,N_7914,N_6787);
nor U8919 (N_8919,N_7140,N_6502);
xor U8920 (N_8920,N_7803,N_7987);
and U8921 (N_8921,N_7142,N_6343);
nand U8922 (N_8922,N_7069,N_6782);
or U8923 (N_8923,N_7180,N_6623);
and U8924 (N_8924,N_6960,N_7829);
and U8925 (N_8925,N_6642,N_6645);
or U8926 (N_8926,N_7092,N_6189);
nand U8927 (N_8927,N_6716,N_7487);
xnor U8928 (N_8928,N_6257,N_7838);
or U8929 (N_8929,N_7035,N_6462);
or U8930 (N_8930,N_6816,N_7083);
nand U8931 (N_8931,N_6748,N_6923);
and U8932 (N_8932,N_7402,N_6722);
nor U8933 (N_8933,N_7801,N_7171);
xor U8934 (N_8934,N_6508,N_6062);
or U8935 (N_8935,N_6904,N_6873);
nand U8936 (N_8936,N_7278,N_7877);
or U8937 (N_8937,N_6671,N_7839);
nand U8938 (N_8938,N_7821,N_6284);
xor U8939 (N_8939,N_6814,N_7272);
xor U8940 (N_8940,N_6305,N_6555);
or U8941 (N_8941,N_6469,N_7454);
nor U8942 (N_8942,N_7420,N_7945);
or U8943 (N_8943,N_6230,N_7485);
xor U8944 (N_8944,N_6010,N_6174);
nor U8945 (N_8945,N_7815,N_7005);
nand U8946 (N_8946,N_6197,N_7038);
nand U8947 (N_8947,N_7053,N_6056);
xnor U8948 (N_8948,N_6504,N_6293);
nor U8949 (N_8949,N_7991,N_7036);
or U8950 (N_8950,N_6300,N_6899);
nor U8951 (N_8951,N_7403,N_7173);
nand U8952 (N_8952,N_7779,N_7161);
or U8953 (N_8953,N_6425,N_6226);
and U8954 (N_8954,N_7516,N_6410);
nand U8955 (N_8955,N_6276,N_7922);
or U8956 (N_8956,N_7160,N_7905);
or U8957 (N_8957,N_7995,N_7842);
xnor U8958 (N_8958,N_7933,N_6685);
and U8959 (N_8959,N_6815,N_6892);
or U8960 (N_8960,N_6160,N_7290);
nor U8961 (N_8961,N_7560,N_6417);
xnor U8962 (N_8962,N_7989,N_7372);
xnor U8963 (N_8963,N_7711,N_7185);
nor U8964 (N_8964,N_6811,N_6379);
xnor U8965 (N_8965,N_6886,N_7880);
or U8966 (N_8966,N_6981,N_6670);
xnor U8967 (N_8967,N_7846,N_7652);
nand U8968 (N_8968,N_7589,N_6388);
nand U8969 (N_8969,N_7003,N_6233);
or U8970 (N_8970,N_7739,N_7322);
and U8971 (N_8971,N_7030,N_6921);
nand U8972 (N_8972,N_7553,N_6691);
or U8973 (N_8973,N_6893,N_6564);
nor U8974 (N_8974,N_6747,N_6674);
xnor U8975 (N_8975,N_7972,N_7958);
or U8976 (N_8976,N_6654,N_6406);
or U8977 (N_8977,N_7970,N_6403);
or U8978 (N_8978,N_6668,N_6399);
nor U8979 (N_8979,N_7358,N_7899);
nand U8980 (N_8980,N_6702,N_7352);
nor U8981 (N_8981,N_6158,N_6256);
and U8982 (N_8982,N_7916,N_7089);
and U8983 (N_8983,N_6254,N_6760);
xor U8984 (N_8984,N_7572,N_7481);
or U8985 (N_8985,N_7507,N_6239);
nand U8986 (N_8986,N_6040,N_6096);
or U8987 (N_8987,N_6351,N_7468);
nor U8988 (N_8988,N_7630,N_7119);
nand U8989 (N_8989,N_6422,N_7496);
and U8990 (N_8990,N_6996,N_7095);
xor U8991 (N_8991,N_6072,N_6218);
nand U8992 (N_8992,N_7443,N_7540);
nand U8993 (N_8993,N_7079,N_6111);
nor U8994 (N_8994,N_6302,N_7361);
nand U8995 (N_8995,N_6009,N_6698);
and U8996 (N_8996,N_7686,N_6552);
nor U8997 (N_8997,N_7329,N_6839);
xnor U8998 (N_8998,N_7044,N_7037);
and U8999 (N_8999,N_7805,N_6213);
nor U9000 (N_9000,N_7854,N_7247);
nand U9001 (N_9001,N_6915,N_6361);
xor U9002 (N_9002,N_7620,N_7775);
or U9003 (N_9003,N_6429,N_7072);
xor U9004 (N_9004,N_7760,N_6411);
or U9005 (N_9005,N_7004,N_6041);
or U9006 (N_9006,N_7987,N_7933);
xnor U9007 (N_9007,N_6549,N_7181);
or U9008 (N_9008,N_7839,N_7014);
nand U9009 (N_9009,N_7871,N_7330);
and U9010 (N_9010,N_6578,N_7733);
nand U9011 (N_9011,N_7111,N_6915);
nand U9012 (N_9012,N_7583,N_6411);
nor U9013 (N_9013,N_6012,N_6528);
and U9014 (N_9014,N_7927,N_7307);
nand U9015 (N_9015,N_6122,N_6532);
xor U9016 (N_9016,N_7485,N_6265);
nor U9017 (N_9017,N_6540,N_7595);
xor U9018 (N_9018,N_7697,N_6099);
nand U9019 (N_9019,N_7888,N_7696);
or U9020 (N_9020,N_6138,N_6227);
or U9021 (N_9021,N_7137,N_7825);
xor U9022 (N_9022,N_6084,N_7700);
and U9023 (N_9023,N_6559,N_7179);
xnor U9024 (N_9024,N_7684,N_6951);
nand U9025 (N_9025,N_6027,N_7441);
xnor U9026 (N_9026,N_6969,N_7683);
nand U9027 (N_9027,N_7941,N_7313);
or U9028 (N_9028,N_6300,N_6099);
nand U9029 (N_9029,N_6749,N_7821);
or U9030 (N_9030,N_7747,N_6938);
nand U9031 (N_9031,N_6121,N_6854);
xnor U9032 (N_9032,N_7358,N_7529);
nand U9033 (N_9033,N_6424,N_6307);
and U9034 (N_9034,N_7700,N_7029);
xor U9035 (N_9035,N_7308,N_6769);
nor U9036 (N_9036,N_7344,N_7830);
nand U9037 (N_9037,N_6598,N_7826);
xnor U9038 (N_9038,N_7340,N_6576);
and U9039 (N_9039,N_7883,N_6939);
nand U9040 (N_9040,N_7181,N_6355);
nor U9041 (N_9041,N_7495,N_7809);
nor U9042 (N_9042,N_6399,N_7886);
nand U9043 (N_9043,N_6649,N_6045);
nand U9044 (N_9044,N_6283,N_7148);
nor U9045 (N_9045,N_7077,N_6689);
nand U9046 (N_9046,N_6802,N_6614);
or U9047 (N_9047,N_6003,N_6670);
xor U9048 (N_9048,N_7207,N_7265);
and U9049 (N_9049,N_7772,N_6322);
or U9050 (N_9050,N_7771,N_7891);
and U9051 (N_9051,N_6174,N_6882);
xor U9052 (N_9052,N_7789,N_7452);
and U9053 (N_9053,N_6276,N_6873);
nand U9054 (N_9054,N_7237,N_7080);
xnor U9055 (N_9055,N_6386,N_6858);
nor U9056 (N_9056,N_6065,N_6600);
nand U9057 (N_9057,N_6367,N_6085);
xnor U9058 (N_9058,N_6549,N_6545);
nand U9059 (N_9059,N_7026,N_7600);
nand U9060 (N_9060,N_7992,N_7875);
xnor U9061 (N_9061,N_7206,N_6246);
xor U9062 (N_9062,N_6324,N_7963);
or U9063 (N_9063,N_6130,N_7908);
nor U9064 (N_9064,N_7407,N_6607);
or U9065 (N_9065,N_7563,N_7884);
xnor U9066 (N_9066,N_7431,N_7985);
nand U9067 (N_9067,N_6803,N_6143);
or U9068 (N_9068,N_7275,N_6618);
and U9069 (N_9069,N_7913,N_6928);
nor U9070 (N_9070,N_6218,N_7026);
nand U9071 (N_9071,N_7890,N_6550);
nand U9072 (N_9072,N_7291,N_7420);
and U9073 (N_9073,N_7327,N_7534);
or U9074 (N_9074,N_7769,N_6341);
nand U9075 (N_9075,N_7762,N_6130);
and U9076 (N_9076,N_7049,N_6231);
nor U9077 (N_9077,N_7152,N_6709);
nor U9078 (N_9078,N_7519,N_7031);
nand U9079 (N_9079,N_6661,N_7430);
xor U9080 (N_9080,N_6245,N_6860);
or U9081 (N_9081,N_7729,N_6734);
and U9082 (N_9082,N_7064,N_6919);
nor U9083 (N_9083,N_7070,N_7695);
xor U9084 (N_9084,N_6326,N_7207);
nor U9085 (N_9085,N_7273,N_6982);
and U9086 (N_9086,N_7527,N_6998);
xnor U9087 (N_9087,N_7374,N_7545);
nand U9088 (N_9088,N_7625,N_6499);
or U9089 (N_9089,N_7884,N_6336);
nor U9090 (N_9090,N_7270,N_7931);
xor U9091 (N_9091,N_6447,N_6718);
or U9092 (N_9092,N_6654,N_7937);
nor U9093 (N_9093,N_7543,N_6208);
xor U9094 (N_9094,N_6271,N_6428);
nand U9095 (N_9095,N_6448,N_6972);
nor U9096 (N_9096,N_6831,N_7578);
nand U9097 (N_9097,N_6497,N_6076);
nor U9098 (N_9098,N_6748,N_7708);
nand U9099 (N_9099,N_7972,N_7279);
nor U9100 (N_9100,N_6962,N_7923);
xnor U9101 (N_9101,N_6834,N_6981);
nand U9102 (N_9102,N_6089,N_7583);
nand U9103 (N_9103,N_6016,N_6556);
or U9104 (N_9104,N_6807,N_7316);
and U9105 (N_9105,N_7676,N_7806);
or U9106 (N_9106,N_7965,N_7250);
or U9107 (N_9107,N_7505,N_7101);
or U9108 (N_9108,N_7939,N_6896);
and U9109 (N_9109,N_6745,N_6999);
or U9110 (N_9110,N_7615,N_7944);
and U9111 (N_9111,N_7832,N_7011);
and U9112 (N_9112,N_6251,N_6146);
or U9113 (N_9113,N_7564,N_7236);
xor U9114 (N_9114,N_7134,N_7357);
and U9115 (N_9115,N_6134,N_6227);
or U9116 (N_9116,N_7479,N_7127);
nor U9117 (N_9117,N_6724,N_7575);
xor U9118 (N_9118,N_6506,N_7917);
and U9119 (N_9119,N_7455,N_6027);
nand U9120 (N_9120,N_7239,N_7719);
or U9121 (N_9121,N_7036,N_6147);
nor U9122 (N_9122,N_7516,N_6714);
nand U9123 (N_9123,N_6451,N_7904);
and U9124 (N_9124,N_6655,N_6130);
nand U9125 (N_9125,N_6750,N_6071);
nor U9126 (N_9126,N_7657,N_7769);
nand U9127 (N_9127,N_7729,N_7585);
nand U9128 (N_9128,N_7172,N_7453);
nand U9129 (N_9129,N_6747,N_6863);
nor U9130 (N_9130,N_6795,N_6861);
and U9131 (N_9131,N_7023,N_6339);
nand U9132 (N_9132,N_6771,N_7807);
nor U9133 (N_9133,N_6772,N_7121);
xor U9134 (N_9134,N_6500,N_7496);
xnor U9135 (N_9135,N_6498,N_7621);
xor U9136 (N_9136,N_6628,N_6763);
and U9137 (N_9137,N_7235,N_6111);
nand U9138 (N_9138,N_7578,N_7130);
nand U9139 (N_9139,N_6299,N_7107);
or U9140 (N_9140,N_6556,N_7457);
and U9141 (N_9141,N_7906,N_6329);
xnor U9142 (N_9142,N_6966,N_6663);
and U9143 (N_9143,N_7943,N_7218);
or U9144 (N_9144,N_7796,N_6279);
nand U9145 (N_9145,N_7258,N_7953);
nor U9146 (N_9146,N_7655,N_7303);
xor U9147 (N_9147,N_7719,N_7963);
or U9148 (N_9148,N_6623,N_6911);
nand U9149 (N_9149,N_7112,N_6407);
xor U9150 (N_9150,N_7415,N_7729);
nand U9151 (N_9151,N_7116,N_7785);
xnor U9152 (N_9152,N_7860,N_7703);
nor U9153 (N_9153,N_7966,N_6986);
nor U9154 (N_9154,N_6615,N_6739);
xor U9155 (N_9155,N_7006,N_6681);
nand U9156 (N_9156,N_7635,N_6067);
nand U9157 (N_9157,N_6608,N_7353);
nor U9158 (N_9158,N_7773,N_6534);
and U9159 (N_9159,N_6770,N_6372);
nand U9160 (N_9160,N_7698,N_6022);
or U9161 (N_9161,N_6977,N_7092);
nand U9162 (N_9162,N_6349,N_6994);
xnor U9163 (N_9163,N_7935,N_7403);
nor U9164 (N_9164,N_6392,N_6400);
nor U9165 (N_9165,N_6179,N_6715);
or U9166 (N_9166,N_6200,N_6149);
or U9167 (N_9167,N_6247,N_7296);
and U9168 (N_9168,N_6313,N_6083);
or U9169 (N_9169,N_6399,N_6894);
nor U9170 (N_9170,N_7513,N_6832);
xor U9171 (N_9171,N_7442,N_6480);
nand U9172 (N_9172,N_7232,N_6974);
nor U9173 (N_9173,N_6073,N_6992);
nor U9174 (N_9174,N_7750,N_6477);
nand U9175 (N_9175,N_6422,N_7190);
xor U9176 (N_9176,N_6471,N_7188);
nand U9177 (N_9177,N_6272,N_7284);
xor U9178 (N_9178,N_7838,N_6958);
xor U9179 (N_9179,N_6599,N_6105);
or U9180 (N_9180,N_6645,N_7203);
nand U9181 (N_9181,N_7588,N_6360);
and U9182 (N_9182,N_6342,N_6217);
xnor U9183 (N_9183,N_6594,N_6221);
nor U9184 (N_9184,N_7867,N_7061);
and U9185 (N_9185,N_7712,N_7410);
nor U9186 (N_9186,N_6078,N_6392);
or U9187 (N_9187,N_6133,N_7649);
nor U9188 (N_9188,N_6455,N_7701);
or U9189 (N_9189,N_7866,N_7668);
or U9190 (N_9190,N_6422,N_7493);
and U9191 (N_9191,N_7372,N_7029);
xor U9192 (N_9192,N_6797,N_6683);
nand U9193 (N_9193,N_6443,N_7606);
nand U9194 (N_9194,N_7348,N_7206);
nor U9195 (N_9195,N_7659,N_6588);
nor U9196 (N_9196,N_7657,N_6237);
nand U9197 (N_9197,N_7215,N_6493);
or U9198 (N_9198,N_7068,N_7295);
and U9199 (N_9199,N_7934,N_7090);
or U9200 (N_9200,N_6509,N_6650);
and U9201 (N_9201,N_7092,N_7327);
nand U9202 (N_9202,N_6727,N_6327);
nand U9203 (N_9203,N_7607,N_6474);
nand U9204 (N_9204,N_6459,N_6177);
nor U9205 (N_9205,N_6249,N_7534);
xor U9206 (N_9206,N_7490,N_7386);
nand U9207 (N_9207,N_7454,N_6369);
and U9208 (N_9208,N_6416,N_7500);
or U9209 (N_9209,N_6345,N_6999);
or U9210 (N_9210,N_7115,N_7498);
or U9211 (N_9211,N_6760,N_7811);
nor U9212 (N_9212,N_6085,N_6712);
and U9213 (N_9213,N_7352,N_6835);
and U9214 (N_9214,N_6792,N_7920);
nand U9215 (N_9215,N_6421,N_6920);
nor U9216 (N_9216,N_7026,N_7741);
xor U9217 (N_9217,N_6799,N_7829);
nor U9218 (N_9218,N_7645,N_7147);
nor U9219 (N_9219,N_7525,N_7716);
and U9220 (N_9220,N_6672,N_7051);
nor U9221 (N_9221,N_6065,N_6603);
nor U9222 (N_9222,N_7103,N_7843);
xor U9223 (N_9223,N_6289,N_6916);
and U9224 (N_9224,N_6375,N_6505);
and U9225 (N_9225,N_7555,N_7282);
or U9226 (N_9226,N_7846,N_6339);
nand U9227 (N_9227,N_7231,N_7034);
nand U9228 (N_9228,N_6270,N_6910);
nor U9229 (N_9229,N_6259,N_6928);
nand U9230 (N_9230,N_7963,N_6468);
nand U9231 (N_9231,N_6875,N_7535);
and U9232 (N_9232,N_7721,N_7948);
nor U9233 (N_9233,N_6227,N_6770);
nor U9234 (N_9234,N_7246,N_7913);
nand U9235 (N_9235,N_7369,N_6662);
and U9236 (N_9236,N_7069,N_6083);
nand U9237 (N_9237,N_6227,N_7718);
xor U9238 (N_9238,N_6968,N_6550);
nor U9239 (N_9239,N_7439,N_6198);
and U9240 (N_9240,N_6312,N_6066);
xnor U9241 (N_9241,N_7105,N_7018);
and U9242 (N_9242,N_6531,N_6208);
nand U9243 (N_9243,N_7409,N_6606);
nand U9244 (N_9244,N_6699,N_6792);
and U9245 (N_9245,N_6185,N_6991);
or U9246 (N_9246,N_6072,N_6247);
nor U9247 (N_9247,N_6197,N_7106);
nor U9248 (N_9248,N_7224,N_7676);
nor U9249 (N_9249,N_7193,N_6799);
nand U9250 (N_9250,N_6616,N_6072);
or U9251 (N_9251,N_7774,N_7005);
xnor U9252 (N_9252,N_6380,N_6126);
or U9253 (N_9253,N_7189,N_7584);
nand U9254 (N_9254,N_6790,N_7449);
nor U9255 (N_9255,N_7542,N_7751);
or U9256 (N_9256,N_6065,N_6123);
xnor U9257 (N_9257,N_6550,N_7160);
nor U9258 (N_9258,N_6814,N_6312);
or U9259 (N_9259,N_6067,N_7772);
nor U9260 (N_9260,N_6671,N_7181);
nand U9261 (N_9261,N_6384,N_7923);
nand U9262 (N_9262,N_7568,N_7334);
xor U9263 (N_9263,N_7539,N_6218);
xor U9264 (N_9264,N_6564,N_6273);
and U9265 (N_9265,N_6388,N_7273);
and U9266 (N_9266,N_7145,N_6837);
nand U9267 (N_9267,N_6164,N_6623);
or U9268 (N_9268,N_7550,N_6656);
xnor U9269 (N_9269,N_7242,N_7076);
nor U9270 (N_9270,N_7318,N_7912);
nand U9271 (N_9271,N_6198,N_6727);
nor U9272 (N_9272,N_6494,N_6236);
xor U9273 (N_9273,N_6940,N_7613);
nand U9274 (N_9274,N_6655,N_7545);
and U9275 (N_9275,N_6677,N_7225);
and U9276 (N_9276,N_7917,N_6180);
and U9277 (N_9277,N_6573,N_6281);
nor U9278 (N_9278,N_6251,N_7813);
nor U9279 (N_9279,N_6066,N_7548);
and U9280 (N_9280,N_7364,N_6097);
and U9281 (N_9281,N_6524,N_6449);
nand U9282 (N_9282,N_7761,N_7946);
xnor U9283 (N_9283,N_6921,N_7958);
or U9284 (N_9284,N_6959,N_7244);
nor U9285 (N_9285,N_6680,N_7882);
xnor U9286 (N_9286,N_6092,N_6983);
nor U9287 (N_9287,N_7184,N_7985);
and U9288 (N_9288,N_7973,N_7179);
nand U9289 (N_9289,N_7619,N_7569);
and U9290 (N_9290,N_6906,N_6201);
and U9291 (N_9291,N_6912,N_6487);
or U9292 (N_9292,N_7334,N_6416);
nor U9293 (N_9293,N_7375,N_6669);
nor U9294 (N_9294,N_7769,N_6167);
and U9295 (N_9295,N_6565,N_6739);
nor U9296 (N_9296,N_6579,N_7926);
nand U9297 (N_9297,N_7861,N_7131);
xnor U9298 (N_9298,N_7212,N_6472);
or U9299 (N_9299,N_7518,N_7170);
xor U9300 (N_9300,N_6330,N_6849);
and U9301 (N_9301,N_6838,N_6985);
xnor U9302 (N_9302,N_6457,N_6727);
or U9303 (N_9303,N_7045,N_6831);
nand U9304 (N_9304,N_6727,N_6368);
xnor U9305 (N_9305,N_6421,N_6707);
xor U9306 (N_9306,N_7859,N_6684);
nor U9307 (N_9307,N_6667,N_7206);
nand U9308 (N_9308,N_7194,N_6586);
nor U9309 (N_9309,N_7316,N_6249);
nor U9310 (N_9310,N_6476,N_6372);
nand U9311 (N_9311,N_7476,N_6736);
nor U9312 (N_9312,N_6114,N_6444);
nand U9313 (N_9313,N_7217,N_7382);
and U9314 (N_9314,N_7116,N_6095);
nor U9315 (N_9315,N_7027,N_7562);
and U9316 (N_9316,N_7497,N_7801);
xor U9317 (N_9317,N_7648,N_6711);
nor U9318 (N_9318,N_6958,N_7212);
xor U9319 (N_9319,N_6081,N_7155);
and U9320 (N_9320,N_6549,N_7146);
nand U9321 (N_9321,N_6676,N_7733);
nor U9322 (N_9322,N_7711,N_6273);
or U9323 (N_9323,N_6417,N_6120);
and U9324 (N_9324,N_6687,N_7090);
nand U9325 (N_9325,N_7310,N_7198);
nand U9326 (N_9326,N_7628,N_7911);
or U9327 (N_9327,N_6829,N_6399);
nor U9328 (N_9328,N_7936,N_7882);
nand U9329 (N_9329,N_6395,N_7693);
xor U9330 (N_9330,N_7200,N_7587);
nand U9331 (N_9331,N_6389,N_6916);
nor U9332 (N_9332,N_6352,N_7716);
or U9333 (N_9333,N_7842,N_6874);
and U9334 (N_9334,N_7763,N_6417);
nor U9335 (N_9335,N_6296,N_6443);
xor U9336 (N_9336,N_7119,N_6958);
nor U9337 (N_9337,N_7549,N_6214);
xor U9338 (N_9338,N_6538,N_6541);
and U9339 (N_9339,N_6527,N_6929);
xor U9340 (N_9340,N_6475,N_7318);
nand U9341 (N_9341,N_7959,N_7997);
or U9342 (N_9342,N_6984,N_7094);
nand U9343 (N_9343,N_6516,N_7710);
or U9344 (N_9344,N_7319,N_6756);
or U9345 (N_9345,N_7218,N_6018);
nand U9346 (N_9346,N_6693,N_7719);
nand U9347 (N_9347,N_7179,N_7050);
or U9348 (N_9348,N_6886,N_7757);
or U9349 (N_9349,N_6277,N_6994);
nor U9350 (N_9350,N_6751,N_6491);
xnor U9351 (N_9351,N_6870,N_7444);
or U9352 (N_9352,N_6503,N_7080);
and U9353 (N_9353,N_7273,N_6672);
or U9354 (N_9354,N_7461,N_6222);
nor U9355 (N_9355,N_6508,N_7164);
and U9356 (N_9356,N_7501,N_6114);
nand U9357 (N_9357,N_7826,N_6203);
xnor U9358 (N_9358,N_7245,N_6134);
nand U9359 (N_9359,N_6747,N_7796);
and U9360 (N_9360,N_6033,N_6456);
nor U9361 (N_9361,N_6807,N_7707);
or U9362 (N_9362,N_6582,N_7497);
and U9363 (N_9363,N_6471,N_6616);
nor U9364 (N_9364,N_6905,N_7248);
nor U9365 (N_9365,N_7170,N_7792);
nand U9366 (N_9366,N_7774,N_7313);
or U9367 (N_9367,N_6759,N_7509);
and U9368 (N_9368,N_6309,N_6167);
nand U9369 (N_9369,N_6191,N_6849);
nor U9370 (N_9370,N_7160,N_7663);
nor U9371 (N_9371,N_6272,N_7155);
nor U9372 (N_9372,N_6538,N_6350);
nand U9373 (N_9373,N_7743,N_7219);
nor U9374 (N_9374,N_6653,N_7410);
or U9375 (N_9375,N_6541,N_6588);
nor U9376 (N_9376,N_7073,N_7605);
or U9377 (N_9377,N_7003,N_7353);
nand U9378 (N_9378,N_7749,N_6693);
nand U9379 (N_9379,N_7739,N_7689);
or U9380 (N_9380,N_6006,N_7679);
or U9381 (N_9381,N_7665,N_7727);
xnor U9382 (N_9382,N_6490,N_6914);
nor U9383 (N_9383,N_7320,N_7078);
and U9384 (N_9384,N_7092,N_6621);
nand U9385 (N_9385,N_7173,N_7960);
nor U9386 (N_9386,N_7660,N_7693);
nand U9387 (N_9387,N_6650,N_7503);
or U9388 (N_9388,N_6754,N_6827);
xnor U9389 (N_9389,N_6545,N_6869);
nor U9390 (N_9390,N_6558,N_7390);
nor U9391 (N_9391,N_6110,N_7043);
nor U9392 (N_9392,N_6270,N_7833);
nor U9393 (N_9393,N_6273,N_7887);
nor U9394 (N_9394,N_6433,N_6441);
nor U9395 (N_9395,N_6750,N_6373);
xor U9396 (N_9396,N_7421,N_7191);
or U9397 (N_9397,N_6067,N_6127);
and U9398 (N_9398,N_7410,N_6400);
xnor U9399 (N_9399,N_6462,N_7419);
or U9400 (N_9400,N_6897,N_7180);
xnor U9401 (N_9401,N_7284,N_6174);
or U9402 (N_9402,N_6018,N_6793);
and U9403 (N_9403,N_6817,N_7700);
xor U9404 (N_9404,N_7797,N_7120);
and U9405 (N_9405,N_7727,N_6445);
and U9406 (N_9406,N_6024,N_7464);
and U9407 (N_9407,N_6750,N_7124);
nor U9408 (N_9408,N_6363,N_6132);
nand U9409 (N_9409,N_6116,N_7080);
or U9410 (N_9410,N_6682,N_6604);
and U9411 (N_9411,N_6440,N_7070);
nand U9412 (N_9412,N_7568,N_7160);
xnor U9413 (N_9413,N_7599,N_6569);
nor U9414 (N_9414,N_6175,N_7847);
nor U9415 (N_9415,N_6074,N_6514);
and U9416 (N_9416,N_6543,N_7045);
and U9417 (N_9417,N_7969,N_7810);
xor U9418 (N_9418,N_7348,N_6691);
and U9419 (N_9419,N_6695,N_7063);
and U9420 (N_9420,N_6551,N_6157);
and U9421 (N_9421,N_6268,N_6691);
nor U9422 (N_9422,N_7930,N_7436);
or U9423 (N_9423,N_7760,N_6659);
nor U9424 (N_9424,N_6218,N_7456);
nand U9425 (N_9425,N_6980,N_7746);
nand U9426 (N_9426,N_6583,N_7020);
nor U9427 (N_9427,N_6867,N_6597);
xnor U9428 (N_9428,N_7092,N_7209);
nand U9429 (N_9429,N_7686,N_7890);
xor U9430 (N_9430,N_6787,N_6369);
or U9431 (N_9431,N_6200,N_6317);
xnor U9432 (N_9432,N_6407,N_7653);
nand U9433 (N_9433,N_6226,N_6782);
nor U9434 (N_9434,N_6980,N_7386);
and U9435 (N_9435,N_6890,N_7316);
and U9436 (N_9436,N_7338,N_6052);
or U9437 (N_9437,N_7299,N_6551);
xnor U9438 (N_9438,N_6219,N_7463);
nor U9439 (N_9439,N_6260,N_7191);
xnor U9440 (N_9440,N_6497,N_6905);
and U9441 (N_9441,N_6079,N_6491);
nand U9442 (N_9442,N_7515,N_6524);
xor U9443 (N_9443,N_6056,N_6423);
nor U9444 (N_9444,N_6901,N_7364);
nor U9445 (N_9445,N_7603,N_6304);
and U9446 (N_9446,N_7138,N_6864);
and U9447 (N_9447,N_7218,N_6237);
nor U9448 (N_9448,N_6461,N_7218);
or U9449 (N_9449,N_6814,N_6402);
xor U9450 (N_9450,N_6511,N_6200);
nand U9451 (N_9451,N_6843,N_6937);
xnor U9452 (N_9452,N_7821,N_7007);
nand U9453 (N_9453,N_7681,N_7228);
or U9454 (N_9454,N_6579,N_6265);
nor U9455 (N_9455,N_7265,N_6327);
and U9456 (N_9456,N_6949,N_7820);
and U9457 (N_9457,N_7592,N_7341);
nor U9458 (N_9458,N_6908,N_7395);
nor U9459 (N_9459,N_6826,N_6310);
and U9460 (N_9460,N_7616,N_7881);
and U9461 (N_9461,N_7572,N_7778);
nor U9462 (N_9462,N_6505,N_7795);
xor U9463 (N_9463,N_6018,N_7894);
and U9464 (N_9464,N_7025,N_6915);
and U9465 (N_9465,N_7698,N_7908);
and U9466 (N_9466,N_7063,N_7488);
and U9467 (N_9467,N_7083,N_7271);
nand U9468 (N_9468,N_7576,N_7366);
nor U9469 (N_9469,N_7042,N_7018);
or U9470 (N_9470,N_6626,N_7086);
and U9471 (N_9471,N_6000,N_6361);
xnor U9472 (N_9472,N_7006,N_7385);
and U9473 (N_9473,N_7566,N_7178);
nor U9474 (N_9474,N_6764,N_7043);
nand U9475 (N_9475,N_7444,N_6693);
xor U9476 (N_9476,N_7512,N_7370);
and U9477 (N_9477,N_7023,N_6928);
nand U9478 (N_9478,N_7978,N_7370);
nor U9479 (N_9479,N_6461,N_6958);
or U9480 (N_9480,N_7139,N_6480);
nand U9481 (N_9481,N_7018,N_6335);
nand U9482 (N_9482,N_6137,N_7822);
nor U9483 (N_9483,N_6724,N_7258);
nand U9484 (N_9484,N_7310,N_6121);
or U9485 (N_9485,N_7363,N_6544);
nor U9486 (N_9486,N_7305,N_6401);
nor U9487 (N_9487,N_7823,N_7011);
xnor U9488 (N_9488,N_6772,N_7659);
or U9489 (N_9489,N_7724,N_6242);
nand U9490 (N_9490,N_6182,N_7791);
nand U9491 (N_9491,N_7669,N_7710);
nand U9492 (N_9492,N_7456,N_6076);
nor U9493 (N_9493,N_6636,N_7694);
nand U9494 (N_9494,N_6648,N_6873);
nor U9495 (N_9495,N_6824,N_7291);
xnor U9496 (N_9496,N_7204,N_6835);
and U9497 (N_9497,N_6531,N_6436);
or U9498 (N_9498,N_6448,N_6400);
and U9499 (N_9499,N_7354,N_6404);
xnor U9500 (N_9500,N_6499,N_7838);
and U9501 (N_9501,N_7415,N_7076);
or U9502 (N_9502,N_7213,N_7705);
nand U9503 (N_9503,N_7862,N_6835);
or U9504 (N_9504,N_7031,N_7526);
xnor U9505 (N_9505,N_7286,N_7063);
and U9506 (N_9506,N_6001,N_6218);
and U9507 (N_9507,N_6408,N_6600);
and U9508 (N_9508,N_7390,N_6944);
nor U9509 (N_9509,N_7938,N_7570);
xnor U9510 (N_9510,N_6241,N_6365);
nor U9511 (N_9511,N_7779,N_6806);
or U9512 (N_9512,N_7330,N_7066);
or U9513 (N_9513,N_7305,N_7553);
and U9514 (N_9514,N_7249,N_7898);
or U9515 (N_9515,N_6446,N_7223);
xnor U9516 (N_9516,N_7736,N_6871);
xnor U9517 (N_9517,N_6367,N_7859);
and U9518 (N_9518,N_6943,N_6859);
nand U9519 (N_9519,N_6582,N_7217);
nand U9520 (N_9520,N_6805,N_7057);
nor U9521 (N_9521,N_7959,N_7531);
or U9522 (N_9522,N_6800,N_7936);
or U9523 (N_9523,N_6874,N_7034);
xnor U9524 (N_9524,N_7788,N_7393);
and U9525 (N_9525,N_7203,N_6057);
or U9526 (N_9526,N_7771,N_6298);
or U9527 (N_9527,N_6860,N_7573);
and U9528 (N_9528,N_6462,N_6305);
and U9529 (N_9529,N_7320,N_7949);
or U9530 (N_9530,N_6331,N_7239);
nand U9531 (N_9531,N_7449,N_7675);
nor U9532 (N_9532,N_6205,N_6015);
and U9533 (N_9533,N_6763,N_7461);
nor U9534 (N_9534,N_7876,N_6506);
nand U9535 (N_9535,N_6220,N_7933);
nor U9536 (N_9536,N_6978,N_6009);
and U9537 (N_9537,N_7639,N_7963);
nand U9538 (N_9538,N_7894,N_6474);
or U9539 (N_9539,N_6261,N_7985);
xnor U9540 (N_9540,N_7970,N_7651);
or U9541 (N_9541,N_6732,N_6316);
xor U9542 (N_9542,N_7485,N_6613);
xnor U9543 (N_9543,N_7794,N_6680);
xor U9544 (N_9544,N_6632,N_7643);
xor U9545 (N_9545,N_6636,N_7735);
nor U9546 (N_9546,N_6358,N_6685);
or U9547 (N_9547,N_6554,N_6364);
nand U9548 (N_9548,N_7263,N_7934);
nand U9549 (N_9549,N_6783,N_6615);
and U9550 (N_9550,N_7517,N_7114);
nor U9551 (N_9551,N_7016,N_6197);
nand U9552 (N_9552,N_7107,N_6906);
nand U9553 (N_9553,N_7165,N_6422);
or U9554 (N_9554,N_7369,N_6688);
or U9555 (N_9555,N_6050,N_7020);
nor U9556 (N_9556,N_7335,N_7285);
or U9557 (N_9557,N_7773,N_7851);
nand U9558 (N_9558,N_7830,N_6011);
or U9559 (N_9559,N_7670,N_6029);
and U9560 (N_9560,N_7684,N_6663);
or U9561 (N_9561,N_7427,N_7284);
nand U9562 (N_9562,N_7968,N_6762);
nor U9563 (N_9563,N_7023,N_6564);
xnor U9564 (N_9564,N_6049,N_7738);
and U9565 (N_9565,N_6565,N_7007);
and U9566 (N_9566,N_6822,N_6751);
xnor U9567 (N_9567,N_7164,N_6169);
nor U9568 (N_9568,N_6493,N_6937);
xor U9569 (N_9569,N_6475,N_6405);
xnor U9570 (N_9570,N_6201,N_6580);
and U9571 (N_9571,N_6317,N_6502);
and U9572 (N_9572,N_7145,N_7709);
nand U9573 (N_9573,N_7376,N_7449);
and U9574 (N_9574,N_6726,N_7737);
nor U9575 (N_9575,N_6797,N_6259);
and U9576 (N_9576,N_7353,N_6640);
and U9577 (N_9577,N_6051,N_6878);
nor U9578 (N_9578,N_6459,N_7180);
or U9579 (N_9579,N_7594,N_7030);
nand U9580 (N_9580,N_6770,N_6159);
and U9581 (N_9581,N_7555,N_6271);
or U9582 (N_9582,N_7411,N_7104);
or U9583 (N_9583,N_6790,N_6798);
xor U9584 (N_9584,N_7026,N_6432);
nor U9585 (N_9585,N_7923,N_7666);
xnor U9586 (N_9586,N_7170,N_6556);
and U9587 (N_9587,N_6958,N_6781);
nor U9588 (N_9588,N_6382,N_6494);
xnor U9589 (N_9589,N_6135,N_6871);
nand U9590 (N_9590,N_7008,N_6702);
nor U9591 (N_9591,N_7605,N_6239);
xnor U9592 (N_9592,N_6730,N_6666);
and U9593 (N_9593,N_7881,N_6517);
nor U9594 (N_9594,N_6851,N_6592);
xnor U9595 (N_9595,N_7417,N_6261);
nand U9596 (N_9596,N_6780,N_7319);
nand U9597 (N_9597,N_6421,N_7116);
nor U9598 (N_9598,N_6309,N_6669);
nand U9599 (N_9599,N_7155,N_7028);
nand U9600 (N_9600,N_7150,N_7745);
xor U9601 (N_9601,N_6385,N_7255);
and U9602 (N_9602,N_7744,N_7989);
and U9603 (N_9603,N_7922,N_7157);
or U9604 (N_9604,N_7442,N_7244);
or U9605 (N_9605,N_6068,N_7596);
nand U9606 (N_9606,N_6625,N_6298);
xnor U9607 (N_9607,N_6290,N_7897);
or U9608 (N_9608,N_6901,N_7035);
nand U9609 (N_9609,N_7648,N_6097);
and U9610 (N_9610,N_6578,N_6587);
nand U9611 (N_9611,N_7382,N_6621);
or U9612 (N_9612,N_7920,N_6253);
and U9613 (N_9613,N_7769,N_6697);
or U9614 (N_9614,N_7466,N_7520);
and U9615 (N_9615,N_6293,N_6536);
and U9616 (N_9616,N_7470,N_7802);
xnor U9617 (N_9617,N_6305,N_6337);
nor U9618 (N_9618,N_7824,N_6708);
and U9619 (N_9619,N_7256,N_7072);
or U9620 (N_9620,N_7398,N_6732);
xor U9621 (N_9621,N_7569,N_7048);
nor U9622 (N_9622,N_6532,N_6775);
xnor U9623 (N_9623,N_7990,N_7092);
and U9624 (N_9624,N_6192,N_6396);
nor U9625 (N_9625,N_6204,N_6155);
nor U9626 (N_9626,N_7580,N_7324);
and U9627 (N_9627,N_7125,N_6386);
xnor U9628 (N_9628,N_7020,N_7312);
or U9629 (N_9629,N_6134,N_6816);
xor U9630 (N_9630,N_7569,N_6809);
xor U9631 (N_9631,N_7101,N_7028);
nor U9632 (N_9632,N_7265,N_6022);
xnor U9633 (N_9633,N_7643,N_7910);
and U9634 (N_9634,N_7709,N_6877);
xnor U9635 (N_9635,N_7067,N_7148);
and U9636 (N_9636,N_6091,N_7970);
and U9637 (N_9637,N_6127,N_7756);
nor U9638 (N_9638,N_7577,N_7374);
nor U9639 (N_9639,N_6298,N_7675);
nand U9640 (N_9640,N_7497,N_6505);
nand U9641 (N_9641,N_7018,N_7787);
xor U9642 (N_9642,N_7454,N_7480);
nor U9643 (N_9643,N_7602,N_6883);
xor U9644 (N_9644,N_7107,N_7173);
nor U9645 (N_9645,N_7596,N_6758);
and U9646 (N_9646,N_7787,N_6041);
xor U9647 (N_9647,N_7850,N_7866);
nor U9648 (N_9648,N_7139,N_7450);
xor U9649 (N_9649,N_7190,N_6891);
xor U9650 (N_9650,N_7382,N_6342);
nand U9651 (N_9651,N_6664,N_6917);
or U9652 (N_9652,N_6436,N_7381);
or U9653 (N_9653,N_7242,N_6183);
and U9654 (N_9654,N_6534,N_6740);
nor U9655 (N_9655,N_7610,N_6420);
nor U9656 (N_9656,N_7364,N_7259);
or U9657 (N_9657,N_6430,N_6824);
and U9658 (N_9658,N_6747,N_6168);
xor U9659 (N_9659,N_7168,N_6800);
and U9660 (N_9660,N_6489,N_7940);
nor U9661 (N_9661,N_7135,N_6374);
or U9662 (N_9662,N_7483,N_6672);
xor U9663 (N_9663,N_6746,N_6146);
and U9664 (N_9664,N_6429,N_7294);
or U9665 (N_9665,N_6179,N_6672);
or U9666 (N_9666,N_6104,N_6144);
or U9667 (N_9667,N_7173,N_6387);
nor U9668 (N_9668,N_6349,N_6741);
nand U9669 (N_9669,N_6536,N_7004);
nand U9670 (N_9670,N_7077,N_6349);
nand U9671 (N_9671,N_7883,N_7910);
xor U9672 (N_9672,N_6669,N_6354);
xor U9673 (N_9673,N_7721,N_6472);
nor U9674 (N_9674,N_7532,N_6489);
xnor U9675 (N_9675,N_6999,N_6746);
and U9676 (N_9676,N_7592,N_7832);
nand U9677 (N_9677,N_6381,N_6880);
xnor U9678 (N_9678,N_7192,N_7564);
nor U9679 (N_9679,N_7721,N_6701);
nand U9680 (N_9680,N_7425,N_6863);
nor U9681 (N_9681,N_7085,N_7615);
nand U9682 (N_9682,N_7344,N_6305);
xnor U9683 (N_9683,N_7526,N_7789);
or U9684 (N_9684,N_6574,N_7851);
nor U9685 (N_9685,N_6780,N_6023);
nand U9686 (N_9686,N_6324,N_7974);
nand U9687 (N_9687,N_6459,N_6908);
nand U9688 (N_9688,N_6729,N_6742);
or U9689 (N_9689,N_7048,N_7643);
or U9690 (N_9690,N_7031,N_6459);
xor U9691 (N_9691,N_6919,N_7725);
nand U9692 (N_9692,N_7859,N_6189);
xor U9693 (N_9693,N_6585,N_6205);
xor U9694 (N_9694,N_7796,N_7237);
nor U9695 (N_9695,N_7524,N_6901);
nand U9696 (N_9696,N_7207,N_7555);
nand U9697 (N_9697,N_7380,N_6880);
nor U9698 (N_9698,N_6380,N_6823);
nand U9699 (N_9699,N_7833,N_6407);
nand U9700 (N_9700,N_7635,N_6688);
nand U9701 (N_9701,N_6425,N_6407);
or U9702 (N_9702,N_6912,N_7545);
or U9703 (N_9703,N_6782,N_7525);
xor U9704 (N_9704,N_7555,N_7999);
xnor U9705 (N_9705,N_7681,N_6761);
or U9706 (N_9706,N_6188,N_6870);
xnor U9707 (N_9707,N_7702,N_6538);
nand U9708 (N_9708,N_6455,N_6939);
xnor U9709 (N_9709,N_7525,N_7160);
nor U9710 (N_9710,N_6653,N_6367);
xor U9711 (N_9711,N_7523,N_7913);
nor U9712 (N_9712,N_7511,N_7189);
nor U9713 (N_9713,N_6579,N_6924);
nor U9714 (N_9714,N_7394,N_7937);
xnor U9715 (N_9715,N_7482,N_7444);
xor U9716 (N_9716,N_6610,N_7133);
nand U9717 (N_9717,N_6132,N_6400);
or U9718 (N_9718,N_6313,N_7215);
nand U9719 (N_9719,N_7339,N_7297);
nor U9720 (N_9720,N_6337,N_6240);
xor U9721 (N_9721,N_7351,N_7668);
nand U9722 (N_9722,N_6591,N_7794);
xnor U9723 (N_9723,N_7000,N_6862);
nor U9724 (N_9724,N_6232,N_6276);
nand U9725 (N_9725,N_6157,N_7289);
xor U9726 (N_9726,N_7273,N_6033);
or U9727 (N_9727,N_7113,N_6666);
xnor U9728 (N_9728,N_7334,N_6688);
nand U9729 (N_9729,N_6287,N_6655);
and U9730 (N_9730,N_7525,N_6218);
xnor U9731 (N_9731,N_7675,N_7937);
or U9732 (N_9732,N_6791,N_6891);
nor U9733 (N_9733,N_7951,N_6709);
nor U9734 (N_9734,N_6202,N_7393);
and U9735 (N_9735,N_7933,N_7946);
xnor U9736 (N_9736,N_6206,N_7129);
nand U9737 (N_9737,N_6166,N_6290);
nor U9738 (N_9738,N_7378,N_7469);
and U9739 (N_9739,N_6602,N_6843);
or U9740 (N_9740,N_6240,N_6814);
nor U9741 (N_9741,N_6740,N_6444);
nand U9742 (N_9742,N_7039,N_6990);
or U9743 (N_9743,N_7293,N_6485);
and U9744 (N_9744,N_7493,N_6921);
and U9745 (N_9745,N_6188,N_7805);
nand U9746 (N_9746,N_7639,N_7156);
or U9747 (N_9747,N_6114,N_6230);
xnor U9748 (N_9748,N_7374,N_6712);
nor U9749 (N_9749,N_7650,N_6016);
nand U9750 (N_9750,N_6778,N_7625);
or U9751 (N_9751,N_6424,N_7912);
nor U9752 (N_9752,N_7816,N_7405);
nor U9753 (N_9753,N_7650,N_7195);
or U9754 (N_9754,N_6275,N_6073);
nor U9755 (N_9755,N_7507,N_7385);
and U9756 (N_9756,N_7960,N_6839);
xor U9757 (N_9757,N_6217,N_7621);
nand U9758 (N_9758,N_6255,N_6879);
or U9759 (N_9759,N_6008,N_6918);
nor U9760 (N_9760,N_7680,N_6653);
nor U9761 (N_9761,N_7285,N_6149);
and U9762 (N_9762,N_6771,N_6778);
or U9763 (N_9763,N_6611,N_6916);
nor U9764 (N_9764,N_7365,N_6896);
or U9765 (N_9765,N_7536,N_6134);
nand U9766 (N_9766,N_6895,N_6386);
nand U9767 (N_9767,N_7451,N_6810);
or U9768 (N_9768,N_7056,N_7070);
nand U9769 (N_9769,N_7689,N_7004);
or U9770 (N_9770,N_7156,N_7744);
or U9771 (N_9771,N_7821,N_6589);
xnor U9772 (N_9772,N_6029,N_6378);
nor U9773 (N_9773,N_6729,N_6472);
and U9774 (N_9774,N_7886,N_6723);
and U9775 (N_9775,N_6944,N_6793);
nand U9776 (N_9776,N_6181,N_7096);
nor U9777 (N_9777,N_7006,N_7273);
and U9778 (N_9778,N_7953,N_6817);
or U9779 (N_9779,N_7265,N_7181);
or U9780 (N_9780,N_7879,N_6476);
and U9781 (N_9781,N_7440,N_7786);
and U9782 (N_9782,N_7173,N_6207);
xnor U9783 (N_9783,N_7830,N_7556);
or U9784 (N_9784,N_6463,N_6007);
nand U9785 (N_9785,N_6533,N_7411);
nand U9786 (N_9786,N_6327,N_6005);
and U9787 (N_9787,N_6754,N_7363);
nor U9788 (N_9788,N_6928,N_7028);
nor U9789 (N_9789,N_7813,N_7105);
and U9790 (N_9790,N_6818,N_7853);
xnor U9791 (N_9791,N_6853,N_7874);
nand U9792 (N_9792,N_7118,N_7019);
nor U9793 (N_9793,N_6921,N_7513);
and U9794 (N_9794,N_6741,N_6619);
or U9795 (N_9795,N_7616,N_7214);
and U9796 (N_9796,N_6583,N_6979);
nor U9797 (N_9797,N_6413,N_7084);
xor U9798 (N_9798,N_7838,N_6464);
nor U9799 (N_9799,N_7546,N_7587);
or U9800 (N_9800,N_7982,N_6432);
nor U9801 (N_9801,N_6793,N_6729);
and U9802 (N_9802,N_6237,N_6574);
nor U9803 (N_9803,N_7430,N_6225);
or U9804 (N_9804,N_7311,N_7945);
xnor U9805 (N_9805,N_7214,N_7325);
and U9806 (N_9806,N_7411,N_7908);
and U9807 (N_9807,N_6858,N_6029);
or U9808 (N_9808,N_7596,N_6117);
xnor U9809 (N_9809,N_6872,N_6458);
xnor U9810 (N_9810,N_6693,N_7370);
nand U9811 (N_9811,N_7059,N_7187);
or U9812 (N_9812,N_7317,N_6242);
or U9813 (N_9813,N_7797,N_7309);
nor U9814 (N_9814,N_6635,N_6585);
nand U9815 (N_9815,N_7653,N_7497);
and U9816 (N_9816,N_7236,N_7124);
nand U9817 (N_9817,N_6754,N_6512);
nand U9818 (N_9818,N_6781,N_7252);
and U9819 (N_9819,N_6665,N_6620);
xor U9820 (N_9820,N_7025,N_6578);
xnor U9821 (N_9821,N_7654,N_7058);
and U9822 (N_9822,N_6712,N_7720);
nor U9823 (N_9823,N_7699,N_6311);
and U9824 (N_9824,N_7957,N_7711);
nor U9825 (N_9825,N_6089,N_7454);
and U9826 (N_9826,N_7254,N_7095);
nor U9827 (N_9827,N_6113,N_7727);
and U9828 (N_9828,N_7493,N_6471);
nor U9829 (N_9829,N_6836,N_7877);
or U9830 (N_9830,N_7152,N_7719);
and U9831 (N_9831,N_6981,N_7270);
xnor U9832 (N_9832,N_7024,N_6098);
nand U9833 (N_9833,N_6291,N_7147);
or U9834 (N_9834,N_7045,N_7918);
nand U9835 (N_9835,N_7105,N_6018);
and U9836 (N_9836,N_7966,N_6265);
nand U9837 (N_9837,N_7574,N_7761);
nand U9838 (N_9838,N_7173,N_7073);
or U9839 (N_9839,N_7274,N_6688);
and U9840 (N_9840,N_6051,N_6059);
and U9841 (N_9841,N_7867,N_7459);
nor U9842 (N_9842,N_6941,N_6444);
xor U9843 (N_9843,N_6190,N_7101);
or U9844 (N_9844,N_6764,N_6883);
and U9845 (N_9845,N_7715,N_6508);
and U9846 (N_9846,N_7580,N_6935);
xor U9847 (N_9847,N_7414,N_6338);
or U9848 (N_9848,N_7454,N_6519);
or U9849 (N_9849,N_6864,N_7928);
xnor U9850 (N_9850,N_6441,N_6105);
nand U9851 (N_9851,N_7512,N_6763);
or U9852 (N_9852,N_6399,N_7044);
nor U9853 (N_9853,N_6830,N_6279);
nor U9854 (N_9854,N_6741,N_7771);
or U9855 (N_9855,N_7813,N_6847);
xnor U9856 (N_9856,N_7234,N_6946);
xnor U9857 (N_9857,N_7752,N_6042);
or U9858 (N_9858,N_6722,N_6407);
or U9859 (N_9859,N_7147,N_6413);
nor U9860 (N_9860,N_6580,N_7500);
nand U9861 (N_9861,N_6619,N_7444);
and U9862 (N_9862,N_7674,N_7163);
nand U9863 (N_9863,N_7844,N_7383);
xor U9864 (N_9864,N_6618,N_7738);
nor U9865 (N_9865,N_6220,N_6882);
nor U9866 (N_9866,N_7342,N_6673);
and U9867 (N_9867,N_7749,N_7542);
or U9868 (N_9868,N_7190,N_7407);
nand U9869 (N_9869,N_6861,N_6010);
nor U9870 (N_9870,N_7840,N_6789);
xnor U9871 (N_9871,N_7152,N_6272);
nand U9872 (N_9872,N_7392,N_6093);
xor U9873 (N_9873,N_7130,N_6801);
or U9874 (N_9874,N_7470,N_6013);
and U9875 (N_9875,N_7181,N_6874);
xnor U9876 (N_9876,N_6030,N_6034);
and U9877 (N_9877,N_6076,N_6388);
nand U9878 (N_9878,N_7003,N_7484);
xnor U9879 (N_9879,N_6081,N_6548);
or U9880 (N_9880,N_7076,N_7934);
and U9881 (N_9881,N_6718,N_7091);
nand U9882 (N_9882,N_6011,N_7926);
or U9883 (N_9883,N_6604,N_6357);
nor U9884 (N_9884,N_7755,N_6955);
or U9885 (N_9885,N_7801,N_7800);
nor U9886 (N_9886,N_6859,N_7862);
nand U9887 (N_9887,N_7203,N_7879);
or U9888 (N_9888,N_6844,N_7887);
and U9889 (N_9889,N_7824,N_7498);
nand U9890 (N_9890,N_6061,N_7204);
xnor U9891 (N_9891,N_7843,N_7638);
xor U9892 (N_9892,N_6226,N_7969);
nor U9893 (N_9893,N_7753,N_7337);
nand U9894 (N_9894,N_7168,N_6469);
and U9895 (N_9895,N_6467,N_6292);
xor U9896 (N_9896,N_6260,N_7146);
nor U9897 (N_9897,N_7897,N_7860);
and U9898 (N_9898,N_7494,N_7040);
nand U9899 (N_9899,N_6654,N_6191);
nor U9900 (N_9900,N_6944,N_6595);
or U9901 (N_9901,N_7247,N_7308);
nor U9902 (N_9902,N_7454,N_7580);
nor U9903 (N_9903,N_6466,N_7533);
xor U9904 (N_9904,N_6803,N_7180);
xor U9905 (N_9905,N_7993,N_6831);
nand U9906 (N_9906,N_6561,N_6366);
xnor U9907 (N_9907,N_7361,N_6404);
nor U9908 (N_9908,N_7985,N_6955);
nor U9909 (N_9909,N_7954,N_7793);
xor U9910 (N_9910,N_6136,N_6296);
nand U9911 (N_9911,N_6763,N_6821);
or U9912 (N_9912,N_7499,N_6381);
or U9913 (N_9913,N_6366,N_6873);
nor U9914 (N_9914,N_7563,N_7941);
nand U9915 (N_9915,N_7825,N_6958);
nand U9916 (N_9916,N_6663,N_7192);
xnor U9917 (N_9917,N_6868,N_7884);
and U9918 (N_9918,N_6489,N_7506);
xor U9919 (N_9919,N_7157,N_7793);
and U9920 (N_9920,N_7526,N_6181);
xnor U9921 (N_9921,N_7291,N_7544);
and U9922 (N_9922,N_7438,N_6423);
and U9923 (N_9923,N_7775,N_7818);
nand U9924 (N_9924,N_6115,N_6944);
xor U9925 (N_9925,N_6682,N_7152);
nor U9926 (N_9926,N_7302,N_6093);
xor U9927 (N_9927,N_7883,N_6746);
nand U9928 (N_9928,N_6371,N_6582);
or U9929 (N_9929,N_6576,N_7056);
xor U9930 (N_9930,N_7989,N_7532);
and U9931 (N_9931,N_6603,N_6616);
xor U9932 (N_9932,N_7217,N_7698);
or U9933 (N_9933,N_7877,N_6602);
nand U9934 (N_9934,N_7266,N_6346);
or U9935 (N_9935,N_7720,N_7745);
nand U9936 (N_9936,N_7265,N_6289);
nor U9937 (N_9937,N_7329,N_7344);
nand U9938 (N_9938,N_6648,N_6139);
nand U9939 (N_9939,N_7327,N_6082);
and U9940 (N_9940,N_7535,N_7016);
nand U9941 (N_9941,N_7928,N_7075);
xor U9942 (N_9942,N_6765,N_6860);
xnor U9943 (N_9943,N_7427,N_7329);
and U9944 (N_9944,N_6577,N_7299);
nor U9945 (N_9945,N_6426,N_6601);
and U9946 (N_9946,N_7775,N_7483);
nand U9947 (N_9947,N_7426,N_6754);
and U9948 (N_9948,N_6105,N_6553);
xnor U9949 (N_9949,N_7948,N_6207);
or U9950 (N_9950,N_7829,N_6599);
nor U9951 (N_9951,N_7270,N_6218);
and U9952 (N_9952,N_6513,N_6392);
and U9953 (N_9953,N_7643,N_7602);
or U9954 (N_9954,N_7658,N_6403);
xnor U9955 (N_9955,N_6431,N_6880);
nor U9956 (N_9956,N_6443,N_6470);
nor U9957 (N_9957,N_6143,N_7554);
or U9958 (N_9958,N_6579,N_7526);
and U9959 (N_9959,N_6509,N_6098);
nor U9960 (N_9960,N_7733,N_6471);
and U9961 (N_9961,N_7558,N_7172);
or U9962 (N_9962,N_7926,N_6455);
nor U9963 (N_9963,N_7484,N_6303);
nor U9964 (N_9964,N_6926,N_6793);
and U9965 (N_9965,N_6472,N_6309);
or U9966 (N_9966,N_6919,N_7366);
xor U9967 (N_9967,N_7885,N_6129);
and U9968 (N_9968,N_6271,N_7310);
xnor U9969 (N_9969,N_7758,N_7911);
xor U9970 (N_9970,N_7676,N_7073);
nor U9971 (N_9971,N_6854,N_6489);
or U9972 (N_9972,N_6610,N_6120);
xor U9973 (N_9973,N_7629,N_7468);
xnor U9974 (N_9974,N_6654,N_7012);
or U9975 (N_9975,N_6700,N_6641);
or U9976 (N_9976,N_6159,N_7800);
and U9977 (N_9977,N_6623,N_6075);
or U9978 (N_9978,N_7600,N_7309);
nor U9979 (N_9979,N_7359,N_7711);
xnor U9980 (N_9980,N_7366,N_7111);
nand U9981 (N_9981,N_6535,N_6072);
xnor U9982 (N_9982,N_6228,N_7892);
nor U9983 (N_9983,N_7071,N_7604);
or U9984 (N_9984,N_7974,N_6010);
xnor U9985 (N_9985,N_6376,N_6445);
xor U9986 (N_9986,N_7811,N_6958);
nand U9987 (N_9987,N_7321,N_6710);
or U9988 (N_9988,N_7397,N_6494);
xnor U9989 (N_9989,N_7034,N_6282);
or U9990 (N_9990,N_6745,N_6812);
and U9991 (N_9991,N_7928,N_6694);
nor U9992 (N_9992,N_6325,N_6036);
xor U9993 (N_9993,N_7692,N_7252);
or U9994 (N_9994,N_7824,N_7859);
nand U9995 (N_9995,N_6365,N_6538);
nand U9996 (N_9996,N_7440,N_6605);
xnor U9997 (N_9997,N_6694,N_7650);
and U9998 (N_9998,N_6501,N_6295);
or U9999 (N_9999,N_7423,N_6229);
and UO_0 (O_0,N_8077,N_9448);
or UO_1 (O_1,N_9904,N_9644);
and UO_2 (O_2,N_8532,N_8316);
nor UO_3 (O_3,N_9376,N_8144);
nor UO_4 (O_4,N_8783,N_9091);
or UO_5 (O_5,N_8707,N_9514);
or UO_6 (O_6,N_8001,N_8305);
nand UO_7 (O_7,N_8009,N_8087);
nor UO_8 (O_8,N_8459,N_9313);
nor UO_9 (O_9,N_8153,N_9931);
xnor UO_10 (O_10,N_8138,N_8996);
or UO_11 (O_11,N_8614,N_8979);
and UO_12 (O_12,N_9192,N_9955);
and UO_13 (O_13,N_9563,N_9092);
xnor UO_14 (O_14,N_9872,N_9315);
nor UO_15 (O_15,N_9000,N_9842);
xnor UO_16 (O_16,N_9981,N_8067);
xnor UO_17 (O_17,N_9673,N_8751);
or UO_18 (O_18,N_9760,N_8274);
and UO_19 (O_19,N_9659,N_9260);
xor UO_20 (O_20,N_9402,N_9160);
or UO_21 (O_21,N_8368,N_9466);
or UO_22 (O_22,N_8580,N_8506);
nand UO_23 (O_23,N_8589,N_9397);
or UO_24 (O_24,N_9609,N_8060);
xnor UO_25 (O_25,N_9972,N_8457);
nor UO_26 (O_26,N_9636,N_8257);
xor UO_27 (O_27,N_8984,N_8334);
xnor UO_28 (O_28,N_9574,N_9196);
or UO_29 (O_29,N_9079,N_9984);
nand UO_30 (O_30,N_9542,N_8466);
xnor UO_31 (O_31,N_9925,N_9068);
nor UO_32 (O_32,N_9915,N_9430);
or UO_33 (O_33,N_9181,N_8072);
and UO_34 (O_34,N_9346,N_8878);
nor UO_35 (O_35,N_8268,N_8544);
nand UO_36 (O_36,N_9861,N_9483);
and UO_37 (O_37,N_8795,N_8727);
nor UO_38 (O_38,N_9982,N_8374);
nand UO_39 (O_39,N_8190,N_8876);
xor UO_40 (O_40,N_8729,N_8345);
and UO_41 (O_41,N_8481,N_9805);
and UO_42 (O_42,N_8218,N_9395);
or UO_43 (O_43,N_9441,N_9611);
nor UO_44 (O_44,N_9713,N_9886);
and UO_45 (O_45,N_9967,N_9628);
xnor UO_46 (O_46,N_9491,N_8447);
and UO_47 (O_47,N_8275,N_9663);
xor UO_48 (O_48,N_9345,N_8663);
nand UO_49 (O_49,N_9794,N_9929);
xor UO_50 (O_50,N_8645,N_9113);
and UO_51 (O_51,N_9490,N_9923);
and UO_52 (O_52,N_8206,N_9961);
nand UO_53 (O_53,N_9950,N_9185);
and UO_54 (O_54,N_9899,N_9729);
or UO_55 (O_55,N_9164,N_8098);
or UO_56 (O_56,N_8145,N_9791);
xor UO_57 (O_57,N_8109,N_9747);
nor UO_58 (O_58,N_9064,N_8562);
nor UO_59 (O_59,N_8255,N_9905);
or UO_60 (O_60,N_9833,N_8025);
and UO_61 (O_61,N_8390,N_8763);
nor UO_62 (O_62,N_8285,N_8664);
and UO_63 (O_63,N_8587,N_9184);
nand UO_64 (O_64,N_9549,N_8963);
nor UO_65 (O_65,N_8628,N_8529);
and UO_66 (O_66,N_9369,N_9204);
and UO_67 (O_67,N_8982,N_8592);
nand UO_68 (O_68,N_9429,N_9567);
and UO_69 (O_69,N_9485,N_8930);
or UO_70 (O_70,N_9585,N_8248);
xor UO_71 (O_71,N_8335,N_9523);
nor UO_72 (O_72,N_9745,N_9414);
nand UO_73 (O_73,N_8643,N_8215);
or UO_74 (O_74,N_9042,N_8995);
or UO_75 (O_75,N_9170,N_9048);
nand UO_76 (O_76,N_9434,N_8759);
and UO_77 (O_77,N_8871,N_9605);
nand UO_78 (O_78,N_9377,N_9386);
or UO_79 (O_79,N_8053,N_8219);
nor UO_80 (O_80,N_9560,N_9634);
nand UO_81 (O_81,N_8208,N_9247);
xor UO_82 (O_82,N_9057,N_8801);
and UO_83 (O_83,N_8442,N_8868);
nand UO_84 (O_84,N_9538,N_8385);
nor UO_85 (O_85,N_9203,N_9056);
nand UO_86 (O_86,N_8910,N_8968);
and UO_87 (O_87,N_9174,N_8292);
xor UO_88 (O_88,N_8678,N_8976);
nand UO_89 (O_89,N_9591,N_9916);
nor UO_90 (O_90,N_8955,N_8843);
nand UO_91 (O_91,N_8071,N_9578);
nor UO_92 (O_92,N_8304,N_9657);
and UO_93 (O_93,N_9069,N_8018);
and UO_94 (O_94,N_8321,N_9977);
nor UO_95 (O_95,N_9324,N_8118);
nor UO_96 (O_96,N_9935,N_8586);
xnor UO_97 (O_97,N_8437,N_9245);
nand UO_98 (O_98,N_8617,N_8943);
xor UO_99 (O_99,N_9654,N_9257);
or UO_100 (O_100,N_8970,N_9444);
nor UO_101 (O_101,N_9703,N_9431);
xor UO_102 (O_102,N_9515,N_8739);
and UO_103 (O_103,N_8822,N_9723);
and UO_104 (O_104,N_9387,N_8119);
nand UO_105 (O_105,N_8012,N_9679);
or UO_106 (O_106,N_9014,N_9843);
nor UO_107 (O_107,N_8901,N_9891);
nor UO_108 (O_108,N_8396,N_9074);
and UO_109 (O_109,N_9734,N_8440);
nand UO_110 (O_110,N_8301,N_8768);
or UO_111 (O_111,N_9777,N_8735);
or UO_112 (O_112,N_8757,N_8567);
nand UO_113 (O_113,N_9357,N_9761);
nor UO_114 (O_114,N_8687,N_8819);
nand UO_115 (O_115,N_8461,N_8046);
or UO_116 (O_116,N_8883,N_8927);
nand UO_117 (O_117,N_9894,N_9642);
nand UO_118 (O_118,N_8836,N_8692);
nor UO_119 (O_119,N_8662,N_8553);
nand UO_120 (O_120,N_8043,N_9507);
xor UO_121 (O_121,N_9613,N_8841);
and UO_122 (O_122,N_9841,N_8343);
nor UO_123 (O_123,N_8900,N_8498);
nor UO_124 (O_124,N_9472,N_8347);
nand UO_125 (O_125,N_9985,N_9211);
nand UO_126 (O_126,N_8517,N_9171);
nand UO_127 (O_127,N_8603,N_8044);
nand UO_128 (O_128,N_9053,N_9695);
and UO_129 (O_129,N_9142,N_9367);
nand UO_130 (O_130,N_9385,N_8887);
nand UO_131 (O_131,N_9090,N_9913);
or UO_132 (O_132,N_8430,N_9311);
xnor UO_133 (O_133,N_8004,N_8752);
xnor UO_134 (O_134,N_8642,N_9329);
or UO_135 (O_135,N_8839,N_9532);
xor UO_136 (O_136,N_9361,N_8547);
and UO_137 (O_137,N_8282,N_9944);
nand UO_138 (O_138,N_9751,N_8740);
xor UO_139 (O_139,N_8624,N_8157);
and UO_140 (O_140,N_9295,N_8113);
nor UO_141 (O_141,N_8496,N_8188);
nand UO_142 (O_142,N_9284,N_8055);
xnor UO_143 (O_143,N_8908,N_9219);
nand UO_144 (O_144,N_9059,N_9946);
nor UO_145 (O_145,N_8332,N_9824);
or UO_146 (O_146,N_9782,N_8658);
xnor UO_147 (O_147,N_9482,N_8407);
and UO_148 (O_148,N_9933,N_9240);
or UO_149 (O_149,N_8639,N_8226);
and UO_150 (O_150,N_9270,N_8837);
or UO_151 (O_151,N_9922,N_9502);
and UO_152 (O_152,N_8370,N_9772);
or UO_153 (O_153,N_9403,N_9648);
nor UO_154 (O_154,N_8400,N_8967);
or UO_155 (O_155,N_9137,N_8718);
xnor UO_156 (O_156,N_9105,N_8183);
nor UO_157 (O_157,N_8748,N_8135);
nor UO_158 (O_158,N_9034,N_9691);
xor UO_159 (O_159,N_9802,N_9653);
and UO_160 (O_160,N_9660,N_8092);
and UO_161 (O_161,N_9023,N_9550);
nand UO_162 (O_162,N_9162,N_8076);
or UO_163 (O_163,N_9312,N_8936);
nor UO_164 (O_164,N_8942,N_8749);
and UO_165 (O_165,N_8129,N_8796);
or UO_166 (O_166,N_8638,N_9154);
or UO_167 (O_167,N_9350,N_8675);
nand UO_168 (O_168,N_9531,N_8328);
nand UO_169 (O_169,N_8480,N_9603);
xor UO_170 (O_170,N_9635,N_8656);
nand UO_171 (O_171,N_9305,N_8916);
xor UO_172 (O_172,N_9117,N_8325);
or UO_173 (O_173,N_9631,N_9697);
and UO_174 (O_174,N_8699,N_8339);
and UO_175 (O_175,N_8929,N_8957);
nand UO_176 (O_176,N_8703,N_8201);
xor UO_177 (O_177,N_8766,N_9216);
xnor UO_178 (O_178,N_9340,N_8753);
or UO_179 (O_179,N_9474,N_8175);
xor UO_180 (O_180,N_8196,N_9980);
or UO_181 (O_181,N_8422,N_8288);
nor UO_182 (O_182,N_8291,N_8170);
nand UO_183 (O_183,N_8243,N_9063);
or UO_184 (O_184,N_8991,N_8512);
xnor UO_185 (O_185,N_8006,N_9365);
nor UO_186 (O_186,N_9363,N_8846);
xor UO_187 (O_187,N_9051,N_8919);
xnor UO_188 (O_188,N_8971,N_9727);
xnor UO_189 (O_189,N_8487,N_9537);
nand UO_190 (O_190,N_8633,N_8915);
or UO_191 (O_191,N_8922,N_9276);
or UO_192 (O_192,N_8682,N_9382);
nor UO_193 (O_193,N_8232,N_9237);
and UO_194 (O_194,N_9986,N_8027);
xor UO_195 (O_195,N_9764,N_9807);
or UO_196 (O_196,N_9853,N_9143);
xnor UO_197 (O_197,N_8572,N_9762);
nor UO_198 (O_198,N_9867,N_9140);
or UO_199 (O_199,N_9887,N_9469);
xnor UO_200 (O_200,N_8420,N_8808);
and UO_201 (O_201,N_8490,N_8371);
xnor UO_202 (O_202,N_8738,N_8398);
or UO_203 (O_203,N_9716,N_8142);
xor UO_204 (O_204,N_9783,N_9880);
xor UO_205 (O_205,N_8786,N_8804);
or UO_206 (O_206,N_9004,N_9597);
xnor UO_207 (O_207,N_8431,N_9138);
and UO_208 (O_208,N_8676,N_8174);
or UO_209 (O_209,N_8668,N_9808);
xor UO_210 (O_210,N_8284,N_8097);
nand UO_211 (O_211,N_8575,N_9581);
and UO_212 (O_212,N_8254,N_8935);
nand UO_213 (O_213,N_8000,N_9683);
nor UO_214 (O_214,N_9266,N_8531);
or UO_215 (O_215,N_9874,N_9306);
or UO_216 (O_216,N_8697,N_9384);
nand UO_217 (O_217,N_9071,N_9655);
nor UO_218 (O_218,N_8404,N_9375);
nand UO_219 (O_219,N_8425,N_8107);
nand UO_220 (O_220,N_8181,N_8228);
and UO_221 (O_221,N_9032,N_9208);
xnor UO_222 (O_222,N_8754,N_9478);
xnor UO_223 (O_223,N_8256,N_8652);
xnor UO_224 (O_224,N_8880,N_8171);
or UO_225 (O_225,N_8485,N_8432);
or UO_226 (O_226,N_9519,N_9975);
xor UO_227 (O_227,N_8148,N_9073);
nand UO_228 (O_228,N_8610,N_8177);
xnor UO_229 (O_229,N_8497,N_8903);
nand UO_230 (O_230,N_8482,N_8378);
nor UO_231 (O_231,N_9547,N_9262);
or UO_232 (O_232,N_9333,N_8261);
and UO_233 (O_233,N_9912,N_8019);
nor UO_234 (O_234,N_8117,N_8478);
and UO_235 (O_235,N_8413,N_9766);
xor UO_236 (O_236,N_8618,N_9493);
xor UO_237 (O_237,N_8913,N_9987);
nand UO_238 (O_238,N_8045,N_8890);
and UO_239 (O_239,N_9393,N_9036);
nor UO_240 (O_240,N_8300,N_8262);
nand UO_241 (O_241,N_9293,N_9152);
nor UO_242 (O_242,N_8665,N_9871);
and UO_243 (O_243,N_8809,N_9030);
nor UO_244 (O_244,N_8124,N_8007);
or UO_245 (O_245,N_8093,N_9383);
xnor UO_246 (O_246,N_9706,N_8221);
and UO_247 (O_247,N_8829,N_8911);
xnor UO_248 (O_248,N_8838,N_8462);
nand UO_249 (O_249,N_9263,N_8015);
or UO_250 (O_250,N_8962,N_8319);
nor UO_251 (O_251,N_9238,N_8975);
or UO_252 (O_252,N_9358,N_8845);
and UO_253 (O_253,N_8944,N_8269);
and UO_254 (O_254,N_9062,N_9755);
and UO_255 (O_255,N_9845,N_9738);
and UO_256 (O_256,N_8778,N_8120);
and UO_257 (O_257,N_8985,N_8090);
nor UO_258 (O_258,N_9781,N_9161);
or UO_259 (O_259,N_8165,N_9684);
nand UO_260 (O_260,N_9167,N_8353);
nor UO_261 (O_261,N_8785,N_9970);
and UO_262 (O_262,N_9918,N_8428);
nand UO_263 (O_263,N_9280,N_8225);
nand UO_264 (O_264,N_8755,N_9480);
xor UO_265 (O_265,N_9804,N_9689);
and UO_266 (O_266,N_9951,N_9509);
or UO_267 (O_267,N_9629,N_9742);
and UO_268 (O_268,N_9598,N_9948);
or UO_269 (O_269,N_9390,N_9910);
nand UO_270 (O_270,N_9331,N_8426);
or UO_271 (O_271,N_9744,N_8460);
or UO_272 (O_272,N_9615,N_9733);
nor UO_273 (O_273,N_9341,N_8094);
or UO_274 (O_274,N_9121,N_9234);
and UO_275 (O_275,N_8777,N_9834);
xor UO_276 (O_276,N_9486,N_9873);
nor UO_277 (O_277,N_9990,N_8865);
nand UO_278 (O_278,N_8105,N_9645);
or UO_279 (O_279,N_8508,N_8861);
and UO_280 (O_280,N_9244,N_8905);
and UO_281 (O_281,N_9667,N_8894);
and UO_282 (O_282,N_8156,N_9038);
nand UO_283 (O_283,N_8810,N_8881);
and UO_284 (O_284,N_9132,N_8688);
nor UO_285 (O_285,N_9811,N_9799);
or UO_286 (O_286,N_9124,N_8561);
nor UO_287 (O_287,N_9296,N_8143);
nor UO_288 (O_288,N_9190,N_9131);
or UO_289 (O_289,N_9666,N_8032);
or UO_290 (O_290,N_8030,N_8443);
nor UO_291 (O_291,N_8276,N_8973);
xor UO_292 (O_292,N_8198,N_8799);
or UO_293 (O_293,N_8635,N_9269);
xor UO_294 (O_294,N_8731,N_9018);
and UO_295 (O_295,N_8978,N_9565);
and UO_296 (O_296,N_8102,N_8702);
nand UO_297 (O_297,N_8691,N_9498);
xor UO_298 (O_298,N_8349,N_9819);
nor UO_299 (O_299,N_9106,N_9649);
nor UO_300 (O_300,N_8902,N_8031);
nand UO_301 (O_301,N_9839,N_8251);
and UO_302 (O_302,N_8684,N_9278);
and UO_303 (O_303,N_8271,N_8560);
or UO_304 (O_304,N_9327,N_8690);
or UO_305 (O_305,N_8059,N_8336);
and UO_306 (O_306,N_9226,N_8010);
nand UO_307 (O_307,N_9086,N_8854);
or UO_308 (O_308,N_9870,N_9854);
and UO_309 (O_309,N_8331,N_8539);
nand UO_310 (O_310,N_9851,N_8577);
or UO_311 (O_311,N_8199,N_9347);
nor UO_312 (O_312,N_9662,N_8281);
xor UO_313 (O_313,N_9878,N_9651);
nor UO_314 (O_314,N_8080,N_8486);
nand UO_315 (O_315,N_9436,N_8303);
xnor UO_316 (O_316,N_8146,N_9176);
or UO_317 (O_317,N_9129,N_9488);
nor UO_318 (O_318,N_9453,N_8619);
nand UO_319 (O_319,N_8666,N_8264);
or UO_320 (O_320,N_9011,N_9020);
and UO_321 (O_321,N_9309,N_9299);
or UO_322 (O_322,N_9909,N_8952);
or UO_323 (O_323,N_9954,N_9594);
xor UO_324 (O_324,N_8403,N_8657);
and UO_325 (O_325,N_9855,N_9089);
nand UO_326 (O_326,N_9774,N_9556);
nand UO_327 (O_327,N_9338,N_9144);
xnor UO_328 (O_328,N_9837,N_9499);
nand UO_329 (O_329,N_9194,N_9731);
and UO_330 (O_330,N_9380,N_9426);
and UO_331 (O_331,N_8949,N_8946);
and UO_332 (O_332,N_8121,N_9463);
and UO_333 (O_333,N_9750,N_8953);
and UO_334 (O_334,N_9516,N_9754);
nand UO_335 (O_335,N_9792,N_8095);
and UO_336 (O_336,N_8528,N_8863);
nand UO_337 (O_337,N_8859,N_8600);
nand UO_338 (O_338,N_9024,N_9302);
nor UO_339 (O_339,N_9103,N_8246);
and UO_340 (O_340,N_9116,N_9720);
or UO_341 (O_341,N_9398,N_8815);
or UO_342 (O_342,N_8802,N_9465);
or UO_343 (O_343,N_8020,N_8858);
nor UO_344 (O_344,N_9107,N_9177);
xor UO_345 (O_345,N_8320,N_9561);
nand UO_346 (O_346,N_9052,N_9520);
nand UO_347 (O_347,N_9054,N_9183);
and UO_348 (O_348,N_9388,N_8834);
or UO_349 (O_349,N_8611,N_9829);
and UO_350 (O_350,N_8653,N_8794);
or UO_351 (O_351,N_8314,N_9566);
xor UO_352 (O_352,N_8200,N_8393);
xnor UO_353 (O_353,N_9087,N_9310);
and UO_354 (O_354,N_9814,N_9971);
nor UO_355 (O_355,N_8523,N_9021);
and UO_356 (O_356,N_8563,N_8989);
nand UO_357 (O_357,N_8601,N_8082);
and UO_358 (O_358,N_9722,N_9902);
and UO_359 (O_359,N_8022,N_8538);
or UO_360 (O_360,N_9707,N_8340);
and UO_361 (O_361,N_8111,N_8698);
and UO_362 (O_362,N_9844,N_8874);
xor UO_363 (O_363,N_8217,N_8453);
and UO_364 (O_364,N_9864,N_9865);
nor UO_365 (O_365,N_9359,N_8917);
xnor UO_366 (O_366,N_9067,N_9608);
and UO_367 (O_367,N_8747,N_9290);
or UO_368 (O_368,N_8667,N_9890);
xnor UO_369 (O_369,N_8886,N_9626);
nand UO_370 (O_370,N_9558,N_8410);
nand UO_371 (O_371,N_9253,N_8730);
and UO_372 (O_372,N_9224,N_9193);
or UO_373 (O_373,N_8279,N_9155);
nand UO_374 (O_374,N_9632,N_9746);
xnor UO_375 (O_375,N_8445,N_8625);
nand UO_376 (O_376,N_9010,N_8631);
nor UO_377 (O_377,N_9885,N_9505);
and UO_378 (O_378,N_8354,N_8849);
and UO_379 (O_379,N_9687,N_8835);
or UO_380 (O_380,N_9786,N_8324);
nand UO_381 (O_381,N_8286,N_9378);
and UO_382 (O_382,N_8184,N_8266);
nand UO_383 (O_383,N_9571,N_9432);
and UO_384 (O_384,N_9039,N_9652);
xnor UO_385 (O_385,N_9371,N_8405);
and UO_386 (O_386,N_8923,N_8632);
and UO_387 (O_387,N_8051,N_9433);
xor UO_388 (O_388,N_9153,N_8724);
nand UO_389 (O_389,N_9801,N_9570);
or UO_390 (O_390,N_9416,N_8524);
nand UO_391 (O_391,N_8627,N_9055);
or UO_392 (O_392,N_8062,N_9267);
and UO_393 (O_393,N_9476,N_9821);
nand UO_394 (O_394,N_8192,N_9647);
nand UO_395 (O_395,N_8709,N_9228);
nand UO_396 (O_396,N_9724,N_9254);
or UO_397 (O_397,N_8502,N_8151);
and UO_398 (O_398,N_9535,N_8693);
or UO_399 (O_399,N_9927,N_8351);
or UO_400 (O_400,N_9941,N_8162);
or UO_401 (O_401,N_8864,N_8745);
and UO_402 (O_402,N_8535,N_9728);
nor UO_403 (O_403,N_9085,N_8411);
nor UO_404 (O_404,N_9188,N_9881);
xor UO_405 (O_405,N_9205,N_8939);
xnor UO_406 (O_406,N_8551,N_9770);
or UO_407 (O_407,N_9404,N_8594);
or UO_408 (O_408,N_9953,N_8770);
nor UO_409 (O_409,N_8756,N_9451);
and UO_410 (O_410,N_8429,N_8714);
and UO_411 (O_411,N_9417,N_9627);
nor UO_412 (O_412,N_9527,N_8623);
xor UO_413 (O_413,N_8089,N_8484);
xor UO_414 (O_414,N_8207,N_9582);
xnor UO_415 (O_415,N_9355,N_9304);
xnor UO_416 (O_416,N_9449,N_9593);
and UO_417 (O_417,N_9209,N_8501);
or UO_418 (O_418,N_9572,N_9119);
and UO_419 (O_419,N_8108,N_9595);
or UO_420 (O_420,N_9856,N_9836);
or UO_421 (O_421,N_9831,N_8602);
xnor UO_422 (O_422,N_9440,N_9037);
nand UO_423 (O_423,N_8290,N_8595);
xor UO_424 (O_424,N_8408,N_9793);
xnor UO_425 (O_425,N_9031,N_9623);
nor UO_426 (O_426,N_9335,N_8193);
xor UO_427 (O_427,N_8161,N_9008);
xnor UO_428 (O_428,N_8115,N_8350);
nor UO_429 (O_429,N_9145,N_8139);
xnor UO_430 (O_430,N_9568,N_8220);
xnor UO_431 (O_431,N_9962,N_8681);
and UO_432 (O_432,N_8541,N_9093);
nand UO_433 (O_433,N_8516,N_8372);
nand UO_434 (O_434,N_9425,N_9464);
and UO_435 (O_435,N_9337,N_8222);
xnor UO_436 (O_436,N_9470,N_9047);
nand UO_437 (O_437,N_8629,N_8655);
nand UO_438 (O_438,N_9100,N_9328);
and UO_439 (O_439,N_8362,N_8140);
or UO_440 (O_440,N_9692,N_9580);
and UO_441 (O_441,N_8850,N_8180);
nand UO_442 (O_442,N_9526,N_9966);
xnor UO_443 (O_443,N_8821,N_9930);
nor UO_444 (O_444,N_9322,N_8298);
nand UO_445 (O_445,N_8186,N_8571);
nand UO_446 (O_446,N_8609,N_9554);
xnor UO_447 (O_447,N_8833,N_9225);
xor UO_448 (O_448,N_8036,N_8084);
or UO_449 (O_449,N_8483,N_8510);
nand UO_450 (O_450,N_9850,N_8659);
and UO_451 (O_451,N_8242,N_9130);
and UO_452 (O_452,N_8473,N_9028);
xor UO_453 (O_453,N_8091,N_8489);
nor UO_454 (O_454,N_8212,N_8211);
and UO_455 (O_455,N_9875,N_9827);
nand UO_456 (O_456,N_8394,N_8898);
and UO_457 (O_457,N_8056,N_8008);
and UO_458 (O_458,N_9848,N_9156);
nor UO_459 (O_459,N_8173,N_8548);
or UO_460 (O_460,N_8178,N_8606);
xnor UO_461 (O_461,N_9230,N_8449);
or UO_462 (O_462,N_9189,N_8003);
nor UO_463 (O_463,N_9896,N_8130);
nor UO_464 (O_464,N_8895,N_9033);
xnor UO_465 (O_465,N_9332,N_9940);
and UO_466 (O_466,N_8818,N_8463);
and UO_467 (O_467,N_8273,N_9114);
or UO_468 (O_468,N_8550,N_9619);
or UO_469 (O_469,N_9678,N_9818);
nor UO_470 (O_470,N_8974,N_8409);
or UO_471 (O_471,N_9249,N_9366);
xor UO_472 (O_472,N_8029,N_8296);
or UO_473 (O_473,N_9275,N_9859);
nor UO_474 (O_474,N_9420,N_8542);
and UO_475 (O_475,N_8790,N_9191);
or UO_476 (O_476,N_8299,N_9529);
and UO_477 (O_477,N_8536,N_9668);
xor UO_478 (O_478,N_8172,N_8585);
xor UO_479 (O_479,N_9095,N_9676);
nand UO_480 (O_480,N_8203,N_8997);
nand UO_481 (O_481,N_8075,N_9442);
and UO_482 (O_482,N_9319,N_9714);
nor UO_483 (O_483,N_9630,N_8424);
or UO_484 (O_484,N_9268,N_8773);
nor UO_485 (O_485,N_8680,N_8406);
and UO_486 (O_486,N_9575,N_8924);
nand UO_487 (O_487,N_9461,N_9040);
and UO_488 (O_488,N_8744,N_9198);
xor UO_489 (O_489,N_9017,N_9298);
nor UO_490 (O_490,N_9229,N_8934);
nand UO_491 (O_491,N_9602,N_8381);
nor UO_492 (O_492,N_9389,N_8357);
and UO_493 (O_493,N_9195,N_9494);
nor UO_494 (O_494,N_9803,N_9825);
xor UO_495 (O_495,N_8722,N_8737);
xor UO_496 (O_496,N_9914,N_9536);
or UO_497 (O_497,N_9412,N_8882);
xnor UO_498 (O_498,N_8505,N_9447);
nor UO_499 (O_499,N_8694,N_8475);
nand UO_500 (O_500,N_9468,N_8302);
nor UO_501 (O_501,N_8848,N_9893);
nor UO_502 (O_502,N_8515,N_9694);
or UO_503 (O_503,N_9638,N_9206);
or UO_504 (O_504,N_8527,N_9806);
nor UO_505 (O_505,N_8582,N_8013);
nand UO_506 (O_506,N_8630,N_9497);
and UO_507 (O_507,N_8041,N_8806);
and UO_508 (O_508,N_8005,N_9500);
and UO_509 (O_509,N_9888,N_8421);
nand UO_510 (O_510,N_9908,N_8956);
nor UO_511 (O_511,N_8504,N_9360);
nand UO_512 (O_512,N_8167,N_9650);
and UO_513 (O_513,N_8518,N_9214);
xnor UO_514 (O_514,N_9307,N_8280);
or UO_515 (O_515,N_9173,N_9533);
nand UO_516 (O_516,N_9272,N_9081);
xor UO_517 (O_517,N_9169,N_8235);
and UO_518 (O_518,N_9699,N_8620);
or UO_519 (O_519,N_8267,N_8427);
or UO_520 (O_520,N_8648,N_8493);
or UO_521 (O_521,N_9796,N_9956);
and UO_522 (O_522,N_8252,N_8596);
and UO_523 (O_523,N_9688,N_9097);
nor UO_524 (O_524,N_9012,N_9539);
and UO_525 (O_525,N_9446,N_9373);
nor UO_526 (O_526,N_9120,N_8471);
nand UO_527 (O_527,N_8725,N_8546);
nand UO_528 (O_528,N_8163,N_9599);
nand UO_529 (O_529,N_8573,N_8327);
xor UO_530 (O_530,N_9976,N_9256);
nand UO_531 (O_531,N_8670,N_8455);
and UO_532 (O_532,N_9624,N_9822);
or UO_533 (O_533,N_9112,N_8965);
xor UO_534 (O_534,N_9920,N_9134);
xor UO_535 (O_535,N_8294,N_8414);
or UO_536 (O_536,N_8369,N_8063);
xor UO_537 (O_537,N_9698,N_9998);
and UO_538 (O_538,N_9146,N_9379);
nor UO_539 (O_539,N_8323,N_8771);
and UO_540 (O_540,N_8862,N_9050);
xnor UO_541 (O_541,N_9199,N_9785);
nand UO_542 (O_542,N_8742,N_8073);
xnor UO_543 (O_543,N_8086,N_9795);
xnor UO_544 (O_544,N_9462,N_8511);
xor UO_545 (O_545,N_8696,N_9484);
or UO_546 (O_546,N_8250,N_8101);
and UO_547 (O_547,N_8125,N_8966);
or UO_548 (O_548,N_9991,N_9323);
xnor UO_549 (O_549,N_9621,N_8704);
and UO_550 (O_550,N_9996,N_9752);
and UO_551 (O_551,N_9938,N_8363);
or UO_552 (O_552,N_9670,N_8784);
nand UO_553 (O_553,N_8495,N_8168);
nand UO_554 (O_554,N_8197,N_9993);
xor UO_555 (O_555,N_8526,N_9960);
nor UO_556 (O_556,N_9610,N_8352);
or UO_557 (O_557,N_8918,N_9400);
nor UO_558 (O_558,N_9919,N_8182);
nor UO_559 (O_559,N_8856,N_8402);
or UO_560 (O_560,N_8064,N_8401);
nor UO_561 (O_561,N_9405,N_9849);
or UO_562 (O_562,N_9368,N_9317);
and UO_563 (O_563,N_9096,N_9789);
and UO_564 (O_564,N_8213,N_9606);
and UO_565 (O_565,N_9150,N_9569);
nand UO_566 (O_566,N_9968,N_9528);
or UO_567 (O_567,N_9473,N_8897);
or UO_568 (O_568,N_9928,N_9576);
and UO_569 (O_569,N_8616,N_9467);
or UO_570 (O_570,N_8451,N_8126);
and UO_571 (O_571,N_8634,N_9439);
xnor UO_572 (O_572,N_9736,N_8581);
nand UO_573 (O_573,N_8456,N_8513);
nand UO_574 (O_574,N_8896,N_8565);
nor UO_575 (O_575,N_9798,N_8686);
xor UO_576 (O_576,N_9243,N_9325);
xnor UO_577 (O_577,N_8491,N_8141);
or UO_578 (O_578,N_8909,N_8448);
or UO_579 (O_579,N_9326,N_8811);
and UO_580 (O_580,N_8237,N_8792);
nand UO_581 (O_581,N_9646,N_9281);
nor UO_582 (O_582,N_9235,N_8509);
nor UO_583 (O_583,N_9303,N_8816);
nand UO_584 (O_584,N_9241,N_9111);
nor UO_585 (O_585,N_8479,N_9637);
or UO_586 (O_586,N_9271,N_8781);
and UO_587 (O_587,N_8103,N_8990);
and UO_588 (O_588,N_8912,N_8187);
or UO_589 (O_589,N_8205,N_8689);
nand UO_590 (O_590,N_8869,N_9737);
and UO_591 (O_591,N_9282,N_8847);
nor UO_592 (O_592,N_8052,N_8817);
or UO_593 (O_593,N_9428,N_9809);
xnor UO_594 (O_594,N_8853,N_9784);
xnor UO_595 (O_595,N_8805,N_8329);
xor UO_596 (O_596,N_8557,N_9330);
nor UO_597 (O_597,N_8104,N_8024);
nor UO_598 (O_598,N_8826,N_8964);
and UO_599 (O_599,N_8476,N_9320);
and UO_600 (O_600,N_8710,N_9496);
nor UO_601 (O_601,N_8674,N_8234);
xor UO_602 (O_602,N_9273,N_9314);
xor UO_603 (O_603,N_9492,N_8941);
xor UO_604 (O_604,N_9555,N_9812);
or UO_605 (O_605,N_9220,N_9525);
and UO_606 (O_606,N_8746,N_8788);
and UO_607 (O_607,N_8721,N_9788);
nand UO_608 (O_608,N_9019,N_8867);
xor UO_609 (O_609,N_9456,N_8277);
and UO_610 (O_610,N_9680,N_9759);
and UO_611 (O_611,N_8700,N_8116);
xor UO_612 (O_612,N_8612,N_9459);
nand UO_613 (O_613,N_8525,N_9725);
nand UO_614 (O_614,N_8272,N_9604);
or UO_615 (O_615,N_9618,N_9810);
nand UO_616 (O_616,N_9702,N_8960);
and UO_617 (O_617,N_9122,N_8947);
or UO_618 (O_618,N_8106,N_9232);
nand UO_619 (O_619,N_9828,N_8258);
or UO_620 (O_620,N_8884,N_8537);
and UO_621 (O_621,N_8240,N_8376);
nand UO_622 (O_622,N_8980,N_9544);
or UO_623 (O_623,N_8166,N_9424);
xor UO_624 (O_624,N_9710,N_9614);
nor UO_625 (O_625,N_8921,N_9588);
and UO_626 (O_626,N_9675,N_9094);
and UO_627 (O_627,N_8202,N_9832);
nand UO_628 (O_628,N_9078,N_8468);
or UO_629 (O_629,N_9900,N_9003);
nand UO_630 (O_630,N_8830,N_8507);
nand UO_631 (O_631,N_9109,N_9215);
and UO_632 (O_632,N_8452,N_8458);
nor UO_633 (O_633,N_9421,N_8860);
and UO_634 (O_634,N_8823,N_9158);
and UO_635 (O_635,N_9876,N_9906);
nand UO_636 (O_636,N_8637,N_9277);
xnor UO_637 (O_637,N_9503,N_8085);
xor UO_638 (O_638,N_9186,N_9664);
nor UO_639 (O_639,N_8002,N_8322);
or UO_640 (O_640,N_9265,N_9126);
and UO_641 (O_641,N_9518,N_8392);
or UO_642 (O_642,N_8543,N_9077);
or UO_643 (O_643,N_9088,N_8937);
nand UO_644 (O_644,N_9983,N_9027);
xor UO_645 (O_645,N_9072,N_9025);
xnor UO_646 (O_646,N_8014,N_9163);
xnor UO_647 (O_647,N_8026,N_9139);
and UO_648 (O_648,N_8814,N_9743);
xnor UO_649 (O_649,N_9076,N_9438);
nor UO_650 (O_650,N_8775,N_9715);
nor UO_651 (O_651,N_9907,N_9708);
and UO_652 (O_652,N_9233,N_9159);
xnor UO_653 (O_653,N_8644,N_8926);
or UO_654 (O_654,N_9172,N_8649);
and UO_655 (O_655,N_9394,N_8433);
nand UO_656 (O_656,N_9712,N_8236);
or UO_657 (O_657,N_9364,N_8134);
and UO_658 (O_658,N_8705,N_8397);
nor UO_659 (O_659,N_8554,N_9513);
or UO_660 (O_660,N_8338,N_9773);
nand UO_661 (O_661,N_8758,N_9251);
xnor UO_662 (O_662,N_9511,N_9207);
or UO_663 (O_663,N_9427,N_9083);
or UO_664 (O_664,N_9577,N_8233);
or UO_665 (O_665,N_8736,N_8959);
nor UO_666 (O_666,N_8608,N_9043);
nand UO_667 (O_667,N_9200,N_9992);
xor UO_668 (O_668,N_8813,N_8673);
and UO_669 (O_669,N_8892,N_8671);
or UO_670 (O_670,N_8342,N_8446);
nor UO_671 (O_671,N_8719,N_9182);
xor UO_672 (O_672,N_8154,N_8034);
and UO_673 (O_673,N_8100,N_8079);
nor UO_674 (O_674,N_8070,N_9596);
or UO_675 (O_675,N_9289,N_8083);
nor UO_676 (O_676,N_9292,N_9965);
nand UO_677 (O_677,N_8477,N_8441);
or UO_678 (O_678,N_8383,N_9753);
xnor UO_679 (O_679,N_8048,N_8499);
or UO_680 (O_680,N_9884,N_9622);
xnor UO_681 (O_681,N_8782,N_8545);
nand UO_682 (O_682,N_8078,N_9672);
xnor UO_683 (O_683,N_9548,N_9830);
nor UO_684 (O_684,N_9274,N_8384);
nand UO_685 (O_685,N_8605,N_8259);
nor UO_686 (O_686,N_9343,N_8954);
or UO_687 (O_687,N_9589,N_9551);
nand UO_688 (O_688,N_9524,N_9013);
xor UO_689 (O_689,N_9959,N_9530);
xor UO_690 (O_690,N_9926,N_9639);
or UO_691 (O_691,N_9301,N_9866);
nor UO_692 (O_692,N_8706,N_8364);
and UO_693 (O_693,N_9717,N_8361);
xor UO_694 (O_694,N_9166,N_8037);
or UO_695 (O_695,N_8017,N_9239);
nor UO_696 (O_696,N_9709,N_8132);
or UO_697 (O_697,N_9740,N_8872);
xor UO_698 (O_698,N_9351,N_9149);
or UO_699 (O_699,N_8313,N_8356);
and UO_700 (O_700,N_8994,N_8650);
nor UO_701 (O_701,N_8717,N_9658);
xor UO_702 (O_702,N_8439,N_8231);
or UO_703 (O_703,N_9553,N_9066);
or UO_704 (O_704,N_8873,N_9118);
xor UO_705 (O_705,N_9392,N_9136);
xor UO_706 (O_706,N_8945,N_8793);
or UO_707 (O_707,N_9732,N_8358);
nor UO_708 (O_708,N_8307,N_8570);
and UO_709 (O_709,N_8764,N_8870);
nor UO_710 (O_710,N_8123,N_9517);
and UO_711 (O_711,N_8247,N_8588);
or UO_712 (O_712,N_8375,N_8743);
or UO_713 (O_713,N_8591,N_8800);
nor UO_714 (O_714,N_8999,N_8866);
nor UO_715 (O_715,N_8054,N_9921);
nand UO_716 (O_716,N_8270,N_9006);
or UO_717 (O_717,N_8685,N_8549);
or UO_718 (O_718,N_8520,N_8578);
and UO_719 (O_719,N_9601,N_9353);
nor UO_720 (O_720,N_9643,N_9590);
or UO_721 (O_721,N_8263,N_8096);
xor UO_722 (O_722,N_8418,N_9979);
xor UO_723 (O_723,N_8147,N_8337);
and UO_724 (O_724,N_9506,N_9797);
or UO_725 (O_725,N_9007,N_8530);
nor UO_726 (O_726,N_8081,N_9815);
nand UO_727 (O_727,N_8708,N_8373);
nand UO_728 (O_728,N_8387,N_8948);
and UO_729 (O_729,N_9127,N_8677);
or UO_730 (O_730,N_9661,N_9259);
and UO_731 (O_731,N_9583,N_9800);
or UO_732 (O_732,N_9450,N_8951);
nor UO_733 (O_733,N_8636,N_9370);
nor UO_734 (O_734,N_9943,N_8391);
or UO_735 (O_735,N_9934,N_9776);
and UO_736 (O_736,N_8640,N_8993);
and UO_737 (O_737,N_8885,N_8604);
nand UO_738 (O_738,N_8734,N_8435);
nor UO_739 (O_739,N_8852,N_8988);
nor UO_740 (O_740,N_8454,N_8265);
and UO_741 (O_741,N_8828,N_9165);
nand UO_742 (O_742,N_8122,N_8992);
or UO_743 (O_743,N_8150,N_8646);
or UO_744 (O_744,N_8711,N_8827);
nor UO_745 (O_745,N_9840,N_8568);
xor UO_746 (O_746,N_8494,N_9665);
xnor UO_747 (O_747,N_9349,N_9846);
xnor UO_748 (O_748,N_9775,N_9080);
xnor UO_749 (O_749,N_9108,N_8556);
and UO_750 (O_750,N_9869,N_8388);
nand UO_751 (O_751,N_8068,N_8906);
or UO_752 (O_752,N_8789,N_9133);
nand UO_753 (O_753,N_8791,N_9820);
xor UO_754 (O_754,N_9437,N_8593);
and UO_755 (O_755,N_8695,N_8474);
or UO_756 (O_756,N_8035,N_9994);
nor UO_757 (O_757,N_8128,N_9508);
nor UO_758 (O_758,N_8137,N_8820);
and UO_759 (O_759,N_9409,N_8185);
or UO_760 (O_760,N_8584,N_8297);
xnor UO_761 (O_761,N_8241,N_8726);
xor UO_762 (O_762,N_8049,N_8932);
xor UO_763 (O_763,N_9236,N_8318);
xor UO_764 (O_764,N_8412,N_9816);
xnor UO_765 (O_765,N_9592,N_9995);
nand UO_766 (O_766,N_9681,N_8038);
or UO_767 (O_767,N_9739,N_8050);
xnor UO_768 (O_768,N_8669,N_8360);
nand UO_769 (O_769,N_9579,N_8950);
or UO_770 (O_770,N_9641,N_9671);
nand UO_771 (O_771,N_8472,N_9719);
xor UO_772 (O_772,N_9339,N_8503);
nand UO_773 (O_773,N_9049,N_8889);
or UO_774 (O_774,N_9104,N_9283);
nor UO_775 (O_775,N_9686,N_9286);
nand UO_776 (O_776,N_9763,N_8260);
nor UO_777 (O_777,N_9110,N_8136);
and UO_778 (O_778,N_8195,N_9082);
nor UO_779 (O_779,N_9250,N_9344);
and UO_780 (O_780,N_8365,N_9210);
nor UO_781 (O_781,N_8540,N_8057);
nor UO_782 (O_782,N_9857,N_9227);
nor UO_783 (O_783,N_9823,N_8607);
or UO_784 (O_784,N_8940,N_8765);
xor UO_785 (O_785,N_9415,N_8127);
or UO_786 (O_786,N_9222,N_8983);
and UO_787 (O_787,N_9559,N_9835);
xor UO_788 (O_788,N_9705,N_8931);
nand UO_789 (O_789,N_9690,N_8249);
nand UO_790 (O_790,N_8521,N_8728);
or UO_791 (O_791,N_9460,N_9391);
nand UO_792 (O_792,N_8131,N_9458);
and UO_793 (O_793,N_8660,N_9963);
or UO_794 (O_794,N_8933,N_9477);
nand UO_795 (O_795,N_8028,N_8444);
or UO_796 (O_796,N_8011,N_9213);
nor UO_797 (O_797,N_8042,N_9041);
and UO_798 (O_798,N_9457,N_9411);
nor UO_799 (O_799,N_8987,N_8733);
xnor UO_800 (O_800,N_9616,N_8780);
nor UO_801 (O_801,N_8230,N_9964);
xor UO_802 (O_802,N_8851,N_8888);
nand UO_803 (O_803,N_8583,N_8732);
xor UO_804 (O_804,N_8194,N_8061);
xor UO_805 (O_805,N_9769,N_9978);
nand UO_806 (O_806,N_8450,N_9084);
nor UO_807 (O_807,N_9674,N_8099);
xor UO_808 (O_808,N_9758,N_9704);
xnor UO_809 (O_809,N_8315,N_8366);
and UO_810 (O_810,N_9046,N_8415);
and UO_811 (O_811,N_9584,N_9128);
and UO_812 (O_812,N_9700,N_8312);
and UO_813 (O_813,N_8158,N_8227);
nand UO_814 (O_814,N_8621,N_8907);
nand UO_815 (O_815,N_8769,N_9600);
nor UO_816 (O_816,N_9749,N_9557);
or UO_817 (O_817,N_8438,N_9826);
nand UO_818 (O_818,N_9435,N_8972);
nand UO_819 (O_819,N_9862,N_8855);
nand UO_820 (O_820,N_9075,N_9633);
nand UO_821 (O_821,N_9787,N_8047);
nand UO_822 (O_822,N_9125,N_8176);
xor UO_823 (O_823,N_8492,N_9479);
and UO_824 (O_824,N_9396,N_8797);
nand UO_825 (O_825,N_9016,N_9974);
or UO_826 (O_826,N_8961,N_8191);
nand UO_827 (O_827,N_9612,N_9101);
xnor UO_828 (O_828,N_8641,N_8750);
or UO_829 (O_829,N_9406,N_9726);
or UO_830 (O_830,N_8465,N_8088);
and UO_831 (O_831,N_9997,N_8938);
nor UO_832 (O_832,N_8359,N_9521);
or UO_833 (O_833,N_8160,N_9454);
xnor UO_834 (O_834,N_9399,N_8857);
or UO_835 (O_835,N_9947,N_9022);
or UO_836 (O_836,N_9099,N_9318);
and UO_837 (O_837,N_9407,N_9711);
nand UO_838 (O_838,N_9002,N_9443);
or UO_839 (O_839,N_8762,N_9898);
nor UO_840 (O_840,N_8981,N_8925);
or UO_841 (O_841,N_8701,N_9218);
or UO_842 (O_842,N_8877,N_8533);
or UO_843 (O_843,N_9264,N_9255);
nand UO_844 (O_844,N_8348,N_8419);
nand UO_845 (O_845,N_9291,N_8114);
or UO_846 (O_846,N_8040,N_8534);
and UO_847 (O_847,N_8904,N_8522);
and UO_848 (O_848,N_9501,N_9607);
xnor UO_849 (O_849,N_8021,N_9718);
nor UO_850 (O_850,N_8058,N_9510);
nand UO_851 (O_851,N_9168,N_9401);
nor UO_852 (O_852,N_9932,N_9860);
or UO_853 (O_853,N_8712,N_8840);
nor UO_854 (O_854,N_9852,N_9098);
and UO_855 (O_855,N_9060,N_8825);
nor UO_856 (O_856,N_9029,N_8377);
and UO_857 (O_857,N_8326,N_9504);
nor UO_858 (O_858,N_9148,N_9882);
xnor UO_859 (O_859,N_9157,N_8416);
nand UO_860 (O_860,N_8720,N_9924);
nor UO_861 (O_861,N_9352,N_9354);
nor UO_862 (O_862,N_9863,N_9573);
nor UO_863 (O_863,N_8772,N_8803);
nor UO_864 (O_864,N_8654,N_9297);
xor UO_865 (O_865,N_8224,N_8647);
nand UO_866 (O_866,N_8555,N_9952);
and UO_867 (O_867,N_9541,N_8355);
nor UO_868 (O_868,N_9552,N_8958);
or UO_869 (O_869,N_8253,N_8399);
and UO_870 (O_870,N_9617,N_9656);
and UO_871 (O_871,N_9640,N_8566);
nor UO_872 (O_872,N_9061,N_9765);
or UO_873 (O_873,N_9540,N_9248);
nand UO_874 (O_874,N_8679,N_8519);
nand UO_875 (O_875,N_9696,N_8564);
or UO_876 (O_876,N_8244,N_9945);
and UO_877 (O_877,N_9562,N_9790);
nor UO_878 (O_878,N_8417,N_8469);
and UO_879 (O_879,N_9969,N_8311);
or UO_880 (O_880,N_8651,N_8155);
nand UO_881 (O_881,N_8289,N_8389);
nor UO_882 (O_882,N_9534,N_9677);
nand UO_883 (O_883,N_9187,N_9942);
nand UO_884 (O_884,N_8558,N_9015);
nand UO_885 (O_885,N_8379,N_8969);
nor UO_886 (O_886,N_9877,N_8514);
or UO_887 (O_887,N_9123,N_9423);
and UO_888 (O_888,N_9246,N_9701);
nand UO_889 (O_889,N_9721,N_8204);
or UO_890 (O_890,N_8330,N_8229);
or UO_891 (O_891,N_9730,N_8723);
nand UO_892 (O_892,N_8245,N_9847);
nor UO_893 (O_893,N_8023,N_9475);
xnor UO_894 (O_894,N_8500,N_8169);
nor UO_895 (O_895,N_8341,N_9348);
and UO_896 (O_896,N_8716,N_9135);
xnor UO_897 (O_897,N_8152,N_8382);
nand UO_898 (O_898,N_8597,N_8779);
or UO_899 (O_899,N_9543,N_8380);
nand UO_900 (O_900,N_9070,N_9564);
nor UO_901 (O_901,N_9321,N_9817);
nor UO_902 (O_902,N_9487,N_8110);
nor UO_903 (O_903,N_9223,N_8309);
nand UO_904 (O_904,N_8216,N_9957);
nand UO_905 (O_905,N_9669,N_9261);
nand UO_906 (O_906,N_9768,N_8189);
nand UO_907 (O_907,N_9858,N_9546);
nand UO_908 (O_908,N_8576,N_8310);
xor UO_909 (O_909,N_8893,N_9231);
xor UO_910 (O_910,N_8436,N_8033);
nand UO_911 (O_911,N_9316,N_9917);
and UO_912 (O_912,N_8613,N_9813);
nand UO_913 (O_913,N_8626,N_8776);
nor UO_914 (O_914,N_9778,N_8579);
xor UO_915 (O_915,N_8767,N_8761);
and UO_916 (O_916,N_9586,N_8598);
xnor UO_917 (O_917,N_9285,N_8112);
nor UO_918 (O_918,N_9300,N_8308);
nand UO_919 (O_919,N_9999,N_9767);
nor UO_920 (O_920,N_8287,N_8552);
and UO_921 (O_921,N_8986,N_9545);
nand UO_922 (O_922,N_8074,N_9901);
nand UO_923 (O_923,N_9336,N_9342);
xnor UO_924 (O_924,N_9445,N_8159);
and UO_925 (O_925,N_9287,N_8149);
or UO_926 (O_926,N_8920,N_9151);
and UO_927 (O_927,N_8223,N_8065);
and UO_928 (O_928,N_9481,N_8423);
nand UO_929 (O_929,N_8133,N_9294);
nor UO_930 (O_930,N_9179,N_9102);
nand UO_931 (O_931,N_9372,N_8434);
nor UO_932 (O_932,N_9334,N_9308);
nor UO_933 (O_933,N_8599,N_8214);
nand UO_934 (O_934,N_8787,N_8488);
nand UO_935 (O_935,N_9410,N_9288);
nor UO_936 (O_936,N_8317,N_9381);
nand UO_937 (O_937,N_9005,N_9748);
nor UO_938 (O_938,N_9937,N_9045);
nand UO_939 (O_939,N_8464,N_9115);
and UO_940 (O_940,N_8590,N_9879);
xor UO_941 (O_941,N_8470,N_9620);
or UO_942 (O_942,N_8278,N_9911);
nand UO_943 (O_943,N_9147,N_8622);
xor UO_944 (O_944,N_9180,N_9197);
xor UO_945 (O_945,N_8807,N_9949);
and UO_946 (O_946,N_8977,N_9279);
nor UO_947 (O_947,N_8306,N_8713);
xor UO_948 (O_948,N_8891,N_9779);
and UO_949 (O_949,N_9838,N_9258);
xnor UO_950 (O_950,N_9175,N_9201);
nor UO_951 (O_951,N_8875,N_8879);
and UO_952 (O_952,N_9422,N_8467);
nor UO_953 (O_953,N_9141,N_9625);
xor UO_954 (O_954,N_8672,N_9455);
nand UO_955 (O_955,N_8683,N_8831);
and UO_956 (O_956,N_9512,N_8039);
or UO_957 (O_957,N_8239,N_9780);
and UO_958 (O_958,N_9212,N_9522);
or UO_959 (O_959,N_8798,N_8574);
nand UO_960 (O_960,N_9883,N_9895);
or UO_961 (O_961,N_8899,N_8928);
nor UO_962 (O_962,N_9735,N_9065);
or UO_963 (O_963,N_9958,N_9757);
and UO_964 (O_964,N_9374,N_8741);
or UO_965 (O_965,N_9362,N_8164);
or UO_966 (O_966,N_9452,N_8179);
nor UO_967 (O_967,N_9202,N_9682);
nand UO_968 (O_968,N_9242,N_9001);
nor UO_969 (O_969,N_8715,N_8842);
and UO_970 (O_970,N_9685,N_8016);
xnor UO_971 (O_971,N_8914,N_9892);
nor UO_972 (O_972,N_8386,N_9903);
nand UO_973 (O_973,N_8760,N_8998);
nand UO_974 (O_974,N_9868,N_9989);
nand UO_975 (O_975,N_8283,N_9939);
or UO_976 (O_976,N_8210,N_8238);
nor UO_977 (O_977,N_8333,N_8209);
or UO_978 (O_978,N_8569,N_8346);
nor UO_979 (O_979,N_8066,N_9741);
xor UO_980 (O_980,N_8295,N_8812);
nor UO_981 (O_981,N_9356,N_8832);
or UO_982 (O_982,N_9413,N_8615);
or UO_983 (O_983,N_9009,N_9221);
nand UO_984 (O_984,N_8774,N_9889);
nand UO_985 (O_985,N_8344,N_9756);
and UO_986 (O_986,N_8069,N_8395);
xor UO_987 (O_987,N_9897,N_8824);
xor UO_988 (O_988,N_8844,N_8661);
and UO_989 (O_989,N_9418,N_9489);
xnor UO_990 (O_990,N_9471,N_8293);
xor UO_991 (O_991,N_9035,N_9419);
nor UO_992 (O_992,N_9058,N_9026);
nand UO_993 (O_993,N_8367,N_9693);
xnor UO_994 (O_994,N_9217,N_9973);
nor UO_995 (O_995,N_9178,N_9252);
nor UO_996 (O_996,N_9988,N_9587);
and UO_997 (O_997,N_9495,N_9771);
or UO_998 (O_998,N_8559,N_9936);
nor UO_999 (O_999,N_9408,N_9044);
xor UO_1000 (O_1000,N_8676,N_9724);
and UO_1001 (O_1001,N_9017,N_8556);
xor UO_1002 (O_1002,N_8550,N_8881);
nor UO_1003 (O_1003,N_9629,N_8365);
nand UO_1004 (O_1004,N_8749,N_9255);
or UO_1005 (O_1005,N_8604,N_9771);
nor UO_1006 (O_1006,N_8339,N_8142);
nand UO_1007 (O_1007,N_9113,N_9443);
nor UO_1008 (O_1008,N_9613,N_9373);
and UO_1009 (O_1009,N_8089,N_9840);
nor UO_1010 (O_1010,N_8485,N_9513);
nor UO_1011 (O_1011,N_8836,N_8597);
xnor UO_1012 (O_1012,N_9744,N_9985);
nor UO_1013 (O_1013,N_9836,N_9154);
xor UO_1014 (O_1014,N_9501,N_9916);
or UO_1015 (O_1015,N_8186,N_9948);
xor UO_1016 (O_1016,N_8567,N_8762);
or UO_1017 (O_1017,N_9720,N_8543);
or UO_1018 (O_1018,N_8980,N_8996);
and UO_1019 (O_1019,N_9916,N_9558);
and UO_1020 (O_1020,N_9193,N_8749);
or UO_1021 (O_1021,N_9064,N_9813);
xor UO_1022 (O_1022,N_8546,N_8876);
xor UO_1023 (O_1023,N_8585,N_9706);
xnor UO_1024 (O_1024,N_9975,N_8959);
xnor UO_1025 (O_1025,N_9941,N_8112);
nand UO_1026 (O_1026,N_9741,N_8223);
xor UO_1027 (O_1027,N_9813,N_9723);
nand UO_1028 (O_1028,N_9269,N_9102);
or UO_1029 (O_1029,N_8735,N_9897);
xnor UO_1030 (O_1030,N_8440,N_8695);
nor UO_1031 (O_1031,N_8585,N_8550);
or UO_1032 (O_1032,N_8797,N_9947);
or UO_1033 (O_1033,N_9670,N_9931);
nand UO_1034 (O_1034,N_9158,N_9340);
xor UO_1035 (O_1035,N_8308,N_9746);
nand UO_1036 (O_1036,N_8139,N_9897);
xor UO_1037 (O_1037,N_8639,N_9367);
nor UO_1038 (O_1038,N_9978,N_8368);
nand UO_1039 (O_1039,N_9795,N_9883);
nor UO_1040 (O_1040,N_8791,N_8611);
xor UO_1041 (O_1041,N_9680,N_9026);
nor UO_1042 (O_1042,N_8196,N_8601);
xnor UO_1043 (O_1043,N_9395,N_8786);
xor UO_1044 (O_1044,N_8627,N_8619);
xor UO_1045 (O_1045,N_8614,N_9617);
xnor UO_1046 (O_1046,N_9129,N_9325);
or UO_1047 (O_1047,N_8350,N_8210);
xnor UO_1048 (O_1048,N_9755,N_8680);
or UO_1049 (O_1049,N_8536,N_9570);
xor UO_1050 (O_1050,N_9411,N_9260);
nor UO_1051 (O_1051,N_8416,N_9053);
xnor UO_1052 (O_1052,N_9023,N_9692);
nand UO_1053 (O_1053,N_9108,N_9566);
or UO_1054 (O_1054,N_9202,N_9100);
and UO_1055 (O_1055,N_8746,N_9502);
nor UO_1056 (O_1056,N_8421,N_9598);
nand UO_1057 (O_1057,N_8625,N_9022);
xor UO_1058 (O_1058,N_9048,N_9437);
xor UO_1059 (O_1059,N_9055,N_9385);
or UO_1060 (O_1060,N_8467,N_9418);
and UO_1061 (O_1061,N_9222,N_8804);
and UO_1062 (O_1062,N_9766,N_9869);
xor UO_1063 (O_1063,N_9819,N_8234);
and UO_1064 (O_1064,N_8439,N_8838);
nor UO_1065 (O_1065,N_9712,N_9375);
xor UO_1066 (O_1066,N_9085,N_8327);
xnor UO_1067 (O_1067,N_9088,N_9129);
and UO_1068 (O_1068,N_8169,N_9414);
nand UO_1069 (O_1069,N_9034,N_9916);
or UO_1070 (O_1070,N_8055,N_8648);
and UO_1071 (O_1071,N_8308,N_8919);
and UO_1072 (O_1072,N_8988,N_8100);
and UO_1073 (O_1073,N_9857,N_9443);
xnor UO_1074 (O_1074,N_9858,N_9209);
and UO_1075 (O_1075,N_9340,N_9461);
or UO_1076 (O_1076,N_8076,N_8678);
nand UO_1077 (O_1077,N_8228,N_8598);
nand UO_1078 (O_1078,N_9647,N_9113);
xnor UO_1079 (O_1079,N_9225,N_8913);
xor UO_1080 (O_1080,N_8129,N_8815);
nor UO_1081 (O_1081,N_8088,N_9467);
xor UO_1082 (O_1082,N_8801,N_8241);
or UO_1083 (O_1083,N_8161,N_8981);
xor UO_1084 (O_1084,N_9968,N_9350);
nor UO_1085 (O_1085,N_8397,N_9124);
and UO_1086 (O_1086,N_9371,N_8321);
or UO_1087 (O_1087,N_8709,N_8643);
and UO_1088 (O_1088,N_8091,N_8058);
nand UO_1089 (O_1089,N_8804,N_8054);
nor UO_1090 (O_1090,N_8859,N_9324);
xor UO_1091 (O_1091,N_8308,N_8157);
nand UO_1092 (O_1092,N_8456,N_8963);
nand UO_1093 (O_1093,N_8514,N_8325);
and UO_1094 (O_1094,N_9187,N_9911);
or UO_1095 (O_1095,N_8252,N_9218);
or UO_1096 (O_1096,N_8234,N_9443);
nand UO_1097 (O_1097,N_9847,N_8448);
xor UO_1098 (O_1098,N_8340,N_8898);
or UO_1099 (O_1099,N_8558,N_8406);
xor UO_1100 (O_1100,N_8450,N_9136);
nand UO_1101 (O_1101,N_8649,N_8642);
and UO_1102 (O_1102,N_8717,N_9270);
nand UO_1103 (O_1103,N_8836,N_8765);
xnor UO_1104 (O_1104,N_8078,N_8322);
xnor UO_1105 (O_1105,N_8113,N_8357);
xor UO_1106 (O_1106,N_9323,N_9741);
nand UO_1107 (O_1107,N_8460,N_9077);
xor UO_1108 (O_1108,N_9750,N_8538);
nand UO_1109 (O_1109,N_9639,N_8022);
nor UO_1110 (O_1110,N_9946,N_8849);
nor UO_1111 (O_1111,N_8103,N_9715);
nor UO_1112 (O_1112,N_9444,N_9699);
and UO_1113 (O_1113,N_9718,N_8188);
nor UO_1114 (O_1114,N_9884,N_8632);
xor UO_1115 (O_1115,N_8237,N_9251);
and UO_1116 (O_1116,N_8110,N_9281);
and UO_1117 (O_1117,N_9465,N_9162);
nand UO_1118 (O_1118,N_9681,N_8506);
xor UO_1119 (O_1119,N_9115,N_9503);
nor UO_1120 (O_1120,N_9880,N_9710);
nor UO_1121 (O_1121,N_9877,N_8031);
or UO_1122 (O_1122,N_8284,N_9128);
nor UO_1123 (O_1123,N_8163,N_8925);
nand UO_1124 (O_1124,N_8489,N_8724);
nor UO_1125 (O_1125,N_9591,N_8935);
and UO_1126 (O_1126,N_8163,N_9021);
and UO_1127 (O_1127,N_9585,N_8769);
nand UO_1128 (O_1128,N_9576,N_8026);
and UO_1129 (O_1129,N_8049,N_8830);
nor UO_1130 (O_1130,N_9951,N_8550);
and UO_1131 (O_1131,N_8922,N_9321);
xnor UO_1132 (O_1132,N_9085,N_8637);
nor UO_1133 (O_1133,N_9264,N_9052);
and UO_1134 (O_1134,N_9200,N_9555);
nor UO_1135 (O_1135,N_9977,N_9910);
nor UO_1136 (O_1136,N_8333,N_8672);
and UO_1137 (O_1137,N_9591,N_8725);
or UO_1138 (O_1138,N_8610,N_9283);
and UO_1139 (O_1139,N_8543,N_9580);
nand UO_1140 (O_1140,N_8592,N_9518);
xor UO_1141 (O_1141,N_9913,N_9105);
or UO_1142 (O_1142,N_8973,N_8090);
xnor UO_1143 (O_1143,N_8279,N_9640);
or UO_1144 (O_1144,N_8692,N_8567);
and UO_1145 (O_1145,N_8458,N_9610);
and UO_1146 (O_1146,N_8607,N_8858);
nor UO_1147 (O_1147,N_8945,N_8084);
nor UO_1148 (O_1148,N_9953,N_8339);
and UO_1149 (O_1149,N_9711,N_9707);
and UO_1150 (O_1150,N_9477,N_8194);
nor UO_1151 (O_1151,N_8371,N_9052);
and UO_1152 (O_1152,N_9852,N_8251);
xor UO_1153 (O_1153,N_9515,N_8718);
xnor UO_1154 (O_1154,N_8519,N_8332);
nor UO_1155 (O_1155,N_8357,N_9665);
and UO_1156 (O_1156,N_9279,N_8845);
and UO_1157 (O_1157,N_9970,N_9094);
or UO_1158 (O_1158,N_9924,N_9651);
nand UO_1159 (O_1159,N_9861,N_8053);
xnor UO_1160 (O_1160,N_8508,N_8418);
xor UO_1161 (O_1161,N_9614,N_8303);
nor UO_1162 (O_1162,N_8391,N_9297);
xnor UO_1163 (O_1163,N_8247,N_8577);
and UO_1164 (O_1164,N_8260,N_8995);
and UO_1165 (O_1165,N_9874,N_9033);
and UO_1166 (O_1166,N_8434,N_9154);
or UO_1167 (O_1167,N_9810,N_8230);
and UO_1168 (O_1168,N_8993,N_9967);
nand UO_1169 (O_1169,N_8091,N_9652);
xor UO_1170 (O_1170,N_8983,N_8964);
or UO_1171 (O_1171,N_8640,N_9337);
xor UO_1172 (O_1172,N_8534,N_9502);
nor UO_1173 (O_1173,N_9938,N_8214);
and UO_1174 (O_1174,N_9055,N_8376);
nor UO_1175 (O_1175,N_8693,N_8907);
or UO_1176 (O_1176,N_8363,N_9902);
xnor UO_1177 (O_1177,N_9088,N_8939);
nand UO_1178 (O_1178,N_9254,N_9058);
nand UO_1179 (O_1179,N_9125,N_8652);
xnor UO_1180 (O_1180,N_9478,N_8311);
xor UO_1181 (O_1181,N_9479,N_8080);
and UO_1182 (O_1182,N_8518,N_8286);
xnor UO_1183 (O_1183,N_9554,N_9332);
and UO_1184 (O_1184,N_8603,N_8492);
and UO_1185 (O_1185,N_8831,N_9302);
xnor UO_1186 (O_1186,N_8284,N_9365);
xor UO_1187 (O_1187,N_9610,N_9042);
nor UO_1188 (O_1188,N_9034,N_8021);
and UO_1189 (O_1189,N_9615,N_8115);
xor UO_1190 (O_1190,N_8785,N_9111);
xnor UO_1191 (O_1191,N_8587,N_9308);
nand UO_1192 (O_1192,N_8473,N_9511);
nand UO_1193 (O_1193,N_9381,N_8158);
nand UO_1194 (O_1194,N_9799,N_9727);
nor UO_1195 (O_1195,N_8023,N_8535);
nand UO_1196 (O_1196,N_9303,N_9525);
and UO_1197 (O_1197,N_8459,N_9028);
nand UO_1198 (O_1198,N_9370,N_8656);
or UO_1199 (O_1199,N_8532,N_9502);
xnor UO_1200 (O_1200,N_8272,N_9722);
xor UO_1201 (O_1201,N_8226,N_8553);
and UO_1202 (O_1202,N_9876,N_9898);
nand UO_1203 (O_1203,N_8869,N_8372);
or UO_1204 (O_1204,N_8177,N_8319);
and UO_1205 (O_1205,N_9654,N_9685);
and UO_1206 (O_1206,N_9554,N_9970);
xnor UO_1207 (O_1207,N_8252,N_8743);
xor UO_1208 (O_1208,N_8898,N_9949);
or UO_1209 (O_1209,N_9966,N_9666);
or UO_1210 (O_1210,N_9390,N_8341);
or UO_1211 (O_1211,N_9862,N_8897);
and UO_1212 (O_1212,N_9116,N_9491);
or UO_1213 (O_1213,N_9309,N_9069);
nand UO_1214 (O_1214,N_9905,N_8061);
nand UO_1215 (O_1215,N_8155,N_9749);
nor UO_1216 (O_1216,N_8333,N_8215);
or UO_1217 (O_1217,N_8623,N_9842);
nand UO_1218 (O_1218,N_9928,N_8443);
or UO_1219 (O_1219,N_8975,N_9623);
and UO_1220 (O_1220,N_8617,N_9289);
xnor UO_1221 (O_1221,N_9051,N_8569);
nand UO_1222 (O_1222,N_9051,N_9207);
and UO_1223 (O_1223,N_9754,N_9100);
nand UO_1224 (O_1224,N_9313,N_9064);
xor UO_1225 (O_1225,N_9522,N_9142);
nor UO_1226 (O_1226,N_8451,N_8749);
nand UO_1227 (O_1227,N_8698,N_9055);
xnor UO_1228 (O_1228,N_9406,N_9287);
nand UO_1229 (O_1229,N_9952,N_9936);
nor UO_1230 (O_1230,N_8563,N_8775);
nand UO_1231 (O_1231,N_8644,N_8758);
nor UO_1232 (O_1232,N_9980,N_9620);
nor UO_1233 (O_1233,N_8273,N_8757);
and UO_1234 (O_1234,N_9497,N_9878);
xor UO_1235 (O_1235,N_8026,N_9317);
or UO_1236 (O_1236,N_9928,N_8666);
nor UO_1237 (O_1237,N_9075,N_8797);
or UO_1238 (O_1238,N_9445,N_8552);
nand UO_1239 (O_1239,N_8291,N_8774);
nor UO_1240 (O_1240,N_8242,N_9342);
or UO_1241 (O_1241,N_8965,N_9446);
nand UO_1242 (O_1242,N_8662,N_9223);
and UO_1243 (O_1243,N_9513,N_9480);
xnor UO_1244 (O_1244,N_9604,N_8265);
xor UO_1245 (O_1245,N_8105,N_9273);
or UO_1246 (O_1246,N_8853,N_9316);
xnor UO_1247 (O_1247,N_8428,N_8352);
and UO_1248 (O_1248,N_9100,N_9358);
or UO_1249 (O_1249,N_8435,N_8582);
xor UO_1250 (O_1250,N_8180,N_8896);
nor UO_1251 (O_1251,N_8799,N_9820);
xnor UO_1252 (O_1252,N_8418,N_9670);
nor UO_1253 (O_1253,N_9097,N_8415);
xor UO_1254 (O_1254,N_9314,N_8963);
and UO_1255 (O_1255,N_8706,N_8026);
nor UO_1256 (O_1256,N_9875,N_9951);
and UO_1257 (O_1257,N_9289,N_9015);
and UO_1258 (O_1258,N_9694,N_8200);
nand UO_1259 (O_1259,N_8966,N_9584);
nor UO_1260 (O_1260,N_8219,N_8101);
nor UO_1261 (O_1261,N_9638,N_9142);
xnor UO_1262 (O_1262,N_8993,N_9858);
and UO_1263 (O_1263,N_9370,N_9618);
xnor UO_1264 (O_1264,N_8173,N_9509);
and UO_1265 (O_1265,N_8970,N_8872);
xor UO_1266 (O_1266,N_8170,N_9510);
or UO_1267 (O_1267,N_9680,N_9989);
nor UO_1268 (O_1268,N_8084,N_8425);
or UO_1269 (O_1269,N_8520,N_8641);
nand UO_1270 (O_1270,N_8514,N_9072);
and UO_1271 (O_1271,N_9343,N_8209);
and UO_1272 (O_1272,N_8870,N_8733);
xor UO_1273 (O_1273,N_8474,N_8997);
xor UO_1274 (O_1274,N_8406,N_8217);
nand UO_1275 (O_1275,N_9820,N_8994);
nand UO_1276 (O_1276,N_8609,N_9126);
nor UO_1277 (O_1277,N_9118,N_9435);
or UO_1278 (O_1278,N_8730,N_8871);
nor UO_1279 (O_1279,N_8281,N_9065);
xor UO_1280 (O_1280,N_9543,N_8376);
nand UO_1281 (O_1281,N_8898,N_9929);
and UO_1282 (O_1282,N_9037,N_8849);
and UO_1283 (O_1283,N_8237,N_8265);
xnor UO_1284 (O_1284,N_9943,N_8039);
and UO_1285 (O_1285,N_8091,N_8409);
nor UO_1286 (O_1286,N_9183,N_8475);
xnor UO_1287 (O_1287,N_9702,N_9918);
xor UO_1288 (O_1288,N_8353,N_9197);
nor UO_1289 (O_1289,N_8478,N_8662);
nor UO_1290 (O_1290,N_9874,N_8279);
and UO_1291 (O_1291,N_8437,N_9519);
or UO_1292 (O_1292,N_8347,N_8703);
nor UO_1293 (O_1293,N_9127,N_9025);
and UO_1294 (O_1294,N_8775,N_8349);
xnor UO_1295 (O_1295,N_8510,N_9673);
xnor UO_1296 (O_1296,N_9578,N_8511);
nor UO_1297 (O_1297,N_8245,N_8660);
nand UO_1298 (O_1298,N_9642,N_9296);
xnor UO_1299 (O_1299,N_8281,N_9916);
nand UO_1300 (O_1300,N_8392,N_8639);
nand UO_1301 (O_1301,N_9490,N_8314);
and UO_1302 (O_1302,N_8471,N_9474);
and UO_1303 (O_1303,N_8402,N_8220);
xor UO_1304 (O_1304,N_9666,N_8864);
and UO_1305 (O_1305,N_9596,N_9479);
nand UO_1306 (O_1306,N_8211,N_9823);
or UO_1307 (O_1307,N_8613,N_8540);
nor UO_1308 (O_1308,N_9692,N_9765);
nand UO_1309 (O_1309,N_9555,N_8322);
nand UO_1310 (O_1310,N_8984,N_8922);
nor UO_1311 (O_1311,N_9241,N_8904);
nand UO_1312 (O_1312,N_8171,N_9036);
nor UO_1313 (O_1313,N_8610,N_8546);
nor UO_1314 (O_1314,N_8116,N_8984);
nor UO_1315 (O_1315,N_8896,N_9154);
nand UO_1316 (O_1316,N_8878,N_9436);
or UO_1317 (O_1317,N_9069,N_9585);
nand UO_1318 (O_1318,N_9654,N_8710);
xnor UO_1319 (O_1319,N_9970,N_9139);
or UO_1320 (O_1320,N_8604,N_8119);
and UO_1321 (O_1321,N_8513,N_8262);
nand UO_1322 (O_1322,N_8614,N_9454);
nand UO_1323 (O_1323,N_9037,N_9420);
or UO_1324 (O_1324,N_8325,N_9063);
nor UO_1325 (O_1325,N_9619,N_8054);
or UO_1326 (O_1326,N_9698,N_9760);
xnor UO_1327 (O_1327,N_9838,N_9048);
nor UO_1328 (O_1328,N_8706,N_8913);
and UO_1329 (O_1329,N_9926,N_8827);
xnor UO_1330 (O_1330,N_8814,N_8574);
or UO_1331 (O_1331,N_9488,N_9088);
xor UO_1332 (O_1332,N_8006,N_9333);
nand UO_1333 (O_1333,N_9691,N_9157);
or UO_1334 (O_1334,N_8719,N_9300);
or UO_1335 (O_1335,N_9731,N_9001);
and UO_1336 (O_1336,N_8939,N_9431);
xor UO_1337 (O_1337,N_8142,N_8696);
xnor UO_1338 (O_1338,N_8678,N_9084);
nand UO_1339 (O_1339,N_9693,N_9446);
or UO_1340 (O_1340,N_8934,N_8444);
xor UO_1341 (O_1341,N_9009,N_8517);
or UO_1342 (O_1342,N_8665,N_8164);
or UO_1343 (O_1343,N_8120,N_9646);
or UO_1344 (O_1344,N_8986,N_9731);
nor UO_1345 (O_1345,N_8257,N_9382);
or UO_1346 (O_1346,N_8581,N_8048);
xnor UO_1347 (O_1347,N_9141,N_8406);
xnor UO_1348 (O_1348,N_8390,N_8400);
nor UO_1349 (O_1349,N_8485,N_9310);
xor UO_1350 (O_1350,N_8576,N_8428);
or UO_1351 (O_1351,N_9889,N_9234);
nand UO_1352 (O_1352,N_8330,N_8023);
or UO_1353 (O_1353,N_9512,N_8736);
and UO_1354 (O_1354,N_9233,N_9374);
and UO_1355 (O_1355,N_9302,N_9611);
nor UO_1356 (O_1356,N_8925,N_9627);
nor UO_1357 (O_1357,N_9547,N_9760);
nand UO_1358 (O_1358,N_8405,N_9132);
nor UO_1359 (O_1359,N_8544,N_8227);
nand UO_1360 (O_1360,N_8632,N_9051);
nor UO_1361 (O_1361,N_9959,N_8124);
or UO_1362 (O_1362,N_8213,N_9887);
xor UO_1363 (O_1363,N_9279,N_8693);
nand UO_1364 (O_1364,N_8606,N_8120);
nor UO_1365 (O_1365,N_8912,N_9233);
nor UO_1366 (O_1366,N_8572,N_8283);
nand UO_1367 (O_1367,N_8396,N_9554);
xnor UO_1368 (O_1368,N_8708,N_8223);
and UO_1369 (O_1369,N_9059,N_9850);
and UO_1370 (O_1370,N_8948,N_8057);
or UO_1371 (O_1371,N_8228,N_8350);
or UO_1372 (O_1372,N_9840,N_8269);
or UO_1373 (O_1373,N_9713,N_8426);
nand UO_1374 (O_1374,N_9614,N_9511);
xor UO_1375 (O_1375,N_9122,N_8672);
or UO_1376 (O_1376,N_8349,N_9355);
xor UO_1377 (O_1377,N_8254,N_8292);
or UO_1378 (O_1378,N_8166,N_8496);
nor UO_1379 (O_1379,N_8024,N_9567);
xnor UO_1380 (O_1380,N_8883,N_9110);
or UO_1381 (O_1381,N_9979,N_9884);
nand UO_1382 (O_1382,N_8180,N_9387);
nand UO_1383 (O_1383,N_8058,N_9578);
nand UO_1384 (O_1384,N_8484,N_8781);
and UO_1385 (O_1385,N_8722,N_8754);
or UO_1386 (O_1386,N_9136,N_9032);
nor UO_1387 (O_1387,N_9006,N_8669);
or UO_1388 (O_1388,N_8910,N_9286);
and UO_1389 (O_1389,N_8918,N_9776);
nor UO_1390 (O_1390,N_9578,N_8332);
nand UO_1391 (O_1391,N_9117,N_9290);
nor UO_1392 (O_1392,N_8131,N_9945);
nor UO_1393 (O_1393,N_8200,N_9991);
nor UO_1394 (O_1394,N_8157,N_8182);
nor UO_1395 (O_1395,N_9137,N_8907);
or UO_1396 (O_1396,N_9991,N_9372);
xor UO_1397 (O_1397,N_8263,N_8419);
or UO_1398 (O_1398,N_8312,N_8426);
xor UO_1399 (O_1399,N_9392,N_8576);
xnor UO_1400 (O_1400,N_8700,N_9244);
xor UO_1401 (O_1401,N_9066,N_9667);
xor UO_1402 (O_1402,N_9973,N_9896);
nand UO_1403 (O_1403,N_8579,N_8777);
nand UO_1404 (O_1404,N_9709,N_9238);
and UO_1405 (O_1405,N_9567,N_8986);
or UO_1406 (O_1406,N_9436,N_8361);
and UO_1407 (O_1407,N_8978,N_9828);
or UO_1408 (O_1408,N_9191,N_9112);
or UO_1409 (O_1409,N_8003,N_8871);
nor UO_1410 (O_1410,N_8830,N_8504);
or UO_1411 (O_1411,N_8952,N_9229);
and UO_1412 (O_1412,N_9761,N_9882);
nand UO_1413 (O_1413,N_8587,N_9794);
xnor UO_1414 (O_1414,N_8153,N_9977);
xnor UO_1415 (O_1415,N_9900,N_8289);
xnor UO_1416 (O_1416,N_8737,N_8996);
nand UO_1417 (O_1417,N_9830,N_8291);
nor UO_1418 (O_1418,N_8462,N_8685);
xnor UO_1419 (O_1419,N_9460,N_9103);
and UO_1420 (O_1420,N_9561,N_8230);
or UO_1421 (O_1421,N_8907,N_9009);
nor UO_1422 (O_1422,N_8078,N_9258);
or UO_1423 (O_1423,N_9553,N_8891);
and UO_1424 (O_1424,N_9319,N_9772);
nand UO_1425 (O_1425,N_9189,N_9329);
nand UO_1426 (O_1426,N_9256,N_9587);
nand UO_1427 (O_1427,N_9717,N_9219);
nor UO_1428 (O_1428,N_9385,N_9946);
xnor UO_1429 (O_1429,N_9604,N_9873);
nor UO_1430 (O_1430,N_9080,N_8286);
nor UO_1431 (O_1431,N_8368,N_9075);
xor UO_1432 (O_1432,N_9952,N_9733);
and UO_1433 (O_1433,N_9471,N_8612);
and UO_1434 (O_1434,N_9252,N_9873);
nand UO_1435 (O_1435,N_8443,N_9585);
and UO_1436 (O_1436,N_8242,N_8576);
and UO_1437 (O_1437,N_8733,N_8221);
nor UO_1438 (O_1438,N_9327,N_8056);
or UO_1439 (O_1439,N_8609,N_9458);
xnor UO_1440 (O_1440,N_8662,N_8446);
and UO_1441 (O_1441,N_8225,N_8322);
and UO_1442 (O_1442,N_8025,N_9418);
nand UO_1443 (O_1443,N_8210,N_8023);
and UO_1444 (O_1444,N_9368,N_9599);
nor UO_1445 (O_1445,N_8719,N_8757);
nand UO_1446 (O_1446,N_9149,N_8725);
or UO_1447 (O_1447,N_9767,N_8799);
and UO_1448 (O_1448,N_9096,N_8118);
and UO_1449 (O_1449,N_9906,N_8512);
and UO_1450 (O_1450,N_8367,N_9043);
nor UO_1451 (O_1451,N_8028,N_9356);
nor UO_1452 (O_1452,N_9285,N_9893);
nor UO_1453 (O_1453,N_9083,N_8273);
xnor UO_1454 (O_1454,N_8518,N_9554);
nor UO_1455 (O_1455,N_8598,N_9897);
nand UO_1456 (O_1456,N_8852,N_9157);
and UO_1457 (O_1457,N_8724,N_9927);
nor UO_1458 (O_1458,N_9457,N_8320);
and UO_1459 (O_1459,N_8176,N_9774);
nand UO_1460 (O_1460,N_9827,N_9786);
nand UO_1461 (O_1461,N_9831,N_9816);
nand UO_1462 (O_1462,N_8326,N_8903);
and UO_1463 (O_1463,N_8179,N_9885);
and UO_1464 (O_1464,N_9471,N_9788);
xnor UO_1465 (O_1465,N_9483,N_8467);
nor UO_1466 (O_1466,N_9161,N_8723);
xor UO_1467 (O_1467,N_9553,N_8615);
and UO_1468 (O_1468,N_8046,N_9481);
xor UO_1469 (O_1469,N_8569,N_9733);
nor UO_1470 (O_1470,N_9839,N_8316);
nor UO_1471 (O_1471,N_8918,N_8038);
nand UO_1472 (O_1472,N_9759,N_8745);
and UO_1473 (O_1473,N_8625,N_9758);
nor UO_1474 (O_1474,N_9447,N_8083);
and UO_1475 (O_1475,N_9830,N_8048);
xnor UO_1476 (O_1476,N_9763,N_8223);
and UO_1477 (O_1477,N_9382,N_8829);
and UO_1478 (O_1478,N_8127,N_8985);
xor UO_1479 (O_1479,N_9994,N_8234);
and UO_1480 (O_1480,N_9485,N_8980);
nand UO_1481 (O_1481,N_8869,N_9272);
and UO_1482 (O_1482,N_8019,N_8987);
xnor UO_1483 (O_1483,N_9958,N_9787);
xor UO_1484 (O_1484,N_8765,N_9988);
and UO_1485 (O_1485,N_8109,N_9245);
nor UO_1486 (O_1486,N_8474,N_9669);
nand UO_1487 (O_1487,N_8578,N_9072);
and UO_1488 (O_1488,N_9346,N_8726);
or UO_1489 (O_1489,N_8461,N_8477);
and UO_1490 (O_1490,N_8089,N_9010);
nand UO_1491 (O_1491,N_8845,N_9715);
xor UO_1492 (O_1492,N_9462,N_9780);
or UO_1493 (O_1493,N_8818,N_8656);
nand UO_1494 (O_1494,N_9932,N_9664);
or UO_1495 (O_1495,N_8899,N_8700);
and UO_1496 (O_1496,N_9832,N_9041);
or UO_1497 (O_1497,N_9094,N_8597);
or UO_1498 (O_1498,N_9559,N_8991);
xor UO_1499 (O_1499,N_9202,N_8522);
endmodule