module basic_500_3000_500_6_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_253,In_4);
xor U1 (N_1,In_192,In_332);
nand U2 (N_2,In_203,In_354);
and U3 (N_3,In_318,In_12);
nor U4 (N_4,In_337,In_47);
nor U5 (N_5,In_52,In_194);
or U6 (N_6,In_496,In_16);
nand U7 (N_7,In_408,In_326);
nand U8 (N_8,In_210,In_145);
nand U9 (N_9,In_417,In_366);
nand U10 (N_10,In_132,In_276);
nand U11 (N_11,In_205,In_365);
and U12 (N_12,In_176,In_11);
nand U13 (N_13,In_445,In_349);
xnor U14 (N_14,In_446,In_219);
and U15 (N_15,In_125,In_225);
nor U16 (N_16,In_469,In_174);
nand U17 (N_17,In_247,In_206);
nand U18 (N_18,In_70,In_135);
nand U19 (N_19,In_239,In_42);
xnor U20 (N_20,In_137,In_472);
nand U21 (N_21,In_155,In_250);
nor U22 (N_22,In_465,In_223);
and U23 (N_23,In_468,In_108);
and U24 (N_24,In_352,In_300);
nand U25 (N_25,In_311,In_343);
or U26 (N_26,In_254,In_249);
nor U27 (N_27,In_395,In_428);
nand U28 (N_28,In_298,In_6);
xnor U29 (N_29,In_296,In_269);
nor U30 (N_30,In_333,In_58);
xnor U31 (N_31,In_435,In_101);
or U32 (N_32,In_84,In_397);
nor U33 (N_33,In_463,In_270);
and U34 (N_34,In_483,In_295);
nand U35 (N_35,In_267,In_350);
nor U36 (N_36,In_30,In_455);
and U37 (N_37,In_238,In_283);
nand U38 (N_38,In_367,In_196);
xor U39 (N_39,In_369,In_44);
nand U40 (N_40,In_466,In_106);
nor U41 (N_41,In_309,In_231);
nor U42 (N_42,In_226,In_118);
or U43 (N_43,In_427,In_447);
nand U44 (N_44,In_178,In_423);
xor U45 (N_45,In_161,In_363);
or U46 (N_46,In_411,In_109);
or U47 (N_47,In_454,In_299);
xnor U48 (N_48,In_379,In_166);
nand U49 (N_49,In_214,In_188);
or U50 (N_50,In_387,In_140);
and U51 (N_51,In_76,In_378);
or U52 (N_52,In_424,In_49);
nor U53 (N_53,In_418,In_248);
nand U54 (N_54,In_464,In_77);
nand U55 (N_55,In_370,In_258);
nor U56 (N_56,In_81,In_360);
nand U57 (N_57,In_20,In_19);
nand U58 (N_58,In_376,In_237);
or U59 (N_59,In_207,In_284);
and U60 (N_60,In_229,In_128);
xnor U61 (N_61,In_124,In_436);
and U62 (N_62,In_22,In_181);
or U63 (N_63,In_215,In_480);
xnor U64 (N_64,In_191,In_69);
or U65 (N_65,In_142,In_51);
and U66 (N_66,In_224,In_55);
nor U67 (N_67,In_230,In_95);
nand U68 (N_68,In_279,In_347);
xor U69 (N_69,In_87,In_195);
and U70 (N_70,In_107,In_285);
and U71 (N_71,In_494,In_104);
nor U72 (N_72,In_38,In_8);
or U73 (N_73,In_96,In_153);
xnor U74 (N_74,In_256,In_273);
or U75 (N_75,In_323,In_425);
nand U76 (N_76,In_272,In_340);
nor U77 (N_77,In_313,In_32);
or U78 (N_78,In_24,In_45);
or U79 (N_79,In_410,In_458);
or U80 (N_80,In_157,In_146);
nor U81 (N_81,In_335,In_110);
xnor U82 (N_82,In_443,In_263);
xor U83 (N_83,In_170,In_438);
and U84 (N_84,In_57,In_26);
xnor U85 (N_85,In_489,In_23);
or U86 (N_86,In_372,In_355);
and U87 (N_87,In_13,In_310);
nand U88 (N_88,In_402,In_131);
xnor U89 (N_89,In_393,In_312);
nor U90 (N_90,In_394,In_162);
or U91 (N_91,In_477,In_232);
nor U92 (N_92,In_34,In_172);
xnor U93 (N_93,In_433,In_136);
and U94 (N_94,In_481,In_92);
nand U95 (N_95,In_86,In_344);
or U96 (N_96,In_260,In_121);
xor U97 (N_97,In_143,In_61);
nor U98 (N_98,In_88,In_327);
nand U99 (N_99,In_396,In_245);
xnor U100 (N_100,In_202,In_325);
and U101 (N_101,In_175,In_189);
or U102 (N_102,In_316,In_241);
or U103 (N_103,In_380,In_97);
and U104 (N_104,In_25,In_53);
or U105 (N_105,In_127,In_287);
nor U106 (N_106,In_83,In_421);
nor U107 (N_107,In_35,In_100);
nand U108 (N_108,In_374,In_193);
xnor U109 (N_109,In_307,In_407);
and U110 (N_110,In_169,In_199);
or U111 (N_111,In_420,In_14);
nor U112 (N_112,In_102,In_17);
xnor U113 (N_113,In_268,In_246);
or U114 (N_114,In_401,In_304);
nand U115 (N_115,In_460,In_452);
xnor U116 (N_116,In_375,In_266);
or U117 (N_117,In_338,In_475);
and U118 (N_118,In_15,In_383);
and U119 (N_119,In_117,In_453);
or U120 (N_120,In_400,In_331);
and U121 (N_121,In_437,In_99);
or U122 (N_122,In_391,In_498);
or U123 (N_123,In_430,In_364);
nand U124 (N_124,In_220,In_5);
or U125 (N_125,In_368,In_67);
or U126 (N_126,In_114,In_150);
xor U127 (N_127,In_21,In_27);
nand U128 (N_128,In_160,In_409);
nor U129 (N_129,In_462,In_474);
xnor U130 (N_130,In_432,In_68);
xor U131 (N_131,In_154,In_186);
xor U132 (N_132,In_493,In_73);
xor U133 (N_133,In_164,In_471);
and U134 (N_134,In_82,In_315);
nor U135 (N_135,In_62,In_209);
or U136 (N_136,In_80,In_257);
nor U137 (N_137,In_37,In_36);
nor U138 (N_138,In_18,In_441);
xor U139 (N_139,In_179,In_426);
or U140 (N_140,In_29,In_294);
or U141 (N_141,In_56,In_54);
nand U142 (N_142,In_324,In_90);
nand U143 (N_143,In_93,In_358);
or U144 (N_144,In_292,In_317);
nand U145 (N_145,In_31,In_242);
xor U146 (N_146,In_373,In_450);
nand U147 (N_147,In_412,In_303);
nand U148 (N_148,In_444,In_329);
xnor U149 (N_149,In_308,In_305);
nor U150 (N_150,In_478,In_200);
nor U151 (N_151,In_159,In_377);
or U152 (N_152,In_28,In_198);
xor U153 (N_153,In_7,In_265);
nand U154 (N_154,In_399,In_322);
xnor U155 (N_155,In_499,In_75);
and U156 (N_156,In_43,In_227);
or U157 (N_157,In_431,In_259);
and U158 (N_158,In_130,In_341);
nand U159 (N_159,In_115,In_281);
or U160 (N_160,In_339,In_385);
nand U161 (N_161,In_217,In_342);
or U162 (N_162,In_334,In_158);
nor U163 (N_163,In_94,In_251);
nand U164 (N_164,In_138,In_415);
nor U165 (N_165,In_359,In_275);
nand U166 (N_166,In_105,In_252);
nor U167 (N_167,In_91,In_320);
nand U168 (N_168,In_497,In_356);
nand U169 (N_169,In_204,In_183);
nor U170 (N_170,In_476,In_488);
nand U171 (N_171,In_171,In_182);
nor U172 (N_172,In_280,In_470);
nand U173 (N_173,In_346,In_277);
nor U174 (N_174,In_2,In_244);
nand U175 (N_175,In_163,In_353);
nor U176 (N_176,In_141,In_216);
or U177 (N_177,In_336,In_9);
nor U178 (N_178,In_213,In_165);
xnor U179 (N_179,In_388,In_235);
and U180 (N_180,In_39,In_149);
xor U181 (N_181,In_293,In_261);
and U182 (N_182,In_167,In_78);
and U183 (N_183,In_405,In_467);
nor U184 (N_184,In_33,In_361);
nand U185 (N_185,In_274,In_222);
xor U186 (N_186,In_74,In_404);
and U187 (N_187,In_10,In_484);
xor U188 (N_188,In_406,In_439);
or U189 (N_189,In_103,In_3);
and U190 (N_190,In_306,In_139);
or U191 (N_191,In_123,In_148);
or U192 (N_192,In_151,In_180);
xor U193 (N_193,In_79,In_113);
and U194 (N_194,In_390,In_384);
xnor U195 (N_195,In_449,In_456);
xnor U196 (N_196,In_398,In_46);
or U197 (N_197,In_282,In_319);
nand U198 (N_198,In_351,In_416);
and U199 (N_199,In_286,In_211);
or U200 (N_200,In_414,In_419);
nor U201 (N_201,In_386,In_168);
nand U202 (N_202,In_64,In_389);
and U203 (N_203,In_490,In_262);
nor U204 (N_204,In_403,In_65);
xnor U205 (N_205,In_392,In_89);
nor U206 (N_206,In_330,In_413);
nor U207 (N_207,In_190,In_461);
or U208 (N_208,In_184,In_278);
or U209 (N_209,In_264,In_212);
nand U210 (N_210,In_156,In_328);
nand U211 (N_211,In_98,In_485);
or U212 (N_212,In_85,In_197);
or U213 (N_213,In_345,In_187);
and U214 (N_214,In_208,In_48);
and U215 (N_215,In_288,In_482);
or U216 (N_216,In_236,In_66);
xor U217 (N_217,In_290,In_50);
nand U218 (N_218,In_134,In_41);
xnor U219 (N_219,In_233,In_381);
xor U220 (N_220,In_301,In_255);
or U221 (N_221,In_357,In_442);
and U222 (N_222,In_243,In_440);
or U223 (N_223,In_116,In_289);
and U224 (N_224,In_459,In_451);
xnor U225 (N_225,In_448,In_147);
and U226 (N_226,In_348,In_120);
nand U227 (N_227,In_434,In_129);
or U228 (N_228,In_60,In_457);
xor U229 (N_229,In_218,In_133);
nor U230 (N_230,In_63,In_302);
nor U231 (N_231,In_1,In_119);
xnor U232 (N_232,In_228,In_177);
nand U233 (N_233,In_234,In_173);
nand U234 (N_234,In_429,In_291);
or U235 (N_235,In_479,In_71);
xor U236 (N_236,In_240,In_122);
and U237 (N_237,In_72,In_321);
nor U238 (N_238,In_112,In_487);
and U239 (N_239,In_473,In_126);
xnor U240 (N_240,In_144,In_152);
and U241 (N_241,In_486,In_185);
or U242 (N_242,In_221,In_422);
nor U243 (N_243,In_382,In_492);
xnor U244 (N_244,In_495,In_59);
xor U245 (N_245,In_40,In_0);
or U246 (N_246,In_371,In_362);
or U247 (N_247,In_201,In_314);
or U248 (N_248,In_297,In_491);
or U249 (N_249,In_271,In_111);
or U250 (N_250,In_177,In_395);
and U251 (N_251,In_313,In_420);
or U252 (N_252,In_93,In_459);
nand U253 (N_253,In_288,In_346);
and U254 (N_254,In_451,In_373);
or U255 (N_255,In_289,In_299);
nor U256 (N_256,In_461,In_319);
or U257 (N_257,In_297,In_472);
and U258 (N_258,In_28,In_122);
nand U259 (N_259,In_377,In_469);
nand U260 (N_260,In_156,In_279);
nand U261 (N_261,In_462,In_414);
and U262 (N_262,In_393,In_52);
nor U263 (N_263,In_430,In_148);
and U264 (N_264,In_83,In_82);
nor U265 (N_265,In_39,In_306);
nor U266 (N_266,In_79,In_171);
nor U267 (N_267,In_139,In_34);
nor U268 (N_268,In_405,In_73);
or U269 (N_269,In_409,In_0);
and U270 (N_270,In_10,In_491);
xor U271 (N_271,In_479,In_111);
or U272 (N_272,In_260,In_392);
nor U273 (N_273,In_249,In_260);
and U274 (N_274,In_339,In_138);
nand U275 (N_275,In_165,In_443);
nor U276 (N_276,In_425,In_413);
nand U277 (N_277,In_200,In_131);
and U278 (N_278,In_163,In_175);
nand U279 (N_279,In_196,In_216);
nor U280 (N_280,In_84,In_494);
nor U281 (N_281,In_54,In_300);
nand U282 (N_282,In_279,In_25);
nand U283 (N_283,In_382,In_299);
nand U284 (N_284,In_116,In_261);
or U285 (N_285,In_18,In_68);
and U286 (N_286,In_226,In_95);
nor U287 (N_287,In_67,In_45);
and U288 (N_288,In_214,In_312);
and U289 (N_289,In_323,In_129);
xnor U290 (N_290,In_482,In_340);
xor U291 (N_291,In_136,In_323);
xor U292 (N_292,In_45,In_497);
and U293 (N_293,In_244,In_175);
or U294 (N_294,In_180,In_341);
and U295 (N_295,In_164,In_175);
or U296 (N_296,In_43,In_236);
or U297 (N_297,In_425,In_440);
and U298 (N_298,In_389,In_140);
nand U299 (N_299,In_81,In_451);
nand U300 (N_300,In_371,In_77);
nand U301 (N_301,In_131,In_79);
nand U302 (N_302,In_422,In_477);
xor U303 (N_303,In_474,In_51);
xor U304 (N_304,In_75,In_159);
nor U305 (N_305,In_170,In_407);
nor U306 (N_306,In_408,In_18);
nor U307 (N_307,In_251,In_447);
xnor U308 (N_308,In_385,In_71);
nand U309 (N_309,In_312,In_245);
and U310 (N_310,In_275,In_380);
xnor U311 (N_311,In_433,In_374);
nand U312 (N_312,In_291,In_496);
xnor U313 (N_313,In_39,In_318);
nand U314 (N_314,In_286,In_380);
and U315 (N_315,In_185,In_339);
xnor U316 (N_316,In_148,In_290);
xnor U317 (N_317,In_280,In_350);
and U318 (N_318,In_371,In_300);
and U319 (N_319,In_390,In_132);
and U320 (N_320,In_76,In_129);
nand U321 (N_321,In_275,In_457);
xnor U322 (N_322,In_306,In_122);
nand U323 (N_323,In_183,In_120);
nor U324 (N_324,In_212,In_332);
and U325 (N_325,In_54,In_400);
xor U326 (N_326,In_97,In_234);
and U327 (N_327,In_291,In_263);
or U328 (N_328,In_29,In_436);
nor U329 (N_329,In_71,In_66);
and U330 (N_330,In_427,In_226);
or U331 (N_331,In_91,In_228);
or U332 (N_332,In_451,In_248);
xnor U333 (N_333,In_477,In_64);
xor U334 (N_334,In_100,In_384);
and U335 (N_335,In_267,In_472);
xor U336 (N_336,In_87,In_224);
and U337 (N_337,In_64,In_32);
nor U338 (N_338,In_136,In_382);
nand U339 (N_339,In_339,In_25);
nor U340 (N_340,In_472,In_445);
nand U341 (N_341,In_12,In_240);
nand U342 (N_342,In_451,In_198);
xor U343 (N_343,In_480,In_244);
nand U344 (N_344,In_307,In_301);
nand U345 (N_345,In_118,In_460);
and U346 (N_346,In_311,In_175);
nand U347 (N_347,In_493,In_242);
nor U348 (N_348,In_417,In_9);
nor U349 (N_349,In_408,In_53);
nand U350 (N_350,In_32,In_404);
nor U351 (N_351,In_306,In_20);
nor U352 (N_352,In_50,In_11);
or U353 (N_353,In_151,In_7);
nor U354 (N_354,In_418,In_284);
and U355 (N_355,In_159,In_305);
or U356 (N_356,In_107,In_422);
and U357 (N_357,In_497,In_36);
or U358 (N_358,In_394,In_493);
and U359 (N_359,In_8,In_203);
or U360 (N_360,In_53,In_92);
and U361 (N_361,In_56,In_166);
nand U362 (N_362,In_439,In_136);
and U363 (N_363,In_420,In_303);
nand U364 (N_364,In_380,In_158);
xnor U365 (N_365,In_274,In_149);
or U366 (N_366,In_441,In_3);
nor U367 (N_367,In_432,In_190);
xnor U368 (N_368,In_121,In_393);
nand U369 (N_369,In_408,In_254);
and U370 (N_370,In_461,In_375);
and U371 (N_371,In_281,In_81);
xor U372 (N_372,In_321,In_207);
nand U373 (N_373,In_471,In_34);
xnor U374 (N_374,In_298,In_16);
xnor U375 (N_375,In_444,In_370);
or U376 (N_376,In_11,In_429);
xor U377 (N_377,In_340,In_11);
xnor U378 (N_378,In_223,In_283);
nor U379 (N_379,In_318,In_31);
and U380 (N_380,In_81,In_290);
or U381 (N_381,In_464,In_479);
nor U382 (N_382,In_243,In_331);
or U383 (N_383,In_296,In_83);
nand U384 (N_384,In_451,In_1);
or U385 (N_385,In_252,In_390);
nand U386 (N_386,In_159,In_77);
or U387 (N_387,In_114,In_358);
nand U388 (N_388,In_477,In_412);
nand U389 (N_389,In_37,In_457);
nand U390 (N_390,In_394,In_10);
nor U391 (N_391,In_5,In_397);
or U392 (N_392,In_22,In_396);
or U393 (N_393,In_116,In_55);
xor U394 (N_394,In_251,In_385);
and U395 (N_395,In_183,In_445);
nor U396 (N_396,In_346,In_345);
or U397 (N_397,In_192,In_317);
or U398 (N_398,In_231,In_426);
or U399 (N_399,In_429,In_378);
nor U400 (N_400,In_10,In_28);
xor U401 (N_401,In_289,In_411);
and U402 (N_402,In_122,In_418);
xnor U403 (N_403,In_484,In_263);
nand U404 (N_404,In_317,In_460);
and U405 (N_405,In_463,In_451);
and U406 (N_406,In_466,In_351);
nand U407 (N_407,In_417,In_260);
and U408 (N_408,In_455,In_112);
or U409 (N_409,In_116,In_71);
nand U410 (N_410,In_240,In_303);
xor U411 (N_411,In_12,In_407);
or U412 (N_412,In_5,In_482);
nand U413 (N_413,In_391,In_138);
and U414 (N_414,In_193,In_207);
xnor U415 (N_415,In_214,In_27);
and U416 (N_416,In_372,In_422);
or U417 (N_417,In_98,In_357);
xor U418 (N_418,In_8,In_350);
or U419 (N_419,In_309,In_426);
xor U420 (N_420,In_50,In_174);
nor U421 (N_421,In_468,In_131);
nor U422 (N_422,In_489,In_93);
nor U423 (N_423,In_208,In_96);
xnor U424 (N_424,In_469,In_384);
nand U425 (N_425,In_455,In_100);
and U426 (N_426,In_183,In_348);
and U427 (N_427,In_223,In_313);
nor U428 (N_428,In_264,In_224);
or U429 (N_429,In_223,In_115);
or U430 (N_430,In_444,In_148);
nor U431 (N_431,In_442,In_152);
or U432 (N_432,In_389,In_164);
xnor U433 (N_433,In_186,In_346);
nor U434 (N_434,In_370,In_421);
or U435 (N_435,In_128,In_47);
xor U436 (N_436,In_152,In_239);
nand U437 (N_437,In_440,In_444);
and U438 (N_438,In_491,In_410);
nand U439 (N_439,In_390,In_388);
or U440 (N_440,In_125,In_401);
or U441 (N_441,In_216,In_213);
nor U442 (N_442,In_329,In_410);
xnor U443 (N_443,In_229,In_53);
or U444 (N_444,In_464,In_284);
nor U445 (N_445,In_1,In_74);
nand U446 (N_446,In_305,In_421);
nor U447 (N_447,In_202,In_239);
or U448 (N_448,In_142,In_364);
nand U449 (N_449,In_207,In_338);
nand U450 (N_450,In_452,In_418);
nor U451 (N_451,In_480,In_8);
nand U452 (N_452,In_409,In_337);
or U453 (N_453,In_137,In_169);
xor U454 (N_454,In_394,In_262);
or U455 (N_455,In_375,In_273);
nor U456 (N_456,In_211,In_42);
nor U457 (N_457,In_116,In_139);
nor U458 (N_458,In_300,In_476);
or U459 (N_459,In_202,In_481);
nand U460 (N_460,In_113,In_65);
and U461 (N_461,In_119,In_145);
xnor U462 (N_462,In_272,In_326);
nand U463 (N_463,In_329,In_228);
xnor U464 (N_464,In_267,In_33);
xnor U465 (N_465,In_149,In_477);
nor U466 (N_466,In_237,In_64);
or U467 (N_467,In_133,In_157);
nand U468 (N_468,In_323,In_376);
xnor U469 (N_469,In_296,In_26);
or U470 (N_470,In_336,In_481);
nand U471 (N_471,In_66,In_101);
nor U472 (N_472,In_102,In_4);
or U473 (N_473,In_330,In_258);
nand U474 (N_474,In_41,In_179);
xor U475 (N_475,In_454,In_414);
nand U476 (N_476,In_334,In_9);
nor U477 (N_477,In_350,In_247);
and U478 (N_478,In_424,In_309);
nand U479 (N_479,In_27,In_332);
and U480 (N_480,In_331,In_256);
nand U481 (N_481,In_55,In_189);
xor U482 (N_482,In_298,In_497);
nor U483 (N_483,In_77,In_246);
or U484 (N_484,In_209,In_122);
nand U485 (N_485,In_156,In_105);
or U486 (N_486,In_133,In_64);
xor U487 (N_487,In_134,In_214);
nor U488 (N_488,In_378,In_398);
nand U489 (N_489,In_321,In_439);
and U490 (N_490,In_215,In_256);
or U491 (N_491,In_62,In_16);
or U492 (N_492,In_358,In_103);
xnor U493 (N_493,In_97,In_312);
and U494 (N_494,In_82,In_58);
or U495 (N_495,In_68,In_365);
xnor U496 (N_496,In_336,In_239);
or U497 (N_497,In_219,In_235);
nand U498 (N_498,In_21,In_319);
nand U499 (N_499,In_49,In_405);
nand U500 (N_500,N_354,N_350);
nand U501 (N_501,N_111,N_389);
xor U502 (N_502,N_16,N_480);
xnor U503 (N_503,N_7,N_273);
and U504 (N_504,N_46,N_171);
and U505 (N_505,N_123,N_318);
or U506 (N_506,N_258,N_378);
nor U507 (N_507,N_260,N_62);
xnor U508 (N_508,N_253,N_78);
xor U509 (N_509,N_150,N_189);
or U510 (N_510,N_328,N_84);
nand U511 (N_511,N_398,N_327);
or U512 (N_512,N_358,N_426);
and U513 (N_513,N_54,N_221);
xor U514 (N_514,N_263,N_160);
and U515 (N_515,N_333,N_77);
nand U516 (N_516,N_270,N_414);
or U517 (N_517,N_347,N_104);
or U518 (N_518,N_365,N_282);
nor U519 (N_519,N_198,N_292);
nor U520 (N_520,N_124,N_24);
nand U521 (N_521,N_34,N_373);
nand U522 (N_522,N_19,N_312);
xnor U523 (N_523,N_22,N_146);
or U524 (N_524,N_473,N_344);
and U525 (N_525,N_453,N_310);
nor U526 (N_526,N_108,N_408);
nand U527 (N_527,N_193,N_174);
or U528 (N_528,N_213,N_413);
nand U529 (N_529,N_116,N_467);
nor U530 (N_530,N_412,N_166);
nand U531 (N_531,N_243,N_313);
nor U532 (N_532,N_12,N_289);
xnor U533 (N_533,N_379,N_52);
xor U534 (N_534,N_307,N_172);
and U535 (N_535,N_141,N_368);
or U536 (N_536,N_291,N_232);
xnor U537 (N_537,N_164,N_406);
nand U538 (N_538,N_457,N_364);
xnor U539 (N_539,N_323,N_251);
nand U540 (N_540,N_149,N_458);
xor U541 (N_541,N_465,N_451);
nor U542 (N_542,N_76,N_380);
nor U543 (N_543,N_167,N_197);
or U544 (N_544,N_227,N_359);
nor U545 (N_545,N_439,N_429);
or U546 (N_546,N_462,N_423);
and U547 (N_547,N_71,N_317);
and U548 (N_548,N_181,N_10);
nor U549 (N_549,N_53,N_95);
xnor U550 (N_550,N_210,N_417);
and U551 (N_551,N_311,N_316);
nor U552 (N_552,N_298,N_67);
xnor U553 (N_553,N_300,N_185);
nand U554 (N_554,N_60,N_231);
nand U555 (N_555,N_262,N_200);
and U556 (N_556,N_397,N_25);
nand U557 (N_557,N_168,N_305);
nor U558 (N_558,N_214,N_450);
nor U559 (N_559,N_91,N_479);
nor U560 (N_560,N_159,N_471);
xnor U561 (N_561,N_395,N_226);
nor U562 (N_562,N_447,N_4);
nand U563 (N_563,N_399,N_348);
nand U564 (N_564,N_88,N_268);
nor U565 (N_565,N_331,N_6);
and U566 (N_566,N_265,N_72);
xnor U567 (N_567,N_446,N_37);
nand U568 (N_568,N_382,N_236);
or U569 (N_569,N_180,N_135);
nor U570 (N_570,N_363,N_217);
and U571 (N_571,N_315,N_51);
nor U572 (N_572,N_448,N_29);
and U573 (N_573,N_411,N_342);
or U574 (N_574,N_83,N_47);
xor U575 (N_575,N_144,N_184);
nor U576 (N_576,N_163,N_470);
nand U577 (N_577,N_341,N_82);
or U578 (N_578,N_267,N_407);
or U579 (N_579,N_339,N_321);
nand U580 (N_580,N_2,N_287);
nor U581 (N_581,N_207,N_9);
nor U582 (N_582,N_374,N_250);
nor U583 (N_583,N_432,N_175);
and U584 (N_584,N_396,N_422);
nor U585 (N_585,N_121,N_301);
and U586 (N_586,N_240,N_427);
xnor U587 (N_587,N_58,N_438);
nor U588 (N_588,N_196,N_367);
or U589 (N_589,N_230,N_103);
nor U590 (N_590,N_375,N_235);
nand U591 (N_591,N_11,N_353);
and U592 (N_592,N_306,N_314);
and U593 (N_593,N_195,N_254);
nand U594 (N_594,N_114,N_370);
xor U595 (N_595,N_122,N_241);
xnor U596 (N_596,N_409,N_154);
and U597 (N_597,N_410,N_387);
and U598 (N_598,N_281,N_393);
nand U599 (N_599,N_170,N_117);
or U600 (N_600,N_418,N_142);
nand U601 (N_601,N_1,N_15);
nand U602 (N_602,N_351,N_415);
and U603 (N_603,N_182,N_452);
or U604 (N_604,N_183,N_404);
xnor U605 (N_605,N_176,N_157);
nor U606 (N_606,N_376,N_120);
nand U607 (N_607,N_107,N_355);
xnor U608 (N_608,N_31,N_86);
nor U609 (N_609,N_188,N_400);
or U610 (N_610,N_464,N_274);
nand U611 (N_611,N_179,N_383);
nor U612 (N_612,N_199,N_224);
and U613 (N_613,N_455,N_105);
or U614 (N_614,N_192,N_303);
nand U615 (N_615,N_162,N_366);
nand U616 (N_616,N_201,N_23);
nor U617 (N_617,N_297,N_456);
and U618 (N_618,N_74,N_57);
nor U619 (N_619,N_324,N_481);
or U620 (N_620,N_486,N_68);
nand U621 (N_621,N_360,N_443);
nor U622 (N_622,N_466,N_206);
or U623 (N_623,N_469,N_81);
or U624 (N_624,N_92,N_186);
nand U625 (N_625,N_238,N_478);
nor U626 (N_626,N_334,N_112);
and U627 (N_627,N_229,N_156);
nand U628 (N_628,N_35,N_33);
nand U629 (N_629,N_336,N_204);
nor U630 (N_630,N_43,N_138);
nand U631 (N_631,N_246,N_442);
nor U632 (N_632,N_290,N_219);
xnor U633 (N_633,N_165,N_346);
and U634 (N_634,N_202,N_209);
nand U635 (N_635,N_484,N_416);
nor U636 (N_636,N_340,N_61);
or U637 (N_637,N_169,N_433);
or U638 (N_638,N_187,N_304);
nand U639 (N_639,N_498,N_237);
nand U640 (N_640,N_132,N_215);
xnor U641 (N_641,N_381,N_128);
and U642 (N_642,N_475,N_284);
and U643 (N_643,N_64,N_269);
xor U644 (N_644,N_492,N_405);
or U645 (N_645,N_216,N_17);
and U646 (N_646,N_110,N_45);
nand U647 (N_647,N_94,N_140);
or U648 (N_648,N_101,N_113);
xnor U649 (N_649,N_26,N_50);
and U650 (N_650,N_444,N_402);
nand U651 (N_651,N_338,N_161);
xor U652 (N_652,N_326,N_220);
xor U653 (N_653,N_30,N_425);
nand U654 (N_654,N_431,N_392);
and U655 (N_655,N_75,N_32);
and U656 (N_656,N_203,N_496);
nor U657 (N_657,N_28,N_255);
xnor U658 (N_658,N_280,N_434);
nand U659 (N_659,N_153,N_391);
nand U660 (N_660,N_39,N_491);
nand U661 (N_661,N_0,N_440);
nand U662 (N_662,N_40,N_386);
and U663 (N_663,N_283,N_394);
or U664 (N_664,N_69,N_79);
nand U665 (N_665,N_463,N_90);
and U666 (N_666,N_56,N_335);
and U667 (N_667,N_8,N_247);
and U668 (N_668,N_41,N_436);
xnor U669 (N_669,N_385,N_158);
and U670 (N_670,N_137,N_131);
nor U671 (N_671,N_489,N_18);
or U672 (N_672,N_278,N_228);
and U673 (N_673,N_279,N_369);
xnor U674 (N_674,N_89,N_190);
nand U675 (N_675,N_99,N_133);
nor U676 (N_676,N_468,N_497);
or U677 (N_677,N_302,N_119);
and U678 (N_678,N_384,N_356);
nor U679 (N_679,N_441,N_118);
or U680 (N_680,N_66,N_377);
nand U681 (N_681,N_460,N_14);
and U682 (N_682,N_372,N_208);
and U683 (N_683,N_225,N_349);
xnor U684 (N_684,N_459,N_257);
nand U685 (N_685,N_143,N_419);
or U686 (N_686,N_3,N_134);
or U687 (N_687,N_97,N_93);
nand U688 (N_688,N_106,N_435);
nand U689 (N_689,N_44,N_309);
nand U690 (N_690,N_294,N_275);
or U691 (N_691,N_211,N_403);
or U692 (N_692,N_177,N_130);
nor U693 (N_693,N_218,N_482);
xnor U694 (N_694,N_65,N_252);
nand U695 (N_695,N_499,N_147);
nor U696 (N_696,N_320,N_286);
nand U697 (N_697,N_80,N_38);
nand U698 (N_698,N_73,N_102);
xnor U699 (N_699,N_299,N_139);
xor U700 (N_700,N_322,N_319);
xor U701 (N_701,N_495,N_249);
xnor U702 (N_702,N_98,N_295);
nor U703 (N_703,N_296,N_485);
or U704 (N_704,N_63,N_454);
and U705 (N_705,N_127,N_420);
and U706 (N_706,N_125,N_362);
and U707 (N_707,N_245,N_388);
xor U708 (N_708,N_87,N_276);
and U709 (N_709,N_48,N_266);
nor U710 (N_710,N_272,N_244);
xnor U711 (N_711,N_477,N_261);
nor U712 (N_712,N_330,N_490);
xnor U713 (N_713,N_194,N_126);
nand U714 (N_714,N_239,N_109);
and U715 (N_715,N_148,N_129);
nand U716 (N_716,N_233,N_325);
and U717 (N_717,N_424,N_449);
xor U718 (N_718,N_488,N_27);
or U719 (N_719,N_332,N_151);
xnor U720 (N_720,N_173,N_96);
nand U721 (N_721,N_430,N_421);
nor U722 (N_722,N_361,N_371);
nor U723 (N_723,N_42,N_248);
nand U724 (N_724,N_483,N_293);
nor U725 (N_725,N_36,N_59);
nor U726 (N_726,N_285,N_55);
and U727 (N_727,N_437,N_205);
nor U728 (N_728,N_242,N_337);
or U729 (N_729,N_308,N_70);
xor U730 (N_730,N_494,N_277);
nand U731 (N_731,N_13,N_390);
and U732 (N_732,N_259,N_136);
or U733 (N_733,N_493,N_145);
nor U734 (N_734,N_445,N_222);
and U735 (N_735,N_223,N_178);
nor U736 (N_736,N_5,N_212);
nand U737 (N_737,N_428,N_155);
and U738 (N_738,N_487,N_264);
or U739 (N_739,N_329,N_357);
nor U740 (N_740,N_256,N_401);
and U741 (N_741,N_21,N_49);
or U742 (N_742,N_288,N_352);
or U743 (N_743,N_345,N_474);
nand U744 (N_744,N_461,N_472);
xnor U745 (N_745,N_115,N_20);
nand U746 (N_746,N_234,N_152);
nor U747 (N_747,N_271,N_85);
nor U748 (N_748,N_100,N_476);
nor U749 (N_749,N_343,N_191);
nand U750 (N_750,N_63,N_276);
nand U751 (N_751,N_459,N_82);
nand U752 (N_752,N_197,N_289);
and U753 (N_753,N_15,N_54);
nand U754 (N_754,N_318,N_347);
or U755 (N_755,N_41,N_61);
xnor U756 (N_756,N_245,N_23);
xor U757 (N_757,N_111,N_41);
nand U758 (N_758,N_408,N_272);
nor U759 (N_759,N_153,N_182);
nor U760 (N_760,N_294,N_408);
and U761 (N_761,N_159,N_278);
nand U762 (N_762,N_235,N_170);
or U763 (N_763,N_371,N_306);
xor U764 (N_764,N_78,N_266);
xnor U765 (N_765,N_192,N_285);
xnor U766 (N_766,N_323,N_256);
or U767 (N_767,N_392,N_293);
nand U768 (N_768,N_413,N_281);
nand U769 (N_769,N_280,N_270);
xnor U770 (N_770,N_322,N_226);
and U771 (N_771,N_462,N_40);
xor U772 (N_772,N_283,N_37);
xnor U773 (N_773,N_400,N_167);
xor U774 (N_774,N_320,N_200);
nor U775 (N_775,N_270,N_430);
nor U776 (N_776,N_106,N_353);
nand U777 (N_777,N_31,N_297);
nor U778 (N_778,N_208,N_394);
and U779 (N_779,N_81,N_265);
nand U780 (N_780,N_162,N_234);
and U781 (N_781,N_11,N_356);
nor U782 (N_782,N_75,N_268);
xor U783 (N_783,N_422,N_291);
nand U784 (N_784,N_169,N_303);
nor U785 (N_785,N_156,N_406);
nor U786 (N_786,N_437,N_421);
xnor U787 (N_787,N_288,N_212);
and U788 (N_788,N_94,N_210);
nor U789 (N_789,N_446,N_175);
and U790 (N_790,N_147,N_82);
and U791 (N_791,N_114,N_298);
nand U792 (N_792,N_59,N_224);
xor U793 (N_793,N_122,N_252);
nor U794 (N_794,N_176,N_48);
nand U795 (N_795,N_111,N_293);
and U796 (N_796,N_273,N_44);
xor U797 (N_797,N_199,N_99);
or U798 (N_798,N_193,N_140);
and U799 (N_799,N_372,N_411);
or U800 (N_800,N_75,N_330);
and U801 (N_801,N_433,N_134);
nor U802 (N_802,N_413,N_67);
xnor U803 (N_803,N_169,N_482);
nand U804 (N_804,N_320,N_479);
or U805 (N_805,N_419,N_85);
and U806 (N_806,N_255,N_330);
or U807 (N_807,N_322,N_449);
or U808 (N_808,N_478,N_488);
and U809 (N_809,N_177,N_420);
xnor U810 (N_810,N_323,N_94);
xor U811 (N_811,N_342,N_0);
nand U812 (N_812,N_355,N_168);
nor U813 (N_813,N_337,N_396);
or U814 (N_814,N_490,N_334);
nor U815 (N_815,N_80,N_130);
and U816 (N_816,N_480,N_366);
and U817 (N_817,N_448,N_58);
nand U818 (N_818,N_43,N_53);
and U819 (N_819,N_32,N_91);
nor U820 (N_820,N_480,N_326);
nand U821 (N_821,N_116,N_357);
nand U822 (N_822,N_321,N_423);
and U823 (N_823,N_14,N_59);
nor U824 (N_824,N_160,N_9);
nor U825 (N_825,N_304,N_172);
xor U826 (N_826,N_170,N_387);
nand U827 (N_827,N_242,N_395);
or U828 (N_828,N_253,N_100);
or U829 (N_829,N_72,N_324);
nor U830 (N_830,N_278,N_108);
xnor U831 (N_831,N_48,N_298);
nor U832 (N_832,N_270,N_96);
nand U833 (N_833,N_114,N_238);
and U834 (N_834,N_311,N_318);
nor U835 (N_835,N_403,N_357);
nor U836 (N_836,N_60,N_8);
xnor U837 (N_837,N_212,N_429);
or U838 (N_838,N_319,N_347);
xnor U839 (N_839,N_269,N_55);
xnor U840 (N_840,N_195,N_296);
xnor U841 (N_841,N_444,N_262);
or U842 (N_842,N_258,N_301);
nand U843 (N_843,N_362,N_55);
xnor U844 (N_844,N_464,N_391);
and U845 (N_845,N_203,N_22);
and U846 (N_846,N_51,N_10);
nand U847 (N_847,N_378,N_463);
xor U848 (N_848,N_97,N_213);
and U849 (N_849,N_443,N_484);
or U850 (N_850,N_280,N_215);
and U851 (N_851,N_464,N_317);
and U852 (N_852,N_233,N_439);
nor U853 (N_853,N_319,N_174);
and U854 (N_854,N_292,N_375);
and U855 (N_855,N_50,N_290);
nor U856 (N_856,N_371,N_80);
nor U857 (N_857,N_325,N_323);
xor U858 (N_858,N_218,N_343);
nor U859 (N_859,N_316,N_294);
xor U860 (N_860,N_345,N_319);
xnor U861 (N_861,N_256,N_281);
nor U862 (N_862,N_156,N_429);
nand U863 (N_863,N_19,N_98);
xnor U864 (N_864,N_493,N_77);
nand U865 (N_865,N_266,N_331);
xor U866 (N_866,N_448,N_66);
xor U867 (N_867,N_439,N_183);
or U868 (N_868,N_183,N_305);
nor U869 (N_869,N_26,N_219);
xor U870 (N_870,N_85,N_46);
xnor U871 (N_871,N_148,N_462);
nand U872 (N_872,N_116,N_317);
nor U873 (N_873,N_488,N_266);
nor U874 (N_874,N_280,N_314);
nor U875 (N_875,N_394,N_189);
or U876 (N_876,N_468,N_362);
xnor U877 (N_877,N_214,N_368);
xor U878 (N_878,N_135,N_159);
nor U879 (N_879,N_443,N_455);
nor U880 (N_880,N_244,N_290);
or U881 (N_881,N_164,N_170);
or U882 (N_882,N_133,N_346);
nor U883 (N_883,N_257,N_133);
and U884 (N_884,N_289,N_205);
xnor U885 (N_885,N_332,N_434);
and U886 (N_886,N_284,N_146);
or U887 (N_887,N_308,N_198);
and U888 (N_888,N_142,N_388);
nor U889 (N_889,N_166,N_432);
nor U890 (N_890,N_8,N_13);
or U891 (N_891,N_153,N_180);
nand U892 (N_892,N_205,N_292);
or U893 (N_893,N_410,N_344);
or U894 (N_894,N_366,N_425);
nor U895 (N_895,N_468,N_329);
xor U896 (N_896,N_213,N_482);
and U897 (N_897,N_226,N_225);
or U898 (N_898,N_95,N_94);
and U899 (N_899,N_470,N_221);
and U900 (N_900,N_88,N_436);
nand U901 (N_901,N_63,N_82);
xor U902 (N_902,N_113,N_490);
nand U903 (N_903,N_208,N_453);
and U904 (N_904,N_46,N_212);
and U905 (N_905,N_204,N_281);
nand U906 (N_906,N_206,N_433);
and U907 (N_907,N_452,N_270);
and U908 (N_908,N_34,N_139);
nand U909 (N_909,N_430,N_458);
or U910 (N_910,N_281,N_406);
nand U911 (N_911,N_458,N_467);
nand U912 (N_912,N_412,N_86);
nor U913 (N_913,N_6,N_148);
or U914 (N_914,N_444,N_171);
nor U915 (N_915,N_91,N_448);
or U916 (N_916,N_79,N_87);
nor U917 (N_917,N_307,N_43);
or U918 (N_918,N_318,N_25);
or U919 (N_919,N_337,N_6);
or U920 (N_920,N_449,N_466);
xnor U921 (N_921,N_350,N_356);
nand U922 (N_922,N_393,N_135);
nor U923 (N_923,N_269,N_210);
nor U924 (N_924,N_367,N_57);
or U925 (N_925,N_476,N_83);
xnor U926 (N_926,N_465,N_337);
nand U927 (N_927,N_308,N_481);
xor U928 (N_928,N_283,N_269);
and U929 (N_929,N_123,N_282);
and U930 (N_930,N_87,N_400);
nor U931 (N_931,N_15,N_491);
and U932 (N_932,N_379,N_141);
nor U933 (N_933,N_54,N_374);
nand U934 (N_934,N_74,N_277);
nand U935 (N_935,N_285,N_222);
xor U936 (N_936,N_255,N_306);
and U937 (N_937,N_306,N_92);
and U938 (N_938,N_186,N_347);
or U939 (N_939,N_300,N_195);
nand U940 (N_940,N_369,N_438);
and U941 (N_941,N_184,N_105);
or U942 (N_942,N_381,N_256);
xnor U943 (N_943,N_353,N_487);
and U944 (N_944,N_259,N_490);
nand U945 (N_945,N_306,N_60);
nor U946 (N_946,N_336,N_330);
nor U947 (N_947,N_1,N_282);
or U948 (N_948,N_131,N_382);
or U949 (N_949,N_148,N_439);
or U950 (N_950,N_385,N_317);
nor U951 (N_951,N_396,N_329);
and U952 (N_952,N_250,N_66);
or U953 (N_953,N_498,N_57);
and U954 (N_954,N_92,N_129);
and U955 (N_955,N_182,N_132);
nor U956 (N_956,N_177,N_91);
xnor U957 (N_957,N_94,N_58);
xor U958 (N_958,N_102,N_8);
and U959 (N_959,N_405,N_171);
xnor U960 (N_960,N_201,N_21);
nand U961 (N_961,N_357,N_377);
or U962 (N_962,N_150,N_7);
xor U963 (N_963,N_444,N_217);
xor U964 (N_964,N_41,N_228);
and U965 (N_965,N_271,N_237);
xor U966 (N_966,N_54,N_292);
xor U967 (N_967,N_440,N_216);
or U968 (N_968,N_115,N_212);
nor U969 (N_969,N_194,N_82);
nand U970 (N_970,N_128,N_106);
xor U971 (N_971,N_336,N_445);
xor U972 (N_972,N_456,N_363);
and U973 (N_973,N_330,N_17);
or U974 (N_974,N_475,N_386);
and U975 (N_975,N_245,N_95);
or U976 (N_976,N_264,N_351);
or U977 (N_977,N_327,N_58);
nand U978 (N_978,N_194,N_23);
or U979 (N_979,N_422,N_156);
xor U980 (N_980,N_434,N_190);
xor U981 (N_981,N_168,N_128);
xnor U982 (N_982,N_180,N_190);
and U983 (N_983,N_103,N_173);
xor U984 (N_984,N_414,N_387);
or U985 (N_985,N_204,N_466);
and U986 (N_986,N_181,N_197);
nor U987 (N_987,N_91,N_242);
nand U988 (N_988,N_49,N_324);
nand U989 (N_989,N_258,N_421);
xor U990 (N_990,N_283,N_420);
xor U991 (N_991,N_289,N_59);
xor U992 (N_992,N_408,N_193);
or U993 (N_993,N_343,N_38);
or U994 (N_994,N_206,N_18);
nor U995 (N_995,N_496,N_366);
and U996 (N_996,N_306,N_472);
or U997 (N_997,N_344,N_90);
nor U998 (N_998,N_182,N_88);
or U999 (N_999,N_17,N_312);
nand U1000 (N_1000,N_982,N_705);
xor U1001 (N_1001,N_624,N_549);
and U1002 (N_1002,N_869,N_584);
or U1003 (N_1003,N_767,N_615);
and U1004 (N_1004,N_632,N_757);
or U1005 (N_1005,N_839,N_822);
and U1006 (N_1006,N_735,N_743);
nor U1007 (N_1007,N_818,N_726);
and U1008 (N_1008,N_708,N_664);
and U1009 (N_1009,N_947,N_628);
and U1010 (N_1010,N_682,N_667);
nor U1011 (N_1011,N_820,N_575);
nor U1012 (N_1012,N_897,N_503);
and U1013 (N_1013,N_826,N_662);
nand U1014 (N_1014,N_540,N_610);
and U1015 (N_1015,N_803,N_773);
nand U1016 (N_1016,N_988,N_514);
nand U1017 (N_1017,N_611,N_999);
or U1018 (N_1018,N_501,N_996);
xor U1019 (N_1019,N_997,N_811);
or U1020 (N_1020,N_921,N_588);
and U1021 (N_1021,N_663,N_945);
nor U1022 (N_1022,N_840,N_910);
nor U1023 (N_1023,N_983,N_967);
xnor U1024 (N_1024,N_768,N_823);
or U1025 (N_1025,N_916,N_530);
and U1026 (N_1026,N_796,N_965);
nand U1027 (N_1027,N_545,N_998);
xnor U1028 (N_1028,N_984,N_860);
xor U1029 (N_1029,N_533,N_737);
nor U1030 (N_1030,N_669,N_802);
xnor U1031 (N_1031,N_631,N_833);
and U1032 (N_1032,N_924,N_824);
nor U1033 (N_1033,N_806,N_793);
xnor U1034 (N_1034,N_932,N_849);
and U1035 (N_1035,N_707,N_755);
and U1036 (N_1036,N_790,N_729);
or U1037 (N_1037,N_504,N_557);
and U1038 (N_1038,N_856,N_966);
nand U1039 (N_1039,N_756,N_646);
xnor U1040 (N_1040,N_629,N_563);
or U1041 (N_1041,N_673,N_571);
xor U1042 (N_1042,N_934,N_854);
xnor U1043 (N_1043,N_569,N_841);
nor U1044 (N_1044,N_905,N_930);
nand U1045 (N_1045,N_969,N_781);
xor U1046 (N_1046,N_780,N_973);
nand U1047 (N_1047,N_509,N_853);
and U1048 (N_1048,N_552,N_799);
or U1049 (N_1049,N_825,N_649);
nand U1050 (N_1050,N_580,N_938);
or U1051 (N_1051,N_689,N_633);
nor U1052 (N_1052,N_694,N_668);
or U1053 (N_1053,N_654,N_920);
or U1054 (N_1054,N_817,N_637);
and U1055 (N_1055,N_522,N_936);
nand U1056 (N_1056,N_902,N_650);
nor U1057 (N_1057,N_890,N_698);
nor U1058 (N_1058,N_837,N_593);
nand U1059 (N_1059,N_625,N_550);
xor U1060 (N_1060,N_622,N_941);
nor U1061 (N_1061,N_714,N_548);
nand U1062 (N_1062,N_518,N_678);
and U1063 (N_1063,N_838,N_888);
xor U1064 (N_1064,N_738,N_538);
and U1065 (N_1065,N_885,N_736);
xnor U1066 (N_1066,N_863,N_543);
nand U1067 (N_1067,N_537,N_872);
nand U1068 (N_1068,N_685,N_570);
or U1069 (N_1069,N_604,N_990);
nand U1070 (N_1070,N_821,N_948);
and U1071 (N_1071,N_568,N_693);
xnor U1072 (N_1072,N_722,N_809);
or U1073 (N_1073,N_683,N_713);
xor U1074 (N_1074,N_894,N_962);
or U1075 (N_1075,N_758,N_532);
and U1076 (N_1076,N_627,N_517);
and U1077 (N_1077,N_715,N_908);
and U1078 (N_1078,N_725,N_659);
nor U1079 (N_1079,N_942,N_977);
nor U1080 (N_1080,N_651,N_778);
nand U1081 (N_1081,N_602,N_808);
or U1082 (N_1082,N_852,N_792);
nor U1083 (N_1083,N_536,N_762);
or U1084 (N_1084,N_697,N_641);
and U1085 (N_1085,N_992,N_787);
or U1086 (N_1086,N_845,N_868);
nand U1087 (N_1087,N_798,N_680);
nor U1088 (N_1088,N_701,N_980);
or U1089 (N_1089,N_579,N_553);
or U1090 (N_1090,N_994,N_674);
and U1091 (N_1091,N_534,N_830);
nor U1092 (N_1092,N_642,N_987);
or U1093 (N_1093,N_857,N_848);
nand U1094 (N_1094,N_859,N_658);
nor U1095 (N_1095,N_547,N_598);
and U1096 (N_1096,N_761,N_525);
xnor U1097 (N_1097,N_789,N_597);
or U1098 (N_1098,N_512,N_587);
and U1099 (N_1099,N_846,N_917);
or U1100 (N_1100,N_972,N_855);
xnor U1101 (N_1101,N_520,N_740);
and U1102 (N_1102,N_727,N_904);
and U1103 (N_1103,N_777,N_832);
nand U1104 (N_1104,N_594,N_929);
nor U1105 (N_1105,N_891,N_724);
xor U1106 (N_1106,N_807,N_576);
nand U1107 (N_1107,N_769,N_591);
nor U1108 (N_1108,N_763,N_609);
nor U1109 (N_1109,N_528,N_524);
and U1110 (N_1110,N_554,N_951);
nor U1111 (N_1111,N_788,N_562);
or U1112 (N_1112,N_559,N_739);
or U1113 (N_1113,N_623,N_665);
nor U1114 (N_1114,N_882,N_546);
or U1115 (N_1115,N_918,N_810);
nor U1116 (N_1116,N_959,N_909);
xor U1117 (N_1117,N_794,N_913);
or U1118 (N_1118,N_935,N_513);
nor U1119 (N_1119,N_883,N_887);
or U1120 (N_1120,N_889,N_523);
or U1121 (N_1121,N_816,N_616);
nor U1122 (N_1122,N_730,N_751);
nand U1123 (N_1123,N_886,N_695);
or U1124 (N_1124,N_986,N_621);
or U1125 (N_1125,N_949,N_679);
and U1126 (N_1126,N_784,N_836);
nor U1127 (N_1127,N_617,N_873);
xnor U1128 (N_1128,N_565,N_521);
xor U1129 (N_1129,N_867,N_898);
nand U1130 (N_1130,N_843,N_764);
nor U1131 (N_1131,N_515,N_690);
nor U1132 (N_1132,N_744,N_880);
nand U1133 (N_1133,N_634,N_989);
and U1134 (N_1134,N_899,N_866);
nand U1135 (N_1135,N_544,N_774);
xor U1136 (N_1136,N_814,N_605);
xor U1137 (N_1137,N_723,N_506);
nor U1138 (N_1138,N_776,N_912);
xor U1139 (N_1139,N_608,N_706);
and U1140 (N_1140,N_733,N_864);
nor U1141 (N_1141,N_970,N_981);
nor U1142 (N_1142,N_635,N_660);
xnor U1143 (N_1143,N_526,N_618);
xnor U1144 (N_1144,N_585,N_719);
nand U1145 (N_1145,N_542,N_516);
and U1146 (N_1146,N_851,N_731);
nor U1147 (N_1147,N_630,N_978);
xor U1148 (N_1148,N_815,N_510);
nand U1149 (N_1149,N_812,N_586);
xnor U1150 (N_1150,N_745,N_879);
and U1151 (N_1151,N_603,N_881);
nand U1152 (N_1152,N_566,N_895);
and U1153 (N_1153,N_960,N_589);
or U1154 (N_1154,N_979,N_871);
nand U1155 (N_1155,N_797,N_993);
xor U1156 (N_1156,N_943,N_675);
or U1157 (N_1157,N_688,N_876);
nor U1158 (N_1158,N_779,N_720);
or U1159 (N_1159,N_963,N_590);
nor U1160 (N_1160,N_567,N_732);
nor U1161 (N_1161,N_974,N_877);
nor U1162 (N_1162,N_944,N_956);
or U1163 (N_1163,N_574,N_734);
xor U1164 (N_1164,N_786,N_946);
nand U1165 (N_1165,N_647,N_861);
nand U1166 (N_1166,N_933,N_813);
nor U1167 (N_1167,N_529,N_581);
xnor U1168 (N_1168,N_907,N_922);
nand U1169 (N_1169,N_749,N_638);
nor U1170 (N_1170,N_639,N_644);
nor U1171 (N_1171,N_752,N_928);
nand U1172 (N_1172,N_502,N_954);
or U1173 (N_1173,N_691,N_539);
nor U1174 (N_1174,N_870,N_927);
and U1175 (N_1175,N_500,N_831);
nand U1176 (N_1176,N_765,N_750);
xnor U1177 (N_1177,N_874,N_896);
or U1178 (N_1178,N_760,N_572);
nor U1179 (N_1179,N_919,N_657);
or U1180 (N_1180,N_561,N_640);
nand U1181 (N_1181,N_710,N_835);
or U1182 (N_1182,N_911,N_865);
xor U1183 (N_1183,N_931,N_976);
xor U1184 (N_1184,N_595,N_901);
and U1185 (N_1185,N_955,N_785);
xnor U1186 (N_1186,N_964,N_653);
xor U1187 (N_1187,N_564,N_711);
nor U1188 (N_1188,N_607,N_925);
or U1189 (N_1189,N_636,N_834);
and U1190 (N_1190,N_703,N_681);
nand U1191 (N_1191,N_555,N_670);
and U1192 (N_1192,N_893,N_709);
and U1193 (N_1193,N_772,N_892);
and U1194 (N_1194,N_878,N_775);
or U1195 (N_1195,N_915,N_612);
xor U1196 (N_1196,N_671,N_782);
nand U1197 (N_1197,N_721,N_712);
and U1198 (N_1198,N_991,N_766);
or U1199 (N_1199,N_957,N_903);
nor U1200 (N_1200,N_661,N_748);
nand U1201 (N_1201,N_620,N_819);
nand U1202 (N_1202,N_702,N_937);
or U1203 (N_1203,N_582,N_583);
and U1204 (N_1204,N_551,N_875);
nand U1205 (N_1205,N_648,N_666);
xnor U1206 (N_1206,N_939,N_741);
and U1207 (N_1207,N_906,N_578);
xnor U1208 (N_1208,N_828,N_596);
xor U1209 (N_1209,N_844,N_656);
nor U1210 (N_1210,N_791,N_884);
xnor U1211 (N_1211,N_696,N_577);
nand U1212 (N_1212,N_771,N_759);
nor U1213 (N_1213,N_687,N_686);
or U1214 (N_1214,N_717,N_795);
or U1215 (N_1215,N_614,N_613);
nand U1216 (N_1216,N_507,N_801);
nor U1217 (N_1217,N_827,N_699);
and U1218 (N_1218,N_804,N_950);
nor U1219 (N_1219,N_953,N_519);
nand U1220 (N_1220,N_684,N_556);
xnor U1221 (N_1221,N_805,N_606);
nand U1222 (N_1222,N_601,N_560);
xor U1223 (N_1223,N_754,N_971);
xnor U1224 (N_1224,N_704,N_783);
nand U1225 (N_1225,N_676,N_655);
and U1226 (N_1226,N_619,N_862);
or U1227 (N_1227,N_858,N_829);
nand U1228 (N_1228,N_511,N_677);
or U1229 (N_1229,N_800,N_961);
or U1230 (N_1230,N_728,N_923);
xor U1231 (N_1231,N_746,N_926);
xor U1232 (N_1232,N_985,N_558);
xor U1233 (N_1233,N_599,N_505);
xor U1234 (N_1234,N_770,N_541);
nand U1235 (N_1235,N_527,N_847);
and U1236 (N_1236,N_952,N_573);
and U1237 (N_1237,N_531,N_535);
or U1238 (N_1238,N_900,N_672);
or U1239 (N_1239,N_718,N_850);
and U1240 (N_1240,N_643,N_975);
nand U1241 (N_1241,N_968,N_914);
or U1242 (N_1242,N_508,N_958);
nor U1243 (N_1243,N_645,N_940);
xor U1244 (N_1244,N_716,N_592);
nand U1245 (N_1245,N_753,N_692);
nor U1246 (N_1246,N_842,N_742);
or U1247 (N_1247,N_747,N_995);
and U1248 (N_1248,N_626,N_700);
and U1249 (N_1249,N_652,N_600);
and U1250 (N_1250,N_612,N_855);
nor U1251 (N_1251,N_933,N_781);
and U1252 (N_1252,N_569,N_691);
nor U1253 (N_1253,N_987,N_572);
nand U1254 (N_1254,N_936,N_536);
and U1255 (N_1255,N_673,N_768);
nand U1256 (N_1256,N_844,N_786);
or U1257 (N_1257,N_663,N_726);
nand U1258 (N_1258,N_797,N_656);
and U1259 (N_1259,N_801,N_809);
nor U1260 (N_1260,N_819,N_999);
nand U1261 (N_1261,N_857,N_940);
nor U1262 (N_1262,N_586,N_849);
and U1263 (N_1263,N_722,N_744);
nand U1264 (N_1264,N_516,N_943);
nor U1265 (N_1265,N_935,N_689);
nor U1266 (N_1266,N_925,N_556);
nand U1267 (N_1267,N_585,N_507);
and U1268 (N_1268,N_728,N_582);
and U1269 (N_1269,N_544,N_972);
nor U1270 (N_1270,N_821,N_740);
and U1271 (N_1271,N_531,N_618);
xnor U1272 (N_1272,N_836,N_841);
nand U1273 (N_1273,N_795,N_699);
or U1274 (N_1274,N_832,N_989);
or U1275 (N_1275,N_593,N_565);
and U1276 (N_1276,N_902,N_921);
and U1277 (N_1277,N_740,N_719);
and U1278 (N_1278,N_598,N_874);
nand U1279 (N_1279,N_814,N_740);
xnor U1280 (N_1280,N_942,N_549);
nor U1281 (N_1281,N_584,N_540);
xnor U1282 (N_1282,N_636,N_810);
or U1283 (N_1283,N_865,N_584);
nand U1284 (N_1284,N_833,N_716);
nand U1285 (N_1285,N_524,N_866);
nand U1286 (N_1286,N_690,N_627);
or U1287 (N_1287,N_744,N_940);
nand U1288 (N_1288,N_643,N_547);
or U1289 (N_1289,N_984,N_610);
xnor U1290 (N_1290,N_997,N_751);
and U1291 (N_1291,N_856,N_826);
nand U1292 (N_1292,N_939,N_545);
nor U1293 (N_1293,N_750,N_594);
nand U1294 (N_1294,N_875,N_501);
and U1295 (N_1295,N_560,N_866);
nor U1296 (N_1296,N_887,N_763);
xor U1297 (N_1297,N_993,N_795);
nand U1298 (N_1298,N_724,N_977);
nor U1299 (N_1299,N_854,N_732);
nor U1300 (N_1300,N_792,N_848);
or U1301 (N_1301,N_607,N_943);
nand U1302 (N_1302,N_786,N_590);
xnor U1303 (N_1303,N_796,N_734);
nand U1304 (N_1304,N_628,N_890);
nand U1305 (N_1305,N_820,N_795);
xor U1306 (N_1306,N_520,N_516);
and U1307 (N_1307,N_629,N_523);
nor U1308 (N_1308,N_504,N_779);
or U1309 (N_1309,N_623,N_543);
and U1310 (N_1310,N_995,N_914);
and U1311 (N_1311,N_657,N_700);
nor U1312 (N_1312,N_620,N_570);
or U1313 (N_1313,N_939,N_759);
xnor U1314 (N_1314,N_742,N_618);
xor U1315 (N_1315,N_699,N_960);
xor U1316 (N_1316,N_794,N_719);
nor U1317 (N_1317,N_892,N_917);
or U1318 (N_1318,N_969,N_924);
or U1319 (N_1319,N_902,N_510);
xnor U1320 (N_1320,N_516,N_710);
and U1321 (N_1321,N_762,N_939);
xor U1322 (N_1322,N_741,N_737);
nand U1323 (N_1323,N_972,N_520);
xor U1324 (N_1324,N_585,N_879);
and U1325 (N_1325,N_507,N_823);
or U1326 (N_1326,N_964,N_597);
nand U1327 (N_1327,N_750,N_525);
xor U1328 (N_1328,N_629,N_506);
xor U1329 (N_1329,N_587,N_674);
and U1330 (N_1330,N_904,N_707);
xor U1331 (N_1331,N_907,N_645);
and U1332 (N_1332,N_549,N_648);
xnor U1333 (N_1333,N_836,N_725);
xnor U1334 (N_1334,N_560,N_899);
nor U1335 (N_1335,N_899,N_774);
nand U1336 (N_1336,N_554,N_670);
or U1337 (N_1337,N_796,N_960);
nand U1338 (N_1338,N_949,N_821);
xnor U1339 (N_1339,N_593,N_798);
nand U1340 (N_1340,N_528,N_906);
or U1341 (N_1341,N_516,N_638);
xnor U1342 (N_1342,N_959,N_886);
and U1343 (N_1343,N_734,N_759);
nand U1344 (N_1344,N_561,N_927);
and U1345 (N_1345,N_921,N_946);
nor U1346 (N_1346,N_863,N_743);
and U1347 (N_1347,N_536,N_990);
or U1348 (N_1348,N_656,N_528);
or U1349 (N_1349,N_988,N_738);
nand U1350 (N_1350,N_511,N_940);
or U1351 (N_1351,N_611,N_996);
nand U1352 (N_1352,N_762,N_524);
xnor U1353 (N_1353,N_788,N_512);
or U1354 (N_1354,N_605,N_925);
nor U1355 (N_1355,N_698,N_818);
or U1356 (N_1356,N_901,N_894);
xor U1357 (N_1357,N_842,N_604);
xor U1358 (N_1358,N_552,N_646);
nand U1359 (N_1359,N_728,N_956);
and U1360 (N_1360,N_682,N_592);
or U1361 (N_1361,N_957,N_901);
nand U1362 (N_1362,N_744,N_658);
or U1363 (N_1363,N_884,N_945);
and U1364 (N_1364,N_643,N_623);
or U1365 (N_1365,N_910,N_734);
and U1366 (N_1366,N_734,N_738);
or U1367 (N_1367,N_526,N_683);
or U1368 (N_1368,N_966,N_651);
nand U1369 (N_1369,N_680,N_975);
nor U1370 (N_1370,N_903,N_555);
and U1371 (N_1371,N_657,N_890);
and U1372 (N_1372,N_900,N_756);
xor U1373 (N_1373,N_930,N_856);
nand U1374 (N_1374,N_544,N_597);
nor U1375 (N_1375,N_676,N_775);
nor U1376 (N_1376,N_682,N_578);
or U1377 (N_1377,N_673,N_725);
or U1378 (N_1378,N_882,N_752);
xnor U1379 (N_1379,N_950,N_686);
nor U1380 (N_1380,N_766,N_647);
xor U1381 (N_1381,N_777,N_670);
nand U1382 (N_1382,N_859,N_607);
or U1383 (N_1383,N_695,N_517);
nand U1384 (N_1384,N_568,N_638);
nand U1385 (N_1385,N_658,N_599);
or U1386 (N_1386,N_576,N_780);
or U1387 (N_1387,N_919,N_777);
and U1388 (N_1388,N_746,N_524);
xnor U1389 (N_1389,N_680,N_967);
or U1390 (N_1390,N_913,N_862);
nand U1391 (N_1391,N_690,N_620);
or U1392 (N_1392,N_782,N_607);
or U1393 (N_1393,N_659,N_814);
and U1394 (N_1394,N_694,N_727);
nor U1395 (N_1395,N_735,N_989);
and U1396 (N_1396,N_645,N_621);
nand U1397 (N_1397,N_614,N_655);
nand U1398 (N_1398,N_860,N_757);
nand U1399 (N_1399,N_788,N_856);
xnor U1400 (N_1400,N_551,N_633);
or U1401 (N_1401,N_791,N_938);
xnor U1402 (N_1402,N_801,N_807);
and U1403 (N_1403,N_937,N_524);
or U1404 (N_1404,N_830,N_593);
and U1405 (N_1405,N_695,N_652);
nor U1406 (N_1406,N_652,N_986);
xor U1407 (N_1407,N_967,N_842);
or U1408 (N_1408,N_509,N_758);
xnor U1409 (N_1409,N_676,N_564);
nor U1410 (N_1410,N_789,N_844);
nor U1411 (N_1411,N_502,N_757);
and U1412 (N_1412,N_533,N_650);
nand U1413 (N_1413,N_890,N_510);
and U1414 (N_1414,N_896,N_958);
or U1415 (N_1415,N_830,N_533);
and U1416 (N_1416,N_782,N_904);
xor U1417 (N_1417,N_580,N_941);
and U1418 (N_1418,N_578,N_716);
and U1419 (N_1419,N_998,N_735);
xnor U1420 (N_1420,N_570,N_699);
or U1421 (N_1421,N_722,N_999);
or U1422 (N_1422,N_704,N_863);
nor U1423 (N_1423,N_952,N_744);
nand U1424 (N_1424,N_955,N_734);
nor U1425 (N_1425,N_625,N_823);
nor U1426 (N_1426,N_500,N_539);
or U1427 (N_1427,N_858,N_552);
nor U1428 (N_1428,N_617,N_637);
and U1429 (N_1429,N_686,N_985);
xnor U1430 (N_1430,N_580,N_574);
and U1431 (N_1431,N_544,N_942);
nand U1432 (N_1432,N_618,N_529);
nand U1433 (N_1433,N_690,N_695);
or U1434 (N_1434,N_571,N_963);
nand U1435 (N_1435,N_848,N_540);
and U1436 (N_1436,N_744,N_626);
and U1437 (N_1437,N_819,N_556);
nand U1438 (N_1438,N_720,N_738);
and U1439 (N_1439,N_626,N_833);
and U1440 (N_1440,N_819,N_939);
and U1441 (N_1441,N_547,N_589);
xnor U1442 (N_1442,N_980,N_765);
and U1443 (N_1443,N_781,N_657);
nor U1444 (N_1444,N_664,N_543);
or U1445 (N_1445,N_845,N_782);
and U1446 (N_1446,N_571,N_734);
nor U1447 (N_1447,N_940,N_864);
and U1448 (N_1448,N_863,N_911);
nor U1449 (N_1449,N_806,N_657);
and U1450 (N_1450,N_649,N_846);
or U1451 (N_1451,N_677,N_560);
nor U1452 (N_1452,N_599,N_982);
and U1453 (N_1453,N_673,N_926);
xnor U1454 (N_1454,N_767,N_674);
xnor U1455 (N_1455,N_552,N_992);
and U1456 (N_1456,N_678,N_908);
or U1457 (N_1457,N_663,N_967);
xnor U1458 (N_1458,N_535,N_676);
xnor U1459 (N_1459,N_556,N_737);
nand U1460 (N_1460,N_576,N_589);
nor U1461 (N_1461,N_908,N_740);
nor U1462 (N_1462,N_620,N_682);
xnor U1463 (N_1463,N_518,N_920);
nor U1464 (N_1464,N_670,N_984);
xnor U1465 (N_1465,N_813,N_834);
nor U1466 (N_1466,N_837,N_943);
nor U1467 (N_1467,N_723,N_579);
and U1468 (N_1468,N_683,N_933);
and U1469 (N_1469,N_684,N_800);
nor U1470 (N_1470,N_890,N_902);
and U1471 (N_1471,N_736,N_650);
nor U1472 (N_1472,N_762,N_842);
xor U1473 (N_1473,N_764,N_745);
nor U1474 (N_1474,N_871,N_821);
or U1475 (N_1475,N_776,N_869);
or U1476 (N_1476,N_547,N_509);
or U1477 (N_1477,N_690,N_944);
nand U1478 (N_1478,N_762,N_647);
or U1479 (N_1479,N_654,N_527);
nor U1480 (N_1480,N_625,N_547);
xor U1481 (N_1481,N_842,N_625);
and U1482 (N_1482,N_714,N_915);
or U1483 (N_1483,N_668,N_632);
or U1484 (N_1484,N_785,N_900);
nor U1485 (N_1485,N_522,N_992);
nor U1486 (N_1486,N_918,N_598);
nand U1487 (N_1487,N_552,N_882);
nand U1488 (N_1488,N_615,N_531);
and U1489 (N_1489,N_814,N_569);
nand U1490 (N_1490,N_752,N_750);
or U1491 (N_1491,N_896,N_742);
and U1492 (N_1492,N_693,N_781);
nand U1493 (N_1493,N_790,N_525);
and U1494 (N_1494,N_635,N_685);
nand U1495 (N_1495,N_882,N_984);
nor U1496 (N_1496,N_866,N_887);
nor U1497 (N_1497,N_633,N_803);
nand U1498 (N_1498,N_949,N_780);
xor U1499 (N_1499,N_778,N_813);
and U1500 (N_1500,N_1417,N_1251);
xor U1501 (N_1501,N_1302,N_1045);
nand U1502 (N_1502,N_1370,N_1361);
nor U1503 (N_1503,N_1062,N_1365);
nor U1504 (N_1504,N_1039,N_1077);
and U1505 (N_1505,N_1168,N_1495);
nor U1506 (N_1506,N_1400,N_1221);
nor U1507 (N_1507,N_1002,N_1223);
nor U1508 (N_1508,N_1281,N_1179);
xnor U1509 (N_1509,N_1430,N_1473);
nor U1510 (N_1510,N_1029,N_1125);
nor U1511 (N_1511,N_1363,N_1023);
nand U1512 (N_1512,N_1409,N_1012);
or U1513 (N_1513,N_1323,N_1314);
and U1514 (N_1514,N_1332,N_1118);
xor U1515 (N_1515,N_1494,N_1044);
xor U1516 (N_1516,N_1170,N_1060);
nand U1517 (N_1517,N_1153,N_1327);
nand U1518 (N_1518,N_1340,N_1064);
nand U1519 (N_1519,N_1116,N_1386);
nor U1520 (N_1520,N_1229,N_1268);
xnor U1521 (N_1521,N_1097,N_1075);
nand U1522 (N_1522,N_1291,N_1066);
and U1523 (N_1523,N_1283,N_1033);
or U1524 (N_1524,N_1198,N_1219);
xnor U1525 (N_1525,N_1000,N_1040);
and U1526 (N_1526,N_1067,N_1286);
nor U1527 (N_1527,N_1137,N_1277);
or U1528 (N_1528,N_1159,N_1036);
nand U1529 (N_1529,N_1249,N_1150);
nand U1530 (N_1530,N_1047,N_1011);
or U1531 (N_1531,N_1015,N_1177);
xor U1532 (N_1532,N_1467,N_1089);
xnor U1533 (N_1533,N_1114,N_1124);
or U1534 (N_1534,N_1410,N_1138);
nor U1535 (N_1535,N_1256,N_1439);
nand U1536 (N_1536,N_1050,N_1109);
and U1537 (N_1537,N_1433,N_1393);
nand U1538 (N_1538,N_1214,N_1376);
or U1539 (N_1539,N_1207,N_1476);
xor U1540 (N_1540,N_1041,N_1282);
xnor U1541 (N_1541,N_1018,N_1427);
nand U1542 (N_1542,N_1173,N_1257);
nand U1543 (N_1543,N_1184,N_1227);
xor U1544 (N_1544,N_1485,N_1298);
xnor U1545 (N_1545,N_1343,N_1127);
and U1546 (N_1546,N_1329,N_1461);
or U1547 (N_1547,N_1341,N_1022);
or U1548 (N_1548,N_1311,N_1348);
nand U1549 (N_1549,N_1247,N_1452);
or U1550 (N_1550,N_1450,N_1358);
nand U1551 (N_1551,N_1471,N_1217);
nand U1552 (N_1552,N_1081,N_1154);
and U1553 (N_1553,N_1420,N_1068);
xnor U1554 (N_1554,N_1253,N_1474);
xnor U1555 (N_1555,N_1367,N_1328);
or U1556 (N_1556,N_1233,N_1026);
xnor U1557 (N_1557,N_1339,N_1218);
nand U1558 (N_1558,N_1470,N_1063);
xor U1559 (N_1559,N_1305,N_1468);
or U1560 (N_1560,N_1111,N_1438);
xnor U1561 (N_1561,N_1028,N_1103);
and U1562 (N_1562,N_1375,N_1083);
nand U1563 (N_1563,N_1326,N_1280);
nor U1564 (N_1564,N_1398,N_1160);
xor U1565 (N_1565,N_1196,N_1053);
nand U1566 (N_1566,N_1491,N_1422);
nand U1567 (N_1567,N_1415,N_1108);
nand U1568 (N_1568,N_1458,N_1180);
nor U1569 (N_1569,N_1086,N_1372);
nand U1570 (N_1570,N_1402,N_1105);
nand U1571 (N_1571,N_1082,N_1020);
or U1572 (N_1572,N_1278,N_1483);
nand U1573 (N_1573,N_1324,N_1297);
xnor U1574 (N_1574,N_1264,N_1009);
xnor U1575 (N_1575,N_1142,N_1197);
nor U1576 (N_1576,N_1013,N_1164);
and U1577 (N_1577,N_1239,N_1094);
nor U1578 (N_1578,N_1019,N_1455);
and U1579 (N_1579,N_1299,N_1122);
xnor U1580 (N_1580,N_1448,N_1371);
xor U1581 (N_1581,N_1065,N_1454);
nand U1582 (N_1582,N_1027,N_1321);
nand U1583 (N_1583,N_1352,N_1319);
and U1584 (N_1584,N_1073,N_1465);
and U1585 (N_1585,N_1347,N_1405);
and U1586 (N_1586,N_1046,N_1148);
xor U1587 (N_1587,N_1443,N_1007);
and U1588 (N_1588,N_1203,N_1300);
xnor U1589 (N_1589,N_1078,N_1354);
or U1590 (N_1590,N_1133,N_1385);
nand U1591 (N_1591,N_1317,N_1056);
and U1592 (N_1592,N_1155,N_1434);
xor U1593 (N_1593,N_1206,N_1342);
or U1594 (N_1594,N_1313,N_1143);
xor U1595 (N_1595,N_1397,N_1374);
xor U1596 (N_1596,N_1295,N_1355);
and U1597 (N_1597,N_1051,N_1091);
and U1598 (N_1598,N_1241,N_1388);
or U1599 (N_1599,N_1212,N_1230);
or U1600 (N_1600,N_1346,N_1185);
nand U1601 (N_1601,N_1453,N_1364);
and U1602 (N_1602,N_1378,N_1382);
or U1603 (N_1603,N_1472,N_1188);
and U1604 (N_1604,N_1449,N_1176);
xnor U1605 (N_1605,N_1131,N_1413);
or U1606 (N_1606,N_1306,N_1416);
and U1607 (N_1607,N_1182,N_1093);
xnor U1608 (N_1608,N_1098,N_1403);
and U1609 (N_1609,N_1254,N_1071);
and U1610 (N_1610,N_1165,N_1469);
xor U1611 (N_1611,N_1404,N_1487);
and U1612 (N_1612,N_1336,N_1310);
nand U1613 (N_1613,N_1238,N_1240);
or U1614 (N_1614,N_1059,N_1477);
nor U1615 (N_1615,N_1231,N_1130);
or U1616 (N_1616,N_1345,N_1090);
nor U1617 (N_1617,N_1481,N_1187);
or U1618 (N_1618,N_1004,N_1200);
nor U1619 (N_1619,N_1243,N_1301);
xor U1620 (N_1620,N_1399,N_1178);
and U1621 (N_1621,N_1003,N_1480);
or U1622 (N_1622,N_1259,N_1275);
nand U1623 (N_1623,N_1102,N_1478);
nand U1624 (N_1624,N_1145,N_1429);
nand U1625 (N_1625,N_1335,N_1161);
and U1626 (N_1626,N_1419,N_1442);
or U1627 (N_1627,N_1387,N_1368);
nor U1628 (N_1628,N_1293,N_1423);
xor U1629 (N_1629,N_1331,N_1204);
nand U1630 (N_1630,N_1392,N_1054);
and U1631 (N_1631,N_1333,N_1010);
nand U1632 (N_1632,N_1279,N_1369);
nand U1633 (N_1633,N_1014,N_1172);
xor U1634 (N_1634,N_1266,N_1107);
nand U1635 (N_1635,N_1490,N_1437);
and U1636 (N_1636,N_1421,N_1016);
and U1637 (N_1637,N_1072,N_1175);
and U1638 (N_1638,N_1289,N_1296);
nand U1639 (N_1639,N_1194,N_1149);
xnor U1640 (N_1640,N_1303,N_1445);
or U1641 (N_1641,N_1447,N_1391);
nand U1642 (N_1642,N_1273,N_1245);
nor U1643 (N_1643,N_1163,N_1489);
nor U1644 (N_1644,N_1113,N_1048);
nand U1645 (N_1645,N_1106,N_1158);
and U1646 (N_1646,N_1463,N_1167);
or U1647 (N_1647,N_1407,N_1287);
and U1648 (N_1648,N_1373,N_1267);
nor U1649 (N_1649,N_1425,N_1320);
nand U1650 (N_1650,N_1244,N_1104);
and U1651 (N_1651,N_1250,N_1436);
or U1652 (N_1652,N_1205,N_1304);
nand U1653 (N_1653,N_1294,N_1353);
nand U1654 (N_1654,N_1069,N_1290);
or U1655 (N_1655,N_1129,N_1431);
nand U1656 (N_1656,N_1276,N_1112);
nand U1657 (N_1657,N_1209,N_1088);
xor U1658 (N_1658,N_1096,N_1265);
nor U1659 (N_1659,N_1488,N_1351);
or U1660 (N_1660,N_1284,N_1460);
and U1661 (N_1661,N_1162,N_1008);
nand U1662 (N_1662,N_1191,N_1043);
or U1663 (N_1663,N_1035,N_1190);
xor U1664 (N_1664,N_1315,N_1322);
and U1665 (N_1665,N_1144,N_1457);
nand U1666 (N_1666,N_1390,N_1334);
xor U1667 (N_1667,N_1225,N_1151);
xor U1668 (N_1668,N_1213,N_1192);
xor U1669 (N_1669,N_1414,N_1349);
nand U1670 (N_1670,N_1424,N_1312);
nand U1671 (N_1671,N_1139,N_1366);
nor U1672 (N_1672,N_1236,N_1171);
nand U1673 (N_1673,N_1497,N_1484);
and U1674 (N_1674,N_1237,N_1486);
xor U1675 (N_1675,N_1132,N_1379);
or U1676 (N_1676,N_1479,N_1441);
nand U1677 (N_1677,N_1255,N_1406);
and U1678 (N_1678,N_1377,N_1202);
nand U1679 (N_1679,N_1380,N_1117);
xor U1680 (N_1680,N_1032,N_1271);
or U1681 (N_1681,N_1232,N_1136);
xor U1682 (N_1682,N_1030,N_1201);
nand U1683 (N_1683,N_1493,N_1252);
and U1684 (N_1684,N_1100,N_1226);
nand U1685 (N_1685,N_1262,N_1087);
nor U1686 (N_1686,N_1466,N_1459);
nand U1687 (N_1687,N_1288,N_1498);
nor U1688 (N_1688,N_1181,N_1263);
nor U1689 (N_1689,N_1099,N_1055);
xnor U1690 (N_1690,N_1381,N_1005);
nor U1691 (N_1691,N_1356,N_1061);
nor U1692 (N_1692,N_1070,N_1384);
nor U1693 (N_1693,N_1195,N_1146);
nand U1694 (N_1694,N_1189,N_1076);
xor U1695 (N_1695,N_1383,N_1049);
xor U1696 (N_1696,N_1446,N_1318);
or U1697 (N_1697,N_1084,N_1101);
or U1698 (N_1698,N_1496,N_1186);
or U1699 (N_1699,N_1428,N_1057);
or U1700 (N_1700,N_1412,N_1440);
nand U1701 (N_1701,N_1344,N_1408);
nor U1702 (N_1702,N_1126,N_1215);
and U1703 (N_1703,N_1147,N_1292);
nand U1704 (N_1704,N_1174,N_1031);
nand U1705 (N_1705,N_1169,N_1362);
nand U1706 (N_1706,N_1451,N_1435);
or U1707 (N_1707,N_1222,N_1258);
xnor U1708 (N_1708,N_1492,N_1135);
nand U1709 (N_1709,N_1156,N_1128);
or U1710 (N_1710,N_1309,N_1034);
nand U1711 (N_1711,N_1183,N_1432);
xor U1712 (N_1712,N_1074,N_1316);
nand U1713 (N_1713,N_1134,N_1396);
or U1714 (N_1714,N_1462,N_1401);
and U1715 (N_1715,N_1079,N_1359);
nor U1716 (N_1716,N_1193,N_1017);
xnor U1717 (N_1717,N_1270,N_1330);
xor U1718 (N_1718,N_1001,N_1025);
and U1719 (N_1719,N_1456,N_1260);
nor U1720 (N_1720,N_1394,N_1261);
nand U1721 (N_1721,N_1308,N_1199);
or U1722 (N_1722,N_1325,N_1085);
and U1723 (N_1723,N_1121,N_1285);
or U1724 (N_1724,N_1357,N_1208);
xnor U1725 (N_1725,N_1152,N_1338);
or U1726 (N_1726,N_1499,N_1140);
nor U1727 (N_1727,N_1235,N_1120);
xnor U1728 (N_1728,N_1037,N_1272);
and U1729 (N_1729,N_1006,N_1210);
nor U1730 (N_1730,N_1242,N_1350);
nand U1731 (N_1731,N_1080,N_1123);
nor U1732 (N_1732,N_1411,N_1475);
nor U1733 (N_1733,N_1274,N_1058);
nor U1734 (N_1734,N_1110,N_1092);
or U1735 (N_1735,N_1444,N_1464);
nor U1736 (N_1736,N_1119,N_1166);
nand U1737 (N_1737,N_1095,N_1042);
and U1738 (N_1738,N_1269,N_1307);
and U1739 (N_1739,N_1052,N_1360);
or U1740 (N_1740,N_1395,N_1211);
and U1741 (N_1741,N_1248,N_1021);
nor U1742 (N_1742,N_1228,N_1141);
nor U1743 (N_1743,N_1426,N_1115);
or U1744 (N_1744,N_1389,N_1418);
and U1745 (N_1745,N_1224,N_1038);
xnor U1746 (N_1746,N_1246,N_1482);
or U1747 (N_1747,N_1337,N_1220);
nor U1748 (N_1748,N_1216,N_1024);
nor U1749 (N_1749,N_1157,N_1234);
nand U1750 (N_1750,N_1157,N_1402);
nor U1751 (N_1751,N_1066,N_1024);
and U1752 (N_1752,N_1176,N_1025);
or U1753 (N_1753,N_1306,N_1209);
and U1754 (N_1754,N_1062,N_1339);
xor U1755 (N_1755,N_1048,N_1262);
nor U1756 (N_1756,N_1046,N_1487);
nand U1757 (N_1757,N_1206,N_1332);
nor U1758 (N_1758,N_1349,N_1231);
nor U1759 (N_1759,N_1423,N_1040);
and U1760 (N_1760,N_1430,N_1248);
or U1761 (N_1761,N_1032,N_1150);
nand U1762 (N_1762,N_1014,N_1070);
nor U1763 (N_1763,N_1341,N_1272);
nand U1764 (N_1764,N_1365,N_1352);
nor U1765 (N_1765,N_1464,N_1468);
and U1766 (N_1766,N_1180,N_1425);
nor U1767 (N_1767,N_1254,N_1180);
or U1768 (N_1768,N_1452,N_1099);
xnor U1769 (N_1769,N_1269,N_1209);
nor U1770 (N_1770,N_1368,N_1149);
nand U1771 (N_1771,N_1036,N_1262);
nand U1772 (N_1772,N_1248,N_1374);
xnor U1773 (N_1773,N_1072,N_1153);
or U1774 (N_1774,N_1008,N_1390);
nor U1775 (N_1775,N_1461,N_1321);
or U1776 (N_1776,N_1188,N_1322);
nor U1777 (N_1777,N_1054,N_1104);
or U1778 (N_1778,N_1487,N_1472);
nor U1779 (N_1779,N_1003,N_1301);
and U1780 (N_1780,N_1161,N_1449);
or U1781 (N_1781,N_1341,N_1355);
or U1782 (N_1782,N_1277,N_1009);
nor U1783 (N_1783,N_1296,N_1060);
nor U1784 (N_1784,N_1473,N_1151);
xor U1785 (N_1785,N_1263,N_1222);
nor U1786 (N_1786,N_1401,N_1343);
or U1787 (N_1787,N_1474,N_1089);
xor U1788 (N_1788,N_1260,N_1067);
or U1789 (N_1789,N_1406,N_1002);
xnor U1790 (N_1790,N_1304,N_1252);
nand U1791 (N_1791,N_1215,N_1227);
nand U1792 (N_1792,N_1137,N_1059);
nand U1793 (N_1793,N_1395,N_1086);
and U1794 (N_1794,N_1398,N_1381);
xor U1795 (N_1795,N_1181,N_1020);
and U1796 (N_1796,N_1280,N_1293);
nand U1797 (N_1797,N_1044,N_1308);
and U1798 (N_1798,N_1077,N_1142);
nand U1799 (N_1799,N_1210,N_1455);
nor U1800 (N_1800,N_1259,N_1341);
xnor U1801 (N_1801,N_1230,N_1341);
nor U1802 (N_1802,N_1169,N_1419);
xor U1803 (N_1803,N_1457,N_1385);
nand U1804 (N_1804,N_1324,N_1173);
and U1805 (N_1805,N_1221,N_1186);
nor U1806 (N_1806,N_1326,N_1053);
nand U1807 (N_1807,N_1408,N_1366);
xor U1808 (N_1808,N_1336,N_1237);
nor U1809 (N_1809,N_1260,N_1228);
nor U1810 (N_1810,N_1435,N_1130);
or U1811 (N_1811,N_1126,N_1324);
nor U1812 (N_1812,N_1222,N_1038);
nor U1813 (N_1813,N_1179,N_1180);
nand U1814 (N_1814,N_1105,N_1244);
nor U1815 (N_1815,N_1298,N_1206);
or U1816 (N_1816,N_1279,N_1345);
nand U1817 (N_1817,N_1288,N_1109);
nor U1818 (N_1818,N_1061,N_1296);
xor U1819 (N_1819,N_1038,N_1269);
xnor U1820 (N_1820,N_1188,N_1386);
and U1821 (N_1821,N_1479,N_1317);
nor U1822 (N_1822,N_1360,N_1287);
and U1823 (N_1823,N_1143,N_1311);
and U1824 (N_1824,N_1196,N_1211);
nand U1825 (N_1825,N_1468,N_1202);
nand U1826 (N_1826,N_1381,N_1034);
or U1827 (N_1827,N_1473,N_1196);
nor U1828 (N_1828,N_1454,N_1003);
nor U1829 (N_1829,N_1114,N_1300);
nor U1830 (N_1830,N_1164,N_1081);
xor U1831 (N_1831,N_1244,N_1238);
nor U1832 (N_1832,N_1372,N_1004);
nand U1833 (N_1833,N_1042,N_1162);
xnor U1834 (N_1834,N_1381,N_1302);
xor U1835 (N_1835,N_1030,N_1268);
and U1836 (N_1836,N_1431,N_1077);
xnor U1837 (N_1837,N_1368,N_1066);
and U1838 (N_1838,N_1036,N_1268);
xnor U1839 (N_1839,N_1339,N_1497);
nor U1840 (N_1840,N_1181,N_1426);
nand U1841 (N_1841,N_1326,N_1095);
xor U1842 (N_1842,N_1273,N_1188);
or U1843 (N_1843,N_1182,N_1340);
or U1844 (N_1844,N_1475,N_1158);
nand U1845 (N_1845,N_1172,N_1195);
nor U1846 (N_1846,N_1342,N_1062);
nand U1847 (N_1847,N_1048,N_1477);
or U1848 (N_1848,N_1079,N_1463);
and U1849 (N_1849,N_1214,N_1367);
nor U1850 (N_1850,N_1243,N_1078);
nor U1851 (N_1851,N_1465,N_1243);
nand U1852 (N_1852,N_1235,N_1076);
nor U1853 (N_1853,N_1280,N_1416);
and U1854 (N_1854,N_1045,N_1464);
or U1855 (N_1855,N_1149,N_1127);
or U1856 (N_1856,N_1382,N_1274);
nand U1857 (N_1857,N_1058,N_1259);
and U1858 (N_1858,N_1437,N_1081);
nor U1859 (N_1859,N_1246,N_1302);
nor U1860 (N_1860,N_1211,N_1436);
and U1861 (N_1861,N_1180,N_1205);
xor U1862 (N_1862,N_1460,N_1432);
or U1863 (N_1863,N_1297,N_1044);
and U1864 (N_1864,N_1101,N_1453);
xor U1865 (N_1865,N_1412,N_1318);
nor U1866 (N_1866,N_1039,N_1203);
nand U1867 (N_1867,N_1431,N_1229);
xnor U1868 (N_1868,N_1203,N_1241);
nor U1869 (N_1869,N_1053,N_1199);
or U1870 (N_1870,N_1238,N_1021);
nor U1871 (N_1871,N_1474,N_1076);
xnor U1872 (N_1872,N_1024,N_1497);
and U1873 (N_1873,N_1435,N_1452);
xnor U1874 (N_1874,N_1017,N_1384);
or U1875 (N_1875,N_1079,N_1107);
and U1876 (N_1876,N_1048,N_1187);
or U1877 (N_1877,N_1251,N_1270);
xor U1878 (N_1878,N_1451,N_1393);
and U1879 (N_1879,N_1149,N_1005);
xor U1880 (N_1880,N_1493,N_1042);
and U1881 (N_1881,N_1315,N_1000);
xnor U1882 (N_1882,N_1143,N_1340);
or U1883 (N_1883,N_1075,N_1247);
nand U1884 (N_1884,N_1318,N_1007);
and U1885 (N_1885,N_1146,N_1445);
xor U1886 (N_1886,N_1072,N_1226);
nand U1887 (N_1887,N_1077,N_1239);
or U1888 (N_1888,N_1449,N_1004);
or U1889 (N_1889,N_1222,N_1243);
xnor U1890 (N_1890,N_1055,N_1293);
nor U1891 (N_1891,N_1403,N_1384);
and U1892 (N_1892,N_1350,N_1136);
nand U1893 (N_1893,N_1259,N_1007);
and U1894 (N_1894,N_1156,N_1164);
nand U1895 (N_1895,N_1368,N_1352);
xnor U1896 (N_1896,N_1297,N_1254);
or U1897 (N_1897,N_1024,N_1087);
nand U1898 (N_1898,N_1398,N_1217);
nor U1899 (N_1899,N_1489,N_1383);
and U1900 (N_1900,N_1403,N_1422);
or U1901 (N_1901,N_1210,N_1291);
and U1902 (N_1902,N_1449,N_1078);
nand U1903 (N_1903,N_1353,N_1378);
nor U1904 (N_1904,N_1112,N_1132);
nand U1905 (N_1905,N_1429,N_1427);
or U1906 (N_1906,N_1109,N_1148);
and U1907 (N_1907,N_1305,N_1425);
nand U1908 (N_1908,N_1444,N_1109);
or U1909 (N_1909,N_1043,N_1246);
nand U1910 (N_1910,N_1026,N_1327);
nand U1911 (N_1911,N_1462,N_1446);
or U1912 (N_1912,N_1403,N_1381);
nor U1913 (N_1913,N_1368,N_1385);
nor U1914 (N_1914,N_1203,N_1106);
nand U1915 (N_1915,N_1172,N_1029);
nor U1916 (N_1916,N_1055,N_1034);
nor U1917 (N_1917,N_1274,N_1423);
and U1918 (N_1918,N_1144,N_1400);
or U1919 (N_1919,N_1067,N_1464);
and U1920 (N_1920,N_1405,N_1062);
and U1921 (N_1921,N_1470,N_1071);
or U1922 (N_1922,N_1272,N_1120);
nand U1923 (N_1923,N_1000,N_1048);
nor U1924 (N_1924,N_1347,N_1465);
and U1925 (N_1925,N_1261,N_1405);
xnor U1926 (N_1926,N_1427,N_1466);
xnor U1927 (N_1927,N_1044,N_1336);
nor U1928 (N_1928,N_1464,N_1185);
nand U1929 (N_1929,N_1003,N_1451);
nand U1930 (N_1930,N_1075,N_1248);
nor U1931 (N_1931,N_1049,N_1089);
or U1932 (N_1932,N_1017,N_1008);
and U1933 (N_1933,N_1324,N_1444);
or U1934 (N_1934,N_1207,N_1347);
or U1935 (N_1935,N_1029,N_1193);
and U1936 (N_1936,N_1476,N_1346);
xor U1937 (N_1937,N_1372,N_1043);
or U1938 (N_1938,N_1342,N_1249);
nand U1939 (N_1939,N_1315,N_1134);
xor U1940 (N_1940,N_1122,N_1484);
nand U1941 (N_1941,N_1138,N_1003);
nor U1942 (N_1942,N_1311,N_1448);
and U1943 (N_1943,N_1245,N_1142);
xor U1944 (N_1944,N_1380,N_1048);
or U1945 (N_1945,N_1490,N_1336);
nand U1946 (N_1946,N_1206,N_1145);
nand U1947 (N_1947,N_1054,N_1238);
xnor U1948 (N_1948,N_1407,N_1457);
nand U1949 (N_1949,N_1226,N_1207);
or U1950 (N_1950,N_1383,N_1263);
or U1951 (N_1951,N_1374,N_1268);
nor U1952 (N_1952,N_1386,N_1076);
xnor U1953 (N_1953,N_1246,N_1171);
or U1954 (N_1954,N_1268,N_1465);
nand U1955 (N_1955,N_1325,N_1408);
and U1956 (N_1956,N_1318,N_1298);
nor U1957 (N_1957,N_1421,N_1376);
nand U1958 (N_1958,N_1050,N_1418);
nand U1959 (N_1959,N_1047,N_1105);
and U1960 (N_1960,N_1273,N_1103);
nand U1961 (N_1961,N_1435,N_1179);
or U1962 (N_1962,N_1325,N_1130);
nand U1963 (N_1963,N_1376,N_1107);
nor U1964 (N_1964,N_1316,N_1428);
nor U1965 (N_1965,N_1377,N_1337);
nor U1966 (N_1966,N_1386,N_1448);
and U1967 (N_1967,N_1112,N_1415);
and U1968 (N_1968,N_1249,N_1270);
nand U1969 (N_1969,N_1095,N_1045);
and U1970 (N_1970,N_1082,N_1060);
xnor U1971 (N_1971,N_1229,N_1321);
and U1972 (N_1972,N_1349,N_1288);
xor U1973 (N_1973,N_1326,N_1232);
nor U1974 (N_1974,N_1193,N_1370);
nor U1975 (N_1975,N_1344,N_1323);
xor U1976 (N_1976,N_1404,N_1206);
nand U1977 (N_1977,N_1343,N_1009);
or U1978 (N_1978,N_1122,N_1259);
or U1979 (N_1979,N_1383,N_1152);
xnor U1980 (N_1980,N_1384,N_1046);
xor U1981 (N_1981,N_1304,N_1381);
or U1982 (N_1982,N_1350,N_1458);
nand U1983 (N_1983,N_1214,N_1263);
and U1984 (N_1984,N_1445,N_1008);
xor U1985 (N_1985,N_1157,N_1498);
and U1986 (N_1986,N_1261,N_1192);
xor U1987 (N_1987,N_1026,N_1253);
xor U1988 (N_1988,N_1290,N_1487);
or U1989 (N_1989,N_1188,N_1081);
nor U1990 (N_1990,N_1194,N_1291);
and U1991 (N_1991,N_1471,N_1029);
or U1992 (N_1992,N_1432,N_1132);
or U1993 (N_1993,N_1389,N_1416);
and U1994 (N_1994,N_1283,N_1318);
nand U1995 (N_1995,N_1037,N_1283);
or U1996 (N_1996,N_1459,N_1077);
xor U1997 (N_1997,N_1297,N_1213);
and U1998 (N_1998,N_1406,N_1182);
xor U1999 (N_1999,N_1468,N_1097);
nand U2000 (N_2000,N_1578,N_1917);
nor U2001 (N_2001,N_1531,N_1563);
or U2002 (N_2002,N_1700,N_1637);
xnor U2003 (N_2003,N_1799,N_1989);
nor U2004 (N_2004,N_1510,N_1522);
nand U2005 (N_2005,N_1733,N_1675);
and U2006 (N_2006,N_1652,N_1624);
or U2007 (N_2007,N_1604,N_1940);
and U2008 (N_2008,N_1718,N_1667);
nor U2009 (N_2009,N_1504,N_1841);
xnor U2010 (N_2010,N_1528,N_1539);
xor U2011 (N_2011,N_1757,N_1827);
nand U2012 (N_2012,N_1872,N_1862);
or U2013 (N_2013,N_1782,N_1889);
xnor U2014 (N_2014,N_1607,N_1612);
nor U2015 (N_2015,N_1664,N_1959);
or U2016 (N_2016,N_1876,N_1738);
and U2017 (N_2017,N_1899,N_1630);
nor U2018 (N_2018,N_1979,N_1880);
or U2019 (N_2019,N_1534,N_1680);
and U2020 (N_2020,N_1789,N_1756);
xor U2021 (N_2021,N_1987,N_1893);
nor U2022 (N_2022,N_1603,N_1566);
and U2023 (N_2023,N_1611,N_1857);
or U2024 (N_2024,N_1980,N_1809);
and U2025 (N_2025,N_1994,N_1649);
xnor U2026 (N_2026,N_1523,N_1546);
nand U2027 (N_2027,N_1844,N_1918);
xnor U2028 (N_2028,N_1877,N_1598);
nand U2029 (N_2029,N_1927,N_1693);
and U2030 (N_2030,N_1725,N_1960);
xor U2031 (N_2031,N_1930,N_1867);
and U2032 (N_2032,N_1922,N_1670);
or U2033 (N_2033,N_1541,N_1682);
xor U2034 (N_2034,N_1879,N_1606);
nand U2035 (N_2035,N_1507,N_1749);
nand U2036 (N_2036,N_1750,N_1813);
and U2037 (N_2037,N_1661,N_1894);
nor U2038 (N_2038,N_1593,N_1945);
nor U2039 (N_2039,N_1638,N_1571);
nand U2040 (N_2040,N_1996,N_1509);
nand U2041 (N_2041,N_1558,N_1990);
nor U2042 (N_2042,N_1678,N_1622);
nor U2043 (N_2043,N_1676,N_1748);
nand U2044 (N_2044,N_1764,N_1503);
nand U2045 (N_2045,N_1714,N_1596);
nand U2046 (N_2046,N_1708,N_1586);
nor U2047 (N_2047,N_1790,N_1795);
nand U2048 (N_2048,N_1920,N_1646);
nor U2049 (N_2049,N_1852,N_1778);
nor U2050 (N_2050,N_1803,N_1962);
xnor U2051 (N_2051,N_1856,N_1614);
nand U2052 (N_2052,N_1936,N_1697);
nor U2053 (N_2053,N_1819,N_1660);
nand U2054 (N_2054,N_1845,N_1814);
xnor U2055 (N_2055,N_1527,N_1617);
and U2056 (N_2056,N_1999,N_1555);
nand U2057 (N_2057,N_1768,N_1535);
nor U2058 (N_2058,N_1974,N_1903);
xnor U2059 (N_2059,N_1923,N_1842);
xnor U2060 (N_2060,N_1836,N_1734);
nor U2061 (N_2061,N_1839,N_1570);
nor U2062 (N_2062,N_1835,N_1643);
xnor U2063 (N_2063,N_1952,N_1538);
xnor U2064 (N_2064,N_1763,N_1656);
or U2065 (N_2065,N_1723,N_1948);
nor U2066 (N_2066,N_1694,N_1984);
nor U2067 (N_2067,N_1545,N_1548);
nand U2068 (N_2068,N_1702,N_1673);
nor U2069 (N_2069,N_1627,N_1797);
or U2070 (N_2070,N_1978,N_1964);
and U2071 (N_2071,N_1710,N_1619);
and U2072 (N_2072,N_1559,N_1901);
xnor U2073 (N_2073,N_1919,N_1726);
nor U2074 (N_2074,N_1599,N_1873);
xnor U2075 (N_2075,N_1791,N_1513);
nor U2076 (N_2076,N_1552,N_1542);
and U2077 (N_2077,N_1985,N_1746);
or U2078 (N_2078,N_1991,N_1776);
xnor U2079 (N_2079,N_1736,N_1592);
nor U2080 (N_2080,N_1701,N_1843);
xor U2081 (N_2081,N_1665,N_1977);
or U2082 (N_2082,N_1932,N_1585);
xor U2083 (N_2083,N_1674,N_1743);
nand U2084 (N_2084,N_1671,N_1762);
xor U2085 (N_2085,N_1773,N_1618);
or U2086 (N_2086,N_1956,N_1672);
or U2087 (N_2087,N_1519,N_1864);
and U2088 (N_2088,N_1645,N_1698);
and U2089 (N_2089,N_1500,N_1657);
nor U2090 (N_2090,N_1760,N_1937);
or U2091 (N_2091,N_1629,N_1915);
and U2092 (N_2092,N_1863,N_1849);
nand U2093 (N_2093,N_1755,N_1635);
nand U2094 (N_2094,N_1717,N_1870);
nor U2095 (N_2095,N_1998,N_1742);
nor U2096 (N_2096,N_1730,N_1754);
and U2097 (N_2097,N_1691,N_1692);
and U2098 (N_2098,N_1982,N_1777);
nand U2099 (N_2099,N_1897,N_1679);
xor U2100 (N_2100,N_1514,N_1866);
xnor U2101 (N_2101,N_1632,N_1851);
or U2102 (N_2102,N_1800,N_1944);
or U2103 (N_2103,N_1560,N_1972);
xnor U2104 (N_2104,N_1688,N_1641);
and U2105 (N_2105,N_1788,N_1767);
nor U2106 (N_2106,N_1798,N_1957);
and U2107 (N_2107,N_1724,N_1687);
or U2108 (N_2108,N_1949,N_1621);
and U2109 (N_2109,N_1533,N_1881);
nor U2110 (N_2110,N_1955,N_1690);
nand U2111 (N_2111,N_1838,N_1913);
nor U2112 (N_2112,N_1954,N_1860);
nor U2113 (N_2113,N_1822,N_1703);
and U2114 (N_2114,N_1713,N_1905);
nand U2115 (N_2115,N_1931,N_1943);
or U2116 (N_2116,N_1547,N_1771);
and U2117 (N_2117,N_1651,N_1644);
xnor U2118 (N_2118,N_1829,N_1885);
and U2119 (N_2119,N_1544,N_1628);
and U2120 (N_2120,N_1647,N_1909);
or U2121 (N_2121,N_1616,N_1769);
xor U2122 (N_2122,N_1961,N_1737);
nor U2123 (N_2123,N_1731,N_1983);
nand U2124 (N_2124,N_1938,N_1766);
nor U2125 (N_2125,N_1820,N_1640);
xnor U2126 (N_2126,N_1779,N_1825);
or U2127 (N_2127,N_1847,N_1796);
nor U2128 (N_2128,N_1793,N_1569);
nand U2129 (N_2129,N_1659,N_1868);
or U2130 (N_2130,N_1941,N_1993);
xnor U2131 (N_2131,N_1840,N_1902);
or U2132 (N_2132,N_1580,N_1556);
xnor U2133 (N_2133,N_1761,N_1615);
and U2134 (N_2134,N_1988,N_1804);
and U2135 (N_2135,N_1506,N_1869);
nand U2136 (N_2136,N_1830,N_1705);
nor U2137 (N_2137,N_1662,N_1582);
or U2138 (N_2138,N_1719,N_1950);
xor U2139 (N_2139,N_1521,N_1807);
or U2140 (N_2140,N_1890,N_1878);
and U2141 (N_2141,N_1741,N_1565);
nor U2142 (N_2142,N_1516,N_1883);
nand U2143 (N_2143,N_1589,N_1801);
or U2144 (N_2144,N_1967,N_1871);
nor U2145 (N_2145,N_1668,N_1861);
and U2146 (N_2146,N_1554,N_1543);
and U2147 (N_2147,N_1526,N_1914);
nand U2148 (N_2148,N_1655,N_1981);
and U2149 (N_2149,N_1574,N_1610);
nand U2150 (N_2150,N_1910,N_1939);
and U2151 (N_2151,N_1787,N_1728);
nand U2152 (N_2152,N_1634,N_1933);
and U2153 (N_2153,N_1564,N_1530);
and U2154 (N_2154,N_1898,N_1745);
nor U2155 (N_2155,N_1576,N_1770);
xor U2156 (N_2156,N_1720,N_1744);
or U2157 (N_2157,N_1602,N_1826);
nand U2158 (N_2158,N_1966,N_1740);
or U2159 (N_2159,N_1846,N_1575);
and U2160 (N_2160,N_1658,N_1573);
or U2161 (N_2161,N_1609,N_1854);
and U2162 (N_2162,N_1524,N_1942);
or U2163 (N_2163,N_1832,N_1568);
nor U2164 (N_2164,N_1946,N_1505);
xor U2165 (N_2165,N_1992,N_1729);
nand U2166 (N_2166,N_1517,N_1613);
or U2167 (N_2167,N_1594,N_1904);
nand U2168 (N_2168,N_1975,N_1824);
or U2169 (N_2169,N_1874,N_1732);
nor U2170 (N_2170,N_1727,N_1550);
nor U2171 (N_2171,N_1951,N_1928);
or U2172 (N_2172,N_1623,N_1677);
or U2173 (N_2173,N_1752,N_1828);
nor U2174 (N_2174,N_1772,N_1625);
and U2175 (N_2175,N_1971,N_1794);
and U2176 (N_2176,N_1907,N_1970);
nand U2177 (N_2177,N_1711,N_1557);
nor U2178 (N_2178,N_1916,N_1642);
nand U2179 (N_2179,N_1620,N_1562);
or U2180 (N_2180,N_1855,N_1811);
or U2181 (N_2181,N_1567,N_1887);
xor U2182 (N_2182,N_1540,N_1986);
or U2183 (N_2183,N_1537,N_1947);
nor U2184 (N_2184,N_1716,N_1818);
and U2185 (N_2185,N_1704,N_1976);
xor U2186 (N_2186,N_1518,N_1626);
and U2187 (N_2187,N_1759,N_1512);
or U2188 (N_2188,N_1806,N_1631);
nor U2189 (N_2189,N_1858,N_1781);
nand U2190 (N_2190,N_1997,N_1888);
and U2191 (N_2191,N_1577,N_1834);
nand U2192 (N_2192,N_1958,N_1605);
or U2193 (N_2193,N_1595,N_1973);
or U2194 (N_2194,N_1925,N_1810);
or U2195 (N_2195,N_1696,N_1587);
nor U2196 (N_2196,N_1508,N_1805);
xor U2197 (N_2197,N_1815,N_1666);
or U2198 (N_2198,N_1681,N_1753);
nand U2199 (N_2199,N_1549,N_1896);
nor U2200 (N_2200,N_1501,N_1895);
or U2201 (N_2201,N_1783,N_1751);
or U2202 (N_2202,N_1817,N_1721);
and U2203 (N_2203,N_1591,N_1929);
xnor U2204 (N_2204,N_1833,N_1900);
nor U2205 (N_2205,N_1886,N_1722);
nand U2206 (N_2206,N_1536,N_1965);
xor U2207 (N_2207,N_1683,N_1709);
xor U2208 (N_2208,N_1875,N_1906);
nor U2209 (N_2209,N_1608,N_1515);
xnor U2210 (N_2210,N_1597,N_1802);
xnor U2211 (N_2211,N_1774,N_1686);
xor U2212 (N_2212,N_1812,N_1853);
and U2213 (N_2213,N_1581,N_1747);
nor U2214 (N_2214,N_1831,N_1633);
xnor U2215 (N_2215,N_1561,N_1511);
or U2216 (N_2216,N_1706,N_1648);
or U2217 (N_2217,N_1639,N_1551);
nor U2218 (N_2218,N_1600,N_1848);
and U2219 (N_2219,N_1953,N_1884);
nor U2220 (N_2220,N_1758,N_1572);
or U2221 (N_2221,N_1821,N_1684);
nand U2222 (N_2222,N_1590,N_1934);
xnor U2223 (N_2223,N_1689,N_1865);
and U2224 (N_2224,N_1735,N_1837);
or U2225 (N_2225,N_1935,N_1529);
nor U2226 (N_2226,N_1775,N_1969);
nor U2227 (N_2227,N_1699,N_1859);
and U2228 (N_2228,N_1921,N_1911);
nor U2229 (N_2229,N_1532,N_1650);
and U2230 (N_2230,N_1601,N_1636);
xnor U2231 (N_2231,N_1695,N_1995);
nor U2232 (N_2232,N_1715,N_1553);
or U2233 (N_2233,N_1892,N_1685);
and U2234 (N_2234,N_1882,N_1968);
nor U2235 (N_2235,N_1712,N_1924);
or U2236 (N_2236,N_1520,N_1926);
nand U2237 (N_2237,N_1525,N_1785);
xnor U2238 (N_2238,N_1792,N_1816);
nand U2239 (N_2239,N_1963,N_1739);
xor U2240 (N_2240,N_1912,N_1654);
or U2241 (N_2241,N_1663,N_1707);
and U2242 (N_2242,N_1823,N_1784);
or U2243 (N_2243,N_1588,N_1583);
and U2244 (N_2244,N_1908,N_1850);
nand U2245 (N_2245,N_1786,N_1780);
nand U2246 (N_2246,N_1669,N_1579);
nand U2247 (N_2247,N_1808,N_1765);
and U2248 (N_2248,N_1584,N_1891);
nand U2249 (N_2249,N_1653,N_1502);
and U2250 (N_2250,N_1868,N_1592);
nand U2251 (N_2251,N_1691,N_1810);
and U2252 (N_2252,N_1578,N_1895);
nor U2253 (N_2253,N_1722,N_1950);
or U2254 (N_2254,N_1978,N_1620);
nor U2255 (N_2255,N_1629,N_1991);
and U2256 (N_2256,N_1767,N_1652);
and U2257 (N_2257,N_1776,N_1590);
and U2258 (N_2258,N_1909,N_1849);
xor U2259 (N_2259,N_1750,N_1970);
xor U2260 (N_2260,N_1786,N_1845);
and U2261 (N_2261,N_1710,N_1976);
or U2262 (N_2262,N_1613,N_1983);
or U2263 (N_2263,N_1546,N_1704);
or U2264 (N_2264,N_1800,N_1851);
xor U2265 (N_2265,N_1832,N_1589);
nor U2266 (N_2266,N_1970,N_1918);
nand U2267 (N_2267,N_1593,N_1759);
or U2268 (N_2268,N_1946,N_1822);
xor U2269 (N_2269,N_1853,N_1728);
nor U2270 (N_2270,N_1955,N_1748);
nor U2271 (N_2271,N_1532,N_1772);
xnor U2272 (N_2272,N_1871,N_1741);
or U2273 (N_2273,N_1890,N_1689);
nand U2274 (N_2274,N_1792,N_1995);
or U2275 (N_2275,N_1620,N_1861);
nand U2276 (N_2276,N_1797,N_1964);
or U2277 (N_2277,N_1944,N_1671);
xor U2278 (N_2278,N_1693,N_1651);
nor U2279 (N_2279,N_1948,N_1960);
or U2280 (N_2280,N_1720,N_1787);
nor U2281 (N_2281,N_1568,N_1686);
nor U2282 (N_2282,N_1709,N_1530);
or U2283 (N_2283,N_1987,N_1600);
and U2284 (N_2284,N_1900,N_1883);
and U2285 (N_2285,N_1574,N_1992);
and U2286 (N_2286,N_1625,N_1673);
nand U2287 (N_2287,N_1653,N_1793);
nor U2288 (N_2288,N_1633,N_1519);
and U2289 (N_2289,N_1843,N_1902);
nor U2290 (N_2290,N_1807,N_1889);
or U2291 (N_2291,N_1883,N_1791);
or U2292 (N_2292,N_1947,N_1842);
nor U2293 (N_2293,N_1589,N_1501);
nand U2294 (N_2294,N_1771,N_1882);
or U2295 (N_2295,N_1740,N_1636);
nor U2296 (N_2296,N_1887,N_1925);
and U2297 (N_2297,N_1825,N_1701);
or U2298 (N_2298,N_1653,N_1990);
and U2299 (N_2299,N_1913,N_1706);
xnor U2300 (N_2300,N_1855,N_1994);
nand U2301 (N_2301,N_1661,N_1904);
or U2302 (N_2302,N_1764,N_1927);
xor U2303 (N_2303,N_1850,N_1903);
or U2304 (N_2304,N_1954,N_1817);
or U2305 (N_2305,N_1891,N_1573);
and U2306 (N_2306,N_1512,N_1931);
nor U2307 (N_2307,N_1604,N_1507);
xnor U2308 (N_2308,N_1708,N_1848);
nor U2309 (N_2309,N_1581,N_1911);
and U2310 (N_2310,N_1778,N_1537);
nor U2311 (N_2311,N_1837,N_1595);
and U2312 (N_2312,N_1857,N_1677);
or U2313 (N_2313,N_1768,N_1833);
nor U2314 (N_2314,N_1612,N_1902);
nand U2315 (N_2315,N_1855,N_1967);
and U2316 (N_2316,N_1880,N_1842);
and U2317 (N_2317,N_1645,N_1999);
nand U2318 (N_2318,N_1908,N_1942);
and U2319 (N_2319,N_1508,N_1851);
xor U2320 (N_2320,N_1619,N_1786);
nor U2321 (N_2321,N_1934,N_1976);
or U2322 (N_2322,N_1670,N_1699);
nand U2323 (N_2323,N_1705,N_1505);
and U2324 (N_2324,N_1767,N_1738);
nor U2325 (N_2325,N_1725,N_1520);
xnor U2326 (N_2326,N_1522,N_1746);
nand U2327 (N_2327,N_1651,N_1880);
or U2328 (N_2328,N_1609,N_1637);
or U2329 (N_2329,N_1682,N_1596);
and U2330 (N_2330,N_1958,N_1729);
and U2331 (N_2331,N_1572,N_1992);
or U2332 (N_2332,N_1996,N_1816);
nor U2333 (N_2333,N_1678,N_1851);
and U2334 (N_2334,N_1687,N_1850);
or U2335 (N_2335,N_1774,N_1816);
and U2336 (N_2336,N_1824,N_1560);
nor U2337 (N_2337,N_1856,N_1641);
or U2338 (N_2338,N_1522,N_1741);
and U2339 (N_2339,N_1541,N_1844);
or U2340 (N_2340,N_1596,N_1700);
xor U2341 (N_2341,N_1531,N_1501);
nor U2342 (N_2342,N_1594,N_1845);
nand U2343 (N_2343,N_1742,N_1991);
nor U2344 (N_2344,N_1990,N_1946);
xnor U2345 (N_2345,N_1542,N_1916);
xnor U2346 (N_2346,N_1965,N_1862);
xnor U2347 (N_2347,N_1745,N_1738);
and U2348 (N_2348,N_1520,N_1855);
nor U2349 (N_2349,N_1996,N_1911);
xnor U2350 (N_2350,N_1740,N_1661);
xnor U2351 (N_2351,N_1993,N_1948);
xnor U2352 (N_2352,N_1994,N_1918);
xnor U2353 (N_2353,N_1869,N_1674);
nand U2354 (N_2354,N_1513,N_1846);
or U2355 (N_2355,N_1574,N_1682);
and U2356 (N_2356,N_1731,N_1773);
nand U2357 (N_2357,N_1888,N_1871);
and U2358 (N_2358,N_1937,N_1933);
nand U2359 (N_2359,N_1809,N_1515);
xnor U2360 (N_2360,N_1983,N_1819);
and U2361 (N_2361,N_1844,N_1553);
nor U2362 (N_2362,N_1583,N_1731);
nor U2363 (N_2363,N_1955,N_1544);
and U2364 (N_2364,N_1519,N_1565);
and U2365 (N_2365,N_1717,N_1910);
xnor U2366 (N_2366,N_1538,N_1579);
nor U2367 (N_2367,N_1674,N_1905);
nor U2368 (N_2368,N_1686,N_1808);
nand U2369 (N_2369,N_1771,N_1930);
nand U2370 (N_2370,N_1936,N_1637);
nor U2371 (N_2371,N_1727,N_1870);
nand U2372 (N_2372,N_1805,N_1533);
xor U2373 (N_2373,N_1675,N_1918);
and U2374 (N_2374,N_1757,N_1936);
or U2375 (N_2375,N_1939,N_1584);
xnor U2376 (N_2376,N_1525,N_1721);
or U2377 (N_2377,N_1977,N_1818);
or U2378 (N_2378,N_1552,N_1991);
and U2379 (N_2379,N_1601,N_1839);
or U2380 (N_2380,N_1815,N_1935);
and U2381 (N_2381,N_1926,N_1613);
nand U2382 (N_2382,N_1610,N_1654);
xor U2383 (N_2383,N_1555,N_1516);
or U2384 (N_2384,N_1520,N_1723);
nor U2385 (N_2385,N_1604,N_1864);
and U2386 (N_2386,N_1764,N_1933);
xor U2387 (N_2387,N_1774,N_1995);
nand U2388 (N_2388,N_1812,N_1847);
xor U2389 (N_2389,N_1504,N_1617);
and U2390 (N_2390,N_1650,N_1927);
or U2391 (N_2391,N_1527,N_1904);
or U2392 (N_2392,N_1735,N_1860);
or U2393 (N_2393,N_1515,N_1856);
and U2394 (N_2394,N_1724,N_1801);
nand U2395 (N_2395,N_1523,N_1680);
nor U2396 (N_2396,N_1616,N_1684);
nor U2397 (N_2397,N_1757,N_1940);
xor U2398 (N_2398,N_1943,N_1932);
and U2399 (N_2399,N_1822,N_1869);
nor U2400 (N_2400,N_1505,N_1778);
nor U2401 (N_2401,N_1506,N_1651);
nand U2402 (N_2402,N_1985,N_1579);
nor U2403 (N_2403,N_1720,N_1689);
xor U2404 (N_2404,N_1658,N_1607);
nand U2405 (N_2405,N_1528,N_1579);
nor U2406 (N_2406,N_1830,N_1741);
or U2407 (N_2407,N_1867,N_1586);
and U2408 (N_2408,N_1935,N_1686);
xnor U2409 (N_2409,N_1701,N_1990);
and U2410 (N_2410,N_1715,N_1916);
and U2411 (N_2411,N_1775,N_1699);
or U2412 (N_2412,N_1721,N_1957);
and U2413 (N_2413,N_1682,N_1885);
or U2414 (N_2414,N_1994,N_1614);
xnor U2415 (N_2415,N_1876,N_1655);
nand U2416 (N_2416,N_1569,N_1525);
and U2417 (N_2417,N_1836,N_1772);
or U2418 (N_2418,N_1717,N_1942);
nand U2419 (N_2419,N_1681,N_1651);
xnor U2420 (N_2420,N_1743,N_1950);
xnor U2421 (N_2421,N_1924,N_1874);
nand U2422 (N_2422,N_1803,N_1583);
and U2423 (N_2423,N_1937,N_1775);
or U2424 (N_2424,N_1771,N_1717);
nor U2425 (N_2425,N_1640,N_1730);
or U2426 (N_2426,N_1951,N_1533);
nor U2427 (N_2427,N_1630,N_1580);
or U2428 (N_2428,N_1944,N_1959);
and U2429 (N_2429,N_1634,N_1728);
nand U2430 (N_2430,N_1784,N_1752);
xor U2431 (N_2431,N_1898,N_1754);
nor U2432 (N_2432,N_1920,N_1509);
and U2433 (N_2433,N_1612,N_1604);
nand U2434 (N_2434,N_1678,N_1977);
and U2435 (N_2435,N_1681,N_1767);
or U2436 (N_2436,N_1621,N_1749);
xnor U2437 (N_2437,N_1860,N_1810);
nand U2438 (N_2438,N_1712,N_1952);
and U2439 (N_2439,N_1805,N_1968);
nor U2440 (N_2440,N_1747,N_1621);
xor U2441 (N_2441,N_1672,N_1647);
nor U2442 (N_2442,N_1541,N_1938);
nand U2443 (N_2443,N_1620,N_1891);
and U2444 (N_2444,N_1687,N_1551);
and U2445 (N_2445,N_1682,N_1579);
xor U2446 (N_2446,N_1830,N_1869);
and U2447 (N_2447,N_1965,N_1764);
xor U2448 (N_2448,N_1907,N_1764);
nor U2449 (N_2449,N_1736,N_1552);
nand U2450 (N_2450,N_1809,N_1725);
nand U2451 (N_2451,N_1686,N_1585);
or U2452 (N_2452,N_1798,N_1570);
xor U2453 (N_2453,N_1573,N_1819);
and U2454 (N_2454,N_1516,N_1614);
and U2455 (N_2455,N_1679,N_1725);
nor U2456 (N_2456,N_1951,N_1585);
nor U2457 (N_2457,N_1529,N_1826);
or U2458 (N_2458,N_1948,N_1611);
xor U2459 (N_2459,N_1965,N_1938);
xnor U2460 (N_2460,N_1581,N_1861);
and U2461 (N_2461,N_1525,N_1631);
xor U2462 (N_2462,N_1653,N_1565);
nand U2463 (N_2463,N_1672,N_1620);
nand U2464 (N_2464,N_1717,N_1599);
nor U2465 (N_2465,N_1620,N_1581);
xnor U2466 (N_2466,N_1677,N_1926);
and U2467 (N_2467,N_1994,N_1688);
nor U2468 (N_2468,N_1920,N_1679);
or U2469 (N_2469,N_1787,N_1618);
or U2470 (N_2470,N_1749,N_1724);
nand U2471 (N_2471,N_1955,N_1521);
nor U2472 (N_2472,N_1828,N_1871);
or U2473 (N_2473,N_1765,N_1876);
nor U2474 (N_2474,N_1839,N_1837);
and U2475 (N_2475,N_1676,N_1542);
xor U2476 (N_2476,N_1888,N_1954);
nand U2477 (N_2477,N_1546,N_1839);
and U2478 (N_2478,N_1892,N_1675);
nor U2479 (N_2479,N_1996,N_1568);
nor U2480 (N_2480,N_1644,N_1641);
and U2481 (N_2481,N_1923,N_1587);
nor U2482 (N_2482,N_1767,N_1628);
nand U2483 (N_2483,N_1799,N_1591);
and U2484 (N_2484,N_1882,N_1884);
nand U2485 (N_2485,N_1875,N_1506);
or U2486 (N_2486,N_1913,N_1917);
or U2487 (N_2487,N_1807,N_1848);
xor U2488 (N_2488,N_1944,N_1514);
or U2489 (N_2489,N_1700,N_1549);
and U2490 (N_2490,N_1540,N_1894);
nor U2491 (N_2491,N_1816,N_1672);
or U2492 (N_2492,N_1685,N_1843);
xnor U2493 (N_2493,N_1584,N_1782);
or U2494 (N_2494,N_1695,N_1594);
nor U2495 (N_2495,N_1655,N_1591);
nor U2496 (N_2496,N_1771,N_1517);
nor U2497 (N_2497,N_1833,N_1550);
or U2498 (N_2498,N_1848,N_1655);
and U2499 (N_2499,N_1666,N_1986);
and U2500 (N_2500,N_2438,N_2179);
or U2501 (N_2501,N_2274,N_2080);
xor U2502 (N_2502,N_2313,N_2340);
nor U2503 (N_2503,N_2498,N_2225);
or U2504 (N_2504,N_2169,N_2445);
or U2505 (N_2505,N_2453,N_2481);
or U2506 (N_2506,N_2330,N_2218);
nand U2507 (N_2507,N_2053,N_2353);
xnor U2508 (N_2508,N_2231,N_2054);
xnor U2509 (N_2509,N_2293,N_2138);
nand U2510 (N_2510,N_2212,N_2206);
nor U2511 (N_2511,N_2027,N_2450);
nand U2512 (N_2512,N_2367,N_2476);
xor U2513 (N_2513,N_2013,N_2331);
nand U2514 (N_2514,N_2074,N_2364);
and U2515 (N_2515,N_2458,N_2076);
nor U2516 (N_2516,N_2121,N_2365);
nand U2517 (N_2517,N_2421,N_2393);
or U2518 (N_2518,N_2485,N_2449);
nor U2519 (N_2519,N_2166,N_2363);
or U2520 (N_2520,N_2203,N_2031);
nand U2521 (N_2521,N_2041,N_2300);
and U2522 (N_2522,N_2046,N_2264);
or U2523 (N_2523,N_2047,N_2327);
and U2524 (N_2524,N_2333,N_2127);
or U2525 (N_2525,N_2226,N_2238);
xnor U2526 (N_2526,N_2192,N_2084);
nor U2527 (N_2527,N_2336,N_2362);
nand U2528 (N_2528,N_2042,N_2297);
nand U2529 (N_2529,N_2168,N_2234);
and U2530 (N_2530,N_2470,N_2173);
nor U2531 (N_2531,N_2093,N_2137);
nand U2532 (N_2532,N_2286,N_2396);
xnor U2533 (N_2533,N_2260,N_2318);
xor U2534 (N_2534,N_2180,N_2237);
or U2535 (N_2535,N_2194,N_2295);
and U2536 (N_2536,N_2221,N_2468);
xor U2537 (N_2537,N_2267,N_2193);
and U2538 (N_2538,N_2029,N_2156);
nand U2539 (N_2539,N_2018,N_2134);
nor U2540 (N_2540,N_2411,N_2355);
xor U2541 (N_2541,N_2435,N_2131);
and U2542 (N_2542,N_2145,N_2250);
nand U2543 (N_2543,N_2429,N_2271);
nor U2544 (N_2544,N_2241,N_2368);
or U2545 (N_2545,N_2125,N_2290);
nand U2546 (N_2546,N_2273,N_2069);
or U2547 (N_2547,N_2142,N_2382);
xnor U2548 (N_2548,N_2437,N_2208);
nand U2549 (N_2549,N_2409,N_2099);
xnor U2550 (N_2550,N_2161,N_2051);
nand U2551 (N_2551,N_2164,N_2083);
xnor U2552 (N_2552,N_2000,N_2104);
and U2553 (N_2553,N_2279,N_2063);
xnor U2554 (N_2554,N_2191,N_2328);
and U2555 (N_2555,N_2348,N_2244);
or U2556 (N_2556,N_2439,N_2281);
xnor U2557 (N_2557,N_2150,N_2268);
xnor U2558 (N_2558,N_2426,N_2052);
and U2559 (N_2559,N_2431,N_2320);
nand U2560 (N_2560,N_2228,N_2397);
xnor U2561 (N_2561,N_2023,N_2332);
nand U2562 (N_2562,N_2072,N_2002);
nor U2563 (N_2563,N_2033,N_2132);
and U2564 (N_2564,N_2466,N_2464);
nor U2565 (N_2565,N_2372,N_2144);
nand U2566 (N_2566,N_2460,N_2189);
nor U2567 (N_2567,N_2098,N_2478);
nor U2568 (N_2568,N_2366,N_2386);
nand U2569 (N_2569,N_2112,N_2287);
and U2570 (N_2570,N_2103,N_2135);
or U2571 (N_2571,N_2389,N_2307);
xnor U2572 (N_2572,N_2178,N_2055);
or U2573 (N_2573,N_2010,N_2339);
nand U2574 (N_2574,N_2251,N_2037);
nand U2575 (N_2575,N_2216,N_2105);
nand U2576 (N_2576,N_2116,N_2067);
and U2577 (N_2577,N_2182,N_2423);
nand U2578 (N_2578,N_2249,N_2489);
nand U2579 (N_2579,N_2130,N_2111);
or U2580 (N_2580,N_2427,N_2197);
xor U2581 (N_2581,N_2494,N_2424);
xnor U2582 (N_2582,N_2443,N_2341);
xor U2583 (N_2583,N_2337,N_2107);
xor U2584 (N_2584,N_2088,N_2275);
xnor U2585 (N_2585,N_2109,N_2085);
or U2586 (N_2586,N_2413,N_2309);
nor U2587 (N_2587,N_2495,N_2172);
xor U2588 (N_2588,N_2209,N_2266);
nor U2589 (N_2589,N_2202,N_2376);
xor U2590 (N_2590,N_2324,N_2378);
xor U2591 (N_2591,N_2402,N_2416);
or U2592 (N_2592,N_2181,N_2422);
nand U2593 (N_2593,N_2484,N_2482);
nand U2594 (N_2594,N_2113,N_2152);
nor U2595 (N_2595,N_2428,N_2448);
nor U2596 (N_2596,N_2154,N_2357);
and U2597 (N_2597,N_2222,N_2346);
and U2598 (N_2598,N_2456,N_2235);
and U2599 (N_2599,N_2361,N_2289);
nor U2600 (N_2600,N_2252,N_2493);
xor U2601 (N_2601,N_2070,N_2284);
and U2602 (N_2602,N_2303,N_2040);
xnor U2603 (N_2603,N_2319,N_2463);
or U2604 (N_2604,N_2308,N_2149);
nand U2605 (N_2605,N_2081,N_2391);
xnor U2606 (N_2606,N_2079,N_2377);
xor U2607 (N_2607,N_2165,N_2020);
or U2608 (N_2608,N_2255,N_2043);
nor U2609 (N_2609,N_2167,N_2269);
nor U2610 (N_2610,N_2342,N_2101);
xnor U2611 (N_2611,N_2242,N_2406);
and U2612 (N_2612,N_2469,N_2133);
xnor U2613 (N_2613,N_2057,N_2270);
or U2614 (N_2614,N_2451,N_2229);
and U2615 (N_2615,N_2188,N_2110);
or U2616 (N_2616,N_2457,N_2487);
nor U2617 (N_2617,N_2227,N_2418);
nor U2618 (N_2618,N_2455,N_2177);
xor U2619 (N_2619,N_2369,N_2210);
nor U2620 (N_2620,N_2347,N_2399);
and U2621 (N_2621,N_2078,N_2232);
nand U2622 (N_2622,N_2442,N_2441);
nand U2623 (N_2623,N_2265,N_2415);
nor U2624 (N_2624,N_2326,N_2459);
nand U2625 (N_2625,N_2499,N_2082);
and U2626 (N_2626,N_2205,N_2021);
or U2627 (N_2627,N_2049,N_2374);
and U2628 (N_2628,N_2417,N_2220);
nand U2629 (N_2629,N_2474,N_2473);
and U2630 (N_2630,N_2350,N_2479);
xor U2631 (N_2631,N_2388,N_2175);
nor U2632 (N_2632,N_2224,N_2146);
xor U2633 (N_2633,N_2400,N_2183);
nor U2634 (N_2634,N_2038,N_2120);
and U2635 (N_2635,N_2017,N_2001);
nand U2636 (N_2636,N_2073,N_2184);
nand U2637 (N_2637,N_2315,N_2176);
or U2638 (N_2638,N_2299,N_2323);
nand U2639 (N_2639,N_2490,N_2405);
and U2640 (N_2640,N_2440,N_2118);
nor U2641 (N_2641,N_2282,N_2061);
and U2642 (N_2642,N_2025,N_2086);
nand U2643 (N_2643,N_2095,N_2026);
and U2644 (N_2644,N_2354,N_2370);
nand U2645 (N_2645,N_2048,N_2199);
xnor U2646 (N_2646,N_2217,N_2153);
nor U2647 (N_2647,N_2301,N_2465);
or U2648 (N_2648,N_2233,N_2062);
or U2649 (N_2649,N_2163,N_2005);
xnor U2650 (N_2650,N_2497,N_2288);
and U2651 (N_2651,N_2028,N_2124);
xnor U2652 (N_2652,N_2343,N_2472);
and U2653 (N_2653,N_2380,N_2012);
nand U2654 (N_2654,N_2059,N_2444);
and U2655 (N_2655,N_2408,N_2296);
or U2656 (N_2656,N_2034,N_2117);
xor U2657 (N_2657,N_2486,N_2345);
nand U2658 (N_2658,N_2185,N_2258);
and U2659 (N_2659,N_2195,N_2174);
nand U2660 (N_2660,N_2066,N_2196);
or U2661 (N_2661,N_2432,N_2285);
or U2662 (N_2662,N_2219,N_2262);
nand U2663 (N_2663,N_2211,N_2283);
xor U2664 (N_2664,N_2036,N_2230);
nand U2665 (N_2665,N_2122,N_2159);
xor U2666 (N_2666,N_2114,N_2214);
nor U2667 (N_2667,N_2058,N_2129);
and U2668 (N_2668,N_2412,N_2089);
and U2669 (N_2669,N_2065,N_2071);
nor U2670 (N_2670,N_2140,N_2280);
nand U2671 (N_2671,N_2024,N_2186);
xnor U2672 (N_2672,N_2371,N_2030);
nand U2673 (N_2673,N_2151,N_2312);
nand U2674 (N_2674,N_2119,N_2011);
nor U2675 (N_2675,N_2141,N_2096);
nor U2676 (N_2676,N_2200,N_2395);
xnor U2677 (N_2677,N_2492,N_2410);
and U2678 (N_2678,N_2007,N_2277);
nor U2679 (N_2679,N_2246,N_2108);
nand U2680 (N_2680,N_2272,N_2204);
nor U2681 (N_2681,N_2436,N_2008);
xnor U2682 (N_2682,N_2398,N_2434);
and U2683 (N_2683,N_2068,N_2321);
xnor U2684 (N_2684,N_2022,N_2128);
nand U2685 (N_2685,N_2394,N_2092);
or U2686 (N_2686,N_2253,N_2006);
or U2687 (N_2687,N_2039,N_2298);
or U2688 (N_2688,N_2254,N_2257);
nor U2689 (N_2689,N_2004,N_2373);
or U2690 (N_2690,N_2091,N_2335);
or U2691 (N_2691,N_2447,N_2452);
or U2692 (N_2692,N_2155,N_2379);
nand U2693 (N_2693,N_2123,N_2462);
nand U2694 (N_2694,N_2467,N_2240);
nor U2695 (N_2695,N_2015,N_2243);
or U2696 (N_2696,N_2259,N_2381);
nand U2697 (N_2697,N_2087,N_2050);
or U2698 (N_2698,N_2414,N_2390);
xnor U2699 (N_2699,N_2094,N_2317);
nand U2700 (N_2700,N_2461,N_2488);
nor U2701 (N_2701,N_2223,N_2344);
nor U2702 (N_2702,N_2170,N_2097);
nand U2703 (N_2703,N_2475,N_2329);
nand U2704 (N_2704,N_2215,N_2322);
or U2705 (N_2705,N_2014,N_2158);
xnor U2706 (N_2706,N_2075,N_2419);
and U2707 (N_2707,N_2292,N_2360);
nand U2708 (N_2708,N_2201,N_2213);
nor U2709 (N_2709,N_2106,N_2157);
xor U2710 (N_2710,N_2198,N_2276);
nand U2711 (N_2711,N_2045,N_2126);
and U2712 (N_2712,N_2143,N_2349);
nand U2713 (N_2713,N_2256,N_2003);
and U2714 (N_2714,N_2060,N_2236);
nand U2715 (N_2715,N_2044,N_2187);
or U2716 (N_2716,N_2139,N_2160);
nor U2717 (N_2717,N_2171,N_2316);
nand U2718 (N_2718,N_2245,N_2190);
nand U2719 (N_2719,N_2404,N_2035);
and U2720 (N_2720,N_2162,N_2403);
nand U2721 (N_2721,N_2306,N_2311);
xor U2722 (N_2722,N_2090,N_2483);
xor U2723 (N_2723,N_2356,N_2147);
nand U2724 (N_2724,N_2294,N_2016);
and U2725 (N_2725,N_2401,N_2302);
xor U2726 (N_2726,N_2064,N_2056);
or U2727 (N_2727,N_2359,N_2310);
nand U2728 (N_2728,N_2358,N_2136);
nor U2729 (N_2729,N_2009,N_2305);
xor U2730 (N_2730,N_2491,N_2351);
nand U2731 (N_2731,N_2115,N_2407);
nor U2732 (N_2732,N_2352,N_2496);
nand U2733 (N_2733,N_2334,N_2263);
xnor U2734 (N_2734,N_2454,N_2019);
xnor U2735 (N_2735,N_2430,N_2239);
or U2736 (N_2736,N_2480,N_2387);
and U2737 (N_2737,N_2477,N_2207);
or U2738 (N_2738,N_2278,N_2314);
or U2739 (N_2739,N_2304,N_2385);
nor U2740 (N_2740,N_2338,N_2392);
or U2741 (N_2741,N_2100,N_2384);
xnor U2742 (N_2742,N_2446,N_2248);
or U2743 (N_2743,N_2325,N_2375);
and U2744 (N_2744,N_2471,N_2077);
nor U2745 (N_2745,N_2261,N_2383);
nor U2746 (N_2746,N_2247,N_2102);
xor U2747 (N_2747,N_2148,N_2433);
nor U2748 (N_2748,N_2291,N_2032);
and U2749 (N_2749,N_2420,N_2425);
or U2750 (N_2750,N_2216,N_2253);
nand U2751 (N_2751,N_2176,N_2368);
nand U2752 (N_2752,N_2023,N_2213);
xnor U2753 (N_2753,N_2176,N_2287);
or U2754 (N_2754,N_2194,N_2234);
and U2755 (N_2755,N_2179,N_2154);
xor U2756 (N_2756,N_2474,N_2383);
xnor U2757 (N_2757,N_2320,N_2258);
and U2758 (N_2758,N_2499,N_2217);
or U2759 (N_2759,N_2012,N_2151);
xnor U2760 (N_2760,N_2348,N_2480);
xor U2761 (N_2761,N_2059,N_2138);
nor U2762 (N_2762,N_2136,N_2427);
nand U2763 (N_2763,N_2072,N_2193);
xor U2764 (N_2764,N_2209,N_2138);
xnor U2765 (N_2765,N_2318,N_2188);
and U2766 (N_2766,N_2054,N_2037);
nand U2767 (N_2767,N_2287,N_2499);
and U2768 (N_2768,N_2155,N_2497);
nor U2769 (N_2769,N_2102,N_2352);
or U2770 (N_2770,N_2447,N_2275);
and U2771 (N_2771,N_2119,N_2316);
nor U2772 (N_2772,N_2361,N_2172);
nor U2773 (N_2773,N_2410,N_2138);
nor U2774 (N_2774,N_2192,N_2010);
nand U2775 (N_2775,N_2044,N_2487);
xor U2776 (N_2776,N_2133,N_2244);
xor U2777 (N_2777,N_2325,N_2063);
nor U2778 (N_2778,N_2069,N_2167);
or U2779 (N_2779,N_2299,N_2129);
or U2780 (N_2780,N_2113,N_2381);
nand U2781 (N_2781,N_2027,N_2439);
nor U2782 (N_2782,N_2227,N_2106);
and U2783 (N_2783,N_2480,N_2136);
nor U2784 (N_2784,N_2322,N_2054);
and U2785 (N_2785,N_2215,N_2420);
nand U2786 (N_2786,N_2419,N_2484);
nor U2787 (N_2787,N_2391,N_2327);
or U2788 (N_2788,N_2135,N_2207);
and U2789 (N_2789,N_2303,N_2338);
xor U2790 (N_2790,N_2287,N_2101);
nand U2791 (N_2791,N_2427,N_2447);
nor U2792 (N_2792,N_2448,N_2115);
nor U2793 (N_2793,N_2265,N_2086);
nor U2794 (N_2794,N_2350,N_2196);
xnor U2795 (N_2795,N_2185,N_2181);
xnor U2796 (N_2796,N_2444,N_2115);
and U2797 (N_2797,N_2227,N_2301);
or U2798 (N_2798,N_2425,N_2331);
xnor U2799 (N_2799,N_2116,N_2315);
and U2800 (N_2800,N_2436,N_2385);
nor U2801 (N_2801,N_2308,N_2051);
and U2802 (N_2802,N_2456,N_2358);
or U2803 (N_2803,N_2171,N_2488);
or U2804 (N_2804,N_2481,N_2035);
nor U2805 (N_2805,N_2074,N_2266);
or U2806 (N_2806,N_2207,N_2415);
and U2807 (N_2807,N_2319,N_2417);
nor U2808 (N_2808,N_2330,N_2235);
xor U2809 (N_2809,N_2261,N_2081);
xnor U2810 (N_2810,N_2014,N_2349);
nor U2811 (N_2811,N_2186,N_2350);
or U2812 (N_2812,N_2385,N_2457);
nand U2813 (N_2813,N_2344,N_2295);
nand U2814 (N_2814,N_2312,N_2419);
nor U2815 (N_2815,N_2478,N_2170);
or U2816 (N_2816,N_2290,N_2133);
nor U2817 (N_2817,N_2130,N_2129);
nand U2818 (N_2818,N_2176,N_2027);
xnor U2819 (N_2819,N_2146,N_2395);
or U2820 (N_2820,N_2425,N_2225);
nor U2821 (N_2821,N_2370,N_2272);
or U2822 (N_2822,N_2335,N_2163);
nand U2823 (N_2823,N_2150,N_2264);
or U2824 (N_2824,N_2382,N_2443);
nor U2825 (N_2825,N_2338,N_2058);
nand U2826 (N_2826,N_2045,N_2469);
or U2827 (N_2827,N_2111,N_2030);
nor U2828 (N_2828,N_2105,N_2360);
and U2829 (N_2829,N_2144,N_2056);
nand U2830 (N_2830,N_2362,N_2381);
and U2831 (N_2831,N_2329,N_2066);
xnor U2832 (N_2832,N_2216,N_2113);
nand U2833 (N_2833,N_2159,N_2475);
xor U2834 (N_2834,N_2157,N_2010);
xnor U2835 (N_2835,N_2370,N_2458);
or U2836 (N_2836,N_2314,N_2223);
and U2837 (N_2837,N_2102,N_2375);
nand U2838 (N_2838,N_2295,N_2304);
xnor U2839 (N_2839,N_2346,N_2401);
xor U2840 (N_2840,N_2383,N_2203);
or U2841 (N_2841,N_2059,N_2279);
nand U2842 (N_2842,N_2067,N_2337);
and U2843 (N_2843,N_2410,N_2158);
or U2844 (N_2844,N_2172,N_2005);
and U2845 (N_2845,N_2000,N_2410);
nand U2846 (N_2846,N_2243,N_2442);
xor U2847 (N_2847,N_2319,N_2267);
xor U2848 (N_2848,N_2196,N_2225);
xor U2849 (N_2849,N_2396,N_2126);
and U2850 (N_2850,N_2304,N_2276);
or U2851 (N_2851,N_2499,N_2040);
or U2852 (N_2852,N_2037,N_2382);
nand U2853 (N_2853,N_2288,N_2295);
or U2854 (N_2854,N_2425,N_2437);
and U2855 (N_2855,N_2496,N_2211);
xnor U2856 (N_2856,N_2089,N_2467);
nand U2857 (N_2857,N_2429,N_2382);
nor U2858 (N_2858,N_2410,N_2238);
xor U2859 (N_2859,N_2240,N_2068);
nand U2860 (N_2860,N_2427,N_2472);
nor U2861 (N_2861,N_2260,N_2418);
nand U2862 (N_2862,N_2113,N_2111);
or U2863 (N_2863,N_2137,N_2261);
or U2864 (N_2864,N_2045,N_2014);
or U2865 (N_2865,N_2173,N_2140);
nand U2866 (N_2866,N_2291,N_2025);
nand U2867 (N_2867,N_2382,N_2317);
nand U2868 (N_2868,N_2134,N_2398);
nor U2869 (N_2869,N_2015,N_2421);
or U2870 (N_2870,N_2334,N_2354);
nor U2871 (N_2871,N_2368,N_2089);
xor U2872 (N_2872,N_2119,N_2498);
nand U2873 (N_2873,N_2209,N_2497);
and U2874 (N_2874,N_2059,N_2392);
and U2875 (N_2875,N_2225,N_2288);
nand U2876 (N_2876,N_2259,N_2484);
nand U2877 (N_2877,N_2282,N_2410);
or U2878 (N_2878,N_2050,N_2452);
nand U2879 (N_2879,N_2406,N_2320);
nor U2880 (N_2880,N_2015,N_2492);
xor U2881 (N_2881,N_2474,N_2231);
nor U2882 (N_2882,N_2365,N_2383);
nand U2883 (N_2883,N_2285,N_2417);
and U2884 (N_2884,N_2164,N_2282);
nand U2885 (N_2885,N_2432,N_2147);
nand U2886 (N_2886,N_2304,N_2498);
xor U2887 (N_2887,N_2263,N_2393);
and U2888 (N_2888,N_2359,N_2339);
or U2889 (N_2889,N_2399,N_2422);
xor U2890 (N_2890,N_2182,N_2171);
xnor U2891 (N_2891,N_2487,N_2390);
nand U2892 (N_2892,N_2310,N_2266);
nor U2893 (N_2893,N_2054,N_2274);
xnor U2894 (N_2894,N_2024,N_2419);
nor U2895 (N_2895,N_2202,N_2002);
nand U2896 (N_2896,N_2320,N_2053);
nor U2897 (N_2897,N_2109,N_2435);
xor U2898 (N_2898,N_2125,N_2166);
xor U2899 (N_2899,N_2416,N_2266);
nand U2900 (N_2900,N_2257,N_2132);
nor U2901 (N_2901,N_2060,N_2201);
and U2902 (N_2902,N_2028,N_2340);
nor U2903 (N_2903,N_2116,N_2217);
xnor U2904 (N_2904,N_2380,N_2057);
or U2905 (N_2905,N_2183,N_2211);
xor U2906 (N_2906,N_2193,N_2482);
xnor U2907 (N_2907,N_2344,N_2066);
or U2908 (N_2908,N_2268,N_2104);
xor U2909 (N_2909,N_2257,N_2117);
nor U2910 (N_2910,N_2029,N_2439);
or U2911 (N_2911,N_2301,N_2031);
xor U2912 (N_2912,N_2014,N_2322);
and U2913 (N_2913,N_2156,N_2259);
and U2914 (N_2914,N_2447,N_2174);
and U2915 (N_2915,N_2263,N_2306);
nand U2916 (N_2916,N_2384,N_2108);
nor U2917 (N_2917,N_2352,N_2067);
xor U2918 (N_2918,N_2090,N_2206);
and U2919 (N_2919,N_2310,N_2027);
and U2920 (N_2920,N_2122,N_2246);
nor U2921 (N_2921,N_2209,N_2219);
nor U2922 (N_2922,N_2060,N_2376);
nor U2923 (N_2923,N_2002,N_2351);
or U2924 (N_2924,N_2485,N_2355);
and U2925 (N_2925,N_2269,N_2462);
nand U2926 (N_2926,N_2074,N_2085);
or U2927 (N_2927,N_2457,N_2144);
or U2928 (N_2928,N_2244,N_2115);
nand U2929 (N_2929,N_2147,N_2338);
and U2930 (N_2930,N_2185,N_2208);
xor U2931 (N_2931,N_2137,N_2005);
nand U2932 (N_2932,N_2387,N_2155);
xor U2933 (N_2933,N_2026,N_2460);
nand U2934 (N_2934,N_2484,N_2100);
nor U2935 (N_2935,N_2258,N_2141);
and U2936 (N_2936,N_2261,N_2027);
or U2937 (N_2937,N_2123,N_2481);
xnor U2938 (N_2938,N_2054,N_2327);
xor U2939 (N_2939,N_2194,N_2167);
nor U2940 (N_2940,N_2019,N_2149);
or U2941 (N_2941,N_2486,N_2379);
xor U2942 (N_2942,N_2255,N_2195);
and U2943 (N_2943,N_2089,N_2243);
xnor U2944 (N_2944,N_2366,N_2284);
xor U2945 (N_2945,N_2050,N_2286);
nand U2946 (N_2946,N_2330,N_2318);
nor U2947 (N_2947,N_2087,N_2252);
and U2948 (N_2948,N_2438,N_2121);
or U2949 (N_2949,N_2074,N_2269);
and U2950 (N_2950,N_2119,N_2051);
xnor U2951 (N_2951,N_2368,N_2346);
nand U2952 (N_2952,N_2430,N_2199);
nor U2953 (N_2953,N_2196,N_2367);
and U2954 (N_2954,N_2044,N_2062);
xnor U2955 (N_2955,N_2060,N_2291);
or U2956 (N_2956,N_2162,N_2236);
and U2957 (N_2957,N_2078,N_2445);
nand U2958 (N_2958,N_2038,N_2176);
nor U2959 (N_2959,N_2451,N_2178);
xor U2960 (N_2960,N_2433,N_2169);
nor U2961 (N_2961,N_2340,N_2072);
nor U2962 (N_2962,N_2371,N_2109);
xor U2963 (N_2963,N_2165,N_2269);
xnor U2964 (N_2964,N_2087,N_2331);
nor U2965 (N_2965,N_2246,N_2197);
or U2966 (N_2966,N_2415,N_2262);
xor U2967 (N_2967,N_2484,N_2363);
and U2968 (N_2968,N_2455,N_2117);
xor U2969 (N_2969,N_2361,N_2311);
and U2970 (N_2970,N_2242,N_2008);
xnor U2971 (N_2971,N_2045,N_2308);
and U2972 (N_2972,N_2061,N_2308);
xor U2973 (N_2973,N_2342,N_2178);
and U2974 (N_2974,N_2466,N_2076);
and U2975 (N_2975,N_2120,N_2365);
nand U2976 (N_2976,N_2071,N_2097);
xor U2977 (N_2977,N_2112,N_2119);
nor U2978 (N_2978,N_2476,N_2308);
xnor U2979 (N_2979,N_2372,N_2443);
nor U2980 (N_2980,N_2123,N_2365);
nor U2981 (N_2981,N_2160,N_2446);
or U2982 (N_2982,N_2244,N_2359);
nand U2983 (N_2983,N_2305,N_2136);
nor U2984 (N_2984,N_2424,N_2464);
or U2985 (N_2985,N_2431,N_2433);
or U2986 (N_2986,N_2066,N_2003);
and U2987 (N_2987,N_2367,N_2483);
and U2988 (N_2988,N_2019,N_2467);
or U2989 (N_2989,N_2382,N_2491);
or U2990 (N_2990,N_2298,N_2258);
xor U2991 (N_2991,N_2346,N_2242);
xnor U2992 (N_2992,N_2368,N_2231);
or U2993 (N_2993,N_2320,N_2497);
or U2994 (N_2994,N_2485,N_2199);
xnor U2995 (N_2995,N_2125,N_2204);
nand U2996 (N_2996,N_2272,N_2183);
nand U2997 (N_2997,N_2383,N_2204);
or U2998 (N_2998,N_2083,N_2416);
or U2999 (N_2999,N_2355,N_2135);
nor UO_0 (O_0,N_2961,N_2713);
nand UO_1 (O_1,N_2987,N_2894);
and UO_2 (O_2,N_2798,N_2827);
nand UO_3 (O_3,N_2862,N_2948);
or UO_4 (O_4,N_2936,N_2910);
nand UO_5 (O_5,N_2912,N_2829);
xor UO_6 (O_6,N_2735,N_2556);
xnor UO_7 (O_7,N_2595,N_2803);
nand UO_8 (O_8,N_2875,N_2665);
nand UO_9 (O_9,N_2833,N_2712);
and UO_10 (O_10,N_2573,N_2797);
nand UO_11 (O_11,N_2820,N_2509);
nand UO_12 (O_12,N_2513,N_2818);
or UO_13 (O_13,N_2680,N_2766);
nor UO_14 (O_14,N_2533,N_2524);
or UO_15 (O_15,N_2577,N_2642);
xor UO_16 (O_16,N_2600,N_2799);
nand UO_17 (O_17,N_2685,N_2704);
nor UO_18 (O_18,N_2622,N_2651);
and UO_19 (O_19,N_2541,N_2944);
and UO_20 (O_20,N_2544,N_2714);
xnor UO_21 (O_21,N_2962,N_2521);
xnor UO_22 (O_22,N_2955,N_2525);
xnor UO_23 (O_23,N_2970,N_2957);
nand UO_24 (O_24,N_2527,N_2647);
xnor UO_25 (O_25,N_2806,N_2539);
nand UO_26 (O_26,N_2674,N_2934);
nor UO_27 (O_27,N_2834,N_2514);
nor UO_28 (O_28,N_2515,N_2971);
nand UO_29 (O_29,N_2660,N_2876);
and UO_30 (O_30,N_2675,N_2777);
or UO_31 (O_31,N_2742,N_2903);
and UO_32 (O_32,N_2588,N_2565);
nor UO_33 (O_33,N_2860,N_2842);
or UO_34 (O_34,N_2796,N_2745);
xnor UO_35 (O_35,N_2931,N_2737);
nor UO_36 (O_36,N_2952,N_2579);
and UO_37 (O_37,N_2789,N_2706);
nand UO_38 (O_38,N_2874,N_2758);
nor UO_39 (O_39,N_2784,N_2867);
nand UO_40 (O_40,N_2709,N_2547);
xnor UO_41 (O_41,N_2967,N_2696);
xor UO_42 (O_42,N_2794,N_2715);
or UO_43 (O_43,N_2840,N_2688);
nand UO_44 (O_44,N_2631,N_2984);
xor UO_45 (O_45,N_2736,N_2972);
and UO_46 (O_46,N_2986,N_2727);
xnor UO_47 (O_47,N_2710,N_2734);
nor UO_48 (O_48,N_2708,N_2590);
nand UO_49 (O_49,N_2873,N_2701);
nor UO_50 (O_50,N_2652,N_2643);
nor UO_51 (O_51,N_2662,N_2639);
nor UO_52 (O_52,N_2943,N_2611);
nor UO_53 (O_53,N_2906,N_2644);
nand UO_54 (O_54,N_2949,N_2606);
nand UO_55 (O_55,N_2612,N_2940);
nor UO_56 (O_56,N_2966,N_2907);
nor UO_57 (O_57,N_2793,N_2786);
and UO_58 (O_58,N_2865,N_2522);
and UO_59 (O_59,N_2693,N_2767);
xor UO_60 (O_60,N_2985,N_2730);
xnor UO_61 (O_61,N_2659,N_2695);
xor UO_62 (O_62,N_2673,N_2536);
nand UO_63 (O_63,N_2650,N_2640);
nand UO_64 (O_64,N_2584,N_2807);
nand UO_65 (O_65,N_2511,N_2995);
xor UO_66 (O_66,N_2633,N_2566);
xnor UO_67 (O_67,N_2591,N_2585);
nor UO_68 (O_68,N_2581,N_2849);
xnor UO_69 (O_69,N_2792,N_2750);
nand UO_70 (O_70,N_2603,N_2838);
and UO_71 (O_71,N_2814,N_2996);
and UO_72 (O_72,N_2619,N_2908);
nor UO_73 (O_73,N_2779,N_2726);
and UO_74 (O_74,N_2604,N_2975);
nand UO_75 (O_75,N_2932,N_2601);
and UO_76 (O_76,N_2679,N_2501);
or UO_77 (O_77,N_2607,N_2773);
or UO_78 (O_78,N_2930,N_2625);
nand UO_79 (O_79,N_2655,N_2756);
nor UO_80 (O_80,N_2580,N_2502);
or UO_81 (O_81,N_2871,N_2848);
and UO_82 (O_82,N_2852,N_2677);
xnor UO_83 (O_83,N_2917,N_2761);
or UO_84 (O_84,N_2725,N_2598);
or UO_85 (O_85,N_2620,N_2641);
nor UO_86 (O_86,N_2999,N_2597);
or UO_87 (O_87,N_2645,N_2783);
xnor UO_88 (O_88,N_2671,N_2589);
nand UO_89 (O_89,N_2769,N_2968);
and UO_90 (O_90,N_2692,N_2764);
nor UO_91 (O_91,N_2535,N_2504);
or UO_92 (O_92,N_2686,N_2902);
and UO_93 (O_93,N_2668,N_2549);
nor UO_94 (O_94,N_2754,N_2516);
and UO_95 (O_95,N_2993,N_2979);
xnor UO_96 (O_96,N_2811,N_2836);
nor UO_97 (O_97,N_2878,N_2855);
xnor UO_98 (O_98,N_2746,N_2921);
xnor UO_99 (O_99,N_2560,N_2672);
nand UO_100 (O_100,N_2628,N_2939);
nor UO_101 (O_101,N_2648,N_2621);
and UO_102 (O_102,N_2594,N_2740);
or UO_103 (O_103,N_2540,N_2815);
or UO_104 (O_104,N_2570,N_2850);
or UO_105 (O_105,N_2744,N_2716);
xnor UO_106 (O_106,N_2583,N_2553);
and UO_107 (O_107,N_2670,N_2884);
or UO_108 (O_108,N_2666,N_2667);
and UO_109 (O_109,N_2663,N_2998);
nand UO_110 (O_110,N_2599,N_2562);
nor UO_111 (O_111,N_2963,N_2636);
nand UO_112 (O_112,N_2518,N_2812);
xnor UO_113 (O_113,N_2572,N_2853);
nor UO_114 (O_114,N_2945,N_2956);
and UO_115 (O_115,N_2881,N_2937);
xor UO_116 (O_116,N_2886,N_2500);
or UO_117 (O_117,N_2697,N_2891);
nor UO_118 (O_118,N_2739,N_2752);
or UO_119 (O_119,N_2809,N_2859);
or UO_120 (O_120,N_2658,N_2960);
xnor UO_121 (O_121,N_2958,N_2879);
or UO_122 (O_122,N_2722,N_2916);
nand UO_123 (O_123,N_2854,N_2578);
or UO_124 (O_124,N_2922,N_2942);
xnor UO_125 (O_125,N_2762,N_2520);
xnor UO_126 (O_126,N_2941,N_2623);
xnor UO_127 (O_127,N_2863,N_2888);
or UO_128 (O_128,N_2523,N_2816);
nand UO_129 (O_129,N_2926,N_2733);
or UO_130 (O_130,N_2691,N_2981);
nor UO_131 (O_131,N_2847,N_2519);
nand UO_132 (O_132,N_2534,N_2757);
and UO_133 (O_133,N_2898,N_2813);
xnor UO_134 (O_134,N_2723,N_2507);
nand UO_135 (O_135,N_2990,N_2669);
and UO_136 (O_136,N_2721,N_2864);
nor UO_137 (O_137,N_2707,N_2749);
nor UO_138 (O_138,N_2569,N_2801);
or UO_139 (O_139,N_2657,N_2732);
nor UO_140 (O_140,N_2915,N_2741);
and UO_141 (O_141,N_2768,N_2743);
nor UO_142 (O_142,N_2637,N_2947);
or UO_143 (O_143,N_2763,N_2543);
nand UO_144 (O_144,N_2989,N_2946);
or UO_145 (O_145,N_2824,N_2738);
nor UO_146 (O_146,N_2983,N_2795);
xor UO_147 (O_147,N_2552,N_2808);
and UO_148 (O_148,N_2653,N_2587);
nand UO_149 (O_149,N_2861,N_2800);
and UO_150 (O_150,N_2823,N_2687);
nand UO_151 (O_151,N_2720,N_2885);
xnor UO_152 (O_152,N_2545,N_2914);
nand UO_153 (O_153,N_2872,N_2775);
nor UO_154 (O_154,N_2615,N_2896);
nor UO_155 (O_155,N_2508,N_2537);
nand UO_156 (O_156,N_2618,N_2959);
nand UO_157 (O_157,N_2719,N_2694);
or UO_158 (O_158,N_2835,N_2822);
and UO_159 (O_159,N_2978,N_2568);
and UO_160 (O_160,N_2555,N_2731);
or UO_161 (O_161,N_2724,N_2909);
and UO_162 (O_162,N_2531,N_2846);
and UO_163 (O_163,N_2574,N_2858);
nand UO_164 (O_164,N_2608,N_2857);
nand UO_165 (O_165,N_2887,N_2748);
nand UO_166 (O_166,N_2832,N_2751);
nand UO_167 (O_167,N_2526,N_2558);
nand UO_168 (O_168,N_2895,N_2557);
nor UO_169 (O_169,N_2774,N_2911);
and UO_170 (O_170,N_2828,N_2528);
nor UO_171 (O_171,N_2866,N_2841);
nor UO_172 (O_172,N_2582,N_2969);
xnor UO_173 (O_173,N_2510,N_2678);
and UO_174 (O_174,N_2602,N_2954);
nand UO_175 (O_175,N_2576,N_2548);
xnor UO_176 (O_176,N_2938,N_2964);
and UO_177 (O_177,N_2626,N_2805);
nand UO_178 (O_178,N_2638,N_2778);
nor UO_179 (O_179,N_2919,N_2933);
nor UO_180 (O_180,N_2851,N_2682);
or UO_181 (O_181,N_2563,N_2654);
nor UO_182 (O_182,N_2571,N_2629);
or UO_183 (O_183,N_2561,N_2771);
and UO_184 (O_184,N_2624,N_2976);
and UO_185 (O_185,N_2689,N_2505);
and UO_186 (O_186,N_2925,N_2924);
xnor UO_187 (O_187,N_2550,N_2920);
nand UO_188 (O_188,N_2593,N_2530);
nand UO_189 (O_189,N_2546,N_2897);
nand UO_190 (O_190,N_2973,N_2927);
and UO_191 (O_191,N_2802,N_2965);
nand UO_192 (O_192,N_2953,N_2883);
or UO_193 (O_193,N_2634,N_2684);
nand UO_194 (O_194,N_2890,N_2656);
xor UO_195 (O_195,N_2772,N_2503);
nor UO_196 (O_196,N_2646,N_2901);
nand UO_197 (O_197,N_2681,N_2649);
nand UO_198 (O_198,N_2951,N_2538);
or UO_199 (O_199,N_2664,N_2564);
nand UO_200 (O_200,N_2991,N_2988);
nor UO_201 (O_201,N_2703,N_2627);
xor UO_202 (O_202,N_2617,N_2843);
and UO_203 (O_203,N_2868,N_2705);
and UO_204 (O_204,N_2870,N_2765);
xor UO_205 (O_205,N_2729,N_2632);
or UO_206 (O_206,N_2782,N_2817);
xnor UO_207 (O_207,N_2974,N_2839);
nand UO_208 (O_208,N_2575,N_2554);
and UO_209 (O_209,N_2529,N_2787);
xor UO_210 (O_210,N_2592,N_2880);
or UO_211 (O_211,N_2770,N_2551);
or UO_212 (O_212,N_2929,N_2517);
nand UO_213 (O_213,N_2747,N_2819);
nand UO_214 (O_214,N_2830,N_2785);
nand UO_215 (O_215,N_2610,N_2781);
or UO_216 (O_216,N_2845,N_2698);
nand UO_217 (O_217,N_2635,N_2702);
xnor UO_218 (O_218,N_2776,N_2804);
and UO_219 (O_219,N_2893,N_2918);
nand UO_220 (O_220,N_2586,N_2596);
or UO_221 (O_221,N_2869,N_2661);
nand UO_222 (O_222,N_2699,N_2791);
nand UO_223 (O_223,N_2837,N_2718);
nand UO_224 (O_224,N_2856,N_2913);
xnor UO_225 (O_225,N_2506,N_2928);
or UO_226 (O_226,N_2882,N_2997);
or UO_227 (O_227,N_2676,N_2605);
and UO_228 (O_228,N_2614,N_2728);
and UO_229 (O_229,N_2900,N_2512);
xor UO_230 (O_230,N_2994,N_2821);
xor UO_231 (O_231,N_2683,N_2790);
nor UO_232 (O_232,N_2613,N_2532);
and UO_233 (O_233,N_2760,N_2899);
nor UO_234 (O_234,N_2717,N_2700);
nand UO_235 (O_235,N_2977,N_2935);
or UO_236 (O_236,N_2616,N_2780);
or UO_237 (O_237,N_2877,N_2992);
or UO_238 (O_238,N_2755,N_2982);
nand UO_239 (O_239,N_2826,N_2844);
xor UO_240 (O_240,N_2904,N_2889);
or UO_241 (O_241,N_2788,N_2753);
nor UO_242 (O_242,N_2892,N_2831);
and UO_243 (O_243,N_2690,N_2810);
nand UO_244 (O_244,N_2980,N_2905);
xnor UO_245 (O_245,N_2825,N_2559);
xnor UO_246 (O_246,N_2609,N_2630);
nand UO_247 (O_247,N_2567,N_2711);
or UO_248 (O_248,N_2759,N_2950);
and UO_249 (O_249,N_2542,N_2923);
nor UO_250 (O_250,N_2899,N_2973);
xor UO_251 (O_251,N_2944,N_2813);
and UO_252 (O_252,N_2699,N_2751);
xor UO_253 (O_253,N_2729,N_2592);
nand UO_254 (O_254,N_2616,N_2848);
xnor UO_255 (O_255,N_2836,N_2995);
xnor UO_256 (O_256,N_2578,N_2522);
xor UO_257 (O_257,N_2919,N_2736);
xnor UO_258 (O_258,N_2848,N_2854);
xor UO_259 (O_259,N_2767,N_2949);
nand UO_260 (O_260,N_2728,N_2594);
and UO_261 (O_261,N_2568,N_2843);
or UO_262 (O_262,N_2636,N_2685);
and UO_263 (O_263,N_2598,N_2897);
xor UO_264 (O_264,N_2618,N_2856);
nand UO_265 (O_265,N_2936,N_2671);
nor UO_266 (O_266,N_2770,N_2975);
or UO_267 (O_267,N_2505,N_2854);
xnor UO_268 (O_268,N_2970,N_2886);
xor UO_269 (O_269,N_2860,N_2947);
xor UO_270 (O_270,N_2655,N_2646);
nor UO_271 (O_271,N_2795,N_2598);
or UO_272 (O_272,N_2963,N_2710);
or UO_273 (O_273,N_2910,N_2673);
nor UO_274 (O_274,N_2786,N_2659);
xnor UO_275 (O_275,N_2635,N_2556);
xor UO_276 (O_276,N_2665,N_2792);
xnor UO_277 (O_277,N_2960,N_2815);
and UO_278 (O_278,N_2533,N_2858);
or UO_279 (O_279,N_2718,N_2742);
xnor UO_280 (O_280,N_2586,N_2610);
nor UO_281 (O_281,N_2985,N_2747);
xor UO_282 (O_282,N_2540,N_2539);
and UO_283 (O_283,N_2751,N_2867);
xnor UO_284 (O_284,N_2936,N_2797);
or UO_285 (O_285,N_2722,N_2831);
xnor UO_286 (O_286,N_2966,N_2792);
xor UO_287 (O_287,N_2599,N_2771);
and UO_288 (O_288,N_2753,N_2717);
nor UO_289 (O_289,N_2531,N_2920);
or UO_290 (O_290,N_2542,N_2543);
and UO_291 (O_291,N_2688,N_2878);
xnor UO_292 (O_292,N_2851,N_2654);
xnor UO_293 (O_293,N_2775,N_2693);
or UO_294 (O_294,N_2855,N_2820);
xor UO_295 (O_295,N_2822,N_2837);
nor UO_296 (O_296,N_2521,N_2640);
xor UO_297 (O_297,N_2894,N_2718);
nor UO_298 (O_298,N_2588,N_2858);
and UO_299 (O_299,N_2957,N_2804);
or UO_300 (O_300,N_2594,N_2533);
and UO_301 (O_301,N_2581,N_2566);
nor UO_302 (O_302,N_2943,N_2819);
nor UO_303 (O_303,N_2806,N_2904);
or UO_304 (O_304,N_2985,N_2847);
xor UO_305 (O_305,N_2834,N_2623);
xor UO_306 (O_306,N_2607,N_2593);
and UO_307 (O_307,N_2952,N_2603);
nand UO_308 (O_308,N_2675,N_2518);
and UO_309 (O_309,N_2785,N_2510);
or UO_310 (O_310,N_2878,N_2922);
nand UO_311 (O_311,N_2533,N_2748);
xnor UO_312 (O_312,N_2695,N_2746);
nor UO_313 (O_313,N_2624,N_2512);
nand UO_314 (O_314,N_2508,N_2788);
nor UO_315 (O_315,N_2549,N_2520);
nor UO_316 (O_316,N_2689,N_2770);
or UO_317 (O_317,N_2540,N_2578);
xor UO_318 (O_318,N_2681,N_2669);
or UO_319 (O_319,N_2758,N_2871);
nand UO_320 (O_320,N_2732,N_2635);
nand UO_321 (O_321,N_2956,N_2962);
nor UO_322 (O_322,N_2551,N_2966);
and UO_323 (O_323,N_2638,N_2533);
nand UO_324 (O_324,N_2594,N_2810);
and UO_325 (O_325,N_2502,N_2669);
xnor UO_326 (O_326,N_2824,N_2723);
nand UO_327 (O_327,N_2679,N_2576);
nand UO_328 (O_328,N_2717,N_2696);
xnor UO_329 (O_329,N_2771,N_2676);
nand UO_330 (O_330,N_2747,N_2505);
xnor UO_331 (O_331,N_2638,N_2979);
nand UO_332 (O_332,N_2593,N_2971);
and UO_333 (O_333,N_2948,N_2591);
nor UO_334 (O_334,N_2618,N_2670);
nor UO_335 (O_335,N_2854,N_2974);
or UO_336 (O_336,N_2932,N_2840);
and UO_337 (O_337,N_2514,N_2775);
xnor UO_338 (O_338,N_2984,N_2987);
nand UO_339 (O_339,N_2901,N_2778);
and UO_340 (O_340,N_2618,N_2699);
or UO_341 (O_341,N_2687,N_2631);
nand UO_342 (O_342,N_2833,N_2763);
xnor UO_343 (O_343,N_2600,N_2843);
nor UO_344 (O_344,N_2721,N_2980);
nand UO_345 (O_345,N_2732,N_2859);
and UO_346 (O_346,N_2817,N_2644);
nand UO_347 (O_347,N_2905,N_2791);
nor UO_348 (O_348,N_2667,N_2555);
and UO_349 (O_349,N_2512,N_2909);
nand UO_350 (O_350,N_2861,N_2815);
or UO_351 (O_351,N_2950,N_2971);
and UO_352 (O_352,N_2808,N_2820);
nand UO_353 (O_353,N_2516,N_2861);
nor UO_354 (O_354,N_2749,N_2906);
nand UO_355 (O_355,N_2638,N_2640);
or UO_356 (O_356,N_2604,N_2962);
nand UO_357 (O_357,N_2696,N_2774);
nand UO_358 (O_358,N_2931,N_2800);
or UO_359 (O_359,N_2554,N_2890);
and UO_360 (O_360,N_2971,N_2934);
xor UO_361 (O_361,N_2606,N_2698);
and UO_362 (O_362,N_2836,N_2707);
xnor UO_363 (O_363,N_2906,N_2973);
nor UO_364 (O_364,N_2747,N_2960);
xor UO_365 (O_365,N_2932,N_2858);
and UO_366 (O_366,N_2523,N_2741);
xor UO_367 (O_367,N_2635,N_2937);
nor UO_368 (O_368,N_2843,N_2696);
or UO_369 (O_369,N_2802,N_2597);
nor UO_370 (O_370,N_2735,N_2533);
and UO_371 (O_371,N_2698,N_2979);
nand UO_372 (O_372,N_2561,N_2649);
and UO_373 (O_373,N_2729,N_2691);
nand UO_374 (O_374,N_2782,N_2906);
nor UO_375 (O_375,N_2792,N_2778);
nand UO_376 (O_376,N_2802,N_2649);
and UO_377 (O_377,N_2964,N_2531);
xor UO_378 (O_378,N_2545,N_2573);
xnor UO_379 (O_379,N_2622,N_2871);
or UO_380 (O_380,N_2563,N_2843);
or UO_381 (O_381,N_2619,N_2503);
and UO_382 (O_382,N_2710,N_2860);
nor UO_383 (O_383,N_2691,N_2872);
nor UO_384 (O_384,N_2590,N_2643);
or UO_385 (O_385,N_2540,N_2689);
xor UO_386 (O_386,N_2787,N_2586);
xnor UO_387 (O_387,N_2781,N_2758);
and UO_388 (O_388,N_2957,N_2574);
nand UO_389 (O_389,N_2612,N_2993);
nor UO_390 (O_390,N_2686,N_2861);
xor UO_391 (O_391,N_2819,N_2916);
xor UO_392 (O_392,N_2914,N_2887);
xnor UO_393 (O_393,N_2732,N_2823);
nor UO_394 (O_394,N_2885,N_2871);
xnor UO_395 (O_395,N_2890,N_2973);
nor UO_396 (O_396,N_2567,N_2610);
nand UO_397 (O_397,N_2910,N_2676);
nor UO_398 (O_398,N_2565,N_2735);
or UO_399 (O_399,N_2931,N_2744);
or UO_400 (O_400,N_2803,N_2701);
or UO_401 (O_401,N_2678,N_2692);
nor UO_402 (O_402,N_2596,N_2858);
xnor UO_403 (O_403,N_2931,N_2556);
nor UO_404 (O_404,N_2850,N_2587);
nor UO_405 (O_405,N_2781,N_2796);
and UO_406 (O_406,N_2993,N_2893);
nand UO_407 (O_407,N_2709,N_2927);
or UO_408 (O_408,N_2879,N_2650);
xnor UO_409 (O_409,N_2818,N_2836);
and UO_410 (O_410,N_2886,N_2940);
nand UO_411 (O_411,N_2645,N_2940);
nor UO_412 (O_412,N_2887,N_2645);
xnor UO_413 (O_413,N_2644,N_2555);
nand UO_414 (O_414,N_2914,N_2961);
nand UO_415 (O_415,N_2976,N_2778);
nor UO_416 (O_416,N_2968,N_2648);
nand UO_417 (O_417,N_2691,N_2532);
nand UO_418 (O_418,N_2731,N_2667);
and UO_419 (O_419,N_2648,N_2874);
nand UO_420 (O_420,N_2533,N_2786);
xor UO_421 (O_421,N_2746,N_2823);
xor UO_422 (O_422,N_2992,N_2678);
xnor UO_423 (O_423,N_2903,N_2585);
and UO_424 (O_424,N_2993,N_2624);
nor UO_425 (O_425,N_2870,N_2924);
and UO_426 (O_426,N_2661,N_2966);
xnor UO_427 (O_427,N_2925,N_2947);
nand UO_428 (O_428,N_2557,N_2990);
and UO_429 (O_429,N_2606,N_2994);
xor UO_430 (O_430,N_2544,N_2799);
nor UO_431 (O_431,N_2654,N_2940);
nand UO_432 (O_432,N_2847,N_2849);
xor UO_433 (O_433,N_2838,N_2873);
xnor UO_434 (O_434,N_2543,N_2628);
nor UO_435 (O_435,N_2532,N_2847);
and UO_436 (O_436,N_2964,N_2755);
or UO_437 (O_437,N_2574,N_2945);
nor UO_438 (O_438,N_2760,N_2845);
nor UO_439 (O_439,N_2535,N_2999);
and UO_440 (O_440,N_2863,N_2577);
nand UO_441 (O_441,N_2889,N_2509);
nand UO_442 (O_442,N_2791,N_2589);
xor UO_443 (O_443,N_2832,N_2918);
xor UO_444 (O_444,N_2986,N_2631);
nor UO_445 (O_445,N_2757,N_2818);
or UO_446 (O_446,N_2758,N_2976);
nand UO_447 (O_447,N_2962,N_2967);
nor UO_448 (O_448,N_2727,N_2800);
xor UO_449 (O_449,N_2779,N_2506);
and UO_450 (O_450,N_2991,N_2918);
nand UO_451 (O_451,N_2549,N_2856);
or UO_452 (O_452,N_2907,N_2609);
nand UO_453 (O_453,N_2625,N_2676);
nand UO_454 (O_454,N_2828,N_2904);
nand UO_455 (O_455,N_2806,N_2520);
xnor UO_456 (O_456,N_2532,N_2869);
xor UO_457 (O_457,N_2835,N_2880);
nand UO_458 (O_458,N_2574,N_2784);
nand UO_459 (O_459,N_2598,N_2974);
and UO_460 (O_460,N_2705,N_2690);
nand UO_461 (O_461,N_2814,N_2793);
nor UO_462 (O_462,N_2802,N_2560);
xor UO_463 (O_463,N_2886,N_2651);
and UO_464 (O_464,N_2620,N_2564);
nor UO_465 (O_465,N_2785,N_2886);
or UO_466 (O_466,N_2895,N_2658);
nor UO_467 (O_467,N_2517,N_2611);
xor UO_468 (O_468,N_2856,N_2665);
nor UO_469 (O_469,N_2976,N_2923);
nor UO_470 (O_470,N_2899,N_2514);
and UO_471 (O_471,N_2511,N_2927);
nor UO_472 (O_472,N_2982,N_2640);
and UO_473 (O_473,N_2891,N_2692);
xnor UO_474 (O_474,N_2823,N_2804);
or UO_475 (O_475,N_2710,N_2945);
nand UO_476 (O_476,N_2850,N_2813);
nor UO_477 (O_477,N_2812,N_2591);
and UO_478 (O_478,N_2996,N_2566);
nand UO_479 (O_479,N_2572,N_2624);
or UO_480 (O_480,N_2519,N_2918);
and UO_481 (O_481,N_2709,N_2572);
or UO_482 (O_482,N_2507,N_2781);
xnor UO_483 (O_483,N_2889,N_2731);
and UO_484 (O_484,N_2507,N_2702);
xnor UO_485 (O_485,N_2571,N_2838);
or UO_486 (O_486,N_2998,N_2512);
nand UO_487 (O_487,N_2710,N_2500);
or UO_488 (O_488,N_2854,N_2630);
nor UO_489 (O_489,N_2711,N_2771);
nor UO_490 (O_490,N_2804,N_2974);
nor UO_491 (O_491,N_2903,N_2624);
nor UO_492 (O_492,N_2528,N_2753);
xor UO_493 (O_493,N_2540,N_2515);
xnor UO_494 (O_494,N_2639,N_2581);
and UO_495 (O_495,N_2934,N_2654);
or UO_496 (O_496,N_2877,N_2902);
xnor UO_497 (O_497,N_2583,N_2813);
or UO_498 (O_498,N_2711,N_2899);
nor UO_499 (O_499,N_2770,N_2724);
endmodule