module basic_1500_15000_2000_20_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_333,In_1356);
nand U1 (N_1,In_1041,In_930);
and U2 (N_2,In_464,In_803);
or U3 (N_3,In_1384,In_828);
and U4 (N_4,In_1125,In_694);
nand U5 (N_5,In_599,In_1251);
or U6 (N_6,In_869,In_782);
or U7 (N_7,In_1083,In_462);
nor U8 (N_8,In_736,In_426);
and U9 (N_9,In_1074,In_872);
or U10 (N_10,In_1218,In_1401);
nand U11 (N_11,In_473,In_961);
nand U12 (N_12,In_495,In_831);
nand U13 (N_13,In_289,In_1367);
and U14 (N_14,In_980,In_1357);
or U15 (N_15,In_695,In_692);
nor U16 (N_16,In_1077,In_487);
nor U17 (N_17,In_28,In_1084);
and U18 (N_18,In_740,In_678);
nor U19 (N_19,In_227,In_423);
nor U20 (N_20,In_475,In_1116);
or U21 (N_21,In_315,In_52);
and U22 (N_22,In_1360,In_349);
xor U23 (N_23,In_712,In_90);
or U24 (N_24,In_545,In_1049);
or U25 (N_25,In_18,In_529);
or U26 (N_26,In_1220,In_975);
or U27 (N_27,In_367,In_1039);
or U28 (N_28,In_1412,In_705);
nand U29 (N_29,In_1051,In_1333);
and U30 (N_30,In_708,In_54);
nand U31 (N_31,In_342,In_1475);
and U32 (N_32,In_382,In_976);
nand U33 (N_33,In_1462,In_179);
nand U34 (N_34,In_196,In_991);
nand U35 (N_35,In_1303,In_1063);
nand U36 (N_36,In_259,In_45);
nor U37 (N_37,In_1155,In_948);
and U38 (N_38,In_900,In_1359);
or U39 (N_39,In_677,In_15);
nand U40 (N_40,In_152,In_1285);
nand U41 (N_41,In_1375,In_911);
nor U42 (N_42,In_628,In_1210);
xor U43 (N_43,In_1238,In_1252);
or U44 (N_44,In_519,In_504);
nand U45 (N_45,In_1326,In_1400);
and U46 (N_46,In_521,In_861);
and U47 (N_47,In_909,In_58);
nand U48 (N_48,In_1054,In_226);
or U49 (N_49,In_143,In_919);
and U50 (N_50,In_36,In_80);
nand U51 (N_51,In_796,In_459);
nor U52 (N_52,In_140,In_1444);
or U53 (N_53,In_542,In_172);
and U54 (N_54,In_664,In_1082);
and U55 (N_55,In_85,In_1436);
nor U56 (N_56,In_697,In_244);
nor U57 (N_57,In_357,In_67);
nand U58 (N_58,In_1270,In_256);
and U59 (N_59,In_79,In_927);
or U60 (N_60,In_543,In_810);
and U61 (N_61,In_937,In_1448);
or U62 (N_62,In_131,In_1354);
or U63 (N_63,In_1045,In_110);
xnor U64 (N_64,In_1102,In_1065);
or U65 (N_65,In_851,In_1260);
and U66 (N_66,In_1193,In_1026);
or U67 (N_67,In_1300,In_277);
nand U68 (N_68,In_1180,In_807);
nand U69 (N_69,In_1114,In_817);
or U70 (N_70,In_578,In_322);
and U71 (N_71,In_1208,In_921);
nand U72 (N_72,In_512,In_1340);
or U73 (N_73,In_1470,In_764);
or U74 (N_74,In_414,In_1186);
and U75 (N_75,In_1046,In_341);
and U76 (N_76,In_653,In_986);
nor U77 (N_77,In_169,In_1241);
nor U78 (N_78,In_1236,In_1403);
and U79 (N_79,In_444,In_449);
nor U80 (N_80,In_1228,In_1129);
nand U81 (N_81,In_1015,In_729);
nor U82 (N_82,In_1295,In_895);
and U83 (N_83,In_1152,In_1262);
or U84 (N_84,In_317,In_270);
nand U85 (N_85,In_1144,In_307);
nor U86 (N_86,In_432,In_1289);
or U87 (N_87,In_1119,In_126);
and U88 (N_88,In_609,In_759);
and U89 (N_89,In_368,In_274);
or U90 (N_90,In_339,In_1321);
nor U91 (N_91,In_321,In_1488);
nor U92 (N_92,In_1154,In_1429);
nand U93 (N_93,In_1227,In_282);
or U94 (N_94,In_1031,In_508);
nand U95 (N_95,In_1104,In_557);
or U96 (N_96,In_1405,In_896);
nand U97 (N_97,In_384,In_556);
or U98 (N_98,In_1336,In_482);
or U99 (N_99,In_555,In_1491);
nand U100 (N_100,In_990,In_239);
and U101 (N_101,In_538,In_1254);
or U102 (N_102,In_515,In_524);
or U103 (N_103,In_478,In_62);
nor U104 (N_104,In_1174,In_460);
nor U105 (N_105,In_1398,In_271);
nand U106 (N_106,In_446,In_48);
and U107 (N_107,In_1131,In_1199);
nand U108 (N_108,In_477,In_290);
or U109 (N_109,In_1040,In_730);
nor U110 (N_110,In_1299,In_252);
nand U111 (N_111,In_1107,In_1120);
or U112 (N_112,In_1277,In_1351);
nand U113 (N_113,In_560,In_607);
or U114 (N_114,In_1346,In_228);
and U115 (N_115,In_928,In_617);
nand U116 (N_116,In_669,In_602);
nand U117 (N_117,In_280,In_343);
and U118 (N_118,In_798,In_157);
xor U119 (N_119,In_1279,In_1173);
and U120 (N_120,In_993,In_1368);
and U121 (N_121,In_217,In_835);
nor U122 (N_122,In_1133,In_1147);
nand U123 (N_123,In_206,In_564);
or U124 (N_124,In_1142,In_588);
and U125 (N_125,In_1485,In_1110);
nand U126 (N_126,In_610,In_758);
and U127 (N_127,In_1467,In_1306);
or U128 (N_128,In_335,In_293);
nand U129 (N_129,In_496,In_1033);
or U130 (N_130,In_885,In_636);
nand U131 (N_131,In_209,In_1290);
or U132 (N_132,In_767,In_1060);
nor U133 (N_133,In_1387,In_950);
and U134 (N_134,In_46,In_979);
nand U135 (N_135,In_88,In_89);
or U136 (N_136,In_591,In_888);
or U137 (N_137,In_940,In_621);
nand U138 (N_138,In_878,In_75);
nand U139 (N_139,In_777,In_198);
nor U140 (N_140,In_1064,In_311);
nand U141 (N_141,In_1059,In_241);
or U142 (N_142,In_1170,In_704);
or U143 (N_143,In_631,In_667);
nand U144 (N_144,In_884,In_283);
and U145 (N_145,In_1474,In_684);
or U146 (N_146,In_313,In_1447);
nand U147 (N_147,In_175,In_1205);
nand U148 (N_148,In_957,In_399);
nand U149 (N_149,In_1006,In_340);
nor U150 (N_150,In_1258,In_64);
and U151 (N_151,In_1003,In_419);
nor U152 (N_152,In_1294,In_845);
or U153 (N_153,In_571,In_1231);
or U154 (N_154,In_405,In_517);
and U155 (N_155,In_800,In_220);
or U156 (N_156,In_467,In_344);
or U157 (N_157,In_520,In_576);
nand U158 (N_158,In_559,In_106);
and U159 (N_159,In_532,In_1394);
or U160 (N_160,In_1203,In_379);
or U161 (N_161,In_424,In_1344);
nand U162 (N_162,In_123,In_395);
and U163 (N_163,In_1292,In_101);
or U164 (N_164,In_371,In_587);
nor U165 (N_165,In_14,In_305);
nor U166 (N_166,In_491,In_431);
and U167 (N_167,In_37,In_332);
or U168 (N_168,In_99,In_943);
or U169 (N_169,In_102,In_505);
or U170 (N_170,In_325,In_73);
nor U171 (N_171,In_665,In_1000);
and U172 (N_172,In_425,In_246);
xor U173 (N_173,In_1349,In_530);
and U174 (N_174,In_49,In_1126);
or U175 (N_175,In_886,In_1420);
and U176 (N_176,In_1019,In_1141);
nand U177 (N_177,In_378,In_1089);
nor U178 (N_178,In_867,In_9);
and U179 (N_179,In_319,In_78);
xnor U180 (N_180,In_1053,In_903);
nor U181 (N_181,In_1092,In_215);
or U182 (N_182,In_369,In_57);
and U183 (N_183,In_1023,In_1156);
xor U184 (N_184,In_563,In_1149);
and U185 (N_185,In_794,In_128);
or U186 (N_186,In_502,In_995);
or U187 (N_187,In_1148,In_375);
and U188 (N_188,In_178,In_1140);
nand U189 (N_189,In_1011,In_1318);
and U190 (N_190,In_1005,In_47);
nand U191 (N_191,In_1305,In_204);
and U192 (N_192,In_871,In_352);
nand U193 (N_193,In_176,In_946);
nor U194 (N_194,In_31,In_1069);
nand U195 (N_195,In_1062,In_1308);
nand U196 (N_196,In_1445,In_522);
nor U197 (N_197,In_1312,In_476);
or U198 (N_198,In_680,In_968);
nor U199 (N_199,In_163,In_1271);
nand U200 (N_200,In_213,In_1438);
and U201 (N_201,In_601,In_744);
nand U202 (N_202,In_233,In_612);
and U203 (N_203,In_1009,In_659);
nor U204 (N_204,In_177,In_651);
or U205 (N_205,In_655,In_523);
nor U206 (N_206,In_774,In_435);
nor U207 (N_207,In_398,In_258);
and U208 (N_208,In_797,In_925);
nor U209 (N_209,In_348,In_201);
nor U210 (N_210,In_168,In_535);
and U211 (N_211,In_565,In_1284);
and U212 (N_212,In_358,In_1109);
or U213 (N_213,In_194,In_267);
nand U214 (N_214,In_922,In_848);
nand U215 (N_215,In_819,In_732);
nand U216 (N_216,In_1150,In_595);
and U217 (N_217,In_1212,In_1386);
and U218 (N_218,In_96,In_967);
and U219 (N_219,In_1449,In_539);
and U220 (N_220,In_1450,In_68);
nor U221 (N_221,In_713,In_1073);
nand U222 (N_222,In_634,In_982);
nor U223 (N_223,In_768,In_639);
nor U224 (N_224,In_1416,In_860);
nor U225 (N_225,In_1087,In_618);
nand U226 (N_226,In_1166,In_753);
or U227 (N_227,In_944,In_1391);
nor U228 (N_228,In_1272,In_722);
or U229 (N_229,In_670,In_159);
or U230 (N_230,In_873,In_323);
nand U231 (N_231,In_623,In_723);
nand U232 (N_232,In_827,In_1280);
nor U233 (N_233,In_1433,In_854);
nor U234 (N_234,In_144,In_686);
and U235 (N_235,In_912,In_361);
and U236 (N_236,In_39,In_370);
or U237 (N_237,In_1377,In_403);
nor U238 (N_238,In_1399,In_81);
or U239 (N_239,In_589,In_908);
nand U240 (N_240,In_973,In_702);
nor U241 (N_241,In_297,In_471);
or U242 (N_242,In_1244,In_897);
or U243 (N_243,In_1163,In_642);
or U244 (N_244,In_996,In_825);
and U245 (N_245,In_799,In_1362);
or U246 (N_246,In_1028,In_404);
xnor U247 (N_247,In_528,In_540);
nand U248 (N_248,In_125,In_1230);
nor U249 (N_249,In_1024,In_1493);
nand U250 (N_250,In_974,In_1437);
or U251 (N_251,In_720,In_1313);
nand U252 (N_252,In_983,In_1421);
and U253 (N_253,In_71,In_372);
or U254 (N_254,In_1101,In_129);
nor U255 (N_255,In_1128,In_770);
and U256 (N_256,In_939,In_314);
and U257 (N_257,In_355,In_436);
nor U258 (N_258,In_1257,In_721);
nand U259 (N_259,In_998,In_1393);
nor U260 (N_260,In_1428,In_813);
and U261 (N_261,In_224,In_422);
or U262 (N_262,In_262,In_468);
nand U263 (N_263,In_97,In_192);
nor U264 (N_264,In_229,In_1130);
nand U265 (N_265,In_119,In_706);
and U266 (N_266,In_386,In_541);
nand U267 (N_267,In_966,In_1188);
xnor U268 (N_268,In_1476,In_1219);
or U269 (N_269,In_1278,In_142);
and U270 (N_270,In_1430,In_812);
or U271 (N_271,In_1389,In_166);
or U272 (N_272,In_1058,In_211);
xnor U273 (N_273,In_1253,In_1309);
nand U274 (N_274,In_23,In_66);
and U275 (N_275,In_626,In_1465);
or U276 (N_276,In_733,In_972);
nor U277 (N_277,In_20,In_98);
or U278 (N_278,In_586,In_572);
nor U279 (N_279,In_509,In_1317);
nand U280 (N_280,In_248,In_132);
and U281 (N_281,In_890,In_296);
nor U282 (N_282,In_445,In_999);
nand U283 (N_283,In_1431,In_29);
and U284 (N_284,In_850,In_1217);
nor U285 (N_285,In_818,In_1160);
and U286 (N_286,In_1079,In_581);
nand U287 (N_287,In_707,In_109);
and U288 (N_288,In_593,In_841);
or U289 (N_289,In_455,In_510);
and U290 (N_290,In_223,In_1392);
or U291 (N_291,In_1406,In_292);
nand U292 (N_292,In_494,In_1464);
and U293 (N_293,In_1135,In_786);
and U294 (N_294,In_1117,In_373);
nor U295 (N_295,In_737,In_329);
nand U296 (N_296,In_795,In_1177);
or U297 (N_297,In_1200,In_1215);
nand U298 (N_298,In_489,In_133);
nor U299 (N_299,In_1407,In_208);
and U300 (N_300,In_676,In_826);
nor U301 (N_301,In_1322,In_42);
and U302 (N_302,In_646,In_1078);
or U303 (N_303,In_1042,In_658);
nand U304 (N_304,In_981,In_1425);
and U305 (N_305,In_225,In_454);
nor U306 (N_306,In_1094,In_934);
nor U307 (N_307,In_690,In_619);
nor U308 (N_308,In_1249,In_624);
and U309 (N_309,In_1432,In_1025);
nor U310 (N_310,In_547,In_1334);
nand U311 (N_311,In_197,In_965);
or U312 (N_312,In_497,In_456);
nand U313 (N_313,In_304,In_1418);
xnor U314 (N_314,In_1029,In_526);
and U315 (N_315,In_881,In_1480);
xnor U316 (N_316,In_1191,In_838);
or U317 (N_317,In_933,In_245);
and U318 (N_318,In_264,In_394);
or U319 (N_319,In_134,In_450);
nand U320 (N_320,In_1224,In_709);
nand U321 (N_321,In_440,In_181);
nand U322 (N_322,In_474,In_108);
and U323 (N_323,In_691,In_1001);
nand U324 (N_324,In_1337,In_117);
nand U325 (N_325,In_1454,In_683);
or U326 (N_326,In_1457,In_410);
nand U327 (N_327,In_1484,In_115);
and U328 (N_328,In_750,In_789);
or U329 (N_329,In_992,In_1380);
or U330 (N_330,In_276,In_387);
nor U331 (N_331,In_429,In_150);
nand U332 (N_332,In_597,In_4);
or U333 (N_333,In_1243,In_1355);
or U334 (N_334,In_657,In_696);
nand U335 (N_335,In_1332,In_1201);
and U336 (N_336,In_1410,In_916);
nor U337 (N_337,In_853,In_785);
nand U338 (N_338,In_1036,In_630);
or U339 (N_339,In_457,In_1211);
or U340 (N_340,In_44,In_592);
or U341 (N_341,In_453,In_779);
or U342 (N_342,In_1497,In_633);
nand U343 (N_343,In_1466,In_230);
or U344 (N_344,In_552,In_420);
or U345 (N_345,In_1273,In_120);
or U346 (N_346,In_1451,In_374);
nor U347 (N_347,In_735,In_407);
nand U348 (N_348,In_151,In_660);
nor U349 (N_349,In_1370,In_920);
nand U350 (N_350,In_865,In_745);
nand U351 (N_351,In_1477,In_1213);
nor U352 (N_352,In_33,In_1250);
or U353 (N_353,In_366,In_30);
nand U354 (N_354,In_682,In_1136);
or U355 (N_355,In_481,In_324);
nand U356 (N_356,In_406,In_354);
nor U357 (N_357,In_441,In_942);
and U358 (N_358,In_913,In_606);
nor U359 (N_359,In_889,In_34);
nor U360 (N_360,In_1283,In_480);
nand U361 (N_361,In_149,In_1434);
or U362 (N_362,In_1175,In_1364);
nor U363 (N_363,In_1441,In_1343);
nor U364 (N_364,In_27,In_1194);
or U365 (N_365,In_433,In_156);
nand U366 (N_366,In_347,In_1293);
and U367 (N_367,In_1132,In_1134);
xor U368 (N_368,In_278,In_611);
nand U369 (N_369,In_275,In_479);
nand U370 (N_370,In_493,In_193);
nor U371 (N_371,In_1324,In_0);
nor U372 (N_372,In_1468,In_629);
or U373 (N_373,In_1323,In_1331);
or U374 (N_374,In_718,In_463);
nor U375 (N_375,In_1106,In_310);
nand U376 (N_376,In_1121,In_671);
or U377 (N_377,In_1288,In_882);
xor U378 (N_378,In_546,In_566);
nand U379 (N_379,In_856,In_364);
and U380 (N_380,In_823,In_1145);
and U381 (N_381,In_1371,In_625);
nand U382 (N_382,In_739,In_235);
and U383 (N_383,In_53,In_362);
nor U384 (N_384,In_1266,In_814);
or U385 (N_385,In_1187,In_1097);
nand U386 (N_386,In_824,In_762);
or U387 (N_387,In_1137,In_1435);
or U388 (N_388,In_1171,In_685);
nand U389 (N_389,In_257,In_183);
nand U390 (N_390,In_174,In_1204);
and U391 (N_391,In_548,In_533);
and U392 (N_392,In_537,In_299);
nand U393 (N_393,In_513,In_579);
nor U394 (N_394,In_1189,In_413);
or U395 (N_395,In_1264,In_331);
nor U396 (N_396,In_1426,In_295);
and U397 (N_397,In_21,In_318);
nand U398 (N_398,In_356,In_842);
or U399 (N_399,In_1460,In_833);
nor U400 (N_400,In_1338,In_1182);
and U401 (N_401,In_139,In_514);
and U402 (N_402,In_1138,In_1027);
and U403 (N_403,In_641,In_288);
and U404 (N_404,In_8,In_1122);
or U405 (N_405,In_815,In_1395);
nand U406 (N_406,In_963,In_162);
nand U407 (N_407,In_931,In_852);
or U408 (N_408,In_839,In_719);
nand U409 (N_409,In_914,In_747);
nand U410 (N_410,In_901,In_346);
nor U411 (N_411,In_917,In_1408);
nor U412 (N_412,In_1030,In_1458);
or U413 (N_413,In_247,In_859);
nor U414 (N_414,In_200,In_1179);
nand U415 (N_415,In_801,In_766);
xnor U416 (N_416,In_350,In_932);
and U417 (N_417,In_742,In_1446);
and U418 (N_418,In_1195,In_1172);
or U419 (N_419,In_613,In_811);
nand U420 (N_420,In_442,In_1055);
or U421 (N_421,In_1178,In_1329);
and U422 (N_422,In_1311,In_1350);
or U423 (N_423,In_1381,In_534);
nand U424 (N_424,In_65,In_844);
and U425 (N_425,In_401,In_1330);
nand U426 (N_426,In_632,In_893);
and U427 (N_427,In_16,In_1268);
xor U428 (N_428,In_112,In_171);
or U429 (N_429,In_647,In_1274);
or U430 (N_430,In_250,In_1452);
or U431 (N_431,In_834,In_1415);
nor U432 (N_432,In_1124,In_752);
nor U433 (N_433,In_1052,In_771);
xor U434 (N_434,In_960,In_124);
or U435 (N_435,In_1383,In_716);
nor U436 (N_436,In_1048,In_905);
and U437 (N_437,In_94,In_924);
nor U438 (N_438,In_418,In_816);
and U439 (N_439,In_1103,In_365);
nor U440 (N_440,In_1081,In_580);
nand U441 (N_441,In_55,In_1453);
or U442 (N_442,In_11,In_121);
xnor U443 (N_443,In_130,In_787);
and U444 (N_444,In_568,In_714);
or U445 (N_445,In_506,In_536);
nand U446 (N_446,In_699,In_72);
nand U447 (N_447,In_91,In_221);
nand U448 (N_448,In_681,In_605);
nor U449 (N_449,In_945,In_644);
nor U450 (N_450,In_302,In_265);
nand U451 (N_451,In_1225,In_427);
and U452 (N_452,In_1255,In_421);
or U453 (N_453,In_1269,In_1198);
and U454 (N_454,In_1265,In_74);
or U455 (N_455,In_428,In_964);
nor U456 (N_456,In_1096,In_666);
or U457 (N_457,In_154,In_1164);
or U458 (N_458,In_465,In_469);
or U459 (N_459,In_87,In_864);
nand U460 (N_460,In_567,In_769);
nor U461 (N_461,In_843,In_281);
nand U462 (N_462,In_32,In_1409);
nand U463 (N_463,In_1276,In_1226);
nand U464 (N_464,In_675,In_1261);
and U465 (N_465,In_391,In_1022);
nand U466 (N_466,In_312,In_955);
nor U467 (N_467,In_689,In_448);
xnor U468 (N_468,In_652,In_847);
or U469 (N_469,In_649,In_158);
nand U470 (N_470,In_59,In_389);
or U471 (N_471,In_748,In_1267);
or U472 (N_472,In_904,In_412);
or U473 (N_473,In_1108,In_439);
or U474 (N_474,In_1115,In_906);
nand U475 (N_475,In_1459,In_978);
and U476 (N_476,In_327,In_1123);
and U477 (N_477,In_791,In_205);
or U478 (N_478,In_1216,In_231);
nor U479 (N_479,In_590,In_415);
nand U480 (N_480,In_701,In_353);
or U481 (N_481,In_531,In_1202);
nor U482 (N_482,In_499,In_1314);
nand U483 (N_483,In_1127,In_584);
nor U484 (N_484,In_1068,In_40);
or U485 (N_485,In_1411,In_1012);
or U486 (N_486,In_821,In_1456);
or U487 (N_487,In_958,In_784);
or U488 (N_488,In_182,In_947);
nand U489 (N_489,In_338,In_594);
and U490 (N_490,In_1043,In_360);
nand U491 (N_491,In_1327,In_254);
nand U492 (N_492,In_635,In_105);
nor U493 (N_493,In_577,In_284);
nand U494 (N_494,In_820,In_69);
nor U495 (N_495,In_77,In_236);
nor U496 (N_496,In_899,In_1146);
nor U497 (N_497,In_483,In_351);
or U498 (N_498,In_243,In_122);
and U499 (N_499,In_727,In_242);
or U500 (N_500,In_381,In_167);
nand U501 (N_501,In_12,In_596);
and U502 (N_502,In_84,In_668);
or U503 (N_503,In_754,In_165);
nor U504 (N_504,In_1017,In_734);
nand U505 (N_505,In_1287,In_1489);
and U506 (N_506,In_760,In_1486);
and U507 (N_507,In_1007,In_604);
and U508 (N_508,In_1099,In_1176);
nor U509 (N_509,In_656,In_443);
nor U510 (N_510,In_806,In_461);
nand U511 (N_511,In_507,In_918);
and U512 (N_512,In_488,In_1157);
or U513 (N_513,In_1328,In_416);
or U514 (N_514,In_376,In_1032);
nor U515 (N_515,In_638,In_114);
or U516 (N_516,In_392,In_1296);
nand U517 (N_517,In_1483,In_1196);
nor U518 (N_518,In_498,In_1192);
or U519 (N_519,In_287,In_56);
nand U520 (N_520,In_837,In_1056);
or U521 (N_521,In_710,In_1353);
and U522 (N_522,In_285,In_1034);
or U523 (N_523,In_778,In_127);
or U524 (N_524,In_396,In_1307);
nor U525 (N_525,In_1365,In_1095);
nand U526 (N_526,In_830,In_1413);
and U527 (N_527,In_189,In_500);
nand U528 (N_528,In_408,In_598);
nand U529 (N_529,In_263,In_1281);
and U530 (N_530,In_393,In_1315);
xor U531 (N_531,In_83,In_954);
nand U532 (N_532,In_765,In_35);
xor U533 (N_533,In_615,In_180);
and U534 (N_534,In_385,In_1348);
nor U535 (N_535,In_1037,In_1378);
nand U536 (N_536,In_1263,In_279);
nand U537 (N_537,In_1209,In_212);
and U538 (N_538,In_1190,In_452);
and U539 (N_539,In_627,In_1259);
nor U540 (N_540,In_1010,In_118);
or U541 (N_541,In_260,In_1158);
or U542 (N_542,In_1221,In_1374);
nor U543 (N_543,In_199,In_775);
or U544 (N_544,In_1206,In_1390);
or U545 (N_545,In_1047,In_291);
nand U546 (N_546,In_472,In_1071);
or U547 (N_547,In_959,In_1085);
or U548 (N_548,In_698,In_1455);
and U549 (N_549,In_300,In_320);
and U550 (N_550,In_334,In_1020);
and U551 (N_551,In_190,In_1361);
nor U552 (N_552,In_447,In_997);
nand U553 (N_553,In_971,In_1345);
nand U554 (N_554,In_808,In_756);
or U555 (N_555,In_987,In_1008);
nand U556 (N_556,In_1018,In_25);
nor U557 (N_557,In_616,In_654);
nand U558 (N_558,In_1479,In_116);
or U559 (N_559,In_1183,In_328);
nand U560 (N_560,In_1478,In_294);
and U561 (N_561,In_527,In_846);
and U562 (N_562,In_1061,In_688);
nor U563 (N_563,In_232,In_863);
nor U564 (N_564,In_146,In_793);
or U565 (N_565,In_561,In_1139);
or U566 (N_566,In_1044,In_1075);
nor U567 (N_567,In_3,In_1297);
nor U568 (N_568,In_1233,In_553);
and U569 (N_569,In_113,In_525);
nor U570 (N_570,In_1050,In_929);
nand U571 (N_571,In_1214,In_1161);
or U572 (N_572,In_1376,In_1067);
nand U573 (N_573,In_822,In_1207);
xnor U574 (N_574,In_1242,In_222);
nand U575 (N_575,In_608,In_1382);
and U576 (N_576,In_783,In_41);
or U577 (N_577,In_952,In_749);
nor U578 (N_578,In_1494,In_216);
or U579 (N_579,In_1235,In_26);
nor U580 (N_580,In_989,In_781);
nand U581 (N_581,In_397,In_1404);
nand U582 (N_582,In_1363,In_6);
nand U583 (N_583,In_17,In_788);
nand U584 (N_584,In_1341,In_700);
and U585 (N_585,In_1417,In_876);
nand U586 (N_586,In_1197,In_1419);
and U587 (N_587,In_490,In_486);
nand U588 (N_588,In_195,In_1245);
or U589 (N_589,In_1492,In_437);
and U590 (N_590,In_191,In_1072);
and U591 (N_591,In_60,In_10);
and U592 (N_592,In_663,In_1397);
and U593 (N_593,In_170,In_234);
nor U594 (N_594,In_614,In_86);
nand U595 (N_595,In_1222,In_1310);
nand U596 (N_596,In_1301,In_1442);
or U597 (N_597,In_907,In_1379);
nand U598 (N_598,In_141,In_1358);
nand U599 (N_599,In_503,In_1165);
nand U600 (N_600,In_269,In_380);
or U601 (N_601,In_1004,In_1090);
nor U602 (N_602,In_544,In_1111);
nand U603 (N_603,In_301,In_400);
or U604 (N_604,In_1237,In_50);
nor U605 (N_605,In_792,In_741);
or U606 (N_606,In_485,In_751);
and U607 (N_607,In_1057,In_1463);
nand U608 (N_608,In_866,In_743);
nor U609 (N_609,In_237,In_188);
nand U610 (N_610,In_249,In_1481);
or U611 (N_611,In_1366,In_309);
and U612 (N_612,In_891,In_910);
nor U613 (N_613,In_253,In_377);
and U614 (N_614,In_466,In_832);
or U615 (N_615,In_1473,In_574);
nor U616 (N_616,In_703,In_969);
or U617 (N_617,In_409,In_516);
and U618 (N_618,In_883,In_214);
and U619 (N_619,In_22,In_1339);
and U620 (N_620,In_725,In_898);
nand U621 (N_621,In_1246,In_1461);
or U622 (N_622,In_111,In_1372);
nor U623 (N_623,In_337,In_207);
nor U624 (N_624,In_155,In_1080);
and U625 (N_625,In_687,In_1427);
or U626 (N_626,In_511,In_1229);
and U627 (N_627,In_390,In_238);
nand U628 (N_628,In_186,In_1091);
and U629 (N_629,In_941,In_518);
and U630 (N_630,In_902,In_1070);
nor U631 (N_631,In_1490,In_363);
nand U632 (N_632,In_1275,In_1184);
nand U633 (N_633,In_870,In_1482);
nand U634 (N_634,In_970,In_1369);
nand U635 (N_635,In_1499,In_603);
nand U636 (N_636,In_1113,In_1240);
nand U637 (N_637,In_829,In_76);
or U638 (N_638,In_438,In_1385);
and U639 (N_639,In_1086,In_773);
and U640 (N_640,In_1002,In_308);
nor U641 (N_641,In_95,In_160);
or U642 (N_642,In_936,In_1347);
nand U643 (N_643,In_138,In_19);
and U644 (N_644,In_1013,In_38);
nor U645 (N_645,In_145,In_877);
nor U646 (N_646,In_585,In_746);
nor U647 (N_647,In_887,In_161);
and U648 (N_648,In_674,In_935);
and U649 (N_649,In_1256,In_104);
and U650 (N_650,In_185,In_763);
or U651 (N_651,In_336,In_92);
and U652 (N_652,In_637,In_549);
nor U653 (N_653,In_1302,In_5);
xor U654 (N_654,In_894,In_724);
and U655 (N_655,In_1422,In_492);
nor U656 (N_656,In_985,In_266);
nand U657 (N_657,In_484,In_728);
or U658 (N_658,In_1496,In_643);
nand U659 (N_659,In_135,In_359);
nor U660 (N_660,In_501,In_451);
nand U661 (N_661,In_1439,In_880);
nand U662 (N_662,In_1498,In_1472);
and U663 (N_663,In_1440,In_662);
and U664 (N_664,In_1291,In_550);
nor U665 (N_665,In_1316,In_956);
and U666 (N_666,In_303,In_43);
and U667 (N_667,In_1402,In_107);
or U668 (N_668,In_272,In_790);
or U669 (N_669,In_776,In_1443);
and U670 (N_670,In_1105,In_836);
nor U671 (N_671,In_458,In_600);
nor U672 (N_672,In_875,In_13);
or U673 (N_673,In_1143,In_148);
nand U674 (N_674,In_383,In_273);
xor U675 (N_675,In_24,In_915);
or U676 (N_676,In_240,In_1388);
nor U677 (N_677,In_757,In_1181);
or U678 (N_678,In_1247,In_137);
nor U679 (N_679,In_645,In_570);
and U680 (N_680,In_218,In_1471);
nand U681 (N_681,In_82,In_1168);
or U682 (N_682,In_780,In_575);
nor U683 (N_683,In_187,In_1088);
nor U684 (N_684,In_330,In_411);
or U685 (N_685,In_804,In_1469);
and U686 (N_686,In_316,In_761);
nand U687 (N_687,In_430,In_2);
or U688 (N_688,In_558,In_93);
and U689 (N_689,In_255,In_717);
nor U690 (N_690,In_672,In_926);
and U691 (N_691,In_840,In_1424);
nor U692 (N_692,In_650,In_136);
or U693 (N_693,In_551,In_715);
and U694 (N_694,In_1373,In_1098);
nand U695 (N_695,In_1066,In_173);
and U696 (N_696,In_620,In_772);
or U697 (N_697,In_953,In_1396);
nand U698 (N_698,In_388,In_147);
nand U699 (N_699,In_984,In_61);
or U700 (N_700,In_1286,In_210);
nand U701 (N_701,In_203,In_1093);
or U702 (N_702,In_202,In_1487);
and U703 (N_703,In_738,In_988);
nand U704 (N_704,In_1325,In_622);
nand U705 (N_705,In_582,In_673);
and U706 (N_706,In_1153,In_1014);
or U707 (N_707,In_858,In_949);
nand U708 (N_708,In_417,In_70);
and U709 (N_709,In_855,In_802);
and U710 (N_710,In_693,In_726);
nand U711 (N_711,In_879,In_1021);
or U712 (N_712,In_268,In_1234);
nor U713 (N_713,In_326,In_1159);
nand U714 (N_714,In_470,In_977);
nor U715 (N_715,In_1232,In_1352);
or U716 (N_716,In_153,In_345);
nor U717 (N_717,In_103,In_1169);
and U718 (N_718,In_1239,In_583);
and U719 (N_719,In_857,In_962);
nor U720 (N_720,In_261,In_1118);
or U721 (N_721,In_640,In_1298);
or U722 (N_722,In_679,In_755);
nand U723 (N_723,In_100,In_562);
or U724 (N_724,In_1,In_1304);
nor U725 (N_725,In_805,In_1162);
and U726 (N_726,In_648,In_298);
or U727 (N_727,In_731,In_1223);
and U728 (N_728,In_219,In_874);
and U729 (N_729,In_1038,In_573);
nor U730 (N_730,In_1076,In_434);
nand U731 (N_731,In_63,In_286);
nand U732 (N_732,In_1016,In_251);
and U733 (N_733,In_1320,In_51);
nor U734 (N_734,In_164,In_1035);
or U735 (N_735,In_868,In_1100);
and U736 (N_736,In_994,In_1335);
nor U737 (N_737,In_661,In_1414);
nor U738 (N_738,In_1319,In_892);
nor U739 (N_739,In_938,In_1495);
and U740 (N_740,In_1185,In_306);
and U741 (N_741,In_849,In_951);
and U742 (N_742,In_1282,In_1342);
nor U743 (N_743,In_7,In_923);
or U744 (N_744,In_1112,In_1167);
or U745 (N_745,In_402,In_1248);
and U746 (N_746,In_862,In_711);
nor U747 (N_747,In_809,In_1151);
nor U748 (N_748,In_554,In_569);
nor U749 (N_749,In_184,In_1423);
nor U750 (N_750,N_393,N_502);
nor U751 (N_751,N_70,N_317);
and U752 (N_752,N_357,N_470);
nor U753 (N_753,N_84,N_630);
or U754 (N_754,N_703,N_244);
and U755 (N_755,N_295,N_658);
nand U756 (N_756,N_566,N_369);
nor U757 (N_757,N_461,N_222);
xnor U758 (N_758,N_367,N_206);
and U759 (N_759,N_426,N_648);
or U760 (N_760,N_26,N_319);
and U761 (N_761,N_72,N_624);
and U762 (N_762,N_52,N_446);
or U763 (N_763,N_242,N_79);
nor U764 (N_764,N_737,N_23);
or U765 (N_765,N_282,N_438);
nand U766 (N_766,N_322,N_452);
or U767 (N_767,N_278,N_730);
and U768 (N_768,N_20,N_439);
nor U769 (N_769,N_371,N_137);
nor U770 (N_770,N_35,N_632);
and U771 (N_771,N_541,N_237);
nand U772 (N_772,N_229,N_734);
nor U773 (N_773,N_126,N_11);
nor U774 (N_774,N_557,N_144);
xor U775 (N_775,N_329,N_447);
xnor U776 (N_776,N_379,N_216);
nor U777 (N_777,N_559,N_299);
or U778 (N_778,N_655,N_440);
nor U779 (N_779,N_611,N_350);
or U780 (N_780,N_238,N_56);
nand U781 (N_781,N_163,N_480);
and U782 (N_782,N_153,N_540);
nand U783 (N_783,N_558,N_594);
or U784 (N_784,N_701,N_610);
or U785 (N_785,N_117,N_489);
or U786 (N_786,N_10,N_335);
nor U787 (N_787,N_492,N_526);
or U788 (N_788,N_529,N_726);
nor U789 (N_789,N_380,N_310);
nand U790 (N_790,N_241,N_622);
nor U791 (N_791,N_58,N_661);
or U792 (N_792,N_285,N_161);
and U793 (N_793,N_75,N_128);
and U794 (N_794,N_93,N_194);
nor U795 (N_795,N_743,N_719);
nor U796 (N_796,N_571,N_81);
nor U797 (N_797,N_520,N_441);
and U798 (N_798,N_16,N_182);
and U799 (N_799,N_718,N_459);
and U800 (N_800,N_479,N_284);
xor U801 (N_801,N_288,N_254);
or U802 (N_802,N_110,N_286);
nand U803 (N_803,N_215,N_3);
and U804 (N_804,N_29,N_454);
or U805 (N_805,N_255,N_619);
and U806 (N_806,N_443,N_564);
and U807 (N_807,N_672,N_149);
and U808 (N_808,N_736,N_381);
or U809 (N_809,N_749,N_108);
or U810 (N_810,N_160,N_606);
nand U811 (N_811,N_535,N_568);
or U812 (N_812,N_677,N_590);
and U813 (N_813,N_476,N_349);
nor U814 (N_814,N_689,N_323);
or U815 (N_815,N_530,N_424);
and U816 (N_816,N_316,N_275);
nand U817 (N_817,N_633,N_145);
nand U818 (N_818,N_266,N_733);
nand U819 (N_819,N_707,N_665);
or U820 (N_820,N_686,N_469);
nand U821 (N_821,N_245,N_724);
nand U822 (N_822,N_198,N_567);
and U823 (N_823,N_748,N_544);
and U824 (N_824,N_217,N_585);
xnor U825 (N_825,N_106,N_577);
and U826 (N_826,N_593,N_346);
nand U827 (N_827,N_490,N_235);
or U828 (N_828,N_265,N_462);
and U829 (N_829,N_385,N_18);
or U830 (N_830,N_460,N_400);
or U831 (N_831,N_192,N_586);
nor U832 (N_832,N_337,N_671);
and U833 (N_833,N_725,N_25);
nand U834 (N_834,N_437,N_642);
and U835 (N_835,N_634,N_220);
nand U836 (N_836,N_214,N_428);
and U837 (N_837,N_212,N_451);
and U838 (N_838,N_236,N_414);
and U839 (N_839,N_727,N_146);
nor U840 (N_840,N_158,N_271);
nor U841 (N_841,N_272,N_30);
xor U842 (N_842,N_488,N_359);
nand U843 (N_843,N_692,N_134);
nor U844 (N_844,N_493,N_184);
nor U845 (N_845,N_289,N_304);
nand U846 (N_846,N_269,N_668);
or U847 (N_847,N_679,N_280);
nor U848 (N_848,N_699,N_496);
and U849 (N_849,N_697,N_739);
nand U850 (N_850,N_458,N_62);
nor U851 (N_851,N_86,N_183);
and U852 (N_852,N_456,N_24);
or U853 (N_853,N_100,N_449);
nand U854 (N_854,N_177,N_711);
and U855 (N_855,N_53,N_616);
and U856 (N_856,N_195,N_42);
or U857 (N_857,N_554,N_178);
and U858 (N_858,N_247,N_200);
nand U859 (N_859,N_687,N_366);
nand U860 (N_860,N_419,N_125);
and U861 (N_861,N_409,N_407);
or U862 (N_862,N_120,N_166);
nand U863 (N_863,N_355,N_98);
and U864 (N_864,N_293,N_170);
nor U865 (N_865,N_623,N_403);
nor U866 (N_866,N_327,N_531);
nor U867 (N_867,N_645,N_67);
nor U868 (N_868,N_64,N_60);
and U869 (N_869,N_475,N_15);
and U870 (N_870,N_6,N_252);
or U871 (N_871,N_342,N_694);
nor U872 (N_872,N_88,N_68);
or U873 (N_873,N_372,N_191);
nor U874 (N_874,N_408,N_429);
or U875 (N_875,N_542,N_172);
xnor U876 (N_876,N_155,N_76);
nand U877 (N_877,N_378,N_308);
nand U878 (N_878,N_651,N_621);
and U879 (N_879,N_71,N_735);
or U880 (N_880,N_270,N_410);
or U881 (N_881,N_2,N_499);
and U882 (N_882,N_225,N_576);
nand U883 (N_883,N_239,N_325);
and U884 (N_884,N_448,N_109);
nor U885 (N_885,N_747,N_599);
or U886 (N_886,N_392,N_620);
and U887 (N_887,N_486,N_313);
and U888 (N_888,N_296,N_165);
or U889 (N_889,N_139,N_545);
nor U890 (N_890,N_706,N_485);
nand U891 (N_891,N_96,N_442);
nor U892 (N_892,N_181,N_376);
or U893 (N_893,N_675,N_133);
or U894 (N_894,N_436,N_267);
xor U895 (N_895,N_107,N_124);
nand U896 (N_896,N_111,N_364);
or U897 (N_897,N_618,N_208);
nor U898 (N_898,N_179,N_387);
or U899 (N_899,N_135,N_383);
nand U900 (N_900,N_80,N_710);
and U901 (N_901,N_274,N_142);
or U902 (N_902,N_151,N_136);
nand U903 (N_903,N_639,N_487);
nand U904 (N_904,N_539,N_202);
nand U905 (N_905,N_48,N_331);
and U906 (N_906,N_22,N_465);
or U907 (N_907,N_547,N_396);
or U908 (N_908,N_92,N_517);
or U909 (N_909,N_680,N_406);
nand U910 (N_910,N_629,N_532);
or U911 (N_911,N_116,N_563);
and U912 (N_912,N_28,N_457);
and U913 (N_913,N_552,N_555);
and U914 (N_914,N_343,N_17);
or U915 (N_915,N_223,N_533);
nand U916 (N_916,N_77,N_249);
or U917 (N_917,N_649,N_123);
and U918 (N_918,N_119,N_625);
and U919 (N_919,N_418,N_481);
and U920 (N_920,N_102,N_505);
and U921 (N_921,N_420,N_678);
or U922 (N_922,N_395,N_314);
nand U923 (N_923,N_180,N_13);
or U924 (N_924,N_497,N_307);
nor U925 (N_925,N_641,N_628);
and U926 (N_926,N_444,N_112);
and U927 (N_927,N_669,N_157);
nand U928 (N_928,N_398,N_549);
and U929 (N_929,N_388,N_46);
nor U930 (N_930,N_213,N_691);
and U931 (N_931,N_613,N_695);
or U932 (N_932,N_352,N_4);
nor U933 (N_933,N_305,N_693);
nor U934 (N_934,N_638,N_173);
nor U935 (N_935,N_9,N_391);
or U936 (N_936,N_91,N_562);
nor U937 (N_937,N_131,N_525);
nand U938 (N_938,N_740,N_527);
and U939 (N_939,N_698,N_127);
and U940 (N_940,N_482,N_666);
nor U941 (N_941,N_696,N_315);
or U942 (N_942,N_176,N_292);
or U943 (N_943,N_528,N_521);
nor U944 (N_944,N_513,N_670);
or U945 (N_945,N_643,N_129);
nand U946 (N_946,N_253,N_187);
nand U947 (N_947,N_647,N_654);
nand U948 (N_948,N_41,N_685);
nand U949 (N_949,N_65,N_591);
nor U950 (N_950,N_411,N_660);
or U951 (N_951,N_581,N_543);
or U952 (N_952,N_263,N_659);
xnor U953 (N_953,N_336,N_326);
nand U954 (N_954,N_574,N_422);
and U955 (N_955,N_636,N_344);
nand U956 (N_956,N_330,N_221);
nor U957 (N_957,N_40,N_312);
nor U958 (N_958,N_511,N_358);
nor U959 (N_959,N_508,N_575);
nor U960 (N_960,N_468,N_14);
and U961 (N_961,N_101,N_273);
and U962 (N_962,N_477,N_104);
nand U963 (N_963,N_328,N_589);
nor U964 (N_964,N_537,N_370);
nand U965 (N_965,N_205,N_193);
or U966 (N_966,N_453,N_425);
nor U967 (N_967,N_397,N_363);
or U968 (N_968,N_536,N_31);
nand U969 (N_969,N_59,N_309);
or U970 (N_970,N_431,N_90);
nand U971 (N_971,N_268,N_97);
or U972 (N_972,N_653,N_61);
or U973 (N_973,N_147,N_612);
nor U974 (N_974,N_467,N_494);
or U975 (N_975,N_471,N_230);
or U976 (N_976,N_729,N_251);
nand U977 (N_977,N_744,N_412);
nand U978 (N_978,N_203,N_503);
xor U979 (N_979,N_168,N_302);
or U980 (N_980,N_1,N_12);
or U981 (N_981,N_207,N_580);
and U982 (N_982,N_650,N_44);
and U983 (N_983,N_548,N_261);
or U984 (N_984,N_617,N_132);
or U985 (N_985,N_401,N_510);
and U986 (N_986,N_673,N_375);
nand U987 (N_987,N_47,N_434);
and U988 (N_988,N_340,N_683);
nand U989 (N_989,N_473,N_538);
nor U990 (N_990,N_54,N_394);
nand U991 (N_991,N_89,N_39);
or U992 (N_992,N_297,N_631);
and U993 (N_993,N_377,N_231);
nor U994 (N_994,N_656,N_209);
nor U995 (N_995,N_514,N_421);
and U996 (N_996,N_676,N_279);
nand U997 (N_997,N_228,N_664);
or U998 (N_998,N_351,N_277);
or U999 (N_999,N_43,N_745);
and U1000 (N_1000,N_602,N_85);
or U1001 (N_1001,N_115,N_347);
and U1002 (N_1002,N_584,N_386);
nand U1003 (N_1003,N_332,N_318);
or U1004 (N_1004,N_78,N_171);
and U1005 (N_1005,N_246,N_704);
nand U1006 (N_1006,N_354,N_495);
nor U1007 (N_1007,N_256,N_657);
or U1008 (N_1008,N_402,N_103);
nor U1009 (N_1009,N_500,N_234);
nor U1010 (N_1010,N_188,N_588);
and U1011 (N_1011,N_652,N_51);
or U1012 (N_1012,N_233,N_615);
nand U1013 (N_1013,N_705,N_311);
nand U1014 (N_1014,N_717,N_360);
and U1015 (N_1015,N_515,N_716);
or U1016 (N_1016,N_95,N_50);
nand U1017 (N_1017,N_644,N_150);
nand U1018 (N_1018,N_321,N_413);
and U1019 (N_1019,N_287,N_356);
or U1020 (N_1020,N_162,N_361);
and U1021 (N_1021,N_723,N_374);
and U1022 (N_1022,N_519,N_637);
nand U1023 (N_1023,N_605,N_262);
nor U1024 (N_1024,N_218,N_715);
nand U1025 (N_1025,N_732,N_523);
nand U1026 (N_1026,N_582,N_573);
nand U1027 (N_1027,N_604,N_587);
nand U1028 (N_1028,N_427,N_201);
and U1029 (N_1029,N_74,N_583);
nor U1030 (N_1030,N_708,N_714);
nor U1031 (N_1031,N_722,N_368);
or U1032 (N_1032,N_635,N_159);
xor U1033 (N_1033,N_399,N_507);
or U1034 (N_1034,N_291,N_560);
nor U1035 (N_1035,N_199,N_682);
and U1036 (N_1036,N_569,N_122);
nand U1037 (N_1037,N_713,N_36);
and U1038 (N_1038,N_169,N_667);
nor U1039 (N_1039,N_324,N_250);
nand U1040 (N_1040,N_73,N_338);
and U1041 (N_1041,N_196,N_373);
or U1042 (N_1042,N_353,N_121);
and U1043 (N_1043,N_281,N_45);
or U1044 (N_1044,N_608,N_259);
nor U1045 (N_1045,N_118,N_721);
nor U1046 (N_1046,N_290,N_435);
nand U1047 (N_1047,N_55,N_546);
and U1048 (N_1048,N_164,N_728);
nand U1049 (N_1049,N_186,N_34);
nor U1050 (N_1050,N_138,N_348);
nand U1051 (N_1051,N_211,N_688);
and U1052 (N_1052,N_82,N_501);
nand U1053 (N_1053,N_140,N_483);
nor U1054 (N_1054,N_614,N_333);
or U1055 (N_1055,N_339,N_175);
nor U1056 (N_1056,N_405,N_143);
and U1057 (N_1057,N_301,N_597);
nor U1058 (N_1058,N_226,N_607);
or U1059 (N_1059,N_5,N_491);
and U1060 (N_1060,N_731,N_570);
and U1061 (N_1061,N_524,N_210);
nor U1062 (N_1062,N_684,N_640);
nor U1063 (N_1063,N_445,N_700);
nand U1064 (N_1064,N_463,N_227);
nand U1065 (N_1065,N_113,N_390);
nor U1066 (N_1066,N_709,N_283);
and U1067 (N_1067,N_276,N_601);
and U1068 (N_1068,N_224,N_592);
nor U1069 (N_1069,N_389,N_99);
nand U1070 (N_1070,N_609,N_720);
nor U1071 (N_1071,N_174,N_94);
or U1072 (N_1072,N_478,N_603);
nor U1073 (N_1073,N_7,N_742);
or U1074 (N_1074,N_432,N_298);
and U1075 (N_1075,N_455,N_306);
nand U1076 (N_1076,N_417,N_257);
nor U1077 (N_1077,N_154,N_232);
or U1078 (N_1078,N_565,N_450);
and U1079 (N_1079,N_0,N_579);
nor U1080 (N_1080,N_551,N_294);
or U1081 (N_1081,N_561,N_362);
xnor U1082 (N_1082,N_105,N_596);
or U1083 (N_1083,N_702,N_189);
and U1084 (N_1084,N_63,N_141);
or U1085 (N_1085,N_260,N_320);
nor U1086 (N_1086,N_148,N_69);
nand U1087 (N_1087,N_433,N_516);
nand U1088 (N_1088,N_382,N_553);
nand U1089 (N_1089,N_345,N_498);
nor U1090 (N_1090,N_464,N_504);
xnor U1091 (N_1091,N_57,N_663);
nand U1092 (N_1092,N_341,N_19);
nor U1093 (N_1093,N_662,N_27);
or U1094 (N_1094,N_506,N_384);
nand U1095 (N_1095,N_240,N_38);
nor U1096 (N_1096,N_243,N_595);
and U1097 (N_1097,N_550,N_219);
or U1098 (N_1098,N_415,N_190);
and U1099 (N_1099,N_472,N_300);
and U1100 (N_1100,N_746,N_600);
and U1101 (N_1101,N_365,N_512);
nand U1102 (N_1102,N_8,N_185);
or U1103 (N_1103,N_156,N_626);
or U1104 (N_1104,N_681,N_416);
or U1105 (N_1105,N_49,N_114);
and U1106 (N_1106,N_741,N_167);
and U1107 (N_1107,N_522,N_197);
and U1108 (N_1108,N_674,N_404);
and U1109 (N_1109,N_258,N_204);
or U1110 (N_1110,N_152,N_130);
xor U1111 (N_1111,N_627,N_37);
nor U1112 (N_1112,N_32,N_474);
and U1113 (N_1113,N_598,N_264);
or U1114 (N_1114,N_738,N_578);
or U1115 (N_1115,N_712,N_303);
and U1116 (N_1116,N_430,N_334);
nor U1117 (N_1117,N_33,N_556);
nand U1118 (N_1118,N_248,N_423);
or U1119 (N_1119,N_572,N_534);
nand U1120 (N_1120,N_66,N_646);
and U1121 (N_1121,N_87,N_21);
and U1122 (N_1122,N_518,N_509);
nand U1123 (N_1123,N_484,N_83);
or U1124 (N_1124,N_466,N_690);
and U1125 (N_1125,N_600,N_47);
and U1126 (N_1126,N_347,N_737);
nor U1127 (N_1127,N_98,N_413);
and U1128 (N_1128,N_441,N_85);
nand U1129 (N_1129,N_586,N_223);
nor U1130 (N_1130,N_225,N_204);
or U1131 (N_1131,N_729,N_49);
or U1132 (N_1132,N_159,N_619);
nand U1133 (N_1133,N_340,N_682);
or U1134 (N_1134,N_57,N_315);
nand U1135 (N_1135,N_36,N_363);
nand U1136 (N_1136,N_277,N_692);
nand U1137 (N_1137,N_457,N_561);
nor U1138 (N_1138,N_12,N_446);
or U1139 (N_1139,N_678,N_15);
or U1140 (N_1140,N_295,N_729);
xnor U1141 (N_1141,N_499,N_572);
or U1142 (N_1142,N_444,N_636);
nand U1143 (N_1143,N_432,N_273);
nand U1144 (N_1144,N_305,N_221);
nor U1145 (N_1145,N_12,N_330);
nand U1146 (N_1146,N_158,N_393);
and U1147 (N_1147,N_705,N_743);
and U1148 (N_1148,N_77,N_595);
nor U1149 (N_1149,N_456,N_128);
nand U1150 (N_1150,N_338,N_566);
nor U1151 (N_1151,N_236,N_234);
or U1152 (N_1152,N_411,N_432);
or U1153 (N_1153,N_179,N_123);
and U1154 (N_1154,N_660,N_381);
or U1155 (N_1155,N_518,N_446);
and U1156 (N_1156,N_737,N_183);
or U1157 (N_1157,N_535,N_239);
and U1158 (N_1158,N_184,N_567);
nor U1159 (N_1159,N_172,N_106);
and U1160 (N_1160,N_344,N_262);
or U1161 (N_1161,N_111,N_266);
nand U1162 (N_1162,N_411,N_638);
and U1163 (N_1163,N_639,N_99);
nor U1164 (N_1164,N_37,N_41);
or U1165 (N_1165,N_604,N_295);
nor U1166 (N_1166,N_515,N_582);
and U1167 (N_1167,N_647,N_278);
or U1168 (N_1168,N_565,N_320);
or U1169 (N_1169,N_378,N_477);
and U1170 (N_1170,N_680,N_278);
or U1171 (N_1171,N_566,N_587);
nor U1172 (N_1172,N_432,N_481);
nor U1173 (N_1173,N_76,N_130);
and U1174 (N_1174,N_676,N_234);
or U1175 (N_1175,N_29,N_140);
nor U1176 (N_1176,N_562,N_224);
nor U1177 (N_1177,N_351,N_297);
nand U1178 (N_1178,N_280,N_690);
nor U1179 (N_1179,N_362,N_110);
xor U1180 (N_1180,N_264,N_612);
and U1181 (N_1181,N_321,N_579);
nand U1182 (N_1182,N_464,N_698);
nor U1183 (N_1183,N_612,N_405);
nand U1184 (N_1184,N_499,N_456);
or U1185 (N_1185,N_118,N_442);
and U1186 (N_1186,N_500,N_237);
or U1187 (N_1187,N_8,N_106);
nand U1188 (N_1188,N_246,N_38);
and U1189 (N_1189,N_679,N_349);
xnor U1190 (N_1190,N_125,N_20);
nor U1191 (N_1191,N_749,N_322);
nand U1192 (N_1192,N_737,N_198);
nand U1193 (N_1193,N_466,N_10);
and U1194 (N_1194,N_276,N_392);
nor U1195 (N_1195,N_721,N_93);
or U1196 (N_1196,N_711,N_477);
and U1197 (N_1197,N_288,N_408);
nor U1198 (N_1198,N_660,N_225);
and U1199 (N_1199,N_529,N_195);
nand U1200 (N_1200,N_1,N_248);
nand U1201 (N_1201,N_707,N_690);
nand U1202 (N_1202,N_566,N_663);
or U1203 (N_1203,N_6,N_491);
nand U1204 (N_1204,N_517,N_17);
and U1205 (N_1205,N_373,N_102);
and U1206 (N_1206,N_469,N_339);
or U1207 (N_1207,N_370,N_589);
and U1208 (N_1208,N_60,N_160);
nand U1209 (N_1209,N_157,N_276);
nand U1210 (N_1210,N_248,N_546);
nand U1211 (N_1211,N_425,N_67);
or U1212 (N_1212,N_636,N_589);
nor U1213 (N_1213,N_478,N_94);
nand U1214 (N_1214,N_147,N_485);
and U1215 (N_1215,N_339,N_15);
nand U1216 (N_1216,N_54,N_84);
nand U1217 (N_1217,N_729,N_292);
or U1218 (N_1218,N_601,N_47);
nand U1219 (N_1219,N_53,N_224);
or U1220 (N_1220,N_280,N_16);
xnor U1221 (N_1221,N_22,N_371);
and U1222 (N_1222,N_89,N_513);
and U1223 (N_1223,N_629,N_452);
nor U1224 (N_1224,N_65,N_163);
nor U1225 (N_1225,N_409,N_743);
or U1226 (N_1226,N_701,N_517);
nor U1227 (N_1227,N_74,N_676);
and U1228 (N_1228,N_423,N_117);
or U1229 (N_1229,N_406,N_259);
and U1230 (N_1230,N_693,N_739);
and U1231 (N_1231,N_280,N_243);
nor U1232 (N_1232,N_661,N_277);
or U1233 (N_1233,N_680,N_319);
and U1234 (N_1234,N_240,N_326);
nor U1235 (N_1235,N_384,N_181);
nor U1236 (N_1236,N_748,N_428);
nand U1237 (N_1237,N_361,N_133);
nand U1238 (N_1238,N_356,N_578);
nor U1239 (N_1239,N_126,N_728);
nor U1240 (N_1240,N_631,N_568);
or U1241 (N_1241,N_345,N_338);
nand U1242 (N_1242,N_44,N_649);
or U1243 (N_1243,N_356,N_482);
and U1244 (N_1244,N_53,N_555);
nand U1245 (N_1245,N_510,N_325);
and U1246 (N_1246,N_744,N_76);
nand U1247 (N_1247,N_683,N_305);
or U1248 (N_1248,N_667,N_105);
or U1249 (N_1249,N_501,N_362);
or U1250 (N_1250,N_610,N_30);
nand U1251 (N_1251,N_482,N_495);
and U1252 (N_1252,N_620,N_533);
or U1253 (N_1253,N_345,N_649);
and U1254 (N_1254,N_408,N_659);
nor U1255 (N_1255,N_348,N_645);
nor U1256 (N_1256,N_225,N_600);
or U1257 (N_1257,N_246,N_115);
and U1258 (N_1258,N_571,N_17);
or U1259 (N_1259,N_186,N_30);
nor U1260 (N_1260,N_470,N_97);
nor U1261 (N_1261,N_152,N_308);
and U1262 (N_1262,N_676,N_726);
or U1263 (N_1263,N_372,N_360);
and U1264 (N_1264,N_507,N_398);
nor U1265 (N_1265,N_602,N_107);
and U1266 (N_1266,N_617,N_137);
nor U1267 (N_1267,N_118,N_666);
or U1268 (N_1268,N_689,N_725);
nor U1269 (N_1269,N_503,N_368);
or U1270 (N_1270,N_648,N_480);
or U1271 (N_1271,N_618,N_334);
nor U1272 (N_1272,N_272,N_322);
and U1273 (N_1273,N_105,N_102);
nor U1274 (N_1274,N_615,N_573);
nor U1275 (N_1275,N_565,N_41);
or U1276 (N_1276,N_727,N_284);
or U1277 (N_1277,N_111,N_395);
or U1278 (N_1278,N_552,N_606);
or U1279 (N_1279,N_112,N_110);
and U1280 (N_1280,N_401,N_239);
or U1281 (N_1281,N_174,N_730);
or U1282 (N_1282,N_431,N_722);
nand U1283 (N_1283,N_672,N_182);
or U1284 (N_1284,N_182,N_490);
nor U1285 (N_1285,N_168,N_474);
or U1286 (N_1286,N_227,N_625);
nor U1287 (N_1287,N_686,N_65);
or U1288 (N_1288,N_192,N_286);
xnor U1289 (N_1289,N_126,N_110);
and U1290 (N_1290,N_357,N_564);
and U1291 (N_1291,N_669,N_587);
nor U1292 (N_1292,N_119,N_539);
nand U1293 (N_1293,N_177,N_361);
xor U1294 (N_1294,N_745,N_146);
or U1295 (N_1295,N_347,N_428);
or U1296 (N_1296,N_397,N_209);
nand U1297 (N_1297,N_270,N_724);
nor U1298 (N_1298,N_99,N_349);
nand U1299 (N_1299,N_314,N_668);
and U1300 (N_1300,N_516,N_645);
or U1301 (N_1301,N_18,N_189);
nor U1302 (N_1302,N_307,N_573);
and U1303 (N_1303,N_167,N_437);
nand U1304 (N_1304,N_712,N_741);
or U1305 (N_1305,N_729,N_427);
or U1306 (N_1306,N_515,N_414);
nand U1307 (N_1307,N_108,N_21);
and U1308 (N_1308,N_54,N_461);
or U1309 (N_1309,N_674,N_257);
nand U1310 (N_1310,N_736,N_297);
and U1311 (N_1311,N_152,N_531);
or U1312 (N_1312,N_573,N_416);
nand U1313 (N_1313,N_177,N_196);
xnor U1314 (N_1314,N_240,N_557);
nand U1315 (N_1315,N_624,N_201);
and U1316 (N_1316,N_743,N_297);
or U1317 (N_1317,N_372,N_565);
nor U1318 (N_1318,N_620,N_490);
or U1319 (N_1319,N_727,N_334);
and U1320 (N_1320,N_711,N_126);
xnor U1321 (N_1321,N_575,N_344);
and U1322 (N_1322,N_670,N_250);
and U1323 (N_1323,N_455,N_738);
nand U1324 (N_1324,N_746,N_473);
and U1325 (N_1325,N_660,N_309);
or U1326 (N_1326,N_505,N_63);
and U1327 (N_1327,N_416,N_448);
nor U1328 (N_1328,N_220,N_421);
nor U1329 (N_1329,N_306,N_397);
nand U1330 (N_1330,N_644,N_480);
xnor U1331 (N_1331,N_659,N_553);
nor U1332 (N_1332,N_261,N_747);
or U1333 (N_1333,N_486,N_629);
nor U1334 (N_1334,N_82,N_232);
or U1335 (N_1335,N_46,N_665);
and U1336 (N_1336,N_295,N_155);
xor U1337 (N_1337,N_375,N_606);
nor U1338 (N_1338,N_20,N_489);
or U1339 (N_1339,N_575,N_567);
nor U1340 (N_1340,N_591,N_686);
nand U1341 (N_1341,N_111,N_620);
nand U1342 (N_1342,N_735,N_26);
or U1343 (N_1343,N_308,N_672);
and U1344 (N_1344,N_330,N_260);
and U1345 (N_1345,N_371,N_315);
nand U1346 (N_1346,N_610,N_79);
or U1347 (N_1347,N_536,N_36);
nand U1348 (N_1348,N_354,N_307);
and U1349 (N_1349,N_582,N_714);
nor U1350 (N_1350,N_617,N_361);
or U1351 (N_1351,N_640,N_542);
and U1352 (N_1352,N_54,N_188);
or U1353 (N_1353,N_607,N_626);
nand U1354 (N_1354,N_178,N_400);
nor U1355 (N_1355,N_28,N_368);
nor U1356 (N_1356,N_714,N_367);
or U1357 (N_1357,N_303,N_101);
nand U1358 (N_1358,N_174,N_184);
nor U1359 (N_1359,N_673,N_404);
nor U1360 (N_1360,N_314,N_366);
nand U1361 (N_1361,N_68,N_350);
nor U1362 (N_1362,N_725,N_428);
or U1363 (N_1363,N_551,N_139);
and U1364 (N_1364,N_132,N_200);
or U1365 (N_1365,N_638,N_257);
nor U1366 (N_1366,N_715,N_381);
nor U1367 (N_1367,N_310,N_209);
nor U1368 (N_1368,N_625,N_86);
nand U1369 (N_1369,N_741,N_354);
nand U1370 (N_1370,N_458,N_101);
nor U1371 (N_1371,N_108,N_623);
and U1372 (N_1372,N_234,N_57);
nor U1373 (N_1373,N_319,N_197);
or U1374 (N_1374,N_515,N_503);
or U1375 (N_1375,N_72,N_158);
and U1376 (N_1376,N_319,N_728);
and U1377 (N_1377,N_706,N_476);
nand U1378 (N_1378,N_484,N_262);
nand U1379 (N_1379,N_478,N_250);
nand U1380 (N_1380,N_594,N_453);
or U1381 (N_1381,N_279,N_742);
nand U1382 (N_1382,N_96,N_105);
nor U1383 (N_1383,N_183,N_166);
and U1384 (N_1384,N_709,N_224);
xnor U1385 (N_1385,N_408,N_511);
nand U1386 (N_1386,N_385,N_229);
and U1387 (N_1387,N_575,N_83);
or U1388 (N_1388,N_223,N_667);
nor U1389 (N_1389,N_372,N_668);
or U1390 (N_1390,N_211,N_573);
nor U1391 (N_1391,N_528,N_566);
or U1392 (N_1392,N_733,N_702);
nand U1393 (N_1393,N_624,N_311);
and U1394 (N_1394,N_553,N_336);
and U1395 (N_1395,N_692,N_737);
nand U1396 (N_1396,N_510,N_265);
and U1397 (N_1397,N_476,N_150);
and U1398 (N_1398,N_514,N_667);
and U1399 (N_1399,N_457,N_190);
or U1400 (N_1400,N_748,N_27);
nand U1401 (N_1401,N_364,N_202);
nand U1402 (N_1402,N_108,N_229);
nand U1403 (N_1403,N_310,N_683);
and U1404 (N_1404,N_388,N_520);
and U1405 (N_1405,N_725,N_377);
and U1406 (N_1406,N_659,N_669);
or U1407 (N_1407,N_433,N_281);
and U1408 (N_1408,N_496,N_319);
and U1409 (N_1409,N_354,N_729);
nand U1410 (N_1410,N_130,N_644);
nor U1411 (N_1411,N_568,N_43);
and U1412 (N_1412,N_346,N_470);
or U1413 (N_1413,N_730,N_665);
nor U1414 (N_1414,N_11,N_467);
nor U1415 (N_1415,N_427,N_619);
or U1416 (N_1416,N_183,N_614);
and U1417 (N_1417,N_391,N_177);
xnor U1418 (N_1418,N_324,N_39);
nor U1419 (N_1419,N_256,N_185);
and U1420 (N_1420,N_629,N_493);
and U1421 (N_1421,N_138,N_450);
nor U1422 (N_1422,N_405,N_87);
nor U1423 (N_1423,N_109,N_677);
nand U1424 (N_1424,N_39,N_144);
or U1425 (N_1425,N_626,N_436);
and U1426 (N_1426,N_647,N_90);
or U1427 (N_1427,N_88,N_89);
nand U1428 (N_1428,N_554,N_427);
nand U1429 (N_1429,N_245,N_640);
and U1430 (N_1430,N_42,N_282);
nand U1431 (N_1431,N_29,N_426);
nor U1432 (N_1432,N_577,N_643);
nand U1433 (N_1433,N_592,N_265);
and U1434 (N_1434,N_486,N_408);
nand U1435 (N_1435,N_37,N_608);
or U1436 (N_1436,N_236,N_274);
nor U1437 (N_1437,N_178,N_356);
nor U1438 (N_1438,N_310,N_383);
or U1439 (N_1439,N_625,N_286);
and U1440 (N_1440,N_476,N_641);
and U1441 (N_1441,N_396,N_427);
or U1442 (N_1442,N_248,N_313);
and U1443 (N_1443,N_746,N_432);
or U1444 (N_1444,N_194,N_610);
nor U1445 (N_1445,N_258,N_588);
nor U1446 (N_1446,N_3,N_411);
nor U1447 (N_1447,N_597,N_592);
nor U1448 (N_1448,N_96,N_741);
nand U1449 (N_1449,N_407,N_382);
or U1450 (N_1450,N_329,N_296);
nor U1451 (N_1451,N_67,N_378);
nand U1452 (N_1452,N_493,N_62);
nand U1453 (N_1453,N_576,N_729);
nor U1454 (N_1454,N_573,N_103);
or U1455 (N_1455,N_499,N_718);
or U1456 (N_1456,N_359,N_566);
or U1457 (N_1457,N_656,N_352);
and U1458 (N_1458,N_150,N_388);
and U1459 (N_1459,N_738,N_240);
or U1460 (N_1460,N_18,N_442);
and U1461 (N_1461,N_663,N_71);
and U1462 (N_1462,N_655,N_138);
or U1463 (N_1463,N_400,N_154);
nand U1464 (N_1464,N_276,N_23);
and U1465 (N_1465,N_290,N_269);
nor U1466 (N_1466,N_571,N_523);
or U1467 (N_1467,N_523,N_491);
nor U1468 (N_1468,N_716,N_739);
nand U1469 (N_1469,N_735,N_210);
nand U1470 (N_1470,N_705,N_123);
or U1471 (N_1471,N_505,N_396);
nand U1472 (N_1472,N_152,N_551);
nor U1473 (N_1473,N_296,N_316);
or U1474 (N_1474,N_747,N_674);
and U1475 (N_1475,N_517,N_5);
nor U1476 (N_1476,N_648,N_82);
nor U1477 (N_1477,N_535,N_445);
and U1478 (N_1478,N_114,N_348);
and U1479 (N_1479,N_97,N_528);
nand U1480 (N_1480,N_726,N_728);
nor U1481 (N_1481,N_82,N_247);
or U1482 (N_1482,N_254,N_460);
nand U1483 (N_1483,N_243,N_582);
nor U1484 (N_1484,N_15,N_194);
or U1485 (N_1485,N_152,N_106);
or U1486 (N_1486,N_101,N_497);
nor U1487 (N_1487,N_297,N_42);
nand U1488 (N_1488,N_702,N_524);
and U1489 (N_1489,N_8,N_635);
and U1490 (N_1490,N_209,N_360);
or U1491 (N_1491,N_437,N_643);
and U1492 (N_1492,N_546,N_711);
and U1493 (N_1493,N_146,N_67);
and U1494 (N_1494,N_584,N_354);
and U1495 (N_1495,N_367,N_202);
nand U1496 (N_1496,N_274,N_446);
nand U1497 (N_1497,N_672,N_625);
nand U1498 (N_1498,N_60,N_420);
or U1499 (N_1499,N_710,N_267);
or U1500 (N_1500,N_1051,N_1010);
or U1501 (N_1501,N_1323,N_821);
nor U1502 (N_1502,N_1150,N_1303);
nor U1503 (N_1503,N_908,N_1141);
nand U1504 (N_1504,N_1153,N_961);
or U1505 (N_1505,N_792,N_1173);
or U1506 (N_1506,N_1252,N_1412);
and U1507 (N_1507,N_1274,N_926);
and U1508 (N_1508,N_1498,N_1122);
nand U1509 (N_1509,N_1129,N_1368);
and U1510 (N_1510,N_857,N_1395);
nor U1511 (N_1511,N_822,N_1367);
or U1512 (N_1512,N_1224,N_1215);
or U1513 (N_1513,N_1040,N_1206);
or U1514 (N_1514,N_1433,N_1483);
or U1515 (N_1515,N_1091,N_1270);
nor U1516 (N_1516,N_900,N_1309);
and U1517 (N_1517,N_913,N_818);
nor U1518 (N_1518,N_1330,N_906);
xor U1519 (N_1519,N_996,N_1351);
and U1520 (N_1520,N_1316,N_1012);
nor U1521 (N_1521,N_804,N_1358);
nand U1522 (N_1522,N_896,N_1280);
nand U1523 (N_1523,N_1095,N_1382);
and U1524 (N_1524,N_915,N_1161);
and U1525 (N_1525,N_1499,N_1468);
or U1526 (N_1526,N_1260,N_1408);
xnor U1527 (N_1527,N_1272,N_838);
nor U1528 (N_1528,N_1453,N_979);
nor U1529 (N_1529,N_1105,N_1221);
nor U1530 (N_1530,N_995,N_1465);
nor U1531 (N_1531,N_1101,N_912);
and U1532 (N_1532,N_847,N_1213);
nor U1533 (N_1533,N_1211,N_1423);
nand U1534 (N_1534,N_1463,N_1293);
and U1535 (N_1535,N_1230,N_820);
or U1536 (N_1536,N_993,N_810);
nand U1537 (N_1537,N_1262,N_795);
nand U1538 (N_1538,N_1456,N_1186);
and U1539 (N_1539,N_1044,N_1132);
and U1540 (N_1540,N_1345,N_1170);
nor U1541 (N_1541,N_1033,N_1043);
or U1542 (N_1542,N_1369,N_895);
nand U1543 (N_1543,N_1302,N_1046);
or U1544 (N_1544,N_919,N_808);
nor U1545 (N_1545,N_1076,N_962);
nand U1546 (N_1546,N_1363,N_1111);
and U1547 (N_1547,N_813,N_902);
nand U1548 (N_1548,N_1269,N_885);
or U1549 (N_1549,N_1344,N_1488);
and U1550 (N_1550,N_863,N_1026);
nand U1551 (N_1551,N_1246,N_866);
and U1552 (N_1552,N_957,N_973);
or U1553 (N_1553,N_1059,N_1304);
nand U1554 (N_1554,N_983,N_1264);
or U1555 (N_1555,N_1257,N_837);
nor U1556 (N_1556,N_1282,N_1157);
or U1557 (N_1557,N_1128,N_1159);
and U1558 (N_1558,N_940,N_1065);
nand U1559 (N_1559,N_811,N_879);
nor U1560 (N_1560,N_765,N_805);
nand U1561 (N_1561,N_1370,N_1396);
and U1562 (N_1562,N_977,N_951);
nor U1563 (N_1563,N_1287,N_815);
or U1564 (N_1564,N_1312,N_1455);
nor U1565 (N_1565,N_1016,N_1376);
nand U1566 (N_1566,N_1255,N_1341);
nor U1567 (N_1567,N_803,N_964);
and U1568 (N_1568,N_1256,N_819);
and U1569 (N_1569,N_781,N_1176);
nand U1570 (N_1570,N_841,N_1019);
or U1571 (N_1571,N_1163,N_757);
and U1572 (N_1572,N_1139,N_901);
nand U1573 (N_1573,N_762,N_1054);
and U1574 (N_1574,N_985,N_776);
nor U1575 (N_1575,N_1003,N_1485);
or U1576 (N_1576,N_1056,N_889);
nor U1577 (N_1577,N_1311,N_1088);
or U1578 (N_1578,N_1049,N_1409);
nor U1579 (N_1579,N_884,N_1015);
nor U1580 (N_1580,N_1177,N_1249);
nand U1581 (N_1581,N_1036,N_1497);
nand U1582 (N_1582,N_959,N_1169);
or U1583 (N_1583,N_1373,N_796);
and U1584 (N_1584,N_945,N_1387);
or U1585 (N_1585,N_759,N_1023);
and U1586 (N_1586,N_1340,N_1209);
or U1587 (N_1587,N_969,N_924);
and U1588 (N_1588,N_1191,N_1394);
and U1589 (N_1589,N_784,N_1310);
and U1590 (N_1590,N_1307,N_1421);
or U1591 (N_1591,N_1354,N_873);
nor U1592 (N_1592,N_914,N_988);
nand U1593 (N_1593,N_1067,N_1145);
nor U1594 (N_1594,N_1188,N_756);
and U1595 (N_1595,N_1377,N_845);
or U1596 (N_1596,N_953,N_785);
and U1597 (N_1597,N_1298,N_862);
and U1598 (N_1598,N_1251,N_1212);
or U1599 (N_1599,N_999,N_1415);
nand U1600 (N_1600,N_1239,N_856);
and U1601 (N_1601,N_1119,N_1347);
and U1602 (N_1602,N_1063,N_771);
nor U1603 (N_1603,N_773,N_1184);
nor U1604 (N_1604,N_1237,N_806);
nor U1605 (N_1605,N_893,N_1000);
and U1606 (N_1606,N_1460,N_1399);
or U1607 (N_1607,N_1028,N_892);
and U1608 (N_1608,N_839,N_1151);
nor U1609 (N_1609,N_1052,N_1108);
nand U1610 (N_1610,N_774,N_894);
nand U1611 (N_1611,N_1178,N_768);
and U1612 (N_1612,N_1086,N_935);
nor U1613 (N_1613,N_1438,N_831);
nor U1614 (N_1614,N_1154,N_760);
or U1615 (N_1615,N_984,N_1374);
nor U1616 (N_1616,N_782,N_1353);
or U1617 (N_1617,N_903,N_1467);
xnor U1618 (N_1618,N_761,N_834);
nand U1619 (N_1619,N_750,N_1275);
or U1620 (N_1620,N_1201,N_1031);
nand U1621 (N_1621,N_1072,N_1068);
and U1622 (N_1622,N_958,N_1286);
and U1623 (N_1623,N_1001,N_764);
and U1624 (N_1624,N_1331,N_974);
and U1625 (N_1625,N_1431,N_770);
or U1626 (N_1626,N_1440,N_1087);
and U1627 (N_1627,N_1407,N_963);
nor U1628 (N_1628,N_1041,N_1048);
nand U1629 (N_1629,N_987,N_1271);
nand U1630 (N_1630,N_1155,N_1491);
nor U1631 (N_1631,N_1143,N_1427);
or U1632 (N_1632,N_1231,N_1118);
or U1633 (N_1633,N_1457,N_992);
nand U1634 (N_1634,N_954,N_767);
nand U1635 (N_1635,N_825,N_1179);
or U1636 (N_1636,N_1100,N_1338);
nand U1637 (N_1637,N_1138,N_1165);
or U1638 (N_1638,N_1225,N_991);
and U1639 (N_1639,N_1417,N_1327);
nand U1640 (N_1640,N_1147,N_1444);
or U1641 (N_1641,N_1320,N_1339);
and U1642 (N_1642,N_1492,N_1240);
or U1643 (N_1643,N_1452,N_1058);
nor U1644 (N_1644,N_1093,N_1069);
nor U1645 (N_1645,N_1416,N_876);
nor U1646 (N_1646,N_1294,N_1217);
or U1647 (N_1647,N_1337,N_971);
nor U1648 (N_1648,N_1356,N_1117);
nand U1649 (N_1649,N_1414,N_1136);
nand U1650 (N_1650,N_1484,N_1328);
nor U1651 (N_1651,N_1386,N_1162);
or U1652 (N_1652,N_981,N_994);
and U1653 (N_1653,N_828,N_1144);
nand U1654 (N_1654,N_1166,N_791);
or U1655 (N_1655,N_1437,N_1247);
and U1656 (N_1656,N_842,N_1442);
or U1657 (N_1657,N_829,N_1352);
nand U1658 (N_1658,N_1443,N_1349);
and U1659 (N_1659,N_1360,N_1329);
or U1660 (N_1660,N_1253,N_1197);
or U1661 (N_1661,N_1299,N_1203);
and U1662 (N_1662,N_869,N_1266);
and U1663 (N_1663,N_1355,N_800);
nor U1664 (N_1664,N_1060,N_1089);
or U1665 (N_1665,N_1276,N_1406);
nand U1666 (N_1666,N_1171,N_1222);
or U1667 (N_1667,N_1400,N_1482);
nand U1668 (N_1668,N_1158,N_970);
nor U1669 (N_1669,N_1167,N_1032);
nor U1670 (N_1670,N_1300,N_1318);
nor U1671 (N_1671,N_1097,N_1478);
and U1672 (N_1672,N_824,N_1005);
nand U1673 (N_1673,N_783,N_1306);
or U1674 (N_1674,N_1446,N_943);
nand U1675 (N_1675,N_1148,N_823);
and U1676 (N_1676,N_1180,N_1495);
nand U1677 (N_1677,N_1198,N_1259);
and U1678 (N_1678,N_1137,N_1200);
nand U1679 (N_1679,N_1418,N_872);
nand U1680 (N_1680,N_1359,N_905);
nor U1681 (N_1681,N_890,N_1420);
or U1682 (N_1682,N_1055,N_1050);
nand U1683 (N_1683,N_1234,N_852);
nor U1684 (N_1684,N_1034,N_934);
and U1685 (N_1685,N_1194,N_1116);
and U1686 (N_1686,N_755,N_1134);
nor U1687 (N_1687,N_1018,N_1017);
nand U1688 (N_1688,N_975,N_1383);
and U1689 (N_1689,N_1125,N_966);
nand U1690 (N_1690,N_1461,N_809);
nand U1691 (N_1691,N_1024,N_1219);
or U1692 (N_1692,N_944,N_1472);
or U1693 (N_1693,N_965,N_1216);
nor U1694 (N_1694,N_1388,N_1285);
nand U1695 (N_1695,N_922,N_1490);
nand U1696 (N_1696,N_882,N_1451);
and U1697 (N_1697,N_799,N_932);
nor U1698 (N_1698,N_763,N_1441);
nand U1699 (N_1699,N_1475,N_836);
nor U1700 (N_1700,N_833,N_1474);
nor U1701 (N_1701,N_1283,N_1301);
or U1702 (N_1702,N_967,N_1466);
nor U1703 (N_1703,N_947,N_858);
nor U1704 (N_1704,N_867,N_1250);
or U1705 (N_1705,N_1322,N_1333);
and U1706 (N_1706,N_1486,N_887);
and U1707 (N_1707,N_1228,N_775);
nor U1708 (N_1708,N_1030,N_1099);
or U1709 (N_1709,N_1413,N_752);
and U1710 (N_1710,N_946,N_1082);
nand U1711 (N_1711,N_1366,N_1432);
or U1712 (N_1712,N_1077,N_1389);
nor U1713 (N_1713,N_1494,N_1190);
nand U1714 (N_1714,N_798,N_1362);
and U1715 (N_1715,N_1061,N_1090);
or U1716 (N_1716,N_1185,N_1254);
and U1717 (N_1717,N_1102,N_978);
nor U1718 (N_1718,N_1326,N_877);
nor U1719 (N_1719,N_1064,N_769);
nor U1720 (N_1720,N_1290,N_917);
nor U1721 (N_1721,N_1021,N_1182);
nand U1722 (N_1722,N_998,N_1480);
or U1723 (N_1723,N_1405,N_1014);
nand U1724 (N_1724,N_1196,N_1039);
nor U1725 (N_1725,N_1164,N_1092);
nor U1726 (N_1726,N_898,N_1245);
or U1727 (N_1727,N_923,N_787);
nor U1728 (N_1728,N_1175,N_1258);
or U1729 (N_1729,N_916,N_1081);
nor U1730 (N_1730,N_1317,N_1291);
and U1731 (N_1731,N_1464,N_1172);
and U1732 (N_1732,N_1229,N_840);
nor U1733 (N_1733,N_1160,N_1103);
and U1734 (N_1734,N_1430,N_1454);
nand U1735 (N_1735,N_1398,N_1227);
or U1736 (N_1736,N_1130,N_1447);
and U1737 (N_1737,N_1127,N_1140);
xnor U1738 (N_1738,N_1419,N_989);
nor U1739 (N_1739,N_1448,N_1357);
and U1740 (N_1740,N_1226,N_950);
xnor U1741 (N_1741,N_972,N_832);
nor U1742 (N_1742,N_1223,N_1078);
nand U1743 (N_1743,N_1288,N_910);
nand U1744 (N_1744,N_1426,N_1403);
nand U1745 (N_1745,N_1434,N_1098);
nand U1746 (N_1746,N_1114,N_1445);
nor U1747 (N_1747,N_1477,N_1348);
nand U1748 (N_1748,N_968,N_1042);
or U1749 (N_1749,N_1273,N_864);
and U1750 (N_1750,N_1401,N_790);
xor U1751 (N_1751,N_955,N_1375);
nand U1752 (N_1752,N_1496,N_1284);
and U1753 (N_1753,N_1361,N_1193);
nand U1754 (N_1754,N_874,N_888);
and U1755 (N_1755,N_982,N_865);
and U1756 (N_1756,N_1047,N_1189);
or U1757 (N_1757,N_1402,N_830);
nand U1758 (N_1758,N_1422,N_844);
nor U1759 (N_1759,N_1070,N_1183);
and U1760 (N_1760,N_1279,N_1008);
or U1761 (N_1761,N_1261,N_1404);
and U1762 (N_1762,N_939,N_1006);
or U1763 (N_1763,N_849,N_1305);
and U1764 (N_1764,N_1109,N_1391);
nor U1765 (N_1765,N_1289,N_930);
or U1766 (N_1766,N_1192,N_1385);
nor U1767 (N_1767,N_911,N_1232);
nor U1768 (N_1768,N_758,N_1007);
nand U1769 (N_1769,N_1263,N_925);
nand U1770 (N_1770,N_929,N_1481);
and U1771 (N_1771,N_937,N_1071);
or U1772 (N_1772,N_1278,N_1002);
nand U1773 (N_1773,N_952,N_1029);
nand U1774 (N_1774,N_1314,N_1424);
and U1775 (N_1775,N_868,N_1364);
and U1776 (N_1776,N_1104,N_1429);
nand U1777 (N_1777,N_1152,N_1009);
nand U1778 (N_1778,N_1233,N_788);
and U1779 (N_1779,N_851,N_1381);
and U1780 (N_1780,N_1149,N_1195);
and U1781 (N_1781,N_1350,N_843);
or U1782 (N_1782,N_1242,N_1207);
or U1783 (N_1783,N_1321,N_1281);
nor U1784 (N_1784,N_1471,N_1074);
nand U1785 (N_1785,N_980,N_1380);
nand U1786 (N_1786,N_1392,N_986);
nor U1787 (N_1787,N_938,N_1297);
and U1788 (N_1788,N_1410,N_1121);
or U1789 (N_1789,N_1210,N_854);
nor U1790 (N_1790,N_1313,N_904);
and U1791 (N_1791,N_1378,N_1390);
and U1792 (N_1792,N_835,N_1372);
or U1793 (N_1793,N_1126,N_1238);
and U1794 (N_1794,N_766,N_1073);
nand U1795 (N_1795,N_1181,N_1135);
or U1796 (N_1796,N_1013,N_1045);
or U1797 (N_1797,N_1123,N_1037);
and U1798 (N_1798,N_1458,N_1397);
nand U1799 (N_1799,N_1493,N_1336);
or U1800 (N_1800,N_1342,N_1425);
or U1801 (N_1801,N_1295,N_909);
and U1802 (N_1802,N_1393,N_1057);
and U1803 (N_1803,N_1462,N_1124);
and U1804 (N_1804,N_918,N_990);
nand U1805 (N_1805,N_949,N_751);
nand U1806 (N_1806,N_1113,N_1084);
or U1807 (N_1807,N_1343,N_880);
and U1808 (N_1808,N_1053,N_1473);
xor U1809 (N_1809,N_1241,N_1435);
and U1810 (N_1810,N_1371,N_794);
and U1811 (N_1811,N_1107,N_1202);
or U1812 (N_1812,N_1079,N_1428);
or U1813 (N_1813,N_1244,N_960);
nand U1814 (N_1814,N_921,N_1075);
or U1815 (N_1815,N_1449,N_997);
or U1816 (N_1816,N_1131,N_772);
nand U1817 (N_1817,N_860,N_1265);
and U1818 (N_1818,N_859,N_1268);
or U1819 (N_1819,N_976,N_1292);
nor U1820 (N_1820,N_1476,N_1110);
and U1821 (N_1821,N_1267,N_1236);
or U1822 (N_1822,N_933,N_753);
nand U1823 (N_1823,N_870,N_1004);
nand U1824 (N_1824,N_861,N_812);
nor U1825 (N_1825,N_1450,N_801);
nor U1826 (N_1826,N_1133,N_814);
or U1827 (N_1827,N_1096,N_1411);
xor U1828 (N_1828,N_1022,N_1035);
nand U1829 (N_1829,N_920,N_1296);
or U1830 (N_1830,N_853,N_1027);
nand U1831 (N_1831,N_1335,N_1325);
nor U1832 (N_1832,N_1020,N_797);
xnor U1833 (N_1833,N_1248,N_1487);
nand U1834 (N_1834,N_883,N_928);
or U1835 (N_1835,N_942,N_1112);
and U1836 (N_1836,N_907,N_1332);
and U1837 (N_1837,N_1365,N_1174);
nor U1838 (N_1838,N_897,N_1106);
or U1839 (N_1839,N_802,N_827);
or U1840 (N_1840,N_1120,N_1436);
and U1841 (N_1841,N_891,N_1235);
nand U1842 (N_1842,N_1146,N_1489);
nor U1843 (N_1843,N_875,N_1346);
or U1844 (N_1844,N_1439,N_878);
or U1845 (N_1845,N_1156,N_817);
nor U1846 (N_1846,N_1115,N_1479);
nor U1847 (N_1847,N_1324,N_931);
nor U1848 (N_1848,N_881,N_1205);
or U1849 (N_1849,N_871,N_789);
nand U1850 (N_1850,N_1208,N_1199);
and U1851 (N_1851,N_1220,N_1469);
nor U1852 (N_1852,N_1459,N_1470);
nor U1853 (N_1853,N_1066,N_786);
or U1854 (N_1854,N_826,N_777);
or U1855 (N_1855,N_936,N_780);
nor U1856 (N_1856,N_1011,N_1080);
or U1857 (N_1857,N_1384,N_779);
or U1858 (N_1858,N_1214,N_816);
or U1859 (N_1859,N_1062,N_1025);
nand U1860 (N_1860,N_1187,N_1038);
or U1861 (N_1861,N_899,N_1142);
and U1862 (N_1862,N_1334,N_855);
nor U1863 (N_1863,N_1218,N_754);
nand U1864 (N_1864,N_1083,N_1308);
or U1865 (N_1865,N_948,N_793);
nand U1866 (N_1866,N_1379,N_1315);
or U1867 (N_1867,N_1277,N_1243);
nor U1868 (N_1868,N_927,N_807);
nand U1869 (N_1869,N_941,N_1168);
and U1870 (N_1870,N_1085,N_846);
nor U1871 (N_1871,N_886,N_1319);
nor U1872 (N_1872,N_778,N_956);
nor U1873 (N_1873,N_848,N_1204);
or U1874 (N_1874,N_1094,N_850);
and U1875 (N_1875,N_1314,N_1176);
nand U1876 (N_1876,N_1334,N_1430);
or U1877 (N_1877,N_1253,N_769);
or U1878 (N_1878,N_1292,N_1314);
or U1879 (N_1879,N_1217,N_1145);
nand U1880 (N_1880,N_978,N_924);
nor U1881 (N_1881,N_964,N_1350);
and U1882 (N_1882,N_1158,N_984);
and U1883 (N_1883,N_850,N_1496);
nand U1884 (N_1884,N_1213,N_1120);
nor U1885 (N_1885,N_1371,N_770);
nor U1886 (N_1886,N_1402,N_1039);
and U1887 (N_1887,N_1025,N_1079);
nand U1888 (N_1888,N_1346,N_1073);
nor U1889 (N_1889,N_1399,N_1282);
nand U1890 (N_1890,N_1442,N_777);
or U1891 (N_1891,N_1410,N_1442);
nand U1892 (N_1892,N_760,N_1280);
or U1893 (N_1893,N_910,N_963);
or U1894 (N_1894,N_1414,N_761);
and U1895 (N_1895,N_1262,N_976);
nand U1896 (N_1896,N_1155,N_1224);
or U1897 (N_1897,N_823,N_1385);
nand U1898 (N_1898,N_1187,N_1277);
and U1899 (N_1899,N_1282,N_1309);
or U1900 (N_1900,N_1186,N_887);
or U1901 (N_1901,N_1125,N_1366);
and U1902 (N_1902,N_1366,N_1430);
nor U1903 (N_1903,N_1361,N_1024);
or U1904 (N_1904,N_1440,N_1105);
nand U1905 (N_1905,N_1438,N_1147);
nor U1906 (N_1906,N_1067,N_1129);
and U1907 (N_1907,N_1410,N_1030);
or U1908 (N_1908,N_812,N_1015);
nand U1909 (N_1909,N_1209,N_1178);
nand U1910 (N_1910,N_1083,N_1406);
and U1911 (N_1911,N_1230,N_1395);
xnor U1912 (N_1912,N_909,N_1471);
nand U1913 (N_1913,N_1212,N_1156);
or U1914 (N_1914,N_1059,N_1021);
and U1915 (N_1915,N_1340,N_902);
or U1916 (N_1916,N_762,N_1217);
nand U1917 (N_1917,N_936,N_1320);
and U1918 (N_1918,N_952,N_913);
nand U1919 (N_1919,N_907,N_981);
nor U1920 (N_1920,N_965,N_1280);
nor U1921 (N_1921,N_1226,N_1362);
nor U1922 (N_1922,N_1259,N_1173);
and U1923 (N_1923,N_1003,N_1388);
nand U1924 (N_1924,N_896,N_1233);
or U1925 (N_1925,N_1138,N_1223);
or U1926 (N_1926,N_807,N_1416);
nand U1927 (N_1927,N_1315,N_1096);
or U1928 (N_1928,N_1238,N_1476);
and U1929 (N_1929,N_1347,N_1441);
nand U1930 (N_1930,N_1073,N_929);
and U1931 (N_1931,N_1471,N_852);
or U1932 (N_1932,N_882,N_1329);
nand U1933 (N_1933,N_1237,N_1175);
or U1934 (N_1934,N_1211,N_1198);
nand U1935 (N_1935,N_1220,N_1155);
nor U1936 (N_1936,N_1103,N_1267);
nor U1937 (N_1937,N_1285,N_967);
or U1938 (N_1938,N_1224,N_965);
or U1939 (N_1939,N_1212,N_906);
and U1940 (N_1940,N_1364,N_754);
nor U1941 (N_1941,N_1127,N_949);
or U1942 (N_1942,N_806,N_931);
or U1943 (N_1943,N_752,N_1308);
or U1944 (N_1944,N_855,N_766);
and U1945 (N_1945,N_992,N_1101);
and U1946 (N_1946,N_795,N_924);
nand U1947 (N_1947,N_1294,N_1282);
or U1948 (N_1948,N_1015,N_1054);
xnor U1949 (N_1949,N_1095,N_883);
xor U1950 (N_1950,N_1251,N_1270);
or U1951 (N_1951,N_1157,N_1299);
or U1952 (N_1952,N_1208,N_1281);
nor U1953 (N_1953,N_849,N_1274);
nand U1954 (N_1954,N_1062,N_961);
and U1955 (N_1955,N_869,N_1074);
nor U1956 (N_1956,N_1172,N_1309);
and U1957 (N_1957,N_813,N_750);
nor U1958 (N_1958,N_903,N_1148);
nor U1959 (N_1959,N_1035,N_1173);
nand U1960 (N_1960,N_1136,N_1436);
nand U1961 (N_1961,N_1186,N_918);
or U1962 (N_1962,N_1363,N_1039);
nor U1963 (N_1963,N_992,N_1092);
and U1964 (N_1964,N_979,N_808);
nor U1965 (N_1965,N_1133,N_1241);
and U1966 (N_1966,N_1079,N_1414);
nor U1967 (N_1967,N_1282,N_1262);
and U1968 (N_1968,N_933,N_1248);
or U1969 (N_1969,N_898,N_1191);
nor U1970 (N_1970,N_1219,N_786);
or U1971 (N_1971,N_1327,N_818);
or U1972 (N_1972,N_1151,N_893);
and U1973 (N_1973,N_1460,N_1126);
nand U1974 (N_1974,N_1011,N_1004);
and U1975 (N_1975,N_1317,N_1000);
nand U1976 (N_1976,N_1409,N_1227);
and U1977 (N_1977,N_978,N_1393);
or U1978 (N_1978,N_1139,N_1294);
nor U1979 (N_1979,N_1273,N_1357);
nand U1980 (N_1980,N_982,N_872);
or U1981 (N_1981,N_796,N_1339);
or U1982 (N_1982,N_943,N_891);
and U1983 (N_1983,N_1210,N_1380);
and U1984 (N_1984,N_923,N_813);
and U1985 (N_1985,N_1094,N_866);
nand U1986 (N_1986,N_1472,N_1148);
and U1987 (N_1987,N_1120,N_909);
nand U1988 (N_1988,N_800,N_1012);
or U1989 (N_1989,N_1184,N_1233);
nand U1990 (N_1990,N_1018,N_1130);
nor U1991 (N_1991,N_1147,N_1468);
or U1992 (N_1992,N_1113,N_851);
nand U1993 (N_1993,N_954,N_985);
nand U1994 (N_1994,N_1357,N_1085);
or U1995 (N_1995,N_833,N_1243);
or U1996 (N_1996,N_851,N_1468);
nor U1997 (N_1997,N_1291,N_940);
nand U1998 (N_1998,N_920,N_943);
or U1999 (N_1999,N_938,N_1275);
nand U2000 (N_2000,N_1252,N_1494);
nor U2001 (N_2001,N_1321,N_1425);
and U2002 (N_2002,N_849,N_1405);
nand U2003 (N_2003,N_1324,N_876);
nor U2004 (N_2004,N_1036,N_1410);
nor U2005 (N_2005,N_860,N_1084);
nand U2006 (N_2006,N_786,N_831);
or U2007 (N_2007,N_1354,N_767);
nor U2008 (N_2008,N_1268,N_751);
nand U2009 (N_2009,N_1430,N_776);
or U2010 (N_2010,N_765,N_1041);
nand U2011 (N_2011,N_1057,N_1328);
nand U2012 (N_2012,N_1048,N_1052);
and U2013 (N_2013,N_1134,N_1499);
and U2014 (N_2014,N_1201,N_1130);
or U2015 (N_2015,N_999,N_772);
nor U2016 (N_2016,N_1468,N_860);
and U2017 (N_2017,N_990,N_794);
nor U2018 (N_2018,N_1393,N_823);
xor U2019 (N_2019,N_920,N_1477);
nand U2020 (N_2020,N_1125,N_1228);
nand U2021 (N_2021,N_1012,N_1330);
or U2022 (N_2022,N_1116,N_856);
xor U2023 (N_2023,N_832,N_1081);
and U2024 (N_2024,N_1460,N_1300);
nor U2025 (N_2025,N_1430,N_1453);
or U2026 (N_2026,N_1081,N_885);
and U2027 (N_2027,N_1183,N_761);
nor U2028 (N_2028,N_1039,N_787);
nand U2029 (N_2029,N_1320,N_1044);
and U2030 (N_2030,N_1287,N_1166);
nor U2031 (N_2031,N_1203,N_988);
nor U2032 (N_2032,N_1033,N_1256);
and U2033 (N_2033,N_958,N_1491);
or U2034 (N_2034,N_1376,N_805);
nor U2035 (N_2035,N_1010,N_828);
or U2036 (N_2036,N_828,N_1322);
or U2037 (N_2037,N_1294,N_1287);
nor U2038 (N_2038,N_881,N_958);
xnor U2039 (N_2039,N_1017,N_1039);
nor U2040 (N_2040,N_1018,N_1206);
nand U2041 (N_2041,N_994,N_841);
nor U2042 (N_2042,N_976,N_1276);
or U2043 (N_2043,N_1275,N_1497);
nor U2044 (N_2044,N_1117,N_1409);
and U2045 (N_2045,N_893,N_1225);
nor U2046 (N_2046,N_1187,N_1316);
nand U2047 (N_2047,N_912,N_1481);
and U2048 (N_2048,N_1381,N_1458);
or U2049 (N_2049,N_801,N_1460);
nand U2050 (N_2050,N_768,N_780);
or U2051 (N_2051,N_1196,N_963);
or U2052 (N_2052,N_1288,N_972);
and U2053 (N_2053,N_1259,N_773);
nand U2054 (N_2054,N_1458,N_1385);
or U2055 (N_2055,N_1446,N_1044);
nor U2056 (N_2056,N_768,N_1063);
nand U2057 (N_2057,N_1050,N_1062);
or U2058 (N_2058,N_978,N_849);
and U2059 (N_2059,N_1044,N_756);
and U2060 (N_2060,N_1242,N_930);
nor U2061 (N_2061,N_835,N_764);
nor U2062 (N_2062,N_1021,N_1017);
nor U2063 (N_2063,N_1395,N_752);
and U2064 (N_2064,N_1392,N_1170);
or U2065 (N_2065,N_1223,N_1095);
and U2066 (N_2066,N_1022,N_1342);
nand U2067 (N_2067,N_963,N_1314);
or U2068 (N_2068,N_1318,N_1075);
nor U2069 (N_2069,N_890,N_784);
xor U2070 (N_2070,N_1458,N_1277);
nor U2071 (N_2071,N_1058,N_817);
nand U2072 (N_2072,N_1255,N_1492);
nor U2073 (N_2073,N_1061,N_1379);
nor U2074 (N_2074,N_1325,N_820);
and U2075 (N_2075,N_1068,N_1353);
nand U2076 (N_2076,N_1333,N_1267);
nor U2077 (N_2077,N_954,N_923);
nor U2078 (N_2078,N_913,N_865);
and U2079 (N_2079,N_957,N_1434);
and U2080 (N_2080,N_880,N_1262);
nand U2081 (N_2081,N_995,N_1082);
nor U2082 (N_2082,N_1007,N_754);
nor U2083 (N_2083,N_1024,N_912);
nand U2084 (N_2084,N_764,N_1437);
nand U2085 (N_2085,N_1076,N_1290);
and U2086 (N_2086,N_1237,N_1456);
nor U2087 (N_2087,N_1232,N_1009);
or U2088 (N_2088,N_1348,N_993);
nor U2089 (N_2089,N_926,N_927);
nand U2090 (N_2090,N_1420,N_1207);
nor U2091 (N_2091,N_1036,N_1463);
or U2092 (N_2092,N_1428,N_1200);
nor U2093 (N_2093,N_1036,N_1043);
or U2094 (N_2094,N_1043,N_1122);
nor U2095 (N_2095,N_1284,N_1371);
or U2096 (N_2096,N_1163,N_859);
and U2097 (N_2097,N_1221,N_981);
and U2098 (N_2098,N_1087,N_1262);
or U2099 (N_2099,N_804,N_1392);
nand U2100 (N_2100,N_870,N_1064);
or U2101 (N_2101,N_1156,N_1293);
nor U2102 (N_2102,N_1382,N_1275);
nor U2103 (N_2103,N_797,N_1459);
and U2104 (N_2104,N_1289,N_1202);
or U2105 (N_2105,N_1153,N_832);
and U2106 (N_2106,N_760,N_1480);
nand U2107 (N_2107,N_1366,N_1127);
or U2108 (N_2108,N_800,N_1457);
nor U2109 (N_2109,N_791,N_1324);
and U2110 (N_2110,N_1095,N_1285);
or U2111 (N_2111,N_948,N_1182);
nand U2112 (N_2112,N_1210,N_888);
and U2113 (N_2113,N_1070,N_956);
xor U2114 (N_2114,N_1392,N_1345);
nor U2115 (N_2115,N_790,N_1320);
or U2116 (N_2116,N_1316,N_1208);
nor U2117 (N_2117,N_1259,N_906);
xnor U2118 (N_2118,N_914,N_1476);
nand U2119 (N_2119,N_1371,N_1055);
nor U2120 (N_2120,N_1183,N_948);
and U2121 (N_2121,N_1114,N_1218);
nor U2122 (N_2122,N_1353,N_1099);
nor U2123 (N_2123,N_1173,N_1056);
or U2124 (N_2124,N_1206,N_833);
and U2125 (N_2125,N_940,N_775);
nor U2126 (N_2126,N_1430,N_933);
or U2127 (N_2127,N_783,N_1359);
and U2128 (N_2128,N_1024,N_1073);
nand U2129 (N_2129,N_814,N_887);
nor U2130 (N_2130,N_1358,N_851);
nand U2131 (N_2131,N_1024,N_1015);
and U2132 (N_2132,N_1406,N_1235);
nor U2133 (N_2133,N_1439,N_959);
or U2134 (N_2134,N_1258,N_1109);
xnor U2135 (N_2135,N_789,N_991);
nor U2136 (N_2136,N_1134,N_1097);
or U2137 (N_2137,N_1016,N_1144);
or U2138 (N_2138,N_1063,N_1489);
and U2139 (N_2139,N_1297,N_1178);
nor U2140 (N_2140,N_807,N_867);
or U2141 (N_2141,N_755,N_916);
or U2142 (N_2142,N_1196,N_1430);
and U2143 (N_2143,N_1404,N_1278);
and U2144 (N_2144,N_929,N_1155);
nor U2145 (N_2145,N_968,N_1027);
and U2146 (N_2146,N_1354,N_1374);
nor U2147 (N_2147,N_1308,N_1142);
and U2148 (N_2148,N_1039,N_1427);
nand U2149 (N_2149,N_1355,N_1448);
nand U2150 (N_2150,N_1274,N_1340);
and U2151 (N_2151,N_972,N_1147);
nor U2152 (N_2152,N_1010,N_796);
or U2153 (N_2153,N_1227,N_1191);
and U2154 (N_2154,N_1038,N_967);
and U2155 (N_2155,N_1266,N_1390);
nor U2156 (N_2156,N_1208,N_1449);
nand U2157 (N_2157,N_895,N_1435);
or U2158 (N_2158,N_1056,N_1044);
and U2159 (N_2159,N_1468,N_1256);
and U2160 (N_2160,N_1472,N_1256);
nand U2161 (N_2161,N_897,N_1062);
nand U2162 (N_2162,N_1254,N_1072);
or U2163 (N_2163,N_781,N_881);
nand U2164 (N_2164,N_1347,N_1019);
nor U2165 (N_2165,N_1431,N_1170);
or U2166 (N_2166,N_1215,N_1163);
xor U2167 (N_2167,N_758,N_1303);
and U2168 (N_2168,N_886,N_1009);
nor U2169 (N_2169,N_1433,N_1166);
nand U2170 (N_2170,N_1422,N_1492);
or U2171 (N_2171,N_1243,N_821);
nor U2172 (N_2172,N_908,N_1408);
nor U2173 (N_2173,N_1338,N_1433);
nor U2174 (N_2174,N_1132,N_1310);
or U2175 (N_2175,N_946,N_801);
or U2176 (N_2176,N_847,N_899);
nor U2177 (N_2177,N_1385,N_1483);
nor U2178 (N_2178,N_1357,N_1070);
or U2179 (N_2179,N_925,N_984);
and U2180 (N_2180,N_1473,N_1127);
nand U2181 (N_2181,N_1128,N_991);
or U2182 (N_2182,N_960,N_768);
nand U2183 (N_2183,N_1314,N_1289);
nor U2184 (N_2184,N_1079,N_773);
or U2185 (N_2185,N_1115,N_883);
and U2186 (N_2186,N_825,N_1273);
nand U2187 (N_2187,N_1263,N_850);
or U2188 (N_2188,N_957,N_817);
and U2189 (N_2189,N_1380,N_1230);
nand U2190 (N_2190,N_1394,N_1092);
or U2191 (N_2191,N_1175,N_1181);
nand U2192 (N_2192,N_1399,N_1046);
nor U2193 (N_2193,N_981,N_1201);
nor U2194 (N_2194,N_867,N_1161);
and U2195 (N_2195,N_1408,N_1183);
and U2196 (N_2196,N_1401,N_923);
nor U2197 (N_2197,N_798,N_1085);
and U2198 (N_2198,N_907,N_1116);
and U2199 (N_2199,N_780,N_783);
and U2200 (N_2200,N_1009,N_1004);
nor U2201 (N_2201,N_967,N_1416);
or U2202 (N_2202,N_1329,N_1138);
and U2203 (N_2203,N_1209,N_1432);
nand U2204 (N_2204,N_961,N_1107);
or U2205 (N_2205,N_961,N_1236);
nor U2206 (N_2206,N_1326,N_1254);
xnor U2207 (N_2207,N_975,N_1405);
nand U2208 (N_2208,N_865,N_929);
or U2209 (N_2209,N_1206,N_1312);
nor U2210 (N_2210,N_1005,N_782);
nor U2211 (N_2211,N_865,N_1374);
nand U2212 (N_2212,N_1013,N_1157);
and U2213 (N_2213,N_1181,N_1491);
or U2214 (N_2214,N_1415,N_922);
xor U2215 (N_2215,N_787,N_897);
or U2216 (N_2216,N_1035,N_1047);
or U2217 (N_2217,N_1088,N_1219);
and U2218 (N_2218,N_963,N_1137);
or U2219 (N_2219,N_1168,N_1294);
or U2220 (N_2220,N_882,N_1415);
or U2221 (N_2221,N_1386,N_1351);
and U2222 (N_2222,N_1357,N_1067);
or U2223 (N_2223,N_1074,N_943);
nor U2224 (N_2224,N_1419,N_1214);
nand U2225 (N_2225,N_924,N_1477);
and U2226 (N_2226,N_1089,N_1473);
nand U2227 (N_2227,N_848,N_1306);
or U2228 (N_2228,N_1420,N_1219);
and U2229 (N_2229,N_1442,N_1432);
nor U2230 (N_2230,N_849,N_1388);
nor U2231 (N_2231,N_1405,N_1268);
nand U2232 (N_2232,N_1349,N_936);
and U2233 (N_2233,N_1438,N_1381);
and U2234 (N_2234,N_1229,N_1496);
nor U2235 (N_2235,N_971,N_1219);
or U2236 (N_2236,N_1424,N_1449);
and U2237 (N_2237,N_751,N_1423);
or U2238 (N_2238,N_844,N_757);
or U2239 (N_2239,N_947,N_1283);
nand U2240 (N_2240,N_1220,N_1450);
nor U2241 (N_2241,N_756,N_1177);
and U2242 (N_2242,N_799,N_1193);
nor U2243 (N_2243,N_1437,N_1283);
and U2244 (N_2244,N_1221,N_794);
and U2245 (N_2245,N_1221,N_785);
nand U2246 (N_2246,N_905,N_1269);
or U2247 (N_2247,N_1264,N_946);
xnor U2248 (N_2248,N_1188,N_987);
or U2249 (N_2249,N_1395,N_965);
nor U2250 (N_2250,N_2021,N_2096);
or U2251 (N_2251,N_2181,N_2142);
xnor U2252 (N_2252,N_2173,N_2090);
and U2253 (N_2253,N_1961,N_1842);
or U2254 (N_2254,N_1881,N_1917);
nand U2255 (N_2255,N_2098,N_2193);
and U2256 (N_2256,N_1970,N_1716);
and U2257 (N_2257,N_1871,N_1965);
and U2258 (N_2258,N_1890,N_1987);
nand U2259 (N_2259,N_2145,N_1927);
nor U2260 (N_2260,N_1990,N_2224);
and U2261 (N_2261,N_2072,N_1648);
or U2262 (N_2262,N_1529,N_1571);
nor U2263 (N_2263,N_2029,N_1734);
nor U2264 (N_2264,N_1682,N_1891);
or U2265 (N_2265,N_2158,N_1999);
nand U2266 (N_2266,N_2019,N_2160);
and U2267 (N_2267,N_2079,N_2244);
or U2268 (N_2268,N_2035,N_1623);
or U2269 (N_2269,N_2034,N_1718);
nor U2270 (N_2270,N_2018,N_1906);
nand U2271 (N_2271,N_1786,N_1502);
and U2272 (N_2272,N_1725,N_1800);
nor U2273 (N_2273,N_1803,N_2107);
nor U2274 (N_2274,N_1962,N_2102);
and U2275 (N_2275,N_2191,N_1821);
nor U2276 (N_2276,N_2188,N_1645);
or U2277 (N_2277,N_2008,N_1951);
nor U2278 (N_2278,N_2056,N_1894);
or U2279 (N_2279,N_1833,N_1986);
nand U2280 (N_2280,N_2123,N_1575);
nand U2281 (N_2281,N_2184,N_1540);
and U2282 (N_2282,N_2016,N_2211);
nor U2283 (N_2283,N_1733,N_1602);
and U2284 (N_2284,N_1925,N_2045);
xor U2285 (N_2285,N_1895,N_1650);
and U2286 (N_2286,N_1554,N_1633);
nor U2287 (N_2287,N_2155,N_1939);
nor U2288 (N_2288,N_1992,N_1688);
or U2289 (N_2289,N_1964,N_1697);
and U2290 (N_2290,N_1875,N_1577);
and U2291 (N_2291,N_1611,N_2076);
or U2292 (N_2292,N_1840,N_1760);
and U2293 (N_2293,N_1983,N_2101);
nor U2294 (N_2294,N_1705,N_2138);
nand U2295 (N_2295,N_1956,N_1810);
or U2296 (N_2296,N_2068,N_1780);
nor U2297 (N_2297,N_1684,N_2215);
nand U2298 (N_2298,N_2206,N_1759);
nor U2299 (N_2299,N_2216,N_2219);
nand U2300 (N_2300,N_1566,N_2063);
nor U2301 (N_2301,N_1740,N_1945);
or U2302 (N_2302,N_2025,N_1896);
and U2303 (N_2303,N_1503,N_1706);
nand U2304 (N_2304,N_1629,N_2024);
or U2305 (N_2305,N_1795,N_1542);
nor U2306 (N_2306,N_1598,N_2128);
nor U2307 (N_2307,N_1715,N_1806);
or U2308 (N_2308,N_1973,N_1910);
and U2309 (N_2309,N_1663,N_2061);
nand U2310 (N_2310,N_2131,N_2065);
or U2311 (N_2311,N_1859,N_2106);
nand U2312 (N_2312,N_2242,N_1724);
or U2313 (N_2313,N_1752,N_2213);
nand U2314 (N_2314,N_1775,N_1589);
or U2315 (N_2315,N_1564,N_1957);
nand U2316 (N_2316,N_1730,N_1915);
or U2317 (N_2317,N_2185,N_2229);
and U2318 (N_2318,N_1664,N_1825);
nor U2319 (N_2319,N_1877,N_2230);
and U2320 (N_2320,N_1827,N_1707);
and U2321 (N_2321,N_1959,N_1818);
or U2322 (N_2322,N_2183,N_2051);
xor U2323 (N_2323,N_2031,N_1549);
or U2324 (N_2324,N_2201,N_2177);
or U2325 (N_2325,N_1860,N_1601);
nor U2326 (N_2326,N_1621,N_2140);
nand U2327 (N_2327,N_2156,N_2124);
nor U2328 (N_2328,N_1782,N_1632);
nor U2329 (N_2329,N_1661,N_2137);
nand U2330 (N_2330,N_1655,N_1704);
nand U2331 (N_2331,N_2148,N_1614);
or U2332 (N_2332,N_1755,N_2190);
or U2333 (N_2333,N_1835,N_1646);
or U2334 (N_2334,N_1527,N_1972);
nor U2335 (N_2335,N_1816,N_2133);
and U2336 (N_2336,N_2174,N_1720);
nand U2337 (N_2337,N_2228,N_1634);
and U2338 (N_2338,N_2146,N_1591);
or U2339 (N_2339,N_1955,N_1873);
and U2340 (N_2340,N_1599,N_1731);
or U2341 (N_2341,N_1558,N_2210);
and U2342 (N_2342,N_1801,N_1644);
and U2343 (N_2343,N_2083,N_2222);
nor U2344 (N_2344,N_2147,N_1659);
and U2345 (N_2345,N_2233,N_2057);
nor U2346 (N_2346,N_1674,N_2014);
and U2347 (N_2347,N_1952,N_1968);
or U2348 (N_2348,N_2087,N_1892);
nor U2349 (N_2349,N_1741,N_1565);
nor U2350 (N_2350,N_1950,N_2084);
nand U2351 (N_2351,N_1582,N_1938);
or U2352 (N_2352,N_1658,N_1605);
nor U2353 (N_2353,N_1905,N_1937);
or U2354 (N_2354,N_2163,N_2020);
nand U2355 (N_2355,N_1631,N_1505);
and U2356 (N_2356,N_1788,N_1732);
and U2357 (N_2357,N_1586,N_2246);
nor U2358 (N_2358,N_1642,N_1769);
or U2359 (N_2359,N_1531,N_2227);
nand U2360 (N_2360,N_2115,N_1792);
and U2361 (N_2361,N_1544,N_2036);
nand U2362 (N_2362,N_2169,N_2209);
nor U2363 (N_2363,N_1675,N_1597);
nor U2364 (N_2364,N_2004,N_2200);
or U2365 (N_2365,N_2129,N_1921);
or U2366 (N_2366,N_2192,N_1899);
nor U2367 (N_2367,N_1757,N_1666);
nand U2368 (N_2368,N_2135,N_1609);
and U2369 (N_2369,N_1504,N_1943);
and U2370 (N_2370,N_1750,N_2226);
nand U2371 (N_2371,N_1814,N_1779);
and U2372 (N_2372,N_2125,N_1912);
or U2373 (N_2373,N_1619,N_1735);
nand U2374 (N_2374,N_1858,N_1539);
xor U2375 (N_2375,N_1712,N_1713);
or U2376 (N_2376,N_1738,N_1668);
nor U2377 (N_2377,N_2232,N_1954);
and U2378 (N_2378,N_1919,N_1533);
nor U2379 (N_2379,N_2122,N_2187);
nand U2380 (N_2380,N_1656,N_1940);
nand U2381 (N_2381,N_1717,N_1880);
nor U2382 (N_2382,N_2127,N_1924);
nand U2383 (N_2383,N_2237,N_2052);
nand U2384 (N_2384,N_1811,N_1887);
and U2385 (N_2385,N_2134,N_1514);
nand U2386 (N_2386,N_1676,N_1883);
nor U2387 (N_2387,N_2104,N_1728);
nand U2388 (N_2388,N_1703,N_1680);
and U2389 (N_2389,N_1907,N_2006);
nor U2390 (N_2390,N_2105,N_2199);
and U2391 (N_2391,N_1702,N_2207);
or U2392 (N_2392,N_1652,N_2015);
and U2393 (N_2393,N_2017,N_1976);
nor U2394 (N_2394,N_1530,N_1861);
or U2395 (N_2395,N_2003,N_1622);
or U2396 (N_2396,N_1626,N_2011);
nand U2397 (N_2397,N_1620,N_1552);
nand U2398 (N_2398,N_1832,N_1984);
nor U2399 (N_2399,N_1721,N_1639);
or U2400 (N_2400,N_1831,N_1600);
nand U2401 (N_2401,N_1635,N_1689);
and U2402 (N_2402,N_1617,N_1926);
and U2403 (N_2403,N_2172,N_1537);
or U2404 (N_2404,N_1572,N_1574);
or U2405 (N_2405,N_2117,N_1903);
or U2406 (N_2406,N_1855,N_1882);
nand U2407 (N_2407,N_1677,N_2223);
and U2408 (N_2408,N_1931,N_1561);
nand U2409 (N_2409,N_1746,N_1590);
or U2410 (N_2410,N_1515,N_2198);
and U2411 (N_2411,N_1579,N_1947);
nand U2412 (N_2412,N_2077,N_1796);
nor U2413 (N_2413,N_2053,N_1603);
nor U2414 (N_2414,N_1773,N_1979);
nand U2415 (N_2415,N_2126,N_1874);
and U2416 (N_2416,N_2103,N_1920);
nand U2417 (N_2417,N_1576,N_2151);
nor U2418 (N_2418,N_1928,N_1908);
nor U2419 (N_2419,N_1616,N_1567);
and U2420 (N_2420,N_1672,N_1797);
nand U2421 (N_2421,N_1607,N_1748);
nand U2422 (N_2422,N_1966,N_1865);
nor U2423 (N_2423,N_2038,N_1798);
and U2424 (N_2424,N_2085,N_2136);
nand U2425 (N_2425,N_2248,N_2054);
nand U2426 (N_2426,N_1808,N_1876);
and U2427 (N_2427,N_1563,N_1555);
nand U2428 (N_2428,N_1692,N_1932);
or U2429 (N_2429,N_1830,N_2153);
or U2430 (N_2430,N_2247,N_2217);
or U2431 (N_2431,N_2075,N_1678);
or U2432 (N_2432,N_1823,N_1868);
nand U2433 (N_2433,N_2152,N_1548);
and U2434 (N_2434,N_2204,N_1596);
or U2435 (N_2435,N_1888,N_1991);
nand U2436 (N_2436,N_1758,N_2108);
nor U2437 (N_2437,N_1649,N_1651);
nand U2438 (N_2438,N_1570,N_1534);
nand U2439 (N_2439,N_2099,N_1606);
and U2440 (N_2440,N_2205,N_1820);
and U2441 (N_2441,N_1739,N_2009);
or U2442 (N_2442,N_1569,N_1517);
nand U2443 (N_2443,N_1995,N_2249);
nand U2444 (N_2444,N_1884,N_2010);
nor U2445 (N_2445,N_1761,N_2040);
or U2446 (N_2446,N_1568,N_2070);
nor U2447 (N_2447,N_1710,N_2157);
and U2448 (N_2448,N_1694,N_2114);
nand U2449 (N_2449,N_1764,N_2120);
or U2450 (N_2450,N_2082,N_1687);
nand U2451 (N_2451,N_1774,N_1793);
nor U2452 (N_2452,N_2243,N_1523);
or U2453 (N_2453,N_1857,N_1847);
nor U2454 (N_2454,N_1893,N_2012);
nand U2455 (N_2455,N_2058,N_1854);
nand U2456 (N_2456,N_2037,N_1749);
and U2457 (N_2457,N_1958,N_1982);
xnor U2458 (N_2458,N_2027,N_2095);
or U2459 (N_2459,N_1993,N_1641);
nand U2460 (N_2460,N_1989,N_1864);
or U2461 (N_2461,N_2071,N_1580);
nand U2462 (N_2462,N_1509,N_1513);
nor U2463 (N_2463,N_2176,N_1777);
and U2464 (N_2464,N_1822,N_1543);
or U2465 (N_2465,N_1998,N_1772);
and U2466 (N_2466,N_1547,N_2033);
and U2467 (N_2467,N_2047,N_1595);
or U2468 (N_2468,N_1671,N_2064);
nor U2469 (N_2469,N_1771,N_1685);
and U2470 (N_2470,N_1546,N_2221);
nor U2471 (N_2471,N_1557,N_1667);
nand U2472 (N_2472,N_2043,N_1980);
nand U2473 (N_2473,N_2195,N_1963);
nor U2474 (N_2474,N_2144,N_1985);
or U2475 (N_2475,N_1695,N_1532);
nand U2476 (N_2476,N_1636,N_1708);
nor U2477 (N_2477,N_2166,N_1785);
and U2478 (N_2478,N_1654,N_1657);
and U2479 (N_2479,N_2225,N_1845);
or U2480 (N_2480,N_1824,N_1754);
nand U2481 (N_2481,N_1693,N_1809);
nor U2482 (N_2482,N_1829,N_2179);
and U2483 (N_2483,N_1977,N_1519);
or U2484 (N_2484,N_1935,N_1528);
nand U2485 (N_2485,N_1813,N_2030);
nor U2486 (N_2486,N_1767,N_2100);
and U2487 (N_2487,N_1608,N_1879);
or U2488 (N_2488,N_1711,N_1747);
nor U2489 (N_2489,N_1851,N_1585);
or U2490 (N_2490,N_1506,N_1904);
or U2491 (N_2491,N_2159,N_2007);
and U2492 (N_2492,N_1518,N_2055);
and U2493 (N_2493,N_1545,N_2202);
and U2494 (N_2494,N_1709,N_1610);
nand U2495 (N_2495,N_2164,N_1913);
nor U2496 (N_2496,N_2121,N_1683);
and U2497 (N_2497,N_1784,N_1743);
nor U2498 (N_2498,N_1897,N_1673);
nand U2499 (N_2499,N_1560,N_2214);
and U2500 (N_2500,N_1768,N_1587);
nand U2501 (N_2501,N_2239,N_2231);
and U2502 (N_2502,N_2039,N_2132);
and U2503 (N_2503,N_1512,N_1719);
or U2504 (N_2504,N_1524,N_1593);
and U2505 (N_2505,N_1878,N_1885);
and U2506 (N_2506,N_2240,N_2212);
nor U2507 (N_2507,N_2118,N_2023);
and U2508 (N_2508,N_1508,N_1604);
and U2509 (N_2509,N_1624,N_2241);
nor U2510 (N_2510,N_2002,N_1838);
nor U2511 (N_2511,N_1948,N_1862);
and U2512 (N_2512,N_1691,N_2026);
and U2513 (N_2513,N_2170,N_1870);
nor U2514 (N_2514,N_2180,N_1553);
nand U2515 (N_2515,N_1933,N_1536);
and U2516 (N_2516,N_1849,N_1812);
nand U2517 (N_2517,N_1776,N_2046);
nor U2518 (N_2518,N_1500,N_1612);
or U2519 (N_2519,N_1722,N_2097);
and U2520 (N_2520,N_2130,N_1974);
xor U2521 (N_2521,N_1791,N_1510);
nor U2522 (N_2522,N_2175,N_1872);
or U2523 (N_2523,N_1916,N_1742);
or U2524 (N_2524,N_1643,N_1936);
and U2525 (N_2525,N_1930,N_1783);
xor U2526 (N_2526,N_1737,N_1686);
and U2527 (N_2527,N_2186,N_1638);
or U2528 (N_2528,N_1751,N_1766);
or U2529 (N_2529,N_1627,N_1846);
or U2530 (N_2530,N_1837,N_2141);
nor U2531 (N_2531,N_2161,N_1844);
nor U2532 (N_2532,N_1898,N_2001);
and U2533 (N_2533,N_1781,N_1994);
nor U2534 (N_2534,N_1807,N_2112);
nor U2535 (N_2535,N_1856,N_1853);
nand U2536 (N_2536,N_1647,N_1852);
nand U2537 (N_2537,N_2032,N_1723);
nand U2538 (N_2538,N_1918,N_1726);
and U2539 (N_2539,N_2208,N_2168);
and U2540 (N_2540,N_1516,N_1714);
nor U2541 (N_2541,N_1802,N_2167);
nand U2542 (N_2542,N_2116,N_2088);
or U2543 (N_2543,N_1690,N_2194);
nor U2544 (N_2544,N_1670,N_2078);
and U2545 (N_2545,N_1628,N_1805);
or U2546 (N_2546,N_2049,N_2091);
nand U2547 (N_2547,N_1573,N_1538);
and U2548 (N_2548,N_1799,N_1848);
nor U2549 (N_2549,N_1615,N_2074);
or U2550 (N_2550,N_1946,N_1637);
nor U2551 (N_2551,N_1909,N_2245);
nand U2552 (N_2552,N_1886,N_1839);
nand U2553 (N_2553,N_1756,N_2109);
or U2554 (N_2554,N_1763,N_2110);
nand U2555 (N_2555,N_1559,N_2189);
or U2556 (N_2556,N_2235,N_1583);
and U2557 (N_2557,N_2220,N_2013);
or U2558 (N_2558,N_2196,N_1790);
nand U2559 (N_2559,N_1618,N_2094);
xnor U2560 (N_2560,N_1975,N_1789);
nand U2561 (N_2561,N_1541,N_1625);
and U2562 (N_2562,N_1902,N_2067);
or U2563 (N_2563,N_2139,N_1841);
nor U2564 (N_2564,N_2028,N_2197);
or U2565 (N_2565,N_1511,N_1679);
or U2566 (N_2566,N_1929,N_2093);
and U2567 (N_2567,N_2238,N_1550);
nor U2568 (N_2568,N_1727,N_1665);
nor U2569 (N_2569,N_1914,N_1949);
or U2570 (N_2570,N_1850,N_1971);
or U2571 (N_2571,N_2182,N_2234);
and U2572 (N_2572,N_2060,N_1526);
and U2573 (N_2573,N_1923,N_2236);
nand U2574 (N_2574,N_1942,N_1501);
and U2575 (N_2575,N_2111,N_1594);
and U2576 (N_2576,N_1815,N_2081);
and U2577 (N_2577,N_2048,N_2162);
nand U2578 (N_2578,N_1765,N_1834);
and U2579 (N_2579,N_1843,N_1869);
or U2580 (N_2580,N_1535,N_2119);
or U2581 (N_2581,N_1522,N_1698);
nor U2582 (N_2582,N_1967,N_1787);
nor U2583 (N_2583,N_1900,N_1969);
and U2584 (N_2584,N_1699,N_1588);
or U2585 (N_2585,N_1520,N_2092);
and U2586 (N_2586,N_1753,N_1669);
and U2587 (N_2587,N_1770,N_2069);
and U2588 (N_2588,N_1613,N_1997);
or U2589 (N_2589,N_1525,N_1662);
nor U2590 (N_2590,N_2022,N_1578);
nor U2591 (N_2591,N_1640,N_2150);
and U2592 (N_2592,N_1701,N_1826);
and U2593 (N_2593,N_2143,N_1867);
and U2594 (N_2594,N_1581,N_1744);
nor U2595 (N_2595,N_1630,N_1817);
nor U2596 (N_2596,N_1729,N_2000);
and U2597 (N_2597,N_1866,N_1863);
and U2598 (N_2598,N_1804,N_1978);
and U2599 (N_2599,N_1551,N_2066);
nand U2600 (N_2600,N_1584,N_1988);
or U2601 (N_2601,N_1922,N_2073);
nor U2602 (N_2602,N_2218,N_1653);
or U2603 (N_2603,N_1521,N_1696);
or U2604 (N_2604,N_1996,N_2005);
and U2605 (N_2605,N_2044,N_2080);
nand U2606 (N_2606,N_1507,N_2154);
nor U2607 (N_2607,N_2178,N_1562);
or U2608 (N_2608,N_1794,N_1778);
and U2609 (N_2609,N_1745,N_1592);
and U2610 (N_2610,N_1736,N_2089);
and U2611 (N_2611,N_1660,N_2171);
nand U2612 (N_2612,N_2050,N_2059);
or U2613 (N_2613,N_2041,N_1556);
nor U2614 (N_2614,N_2203,N_1836);
nand U2615 (N_2615,N_1828,N_1901);
nand U2616 (N_2616,N_1981,N_1953);
and U2617 (N_2617,N_1944,N_2149);
nor U2618 (N_2618,N_1681,N_1762);
nand U2619 (N_2619,N_2113,N_1700);
and U2620 (N_2620,N_1911,N_1941);
or U2621 (N_2621,N_1819,N_2042);
or U2622 (N_2622,N_1889,N_2165);
and U2623 (N_2623,N_1934,N_1960);
or U2624 (N_2624,N_2086,N_2062);
nand U2625 (N_2625,N_1665,N_2174);
nand U2626 (N_2626,N_1739,N_2071);
and U2627 (N_2627,N_1532,N_1725);
or U2628 (N_2628,N_1933,N_1505);
nor U2629 (N_2629,N_1838,N_1753);
nand U2630 (N_2630,N_2018,N_2237);
nand U2631 (N_2631,N_1672,N_1521);
nand U2632 (N_2632,N_2015,N_1527);
and U2633 (N_2633,N_2029,N_2025);
nand U2634 (N_2634,N_1832,N_1991);
nor U2635 (N_2635,N_1835,N_1596);
nor U2636 (N_2636,N_2037,N_1904);
or U2637 (N_2637,N_2210,N_1634);
nand U2638 (N_2638,N_2195,N_1932);
nand U2639 (N_2639,N_1984,N_2139);
nand U2640 (N_2640,N_1970,N_1991);
nor U2641 (N_2641,N_1942,N_1878);
and U2642 (N_2642,N_1754,N_1998);
or U2643 (N_2643,N_1550,N_2224);
or U2644 (N_2644,N_1943,N_1958);
or U2645 (N_2645,N_1845,N_2108);
or U2646 (N_2646,N_2132,N_1802);
or U2647 (N_2647,N_2077,N_1652);
xnor U2648 (N_2648,N_1589,N_2145);
nor U2649 (N_2649,N_1878,N_1755);
nand U2650 (N_2650,N_1807,N_2181);
and U2651 (N_2651,N_1791,N_2142);
nor U2652 (N_2652,N_1533,N_2176);
or U2653 (N_2653,N_2156,N_2088);
and U2654 (N_2654,N_1604,N_1876);
nor U2655 (N_2655,N_1886,N_2242);
nand U2656 (N_2656,N_1659,N_1618);
or U2657 (N_2657,N_2030,N_1613);
and U2658 (N_2658,N_1699,N_2147);
nand U2659 (N_2659,N_1990,N_1913);
nand U2660 (N_2660,N_2020,N_1661);
nand U2661 (N_2661,N_2235,N_1760);
nand U2662 (N_2662,N_2038,N_2004);
nor U2663 (N_2663,N_2016,N_2088);
nor U2664 (N_2664,N_1533,N_2164);
or U2665 (N_2665,N_1997,N_2029);
nor U2666 (N_2666,N_1888,N_1734);
or U2667 (N_2667,N_2200,N_2050);
xnor U2668 (N_2668,N_1683,N_2044);
nand U2669 (N_2669,N_2111,N_2244);
nand U2670 (N_2670,N_2072,N_1723);
nor U2671 (N_2671,N_1536,N_1502);
nand U2672 (N_2672,N_1924,N_1708);
and U2673 (N_2673,N_1911,N_2140);
or U2674 (N_2674,N_1883,N_1579);
and U2675 (N_2675,N_1541,N_2051);
and U2676 (N_2676,N_1957,N_2018);
nor U2677 (N_2677,N_1947,N_1605);
or U2678 (N_2678,N_2171,N_1732);
and U2679 (N_2679,N_1788,N_1632);
and U2680 (N_2680,N_1873,N_1740);
or U2681 (N_2681,N_1967,N_1685);
nor U2682 (N_2682,N_2097,N_2121);
nor U2683 (N_2683,N_2246,N_1812);
or U2684 (N_2684,N_2195,N_1637);
and U2685 (N_2685,N_1647,N_2128);
nand U2686 (N_2686,N_2187,N_2103);
xnor U2687 (N_2687,N_1503,N_1658);
nor U2688 (N_2688,N_2066,N_2027);
or U2689 (N_2689,N_2097,N_1704);
and U2690 (N_2690,N_2091,N_1724);
and U2691 (N_2691,N_1624,N_2164);
nand U2692 (N_2692,N_1934,N_1551);
nor U2693 (N_2693,N_2019,N_2062);
nand U2694 (N_2694,N_1700,N_1546);
and U2695 (N_2695,N_1734,N_2025);
or U2696 (N_2696,N_1673,N_1941);
nor U2697 (N_2697,N_1757,N_1637);
nor U2698 (N_2698,N_2188,N_1992);
and U2699 (N_2699,N_1537,N_1727);
nor U2700 (N_2700,N_2082,N_2025);
and U2701 (N_2701,N_2011,N_1757);
or U2702 (N_2702,N_1501,N_1758);
and U2703 (N_2703,N_1590,N_2109);
nand U2704 (N_2704,N_2227,N_2179);
and U2705 (N_2705,N_2118,N_1592);
or U2706 (N_2706,N_2066,N_2079);
or U2707 (N_2707,N_1715,N_1712);
and U2708 (N_2708,N_1706,N_2112);
nand U2709 (N_2709,N_1800,N_1784);
and U2710 (N_2710,N_1706,N_1879);
nand U2711 (N_2711,N_1861,N_1600);
nand U2712 (N_2712,N_2130,N_1946);
nor U2713 (N_2713,N_1800,N_1521);
or U2714 (N_2714,N_2140,N_1977);
xnor U2715 (N_2715,N_1778,N_1702);
nor U2716 (N_2716,N_1786,N_1906);
nand U2717 (N_2717,N_2240,N_1932);
nor U2718 (N_2718,N_1779,N_1578);
nor U2719 (N_2719,N_1680,N_1561);
nor U2720 (N_2720,N_1702,N_1516);
xnor U2721 (N_2721,N_2193,N_2003);
and U2722 (N_2722,N_2021,N_1872);
and U2723 (N_2723,N_1809,N_1772);
and U2724 (N_2724,N_1893,N_2142);
nand U2725 (N_2725,N_1621,N_1673);
nand U2726 (N_2726,N_1858,N_1660);
nand U2727 (N_2727,N_2167,N_1874);
nor U2728 (N_2728,N_1529,N_1942);
nor U2729 (N_2729,N_1531,N_1625);
nand U2730 (N_2730,N_1663,N_1566);
and U2731 (N_2731,N_1664,N_1557);
and U2732 (N_2732,N_1881,N_2131);
and U2733 (N_2733,N_1748,N_2026);
or U2734 (N_2734,N_1576,N_1695);
nor U2735 (N_2735,N_1513,N_1829);
nor U2736 (N_2736,N_1870,N_1954);
or U2737 (N_2737,N_1990,N_1897);
and U2738 (N_2738,N_1958,N_2017);
or U2739 (N_2739,N_2005,N_1520);
or U2740 (N_2740,N_1546,N_1773);
and U2741 (N_2741,N_1828,N_2063);
or U2742 (N_2742,N_2103,N_1583);
nor U2743 (N_2743,N_1715,N_1601);
and U2744 (N_2744,N_1510,N_1683);
and U2745 (N_2745,N_1911,N_1815);
nor U2746 (N_2746,N_1533,N_1806);
or U2747 (N_2747,N_2159,N_1505);
or U2748 (N_2748,N_1950,N_2065);
nor U2749 (N_2749,N_2000,N_1846);
or U2750 (N_2750,N_2036,N_2144);
and U2751 (N_2751,N_1522,N_2129);
and U2752 (N_2752,N_1529,N_1778);
and U2753 (N_2753,N_1719,N_1703);
nand U2754 (N_2754,N_1677,N_1705);
or U2755 (N_2755,N_2153,N_1650);
or U2756 (N_2756,N_1864,N_1979);
xnor U2757 (N_2757,N_1618,N_2063);
or U2758 (N_2758,N_2002,N_1770);
nand U2759 (N_2759,N_2239,N_1560);
or U2760 (N_2760,N_1729,N_1642);
or U2761 (N_2761,N_2015,N_2160);
or U2762 (N_2762,N_2202,N_2064);
nand U2763 (N_2763,N_1817,N_2164);
nor U2764 (N_2764,N_1680,N_1817);
nor U2765 (N_2765,N_1508,N_2028);
or U2766 (N_2766,N_1742,N_1868);
nor U2767 (N_2767,N_1529,N_1784);
and U2768 (N_2768,N_2063,N_1865);
or U2769 (N_2769,N_2143,N_1935);
and U2770 (N_2770,N_1671,N_2027);
nor U2771 (N_2771,N_2072,N_1789);
nor U2772 (N_2772,N_2119,N_1600);
nor U2773 (N_2773,N_1881,N_1814);
and U2774 (N_2774,N_1692,N_1513);
nand U2775 (N_2775,N_1645,N_1643);
nor U2776 (N_2776,N_1661,N_2120);
and U2777 (N_2777,N_1904,N_1533);
nand U2778 (N_2778,N_1647,N_1788);
nand U2779 (N_2779,N_1671,N_1634);
nand U2780 (N_2780,N_1672,N_1917);
or U2781 (N_2781,N_1778,N_1701);
nor U2782 (N_2782,N_2001,N_1807);
nand U2783 (N_2783,N_1818,N_1624);
and U2784 (N_2784,N_2169,N_1874);
and U2785 (N_2785,N_2184,N_2138);
and U2786 (N_2786,N_1813,N_2218);
nand U2787 (N_2787,N_2054,N_2122);
or U2788 (N_2788,N_1965,N_1814);
or U2789 (N_2789,N_1560,N_1703);
or U2790 (N_2790,N_1933,N_1994);
or U2791 (N_2791,N_2071,N_1782);
nand U2792 (N_2792,N_1518,N_1554);
or U2793 (N_2793,N_1806,N_1816);
or U2794 (N_2794,N_1868,N_1599);
or U2795 (N_2795,N_2018,N_1530);
and U2796 (N_2796,N_1960,N_2100);
nor U2797 (N_2797,N_1998,N_1755);
nor U2798 (N_2798,N_1772,N_1831);
and U2799 (N_2799,N_1714,N_2135);
nand U2800 (N_2800,N_2145,N_2049);
and U2801 (N_2801,N_1945,N_1794);
nor U2802 (N_2802,N_1995,N_1501);
or U2803 (N_2803,N_1911,N_1622);
and U2804 (N_2804,N_1679,N_1988);
and U2805 (N_2805,N_2234,N_1696);
and U2806 (N_2806,N_1618,N_1603);
and U2807 (N_2807,N_2187,N_2005);
and U2808 (N_2808,N_2164,N_2046);
and U2809 (N_2809,N_1747,N_2144);
or U2810 (N_2810,N_1868,N_1531);
and U2811 (N_2811,N_2196,N_1743);
nand U2812 (N_2812,N_1534,N_1967);
nand U2813 (N_2813,N_2074,N_1764);
nor U2814 (N_2814,N_1860,N_1923);
and U2815 (N_2815,N_1510,N_1639);
nand U2816 (N_2816,N_1556,N_1812);
and U2817 (N_2817,N_1861,N_2218);
or U2818 (N_2818,N_1884,N_2125);
nor U2819 (N_2819,N_1534,N_1852);
or U2820 (N_2820,N_2190,N_1861);
nor U2821 (N_2821,N_2110,N_1992);
and U2822 (N_2822,N_2049,N_1986);
nor U2823 (N_2823,N_1969,N_2219);
and U2824 (N_2824,N_1500,N_2172);
nor U2825 (N_2825,N_1573,N_1860);
nand U2826 (N_2826,N_2089,N_1678);
and U2827 (N_2827,N_1791,N_2202);
nor U2828 (N_2828,N_2107,N_1888);
or U2829 (N_2829,N_1788,N_1882);
nand U2830 (N_2830,N_1621,N_1797);
or U2831 (N_2831,N_1602,N_2034);
or U2832 (N_2832,N_1663,N_1719);
and U2833 (N_2833,N_1661,N_1565);
or U2834 (N_2834,N_1838,N_1892);
or U2835 (N_2835,N_1702,N_2112);
nor U2836 (N_2836,N_2093,N_1835);
and U2837 (N_2837,N_2207,N_1719);
or U2838 (N_2838,N_1642,N_2135);
nor U2839 (N_2839,N_1905,N_1623);
and U2840 (N_2840,N_1757,N_2010);
nor U2841 (N_2841,N_1643,N_2180);
nor U2842 (N_2842,N_1762,N_1724);
or U2843 (N_2843,N_2226,N_1543);
and U2844 (N_2844,N_2015,N_1695);
or U2845 (N_2845,N_2131,N_2145);
nor U2846 (N_2846,N_1812,N_2057);
nand U2847 (N_2847,N_2139,N_2002);
and U2848 (N_2848,N_2118,N_1965);
and U2849 (N_2849,N_1704,N_1873);
and U2850 (N_2850,N_1991,N_1543);
or U2851 (N_2851,N_1806,N_1981);
and U2852 (N_2852,N_1533,N_1862);
nor U2853 (N_2853,N_1883,N_1525);
or U2854 (N_2854,N_1917,N_1555);
nand U2855 (N_2855,N_2225,N_2176);
nand U2856 (N_2856,N_2030,N_2165);
and U2857 (N_2857,N_2242,N_2217);
nor U2858 (N_2858,N_1671,N_1517);
nor U2859 (N_2859,N_2005,N_1723);
or U2860 (N_2860,N_1870,N_1716);
nand U2861 (N_2861,N_1625,N_1816);
xnor U2862 (N_2862,N_1649,N_2227);
nand U2863 (N_2863,N_1909,N_1826);
and U2864 (N_2864,N_1932,N_2208);
and U2865 (N_2865,N_1699,N_1689);
nor U2866 (N_2866,N_1921,N_2080);
and U2867 (N_2867,N_1934,N_2123);
and U2868 (N_2868,N_1951,N_1853);
nand U2869 (N_2869,N_2123,N_1859);
or U2870 (N_2870,N_1547,N_1783);
nand U2871 (N_2871,N_1930,N_1819);
and U2872 (N_2872,N_1669,N_2231);
nand U2873 (N_2873,N_1958,N_1863);
or U2874 (N_2874,N_1840,N_2173);
nor U2875 (N_2875,N_1723,N_1604);
nor U2876 (N_2876,N_1643,N_1980);
nand U2877 (N_2877,N_2020,N_1819);
nor U2878 (N_2878,N_1796,N_2199);
nor U2879 (N_2879,N_2113,N_1840);
or U2880 (N_2880,N_1646,N_2130);
or U2881 (N_2881,N_2213,N_2010);
or U2882 (N_2882,N_1642,N_1672);
and U2883 (N_2883,N_2216,N_1749);
and U2884 (N_2884,N_1504,N_1817);
or U2885 (N_2885,N_2093,N_1695);
or U2886 (N_2886,N_1647,N_1523);
nor U2887 (N_2887,N_2063,N_1636);
nand U2888 (N_2888,N_2112,N_1811);
nand U2889 (N_2889,N_1843,N_1637);
nor U2890 (N_2890,N_1846,N_2173);
nor U2891 (N_2891,N_2059,N_1837);
and U2892 (N_2892,N_1824,N_2129);
nand U2893 (N_2893,N_1566,N_1744);
nor U2894 (N_2894,N_1535,N_1661);
nor U2895 (N_2895,N_1668,N_2102);
or U2896 (N_2896,N_1716,N_2032);
and U2897 (N_2897,N_1979,N_2025);
nand U2898 (N_2898,N_1551,N_2101);
nor U2899 (N_2899,N_2198,N_1604);
nor U2900 (N_2900,N_2088,N_1732);
nand U2901 (N_2901,N_1560,N_2201);
or U2902 (N_2902,N_2141,N_2087);
or U2903 (N_2903,N_2066,N_1855);
nor U2904 (N_2904,N_1821,N_1711);
or U2905 (N_2905,N_1926,N_2149);
nor U2906 (N_2906,N_1651,N_2003);
or U2907 (N_2907,N_1630,N_1632);
nor U2908 (N_2908,N_1895,N_1568);
nand U2909 (N_2909,N_1930,N_1914);
nor U2910 (N_2910,N_1691,N_2002);
xnor U2911 (N_2911,N_1813,N_1545);
nand U2912 (N_2912,N_1754,N_1513);
or U2913 (N_2913,N_1971,N_1840);
nand U2914 (N_2914,N_2153,N_1987);
nor U2915 (N_2915,N_1823,N_1712);
xor U2916 (N_2916,N_1925,N_1843);
or U2917 (N_2917,N_1941,N_1777);
nor U2918 (N_2918,N_1666,N_2132);
or U2919 (N_2919,N_2188,N_2008);
nor U2920 (N_2920,N_2056,N_2023);
nand U2921 (N_2921,N_1834,N_2157);
nor U2922 (N_2922,N_1559,N_1916);
and U2923 (N_2923,N_1702,N_1635);
nor U2924 (N_2924,N_1836,N_1904);
nand U2925 (N_2925,N_2197,N_1874);
nor U2926 (N_2926,N_1592,N_1958);
and U2927 (N_2927,N_1937,N_1876);
or U2928 (N_2928,N_2178,N_2157);
and U2929 (N_2929,N_1786,N_1630);
or U2930 (N_2930,N_1829,N_1559);
or U2931 (N_2931,N_1917,N_1592);
nand U2932 (N_2932,N_2011,N_2168);
and U2933 (N_2933,N_1782,N_2049);
or U2934 (N_2934,N_2213,N_1620);
or U2935 (N_2935,N_2215,N_2001);
or U2936 (N_2936,N_2127,N_1661);
or U2937 (N_2937,N_2150,N_1599);
and U2938 (N_2938,N_1526,N_2225);
or U2939 (N_2939,N_1556,N_2236);
nor U2940 (N_2940,N_1993,N_1965);
or U2941 (N_2941,N_1848,N_1701);
or U2942 (N_2942,N_2036,N_1730);
and U2943 (N_2943,N_1937,N_1955);
and U2944 (N_2944,N_1974,N_1511);
and U2945 (N_2945,N_1888,N_1708);
or U2946 (N_2946,N_1889,N_1818);
or U2947 (N_2947,N_2071,N_1525);
nor U2948 (N_2948,N_1626,N_2186);
or U2949 (N_2949,N_2230,N_1552);
nor U2950 (N_2950,N_1608,N_1681);
nand U2951 (N_2951,N_1578,N_1754);
or U2952 (N_2952,N_2170,N_1862);
nor U2953 (N_2953,N_2146,N_2188);
or U2954 (N_2954,N_1580,N_1999);
and U2955 (N_2955,N_1768,N_1630);
nor U2956 (N_2956,N_2051,N_1708);
xnor U2957 (N_2957,N_1593,N_1713);
nor U2958 (N_2958,N_1665,N_1952);
nand U2959 (N_2959,N_1677,N_1920);
and U2960 (N_2960,N_2150,N_1603);
and U2961 (N_2961,N_1631,N_1822);
or U2962 (N_2962,N_2183,N_1601);
nand U2963 (N_2963,N_2206,N_2064);
nor U2964 (N_2964,N_1929,N_2104);
nor U2965 (N_2965,N_1716,N_1932);
and U2966 (N_2966,N_1587,N_1559);
or U2967 (N_2967,N_2174,N_1788);
or U2968 (N_2968,N_1897,N_2226);
and U2969 (N_2969,N_2249,N_1559);
nor U2970 (N_2970,N_2201,N_1982);
or U2971 (N_2971,N_2094,N_1687);
and U2972 (N_2972,N_2142,N_2121);
nand U2973 (N_2973,N_2052,N_1579);
or U2974 (N_2974,N_2142,N_1735);
and U2975 (N_2975,N_1730,N_1645);
nor U2976 (N_2976,N_1889,N_1759);
nor U2977 (N_2977,N_2098,N_1846);
xor U2978 (N_2978,N_1786,N_1700);
nor U2979 (N_2979,N_1719,N_2129);
nand U2980 (N_2980,N_2015,N_1971);
nand U2981 (N_2981,N_1713,N_1510);
and U2982 (N_2982,N_1585,N_1745);
or U2983 (N_2983,N_1763,N_2247);
nor U2984 (N_2984,N_2147,N_2034);
and U2985 (N_2985,N_2006,N_2054);
or U2986 (N_2986,N_1548,N_1532);
or U2987 (N_2987,N_1685,N_1868);
and U2988 (N_2988,N_2114,N_1549);
and U2989 (N_2989,N_1988,N_1738);
and U2990 (N_2990,N_2096,N_1798);
or U2991 (N_2991,N_2172,N_1631);
nand U2992 (N_2992,N_2149,N_2208);
nor U2993 (N_2993,N_2095,N_2199);
nand U2994 (N_2994,N_2236,N_2042);
nor U2995 (N_2995,N_1678,N_1565);
nand U2996 (N_2996,N_1756,N_1766);
and U2997 (N_2997,N_1868,N_1550);
or U2998 (N_2998,N_2215,N_1671);
or U2999 (N_2999,N_2051,N_1527);
or U3000 (N_3000,N_2915,N_2415);
or U3001 (N_3001,N_2457,N_2344);
or U3002 (N_3002,N_2724,N_2660);
or U3003 (N_3003,N_2402,N_2866);
nor U3004 (N_3004,N_2341,N_2364);
or U3005 (N_3005,N_2510,N_2285);
and U3006 (N_3006,N_2560,N_2908);
or U3007 (N_3007,N_2472,N_2338);
nand U3008 (N_3008,N_2808,N_2625);
nor U3009 (N_3009,N_2500,N_2283);
nand U3010 (N_3010,N_2569,N_2925);
or U3011 (N_3011,N_2731,N_2685);
or U3012 (N_3012,N_2888,N_2860);
or U3013 (N_3013,N_2922,N_2273);
nor U3014 (N_3014,N_2811,N_2828);
nor U3015 (N_3015,N_2679,N_2920);
and U3016 (N_3016,N_2473,N_2862);
and U3017 (N_3017,N_2382,N_2841);
xor U3018 (N_3018,N_2825,N_2947);
or U3019 (N_3019,N_2969,N_2881);
nand U3020 (N_3020,N_2777,N_2766);
and U3021 (N_3021,N_2697,N_2883);
nand U3022 (N_3022,N_2315,N_2870);
or U3023 (N_3023,N_2640,N_2501);
nor U3024 (N_3024,N_2840,N_2691);
or U3025 (N_3025,N_2366,N_2821);
or U3026 (N_3026,N_2662,N_2555);
nor U3027 (N_3027,N_2573,N_2700);
and U3028 (N_3028,N_2842,N_2683);
or U3029 (N_3029,N_2369,N_2716);
nand U3030 (N_3030,N_2463,N_2894);
or U3031 (N_3031,N_2796,N_2781);
and U3032 (N_3032,N_2865,N_2688);
nor U3033 (N_3033,N_2748,N_2753);
or U3034 (N_3034,N_2970,N_2447);
and U3035 (N_3035,N_2985,N_2306);
nor U3036 (N_3036,N_2563,N_2764);
nand U3037 (N_3037,N_2876,N_2327);
and U3038 (N_3038,N_2790,N_2751);
nand U3039 (N_3039,N_2289,N_2899);
and U3040 (N_3040,N_2643,N_2971);
and U3041 (N_3041,N_2331,N_2257);
or U3042 (N_3042,N_2897,N_2519);
and U3043 (N_3043,N_2852,N_2532);
and U3044 (N_3044,N_2547,N_2775);
and U3045 (N_3045,N_2823,N_2779);
nand U3046 (N_3046,N_2851,N_2301);
and U3047 (N_3047,N_2475,N_2795);
nor U3048 (N_3048,N_2641,N_2690);
and U3049 (N_3049,N_2395,N_2809);
and U3050 (N_3050,N_2658,N_2638);
nor U3051 (N_3051,N_2416,N_2522);
nand U3052 (N_3052,N_2845,N_2835);
and U3053 (N_3053,N_2846,N_2495);
nand U3054 (N_3054,N_2623,N_2564);
nor U3055 (N_3055,N_2998,N_2986);
nand U3056 (N_3056,N_2437,N_2448);
or U3057 (N_3057,N_2304,N_2916);
and U3058 (N_3058,N_2652,N_2667);
nor U3059 (N_3059,N_2379,N_2820);
nand U3060 (N_3060,N_2722,N_2614);
nand U3061 (N_3061,N_2601,N_2740);
and U3062 (N_3062,N_2539,N_2630);
nand U3063 (N_3063,N_2413,N_2520);
and U3064 (N_3064,N_2831,N_2956);
and U3065 (N_3065,N_2405,N_2784);
nand U3066 (N_3066,N_2387,N_2720);
or U3067 (N_3067,N_2441,N_2913);
nand U3068 (N_3068,N_2446,N_2732);
nand U3069 (N_3069,N_2455,N_2414);
or U3070 (N_3070,N_2390,N_2941);
and U3071 (N_3071,N_2468,N_2791);
nand U3072 (N_3072,N_2773,N_2967);
nor U3073 (N_3073,N_2817,N_2517);
nor U3074 (N_3074,N_2856,N_2543);
nor U3075 (N_3075,N_2478,N_2297);
nand U3076 (N_3076,N_2318,N_2933);
or U3077 (N_3077,N_2368,N_2258);
xnor U3078 (N_3078,N_2803,N_2738);
or U3079 (N_3079,N_2848,N_2788);
nand U3080 (N_3080,N_2620,N_2325);
nand U3081 (N_3081,N_2943,N_2878);
and U3082 (N_3082,N_2276,N_2471);
nand U3083 (N_3083,N_2617,N_2747);
and U3084 (N_3084,N_2271,N_2698);
nor U3085 (N_3085,N_2714,N_2587);
nand U3086 (N_3086,N_2359,N_2787);
nor U3087 (N_3087,N_2893,N_2567);
or U3088 (N_3088,N_2919,N_2435);
and U3089 (N_3089,N_2749,N_2905);
and U3090 (N_3090,N_2636,N_2383);
nand U3091 (N_3091,N_2308,N_2671);
or U3092 (N_3092,N_2330,N_2909);
nor U3093 (N_3093,N_2678,N_2511);
nand U3094 (N_3094,N_2651,N_2333);
and U3095 (N_3095,N_2657,N_2419);
and U3096 (N_3096,N_2769,N_2509);
nand U3097 (N_3097,N_2484,N_2812);
or U3098 (N_3098,N_2928,N_2586);
or U3099 (N_3099,N_2499,N_2439);
nor U3100 (N_3100,N_2357,N_2299);
or U3101 (N_3101,N_2844,N_2406);
and U3102 (N_3102,N_2372,N_2332);
or U3103 (N_3103,N_2901,N_2994);
nand U3104 (N_3104,N_2482,N_2252);
nand U3105 (N_3105,N_2502,N_2523);
or U3106 (N_3106,N_2912,N_2950);
and U3107 (N_3107,N_2515,N_2827);
and U3108 (N_3108,N_2403,N_2793);
or U3109 (N_3109,N_2497,N_2378);
nor U3110 (N_3110,N_2409,N_2269);
or U3111 (N_3111,N_2734,N_2622);
or U3112 (N_3112,N_2952,N_2995);
or U3113 (N_3113,N_2774,N_2742);
or U3114 (N_3114,N_2351,N_2572);
nand U3115 (N_3115,N_2559,N_2843);
nor U3116 (N_3116,N_2613,N_2918);
nand U3117 (N_3117,N_2427,N_2672);
nor U3118 (N_3118,N_2602,N_2320);
nand U3119 (N_3119,N_2397,N_2902);
nor U3120 (N_3120,N_2728,N_2668);
nor U3121 (N_3121,N_2705,N_2674);
nor U3122 (N_3122,N_2713,N_2605);
or U3123 (N_3123,N_2615,N_2599);
and U3124 (N_3124,N_2675,N_2806);
and U3125 (N_3125,N_2887,N_2488);
nand U3126 (N_3126,N_2340,N_2485);
nor U3127 (N_3127,N_2417,N_2305);
and U3128 (N_3128,N_2254,N_2489);
nor U3129 (N_3129,N_2661,N_2975);
nor U3130 (N_3130,N_2810,N_2470);
nor U3131 (N_3131,N_2834,N_2343);
nor U3132 (N_3132,N_2972,N_2339);
or U3133 (N_3133,N_2503,N_2365);
nor U3134 (N_3134,N_2531,N_2381);
xnor U3135 (N_3135,N_2477,N_2959);
or U3136 (N_3136,N_2858,N_2380);
or U3137 (N_3137,N_2303,N_2999);
nand U3138 (N_3138,N_2363,N_2644);
nand U3139 (N_3139,N_2634,N_2253);
nand U3140 (N_3140,N_2780,N_2818);
and U3141 (N_3141,N_2256,N_2314);
nor U3142 (N_3142,N_2725,N_2677);
and U3143 (N_3143,N_2294,N_2910);
nand U3144 (N_3144,N_2923,N_2861);
xnor U3145 (N_3145,N_2872,N_2752);
or U3146 (N_3146,N_2792,N_2545);
and U3147 (N_3147,N_2576,N_2839);
nand U3148 (N_3148,N_2693,N_2896);
nand U3149 (N_3149,N_2418,N_2836);
and U3150 (N_3150,N_2371,N_2807);
nor U3151 (N_3151,N_2884,N_2443);
nor U3152 (N_3152,N_2431,N_2938);
or U3153 (N_3153,N_2760,N_2832);
or U3154 (N_3154,N_2541,N_2715);
nand U3155 (N_3155,N_2624,N_2251);
and U3156 (N_3156,N_2370,N_2592);
nor U3157 (N_3157,N_2430,N_2882);
or U3158 (N_3158,N_2954,N_2260);
xnor U3159 (N_3159,N_2566,N_2830);
nor U3160 (N_3160,N_2507,N_2648);
and U3161 (N_3161,N_2857,N_2581);
and U3162 (N_3162,N_2879,N_2346);
and U3163 (N_3163,N_2570,N_2534);
nor U3164 (N_3164,N_2445,N_2467);
and U3165 (N_3165,N_2649,N_2293);
or U3166 (N_3166,N_2440,N_2927);
xor U3167 (N_3167,N_2756,N_2323);
and U3168 (N_3168,N_2645,N_2428);
or U3169 (N_3169,N_2782,N_2266);
and U3170 (N_3170,N_2525,N_2274);
and U3171 (N_3171,N_2450,N_2490);
or U3172 (N_3172,N_2837,N_2518);
or U3173 (N_3173,N_2895,N_2981);
nand U3174 (N_3174,N_2931,N_2707);
nand U3175 (N_3175,N_2578,N_2960);
nand U3176 (N_3176,N_2596,N_2921);
or U3177 (N_3177,N_2527,N_2891);
or U3178 (N_3178,N_2957,N_2802);
xor U3179 (N_3179,N_2361,N_2637);
or U3180 (N_3180,N_2976,N_2337);
nor U3181 (N_3181,N_2528,N_2384);
or U3182 (N_3182,N_2549,N_2655);
nor U3183 (N_3183,N_2873,N_2942);
and U3184 (N_3184,N_2633,N_2530);
or U3185 (N_3185,N_2642,N_2480);
nor U3186 (N_3186,N_2562,N_2375);
and U3187 (N_3187,N_2262,N_2659);
or U3188 (N_3188,N_2483,N_2557);
nand U3189 (N_3189,N_2438,N_2612);
and U3190 (N_3190,N_2295,N_2907);
xor U3191 (N_3191,N_2783,N_2568);
nor U3192 (N_3192,N_2514,N_2492);
nand U3193 (N_3193,N_2750,N_2864);
nor U3194 (N_3194,N_2374,N_2466);
nor U3195 (N_3195,N_2757,N_2561);
and U3196 (N_3196,N_2816,N_2513);
nand U3197 (N_3197,N_2553,N_2699);
and U3198 (N_3198,N_2287,N_2310);
or U3199 (N_3199,N_2506,N_2673);
nand U3200 (N_3200,N_2964,N_2996);
or U3201 (N_3201,N_2974,N_2867);
and U3202 (N_3202,N_2548,N_2611);
nor U3203 (N_3203,N_2465,N_2930);
or U3204 (N_3204,N_2727,N_2741);
nand U3205 (N_3205,N_2983,N_2444);
or U3206 (N_3206,N_2328,N_2604);
nor U3207 (N_3207,N_2647,N_2453);
or U3208 (N_3208,N_2593,N_2469);
nor U3209 (N_3209,N_2393,N_2542);
nor U3210 (N_3210,N_2433,N_2755);
or U3211 (N_3211,N_2735,N_2953);
and U3212 (N_3212,N_2934,N_2311);
and U3213 (N_3213,N_2639,N_2982);
nand U3214 (N_3214,N_2966,N_2595);
and U3215 (N_3215,N_2342,N_2476);
and U3216 (N_3216,N_2424,N_2425);
nand U3217 (N_3217,N_2278,N_2298);
or U3218 (N_3218,N_2399,N_2436);
nor U3219 (N_3219,N_2516,N_2877);
and U3220 (N_3220,N_2389,N_2377);
nand U3221 (N_3221,N_2400,N_2461);
or U3222 (N_3222,N_2263,N_2524);
or U3223 (N_3223,N_2869,N_2504);
nor U3224 (N_3224,N_2550,N_2412);
nor U3225 (N_3225,N_2616,N_2558);
nor U3226 (N_3226,N_2854,N_2676);
or U3227 (N_3227,N_2664,N_2776);
nor U3228 (N_3228,N_2376,N_2656);
or U3229 (N_3229,N_2434,N_2458);
nor U3230 (N_3230,N_2594,N_2733);
nand U3231 (N_3231,N_2556,N_2474);
or U3232 (N_3232,N_2307,N_2900);
nand U3233 (N_3233,N_2432,N_2978);
or U3234 (N_3234,N_2980,N_2984);
and U3235 (N_3235,N_2682,N_2423);
nor U3236 (N_3236,N_2702,N_2706);
and U3237 (N_3237,N_2987,N_2597);
nor U3238 (N_3238,N_2906,N_2917);
nor U3239 (N_3239,N_2336,N_2739);
and U3240 (N_3240,N_2498,N_2388);
or U3241 (N_3241,N_2926,N_2772);
nand U3242 (N_3242,N_2759,N_2798);
nor U3243 (N_3243,N_2335,N_2356);
nand U3244 (N_3244,N_2398,N_2627);
nand U3245 (N_3245,N_2829,N_2822);
and U3246 (N_3246,N_2259,N_2603);
or U3247 (N_3247,N_2540,N_2686);
or U3248 (N_3248,N_2704,N_2701);
nor U3249 (N_3249,N_2746,N_2826);
nand U3250 (N_3250,N_2762,N_2929);
and U3251 (N_3251,N_2600,N_2847);
nand U3252 (N_3252,N_2312,N_2521);
and U3253 (N_3253,N_2533,N_2936);
and U3254 (N_3254,N_2481,N_2815);
and U3255 (N_3255,N_2373,N_2695);
nor U3256 (N_3256,N_2407,N_2408);
nand U3257 (N_3257,N_2394,N_2813);
nand U3258 (N_3258,N_2850,N_2279);
nand U3259 (N_3259,N_2348,N_2537);
and U3260 (N_3260,N_2347,N_2723);
nor U3261 (N_3261,N_2281,N_2708);
nor U3262 (N_3262,N_2512,N_2744);
nor U3263 (N_3263,N_2349,N_2946);
or U3264 (N_3264,N_2681,N_2729);
xor U3265 (N_3265,N_2955,N_2385);
or U3266 (N_3266,N_2606,N_2988);
nor U3267 (N_3267,N_2386,N_2949);
or U3268 (N_3268,N_2653,N_2302);
nor U3269 (N_3269,N_2635,N_2786);
nor U3270 (N_3270,N_2591,N_2529);
nand U3271 (N_3271,N_2932,N_2609);
nor U3272 (N_3272,N_2886,N_2871);
nor U3273 (N_3273,N_2626,N_2940);
nand U3274 (N_3274,N_2284,N_2280);
nor U3275 (N_3275,N_2824,N_2621);
nand U3276 (N_3276,N_2789,N_2666);
or U3277 (N_3277,N_2401,N_2300);
and U3278 (N_3278,N_2863,N_2265);
nand U3279 (N_3279,N_2442,N_2354);
and U3280 (N_3280,N_2317,N_2629);
nand U3281 (N_3281,N_2277,N_2687);
nand U3282 (N_3282,N_2571,N_2487);
and U3283 (N_3283,N_2801,N_2296);
and U3284 (N_3284,N_2853,N_2508);
or U3285 (N_3285,N_2610,N_2316);
nor U3286 (N_3286,N_2631,N_2794);
nor U3287 (N_3287,N_2355,N_2768);
or U3288 (N_3288,N_2703,N_2745);
nand U3289 (N_3289,N_2404,N_2582);
and U3290 (N_3290,N_2804,N_2546);
or U3291 (N_3291,N_2903,N_2282);
xnor U3292 (N_3292,N_2948,N_2579);
nor U3293 (N_3293,N_2460,N_2805);
nand U3294 (N_3294,N_2632,N_2990);
nor U3295 (N_3295,N_2650,N_2669);
and U3296 (N_3296,N_2710,N_2554);
nand U3297 (N_3297,N_2654,N_2585);
nor U3298 (N_3298,N_2754,N_2267);
and U3299 (N_3299,N_2989,N_2991);
and U3300 (N_3300,N_2684,N_2680);
and U3301 (N_3301,N_2329,N_2565);
nor U3302 (N_3302,N_2665,N_2574);
nand U3303 (N_3303,N_2914,N_2904);
or U3304 (N_3304,N_2721,N_2456);
and U3305 (N_3305,N_2997,N_2945);
nor U3306 (N_3306,N_2717,N_2493);
or U3307 (N_3307,N_2291,N_2993);
nand U3308 (N_3308,N_2410,N_2924);
and U3309 (N_3309,N_2799,N_2771);
or U3310 (N_3310,N_2580,N_2689);
and U3311 (N_3311,N_2965,N_2968);
or U3312 (N_3312,N_2855,N_2309);
nor U3313 (N_3313,N_2345,N_2646);
nor U3314 (N_3314,N_2885,N_2743);
nand U3315 (N_3315,N_2551,N_2973);
nor U3316 (N_3316,N_2961,N_2421);
or U3317 (N_3317,N_2628,N_2736);
and U3318 (N_3318,N_2761,N_2319);
or U3319 (N_3319,N_2286,N_2618);
and U3320 (N_3320,N_2778,N_2712);
or U3321 (N_3321,N_2583,N_2911);
nor U3322 (N_3322,N_2326,N_2429);
nand U3323 (N_3323,N_2577,N_2880);
nor U3324 (N_3324,N_2607,N_2767);
nor U3325 (N_3325,N_2449,N_2892);
and U3326 (N_3326,N_2939,N_2890);
or U3327 (N_3327,N_2353,N_2526);
xnor U3328 (N_3328,N_2958,N_2367);
and U3329 (N_3329,N_2544,N_2692);
nor U3330 (N_3330,N_2575,N_2819);
or U3331 (N_3331,N_2426,N_2770);
nand U3332 (N_3332,N_2536,N_2889);
nand U3333 (N_3333,N_2874,N_2737);
or U3334 (N_3334,N_2264,N_2288);
nand U3335 (N_3335,N_2250,N_2833);
and U3336 (N_3336,N_2491,N_2875);
nand U3337 (N_3337,N_2718,N_2962);
or U3338 (N_3338,N_2709,N_2505);
and U3339 (N_3339,N_2270,N_2590);
and U3340 (N_3340,N_2494,N_2937);
xor U3341 (N_3341,N_2694,N_2992);
or U3342 (N_3342,N_2479,N_2464);
and U3343 (N_3343,N_2552,N_2451);
nor U3344 (N_3344,N_2261,N_2538);
nand U3345 (N_3345,N_2352,N_2350);
and U3346 (N_3346,N_2462,N_2292);
nand U3347 (N_3347,N_2696,N_2944);
nand U3348 (N_3348,N_2963,N_2459);
or U3349 (N_3349,N_2454,N_2838);
nor U3350 (N_3350,N_2411,N_2979);
nor U3351 (N_3351,N_2726,N_2898);
or U3352 (N_3352,N_2422,N_2275);
nor U3353 (N_3353,N_2977,N_2496);
or U3354 (N_3354,N_2588,N_2324);
and U3355 (N_3355,N_2360,N_2797);
or U3356 (N_3356,N_2322,N_2619);
nand U3357 (N_3357,N_2859,N_2663);
nand U3358 (N_3358,N_2358,N_2951);
nand U3359 (N_3359,N_2719,N_2321);
nand U3360 (N_3360,N_2598,N_2758);
and U3361 (N_3361,N_2711,N_2763);
and U3362 (N_3362,N_2849,N_2785);
nand U3363 (N_3363,N_2420,N_2396);
nor U3364 (N_3364,N_2391,N_2486);
nand U3365 (N_3365,N_2935,N_2268);
or U3366 (N_3366,N_2800,N_2608);
or U3367 (N_3367,N_2452,N_2730);
or U3368 (N_3368,N_2814,N_2670);
or U3369 (N_3369,N_2290,N_2868);
and U3370 (N_3370,N_2535,N_2272);
or U3371 (N_3371,N_2313,N_2765);
xor U3372 (N_3372,N_2392,N_2589);
xnor U3373 (N_3373,N_2362,N_2255);
nand U3374 (N_3374,N_2584,N_2334);
nor U3375 (N_3375,N_2923,N_2853);
nand U3376 (N_3376,N_2863,N_2887);
nand U3377 (N_3377,N_2969,N_2833);
nor U3378 (N_3378,N_2551,N_2501);
and U3379 (N_3379,N_2724,N_2558);
and U3380 (N_3380,N_2717,N_2845);
nand U3381 (N_3381,N_2879,N_2327);
xnor U3382 (N_3382,N_2994,N_2887);
xor U3383 (N_3383,N_2785,N_2807);
nand U3384 (N_3384,N_2954,N_2474);
nor U3385 (N_3385,N_2600,N_2263);
and U3386 (N_3386,N_2939,N_2897);
nand U3387 (N_3387,N_2316,N_2293);
nand U3388 (N_3388,N_2989,N_2488);
nor U3389 (N_3389,N_2491,N_2852);
nor U3390 (N_3390,N_2592,N_2303);
nand U3391 (N_3391,N_2881,N_2293);
nor U3392 (N_3392,N_2423,N_2945);
nor U3393 (N_3393,N_2983,N_2922);
nor U3394 (N_3394,N_2929,N_2973);
nand U3395 (N_3395,N_2948,N_2842);
or U3396 (N_3396,N_2894,N_2356);
or U3397 (N_3397,N_2725,N_2546);
or U3398 (N_3398,N_2288,N_2986);
nand U3399 (N_3399,N_2495,N_2880);
nor U3400 (N_3400,N_2629,N_2568);
and U3401 (N_3401,N_2863,N_2945);
and U3402 (N_3402,N_2340,N_2772);
and U3403 (N_3403,N_2878,N_2811);
nor U3404 (N_3404,N_2764,N_2365);
and U3405 (N_3405,N_2502,N_2915);
and U3406 (N_3406,N_2435,N_2426);
nor U3407 (N_3407,N_2535,N_2496);
and U3408 (N_3408,N_2925,N_2857);
and U3409 (N_3409,N_2546,N_2398);
or U3410 (N_3410,N_2250,N_2557);
nor U3411 (N_3411,N_2299,N_2318);
or U3412 (N_3412,N_2761,N_2437);
nand U3413 (N_3413,N_2699,N_2331);
nand U3414 (N_3414,N_2267,N_2575);
or U3415 (N_3415,N_2767,N_2649);
and U3416 (N_3416,N_2734,N_2392);
or U3417 (N_3417,N_2599,N_2449);
xor U3418 (N_3418,N_2462,N_2575);
or U3419 (N_3419,N_2680,N_2292);
nor U3420 (N_3420,N_2519,N_2324);
nand U3421 (N_3421,N_2487,N_2486);
nor U3422 (N_3422,N_2629,N_2626);
or U3423 (N_3423,N_2512,N_2506);
nor U3424 (N_3424,N_2716,N_2827);
nor U3425 (N_3425,N_2687,N_2344);
nor U3426 (N_3426,N_2875,N_2425);
or U3427 (N_3427,N_2952,N_2321);
nor U3428 (N_3428,N_2839,N_2824);
and U3429 (N_3429,N_2399,N_2999);
nor U3430 (N_3430,N_2741,N_2323);
or U3431 (N_3431,N_2362,N_2293);
nand U3432 (N_3432,N_2343,N_2942);
nor U3433 (N_3433,N_2380,N_2831);
nand U3434 (N_3434,N_2797,N_2665);
and U3435 (N_3435,N_2385,N_2505);
and U3436 (N_3436,N_2963,N_2812);
nand U3437 (N_3437,N_2746,N_2742);
or U3438 (N_3438,N_2748,N_2581);
and U3439 (N_3439,N_2556,N_2276);
and U3440 (N_3440,N_2447,N_2357);
nor U3441 (N_3441,N_2734,N_2821);
nand U3442 (N_3442,N_2791,N_2890);
nand U3443 (N_3443,N_2945,N_2695);
and U3444 (N_3444,N_2479,N_2345);
and U3445 (N_3445,N_2704,N_2659);
or U3446 (N_3446,N_2606,N_2299);
or U3447 (N_3447,N_2493,N_2778);
or U3448 (N_3448,N_2561,N_2267);
nor U3449 (N_3449,N_2371,N_2789);
nand U3450 (N_3450,N_2959,N_2982);
and U3451 (N_3451,N_2890,N_2902);
nand U3452 (N_3452,N_2335,N_2483);
or U3453 (N_3453,N_2509,N_2627);
or U3454 (N_3454,N_2408,N_2838);
xor U3455 (N_3455,N_2764,N_2879);
nor U3456 (N_3456,N_2660,N_2296);
and U3457 (N_3457,N_2868,N_2943);
and U3458 (N_3458,N_2975,N_2422);
or U3459 (N_3459,N_2400,N_2469);
nand U3460 (N_3460,N_2846,N_2418);
nor U3461 (N_3461,N_2584,N_2682);
nand U3462 (N_3462,N_2874,N_2518);
nand U3463 (N_3463,N_2329,N_2417);
nand U3464 (N_3464,N_2573,N_2842);
or U3465 (N_3465,N_2789,N_2762);
and U3466 (N_3466,N_2766,N_2840);
or U3467 (N_3467,N_2502,N_2653);
nand U3468 (N_3468,N_2351,N_2483);
nand U3469 (N_3469,N_2504,N_2518);
or U3470 (N_3470,N_2455,N_2418);
nand U3471 (N_3471,N_2304,N_2293);
nand U3472 (N_3472,N_2934,N_2403);
or U3473 (N_3473,N_2950,N_2621);
nor U3474 (N_3474,N_2809,N_2337);
or U3475 (N_3475,N_2372,N_2545);
nor U3476 (N_3476,N_2990,N_2647);
nand U3477 (N_3477,N_2767,N_2987);
or U3478 (N_3478,N_2590,N_2523);
and U3479 (N_3479,N_2378,N_2648);
and U3480 (N_3480,N_2464,N_2393);
nor U3481 (N_3481,N_2404,N_2853);
or U3482 (N_3482,N_2622,N_2286);
nor U3483 (N_3483,N_2796,N_2335);
and U3484 (N_3484,N_2385,N_2535);
or U3485 (N_3485,N_2778,N_2706);
nand U3486 (N_3486,N_2338,N_2820);
and U3487 (N_3487,N_2921,N_2266);
nor U3488 (N_3488,N_2545,N_2258);
and U3489 (N_3489,N_2427,N_2770);
nor U3490 (N_3490,N_2925,N_2738);
or U3491 (N_3491,N_2569,N_2397);
and U3492 (N_3492,N_2629,N_2394);
nor U3493 (N_3493,N_2595,N_2786);
and U3494 (N_3494,N_2601,N_2258);
and U3495 (N_3495,N_2520,N_2344);
nand U3496 (N_3496,N_2285,N_2396);
and U3497 (N_3497,N_2852,N_2474);
and U3498 (N_3498,N_2366,N_2454);
and U3499 (N_3499,N_2592,N_2669);
nor U3500 (N_3500,N_2974,N_2958);
and U3501 (N_3501,N_2518,N_2369);
nand U3502 (N_3502,N_2344,N_2992);
nor U3503 (N_3503,N_2831,N_2737);
nor U3504 (N_3504,N_2910,N_2984);
and U3505 (N_3505,N_2747,N_2293);
or U3506 (N_3506,N_2866,N_2615);
or U3507 (N_3507,N_2414,N_2953);
and U3508 (N_3508,N_2264,N_2801);
nor U3509 (N_3509,N_2303,N_2639);
and U3510 (N_3510,N_2467,N_2565);
or U3511 (N_3511,N_2447,N_2367);
nand U3512 (N_3512,N_2807,N_2753);
or U3513 (N_3513,N_2630,N_2948);
or U3514 (N_3514,N_2388,N_2480);
nor U3515 (N_3515,N_2511,N_2858);
nor U3516 (N_3516,N_2255,N_2366);
and U3517 (N_3517,N_2515,N_2718);
or U3518 (N_3518,N_2503,N_2808);
or U3519 (N_3519,N_2313,N_2376);
nor U3520 (N_3520,N_2755,N_2903);
nor U3521 (N_3521,N_2341,N_2801);
or U3522 (N_3522,N_2902,N_2479);
nor U3523 (N_3523,N_2449,N_2299);
nand U3524 (N_3524,N_2998,N_2881);
xor U3525 (N_3525,N_2536,N_2376);
nor U3526 (N_3526,N_2408,N_2621);
and U3527 (N_3527,N_2967,N_2335);
or U3528 (N_3528,N_2386,N_2983);
nor U3529 (N_3529,N_2501,N_2350);
and U3530 (N_3530,N_2772,N_2835);
xor U3531 (N_3531,N_2303,N_2426);
nor U3532 (N_3532,N_2287,N_2609);
nand U3533 (N_3533,N_2433,N_2863);
and U3534 (N_3534,N_2533,N_2445);
or U3535 (N_3535,N_2873,N_2856);
and U3536 (N_3536,N_2738,N_2455);
nor U3537 (N_3537,N_2366,N_2705);
nor U3538 (N_3538,N_2964,N_2310);
and U3539 (N_3539,N_2459,N_2657);
nand U3540 (N_3540,N_2936,N_2518);
and U3541 (N_3541,N_2516,N_2340);
nand U3542 (N_3542,N_2378,N_2721);
nor U3543 (N_3543,N_2410,N_2395);
or U3544 (N_3544,N_2814,N_2349);
nor U3545 (N_3545,N_2657,N_2546);
nor U3546 (N_3546,N_2511,N_2549);
nor U3547 (N_3547,N_2378,N_2772);
nor U3548 (N_3548,N_2596,N_2413);
or U3549 (N_3549,N_2537,N_2417);
and U3550 (N_3550,N_2549,N_2697);
or U3551 (N_3551,N_2786,N_2412);
or U3552 (N_3552,N_2310,N_2405);
nand U3553 (N_3553,N_2268,N_2561);
and U3554 (N_3554,N_2792,N_2964);
and U3555 (N_3555,N_2857,N_2773);
nor U3556 (N_3556,N_2502,N_2591);
nand U3557 (N_3557,N_2738,N_2620);
nand U3558 (N_3558,N_2492,N_2489);
and U3559 (N_3559,N_2853,N_2735);
or U3560 (N_3560,N_2922,N_2513);
nor U3561 (N_3561,N_2357,N_2378);
nand U3562 (N_3562,N_2830,N_2376);
nand U3563 (N_3563,N_2754,N_2923);
nand U3564 (N_3564,N_2796,N_2669);
and U3565 (N_3565,N_2777,N_2475);
or U3566 (N_3566,N_2813,N_2908);
nor U3567 (N_3567,N_2598,N_2634);
or U3568 (N_3568,N_2277,N_2498);
or U3569 (N_3569,N_2895,N_2871);
or U3570 (N_3570,N_2339,N_2781);
nor U3571 (N_3571,N_2688,N_2554);
nor U3572 (N_3572,N_2908,N_2712);
nor U3573 (N_3573,N_2309,N_2919);
nor U3574 (N_3574,N_2827,N_2751);
nand U3575 (N_3575,N_2449,N_2323);
or U3576 (N_3576,N_2525,N_2430);
xnor U3577 (N_3577,N_2473,N_2940);
nand U3578 (N_3578,N_2440,N_2578);
nor U3579 (N_3579,N_2904,N_2300);
and U3580 (N_3580,N_2707,N_2981);
nor U3581 (N_3581,N_2866,N_2380);
nand U3582 (N_3582,N_2381,N_2577);
nor U3583 (N_3583,N_2436,N_2276);
or U3584 (N_3584,N_2751,N_2894);
nor U3585 (N_3585,N_2713,N_2334);
nand U3586 (N_3586,N_2547,N_2372);
nand U3587 (N_3587,N_2825,N_2817);
and U3588 (N_3588,N_2338,N_2939);
or U3589 (N_3589,N_2546,N_2676);
xor U3590 (N_3590,N_2478,N_2271);
or U3591 (N_3591,N_2804,N_2664);
nand U3592 (N_3592,N_2487,N_2943);
nand U3593 (N_3593,N_2468,N_2703);
nand U3594 (N_3594,N_2318,N_2273);
nor U3595 (N_3595,N_2333,N_2836);
or U3596 (N_3596,N_2824,N_2740);
or U3597 (N_3597,N_2528,N_2622);
nor U3598 (N_3598,N_2320,N_2537);
xnor U3599 (N_3599,N_2441,N_2303);
or U3600 (N_3600,N_2419,N_2969);
nand U3601 (N_3601,N_2702,N_2866);
and U3602 (N_3602,N_2908,N_2816);
xor U3603 (N_3603,N_2769,N_2566);
or U3604 (N_3604,N_2445,N_2700);
and U3605 (N_3605,N_2799,N_2923);
nand U3606 (N_3606,N_2391,N_2675);
xor U3607 (N_3607,N_2401,N_2526);
and U3608 (N_3608,N_2572,N_2808);
nor U3609 (N_3609,N_2362,N_2764);
xor U3610 (N_3610,N_2396,N_2963);
and U3611 (N_3611,N_2852,N_2686);
nor U3612 (N_3612,N_2554,N_2374);
or U3613 (N_3613,N_2567,N_2328);
nand U3614 (N_3614,N_2344,N_2954);
and U3615 (N_3615,N_2986,N_2962);
nor U3616 (N_3616,N_2963,N_2888);
or U3617 (N_3617,N_2593,N_2743);
nand U3618 (N_3618,N_2746,N_2939);
nand U3619 (N_3619,N_2632,N_2285);
xnor U3620 (N_3620,N_2753,N_2367);
and U3621 (N_3621,N_2498,N_2681);
or U3622 (N_3622,N_2885,N_2883);
nand U3623 (N_3623,N_2819,N_2481);
nor U3624 (N_3624,N_2756,N_2737);
nor U3625 (N_3625,N_2458,N_2828);
nor U3626 (N_3626,N_2884,N_2848);
nand U3627 (N_3627,N_2648,N_2820);
or U3628 (N_3628,N_2756,N_2874);
nand U3629 (N_3629,N_2712,N_2258);
nand U3630 (N_3630,N_2722,N_2877);
or U3631 (N_3631,N_2279,N_2518);
nor U3632 (N_3632,N_2929,N_2362);
and U3633 (N_3633,N_2495,N_2732);
nor U3634 (N_3634,N_2874,N_2971);
and U3635 (N_3635,N_2979,N_2522);
or U3636 (N_3636,N_2872,N_2472);
nor U3637 (N_3637,N_2330,N_2523);
and U3638 (N_3638,N_2405,N_2823);
nand U3639 (N_3639,N_2525,N_2317);
or U3640 (N_3640,N_2266,N_2877);
nor U3641 (N_3641,N_2890,N_2542);
nand U3642 (N_3642,N_2510,N_2840);
xnor U3643 (N_3643,N_2871,N_2499);
or U3644 (N_3644,N_2866,N_2677);
nor U3645 (N_3645,N_2721,N_2391);
or U3646 (N_3646,N_2332,N_2864);
nor U3647 (N_3647,N_2989,N_2515);
nand U3648 (N_3648,N_2403,N_2559);
and U3649 (N_3649,N_2558,N_2283);
and U3650 (N_3650,N_2359,N_2283);
nor U3651 (N_3651,N_2526,N_2537);
nand U3652 (N_3652,N_2489,N_2817);
xnor U3653 (N_3653,N_2922,N_2658);
and U3654 (N_3654,N_2871,N_2384);
or U3655 (N_3655,N_2909,N_2960);
or U3656 (N_3656,N_2808,N_2694);
or U3657 (N_3657,N_2881,N_2856);
or U3658 (N_3658,N_2443,N_2348);
nor U3659 (N_3659,N_2966,N_2933);
nand U3660 (N_3660,N_2271,N_2568);
nor U3661 (N_3661,N_2374,N_2445);
nand U3662 (N_3662,N_2381,N_2647);
or U3663 (N_3663,N_2804,N_2448);
nand U3664 (N_3664,N_2934,N_2985);
nor U3665 (N_3665,N_2665,N_2930);
and U3666 (N_3666,N_2488,N_2656);
and U3667 (N_3667,N_2784,N_2825);
nor U3668 (N_3668,N_2612,N_2624);
and U3669 (N_3669,N_2493,N_2613);
nor U3670 (N_3670,N_2541,N_2633);
nor U3671 (N_3671,N_2454,N_2773);
nor U3672 (N_3672,N_2371,N_2741);
and U3673 (N_3673,N_2705,N_2421);
or U3674 (N_3674,N_2279,N_2507);
or U3675 (N_3675,N_2296,N_2422);
nand U3676 (N_3676,N_2673,N_2642);
nand U3677 (N_3677,N_2896,N_2561);
nor U3678 (N_3678,N_2521,N_2572);
and U3679 (N_3679,N_2587,N_2623);
xnor U3680 (N_3680,N_2762,N_2654);
nand U3681 (N_3681,N_2573,N_2463);
nor U3682 (N_3682,N_2880,N_2945);
and U3683 (N_3683,N_2354,N_2329);
or U3684 (N_3684,N_2837,N_2636);
xor U3685 (N_3685,N_2281,N_2397);
or U3686 (N_3686,N_2575,N_2929);
or U3687 (N_3687,N_2756,N_2898);
nor U3688 (N_3688,N_2710,N_2794);
nor U3689 (N_3689,N_2968,N_2489);
nor U3690 (N_3690,N_2511,N_2470);
nor U3691 (N_3691,N_2282,N_2317);
or U3692 (N_3692,N_2807,N_2630);
and U3693 (N_3693,N_2490,N_2714);
or U3694 (N_3694,N_2485,N_2751);
nor U3695 (N_3695,N_2946,N_2465);
nor U3696 (N_3696,N_2746,N_2719);
nand U3697 (N_3697,N_2953,N_2995);
and U3698 (N_3698,N_2392,N_2744);
nor U3699 (N_3699,N_2463,N_2354);
nor U3700 (N_3700,N_2925,N_2434);
nand U3701 (N_3701,N_2607,N_2419);
and U3702 (N_3702,N_2419,N_2253);
nor U3703 (N_3703,N_2276,N_2708);
or U3704 (N_3704,N_2328,N_2989);
nand U3705 (N_3705,N_2419,N_2988);
or U3706 (N_3706,N_2912,N_2828);
nor U3707 (N_3707,N_2936,N_2590);
nand U3708 (N_3708,N_2853,N_2301);
nor U3709 (N_3709,N_2681,N_2906);
or U3710 (N_3710,N_2882,N_2907);
nand U3711 (N_3711,N_2484,N_2323);
and U3712 (N_3712,N_2953,N_2944);
nor U3713 (N_3713,N_2490,N_2677);
nor U3714 (N_3714,N_2670,N_2750);
and U3715 (N_3715,N_2990,N_2505);
xor U3716 (N_3716,N_2749,N_2570);
nor U3717 (N_3717,N_2431,N_2364);
nand U3718 (N_3718,N_2929,N_2999);
nand U3719 (N_3719,N_2671,N_2323);
and U3720 (N_3720,N_2561,N_2395);
nor U3721 (N_3721,N_2293,N_2757);
or U3722 (N_3722,N_2570,N_2304);
or U3723 (N_3723,N_2808,N_2525);
or U3724 (N_3724,N_2852,N_2902);
or U3725 (N_3725,N_2404,N_2852);
and U3726 (N_3726,N_2871,N_2423);
nor U3727 (N_3727,N_2595,N_2521);
and U3728 (N_3728,N_2421,N_2947);
nand U3729 (N_3729,N_2771,N_2948);
nand U3730 (N_3730,N_2322,N_2372);
xnor U3731 (N_3731,N_2825,N_2632);
nor U3732 (N_3732,N_2384,N_2731);
and U3733 (N_3733,N_2347,N_2317);
nand U3734 (N_3734,N_2610,N_2663);
nor U3735 (N_3735,N_2873,N_2643);
nand U3736 (N_3736,N_2759,N_2881);
nand U3737 (N_3737,N_2551,N_2450);
nand U3738 (N_3738,N_2761,N_2635);
or U3739 (N_3739,N_2760,N_2999);
nor U3740 (N_3740,N_2463,N_2263);
nor U3741 (N_3741,N_2387,N_2834);
and U3742 (N_3742,N_2316,N_2893);
nand U3743 (N_3743,N_2588,N_2925);
or U3744 (N_3744,N_2345,N_2961);
and U3745 (N_3745,N_2812,N_2385);
or U3746 (N_3746,N_2341,N_2394);
or U3747 (N_3747,N_2876,N_2309);
nor U3748 (N_3748,N_2318,N_2295);
xor U3749 (N_3749,N_2428,N_2967);
or U3750 (N_3750,N_3451,N_3233);
or U3751 (N_3751,N_3427,N_3621);
or U3752 (N_3752,N_3551,N_3381);
or U3753 (N_3753,N_3498,N_3740);
and U3754 (N_3754,N_3473,N_3076);
or U3755 (N_3755,N_3595,N_3619);
nand U3756 (N_3756,N_3351,N_3736);
or U3757 (N_3757,N_3541,N_3463);
or U3758 (N_3758,N_3548,N_3386);
or U3759 (N_3759,N_3031,N_3558);
and U3760 (N_3760,N_3467,N_3057);
and U3761 (N_3761,N_3734,N_3329);
or U3762 (N_3762,N_3020,N_3586);
nand U3763 (N_3763,N_3108,N_3030);
nand U3764 (N_3764,N_3468,N_3025);
nand U3765 (N_3765,N_3681,N_3490);
nand U3766 (N_3766,N_3379,N_3338);
and U3767 (N_3767,N_3477,N_3152);
nand U3768 (N_3768,N_3245,N_3589);
nand U3769 (N_3769,N_3109,N_3482);
nand U3770 (N_3770,N_3633,N_3056);
nand U3771 (N_3771,N_3142,N_3275);
or U3772 (N_3772,N_3083,N_3287);
or U3773 (N_3773,N_3531,N_3724);
and U3774 (N_3774,N_3378,N_3235);
xor U3775 (N_3775,N_3702,N_3113);
nand U3776 (N_3776,N_3550,N_3018);
xor U3777 (N_3777,N_3085,N_3708);
and U3778 (N_3778,N_3514,N_3191);
or U3779 (N_3779,N_3010,N_3087);
or U3780 (N_3780,N_3368,N_3657);
nand U3781 (N_3781,N_3178,N_3471);
or U3782 (N_3782,N_3455,N_3073);
and U3783 (N_3783,N_3183,N_3453);
or U3784 (N_3784,N_3003,N_3642);
nand U3785 (N_3785,N_3554,N_3487);
nand U3786 (N_3786,N_3277,N_3655);
nor U3787 (N_3787,N_3549,N_3699);
nand U3788 (N_3788,N_3236,N_3685);
nand U3789 (N_3789,N_3501,N_3315);
nand U3790 (N_3790,N_3211,N_3229);
and U3791 (N_3791,N_3251,N_3643);
and U3792 (N_3792,N_3735,N_3268);
or U3793 (N_3793,N_3524,N_3330);
and U3794 (N_3794,N_3074,N_3475);
and U3795 (N_3795,N_3224,N_3278);
and U3796 (N_3796,N_3500,N_3441);
or U3797 (N_3797,N_3340,N_3510);
nand U3798 (N_3798,N_3372,N_3544);
and U3799 (N_3799,N_3469,N_3300);
and U3800 (N_3800,N_3144,N_3119);
and U3801 (N_3801,N_3247,N_3506);
nor U3802 (N_3802,N_3127,N_3201);
nor U3803 (N_3803,N_3611,N_3215);
xnor U3804 (N_3804,N_3722,N_3089);
and U3805 (N_3805,N_3060,N_3519);
nor U3806 (N_3806,N_3175,N_3373);
nand U3807 (N_3807,N_3632,N_3527);
and U3808 (N_3808,N_3522,N_3069);
or U3809 (N_3809,N_3009,N_3384);
nor U3810 (N_3810,N_3555,N_3179);
nor U3811 (N_3811,N_3623,N_3682);
xnor U3812 (N_3812,N_3440,N_3709);
and U3813 (N_3813,N_3326,N_3604);
or U3814 (N_3814,N_3557,N_3364);
or U3815 (N_3815,N_3129,N_3537);
or U3816 (N_3816,N_3303,N_3237);
and U3817 (N_3817,N_3147,N_3645);
and U3818 (N_3818,N_3322,N_3264);
or U3819 (N_3819,N_3267,N_3584);
or U3820 (N_3820,N_3285,N_3148);
nand U3821 (N_3821,N_3374,N_3513);
or U3822 (N_3822,N_3156,N_3663);
nor U3823 (N_3823,N_3099,N_3265);
and U3824 (N_3824,N_3496,N_3637);
and U3825 (N_3825,N_3096,N_3166);
nand U3826 (N_3826,N_3036,N_3518);
or U3827 (N_3827,N_3594,N_3483);
nand U3828 (N_3828,N_3197,N_3344);
nor U3829 (N_3829,N_3098,N_3260);
and U3830 (N_3830,N_3239,N_3610);
nand U3831 (N_3831,N_3337,N_3577);
nand U3832 (N_3832,N_3700,N_3556);
nand U3833 (N_3833,N_3291,N_3058);
nor U3834 (N_3834,N_3054,N_3669);
nor U3835 (N_3835,N_3647,N_3240);
or U3836 (N_3836,N_3488,N_3667);
or U3837 (N_3837,N_3213,N_3413);
or U3838 (N_3838,N_3732,N_3746);
or U3839 (N_3839,N_3184,N_3234);
nand U3840 (N_3840,N_3005,N_3635);
and U3841 (N_3841,N_3401,N_3420);
and U3842 (N_3842,N_3695,N_3404);
or U3843 (N_3843,N_3186,N_3082);
nor U3844 (N_3844,N_3327,N_3043);
nor U3845 (N_3845,N_3684,N_3218);
or U3846 (N_3846,N_3116,N_3172);
and U3847 (N_3847,N_3047,N_3388);
and U3848 (N_3848,N_3414,N_3159);
and U3849 (N_3849,N_3542,N_3192);
or U3850 (N_3850,N_3336,N_3041);
nand U3851 (N_3851,N_3103,N_3707);
or U3852 (N_3852,N_3567,N_3389);
or U3853 (N_3853,N_3301,N_3081);
nor U3854 (N_3854,N_3442,N_3161);
or U3855 (N_3855,N_3155,N_3366);
or U3856 (N_3856,N_3072,N_3320);
and U3857 (N_3857,N_3662,N_3710);
nand U3858 (N_3858,N_3546,N_3097);
and U3859 (N_3859,N_3661,N_3507);
or U3860 (N_3860,N_3634,N_3450);
nor U3861 (N_3861,N_3295,N_3261);
or U3862 (N_3862,N_3292,N_3288);
nand U3863 (N_3863,N_3680,N_3607);
xor U3864 (N_3864,N_3508,N_3377);
nor U3865 (N_3865,N_3590,N_3572);
or U3866 (N_3866,N_3703,N_3525);
and U3867 (N_3867,N_3733,N_3310);
and U3868 (N_3868,N_3023,N_3484);
xnor U3869 (N_3869,N_3398,N_3445);
or U3870 (N_3870,N_3297,N_3137);
nand U3871 (N_3871,N_3094,N_3606);
and U3872 (N_3872,N_3321,N_3491);
and U3873 (N_3873,N_3687,N_3438);
nand U3874 (N_3874,N_3363,N_3408);
nor U3875 (N_3875,N_3112,N_3578);
nand U3876 (N_3876,N_3013,N_3139);
or U3877 (N_3877,N_3253,N_3199);
nand U3878 (N_3878,N_3658,N_3106);
or U3879 (N_3879,N_3561,N_3162);
nand U3880 (N_3880,N_3512,N_3101);
xnor U3881 (N_3881,N_3715,N_3362);
or U3882 (N_3882,N_3086,N_3304);
nor U3883 (N_3883,N_3696,N_3560);
or U3884 (N_3884,N_3638,N_3651);
nor U3885 (N_3885,N_3169,N_3311);
nand U3886 (N_3886,N_3221,N_3002);
and U3887 (N_3887,N_3314,N_3676);
and U3888 (N_3888,N_3480,N_3367);
nor U3889 (N_3889,N_3472,N_3180);
nand U3890 (N_3890,N_3656,N_3004);
and U3891 (N_3891,N_3104,N_3185);
nor U3892 (N_3892,N_3448,N_3489);
nand U3893 (N_3893,N_3418,N_3318);
nor U3894 (N_3894,N_3145,N_3565);
or U3895 (N_3895,N_3628,N_3284);
or U3896 (N_3896,N_3063,N_3254);
xnor U3897 (N_3897,N_3032,N_3380);
or U3898 (N_3898,N_3517,N_3189);
nand U3899 (N_3899,N_3605,N_3259);
and U3900 (N_3900,N_3202,N_3037);
xor U3901 (N_3901,N_3255,N_3190);
nor U3902 (N_3902,N_3598,N_3402);
nor U3903 (N_3903,N_3346,N_3207);
or U3904 (N_3904,N_3552,N_3280);
nor U3905 (N_3905,N_3121,N_3017);
or U3906 (N_3906,N_3353,N_3624);
and U3907 (N_3907,N_3744,N_3614);
nand U3908 (N_3908,N_3133,N_3677);
nand U3909 (N_3909,N_3585,N_3516);
nand U3910 (N_3910,N_3026,N_3006);
nor U3911 (N_3911,N_3485,N_3217);
and U3912 (N_3912,N_3028,N_3620);
and U3913 (N_3913,N_3686,N_3443);
nand U3914 (N_3914,N_3130,N_3205);
or U3915 (N_3915,N_3067,N_3460);
and U3916 (N_3916,N_3212,N_3547);
and U3917 (N_3917,N_3583,N_3536);
or U3918 (N_3918,N_3171,N_3726);
xnor U3919 (N_3919,N_3563,N_3066);
nand U3920 (N_3920,N_3694,N_3078);
nor U3921 (N_3921,N_3208,N_3738);
xor U3922 (N_3922,N_3256,N_3281);
or U3923 (N_3923,N_3163,N_3742);
nor U3924 (N_3924,N_3357,N_3027);
nor U3925 (N_3925,N_3262,N_3024);
or U3926 (N_3926,N_3350,N_3574);
and U3927 (N_3927,N_3048,N_3530);
nand U3928 (N_3928,N_3126,N_3434);
or U3929 (N_3929,N_3706,N_3494);
and U3930 (N_3930,N_3629,N_3135);
or U3931 (N_3931,N_3691,N_3195);
nor U3932 (N_3932,N_3231,N_3328);
and U3933 (N_3933,N_3335,N_3409);
nor U3934 (N_3934,N_3117,N_3627);
and U3935 (N_3935,N_3421,N_3334);
or U3936 (N_3936,N_3021,N_3071);
or U3937 (N_3937,N_3204,N_3428);
or U3938 (N_3938,N_3114,N_3059);
and U3939 (N_3939,N_3739,N_3219);
or U3940 (N_3940,N_3419,N_3406);
and U3941 (N_3941,N_3743,N_3602);
nor U3942 (N_3942,N_3616,N_3214);
nand U3943 (N_3943,N_3248,N_3729);
and U3944 (N_3944,N_3539,N_3433);
and U3945 (N_3945,N_3431,N_3052);
and U3946 (N_3946,N_3196,N_3592);
and U3947 (N_3947,N_3405,N_3216);
nor U3948 (N_3948,N_3014,N_3065);
nand U3949 (N_3949,N_3690,N_3257);
and U3950 (N_3950,N_3515,N_3478);
nand U3951 (N_3951,N_3150,N_3307);
nand U3952 (N_3952,N_3609,N_3603);
or U3953 (N_3953,N_3348,N_3022);
and U3954 (N_3954,N_3430,N_3631);
or U3955 (N_3955,N_3587,N_3200);
nand U3956 (N_3956,N_3151,N_3429);
or U3957 (N_3957,N_3193,N_3535);
or U3958 (N_3958,N_3416,N_3134);
nor U3959 (N_3959,N_3387,N_3673);
nor U3960 (N_3960,N_3283,N_3276);
nor U3961 (N_3961,N_3395,N_3597);
or U3962 (N_3962,N_3678,N_3458);
and U3963 (N_3963,N_3170,N_3062);
nor U3964 (N_3964,N_3138,N_3679);
and U3965 (N_3965,N_3035,N_3149);
or U3966 (N_3966,N_3039,N_3741);
and U3967 (N_3967,N_3258,N_3465);
nor U3968 (N_3968,N_3720,N_3222);
nor U3969 (N_3969,N_3444,N_3349);
nand U3970 (N_3970,N_3748,N_3615);
or U3971 (N_3971,N_3410,N_3432);
or U3972 (N_3972,N_3051,N_3061);
nand U3973 (N_3973,N_3447,N_3683);
nor U3974 (N_3974,N_3644,N_3626);
or U3975 (N_3975,N_3529,N_3566);
or U3976 (N_3976,N_3641,N_3526);
and U3977 (N_3977,N_3665,N_3157);
nand U3978 (N_3978,N_3470,N_3012);
and U3979 (N_3979,N_3077,N_3294);
or U3980 (N_3980,N_3618,N_3481);
or U3981 (N_3981,N_3625,N_3737);
nand U3982 (N_3982,N_3040,N_3165);
nand U3983 (N_3983,N_3100,N_3523);
nor U3984 (N_3984,N_3671,N_3596);
nor U3985 (N_3985,N_3309,N_3140);
and U3986 (N_3986,N_3639,N_3299);
or U3987 (N_3987,N_3308,N_3164);
and U3988 (N_3988,N_3728,N_3497);
and U3989 (N_3989,N_3370,N_3209);
or U3990 (N_3990,N_3712,N_3323);
and U3991 (N_3991,N_3600,N_3332);
or U3992 (N_3992,N_3225,N_3242);
or U3993 (N_3993,N_3227,N_3286);
xor U3994 (N_3994,N_3582,N_3007);
nor U3995 (N_3995,N_3452,N_3579);
nand U3996 (N_3996,N_3653,N_3115);
or U3997 (N_3997,N_3437,N_3403);
nor U3998 (N_3998,N_3391,N_3666);
or U3999 (N_3999,N_3581,N_3459);
nor U4000 (N_4000,N_3474,N_3385);
nand U4001 (N_4001,N_3358,N_3016);
and U4002 (N_4002,N_3553,N_3727);
nor U4003 (N_4003,N_3075,N_3650);
and U4004 (N_4004,N_3559,N_3479);
nand U4005 (N_4005,N_3203,N_3461);
nand U4006 (N_4006,N_3198,N_3399);
or U4007 (N_4007,N_3352,N_3648);
nand U4008 (N_4008,N_3033,N_3716);
and U4009 (N_4009,N_3446,N_3688);
and U4010 (N_4010,N_3593,N_3569);
nand U4011 (N_4011,N_3230,N_3376);
and U4012 (N_4012,N_3210,N_3533);
or U4013 (N_4013,N_3123,N_3102);
and U4014 (N_4014,N_3664,N_3731);
nand U4015 (N_4015,N_3070,N_3576);
nand U4016 (N_4016,N_3341,N_3146);
nor U4017 (N_4017,N_3091,N_3136);
nand U4018 (N_4018,N_3704,N_3528);
nor U4019 (N_4019,N_3718,N_3319);
nor U4020 (N_4020,N_3289,N_3206);
nand U4021 (N_4021,N_3331,N_3564);
and U4022 (N_4022,N_3668,N_3282);
nand U4023 (N_4023,N_3670,N_3355);
and U4024 (N_4024,N_3545,N_3001);
or U4025 (N_4025,N_3591,N_3272);
and U4026 (N_4026,N_3354,N_3263);
and U4027 (N_4027,N_3243,N_3049);
and U4028 (N_4028,N_3375,N_3055);
and U4029 (N_4029,N_3568,N_3649);
or U4030 (N_4030,N_3383,N_3273);
nor U4031 (N_4031,N_3534,N_3693);
or U4032 (N_4032,N_3466,N_3521);
or U4033 (N_4033,N_3270,N_3698);
and U4034 (N_4034,N_3697,N_3502);
or U4035 (N_4035,N_3660,N_3120);
and U4036 (N_4036,N_3356,N_3714);
or U4037 (N_4037,N_3371,N_3228);
and U4038 (N_4038,N_3493,N_3168);
xor U4039 (N_4039,N_3659,N_3347);
nand U4040 (N_4040,N_3045,N_3423);
nand U4041 (N_4041,N_3511,N_3630);
nand U4042 (N_4042,N_3293,N_3095);
and U4043 (N_4043,N_3365,N_3141);
or U4044 (N_4044,N_3462,N_3343);
nor U4045 (N_4045,N_3359,N_3575);
or U4046 (N_4046,N_3617,N_3132);
or U4047 (N_4047,N_3317,N_3125);
and U4048 (N_4048,N_3279,N_3654);
and U4049 (N_4049,N_3580,N_3232);
and U4050 (N_4050,N_3411,N_3407);
nand U4051 (N_4051,N_3090,N_3177);
nand U4052 (N_4052,N_3305,N_3093);
or U4053 (N_4053,N_3296,N_3298);
nand U4054 (N_4054,N_3187,N_3053);
nand U4055 (N_4055,N_3713,N_3652);
or U4056 (N_4056,N_3034,N_3570);
nand U4057 (N_4057,N_3425,N_3249);
xnor U4058 (N_4058,N_3194,N_3417);
and U4059 (N_4059,N_3339,N_3562);
nand U4060 (N_4060,N_3543,N_3705);
nand U4061 (N_4061,N_3080,N_3042);
and U4062 (N_4062,N_3672,N_3333);
and U4063 (N_4063,N_3717,N_3613);
nor U4064 (N_4064,N_3701,N_3505);
nor U4065 (N_4065,N_3495,N_3223);
nand U4066 (N_4066,N_3176,N_3008);
nand U4067 (N_4067,N_3079,N_3622);
or U4068 (N_4068,N_3252,N_3044);
and U4069 (N_4069,N_3312,N_3345);
or U4070 (N_4070,N_3456,N_3068);
nor U4071 (N_4071,N_3173,N_3244);
nor U4072 (N_4072,N_3689,N_3181);
and U4073 (N_4073,N_3675,N_3599);
nand U4074 (N_4074,N_3730,N_3725);
nor U4075 (N_4075,N_3153,N_3306);
nand U4076 (N_4076,N_3154,N_3723);
or U4077 (N_4077,N_3226,N_3392);
nand U4078 (N_4078,N_3390,N_3105);
or U4079 (N_4079,N_3509,N_3360);
or U4080 (N_4080,N_3636,N_3143);
nand U4081 (N_4081,N_3342,N_3158);
and U4082 (N_4082,N_3118,N_3532);
or U4083 (N_4083,N_3464,N_3504);
nor U4084 (N_4084,N_3111,N_3241);
nand U4085 (N_4085,N_3238,N_3011);
nor U4086 (N_4086,N_3426,N_3361);
and U4087 (N_4087,N_3038,N_3454);
or U4088 (N_4088,N_3188,N_3499);
or U4089 (N_4089,N_3612,N_3015);
nor U4090 (N_4090,N_3588,N_3747);
and U4091 (N_4091,N_3692,N_3721);
xor U4092 (N_4092,N_3324,N_3424);
xnor U4093 (N_4093,N_3711,N_3271);
nand U4094 (N_4094,N_3000,N_3131);
nor U4095 (N_4095,N_3422,N_3503);
nand U4096 (N_4096,N_3246,N_3325);
nand U4097 (N_4097,N_3538,N_3290);
or U4098 (N_4098,N_3220,N_3573);
nand U4099 (N_4099,N_3160,N_3313);
nand U4100 (N_4100,N_3182,N_3092);
or U4101 (N_4101,N_3122,N_3174);
nand U4102 (N_4102,N_3492,N_3266);
nor U4103 (N_4103,N_3640,N_3400);
or U4104 (N_4104,N_3435,N_3302);
and U4105 (N_4105,N_3167,N_3415);
or U4106 (N_4106,N_3029,N_3250);
nand U4107 (N_4107,N_3608,N_3274);
nand U4108 (N_4108,N_3393,N_3394);
or U4109 (N_4109,N_3046,N_3397);
or U4110 (N_4110,N_3369,N_3476);
nand U4111 (N_4111,N_3457,N_3540);
or U4112 (N_4112,N_3439,N_3064);
nor U4113 (N_4113,N_3050,N_3382);
or U4114 (N_4114,N_3019,N_3110);
nand U4115 (N_4115,N_3601,N_3128);
and U4116 (N_4116,N_3486,N_3412);
nor U4117 (N_4117,N_3745,N_3084);
nor U4118 (N_4118,N_3269,N_3674);
or U4119 (N_4119,N_3107,N_3124);
or U4120 (N_4120,N_3088,N_3571);
nand U4121 (N_4121,N_3646,N_3396);
and U4122 (N_4122,N_3436,N_3316);
nand U4123 (N_4123,N_3719,N_3449);
or U4124 (N_4124,N_3520,N_3749);
nand U4125 (N_4125,N_3592,N_3326);
nor U4126 (N_4126,N_3481,N_3624);
nand U4127 (N_4127,N_3424,N_3380);
nor U4128 (N_4128,N_3400,N_3635);
nand U4129 (N_4129,N_3200,N_3340);
or U4130 (N_4130,N_3624,N_3156);
nor U4131 (N_4131,N_3423,N_3515);
and U4132 (N_4132,N_3076,N_3381);
or U4133 (N_4133,N_3565,N_3749);
nand U4134 (N_4134,N_3680,N_3145);
and U4135 (N_4135,N_3475,N_3272);
and U4136 (N_4136,N_3052,N_3588);
nand U4137 (N_4137,N_3295,N_3077);
nand U4138 (N_4138,N_3238,N_3738);
or U4139 (N_4139,N_3172,N_3225);
nand U4140 (N_4140,N_3230,N_3535);
or U4141 (N_4141,N_3458,N_3572);
or U4142 (N_4142,N_3181,N_3379);
nand U4143 (N_4143,N_3282,N_3386);
and U4144 (N_4144,N_3066,N_3647);
and U4145 (N_4145,N_3215,N_3316);
nand U4146 (N_4146,N_3551,N_3031);
or U4147 (N_4147,N_3565,N_3164);
nor U4148 (N_4148,N_3635,N_3409);
xor U4149 (N_4149,N_3223,N_3392);
nor U4150 (N_4150,N_3388,N_3409);
or U4151 (N_4151,N_3597,N_3679);
nor U4152 (N_4152,N_3297,N_3235);
or U4153 (N_4153,N_3065,N_3551);
nand U4154 (N_4154,N_3177,N_3415);
nor U4155 (N_4155,N_3268,N_3574);
or U4156 (N_4156,N_3674,N_3430);
and U4157 (N_4157,N_3197,N_3113);
or U4158 (N_4158,N_3369,N_3196);
nor U4159 (N_4159,N_3314,N_3416);
and U4160 (N_4160,N_3689,N_3749);
xor U4161 (N_4161,N_3695,N_3214);
and U4162 (N_4162,N_3504,N_3049);
or U4163 (N_4163,N_3304,N_3731);
xnor U4164 (N_4164,N_3517,N_3098);
or U4165 (N_4165,N_3325,N_3111);
nand U4166 (N_4166,N_3652,N_3504);
or U4167 (N_4167,N_3392,N_3043);
and U4168 (N_4168,N_3437,N_3234);
or U4169 (N_4169,N_3601,N_3257);
xor U4170 (N_4170,N_3249,N_3657);
xor U4171 (N_4171,N_3694,N_3347);
and U4172 (N_4172,N_3153,N_3032);
and U4173 (N_4173,N_3707,N_3503);
nand U4174 (N_4174,N_3720,N_3310);
or U4175 (N_4175,N_3478,N_3339);
and U4176 (N_4176,N_3017,N_3160);
xor U4177 (N_4177,N_3025,N_3124);
or U4178 (N_4178,N_3711,N_3654);
and U4179 (N_4179,N_3646,N_3383);
and U4180 (N_4180,N_3131,N_3196);
and U4181 (N_4181,N_3323,N_3304);
or U4182 (N_4182,N_3028,N_3434);
nand U4183 (N_4183,N_3624,N_3334);
nand U4184 (N_4184,N_3336,N_3015);
nand U4185 (N_4185,N_3698,N_3227);
nand U4186 (N_4186,N_3301,N_3487);
and U4187 (N_4187,N_3045,N_3419);
nand U4188 (N_4188,N_3662,N_3042);
or U4189 (N_4189,N_3328,N_3465);
or U4190 (N_4190,N_3730,N_3652);
or U4191 (N_4191,N_3677,N_3450);
and U4192 (N_4192,N_3492,N_3475);
nand U4193 (N_4193,N_3725,N_3178);
and U4194 (N_4194,N_3667,N_3109);
nand U4195 (N_4195,N_3022,N_3626);
and U4196 (N_4196,N_3579,N_3652);
nand U4197 (N_4197,N_3019,N_3618);
or U4198 (N_4198,N_3554,N_3000);
and U4199 (N_4199,N_3473,N_3659);
nor U4200 (N_4200,N_3736,N_3221);
nand U4201 (N_4201,N_3675,N_3121);
nand U4202 (N_4202,N_3191,N_3074);
nand U4203 (N_4203,N_3000,N_3621);
and U4204 (N_4204,N_3556,N_3076);
nand U4205 (N_4205,N_3739,N_3068);
nand U4206 (N_4206,N_3526,N_3655);
and U4207 (N_4207,N_3034,N_3117);
nor U4208 (N_4208,N_3299,N_3208);
and U4209 (N_4209,N_3620,N_3661);
and U4210 (N_4210,N_3557,N_3230);
or U4211 (N_4211,N_3649,N_3010);
and U4212 (N_4212,N_3003,N_3631);
nand U4213 (N_4213,N_3326,N_3572);
nand U4214 (N_4214,N_3091,N_3643);
and U4215 (N_4215,N_3049,N_3664);
xor U4216 (N_4216,N_3516,N_3746);
nor U4217 (N_4217,N_3635,N_3063);
nand U4218 (N_4218,N_3335,N_3087);
xnor U4219 (N_4219,N_3634,N_3188);
nand U4220 (N_4220,N_3311,N_3250);
and U4221 (N_4221,N_3197,N_3520);
or U4222 (N_4222,N_3146,N_3019);
nand U4223 (N_4223,N_3316,N_3219);
or U4224 (N_4224,N_3317,N_3189);
and U4225 (N_4225,N_3355,N_3010);
or U4226 (N_4226,N_3351,N_3553);
nor U4227 (N_4227,N_3249,N_3159);
nand U4228 (N_4228,N_3353,N_3468);
and U4229 (N_4229,N_3434,N_3341);
and U4230 (N_4230,N_3028,N_3299);
nand U4231 (N_4231,N_3022,N_3267);
nor U4232 (N_4232,N_3604,N_3656);
or U4233 (N_4233,N_3045,N_3193);
nor U4234 (N_4234,N_3172,N_3031);
nor U4235 (N_4235,N_3673,N_3555);
or U4236 (N_4236,N_3742,N_3048);
nand U4237 (N_4237,N_3743,N_3192);
or U4238 (N_4238,N_3469,N_3184);
or U4239 (N_4239,N_3483,N_3655);
or U4240 (N_4240,N_3574,N_3084);
nand U4241 (N_4241,N_3539,N_3417);
nand U4242 (N_4242,N_3593,N_3182);
or U4243 (N_4243,N_3567,N_3470);
and U4244 (N_4244,N_3737,N_3121);
or U4245 (N_4245,N_3527,N_3216);
nor U4246 (N_4246,N_3555,N_3477);
nand U4247 (N_4247,N_3084,N_3700);
nand U4248 (N_4248,N_3313,N_3721);
and U4249 (N_4249,N_3641,N_3419);
and U4250 (N_4250,N_3647,N_3229);
or U4251 (N_4251,N_3434,N_3199);
and U4252 (N_4252,N_3611,N_3046);
and U4253 (N_4253,N_3507,N_3330);
or U4254 (N_4254,N_3333,N_3067);
or U4255 (N_4255,N_3038,N_3394);
and U4256 (N_4256,N_3086,N_3601);
and U4257 (N_4257,N_3603,N_3401);
nor U4258 (N_4258,N_3436,N_3241);
nand U4259 (N_4259,N_3148,N_3427);
nand U4260 (N_4260,N_3343,N_3214);
or U4261 (N_4261,N_3535,N_3333);
and U4262 (N_4262,N_3734,N_3738);
or U4263 (N_4263,N_3546,N_3141);
nand U4264 (N_4264,N_3548,N_3439);
or U4265 (N_4265,N_3593,N_3463);
nand U4266 (N_4266,N_3499,N_3226);
nor U4267 (N_4267,N_3742,N_3533);
and U4268 (N_4268,N_3067,N_3345);
nor U4269 (N_4269,N_3161,N_3477);
and U4270 (N_4270,N_3572,N_3171);
or U4271 (N_4271,N_3077,N_3603);
or U4272 (N_4272,N_3332,N_3224);
xor U4273 (N_4273,N_3629,N_3336);
nor U4274 (N_4274,N_3232,N_3094);
or U4275 (N_4275,N_3242,N_3611);
and U4276 (N_4276,N_3120,N_3633);
nand U4277 (N_4277,N_3588,N_3428);
and U4278 (N_4278,N_3165,N_3254);
xnor U4279 (N_4279,N_3501,N_3742);
and U4280 (N_4280,N_3072,N_3210);
or U4281 (N_4281,N_3532,N_3522);
nor U4282 (N_4282,N_3571,N_3476);
or U4283 (N_4283,N_3422,N_3403);
nor U4284 (N_4284,N_3110,N_3244);
nor U4285 (N_4285,N_3260,N_3273);
and U4286 (N_4286,N_3586,N_3489);
nor U4287 (N_4287,N_3092,N_3542);
and U4288 (N_4288,N_3656,N_3277);
or U4289 (N_4289,N_3712,N_3321);
and U4290 (N_4290,N_3007,N_3549);
xnor U4291 (N_4291,N_3005,N_3123);
and U4292 (N_4292,N_3396,N_3067);
xor U4293 (N_4293,N_3684,N_3183);
and U4294 (N_4294,N_3078,N_3286);
nor U4295 (N_4295,N_3363,N_3111);
and U4296 (N_4296,N_3070,N_3430);
nand U4297 (N_4297,N_3518,N_3395);
nand U4298 (N_4298,N_3163,N_3318);
nor U4299 (N_4299,N_3067,N_3246);
and U4300 (N_4300,N_3498,N_3608);
nor U4301 (N_4301,N_3292,N_3221);
or U4302 (N_4302,N_3009,N_3327);
and U4303 (N_4303,N_3605,N_3371);
nor U4304 (N_4304,N_3398,N_3324);
nand U4305 (N_4305,N_3644,N_3103);
nor U4306 (N_4306,N_3558,N_3614);
nor U4307 (N_4307,N_3152,N_3559);
nor U4308 (N_4308,N_3454,N_3631);
or U4309 (N_4309,N_3502,N_3293);
or U4310 (N_4310,N_3032,N_3210);
nor U4311 (N_4311,N_3185,N_3378);
and U4312 (N_4312,N_3305,N_3029);
nor U4313 (N_4313,N_3340,N_3737);
and U4314 (N_4314,N_3398,N_3568);
and U4315 (N_4315,N_3585,N_3380);
or U4316 (N_4316,N_3297,N_3293);
nor U4317 (N_4317,N_3177,N_3329);
and U4318 (N_4318,N_3522,N_3652);
nand U4319 (N_4319,N_3171,N_3241);
and U4320 (N_4320,N_3535,N_3489);
and U4321 (N_4321,N_3202,N_3402);
nand U4322 (N_4322,N_3175,N_3257);
nor U4323 (N_4323,N_3610,N_3496);
and U4324 (N_4324,N_3583,N_3537);
and U4325 (N_4325,N_3695,N_3722);
and U4326 (N_4326,N_3178,N_3170);
and U4327 (N_4327,N_3551,N_3529);
nand U4328 (N_4328,N_3625,N_3518);
or U4329 (N_4329,N_3313,N_3106);
and U4330 (N_4330,N_3578,N_3741);
and U4331 (N_4331,N_3691,N_3541);
nor U4332 (N_4332,N_3371,N_3741);
and U4333 (N_4333,N_3282,N_3358);
and U4334 (N_4334,N_3248,N_3174);
and U4335 (N_4335,N_3579,N_3418);
nor U4336 (N_4336,N_3127,N_3540);
nor U4337 (N_4337,N_3739,N_3101);
and U4338 (N_4338,N_3018,N_3135);
nand U4339 (N_4339,N_3590,N_3319);
xnor U4340 (N_4340,N_3109,N_3012);
nand U4341 (N_4341,N_3709,N_3520);
nand U4342 (N_4342,N_3736,N_3089);
nand U4343 (N_4343,N_3299,N_3529);
nor U4344 (N_4344,N_3470,N_3071);
nor U4345 (N_4345,N_3490,N_3350);
or U4346 (N_4346,N_3669,N_3290);
nand U4347 (N_4347,N_3633,N_3747);
nand U4348 (N_4348,N_3209,N_3077);
nand U4349 (N_4349,N_3323,N_3050);
nand U4350 (N_4350,N_3367,N_3485);
or U4351 (N_4351,N_3058,N_3718);
xor U4352 (N_4352,N_3069,N_3147);
and U4353 (N_4353,N_3675,N_3369);
or U4354 (N_4354,N_3251,N_3262);
or U4355 (N_4355,N_3681,N_3058);
or U4356 (N_4356,N_3515,N_3736);
nand U4357 (N_4357,N_3740,N_3061);
nand U4358 (N_4358,N_3448,N_3388);
nor U4359 (N_4359,N_3670,N_3531);
nand U4360 (N_4360,N_3256,N_3308);
nor U4361 (N_4361,N_3183,N_3081);
nor U4362 (N_4362,N_3567,N_3575);
nand U4363 (N_4363,N_3688,N_3171);
or U4364 (N_4364,N_3361,N_3132);
nor U4365 (N_4365,N_3509,N_3331);
and U4366 (N_4366,N_3363,N_3583);
nor U4367 (N_4367,N_3331,N_3642);
xor U4368 (N_4368,N_3083,N_3000);
nand U4369 (N_4369,N_3492,N_3349);
and U4370 (N_4370,N_3393,N_3530);
or U4371 (N_4371,N_3058,N_3257);
nand U4372 (N_4372,N_3504,N_3011);
and U4373 (N_4373,N_3335,N_3258);
nor U4374 (N_4374,N_3288,N_3198);
and U4375 (N_4375,N_3427,N_3744);
nor U4376 (N_4376,N_3034,N_3507);
or U4377 (N_4377,N_3203,N_3497);
and U4378 (N_4378,N_3467,N_3051);
or U4379 (N_4379,N_3467,N_3551);
nand U4380 (N_4380,N_3401,N_3512);
nand U4381 (N_4381,N_3572,N_3280);
and U4382 (N_4382,N_3260,N_3087);
or U4383 (N_4383,N_3064,N_3649);
nor U4384 (N_4384,N_3059,N_3146);
nor U4385 (N_4385,N_3138,N_3420);
or U4386 (N_4386,N_3642,N_3111);
nand U4387 (N_4387,N_3511,N_3748);
xor U4388 (N_4388,N_3146,N_3202);
nor U4389 (N_4389,N_3696,N_3095);
or U4390 (N_4390,N_3382,N_3145);
and U4391 (N_4391,N_3095,N_3114);
nor U4392 (N_4392,N_3262,N_3218);
or U4393 (N_4393,N_3243,N_3183);
nor U4394 (N_4394,N_3439,N_3616);
or U4395 (N_4395,N_3534,N_3688);
and U4396 (N_4396,N_3103,N_3312);
nand U4397 (N_4397,N_3088,N_3321);
nand U4398 (N_4398,N_3086,N_3305);
or U4399 (N_4399,N_3183,N_3156);
nand U4400 (N_4400,N_3466,N_3681);
nand U4401 (N_4401,N_3535,N_3683);
nor U4402 (N_4402,N_3474,N_3700);
or U4403 (N_4403,N_3322,N_3522);
nor U4404 (N_4404,N_3050,N_3247);
and U4405 (N_4405,N_3674,N_3390);
nor U4406 (N_4406,N_3127,N_3059);
nor U4407 (N_4407,N_3061,N_3718);
nor U4408 (N_4408,N_3348,N_3651);
nor U4409 (N_4409,N_3202,N_3247);
nand U4410 (N_4410,N_3167,N_3197);
and U4411 (N_4411,N_3675,N_3638);
nor U4412 (N_4412,N_3026,N_3333);
or U4413 (N_4413,N_3373,N_3522);
and U4414 (N_4414,N_3293,N_3617);
or U4415 (N_4415,N_3470,N_3676);
or U4416 (N_4416,N_3085,N_3047);
and U4417 (N_4417,N_3598,N_3321);
or U4418 (N_4418,N_3126,N_3236);
and U4419 (N_4419,N_3034,N_3551);
or U4420 (N_4420,N_3627,N_3615);
nand U4421 (N_4421,N_3350,N_3487);
nand U4422 (N_4422,N_3667,N_3197);
nor U4423 (N_4423,N_3099,N_3631);
nor U4424 (N_4424,N_3180,N_3392);
or U4425 (N_4425,N_3616,N_3395);
nor U4426 (N_4426,N_3404,N_3585);
and U4427 (N_4427,N_3250,N_3481);
nor U4428 (N_4428,N_3372,N_3580);
and U4429 (N_4429,N_3646,N_3257);
or U4430 (N_4430,N_3004,N_3540);
nand U4431 (N_4431,N_3133,N_3561);
nand U4432 (N_4432,N_3128,N_3530);
and U4433 (N_4433,N_3557,N_3334);
or U4434 (N_4434,N_3604,N_3064);
nand U4435 (N_4435,N_3519,N_3489);
nand U4436 (N_4436,N_3598,N_3407);
or U4437 (N_4437,N_3045,N_3137);
nand U4438 (N_4438,N_3418,N_3135);
and U4439 (N_4439,N_3683,N_3603);
or U4440 (N_4440,N_3322,N_3435);
xnor U4441 (N_4441,N_3129,N_3616);
and U4442 (N_4442,N_3481,N_3109);
and U4443 (N_4443,N_3336,N_3443);
and U4444 (N_4444,N_3451,N_3637);
nand U4445 (N_4445,N_3591,N_3435);
nand U4446 (N_4446,N_3001,N_3060);
nand U4447 (N_4447,N_3507,N_3445);
or U4448 (N_4448,N_3232,N_3604);
nand U4449 (N_4449,N_3407,N_3029);
nand U4450 (N_4450,N_3414,N_3027);
nor U4451 (N_4451,N_3303,N_3615);
nor U4452 (N_4452,N_3416,N_3067);
nand U4453 (N_4453,N_3205,N_3714);
xor U4454 (N_4454,N_3101,N_3697);
nor U4455 (N_4455,N_3526,N_3253);
and U4456 (N_4456,N_3614,N_3508);
and U4457 (N_4457,N_3498,N_3731);
or U4458 (N_4458,N_3719,N_3101);
or U4459 (N_4459,N_3298,N_3265);
xor U4460 (N_4460,N_3520,N_3746);
or U4461 (N_4461,N_3462,N_3116);
nor U4462 (N_4462,N_3361,N_3316);
nor U4463 (N_4463,N_3406,N_3281);
or U4464 (N_4464,N_3183,N_3509);
nand U4465 (N_4465,N_3103,N_3118);
xor U4466 (N_4466,N_3677,N_3660);
xor U4467 (N_4467,N_3476,N_3309);
and U4468 (N_4468,N_3387,N_3488);
or U4469 (N_4469,N_3060,N_3729);
nor U4470 (N_4470,N_3693,N_3332);
or U4471 (N_4471,N_3309,N_3011);
xnor U4472 (N_4472,N_3309,N_3479);
nor U4473 (N_4473,N_3005,N_3383);
or U4474 (N_4474,N_3154,N_3556);
and U4475 (N_4475,N_3660,N_3457);
and U4476 (N_4476,N_3001,N_3391);
or U4477 (N_4477,N_3587,N_3127);
or U4478 (N_4478,N_3453,N_3436);
nand U4479 (N_4479,N_3093,N_3177);
nor U4480 (N_4480,N_3636,N_3111);
and U4481 (N_4481,N_3349,N_3115);
nand U4482 (N_4482,N_3146,N_3217);
or U4483 (N_4483,N_3009,N_3470);
nand U4484 (N_4484,N_3561,N_3400);
and U4485 (N_4485,N_3162,N_3385);
nor U4486 (N_4486,N_3497,N_3143);
and U4487 (N_4487,N_3171,N_3158);
and U4488 (N_4488,N_3719,N_3732);
nand U4489 (N_4489,N_3006,N_3152);
or U4490 (N_4490,N_3110,N_3589);
nor U4491 (N_4491,N_3601,N_3407);
or U4492 (N_4492,N_3426,N_3739);
or U4493 (N_4493,N_3569,N_3437);
and U4494 (N_4494,N_3609,N_3541);
or U4495 (N_4495,N_3553,N_3394);
and U4496 (N_4496,N_3656,N_3224);
and U4497 (N_4497,N_3296,N_3254);
and U4498 (N_4498,N_3661,N_3714);
nor U4499 (N_4499,N_3265,N_3005);
xor U4500 (N_4500,N_3768,N_3964);
and U4501 (N_4501,N_4319,N_3841);
nor U4502 (N_4502,N_4169,N_4391);
and U4503 (N_4503,N_4092,N_4235);
and U4504 (N_4504,N_4332,N_4250);
or U4505 (N_4505,N_4167,N_4443);
and U4506 (N_4506,N_4165,N_3829);
nor U4507 (N_4507,N_3984,N_4344);
xor U4508 (N_4508,N_4038,N_4121);
or U4509 (N_4509,N_4021,N_4042);
and U4510 (N_4510,N_4425,N_4362);
nor U4511 (N_4511,N_4124,N_4017);
nor U4512 (N_4512,N_4420,N_4396);
nand U4513 (N_4513,N_4211,N_4137);
or U4514 (N_4514,N_4227,N_4143);
nand U4515 (N_4515,N_3896,N_3949);
nor U4516 (N_4516,N_4263,N_3876);
xnor U4517 (N_4517,N_3756,N_4252);
nand U4518 (N_4518,N_3918,N_4027);
or U4519 (N_4519,N_4113,N_3921);
nand U4520 (N_4520,N_4437,N_4152);
or U4521 (N_4521,N_4091,N_4019);
or U4522 (N_4522,N_4482,N_3831);
nor U4523 (N_4523,N_3989,N_4216);
and U4524 (N_4524,N_4006,N_4142);
nand U4525 (N_4525,N_4457,N_3889);
or U4526 (N_4526,N_4181,N_3995);
nor U4527 (N_4527,N_3827,N_4005);
or U4528 (N_4528,N_4179,N_3779);
nand U4529 (N_4529,N_3903,N_4034);
or U4530 (N_4530,N_4207,N_4088);
and U4531 (N_4531,N_4046,N_3913);
and U4532 (N_4532,N_3825,N_4233);
and U4533 (N_4533,N_4444,N_3856);
nand U4534 (N_4534,N_4246,N_3833);
and U4535 (N_4535,N_4297,N_4101);
nor U4536 (N_4536,N_4369,N_3867);
nor U4537 (N_4537,N_4161,N_4056);
and U4538 (N_4538,N_3920,N_4162);
nor U4539 (N_4539,N_3917,N_4083);
nor U4540 (N_4540,N_4125,N_3916);
and U4541 (N_4541,N_4203,N_3847);
or U4542 (N_4542,N_4397,N_4290);
nor U4543 (N_4543,N_3800,N_4377);
nor U4544 (N_4544,N_3873,N_4243);
nand U4545 (N_4545,N_4172,N_4331);
or U4546 (N_4546,N_3753,N_4469);
nand U4547 (N_4547,N_4176,N_4132);
nand U4548 (N_4548,N_4418,N_4385);
nor U4549 (N_4549,N_3990,N_4007);
nor U4550 (N_4550,N_4242,N_3924);
nand U4551 (N_4551,N_4256,N_4366);
nand U4552 (N_4552,N_4423,N_4388);
nor U4553 (N_4553,N_3801,N_4177);
and U4554 (N_4554,N_3969,N_4382);
nand U4555 (N_4555,N_4085,N_4342);
nor U4556 (N_4556,N_3868,N_4267);
nor U4557 (N_4557,N_4004,N_3946);
nor U4558 (N_4558,N_4470,N_3793);
nor U4559 (N_4559,N_4458,N_4001);
nand U4560 (N_4560,N_3872,N_3846);
nand U4561 (N_4561,N_4071,N_4089);
or U4562 (N_4562,N_4214,N_4310);
and U4563 (N_4563,N_3851,N_4410);
nand U4564 (N_4564,N_4052,N_3863);
nand U4565 (N_4565,N_4221,N_4253);
or U4566 (N_4566,N_3790,N_3798);
nand U4567 (N_4567,N_4066,N_4183);
nand U4568 (N_4568,N_4130,N_3973);
nand U4569 (N_4569,N_4204,N_4341);
xnor U4570 (N_4570,N_4449,N_3882);
nand U4571 (N_4571,N_3776,N_4020);
xor U4572 (N_4572,N_4286,N_4481);
xnor U4573 (N_4573,N_4412,N_4315);
nand U4574 (N_4574,N_3771,N_3997);
nand U4575 (N_4575,N_4333,N_4273);
or U4576 (N_4576,N_3961,N_4245);
nor U4577 (N_4577,N_3774,N_4055);
and U4578 (N_4578,N_3762,N_3783);
nand U4579 (N_4579,N_3957,N_4431);
and U4580 (N_4580,N_4447,N_3862);
nand U4581 (N_4581,N_4467,N_3906);
nor U4582 (N_4582,N_4129,N_4300);
or U4583 (N_4583,N_4257,N_3926);
nand U4584 (N_4584,N_3815,N_4361);
and U4585 (N_4585,N_4039,N_4475);
or U4586 (N_4586,N_4115,N_4002);
nor U4587 (N_4587,N_4059,N_4346);
and U4588 (N_4588,N_4483,N_3781);
and U4589 (N_4589,N_4240,N_4160);
or U4590 (N_4590,N_3871,N_4474);
and U4591 (N_4591,N_4477,N_4280);
nand U4592 (N_4592,N_3999,N_4304);
nand U4593 (N_4593,N_4104,N_4394);
or U4594 (N_4594,N_3890,N_3767);
and U4595 (N_4595,N_4222,N_4419);
and U4596 (N_4596,N_4186,N_4248);
and U4597 (N_4597,N_4368,N_4321);
and U4598 (N_4598,N_4069,N_4223);
nor U4599 (N_4599,N_3757,N_4175);
nand U4600 (N_4600,N_3760,N_4465);
and U4601 (N_4601,N_4239,N_3881);
or U4602 (N_4602,N_3861,N_4359);
xnor U4603 (N_4603,N_4099,N_3939);
nand U4604 (N_4604,N_4312,N_4429);
or U4605 (N_4605,N_3859,N_4164);
nor U4606 (N_4606,N_4105,N_4014);
and U4607 (N_4607,N_3884,N_4276);
nand U4608 (N_4608,N_3979,N_4451);
or U4609 (N_4609,N_4070,N_3848);
and U4610 (N_4610,N_4249,N_4217);
or U4611 (N_4611,N_3796,N_3845);
and U4612 (N_4612,N_4330,N_4324);
nor U4613 (N_4613,N_3799,N_3971);
xor U4614 (N_4614,N_4422,N_4180);
nor U4615 (N_4615,N_3943,N_3895);
and U4616 (N_4616,N_4343,N_4018);
nand U4617 (N_4617,N_3878,N_3934);
or U4618 (N_4618,N_3883,N_4197);
nor U4619 (N_4619,N_4277,N_4023);
and U4620 (N_4620,N_3816,N_4199);
nand U4621 (N_4621,N_4490,N_3817);
nand U4622 (N_4622,N_4148,N_3879);
nand U4623 (N_4623,N_3955,N_3803);
and U4624 (N_4624,N_4141,N_4285);
or U4625 (N_4625,N_4212,N_4426);
nand U4626 (N_4626,N_4287,N_3849);
nor U4627 (N_4627,N_4261,N_4030);
or U4628 (N_4628,N_4355,N_4358);
nor U4629 (N_4629,N_4062,N_3870);
nor U4630 (N_4630,N_4053,N_4238);
or U4631 (N_4631,N_4182,N_4436);
nand U4632 (N_4632,N_4380,N_4260);
and U4633 (N_4633,N_3869,N_4283);
and U4634 (N_4634,N_4155,N_4201);
and U4635 (N_4635,N_4045,N_3897);
nor U4636 (N_4636,N_3818,N_4026);
nand U4637 (N_4637,N_4365,N_4299);
nand U4638 (N_4638,N_4131,N_4356);
and U4639 (N_4639,N_4414,N_3789);
nor U4640 (N_4640,N_4051,N_4371);
or U4641 (N_4641,N_4008,N_3919);
or U4642 (N_4642,N_3925,N_3852);
or U4643 (N_4643,N_3810,N_3911);
or U4644 (N_4644,N_3751,N_4270);
and U4645 (N_4645,N_4320,N_3900);
and U4646 (N_4646,N_4236,N_3770);
nor U4647 (N_4647,N_4398,N_3907);
or U4648 (N_4648,N_4405,N_3891);
and U4649 (N_4649,N_3759,N_4067);
nor U4650 (N_4650,N_4033,N_3953);
or U4651 (N_4651,N_4171,N_4284);
and U4652 (N_4652,N_4488,N_3940);
or U4653 (N_4653,N_4140,N_4135);
or U4654 (N_4654,N_3806,N_4118);
and U4655 (N_4655,N_3865,N_4448);
nor U4656 (N_4656,N_4090,N_4187);
nand U4657 (N_4657,N_4413,N_4439);
nand U4658 (N_4658,N_4190,N_3792);
nor U4659 (N_4659,N_4074,N_4213);
and U4660 (N_4660,N_4079,N_3755);
nor U4661 (N_4661,N_4219,N_4076);
and U4662 (N_4662,N_3763,N_3772);
nand U4663 (N_4663,N_4293,N_4499);
nor U4664 (N_4664,N_4100,N_4068);
nor U4665 (N_4665,N_4146,N_3786);
nand U4666 (N_4666,N_4196,N_4226);
and U4667 (N_4667,N_3923,N_4268);
nand U4668 (N_4668,N_4220,N_4145);
or U4669 (N_4669,N_4061,N_3823);
nor U4670 (N_4670,N_4072,N_4107);
nor U4671 (N_4671,N_3858,N_4188);
and U4672 (N_4672,N_3974,N_4112);
or U4673 (N_4673,N_4054,N_4440);
or U4674 (N_4674,N_3758,N_4336);
nand U4675 (N_4675,N_3909,N_3777);
nor U4676 (N_4676,N_3780,N_4254);
and U4677 (N_4677,N_3988,N_3855);
nor U4678 (N_4678,N_4339,N_4379);
and U4679 (N_4679,N_3922,N_4210);
or U4680 (N_4680,N_4228,N_3993);
nand U4681 (N_4681,N_3931,N_4328);
nand U4682 (N_4682,N_3854,N_4127);
and U4683 (N_4683,N_3945,N_3965);
or U4684 (N_4684,N_4114,N_4464);
or U4685 (N_4685,N_4432,N_4073);
nor U4686 (N_4686,N_4064,N_4029);
nand U4687 (N_4687,N_3936,N_4375);
and U4688 (N_4688,N_4109,N_4258);
nor U4689 (N_4689,N_4275,N_4234);
and U4690 (N_4690,N_4103,N_4364);
nor U4691 (N_4691,N_4279,N_3933);
nand U4692 (N_4692,N_3832,N_4349);
nor U4693 (N_4693,N_3948,N_4274);
or U4694 (N_4694,N_3912,N_3941);
or U4695 (N_4695,N_3814,N_4435);
nor U4696 (N_4696,N_4392,N_4462);
and U4697 (N_4697,N_4357,N_4360);
nand U4698 (N_4698,N_4408,N_4494);
and U4699 (N_4699,N_4496,N_3812);
and U4700 (N_4700,N_4466,N_3932);
nand U4701 (N_4701,N_4136,N_4093);
nand U4702 (N_4702,N_4097,N_3788);
nand U4703 (N_4703,N_4173,N_3977);
or U4704 (N_4704,N_3985,N_4215);
or U4705 (N_4705,N_3902,N_3966);
nand U4706 (N_4706,N_4126,N_4191);
nand U4707 (N_4707,N_4024,N_3915);
nand U4708 (N_4708,N_4086,N_4230);
and U4709 (N_4709,N_4291,N_4484);
or U4710 (N_4710,N_4278,N_4325);
and U4711 (N_4711,N_4307,N_4225);
or U4712 (N_4712,N_3886,N_3835);
nor U4713 (N_4713,N_4170,N_4015);
or U4714 (N_4714,N_4031,N_4348);
or U4715 (N_4715,N_4306,N_4195);
nor U4716 (N_4716,N_4208,N_3982);
nor U4717 (N_4717,N_4163,N_3842);
nor U4718 (N_4718,N_3824,N_4317);
nor U4719 (N_4719,N_4049,N_4157);
and U4720 (N_4720,N_4446,N_4495);
or U4721 (N_4721,N_3782,N_4288);
or U4722 (N_4722,N_4231,N_4373);
nor U4723 (N_4723,N_4037,N_3766);
or U4724 (N_4724,N_3938,N_4400);
xnor U4725 (N_4725,N_4032,N_4116);
or U4726 (N_4726,N_4158,N_4036);
and U4727 (N_4727,N_4292,N_4189);
nand U4728 (N_4728,N_4117,N_4282);
and U4729 (N_4729,N_4318,N_4184);
nor U4730 (N_4730,N_4119,N_4266);
and U4731 (N_4731,N_3797,N_4430);
nand U4732 (N_4732,N_4347,N_3983);
and U4733 (N_4733,N_4156,N_4218);
or U4734 (N_4734,N_4301,N_4308);
or U4735 (N_4735,N_3956,N_4095);
nor U4736 (N_4736,N_4147,N_4383);
or U4737 (N_4737,N_4337,N_3980);
or U4738 (N_4738,N_3765,N_4192);
or U4739 (N_4739,N_3857,N_4098);
nand U4740 (N_4740,N_4200,N_4402);
or U4741 (N_4741,N_4372,N_3795);
nor U4742 (N_4742,N_3761,N_3996);
nand U4743 (N_4743,N_3877,N_3808);
xnor U4744 (N_4744,N_3785,N_3944);
and U4745 (N_4745,N_4271,N_4123);
and U4746 (N_4746,N_4351,N_4247);
and U4747 (N_4747,N_3950,N_4009);
and U4748 (N_4748,N_4133,N_3844);
and U4749 (N_4749,N_4237,N_3826);
and U4750 (N_4750,N_3910,N_4012);
or U4751 (N_4751,N_4498,N_4106);
nand U4752 (N_4752,N_4082,N_4077);
or U4753 (N_4753,N_3853,N_3998);
nand U4754 (N_4754,N_4434,N_4111);
or U4755 (N_4755,N_3930,N_4013);
nand U4756 (N_4756,N_3821,N_4178);
and U4757 (N_4757,N_3894,N_4416);
or U4758 (N_4758,N_3874,N_4326);
nor U4759 (N_4759,N_3764,N_3811);
or U4760 (N_4760,N_3914,N_3836);
nand U4761 (N_4761,N_4108,N_4417);
and U4762 (N_4762,N_4468,N_3843);
or U4763 (N_4763,N_4194,N_4244);
and U4764 (N_4764,N_4303,N_4340);
and U4765 (N_4765,N_4487,N_4120);
or U4766 (N_4766,N_4035,N_4044);
and U4767 (N_4767,N_3794,N_4472);
nand U4768 (N_4768,N_4370,N_3834);
nand U4769 (N_4769,N_4314,N_3840);
nor U4770 (N_4770,N_4043,N_4265);
nand U4771 (N_4771,N_4353,N_4491);
or U4772 (N_4772,N_4471,N_3850);
nor U4773 (N_4773,N_4463,N_3970);
nor U4774 (N_4774,N_4084,N_4493);
and U4775 (N_4775,N_4305,N_4461);
nand U4776 (N_4776,N_3937,N_3864);
or U4777 (N_4777,N_3986,N_3975);
nand U4778 (N_4778,N_3991,N_4048);
or U4779 (N_4779,N_4205,N_4322);
xor U4780 (N_4780,N_4080,N_3830);
nand U4781 (N_4781,N_4150,N_3901);
nor U4782 (N_4782,N_4441,N_3787);
and U4783 (N_4783,N_4010,N_4040);
and U4784 (N_4784,N_4241,N_4232);
nand U4785 (N_4785,N_4486,N_3750);
or U4786 (N_4786,N_3822,N_4403);
nand U4787 (N_4787,N_4011,N_3778);
nand U4788 (N_4788,N_4294,N_4153);
nor U4789 (N_4789,N_4445,N_4255);
nor U4790 (N_4790,N_4442,N_3981);
and U4791 (N_4791,N_4473,N_4058);
nand U4792 (N_4792,N_4309,N_3875);
or U4793 (N_4793,N_4025,N_3813);
nand U4794 (N_4794,N_3898,N_3976);
and U4795 (N_4795,N_4295,N_4262);
or U4796 (N_4796,N_4453,N_4259);
nand U4797 (N_4797,N_4063,N_4459);
nor U4798 (N_4798,N_3828,N_4438);
and U4799 (N_4799,N_4057,N_3942);
nor U4800 (N_4800,N_3805,N_3978);
or U4801 (N_4801,N_4381,N_4193);
xnor U4802 (N_4802,N_3807,N_4404);
nor U4803 (N_4803,N_4128,N_4393);
and U4804 (N_4804,N_4311,N_4354);
or U4805 (N_4805,N_3947,N_4078);
and U4806 (N_4806,N_4159,N_4428);
or U4807 (N_4807,N_4485,N_4022);
nand U4808 (N_4808,N_4229,N_3804);
nand U4809 (N_4809,N_4352,N_4289);
nor U4810 (N_4810,N_3866,N_3809);
xnor U4811 (N_4811,N_3927,N_3928);
and U4812 (N_4812,N_4345,N_4478);
or U4813 (N_4813,N_3954,N_3880);
nand U4814 (N_4814,N_4224,N_4096);
nor U4815 (N_4815,N_4387,N_4350);
nand U4816 (N_4816,N_3754,N_3992);
nand U4817 (N_4817,N_4406,N_3987);
nand U4818 (N_4818,N_3962,N_3820);
nor U4819 (N_4819,N_4047,N_4313);
and U4820 (N_4820,N_4401,N_4122);
and U4821 (N_4821,N_4087,N_4094);
and U4822 (N_4822,N_4427,N_4460);
nor U4823 (N_4823,N_3838,N_4492);
nor U4824 (N_4824,N_4302,N_4003);
and U4825 (N_4825,N_4075,N_3802);
nor U4826 (N_4826,N_4338,N_3752);
nand U4827 (N_4827,N_4264,N_3887);
or U4828 (N_4828,N_4378,N_4479);
nor U4829 (N_4829,N_4110,N_4102);
nor U4830 (N_4830,N_4407,N_4415);
or U4831 (N_4831,N_4480,N_3784);
nor U4832 (N_4832,N_4386,N_4395);
nand U4833 (N_4833,N_3905,N_4376);
or U4834 (N_4834,N_4296,N_4489);
or U4835 (N_4835,N_4456,N_3791);
or U4836 (N_4836,N_3769,N_3908);
xor U4837 (N_4837,N_4041,N_4198);
nor U4838 (N_4838,N_4455,N_4374);
nor U4839 (N_4839,N_4327,N_3929);
nor U4840 (N_4840,N_3958,N_4334);
or U4841 (N_4841,N_3960,N_3967);
nor U4842 (N_4842,N_3952,N_4272);
or U4843 (N_4843,N_4185,N_4450);
nand U4844 (N_4844,N_4433,N_4138);
xnor U4845 (N_4845,N_4166,N_4316);
nor U4846 (N_4846,N_4060,N_4174);
or U4847 (N_4847,N_3968,N_3963);
and U4848 (N_4848,N_3775,N_3892);
nor U4849 (N_4849,N_3994,N_4421);
or U4850 (N_4850,N_4452,N_4298);
nor U4851 (N_4851,N_3839,N_4390);
and U4852 (N_4852,N_3837,N_4281);
or U4853 (N_4853,N_4454,N_4335);
or U4854 (N_4854,N_4144,N_4363);
nand U4855 (N_4855,N_3819,N_3959);
nor U4856 (N_4856,N_3888,N_3773);
and U4857 (N_4857,N_3972,N_4389);
nor U4858 (N_4858,N_4497,N_4168);
or U4859 (N_4859,N_3899,N_4134);
and U4860 (N_4860,N_4323,N_4139);
or U4861 (N_4861,N_3904,N_3885);
and U4862 (N_4862,N_3951,N_4409);
and U4863 (N_4863,N_3935,N_4028);
and U4864 (N_4864,N_4411,N_4384);
xnor U4865 (N_4865,N_4269,N_4000);
xor U4866 (N_4866,N_4050,N_4154);
nand U4867 (N_4867,N_4151,N_4016);
and U4868 (N_4868,N_4399,N_4424);
or U4869 (N_4869,N_4476,N_4081);
nand U4870 (N_4870,N_3860,N_4251);
or U4871 (N_4871,N_4367,N_4149);
and U4872 (N_4872,N_4065,N_4209);
nand U4873 (N_4873,N_4206,N_3893);
or U4874 (N_4874,N_4202,N_4329);
and U4875 (N_4875,N_3838,N_3871);
and U4876 (N_4876,N_4024,N_3768);
nor U4877 (N_4877,N_4388,N_3896);
nor U4878 (N_4878,N_3934,N_4247);
nand U4879 (N_4879,N_4265,N_4139);
nor U4880 (N_4880,N_3928,N_4432);
nor U4881 (N_4881,N_3922,N_3851);
nand U4882 (N_4882,N_4336,N_4273);
nor U4883 (N_4883,N_4167,N_4157);
nor U4884 (N_4884,N_4251,N_4057);
and U4885 (N_4885,N_4231,N_4406);
or U4886 (N_4886,N_4297,N_4177);
and U4887 (N_4887,N_4036,N_3898);
nor U4888 (N_4888,N_4438,N_4435);
and U4889 (N_4889,N_4392,N_4194);
nand U4890 (N_4890,N_4382,N_4246);
or U4891 (N_4891,N_3837,N_4118);
or U4892 (N_4892,N_4408,N_4431);
nand U4893 (N_4893,N_4169,N_4233);
nand U4894 (N_4894,N_4460,N_3914);
nand U4895 (N_4895,N_4292,N_4225);
nand U4896 (N_4896,N_4221,N_3944);
nand U4897 (N_4897,N_3933,N_4433);
nand U4898 (N_4898,N_4037,N_4265);
nand U4899 (N_4899,N_4036,N_4379);
nor U4900 (N_4900,N_4309,N_4477);
and U4901 (N_4901,N_4089,N_4416);
or U4902 (N_4902,N_4046,N_3944);
or U4903 (N_4903,N_4207,N_3803);
nor U4904 (N_4904,N_4296,N_4412);
or U4905 (N_4905,N_4305,N_4360);
nand U4906 (N_4906,N_3948,N_4016);
or U4907 (N_4907,N_4410,N_4007);
nor U4908 (N_4908,N_3849,N_3775);
nor U4909 (N_4909,N_3993,N_4039);
or U4910 (N_4910,N_4152,N_3764);
nand U4911 (N_4911,N_4009,N_4333);
nor U4912 (N_4912,N_3857,N_3908);
or U4913 (N_4913,N_4360,N_4183);
or U4914 (N_4914,N_4133,N_4034);
and U4915 (N_4915,N_4332,N_4122);
nor U4916 (N_4916,N_3813,N_4206);
xnor U4917 (N_4917,N_3999,N_4080);
nand U4918 (N_4918,N_4181,N_4363);
or U4919 (N_4919,N_4360,N_4001);
nand U4920 (N_4920,N_4454,N_4266);
nor U4921 (N_4921,N_4428,N_3905);
nor U4922 (N_4922,N_3911,N_4125);
nand U4923 (N_4923,N_4020,N_4285);
nor U4924 (N_4924,N_4059,N_4094);
nor U4925 (N_4925,N_4192,N_3934);
nand U4926 (N_4926,N_4030,N_4045);
nand U4927 (N_4927,N_3840,N_4378);
nor U4928 (N_4928,N_4462,N_3875);
nor U4929 (N_4929,N_3870,N_4140);
nand U4930 (N_4930,N_4148,N_4341);
nand U4931 (N_4931,N_4047,N_4212);
and U4932 (N_4932,N_4316,N_3863);
nor U4933 (N_4933,N_4170,N_3890);
nand U4934 (N_4934,N_3873,N_3984);
and U4935 (N_4935,N_4138,N_3992);
nand U4936 (N_4936,N_4136,N_4478);
or U4937 (N_4937,N_3853,N_4361);
or U4938 (N_4938,N_4139,N_4045);
nor U4939 (N_4939,N_3885,N_3864);
nand U4940 (N_4940,N_4049,N_4484);
nor U4941 (N_4941,N_4077,N_4499);
xor U4942 (N_4942,N_4329,N_3759);
nor U4943 (N_4943,N_4427,N_3756);
or U4944 (N_4944,N_3820,N_4261);
nand U4945 (N_4945,N_3865,N_3948);
or U4946 (N_4946,N_4257,N_3900);
or U4947 (N_4947,N_4140,N_3856);
nand U4948 (N_4948,N_4194,N_4309);
or U4949 (N_4949,N_4259,N_4083);
or U4950 (N_4950,N_3967,N_4455);
nor U4951 (N_4951,N_3929,N_3816);
or U4952 (N_4952,N_4322,N_4365);
nor U4953 (N_4953,N_4081,N_3959);
and U4954 (N_4954,N_4034,N_3909);
nor U4955 (N_4955,N_3839,N_3797);
or U4956 (N_4956,N_4448,N_4110);
or U4957 (N_4957,N_4107,N_4337);
nand U4958 (N_4958,N_4359,N_3810);
nor U4959 (N_4959,N_3917,N_3970);
and U4960 (N_4960,N_3860,N_4388);
nor U4961 (N_4961,N_4445,N_3890);
nand U4962 (N_4962,N_4491,N_3873);
nand U4963 (N_4963,N_4366,N_4143);
and U4964 (N_4964,N_4413,N_4448);
and U4965 (N_4965,N_4498,N_4405);
and U4966 (N_4966,N_4165,N_4467);
or U4967 (N_4967,N_3962,N_3904);
or U4968 (N_4968,N_4269,N_4285);
nand U4969 (N_4969,N_4427,N_4122);
and U4970 (N_4970,N_3928,N_4191);
or U4971 (N_4971,N_4350,N_4354);
or U4972 (N_4972,N_4478,N_4053);
nand U4973 (N_4973,N_4408,N_4352);
or U4974 (N_4974,N_3847,N_4083);
and U4975 (N_4975,N_3771,N_4220);
nand U4976 (N_4976,N_4327,N_4194);
and U4977 (N_4977,N_3958,N_4367);
or U4978 (N_4978,N_4433,N_4019);
nand U4979 (N_4979,N_4429,N_4476);
or U4980 (N_4980,N_4078,N_4250);
or U4981 (N_4981,N_4362,N_3878);
nor U4982 (N_4982,N_3770,N_3922);
and U4983 (N_4983,N_3958,N_3966);
xnor U4984 (N_4984,N_4189,N_4241);
nand U4985 (N_4985,N_4318,N_3925);
nand U4986 (N_4986,N_4048,N_4147);
nand U4987 (N_4987,N_3811,N_3912);
nand U4988 (N_4988,N_3844,N_3951);
or U4989 (N_4989,N_3810,N_4435);
xor U4990 (N_4990,N_4147,N_4404);
and U4991 (N_4991,N_4455,N_4498);
nand U4992 (N_4992,N_4443,N_4415);
nor U4993 (N_4993,N_3969,N_3984);
or U4994 (N_4994,N_3825,N_4473);
nor U4995 (N_4995,N_4169,N_4017);
nand U4996 (N_4996,N_3861,N_4268);
nor U4997 (N_4997,N_3891,N_4477);
nand U4998 (N_4998,N_3875,N_4242);
or U4999 (N_4999,N_4106,N_4192);
nand U5000 (N_5000,N_4413,N_4014);
and U5001 (N_5001,N_4031,N_4230);
and U5002 (N_5002,N_3761,N_4253);
nand U5003 (N_5003,N_4251,N_3869);
and U5004 (N_5004,N_4073,N_4124);
or U5005 (N_5005,N_4211,N_3798);
and U5006 (N_5006,N_4159,N_4498);
nor U5007 (N_5007,N_4149,N_4315);
nor U5008 (N_5008,N_3789,N_4027);
or U5009 (N_5009,N_3900,N_4117);
nor U5010 (N_5010,N_4310,N_3966);
nand U5011 (N_5011,N_4320,N_4104);
nand U5012 (N_5012,N_4111,N_4474);
and U5013 (N_5013,N_3822,N_4067);
and U5014 (N_5014,N_3878,N_3767);
and U5015 (N_5015,N_3913,N_4226);
nor U5016 (N_5016,N_4264,N_4159);
nor U5017 (N_5017,N_4130,N_4087);
or U5018 (N_5018,N_4474,N_3835);
nor U5019 (N_5019,N_3802,N_3941);
and U5020 (N_5020,N_4420,N_4049);
and U5021 (N_5021,N_4071,N_3831);
nand U5022 (N_5022,N_4334,N_4152);
xor U5023 (N_5023,N_4252,N_3800);
nand U5024 (N_5024,N_3916,N_4231);
or U5025 (N_5025,N_4044,N_4477);
and U5026 (N_5026,N_3794,N_4459);
nand U5027 (N_5027,N_4022,N_4225);
or U5028 (N_5028,N_3861,N_3889);
nor U5029 (N_5029,N_3869,N_3806);
nand U5030 (N_5030,N_3920,N_4103);
and U5031 (N_5031,N_3945,N_4475);
nor U5032 (N_5032,N_4063,N_3980);
and U5033 (N_5033,N_3752,N_4262);
and U5034 (N_5034,N_4409,N_4461);
and U5035 (N_5035,N_4419,N_3818);
nor U5036 (N_5036,N_4020,N_4198);
nand U5037 (N_5037,N_3916,N_4178);
nor U5038 (N_5038,N_3868,N_4198);
nor U5039 (N_5039,N_4267,N_4016);
nor U5040 (N_5040,N_3895,N_4299);
nor U5041 (N_5041,N_4465,N_4091);
or U5042 (N_5042,N_4206,N_4345);
and U5043 (N_5043,N_4118,N_3809);
and U5044 (N_5044,N_3756,N_4304);
and U5045 (N_5045,N_3862,N_3961);
or U5046 (N_5046,N_4084,N_4019);
or U5047 (N_5047,N_4305,N_4265);
and U5048 (N_5048,N_4263,N_3985);
or U5049 (N_5049,N_3802,N_4324);
nand U5050 (N_5050,N_4327,N_3990);
or U5051 (N_5051,N_4064,N_4059);
or U5052 (N_5052,N_3916,N_4027);
nor U5053 (N_5053,N_4063,N_4193);
nor U5054 (N_5054,N_4150,N_4406);
and U5055 (N_5055,N_4085,N_4182);
and U5056 (N_5056,N_4183,N_4243);
nand U5057 (N_5057,N_4182,N_4462);
xnor U5058 (N_5058,N_4304,N_4483);
and U5059 (N_5059,N_4129,N_3972);
nand U5060 (N_5060,N_4421,N_4156);
or U5061 (N_5061,N_4060,N_3988);
and U5062 (N_5062,N_4472,N_3964);
and U5063 (N_5063,N_4403,N_3798);
and U5064 (N_5064,N_3764,N_4416);
nor U5065 (N_5065,N_4402,N_3771);
nor U5066 (N_5066,N_4367,N_4228);
nand U5067 (N_5067,N_3839,N_4038);
and U5068 (N_5068,N_4499,N_4183);
or U5069 (N_5069,N_4118,N_3984);
and U5070 (N_5070,N_3765,N_4422);
and U5071 (N_5071,N_4014,N_4132);
or U5072 (N_5072,N_4122,N_4013);
nor U5073 (N_5073,N_4244,N_3811);
nor U5074 (N_5074,N_4280,N_4485);
xor U5075 (N_5075,N_4007,N_4199);
or U5076 (N_5076,N_4342,N_4163);
nand U5077 (N_5077,N_4083,N_3831);
and U5078 (N_5078,N_4018,N_4192);
or U5079 (N_5079,N_4335,N_4025);
and U5080 (N_5080,N_4291,N_4367);
nor U5081 (N_5081,N_4174,N_3932);
nand U5082 (N_5082,N_3758,N_4223);
nor U5083 (N_5083,N_4406,N_3775);
and U5084 (N_5084,N_3820,N_3927);
and U5085 (N_5085,N_4306,N_4373);
and U5086 (N_5086,N_3895,N_3887);
nand U5087 (N_5087,N_4287,N_4242);
nor U5088 (N_5088,N_3896,N_4243);
and U5089 (N_5089,N_3760,N_4345);
nor U5090 (N_5090,N_4098,N_4307);
and U5091 (N_5091,N_4233,N_4269);
nand U5092 (N_5092,N_4471,N_4425);
nor U5093 (N_5093,N_3956,N_4048);
nand U5094 (N_5094,N_4262,N_4068);
and U5095 (N_5095,N_4263,N_4388);
or U5096 (N_5096,N_3935,N_4021);
and U5097 (N_5097,N_4498,N_4458);
nand U5098 (N_5098,N_4083,N_4043);
xnor U5099 (N_5099,N_4170,N_4337);
nor U5100 (N_5100,N_4373,N_4269);
nand U5101 (N_5101,N_4170,N_4387);
nor U5102 (N_5102,N_4156,N_4328);
or U5103 (N_5103,N_3770,N_4165);
nand U5104 (N_5104,N_4262,N_3814);
nor U5105 (N_5105,N_4198,N_3912);
or U5106 (N_5106,N_4468,N_3851);
nor U5107 (N_5107,N_4161,N_4242);
and U5108 (N_5108,N_3771,N_3878);
nor U5109 (N_5109,N_4027,N_4113);
or U5110 (N_5110,N_3817,N_3872);
and U5111 (N_5111,N_4116,N_4151);
and U5112 (N_5112,N_4402,N_4011);
nand U5113 (N_5113,N_3969,N_3806);
nor U5114 (N_5114,N_4128,N_4113);
and U5115 (N_5115,N_4028,N_4259);
and U5116 (N_5116,N_3949,N_3830);
and U5117 (N_5117,N_4073,N_3825);
nand U5118 (N_5118,N_3960,N_4302);
and U5119 (N_5119,N_3935,N_3758);
and U5120 (N_5120,N_3786,N_4019);
xor U5121 (N_5121,N_3982,N_4024);
and U5122 (N_5122,N_3830,N_4461);
nand U5123 (N_5123,N_3873,N_4309);
nand U5124 (N_5124,N_4095,N_4259);
nor U5125 (N_5125,N_3822,N_4095);
nand U5126 (N_5126,N_4393,N_4373);
nor U5127 (N_5127,N_3877,N_4285);
or U5128 (N_5128,N_4037,N_4395);
nor U5129 (N_5129,N_3998,N_3818);
nand U5130 (N_5130,N_4043,N_4349);
nor U5131 (N_5131,N_4435,N_4322);
and U5132 (N_5132,N_4460,N_3838);
xnor U5133 (N_5133,N_4173,N_4196);
or U5134 (N_5134,N_4383,N_4156);
and U5135 (N_5135,N_4114,N_3825);
and U5136 (N_5136,N_4090,N_3809);
nand U5137 (N_5137,N_4112,N_4090);
and U5138 (N_5138,N_4257,N_3784);
nor U5139 (N_5139,N_4058,N_4438);
nand U5140 (N_5140,N_4464,N_3821);
or U5141 (N_5141,N_4441,N_4450);
nand U5142 (N_5142,N_4257,N_4485);
and U5143 (N_5143,N_3923,N_3866);
and U5144 (N_5144,N_3799,N_3976);
and U5145 (N_5145,N_4045,N_3882);
and U5146 (N_5146,N_3779,N_4254);
nand U5147 (N_5147,N_3762,N_4481);
nor U5148 (N_5148,N_3777,N_4106);
nor U5149 (N_5149,N_4361,N_3982);
nand U5150 (N_5150,N_4053,N_3841);
nor U5151 (N_5151,N_4440,N_4005);
nand U5152 (N_5152,N_3837,N_4081);
and U5153 (N_5153,N_4099,N_3883);
nand U5154 (N_5154,N_3758,N_4490);
nand U5155 (N_5155,N_4021,N_4014);
and U5156 (N_5156,N_4224,N_4380);
and U5157 (N_5157,N_3912,N_4441);
or U5158 (N_5158,N_4277,N_4034);
or U5159 (N_5159,N_4095,N_4103);
nand U5160 (N_5160,N_4022,N_3996);
nor U5161 (N_5161,N_4341,N_4038);
and U5162 (N_5162,N_3857,N_4418);
and U5163 (N_5163,N_4260,N_3882);
nand U5164 (N_5164,N_4301,N_4097);
nor U5165 (N_5165,N_4301,N_4061);
nor U5166 (N_5166,N_4034,N_4322);
nand U5167 (N_5167,N_3899,N_4001);
nor U5168 (N_5168,N_3760,N_3908);
nand U5169 (N_5169,N_4095,N_4045);
nor U5170 (N_5170,N_4179,N_4056);
or U5171 (N_5171,N_3845,N_3843);
or U5172 (N_5172,N_4420,N_4479);
or U5173 (N_5173,N_3767,N_4432);
nand U5174 (N_5174,N_4106,N_3758);
nor U5175 (N_5175,N_4038,N_4245);
xor U5176 (N_5176,N_3822,N_4250);
nor U5177 (N_5177,N_4170,N_3888);
nor U5178 (N_5178,N_3855,N_4402);
and U5179 (N_5179,N_4399,N_3772);
and U5180 (N_5180,N_4203,N_4254);
nand U5181 (N_5181,N_4470,N_4407);
nor U5182 (N_5182,N_4193,N_4333);
or U5183 (N_5183,N_3967,N_3998);
nor U5184 (N_5184,N_4113,N_4173);
or U5185 (N_5185,N_4047,N_4185);
nand U5186 (N_5186,N_4276,N_4203);
and U5187 (N_5187,N_3923,N_3962);
nor U5188 (N_5188,N_4211,N_4175);
nand U5189 (N_5189,N_4052,N_4197);
nand U5190 (N_5190,N_4175,N_4342);
and U5191 (N_5191,N_4457,N_4207);
nand U5192 (N_5192,N_4424,N_4435);
nor U5193 (N_5193,N_4005,N_3891);
and U5194 (N_5194,N_4249,N_4197);
or U5195 (N_5195,N_3932,N_4355);
nor U5196 (N_5196,N_3778,N_4332);
or U5197 (N_5197,N_4165,N_4292);
nor U5198 (N_5198,N_4463,N_3993);
nor U5199 (N_5199,N_4292,N_4034);
and U5200 (N_5200,N_3751,N_4243);
and U5201 (N_5201,N_4370,N_4259);
nand U5202 (N_5202,N_3951,N_4200);
nand U5203 (N_5203,N_4110,N_4365);
nor U5204 (N_5204,N_4420,N_4070);
nand U5205 (N_5205,N_4320,N_3928);
and U5206 (N_5206,N_3874,N_4183);
nor U5207 (N_5207,N_4347,N_3941);
and U5208 (N_5208,N_4197,N_4260);
nand U5209 (N_5209,N_4422,N_4445);
nand U5210 (N_5210,N_3877,N_4034);
nor U5211 (N_5211,N_3942,N_4285);
nor U5212 (N_5212,N_3975,N_4218);
and U5213 (N_5213,N_4437,N_3851);
or U5214 (N_5214,N_4103,N_3817);
and U5215 (N_5215,N_4202,N_4257);
or U5216 (N_5216,N_4245,N_4045);
nor U5217 (N_5217,N_3750,N_4240);
nand U5218 (N_5218,N_4004,N_4391);
or U5219 (N_5219,N_3809,N_4236);
nor U5220 (N_5220,N_3766,N_4312);
nand U5221 (N_5221,N_4182,N_4194);
and U5222 (N_5222,N_4467,N_4129);
nand U5223 (N_5223,N_4409,N_4339);
nand U5224 (N_5224,N_3773,N_4421);
nor U5225 (N_5225,N_4367,N_3754);
or U5226 (N_5226,N_4129,N_4254);
nand U5227 (N_5227,N_4173,N_4096);
and U5228 (N_5228,N_3927,N_4088);
nor U5229 (N_5229,N_4019,N_4069);
nor U5230 (N_5230,N_4370,N_4034);
and U5231 (N_5231,N_3750,N_3821);
nand U5232 (N_5232,N_4287,N_4381);
xor U5233 (N_5233,N_4261,N_3856);
or U5234 (N_5234,N_4345,N_3842);
nand U5235 (N_5235,N_4041,N_4492);
or U5236 (N_5236,N_4451,N_3868);
and U5237 (N_5237,N_4476,N_3897);
nand U5238 (N_5238,N_4087,N_4098);
or U5239 (N_5239,N_4119,N_4207);
and U5240 (N_5240,N_4415,N_4316);
nor U5241 (N_5241,N_4326,N_4259);
xor U5242 (N_5242,N_4163,N_3818);
or U5243 (N_5243,N_4264,N_4416);
or U5244 (N_5244,N_4260,N_4491);
nor U5245 (N_5245,N_4382,N_4494);
and U5246 (N_5246,N_3929,N_4311);
and U5247 (N_5247,N_4062,N_4073);
xor U5248 (N_5248,N_3790,N_3857);
or U5249 (N_5249,N_4205,N_4105);
and U5250 (N_5250,N_5034,N_4863);
and U5251 (N_5251,N_4789,N_4775);
or U5252 (N_5252,N_4866,N_5045);
and U5253 (N_5253,N_4677,N_4714);
nand U5254 (N_5254,N_4596,N_5191);
and U5255 (N_5255,N_4826,N_4962);
xnor U5256 (N_5256,N_4629,N_4665);
nand U5257 (N_5257,N_5136,N_5100);
nand U5258 (N_5258,N_4529,N_4817);
nor U5259 (N_5259,N_5149,N_4813);
nand U5260 (N_5260,N_5108,N_4907);
and U5261 (N_5261,N_4965,N_4786);
nand U5262 (N_5262,N_4883,N_5084);
nor U5263 (N_5263,N_5031,N_5114);
nand U5264 (N_5264,N_4622,N_4741);
nor U5265 (N_5265,N_5088,N_5003);
and U5266 (N_5266,N_4570,N_5197);
nand U5267 (N_5267,N_5247,N_4598);
nor U5268 (N_5268,N_4824,N_5192);
nand U5269 (N_5269,N_4545,N_4736);
xnor U5270 (N_5270,N_4502,N_4692);
or U5271 (N_5271,N_5015,N_5023);
and U5272 (N_5272,N_5182,N_4788);
or U5273 (N_5273,N_4847,N_4891);
nor U5274 (N_5274,N_4770,N_4902);
and U5275 (N_5275,N_4657,N_5041);
or U5276 (N_5276,N_5178,N_4509);
or U5277 (N_5277,N_4604,N_5081);
and U5278 (N_5278,N_4553,N_4676);
or U5279 (N_5279,N_4758,N_4739);
nand U5280 (N_5280,N_4892,N_5086);
or U5281 (N_5281,N_4681,N_4840);
nor U5282 (N_5282,N_5121,N_4979);
nor U5283 (N_5283,N_4548,N_5133);
nand U5284 (N_5284,N_5066,N_4627);
nand U5285 (N_5285,N_4594,N_5240);
xor U5286 (N_5286,N_4790,N_4765);
or U5287 (N_5287,N_5189,N_4887);
and U5288 (N_5288,N_4792,N_5057);
or U5289 (N_5289,N_4696,N_4998);
and U5290 (N_5290,N_5026,N_5172);
nand U5291 (N_5291,N_5190,N_5120);
nand U5292 (N_5292,N_4935,N_4514);
and U5293 (N_5293,N_5028,N_4833);
and U5294 (N_5294,N_5225,N_4601);
nor U5295 (N_5295,N_5193,N_5201);
nand U5296 (N_5296,N_4724,N_4787);
nand U5297 (N_5297,N_4993,N_4726);
and U5298 (N_5298,N_4712,N_4874);
or U5299 (N_5299,N_4649,N_5165);
nand U5300 (N_5300,N_4504,N_4723);
nand U5301 (N_5301,N_4635,N_4842);
nand U5302 (N_5302,N_5082,N_4720);
and U5303 (N_5303,N_4513,N_4803);
nand U5304 (N_5304,N_5221,N_5228);
and U5305 (N_5305,N_4701,N_4634);
nand U5306 (N_5306,N_4631,N_4961);
and U5307 (N_5307,N_5118,N_5224);
and U5308 (N_5308,N_4898,N_4808);
or U5309 (N_5309,N_4702,N_5176);
and U5310 (N_5310,N_4688,N_4507);
nand U5311 (N_5311,N_4849,N_5127);
or U5312 (N_5312,N_5206,N_4869);
nand U5313 (N_5313,N_5115,N_4916);
nand U5314 (N_5314,N_4919,N_5154);
nand U5315 (N_5315,N_5142,N_4825);
nor U5316 (N_5316,N_4949,N_4515);
nor U5317 (N_5317,N_4872,N_5239);
nor U5318 (N_5318,N_4621,N_5187);
nand U5319 (N_5319,N_4839,N_4699);
nor U5320 (N_5320,N_4587,N_4953);
nand U5321 (N_5321,N_4615,N_4608);
and U5322 (N_5322,N_5113,N_4603);
and U5323 (N_5323,N_5055,N_5091);
nor U5324 (N_5324,N_4865,N_4917);
or U5325 (N_5325,N_4547,N_4915);
nand U5326 (N_5326,N_5242,N_5029);
nand U5327 (N_5327,N_5020,N_4695);
nand U5328 (N_5328,N_5185,N_4988);
and U5329 (N_5329,N_4828,N_5156);
nor U5330 (N_5330,N_5032,N_4894);
nand U5331 (N_5331,N_5148,N_5209);
nand U5332 (N_5332,N_4805,N_4607);
xnor U5333 (N_5333,N_5202,N_4852);
or U5334 (N_5334,N_4855,N_4745);
and U5335 (N_5335,N_4815,N_4936);
nand U5336 (N_5336,N_4801,N_4860);
and U5337 (N_5337,N_4749,N_5038);
nor U5338 (N_5338,N_5013,N_4862);
and U5339 (N_5339,N_5109,N_4997);
nor U5340 (N_5340,N_4861,N_5203);
nand U5341 (N_5341,N_5128,N_5174);
nand U5342 (N_5342,N_5147,N_4644);
nand U5343 (N_5343,N_4523,N_4811);
nor U5344 (N_5344,N_4734,N_5137);
nor U5345 (N_5345,N_5145,N_4978);
or U5346 (N_5346,N_5094,N_4595);
nor U5347 (N_5347,N_5087,N_4882);
nand U5348 (N_5348,N_4572,N_4776);
or U5349 (N_5349,N_4851,N_4521);
nor U5350 (N_5350,N_5179,N_4777);
or U5351 (N_5351,N_4571,N_5162);
nand U5352 (N_5352,N_5143,N_4531);
nand U5353 (N_5353,N_5076,N_4864);
nand U5354 (N_5354,N_5073,N_4686);
nor U5355 (N_5355,N_4643,N_4633);
nor U5356 (N_5356,N_4886,N_4524);
and U5357 (N_5357,N_4551,N_4605);
and U5358 (N_5358,N_4698,N_4810);
or U5359 (N_5359,N_4556,N_4655);
nand U5360 (N_5360,N_4654,N_5208);
nor U5361 (N_5361,N_5213,N_5093);
nor U5362 (N_5362,N_4857,N_4667);
nand U5363 (N_5363,N_4592,N_4661);
nand U5364 (N_5364,N_5096,N_4975);
and U5365 (N_5365,N_4967,N_5047);
or U5366 (N_5366,N_5204,N_4602);
xnor U5367 (N_5367,N_5234,N_5027);
or U5368 (N_5368,N_4517,N_4818);
nand U5369 (N_5369,N_5233,N_4672);
and U5370 (N_5370,N_4729,N_5144);
nor U5371 (N_5371,N_5021,N_4740);
or U5372 (N_5372,N_4500,N_5004);
and U5373 (N_5373,N_4530,N_4853);
nand U5374 (N_5374,N_4926,N_5188);
nor U5375 (N_5375,N_4518,N_4744);
xor U5376 (N_5376,N_4774,N_4573);
or U5377 (N_5377,N_4673,N_4870);
or U5378 (N_5378,N_4728,N_4831);
nor U5379 (N_5379,N_4766,N_4632);
or U5380 (N_5380,N_4558,N_5155);
and U5381 (N_5381,N_5069,N_4911);
xnor U5382 (N_5382,N_4799,N_4528);
nand U5383 (N_5383,N_5006,N_4837);
nand U5384 (N_5384,N_4893,N_5037);
nand U5385 (N_5385,N_4793,N_4683);
and U5386 (N_5386,N_4945,N_4764);
nand U5387 (N_5387,N_4568,N_4954);
nand U5388 (N_5388,N_4501,N_4536);
nand U5389 (N_5389,N_4956,N_4611);
or U5390 (N_5390,N_5060,N_5195);
nor U5391 (N_5391,N_5241,N_4743);
or U5392 (N_5392,N_5227,N_5077);
nand U5393 (N_5393,N_5150,N_4964);
nand U5394 (N_5394,N_4854,N_4832);
or U5395 (N_5395,N_4938,N_5001);
and U5396 (N_5396,N_4829,N_4693);
or U5397 (N_5397,N_5070,N_5168);
and U5398 (N_5398,N_4779,N_4640);
nor U5399 (N_5399,N_5175,N_4848);
or U5400 (N_5400,N_4559,N_4981);
nor U5401 (N_5401,N_4951,N_4535);
nor U5402 (N_5402,N_5033,N_4700);
and U5403 (N_5403,N_4760,N_4527);
nand U5404 (N_5404,N_5056,N_4983);
or U5405 (N_5405,N_4538,N_4576);
nor U5406 (N_5406,N_4966,N_5123);
nand U5407 (N_5407,N_4580,N_4973);
and U5408 (N_5408,N_4735,N_4952);
and U5409 (N_5409,N_4922,N_5092);
nand U5410 (N_5410,N_4880,N_5223);
or U5411 (N_5411,N_4526,N_5078);
nor U5412 (N_5412,N_4985,N_4937);
and U5413 (N_5413,N_4694,N_4947);
nor U5414 (N_5414,N_5152,N_4540);
nor U5415 (N_5415,N_4708,N_4843);
nand U5416 (N_5416,N_4890,N_4913);
nor U5417 (N_5417,N_5217,N_4543);
and U5418 (N_5418,N_4606,N_4617);
nor U5419 (N_5419,N_4550,N_4943);
xnor U5420 (N_5420,N_4946,N_4995);
and U5421 (N_5421,N_4583,N_4958);
and U5422 (N_5422,N_5124,N_5009);
and U5423 (N_5423,N_5141,N_4940);
nand U5424 (N_5424,N_5072,N_5160);
xnor U5425 (N_5425,N_4955,N_5181);
and U5426 (N_5426,N_5059,N_4679);
nand U5427 (N_5427,N_4999,N_4822);
or U5428 (N_5428,N_4960,N_4932);
nor U5429 (N_5429,N_4845,N_4821);
nand U5430 (N_5430,N_5043,N_4508);
nor U5431 (N_5431,N_4616,N_5122);
nand U5432 (N_5432,N_4650,N_4578);
nor U5433 (N_5433,N_4563,N_4641);
and U5434 (N_5434,N_4674,N_5132);
nor U5435 (N_5435,N_5210,N_4669);
xor U5436 (N_5436,N_4838,N_4612);
or U5437 (N_5437,N_4511,N_4969);
nand U5438 (N_5438,N_4706,N_4888);
and U5439 (N_5439,N_5157,N_4727);
nor U5440 (N_5440,N_4647,N_4668);
nand U5441 (N_5441,N_4546,N_4948);
or U5442 (N_5442,N_5139,N_4586);
or U5443 (N_5443,N_5130,N_5112);
or U5444 (N_5444,N_5110,N_4769);
nor U5445 (N_5445,N_4797,N_4772);
nand U5446 (N_5446,N_4533,N_4780);
or U5447 (N_5447,N_4717,N_4972);
nor U5448 (N_5448,N_4755,N_4625);
and U5449 (N_5449,N_4812,N_4889);
or U5450 (N_5450,N_5039,N_4737);
and U5451 (N_5451,N_5211,N_4980);
nand U5452 (N_5452,N_4957,N_4623);
or U5453 (N_5453,N_5198,N_5207);
and U5454 (N_5454,N_4747,N_5177);
nand U5455 (N_5455,N_4512,N_4597);
nor U5456 (N_5456,N_5062,N_4703);
or U5457 (N_5457,N_5054,N_4516);
nand U5458 (N_5458,N_4850,N_4575);
nand U5459 (N_5459,N_4711,N_4716);
or U5460 (N_5460,N_4505,N_4930);
nand U5461 (N_5461,N_4705,N_4564);
and U5462 (N_5462,N_4784,N_5249);
or U5463 (N_5463,N_4900,N_5111);
nand U5464 (N_5464,N_5117,N_4732);
and U5465 (N_5465,N_4725,N_4794);
nand U5466 (N_5466,N_5102,N_5010);
and U5467 (N_5467,N_4549,N_5017);
or U5468 (N_5468,N_5105,N_5216);
and U5469 (N_5469,N_4544,N_5083);
nor U5470 (N_5470,N_4816,N_5245);
nand U5471 (N_5471,N_5237,N_4555);
nor U5472 (N_5472,N_4520,N_4925);
nand U5473 (N_5473,N_5158,N_4798);
nor U5474 (N_5474,N_4722,N_5166);
nand U5475 (N_5475,N_5229,N_5050);
or U5476 (N_5476,N_4820,N_5097);
and U5477 (N_5477,N_4684,N_5061);
or U5478 (N_5478,N_5014,N_4614);
and U5479 (N_5479,N_4680,N_5226);
nor U5480 (N_5480,N_4778,N_5095);
nand U5481 (N_5481,N_5186,N_4748);
and U5482 (N_5482,N_5135,N_4773);
nor U5483 (N_5483,N_4678,N_5184);
or U5484 (N_5484,N_4600,N_4942);
nand U5485 (N_5485,N_5074,N_4590);
and U5486 (N_5486,N_4675,N_5214);
nand U5487 (N_5487,N_4918,N_4809);
nor U5488 (N_5488,N_4991,N_4934);
nor U5489 (N_5489,N_5212,N_4565);
nor U5490 (N_5490,N_4931,N_5008);
or U5491 (N_5491,N_4613,N_5067);
nor U5492 (N_5492,N_5196,N_5053);
nor U5493 (N_5493,N_4519,N_5035);
and U5494 (N_5494,N_5146,N_5243);
nand U5495 (N_5495,N_5180,N_5119);
nand U5496 (N_5496,N_5002,N_4620);
or U5497 (N_5497,N_5071,N_4933);
nand U5498 (N_5498,N_5171,N_4733);
nor U5499 (N_5499,N_5220,N_4771);
or U5500 (N_5500,N_4658,N_4731);
nand U5501 (N_5501,N_4835,N_4992);
nand U5502 (N_5502,N_4582,N_4690);
and U5503 (N_5503,N_4532,N_5131);
or U5504 (N_5504,N_4626,N_5005);
and U5505 (N_5505,N_4841,N_5215);
nor U5506 (N_5506,N_5246,N_4730);
nor U5507 (N_5507,N_5051,N_4867);
and U5508 (N_5508,N_4687,N_4567);
and U5509 (N_5509,N_4920,N_4762);
and U5510 (N_5510,N_4871,N_4796);
nand U5511 (N_5511,N_4539,N_4989);
nand U5512 (N_5512,N_4659,N_5248);
or U5513 (N_5513,N_4827,N_4908);
nor U5514 (N_5514,N_4795,N_5000);
nand U5515 (N_5515,N_4697,N_4753);
nand U5516 (N_5516,N_4782,N_5089);
nor U5517 (N_5517,N_5183,N_4971);
nand U5518 (N_5518,N_4651,N_4719);
nor U5519 (N_5519,N_4987,N_4858);
nor U5520 (N_5520,N_4944,N_4904);
or U5521 (N_5521,N_5104,N_4646);
and U5522 (N_5522,N_5194,N_4666);
xnor U5523 (N_5523,N_4856,N_5164);
and U5524 (N_5524,N_4763,N_4588);
nor U5525 (N_5525,N_4756,N_4976);
nand U5526 (N_5526,N_5064,N_5238);
and U5527 (N_5527,N_5219,N_5036);
or U5528 (N_5528,N_4912,N_4653);
nor U5529 (N_5529,N_4767,N_4802);
or U5530 (N_5530,N_4759,N_4639);
xnor U5531 (N_5531,N_4721,N_5065);
or U5532 (N_5532,N_4844,N_4868);
or U5533 (N_5533,N_4791,N_5151);
and U5534 (N_5534,N_5163,N_5048);
nor U5535 (N_5535,N_4859,N_4591);
and U5536 (N_5536,N_5058,N_5140);
nand U5537 (N_5537,N_4897,N_5103);
and U5538 (N_5538,N_4990,N_4662);
and U5539 (N_5539,N_4636,N_4645);
nor U5540 (N_5540,N_4846,N_5046);
nor U5541 (N_5541,N_5199,N_4746);
nand U5542 (N_5542,N_4610,N_4814);
nor U5543 (N_5543,N_4879,N_5080);
or U5544 (N_5544,N_4510,N_4609);
or U5545 (N_5545,N_4671,N_4781);
and U5546 (N_5546,N_4750,N_4878);
and U5547 (N_5547,N_5159,N_4977);
and U5548 (N_5548,N_5244,N_4618);
nand U5549 (N_5549,N_4910,N_4642);
or U5550 (N_5550,N_4589,N_4986);
nand U5551 (N_5551,N_4909,N_4819);
nand U5552 (N_5552,N_4941,N_4823);
nand U5553 (N_5553,N_4566,N_5012);
or U5554 (N_5554,N_4785,N_4994);
or U5555 (N_5555,N_4921,N_5235);
nand U5556 (N_5556,N_4877,N_4561);
nor U5557 (N_5557,N_5232,N_4619);
or U5558 (N_5558,N_4709,N_5101);
nand U5559 (N_5559,N_4542,N_5205);
or U5560 (N_5560,N_4836,N_4710);
and U5561 (N_5561,N_4593,N_5098);
nand U5562 (N_5562,N_5231,N_5011);
and U5563 (N_5563,N_5099,N_5018);
nor U5564 (N_5564,N_4939,N_5170);
nand U5565 (N_5565,N_5218,N_4577);
nand U5566 (N_5566,N_4670,N_4638);
nand U5567 (N_5567,N_4534,N_5236);
nor U5568 (N_5568,N_4761,N_4599);
nor U5569 (N_5569,N_4968,N_4884);
xnor U5570 (N_5570,N_4503,N_4574);
or U5571 (N_5571,N_4682,N_4982);
and U5572 (N_5572,N_4876,N_5019);
and U5573 (N_5573,N_4704,N_5090);
and U5574 (N_5574,N_4685,N_4751);
and U5575 (N_5575,N_4664,N_5052);
and U5576 (N_5576,N_4901,N_4974);
and U5577 (N_5577,N_4754,N_4660);
or U5578 (N_5578,N_4560,N_4924);
or U5579 (N_5579,N_4637,N_4885);
nand U5580 (N_5580,N_4624,N_4738);
nor U5581 (N_5581,N_4807,N_4914);
or U5582 (N_5582,N_4630,N_5063);
nor U5583 (N_5583,N_4928,N_5126);
and U5584 (N_5584,N_5022,N_5025);
nor U5585 (N_5585,N_4691,N_4707);
or U5586 (N_5586,N_5125,N_5106);
or U5587 (N_5587,N_5042,N_4895);
nor U5588 (N_5588,N_4896,N_5116);
nor U5589 (N_5589,N_4929,N_4984);
xor U5590 (N_5590,N_4800,N_5167);
nand U5591 (N_5591,N_4742,N_5075);
nor U5592 (N_5592,N_5153,N_4873);
nand U5593 (N_5593,N_4628,N_4713);
and U5594 (N_5594,N_4875,N_4522);
nand U5595 (N_5595,N_4554,N_5169);
and U5596 (N_5596,N_5129,N_4584);
nor U5597 (N_5597,N_5085,N_5007);
and U5598 (N_5598,N_4585,N_5134);
nor U5599 (N_5599,N_4950,N_4541);
or U5600 (N_5600,N_4579,N_4537);
nor U5601 (N_5601,N_4569,N_5138);
nand U5602 (N_5602,N_4689,N_4881);
and U5603 (N_5603,N_4562,N_4834);
nor U5604 (N_5604,N_4768,N_4648);
nor U5605 (N_5605,N_4757,N_5049);
nor U5606 (N_5606,N_4552,N_4903);
or U5607 (N_5607,N_4656,N_4752);
nand U5608 (N_5608,N_5222,N_5040);
nor U5609 (N_5609,N_4959,N_4927);
and U5610 (N_5610,N_4963,N_4923);
nor U5611 (N_5611,N_5200,N_5161);
or U5612 (N_5612,N_4830,N_4506);
nor U5613 (N_5613,N_5024,N_4906);
or U5614 (N_5614,N_4525,N_4652);
xor U5615 (N_5615,N_4718,N_4970);
nor U5616 (N_5616,N_4804,N_4905);
and U5617 (N_5617,N_4806,N_5068);
and U5618 (N_5618,N_5044,N_5030);
and U5619 (N_5619,N_4557,N_4663);
nand U5620 (N_5620,N_4581,N_5079);
nand U5621 (N_5621,N_4783,N_4996);
nand U5622 (N_5622,N_5016,N_5230);
or U5623 (N_5623,N_4715,N_4899);
and U5624 (N_5624,N_5107,N_5173);
nor U5625 (N_5625,N_4772,N_5130);
nor U5626 (N_5626,N_4540,N_4763);
nand U5627 (N_5627,N_5152,N_4719);
or U5628 (N_5628,N_4630,N_4604);
nor U5629 (N_5629,N_5091,N_4534);
or U5630 (N_5630,N_5110,N_5199);
and U5631 (N_5631,N_4921,N_5188);
nor U5632 (N_5632,N_5002,N_4529);
nand U5633 (N_5633,N_4998,N_5067);
nor U5634 (N_5634,N_4879,N_4942);
nand U5635 (N_5635,N_5147,N_5175);
nor U5636 (N_5636,N_4694,N_4776);
nand U5637 (N_5637,N_5203,N_5103);
or U5638 (N_5638,N_5023,N_4937);
nand U5639 (N_5639,N_4963,N_4798);
nand U5640 (N_5640,N_5118,N_4806);
nand U5641 (N_5641,N_4663,N_5073);
nand U5642 (N_5642,N_4701,N_4616);
and U5643 (N_5643,N_4734,N_4832);
nor U5644 (N_5644,N_4819,N_5215);
nor U5645 (N_5645,N_4538,N_4756);
or U5646 (N_5646,N_4627,N_4507);
nor U5647 (N_5647,N_4846,N_4569);
nor U5648 (N_5648,N_5007,N_5151);
or U5649 (N_5649,N_5042,N_4745);
nor U5650 (N_5650,N_4512,N_5199);
or U5651 (N_5651,N_4750,N_4591);
or U5652 (N_5652,N_4933,N_5144);
nor U5653 (N_5653,N_5140,N_4561);
or U5654 (N_5654,N_4626,N_4855);
or U5655 (N_5655,N_4811,N_4748);
nand U5656 (N_5656,N_4724,N_4682);
nand U5657 (N_5657,N_5145,N_5023);
nor U5658 (N_5658,N_5159,N_4711);
nor U5659 (N_5659,N_5185,N_4712);
and U5660 (N_5660,N_4942,N_5129);
and U5661 (N_5661,N_4784,N_4650);
and U5662 (N_5662,N_4826,N_4873);
and U5663 (N_5663,N_4506,N_4910);
and U5664 (N_5664,N_4866,N_4728);
nor U5665 (N_5665,N_4693,N_4652);
and U5666 (N_5666,N_4689,N_5038);
nor U5667 (N_5667,N_4831,N_4826);
nor U5668 (N_5668,N_4950,N_5057);
nor U5669 (N_5669,N_4577,N_4676);
and U5670 (N_5670,N_5150,N_4912);
nor U5671 (N_5671,N_5032,N_4668);
or U5672 (N_5672,N_4833,N_5207);
and U5673 (N_5673,N_5198,N_5223);
nand U5674 (N_5674,N_5112,N_4711);
nand U5675 (N_5675,N_4916,N_5160);
nor U5676 (N_5676,N_5179,N_5135);
nor U5677 (N_5677,N_5155,N_4560);
nor U5678 (N_5678,N_4689,N_4604);
nor U5679 (N_5679,N_5144,N_5215);
nand U5680 (N_5680,N_4540,N_4975);
nand U5681 (N_5681,N_4753,N_5212);
or U5682 (N_5682,N_5117,N_4694);
or U5683 (N_5683,N_4731,N_4637);
and U5684 (N_5684,N_4975,N_4635);
nand U5685 (N_5685,N_5080,N_5004);
and U5686 (N_5686,N_5229,N_4904);
or U5687 (N_5687,N_4873,N_4803);
and U5688 (N_5688,N_4641,N_5122);
nor U5689 (N_5689,N_4868,N_4988);
nor U5690 (N_5690,N_5066,N_4972);
or U5691 (N_5691,N_4946,N_5139);
nor U5692 (N_5692,N_4688,N_5165);
and U5693 (N_5693,N_4901,N_5028);
and U5694 (N_5694,N_4661,N_4505);
nor U5695 (N_5695,N_5118,N_5019);
nand U5696 (N_5696,N_4857,N_5067);
nand U5697 (N_5697,N_4616,N_4629);
and U5698 (N_5698,N_4972,N_4848);
nand U5699 (N_5699,N_5147,N_5106);
xor U5700 (N_5700,N_5005,N_5153);
and U5701 (N_5701,N_4643,N_4796);
and U5702 (N_5702,N_4967,N_4848);
and U5703 (N_5703,N_4560,N_4519);
nor U5704 (N_5704,N_4801,N_4639);
nor U5705 (N_5705,N_5218,N_4546);
nand U5706 (N_5706,N_4672,N_4580);
and U5707 (N_5707,N_5210,N_5014);
or U5708 (N_5708,N_4697,N_5201);
and U5709 (N_5709,N_4634,N_5224);
and U5710 (N_5710,N_4531,N_4535);
xnor U5711 (N_5711,N_5094,N_4651);
and U5712 (N_5712,N_4909,N_4820);
or U5713 (N_5713,N_4618,N_5168);
nor U5714 (N_5714,N_4534,N_4515);
nand U5715 (N_5715,N_5148,N_4995);
nand U5716 (N_5716,N_4657,N_4984);
and U5717 (N_5717,N_4740,N_4618);
or U5718 (N_5718,N_5189,N_4779);
nor U5719 (N_5719,N_4621,N_4957);
xor U5720 (N_5720,N_5090,N_4983);
and U5721 (N_5721,N_5003,N_4527);
nor U5722 (N_5722,N_4956,N_4556);
or U5723 (N_5723,N_5164,N_5013);
nor U5724 (N_5724,N_5104,N_5115);
nand U5725 (N_5725,N_4979,N_4641);
nor U5726 (N_5726,N_4832,N_4924);
xnor U5727 (N_5727,N_4779,N_4635);
and U5728 (N_5728,N_4991,N_4650);
nor U5729 (N_5729,N_4742,N_5180);
nor U5730 (N_5730,N_4835,N_4887);
and U5731 (N_5731,N_5110,N_5205);
and U5732 (N_5732,N_4925,N_4587);
or U5733 (N_5733,N_4854,N_5058);
and U5734 (N_5734,N_4645,N_5204);
nor U5735 (N_5735,N_5155,N_4849);
and U5736 (N_5736,N_5098,N_5216);
nand U5737 (N_5737,N_5141,N_4855);
nand U5738 (N_5738,N_4505,N_4823);
or U5739 (N_5739,N_4838,N_4649);
nand U5740 (N_5740,N_4618,N_4578);
and U5741 (N_5741,N_4589,N_4696);
nor U5742 (N_5742,N_4598,N_4581);
or U5743 (N_5743,N_4811,N_4880);
or U5744 (N_5744,N_4647,N_4801);
nor U5745 (N_5745,N_4847,N_4700);
nand U5746 (N_5746,N_5173,N_4688);
nor U5747 (N_5747,N_5127,N_5017);
nand U5748 (N_5748,N_5199,N_4511);
nand U5749 (N_5749,N_4654,N_4530);
nand U5750 (N_5750,N_4757,N_5080);
nand U5751 (N_5751,N_4778,N_5203);
or U5752 (N_5752,N_4651,N_4827);
and U5753 (N_5753,N_5086,N_4983);
or U5754 (N_5754,N_4611,N_4607);
and U5755 (N_5755,N_4662,N_4737);
nand U5756 (N_5756,N_5095,N_5026);
and U5757 (N_5757,N_4990,N_4873);
or U5758 (N_5758,N_4656,N_5201);
or U5759 (N_5759,N_4980,N_4708);
or U5760 (N_5760,N_4594,N_5159);
nand U5761 (N_5761,N_4653,N_4528);
and U5762 (N_5762,N_4909,N_4604);
or U5763 (N_5763,N_4907,N_4565);
or U5764 (N_5764,N_5164,N_4844);
nand U5765 (N_5765,N_4741,N_5231);
xor U5766 (N_5766,N_4931,N_4721);
nand U5767 (N_5767,N_5032,N_4577);
nor U5768 (N_5768,N_4818,N_4992);
or U5769 (N_5769,N_5075,N_4724);
or U5770 (N_5770,N_4584,N_5197);
nor U5771 (N_5771,N_5020,N_4634);
nor U5772 (N_5772,N_5233,N_4674);
nor U5773 (N_5773,N_5134,N_4867);
and U5774 (N_5774,N_4515,N_5120);
nor U5775 (N_5775,N_4615,N_5031);
nand U5776 (N_5776,N_5008,N_4870);
and U5777 (N_5777,N_4778,N_4827);
and U5778 (N_5778,N_4752,N_5021);
and U5779 (N_5779,N_4828,N_4904);
or U5780 (N_5780,N_4727,N_5091);
and U5781 (N_5781,N_4972,N_4863);
or U5782 (N_5782,N_4879,N_5033);
nor U5783 (N_5783,N_5031,N_4748);
and U5784 (N_5784,N_4671,N_4522);
and U5785 (N_5785,N_4559,N_4584);
nor U5786 (N_5786,N_4597,N_4611);
nand U5787 (N_5787,N_4743,N_4851);
and U5788 (N_5788,N_5172,N_4773);
nand U5789 (N_5789,N_4926,N_5083);
or U5790 (N_5790,N_4512,N_4643);
nand U5791 (N_5791,N_4722,N_4549);
and U5792 (N_5792,N_4886,N_4991);
nand U5793 (N_5793,N_5115,N_4806);
and U5794 (N_5794,N_5092,N_5211);
and U5795 (N_5795,N_4942,N_5182);
and U5796 (N_5796,N_4534,N_4946);
nand U5797 (N_5797,N_5242,N_5132);
or U5798 (N_5798,N_5143,N_4862);
or U5799 (N_5799,N_4836,N_4684);
nor U5800 (N_5800,N_4916,N_4716);
nand U5801 (N_5801,N_5192,N_5118);
or U5802 (N_5802,N_5203,N_4717);
or U5803 (N_5803,N_4946,N_5029);
or U5804 (N_5804,N_4533,N_4730);
and U5805 (N_5805,N_5102,N_5052);
or U5806 (N_5806,N_5105,N_5094);
and U5807 (N_5807,N_4659,N_4881);
nor U5808 (N_5808,N_4828,N_4537);
and U5809 (N_5809,N_4920,N_4895);
and U5810 (N_5810,N_4872,N_4875);
and U5811 (N_5811,N_4528,N_5105);
or U5812 (N_5812,N_4584,N_5037);
nand U5813 (N_5813,N_4833,N_4795);
nand U5814 (N_5814,N_5097,N_5115);
nand U5815 (N_5815,N_4909,N_4874);
nand U5816 (N_5816,N_4685,N_4524);
or U5817 (N_5817,N_5064,N_4569);
nand U5818 (N_5818,N_5002,N_5200);
nand U5819 (N_5819,N_4759,N_4555);
nand U5820 (N_5820,N_4995,N_4924);
or U5821 (N_5821,N_4705,N_4749);
and U5822 (N_5822,N_4594,N_5166);
nor U5823 (N_5823,N_5203,N_4964);
xor U5824 (N_5824,N_4734,N_4639);
xnor U5825 (N_5825,N_4984,N_5125);
and U5826 (N_5826,N_4504,N_4670);
nand U5827 (N_5827,N_5040,N_4682);
and U5828 (N_5828,N_4813,N_4944);
or U5829 (N_5829,N_4941,N_4524);
and U5830 (N_5830,N_5030,N_4976);
nor U5831 (N_5831,N_4981,N_4537);
or U5832 (N_5832,N_4910,N_4753);
nor U5833 (N_5833,N_4659,N_4633);
and U5834 (N_5834,N_4988,N_5067);
or U5835 (N_5835,N_4616,N_4729);
nor U5836 (N_5836,N_4548,N_4704);
nand U5837 (N_5837,N_4823,N_4813);
or U5838 (N_5838,N_5227,N_4519);
xnor U5839 (N_5839,N_4797,N_4790);
and U5840 (N_5840,N_4538,N_5220);
nor U5841 (N_5841,N_5216,N_4744);
nor U5842 (N_5842,N_4853,N_4781);
or U5843 (N_5843,N_4550,N_5035);
and U5844 (N_5844,N_4728,N_4528);
or U5845 (N_5845,N_4830,N_4934);
nand U5846 (N_5846,N_5079,N_4987);
nor U5847 (N_5847,N_4595,N_5096);
nand U5848 (N_5848,N_4976,N_5018);
nor U5849 (N_5849,N_4922,N_5050);
and U5850 (N_5850,N_4972,N_5071);
nand U5851 (N_5851,N_5156,N_4708);
and U5852 (N_5852,N_5177,N_5055);
or U5853 (N_5853,N_4746,N_4822);
or U5854 (N_5854,N_5093,N_4828);
and U5855 (N_5855,N_4754,N_5153);
nand U5856 (N_5856,N_5071,N_4796);
or U5857 (N_5857,N_5091,N_4527);
or U5858 (N_5858,N_4882,N_5079);
nor U5859 (N_5859,N_5011,N_4500);
and U5860 (N_5860,N_5102,N_4530);
nand U5861 (N_5861,N_4523,N_4585);
or U5862 (N_5862,N_4981,N_5225);
and U5863 (N_5863,N_4550,N_4970);
nor U5864 (N_5864,N_4931,N_4534);
nand U5865 (N_5865,N_4724,N_5012);
and U5866 (N_5866,N_4887,N_4703);
nor U5867 (N_5867,N_4608,N_4734);
nor U5868 (N_5868,N_4913,N_5055);
or U5869 (N_5869,N_4616,N_4782);
nand U5870 (N_5870,N_4812,N_4508);
nand U5871 (N_5871,N_5076,N_5235);
or U5872 (N_5872,N_5208,N_4683);
nand U5873 (N_5873,N_4933,N_4880);
nand U5874 (N_5874,N_5132,N_4717);
nor U5875 (N_5875,N_4600,N_4597);
and U5876 (N_5876,N_5188,N_5242);
or U5877 (N_5877,N_4766,N_4993);
nand U5878 (N_5878,N_5089,N_4616);
and U5879 (N_5879,N_4577,N_4907);
or U5880 (N_5880,N_4515,N_5163);
nor U5881 (N_5881,N_4518,N_4508);
nand U5882 (N_5882,N_4911,N_5019);
nor U5883 (N_5883,N_4993,N_4836);
and U5884 (N_5884,N_4866,N_5030);
or U5885 (N_5885,N_5079,N_4738);
nand U5886 (N_5886,N_4833,N_4860);
nor U5887 (N_5887,N_4728,N_4799);
nor U5888 (N_5888,N_4556,N_5217);
xor U5889 (N_5889,N_4513,N_5037);
nand U5890 (N_5890,N_4738,N_5122);
or U5891 (N_5891,N_4775,N_5137);
nand U5892 (N_5892,N_4623,N_4670);
or U5893 (N_5893,N_5166,N_4998);
nor U5894 (N_5894,N_5093,N_4549);
or U5895 (N_5895,N_5176,N_4750);
or U5896 (N_5896,N_4600,N_5127);
nand U5897 (N_5897,N_4539,N_5079);
or U5898 (N_5898,N_5234,N_4676);
nor U5899 (N_5899,N_4628,N_4879);
and U5900 (N_5900,N_4609,N_5032);
and U5901 (N_5901,N_5064,N_5178);
or U5902 (N_5902,N_5086,N_5080);
nand U5903 (N_5903,N_5159,N_4891);
nand U5904 (N_5904,N_4921,N_4855);
nand U5905 (N_5905,N_4910,N_5198);
or U5906 (N_5906,N_4620,N_4849);
xnor U5907 (N_5907,N_5065,N_4811);
nand U5908 (N_5908,N_4513,N_5151);
nor U5909 (N_5909,N_4872,N_5073);
or U5910 (N_5910,N_4990,N_4634);
and U5911 (N_5911,N_4636,N_5234);
nor U5912 (N_5912,N_4797,N_5067);
and U5913 (N_5913,N_4635,N_5103);
or U5914 (N_5914,N_4882,N_4978);
nand U5915 (N_5915,N_5036,N_5152);
and U5916 (N_5916,N_4671,N_4736);
nand U5917 (N_5917,N_4713,N_4749);
and U5918 (N_5918,N_4801,N_4815);
nor U5919 (N_5919,N_4857,N_5142);
or U5920 (N_5920,N_4686,N_5220);
nand U5921 (N_5921,N_4564,N_4599);
or U5922 (N_5922,N_5042,N_4587);
xor U5923 (N_5923,N_5062,N_4851);
and U5924 (N_5924,N_5031,N_4654);
nor U5925 (N_5925,N_4655,N_5207);
nor U5926 (N_5926,N_4504,N_4754);
nor U5927 (N_5927,N_4858,N_4647);
and U5928 (N_5928,N_4502,N_5209);
or U5929 (N_5929,N_4970,N_4580);
nor U5930 (N_5930,N_5133,N_4566);
nand U5931 (N_5931,N_4805,N_4553);
nor U5932 (N_5932,N_4585,N_4518);
or U5933 (N_5933,N_4928,N_4997);
nor U5934 (N_5934,N_4553,N_4674);
xnor U5935 (N_5935,N_4944,N_5145);
and U5936 (N_5936,N_4986,N_4806);
and U5937 (N_5937,N_4684,N_5145);
nor U5938 (N_5938,N_4638,N_5118);
nor U5939 (N_5939,N_5193,N_4507);
or U5940 (N_5940,N_4799,N_4698);
nand U5941 (N_5941,N_4934,N_4583);
or U5942 (N_5942,N_5099,N_4586);
nor U5943 (N_5943,N_5022,N_4589);
or U5944 (N_5944,N_4598,N_5089);
or U5945 (N_5945,N_5058,N_4695);
or U5946 (N_5946,N_5047,N_4798);
nor U5947 (N_5947,N_4753,N_4811);
nor U5948 (N_5948,N_4677,N_4573);
nor U5949 (N_5949,N_5103,N_5086);
nand U5950 (N_5950,N_4790,N_4739);
nor U5951 (N_5951,N_4509,N_4978);
nor U5952 (N_5952,N_4518,N_4912);
nor U5953 (N_5953,N_4802,N_4928);
or U5954 (N_5954,N_5045,N_4767);
or U5955 (N_5955,N_4524,N_4651);
and U5956 (N_5956,N_4890,N_4731);
and U5957 (N_5957,N_4826,N_5039);
nor U5958 (N_5958,N_5187,N_5012);
nor U5959 (N_5959,N_4796,N_4855);
or U5960 (N_5960,N_4733,N_4643);
nor U5961 (N_5961,N_5178,N_4584);
and U5962 (N_5962,N_4944,N_4603);
nor U5963 (N_5963,N_4887,N_4708);
nand U5964 (N_5964,N_4872,N_4771);
nand U5965 (N_5965,N_4887,N_4634);
and U5966 (N_5966,N_4671,N_5167);
or U5967 (N_5967,N_4782,N_4506);
or U5968 (N_5968,N_4846,N_4591);
and U5969 (N_5969,N_4966,N_5099);
nand U5970 (N_5970,N_5190,N_5014);
nor U5971 (N_5971,N_4986,N_5037);
nor U5972 (N_5972,N_4795,N_5057);
or U5973 (N_5973,N_5113,N_4608);
nor U5974 (N_5974,N_4855,N_5068);
or U5975 (N_5975,N_4782,N_4621);
nand U5976 (N_5976,N_4803,N_4549);
or U5977 (N_5977,N_5247,N_4688);
and U5978 (N_5978,N_4952,N_4935);
nor U5979 (N_5979,N_5122,N_4640);
nor U5980 (N_5980,N_5020,N_4712);
or U5981 (N_5981,N_5163,N_5034);
nand U5982 (N_5982,N_5016,N_4702);
nor U5983 (N_5983,N_4609,N_4590);
and U5984 (N_5984,N_4843,N_4815);
or U5985 (N_5985,N_4562,N_4902);
nand U5986 (N_5986,N_4553,N_4736);
and U5987 (N_5987,N_5103,N_4733);
nor U5988 (N_5988,N_4741,N_4809);
nor U5989 (N_5989,N_5156,N_5194);
and U5990 (N_5990,N_4749,N_4899);
nand U5991 (N_5991,N_4929,N_5212);
nand U5992 (N_5992,N_4538,N_4557);
nor U5993 (N_5993,N_5195,N_5108);
or U5994 (N_5994,N_4722,N_4876);
and U5995 (N_5995,N_5087,N_4640);
or U5996 (N_5996,N_5074,N_4565);
nor U5997 (N_5997,N_4612,N_4545);
nand U5998 (N_5998,N_5222,N_5139);
nor U5999 (N_5999,N_4649,N_5077);
and U6000 (N_6000,N_5807,N_5912);
or U6001 (N_6001,N_5888,N_5838);
or U6002 (N_6002,N_5868,N_5435);
or U6003 (N_6003,N_5731,N_5593);
nor U6004 (N_6004,N_5942,N_5257);
or U6005 (N_6005,N_5867,N_5330);
xnor U6006 (N_6006,N_5957,N_5745);
or U6007 (N_6007,N_5672,N_5417);
nor U6008 (N_6008,N_5414,N_5560);
nor U6009 (N_6009,N_5752,N_5946);
or U6010 (N_6010,N_5970,N_5284);
and U6011 (N_6011,N_5810,N_5921);
nor U6012 (N_6012,N_5539,N_5675);
and U6013 (N_6013,N_5448,N_5334);
and U6014 (N_6014,N_5835,N_5483);
and U6015 (N_6015,N_5359,N_5447);
nor U6016 (N_6016,N_5380,N_5580);
nand U6017 (N_6017,N_5842,N_5777);
nand U6018 (N_6018,N_5616,N_5324);
nor U6019 (N_6019,N_5335,N_5931);
xor U6020 (N_6020,N_5582,N_5882);
and U6021 (N_6021,N_5609,N_5613);
and U6022 (N_6022,N_5900,N_5724);
nor U6023 (N_6023,N_5309,N_5503);
nor U6024 (N_6024,N_5697,N_5293);
or U6025 (N_6025,N_5977,N_5951);
nand U6026 (N_6026,N_5276,N_5678);
nor U6027 (N_6027,N_5420,N_5575);
and U6028 (N_6028,N_5432,N_5328);
or U6029 (N_6029,N_5500,N_5327);
nor U6030 (N_6030,N_5389,N_5578);
or U6031 (N_6031,N_5894,N_5450);
and U6032 (N_6032,N_5656,N_5401);
or U6033 (N_6033,N_5669,N_5258);
or U6034 (N_6034,N_5784,N_5344);
and U6035 (N_6035,N_5331,N_5909);
and U6036 (N_6036,N_5962,N_5918);
nor U6037 (N_6037,N_5445,N_5374);
nand U6038 (N_6038,N_5915,N_5287);
nor U6039 (N_6039,N_5457,N_5819);
nand U6040 (N_6040,N_5851,N_5727);
and U6041 (N_6041,N_5855,N_5289);
nand U6042 (N_6042,N_5310,N_5622);
nand U6043 (N_6043,N_5419,N_5744);
and U6044 (N_6044,N_5674,N_5824);
and U6045 (N_6045,N_5710,N_5252);
and U6046 (N_6046,N_5464,N_5550);
nand U6047 (N_6047,N_5403,N_5852);
nand U6048 (N_6048,N_5364,N_5486);
or U6049 (N_6049,N_5812,N_5920);
nand U6050 (N_6050,N_5617,N_5573);
nor U6051 (N_6051,N_5633,N_5863);
or U6052 (N_6052,N_5989,N_5716);
nand U6053 (N_6053,N_5369,N_5570);
or U6054 (N_6054,N_5387,N_5526);
and U6055 (N_6055,N_5636,N_5995);
or U6056 (N_6056,N_5907,N_5877);
or U6057 (N_6057,N_5911,N_5879);
or U6058 (N_6058,N_5964,N_5528);
and U6059 (N_6059,N_5822,N_5925);
nand U6060 (N_6060,N_5686,N_5471);
and U6061 (N_6061,N_5607,N_5568);
or U6062 (N_6062,N_5265,N_5983);
and U6063 (N_6063,N_5999,N_5634);
xor U6064 (N_6064,N_5549,N_5308);
nand U6065 (N_6065,N_5288,N_5396);
or U6066 (N_6066,N_5699,N_5996);
nor U6067 (N_6067,N_5735,N_5924);
nand U6068 (N_6068,N_5532,N_5520);
and U6069 (N_6069,N_5495,N_5864);
or U6070 (N_6070,N_5994,N_5552);
nand U6071 (N_6071,N_5981,N_5950);
nor U6072 (N_6072,N_5277,N_5415);
or U6073 (N_6073,N_5423,N_5839);
or U6074 (N_6074,N_5299,N_5829);
nor U6075 (N_6075,N_5397,N_5787);
nor U6076 (N_6076,N_5885,N_5569);
or U6077 (N_6077,N_5251,N_5908);
or U6078 (N_6078,N_5466,N_5395);
and U6079 (N_6079,N_5732,N_5714);
and U6080 (N_6080,N_5998,N_5778);
and U6081 (N_6081,N_5755,N_5934);
nor U6082 (N_6082,N_5943,N_5834);
nor U6083 (N_6083,N_5960,N_5282);
nor U6084 (N_6084,N_5562,N_5640);
nand U6085 (N_6085,N_5291,N_5456);
and U6086 (N_6086,N_5747,N_5583);
nor U6087 (N_6087,N_5704,N_5592);
or U6088 (N_6088,N_5788,N_5507);
or U6089 (N_6089,N_5262,N_5345);
nand U6090 (N_6090,N_5626,N_5661);
and U6091 (N_6091,N_5698,N_5837);
and U6092 (N_6092,N_5862,N_5679);
and U6093 (N_6093,N_5692,N_5270);
or U6094 (N_6094,N_5875,N_5805);
and U6095 (N_6095,N_5988,N_5431);
nor U6096 (N_6096,N_5889,N_5843);
or U6097 (N_6097,N_5748,N_5430);
nor U6098 (N_6098,N_5774,N_5587);
nor U6099 (N_6099,N_5358,N_5904);
nand U6100 (N_6100,N_5687,N_5256);
and U6101 (N_6101,N_5976,N_5429);
or U6102 (N_6102,N_5482,N_5725);
or U6103 (N_6103,N_5991,N_5689);
and U6104 (N_6104,N_5406,N_5901);
nand U6105 (N_6105,N_5368,N_5947);
nand U6106 (N_6106,N_5659,N_5576);
or U6107 (N_6107,N_5497,N_5623);
and U6108 (N_6108,N_5969,N_5340);
or U6109 (N_6109,N_5315,N_5638);
and U6110 (N_6110,N_5425,N_5489);
and U6111 (N_6111,N_5349,N_5555);
and U6112 (N_6112,N_5402,N_5565);
and U6113 (N_6113,N_5399,N_5467);
nor U6114 (N_6114,N_5458,N_5690);
or U6115 (N_6115,N_5440,N_5726);
nand U6116 (N_6116,N_5913,N_5491);
nand U6117 (N_6117,N_5876,N_5292);
or U6118 (N_6118,N_5860,N_5512);
nand U6119 (N_6119,N_5770,N_5800);
nor U6120 (N_6120,N_5502,N_5438);
nor U6121 (N_6121,N_5342,N_5294);
and U6122 (N_6122,N_5619,N_5871);
nor U6123 (N_6123,N_5346,N_5356);
nor U6124 (N_6124,N_5274,N_5741);
nand U6125 (N_6125,N_5514,N_5412);
or U6126 (N_6126,N_5295,N_5769);
or U6127 (N_6127,N_5785,N_5814);
or U6128 (N_6128,N_5685,N_5465);
or U6129 (N_6129,N_5479,N_5338);
nand U6130 (N_6130,N_5606,N_5910);
and U6131 (N_6131,N_5544,N_5645);
nor U6132 (N_6132,N_5985,N_5708);
and U6133 (N_6133,N_5314,N_5574);
nand U6134 (N_6134,N_5798,N_5662);
or U6135 (N_6135,N_5605,N_5844);
and U6136 (N_6136,N_5641,N_5442);
nor U6137 (N_6137,N_5736,N_5452);
nand U6138 (N_6138,N_5892,N_5618);
xnor U6139 (N_6139,N_5786,N_5967);
nand U6140 (N_6140,N_5341,N_5980);
nand U6141 (N_6141,N_5475,N_5493);
and U6142 (N_6142,N_5766,N_5696);
or U6143 (N_6143,N_5504,N_5566);
xnor U6144 (N_6144,N_5557,N_5279);
nand U6145 (N_6145,N_5906,N_5540);
or U6146 (N_6146,N_5953,N_5802);
nor U6147 (N_6147,N_5955,N_5945);
nor U6148 (N_6148,N_5597,N_5360);
nor U6149 (N_6149,N_5776,N_5488);
nand U6150 (N_6150,N_5460,N_5316);
nor U6151 (N_6151,N_5472,N_5434);
nand U6152 (N_6152,N_5377,N_5836);
nand U6153 (N_6153,N_5905,N_5300);
nor U6154 (N_6154,N_5273,N_5919);
and U6155 (N_6155,N_5336,N_5581);
or U6156 (N_6156,N_5719,N_5343);
or U6157 (N_6157,N_5891,N_5433);
nor U6158 (N_6158,N_5803,N_5840);
or U6159 (N_6159,N_5703,N_5268);
and U6160 (N_6160,N_5984,N_5937);
nor U6161 (N_6161,N_5280,N_5372);
and U6162 (N_6162,N_5612,N_5519);
nand U6163 (N_6163,N_5437,N_5305);
or U6164 (N_6164,N_5796,N_5477);
nand U6165 (N_6165,N_5954,N_5362);
and U6166 (N_6166,N_5644,N_5753);
or U6167 (N_6167,N_5734,N_5987);
nor U6168 (N_6168,N_5376,N_5302);
nor U6169 (N_6169,N_5792,N_5333);
xor U6170 (N_6170,N_5663,N_5761);
and U6171 (N_6171,N_5728,N_5285);
or U6172 (N_6172,N_5743,N_5700);
and U6173 (N_6173,N_5563,N_5702);
nand U6174 (N_6174,N_5722,N_5642);
or U6175 (N_6175,N_5628,N_5453);
or U6176 (N_6176,N_5264,N_5579);
or U6177 (N_6177,N_5311,N_5712);
nor U6178 (N_6178,N_5478,N_5409);
and U6179 (N_6179,N_5325,N_5339);
or U6180 (N_6180,N_5610,N_5694);
nand U6181 (N_6181,N_5537,N_5643);
xnor U6182 (N_6182,N_5978,N_5831);
nand U6183 (N_6183,N_5968,N_5365);
and U6184 (N_6184,N_5366,N_5533);
nand U6185 (N_6185,N_5923,N_5706);
and U6186 (N_6186,N_5313,N_5329);
nor U6187 (N_6187,N_5883,N_5808);
nand U6188 (N_6188,N_5804,N_5564);
and U6189 (N_6189,N_5992,N_5518);
or U6190 (N_6190,N_5385,N_5378);
and U6191 (N_6191,N_5383,N_5832);
xor U6192 (N_6192,N_5966,N_5271);
nor U6193 (N_6193,N_5269,N_5446);
and U6194 (N_6194,N_5427,N_5681);
nor U6195 (N_6195,N_5585,N_5426);
nand U6196 (N_6196,N_5870,N_5506);
or U6197 (N_6197,N_5768,N_5469);
nor U6198 (N_6198,N_5749,N_5684);
or U6199 (N_6199,N_5750,N_5283);
or U6200 (N_6200,N_5757,N_5758);
nand U6201 (N_6201,N_5547,N_5599);
nand U6202 (N_6202,N_5650,N_5683);
and U6203 (N_6203,N_5933,N_5290);
or U6204 (N_6204,N_5858,N_5281);
or U6205 (N_6205,N_5668,N_5973);
xnor U6206 (N_6206,N_5790,N_5789);
nor U6207 (N_6207,N_5411,N_5746);
xor U6208 (N_6208,N_5772,N_5737);
and U6209 (N_6209,N_5721,N_5454);
nand U6210 (N_6210,N_5306,N_5880);
and U6211 (N_6211,N_5637,N_5523);
xor U6212 (N_6212,N_5588,N_5941);
nand U6213 (N_6213,N_5986,N_5887);
and U6214 (N_6214,N_5494,N_5261);
nand U6215 (N_6215,N_5938,N_5490);
nand U6216 (N_6216,N_5404,N_5455);
or U6217 (N_6217,N_5484,N_5348);
nand U6218 (N_6218,N_5538,N_5598);
nand U6219 (N_6219,N_5370,N_5701);
nor U6220 (N_6220,N_5765,N_5474);
and U6221 (N_6221,N_5559,N_5558);
or U6222 (N_6222,N_5793,N_5630);
or U6223 (N_6223,N_5958,N_5361);
and U6224 (N_6224,N_5801,N_5853);
or U6225 (N_6225,N_5711,N_5422);
nor U6226 (N_6226,N_5903,N_5817);
nand U6227 (N_6227,N_5823,N_5825);
nor U6228 (N_6228,N_5647,N_5254);
and U6229 (N_6229,N_5929,N_5255);
and U6230 (N_6230,N_5393,N_5548);
nand U6231 (N_6231,N_5917,N_5354);
or U6232 (N_6232,N_5556,N_5449);
nand U6233 (N_6233,N_5657,N_5517);
or U6234 (N_6234,N_5818,N_5317);
and U6235 (N_6235,N_5615,N_5390);
or U6236 (N_6236,N_5625,N_5729);
and U6237 (N_6237,N_5384,N_5531);
xor U6238 (N_6238,N_5353,N_5854);
or U6239 (N_6239,N_5667,N_5516);
and U6240 (N_6240,N_5884,N_5705);
nor U6241 (N_6241,N_5660,N_5527);
nor U6242 (N_6242,N_5845,N_5545);
and U6243 (N_6243,N_5461,N_5443);
nor U6244 (N_6244,N_5791,N_5990);
nand U6245 (N_6245,N_5982,N_5253);
and U6246 (N_6246,N_5682,N_5873);
nor U6247 (N_6247,N_5751,N_5898);
and U6248 (N_6248,N_5730,N_5820);
nor U6249 (N_6249,N_5602,N_5723);
and U6250 (N_6250,N_5809,N_5351);
and U6251 (N_6251,N_5930,N_5653);
and U6252 (N_6252,N_5782,N_5421);
or U6253 (N_6253,N_5505,N_5286);
nor U6254 (N_6254,N_5577,N_5902);
nor U6255 (N_6255,N_5866,N_5848);
nand U6256 (N_6256,N_5767,N_5522);
and U6257 (N_6257,N_5974,N_5468);
nand U6258 (N_6258,N_5551,N_5715);
or U6259 (N_6259,N_5304,N_5811);
or U6260 (N_6260,N_5997,N_5826);
nand U6261 (N_6261,N_5590,N_5267);
or U6262 (N_6262,N_5754,N_5611);
xnor U6263 (N_6263,N_5677,N_5398);
nor U6264 (N_6264,N_5707,N_5546);
nor U6265 (N_6265,N_5509,N_5895);
nand U6266 (N_6266,N_5652,N_5524);
nor U6267 (N_6267,N_5830,N_5441);
nand U6268 (N_6268,N_5897,N_5312);
or U6269 (N_6269,N_5260,N_5932);
or U6270 (N_6270,N_5266,N_5779);
nor U6271 (N_6271,N_5865,N_5673);
nor U6272 (N_6272,N_5428,N_5525);
nor U6273 (N_6273,N_5529,N_5319);
and U6274 (N_6274,N_5410,N_5595);
nand U6275 (N_6275,N_5498,N_5718);
or U6276 (N_6276,N_5407,N_5499);
or U6277 (N_6277,N_5496,N_5381);
nor U6278 (N_6278,N_5713,N_5740);
or U6279 (N_6279,N_5648,N_5815);
nor U6280 (N_6280,N_5326,N_5795);
nor U6281 (N_6281,N_5553,N_5695);
nand U6282 (N_6282,N_5927,N_5600);
and U6283 (N_6283,N_5914,N_5688);
nand U6284 (N_6284,N_5841,N_5806);
nand U6285 (N_6285,N_5510,N_5307);
nor U6286 (N_6286,N_5965,N_5391);
or U6287 (N_6287,N_5275,N_5534);
nor U6288 (N_6288,N_5298,N_5416);
xor U6289 (N_6289,N_5926,N_5896);
nor U6290 (N_6290,N_5386,N_5463);
nand U6291 (N_6291,N_5589,N_5691);
and U6292 (N_6292,N_5367,N_5278);
or U6293 (N_6293,N_5530,N_5709);
nor U6294 (N_6294,N_5554,N_5763);
or U6295 (N_6295,N_5813,N_5759);
nand U6296 (N_6296,N_5665,N_5733);
and U6297 (N_6297,N_5318,N_5601);
or U6298 (N_6298,N_5881,N_5572);
nor U6299 (N_6299,N_5424,N_5408);
and U6300 (N_6300,N_5827,N_5833);
nor U6301 (N_6301,N_5620,N_5451);
nand U6302 (N_6302,N_5671,N_5541);
or U6303 (N_6303,N_5487,N_5939);
nor U6304 (N_6304,N_5462,N_5869);
or U6305 (N_6305,N_5664,N_5571);
nor U6306 (N_6306,N_5321,N_5756);
or U6307 (N_6307,N_5821,N_5961);
and U6308 (N_6308,N_5670,N_5739);
nor U6309 (N_6309,N_5259,N_5676);
nand U6310 (N_6310,N_5392,N_5413);
and U6311 (N_6311,N_5631,N_5492);
nand U6312 (N_6312,N_5485,N_5418);
nand U6313 (N_6313,N_5476,N_5388);
nand U6314 (N_6314,N_5543,N_5720);
nor U6315 (N_6315,N_5979,N_5762);
nor U6316 (N_6316,N_5297,N_5649);
nand U6317 (N_6317,N_5470,N_5473);
nand U6318 (N_6318,N_5874,N_5935);
nor U6319 (N_6319,N_5263,N_5373);
nor U6320 (N_6320,N_5603,N_5760);
nand U6321 (N_6321,N_5511,N_5515);
and U6322 (N_6322,N_5629,N_5347);
nand U6323 (N_6323,N_5379,N_5856);
nor U6324 (N_6324,N_5849,N_5890);
nand U6325 (N_6325,N_5742,N_5561);
nor U6326 (N_6326,N_5738,N_5439);
and U6327 (N_6327,N_5480,N_5847);
and U6328 (N_6328,N_5627,N_5651);
or U6329 (N_6329,N_5371,N_5899);
or U6330 (N_6330,N_5680,N_5624);
or U6331 (N_6331,N_5355,N_5944);
or U6332 (N_6332,N_5591,N_5352);
nor U6333 (N_6333,N_5952,N_5350);
and U6334 (N_6334,N_5357,N_5646);
nor U6335 (N_6335,N_5521,N_5322);
nand U6336 (N_6336,N_5621,N_5382);
or U6337 (N_6337,N_5303,N_5272);
or U6338 (N_6338,N_5872,N_5963);
xor U6339 (N_6339,N_5586,N_5916);
or U6340 (N_6340,N_5584,N_5535);
and U6341 (N_6341,N_5949,N_5693);
and U6342 (N_6342,N_5956,N_5596);
nand U6343 (N_6343,N_5857,N_5501);
or U6344 (N_6344,N_5928,N_5594);
nand U6345 (N_6345,N_5773,N_5614);
nor U6346 (N_6346,N_5717,N_5783);
nand U6347 (N_6347,N_5323,N_5508);
nor U6348 (N_6348,N_5799,N_5828);
nand U6349 (N_6349,N_5797,N_5886);
and U6350 (N_6350,N_5405,N_5363);
nor U6351 (N_6351,N_5301,N_5250);
nand U6352 (N_6352,N_5893,N_5536);
and U6353 (N_6353,N_5608,N_5513);
and U6354 (N_6354,N_5993,N_5972);
or U6355 (N_6355,N_5332,N_5604);
nor U6356 (N_6356,N_5337,N_5859);
or U6357 (N_6357,N_5444,N_5436);
and U6358 (N_6358,N_5775,N_5794);
nand U6359 (N_6359,N_5816,N_5959);
nand U6360 (N_6360,N_5781,N_5481);
nand U6361 (N_6361,N_5971,N_5400);
and U6362 (N_6362,N_5394,N_5654);
nor U6363 (N_6363,N_5846,N_5940);
nor U6364 (N_6364,N_5666,N_5780);
nand U6365 (N_6365,N_5861,N_5655);
and U6366 (N_6366,N_5459,N_5936);
or U6367 (N_6367,N_5922,N_5542);
nor U6368 (N_6368,N_5567,N_5658);
and U6369 (N_6369,N_5975,N_5632);
and U6370 (N_6370,N_5771,N_5296);
or U6371 (N_6371,N_5375,N_5635);
and U6372 (N_6372,N_5639,N_5878);
nor U6373 (N_6373,N_5948,N_5320);
nand U6374 (N_6374,N_5764,N_5850);
and U6375 (N_6375,N_5963,N_5810);
nor U6376 (N_6376,N_5751,N_5445);
nor U6377 (N_6377,N_5812,N_5599);
xor U6378 (N_6378,N_5637,N_5380);
and U6379 (N_6379,N_5272,N_5453);
nor U6380 (N_6380,N_5808,N_5858);
nor U6381 (N_6381,N_5696,N_5611);
nand U6382 (N_6382,N_5595,N_5838);
xnor U6383 (N_6383,N_5902,N_5728);
nor U6384 (N_6384,N_5889,N_5982);
nor U6385 (N_6385,N_5380,N_5482);
and U6386 (N_6386,N_5882,N_5414);
nor U6387 (N_6387,N_5809,N_5726);
nand U6388 (N_6388,N_5344,N_5297);
and U6389 (N_6389,N_5653,N_5909);
or U6390 (N_6390,N_5488,N_5578);
nor U6391 (N_6391,N_5854,N_5922);
and U6392 (N_6392,N_5669,N_5597);
or U6393 (N_6393,N_5683,N_5267);
nor U6394 (N_6394,N_5873,N_5728);
or U6395 (N_6395,N_5533,N_5545);
nor U6396 (N_6396,N_5870,N_5343);
nand U6397 (N_6397,N_5444,N_5661);
nand U6398 (N_6398,N_5941,N_5333);
or U6399 (N_6399,N_5552,N_5371);
nor U6400 (N_6400,N_5361,N_5787);
nand U6401 (N_6401,N_5504,N_5909);
nand U6402 (N_6402,N_5837,N_5490);
or U6403 (N_6403,N_5740,N_5599);
nand U6404 (N_6404,N_5376,N_5700);
nor U6405 (N_6405,N_5837,N_5354);
or U6406 (N_6406,N_5255,N_5922);
nand U6407 (N_6407,N_5661,N_5680);
and U6408 (N_6408,N_5741,N_5563);
nand U6409 (N_6409,N_5337,N_5685);
or U6410 (N_6410,N_5779,N_5259);
nand U6411 (N_6411,N_5480,N_5473);
nor U6412 (N_6412,N_5321,N_5806);
nor U6413 (N_6413,N_5784,N_5450);
and U6414 (N_6414,N_5892,N_5634);
or U6415 (N_6415,N_5275,N_5586);
or U6416 (N_6416,N_5820,N_5883);
nand U6417 (N_6417,N_5280,N_5858);
nor U6418 (N_6418,N_5690,N_5891);
or U6419 (N_6419,N_5401,N_5469);
nor U6420 (N_6420,N_5356,N_5362);
and U6421 (N_6421,N_5860,N_5287);
or U6422 (N_6422,N_5877,N_5601);
nor U6423 (N_6423,N_5804,N_5701);
and U6424 (N_6424,N_5768,N_5905);
or U6425 (N_6425,N_5516,N_5813);
and U6426 (N_6426,N_5515,N_5757);
or U6427 (N_6427,N_5823,N_5583);
and U6428 (N_6428,N_5473,N_5491);
and U6429 (N_6429,N_5460,N_5949);
or U6430 (N_6430,N_5631,N_5481);
xnor U6431 (N_6431,N_5666,N_5352);
nor U6432 (N_6432,N_5937,N_5903);
and U6433 (N_6433,N_5312,N_5539);
or U6434 (N_6434,N_5883,N_5669);
or U6435 (N_6435,N_5862,N_5520);
nand U6436 (N_6436,N_5810,N_5385);
nand U6437 (N_6437,N_5925,N_5509);
nor U6438 (N_6438,N_5822,N_5940);
and U6439 (N_6439,N_5825,N_5434);
and U6440 (N_6440,N_5966,N_5438);
nand U6441 (N_6441,N_5907,N_5717);
and U6442 (N_6442,N_5325,N_5546);
or U6443 (N_6443,N_5785,N_5676);
nor U6444 (N_6444,N_5868,N_5490);
nand U6445 (N_6445,N_5458,N_5790);
and U6446 (N_6446,N_5662,N_5547);
or U6447 (N_6447,N_5979,N_5854);
nand U6448 (N_6448,N_5812,N_5660);
or U6449 (N_6449,N_5282,N_5263);
nand U6450 (N_6450,N_5923,N_5398);
and U6451 (N_6451,N_5829,N_5663);
xor U6452 (N_6452,N_5901,N_5993);
nor U6453 (N_6453,N_5338,N_5545);
and U6454 (N_6454,N_5288,N_5259);
and U6455 (N_6455,N_5591,N_5280);
and U6456 (N_6456,N_5894,N_5489);
nor U6457 (N_6457,N_5288,N_5535);
and U6458 (N_6458,N_5808,N_5485);
and U6459 (N_6459,N_5411,N_5529);
nor U6460 (N_6460,N_5883,N_5578);
nor U6461 (N_6461,N_5303,N_5302);
or U6462 (N_6462,N_5953,N_5667);
nor U6463 (N_6463,N_5400,N_5604);
or U6464 (N_6464,N_5755,N_5853);
nand U6465 (N_6465,N_5360,N_5767);
nor U6466 (N_6466,N_5419,N_5612);
nor U6467 (N_6467,N_5750,N_5809);
and U6468 (N_6468,N_5802,N_5568);
or U6469 (N_6469,N_5971,N_5545);
nor U6470 (N_6470,N_5468,N_5582);
or U6471 (N_6471,N_5277,N_5615);
nand U6472 (N_6472,N_5897,N_5431);
nor U6473 (N_6473,N_5847,N_5491);
or U6474 (N_6474,N_5372,N_5497);
or U6475 (N_6475,N_5559,N_5833);
nor U6476 (N_6476,N_5866,N_5760);
or U6477 (N_6477,N_5528,N_5400);
nor U6478 (N_6478,N_5965,N_5657);
nand U6479 (N_6479,N_5364,N_5554);
and U6480 (N_6480,N_5756,N_5802);
and U6481 (N_6481,N_5471,N_5345);
nor U6482 (N_6482,N_5384,N_5936);
and U6483 (N_6483,N_5430,N_5373);
or U6484 (N_6484,N_5358,N_5907);
and U6485 (N_6485,N_5740,N_5730);
nor U6486 (N_6486,N_5313,N_5510);
nor U6487 (N_6487,N_5468,N_5341);
and U6488 (N_6488,N_5294,N_5648);
nand U6489 (N_6489,N_5372,N_5882);
nor U6490 (N_6490,N_5261,N_5784);
and U6491 (N_6491,N_5977,N_5749);
or U6492 (N_6492,N_5684,N_5739);
and U6493 (N_6493,N_5833,N_5752);
nand U6494 (N_6494,N_5973,N_5747);
nand U6495 (N_6495,N_5639,N_5251);
nor U6496 (N_6496,N_5860,N_5703);
or U6497 (N_6497,N_5563,N_5899);
nor U6498 (N_6498,N_5462,N_5753);
and U6499 (N_6499,N_5316,N_5855);
xor U6500 (N_6500,N_5536,N_5433);
xor U6501 (N_6501,N_5597,N_5774);
nor U6502 (N_6502,N_5725,N_5952);
nand U6503 (N_6503,N_5821,N_5928);
nand U6504 (N_6504,N_5679,N_5476);
nand U6505 (N_6505,N_5546,N_5981);
nand U6506 (N_6506,N_5377,N_5333);
or U6507 (N_6507,N_5564,N_5837);
xor U6508 (N_6508,N_5553,N_5668);
nor U6509 (N_6509,N_5909,N_5328);
xor U6510 (N_6510,N_5919,N_5423);
nand U6511 (N_6511,N_5736,N_5361);
nand U6512 (N_6512,N_5282,N_5387);
nor U6513 (N_6513,N_5912,N_5741);
and U6514 (N_6514,N_5930,N_5497);
or U6515 (N_6515,N_5684,N_5573);
and U6516 (N_6516,N_5569,N_5598);
nand U6517 (N_6517,N_5411,N_5630);
nand U6518 (N_6518,N_5789,N_5335);
nand U6519 (N_6519,N_5654,N_5570);
and U6520 (N_6520,N_5753,N_5376);
and U6521 (N_6521,N_5830,N_5292);
and U6522 (N_6522,N_5888,N_5755);
nor U6523 (N_6523,N_5857,N_5890);
and U6524 (N_6524,N_5837,N_5364);
nor U6525 (N_6525,N_5426,N_5937);
nand U6526 (N_6526,N_5871,N_5491);
nand U6527 (N_6527,N_5531,N_5449);
and U6528 (N_6528,N_5379,N_5777);
nor U6529 (N_6529,N_5296,N_5288);
or U6530 (N_6530,N_5885,N_5478);
and U6531 (N_6531,N_5533,N_5856);
and U6532 (N_6532,N_5502,N_5529);
nand U6533 (N_6533,N_5846,N_5856);
or U6534 (N_6534,N_5443,N_5292);
or U6535 (N_6535,N_5745,N_5542);
nand U6536 (N_6536,N_5446,N_5284);
nor U6537 (N_6537,N_5750,N_5345);
and U6538 (N_6538,N_5747,N_5399);
nor U6539 (N_6539,N_5405,N_5481);
or U6540 (N_6540,N_5425,N_5494);
nor U6541 (N_6541,N_5702,N_5285);
nor U6542 (N_6542,N_5913,N_5498);
or U6543 (N_6543,N_5261,N_5601);
and U6544 (N_6544,N_5719,N_5835);
or U6545 (N_6545,N_5896,N_5423);
or U6546 (N_6546,N_5708,N_5346);
and U6547 (N_6547,N_5774,N_5877);
nand U6548 (N_6548,N_5848,N_5537);
nor U6549 (N_6549,N_5776,N_5947);
or U6550 (N_6550,N_5267,N_5900);
and U6551 (N_6551,N_5562,N_5870);
nand U6552 (N_6552,N_5988,N_5777);
and U6553 (N_6553,N_5298,N_5532);
or U6554 (N_6554,N_5357,N_5490);
and U6555 (N_6555,N_5992,N_5430);
and U6556 (N_6556,N_5777,N_5946);
nor U6557 (N_6557,N_5984,N_5914);
nand U6558 (N_6558,N_5641,N_5723);
nor U6559 (N_6559,N_5427,N_5692);
and U6560 (N_6560,N_5507,N_5484);
nor U6561 (N_6561,N_5369,N_5355);
nand U6562 (N_6562,N_5718,N_5731);
nand U6563 (N_6563,N_5530,N_5726);
nand U6564 (N_6564,N_5904,N_5948);
nand U6565 (N_6565,N_5544,N_5888);
or U6566 (N_6566,N_5559,N_5668);
or U6567 (N_6567,N_5830,N_5554);
or U6568 (N_6568,N_5824,N_5945);
and U6569 (N_6569,N_5725,N_5611);
nor U6570 (N_6570,N_5306,N_5715);
or U6571 (N_6571,N_5872,N_5727);
nand U6572 (N_6572,N_5534,N_5777);
nor U6573 (N_6573,N_5629,N_5276);
nand U6574 (N_6574,N_5516,N_5606);
or U6575 (N_6575,N_5853,N_5821);
and U6576 (N_6576,N_5560,N_5292);
or U6577 (N_6577,N_5579,N_5559);
nor U6578 (N_6578,N_5777,N_5301);
xnor U6579 (N_6579,N_5966,N_5652);
or U6580 (N_6580,N_5786,N_5383);
nand U6581 (N_6581,N_5561,N_5569);
or U6582 (N_6582,N_5593,N_5295);
nand U6583 (N_6583,N_5801,N_5980);
or U6584 (N_6584,N_5827,N_5317);
or U6585 (N_6585,N_5713,N_5954);
and U6586 (N_6586,N_5899,N_5455);
nand U6587 (N_6587,N_5428,N_5489);
or U6588 (N_6588,N_5358,N_5678);
nand U6589 (N_6589,N_5407,N_5683);
or U6590 (N_6590,N_5774,N_5860);
or U6591 (N_6591,N_5946,N_5698);
or U6592 (N_6592,N_5968,N_5871);
xor U6593 (N_6593,N_5284,N_5393);
or U6594 (N_6594,N_5399,N_5721);
or U6595 (N_6595,N_5799,N_5810);
and U6596 (N_6596,N_5955,N_5345);
or U6597 (N_6597,N_5844,N_5615);
nor U6598 (N_6598,N_5746,N_5817);
or U6599 (N_6599,N_5525,N_5816);
and U6600 (N_6600,N_5368,N_5325);
or U6601 (N_6601,N_5724,N_5881);
or U6602 (N_6602,N_5825,N_5759);
and U6603 (N_6603,N_5972,N_5468);
xnor U6604 (N_6604,N_5317,N_5725);
and U6605 (N_6605,N_5345,N_5304);
and U6606 (N_6606,N_5544,N_5844);
and U6607 (N_6607,N_5777,N_5891);
or U6608 (N_6608,N_5452,N_5565);
or U6609 (N_6609,N_5636,N_5913);
and U6610 (N_6610,N_5665,N_5520);
and U6611 (N_6611,N_5582,N_5465);
nand U6612 (N_6612,N_5691,N_5710);
and U6613 (N_6613,N_5346,N_5459);
nor U6614 (N_6614,N_5842,N_5479);
nor U6615 (N_6615,N_5582,N_5358);
nand U6616 (N_6616,N_5948,N_5424);
nand U6617 (N_6617,N_5277,N_5611);
nand U6618 (N_6618,N_5788,N_5305);
or U6619 (N_6619,N_5483,N_5976);
nor U6620 (N_6620,N_5802,N_5670);
nand U6621 (N_6621,N_5592,N_5948);
or U6622 (N_6622,N_5427,N_5400);
or U6623 (N_6623,N_5894,N_5934);
xor U6624 (N_6624,N_5450,N_5799);
nand U6625 (N_6625,N_5849,N_5258);
xnor U6626 (N_6626,N_5342,N_5322);
and U6627 (N_6627,N_5355,N_5915);
nor U6628 (N_6628,N_5766,N_5577);
or U6629 (N_6629,N_5493,N_5750);
and U6630 (N_6630,N_5967,N_5673);
nor U6631 (N_6631,N_5498,N_5416);
or U6632 (N_6632,N_5846,N_5602);
and U6633 (N_6633,N_5933,N_5379);
and U6634 (N_6634,N_5583,N_5810);
nor U6635 (N_6635,N_5514,N_5963);
nand U6636 (N_6636,N_5599,N_5417);
or U6637 (N_6637,N_5987,N_5849);
nand U6638 (N_6638,N_5751,N_5733);
nor U6639 (N_6639,N_5362,N_5704);
or U6640 (N_6640,N_5744,N_5705);
or U6641 (N_6641,N_5398,N_5942);
nand U6642 (N_6642,N_5627,N_5884);
and U6643 (N_6643,N_5634,N_5642);
nor U6644 (N_6644,N_5743,N_5542);
or U6645 (N_6645,N_5771,N_5376);
nand U6646 (N_6646,N_5549,N_5812);
xor U6647 (N_6647,N_5666,N_5827);
and U6648 (N_6648,N_5655,N_5304);
xor U6649 (N_6649,N_5771,N_5617);
or U6650 (N_6650,N_5568,N_5709);
nor U6651 (N_6651,N_5475,N_5893);
or U6652 (N_6652,N_5739,N_5877);
and U6653 (N_6653,N_5982,N_5361);
nor U6654 (N_6654,N_5775,N_5415);
and U6655 (N_6655,N_5631,N_5675);
nand U6656 (N_6656,N_5755,N_5287);
or U6657 (N_6657,N_5960,N_5424);
or U6658 (N_6658,N_5813,N_5475);
or U6659 (N_6659,N_5485,N_5483);
nand U6660 (N_6660,N_5747,N_5676);
or U6661 (N_6661,N_5480,N_5603);
nor U6662 (N_6662,N_5528,N_5745);
or U6663 (N_6663,N_5717,N_5655);
nor U6664 (N_6664,N_5847,N_5667);
nor U6665 (N_6665,N_5651,N_5811);
or U6666 (N_6666,N_5699,N_5940);
nand U6667 (N_6667,N_5716,N_5813);
nand U6668 (N_6668,N_5584,N_5469);
nor U6669 (N_6669,N_5459,N_5554);
and U6670 (N_6670,N_5683,N_5435);
and U6671 (N_6671,N_5927,N_5696);
nand U6672 (N_6672,N_5383,N_5520);
or U6673 (N_6673,N_5915,N_5866);
or U6674 (N_6674,N_5997,N_5615);
nor U6675 (N_6675,N_5619,N_5900);
xor U6676 (N_6676,N_5722,N_5686);
and U6677 (N_6677,N_5383,N_5572);
and U6678 (N_6678,N_5850,N_5988);
nand U6679 (N_6679,N_5652,N_5826);
nor U6680 (N_6680,N_5261,N_5961);
nor U6681 (N_6681,N_5931,N_5259);
or U6682 (N_6682,N_5480,N_5837);
or U6683 (N_6683,N_5577,N_5555);
and U6684 (N_6684,N_5254,N_5435);
and U6685 (N_6685,N_5376,N_5387);
nor U6686 (N_6686,N_5775,N_5276);
and U6687 (N_6687,N_5799,N_5642);
nor U6688 (N_6688,N_5808,N_5818);
or U6689 (N_6689,N_5593,N_5360);
nand U6690 (N_6690,N_5390,N_5715);
nand U6691 (N_6691,N_5899,N_5268);
or U6692 (N_6692,N_5472,N_5984);
xor U6693 (N_6693,N_5829,N_5447);
or U6694 (N_6694,N_5858,N_5667);
nand U6695 (N_6695,N_5428,N_5554);
nor U6696 (N_6696,N_5626,N_5292);
nor U6697 (N_6697,N_5702,N_5348);
and U6698 (N_6698,N_5686,N_5314);
nand U6699 (N_6699,N_5571,N_5823);
nor U6700 (N_6700,N_5596,N_5570);
and U6701 (N_6701,N_5859,N_5837);
or U6702 (N_6702,N_5994,N_5933);
nand U6703 (N_6703,N_5369,N_5702);
nor U6704 (N_6704,N_5367,N_5287);
xor U6705 (N_6705,N_5738,N_5786);
nand U6706 (N_6706,N_5435,N_5899);
or U6707 (N_6707,N_5888,N_5795);
nand U6708 (N_6708,N_5720,N_5299);
or U6709 (N_6709,N_5864,N_5852);
nor U6710 (N_6710,N_5743,N_5267);
or U6711 (N_6711,N_5631,N_5600);
nor U6712 (N_6712,N_5776,N_5748);
nand U6713 (N_6713,N_5637,N_5853);
nor U6714 (N_6714,N_5810,N_5339);
and U6715 (N_6715,N_5423,N_5520);
nor U6716 (N_6716,N_5864,N_5456);
or U6717 (N_6717,N_5756,N_5960);
and U6718 (N_6718,N_5630,N_5525);
or U6719 (N_6719,N_5964,N_5911);
and U6720 (N_6720,N_5650,N_5492);
and U6721 (N_6721,N_5266,N_5410);
and U6722 (N_6722,N_5876,N_5542);
nor U6723 (N_6723,N_5551,N_5397);
nand U6724 (N_6724,N_5940,N_5371);
or U6725 (N_6725,N_5491,N_5465);
nor U6726 (N_6726,N_5350,N_5405);
nor U6727 (N_6727,N_5462,N_5331);
and U6728 (N_6728,N_5633,N_5700);
and U6729 (N_6729,N_5683,N_5410);
nand U6730 (N_6730,N_5706,N_5352);
nand U6731 (N_6731,N_5987,N_5373);
nand U6732 (N_6732,N_5451,N_5691);
and U6733 (N_6733,N_5963,N_5814);
and U6734 (N_6734,N_5595,N_5946);
nand U6735 (N_6735,N_5509,N_5965);
nand U6736 (N_6736,N_5666,N_5826);
and U6737 (N_6737,N_5267,N_5286);
nand U6738 (N_6738,N_5662,N_5463);
or U6739 (N_6739,N_5782,N_5956);
nor U6740 (N_6740,N_5579,N_5943);
nor U6741 (N_6741,N_5683,N_5569);
xnor U6742 (N_6742,N_5338,N_5603);
or U6743 (N_6743,N_5598,N_5980);
and U6744 (N_6744,N_5952,N_5964);
or U6745 (N_6745,N_5280,N_5575);
nand U6746 (N_6746,N_5342,N_5368);
and U6747 (N_6747,N_5310,N_5737);
nand U6748 (N_6748,N_5720,N_5964);
nand U6749 (N_6749,N_5598,N_5820);
and U6750 (N_6750,N_6010,N_6506);
or U6751 (N_6751,N_6655,N_6077);
nor U6752 (N_6752,N_6423,N_6610);
or U6753 (N_6753,N_6226,N_6576);
nor U6754 (N_6754,N_6570,N_6253);
or U6755 (N_6755,N_6460,N_6478);
or U6756 (N_6756,N_6186,N_6062);
or U6757 (N_6757,N_6304,N_6048);
or U6758 (N_6758,N_6428,N_6211);
or U6759 (N_6759,N_6337,N_6422);
or U6760 (N_6760,N_6325,N_6220);
and U6761 (N_6761,N_6547,N_6736);
nand U6762 (N_6762,N_6013,N_6002);
nor U6763 (N_6763,N_6335,N_6394);
nand U6764 (N_6764,N_6266,N_6030);
nor U6765 (N_6765,N_6638,N_6140);
or U6766 (N_6766,N_6119,N_6381);
or U6767 (N_6767,N_6678,N_6364);
nor U6768 (N_6768,N_6214,N_6050);
and U6769 (N_6769,N_6219,N_6651);
xnor U6770 (N_6770,N_6730,N_6668);
or U6771 (N_6771,N_6566,N_6522);
nor U6772 (N_6772,N_6090,N_6221);
nand U6773 (N_6773,N_6291,N_6306);
nand U6774 (N_6774,N_6380,N_6127);
and U6775 (N_6775,N_6677,N_6145);
nand U6776 (N_6776,N_6182,N_6404);
nand U6777 (N_6777,N_6009,N_6698);
nor U6778 (N_6778,N_6323,N_6473);
nor U6779 (N_6779,N_6063,N_6372);
xor U6780 (N_6780,N_6016,N_6263);
or U6781 (N_6781,N_6113,N_6560);
and U6782 (N_6782,N_6561,N_6539);
xor U6783 (N_6783,N_6684,N_6542);
or U6784 (N_6784,N_6005,N_6284);
nand U6785 (N_6785,N_6187,N_6289);
nand U6786 (N_6786,N_6258,N_6511);
nand U6787 (N_6787,N_6400,N_6331);
or U6788 (N_6788,N_6744,N_6327);
or U6789 (N_6789,N_6254,N_6321);
and U6790 (N_6790,N_6554,N_6636);
and U6791 (N_6791,N_6704,N_6023);
or U6792 (N_6792,N_6061,N_6671);
and U6793 (N_6793,N_6732,N_6098);
or U6794 (N_6794,N_6371,N_6456);
nand U6795 (N_6795,N_6541,N_6477);
and U6796 (N_6796,N_6339,N_6660);
and U6797 (N_6797,N_6000,N_6348);
and U6798 (N_6798,N_6224,N_6682);
or U6799 (N_6799,N_6095,N_6611);
nor U6800 (N_6800,N_6391,N_6599);
and U6801 (N_6801,N_6232,N_6108);
or U6802 (N_6802,N_6410,N_6315);
or U6803 (N_6803,N_6305,N_6267);
xnor U6804 (N_6804,N_6406,N_6279);
nor U6805 (N_6805,N_6157,N_6720);
and U6806 (N_6806,N_6256,N_6713);
or U6807 (N_6807,N_6303,N_6045);
nor U6808 (N_6808,N_6646,N_6012);
or U6809 (N_6809,N_6618,N_6594);
nand U6810 (N_6810,N_6626,N_6625);
nand U6811 (N_6811,N_6234,N_6426);
nor U6812 (N_6812,N_6096,N_6044);
and U6813 (N_6813,N_6616,N_6179);
and U6814 (N_6814,N_6637,N_6197);
nand U6815 (N_6815,N_6240,N_6430);
nand U6816 (N_6816,N_6553,N_6395);
nor U6817 (N_6817,N_6535,N_6326);
nand U6818 (N_6818,N_6270,N_6347);
or U6819 (N_6819,N_6213,N_6021);
xor U6820 (N_6820,N_6297,N_6557);
or U6821 (N_6821,N_6417,N_6414);
and U6822 (N_6822,N_6549,N_6078);
and U6823 (N_6823,N_6527,N_6679);
and U6824 (N_6824,N_6196,N_6368);
nor U6825 (N_6825,N_6249,N_6248);
nor U6826 (N_6826,N_6536,N_6362);
or U6827 (N_6827,N_6559,N_6401);
nor U6828 (N_6828,N_6114,N_6302);
nand U6829 (N_6829,N_6017,N_6738);
nand U6830 (N_6830,N_6568,N_6386);
and U6831 (N_6831,N_6603,N_6105);
nor U6832 (N_6832,N_6457,N_6107);
nor U6833 (N_6833,N_6295,N_6491);
and U6834 (N_6834,N_6130,N_6701);
nand U6835 (N_6835,N_6168,N_6237);
or U6836 (N_6836,N_6470,N_6039);
or U6837 (N_6837,N_6116,N_6055);
and U6838 (N_6838,N_6508,N_6669);
nand U6839 (N_6839,N_6408,N_6700);
nor U6840 (N_6840,N_6181,N_6641);
nand U6841 (N_6841,N_6383,N_6461);
nor U6842 (N_6842,N_6313,N_6605);
or U6843 (N_6843,N_6149,N_6433);
or U6844 (N_6844,N_6654,N_6658);
nor U6845 (N_6845,N_6006,N_6402);
nand U6846 (N_6846,N_6523,N_6645);
or U6847 (N_6847,N_6358,N_6345);
nor U6848 (N_6848,N_6271,N_6117);
and U6849 (N_6849,N_6265,N_6354);
or U6850 (N_6850,N_6630,N_6622);
or U6851 (N_6851,N_6094,N_6106);
nor U6852 (N_6852,N_6390,N_6280);
nor U6853 (N_6853,N_6397,N_6312);
or U6854 (N_6854,N_6393,N_6307);
xor U6855 (N_6855,N_6259,N_6388);
nand U6856 (N_6856,N_6509,N_6466);
nand U6857 (N_6857,N_6631,N_6514);
nand U6858 (N_6858,N_6132,N_6378);
and U6859 (N_6859,N_6215,N_6501);
and U6860 (N_6860,N_6450,N_6657);
or U6861 (N_6861,N_6073,N_6420);
or U6862 (N_6862,N_6178,N_6099);
and U6863 (N_6863,N_6115,N_6136);
and U6864 (N_6864,N_6126,N_6047);
nand U6865 (N_6865,N_6018,N_6382);
nor U6866 (N_6866,N_6148,N_6238);
nor U6867 (N_6867,N_6218,N_6696);
and U6868 (N_6868,N_6144,N_6502);
and U6869 (N_6869,N_6529,N_6524);
xor U6870 (N_6870,N_6212,N_6160);
and U6871 (N_6871,N_6617,N_6723);
nor U6872 (N_6872,N_6556,N_6193);
nand U6873 (N_6873,N_6424,N_6276);
nor U6874 (N_6874,N_6169,N_6076);
and U6875 (N_6875,N_6442,N_6642);
and U6876 (N_6876,N_6142,N_6405);
and U6877 (N_6877,N_6356,N_6463);
nand U6878 (N_6878,N_6747,N_6582);
and U6879 (N_6879,N_6471,N_6085);
or U6880 (N_6880,N_6448,N_6665);
or U6881 (N_6881,N_6092,N_6166);
nand U6882 (N_6882,N_6161,N_6086);
nor U6883 (N_6883,N_6025,N_6071);
xnor U6884 (N_6884,N_6320,N_6718);
nor U6885 (N_6885,N_6328,N_6046);
and U6886 (N_6886,N_6319,N_6596);
nand U6887 (N_6887,N_6282,N_6745);
nor U6888 (N_6888,N_6703,N_6585);
or U6889 (N_6889,N_6573,N_6014);
or U6890 (N_6890,N_6139,N_6588);
nor U6891 (N_6891,N_6667,N_6674);
nor U6892 (N_6892,N_6070,N_6278);
and U6893 (N_6893,N_6209,N_6162);
nor U6894 (N_6894,N_6188,N_6043);
nor U6895 (N_6895,N_6299,N_6118);
and U6896 (N_6896,N_6264,N_6474);
and U6897 (N_6897,N_6515,N_6741);
or U6898 (N_6898,N_6710,N_6203);
nor U6899 (N_6899,N_6101,N_6038);
nor U6900 (N_6900,N_6493,N_6512);
nor U6901 (N_6901,N_6399,N_6749);
nand U6902 (N_6902,N_6469,N_6322);
and U6903 (N_6903,N_6223,N_6639);
and U6904 (N_6904,N_6398,N_6233);
xor U6905 (N_6905,N_6274,N_6505);
and U6906 (N_6906,N_6643,N_6513);
nand U6907 (N_6907,N_6396,N_6740);
nor U6908 (N_6908,N_6575,N_6034);
nor U6909 (N_6909,N_6421,N_6155);
or U6910 (N_6910,N_6141,N_6200);
nand U6911 (N_6911,N_6434,N_6739);
nand U6912 (N_6912,N_6174,N_6462);
nand U6913 (N_6913,N_6122,N_6445);
or U6914 (N_6914,N_6656,N_6375);
and U6915 (N_6915,N_6123,N_6748);
and U6916 (N_6916,N_6459,N_6673);
and U6917 (N_6917,N_6330,N_6392);
nand U6918 (N_6918,N_6247,N_6563);
and U6919 (N_6919,N_6171,N_6510);
and U6920 (N_6920,N_6647,N_6498);
and U6921 (N_6921,N_6734,N_6578);
nand U6922 (N_6922,N_6571,N_6694);
xnor U6923 (N_6923,N_6614,N_6332);
and U6924 (N_6924,N_6379,N_6693);
or U6925 (N_6925,N_6222,N_6706);
or U6926 (N_6926,N_6341,N_6608);
nand U6927 (N_6927,N_6198,N_6389);
nand U6928 (N_6928,N_6022,N_6598);
nor U6929 (N_6929,N_6154,N_6587);
nand U6930 (N_6930,N_6054,N_6208);
xnor U6931 (N_6931,N_6191,N_6444);
nand U6932 (N_6932,N_6579,N_6300);
or U6933 (N_6933,N_6082,N_6661);
or U6934 (N_6934,N_6285,N_6439);
and U6935 (N_6935,N_6480,N_6727);
nand U6936 (N_6936,N_6065,N_6467);
and U6937 (N_6937,N_6488,N_6164);
or U6938 (N_6938,N_6202,N_6296);
nor U6939 (N_6939,N_6530,N_6194);
nand U6940 (N_6940,N_6053,N_6580);
and U6941 (N_6941,N_6702,N_6093);
or U6942 (N_6942,N_6534,N_6275);
or U6943 (N_6943,N_6409,N_6125);
nor U6944 (N_6944,N_6489,N_6416);
and U6945 (N_6945,N_6260,N_6419);
or U6946 (N_6946,N_6359,N_6360);
nor U6947 (N_6947,N_6283,N_6242);
and U6948 (N_6948,N_6310,N_6726);
xnor U6949 (N_6949,N_6365,N_6464);
nor U6950 (N_6950,N_6120,N_6102);
nand U6951 (N_6951,N_6342,N_6066);
or U6952 (N_6952,N_6699,N_6562);
or U6953 (N_6953,N_6227,N_6583);
or U6954 (N_6954,N_6104,N_6019);
and U6955 (N_6955,N_6546,N_6255);
or U6956 (N_6956,N_6431,N_6543);
or U6957 (N_6957,N_6293,N_6733);
nor U6958 (N_6958,N_6499,N_6644);
nor U6959 (N_6959,N_6716,N_6432);
and U6960 (N_6960,N_6204,N_6349);
nand U6961 (N_6961,N_6151,N_6056);
or U6962 (N_6962,N_6294,N_6369);
nor U6963 (N_6963,N_6150,N_6001);
and U6964 (N_6964,N_6652,N_6052);
and U6965 (N_6965,N_6173,N_6340);
nand U6966 (N_6966,N_6176,N_6632);
and U6967 (N_6967,N_6621,N_6192);
or U6968 (N_6968,N_6245,N_6552);
or U6969 (N_6969,N_6027,N_6243);
and U6970 (N_6970,N_6681,N_6059);
nor U6971 (N_6971,N_6334,N_6361);
and U6972 (N_6972,N_6229,N_6346);
nor U6973 (N_6973,N_6485,N_6298);
and U6974 (N_6974,N_6020,N_6446);
or U6975 (N_6975,N_6069,N_6314);
nor U6976 (N_6976,N_6691,N_6533);
nand U6977 (N_6977,N_6504,N_6447);
and U6978 (N_6978,N_6207,N_6683);
or U6979 (N_6979,N_6281,N_6412);
or U6980 (N_6980,N_6475,N_6355);
nor U6981 (N_6981,N_6627,N_6411);
nand U6982 (N_6982,N_6558,N_6152);
nor U6983 (N_6983,N_6074,N_6483);
xor U6984 (N_6984,N_6600,N_6590);
or U6985 (N_6985,N_6028,N_6137);
or U6986 (N_6986,N_6550,N_6484);
nand U6987 (N_6987,N_6228,N_6135);
nor U6988 (N_6988,N_6476,N_6079);
or U6989 (N_6989,N_6743,N_6165);
and U6990 (N_6990,N_6317,N_6520);
nand U6991 (N_6991,N_6067,N_6257);
and U6992 (N_6992,N_6607,N_6440);
or U6993 (N_6993,N_6269,N_6680);
xor U6994 (N_6994,N_6068,N_6338);
xnor U6995 (N_6995,N_6324,N_6635);
and U6996 (N_6996,N_6468,N_6692);
nor U6997 (N_6997,N_6190,N_6205);
and U6998 (N_6998,N_6235,N_6538);
or U6999 (N_6999,N_6131,N_6687);
and U7000 (N_7000,N_6103,N_6717);
nor U7001 (N_7001,N_6072,N_6250);
nor U7002 (N_7002,N_6521,N_6670);
or U7003 (N_7003,N_6251,N_6620);
or U7004 (N_7004,N_6413,N_6403);
nand U7005 (N_7005,N_6236,N_6089);
nor U7006 (N_7006,N_6666,N_6128);
nor U7007 (N_7007,N_6437,N_6316);
nor U7008 (N_7008,N_6367,N_6415);
or U7009 (N_7009,N_6244,N_6597);
or U7010 (N_7010,N_6516,N_6185);
and U7011 (N_7011,N_6363,N_6517);
and U7012 (N_7012,N_6567,N_6377);
nor U7013 (N_7013,N_6490,N_6574);
and U7014 (N_7014,N_6532,N_6343);
nor U7015 (N_7015,N_6586,N_6374);
nor U7016 (N_7016,N_6177,N_6357);
nand U7017 (N_7017,N_6252,N_6719);
nor U7018 (N_7018,N_6629,N_6551);
and U7019 (N_7019,N_6569,N_6036);
and U7020 (N_7020,N_6675,N_6714);
nor U7021 (N_7021,N_6272,N_6147);
and U7022 (N_7022,N_6385,N_6453);
nand U7023 (N_7023,N_6449,N_6662);
nor U7024 (N_7024,N_6648,N_6602);
and U7025 (N_7025,N_6540,N_6309);
and U7026 (N_7026,N_6715,N_6081);
and U7027 (N_7027,N_6729,N_6159);
or U7028 (N_7028,N_6091,N_6619);
nor U7029 (N_7029,N_6492,N_6087);
nand U7030 (N_7030,N_6592,N_6436);
nor U7031 (N_7031,N_6058,N_6109);
nor U7032 (N_7032,N_6040,N_6685);
or U7033 (N_7033,N_6344,N_6725);
nand U7034 (N_7034,N_6370,N_6261);
nand U7035 (N_7035,N_6042,N_6311);
nor U7036 (N_7036,N_6545,N_6451);
nand U7037 (N_7037,N_6287,N_6507);
nand U7038 (N_7038,N_6146,N_6465);
and U7039 (N_7039,N_6031,N_6143);
or U7040 (N_7040,N_6084,N_6007);
nor U7041 (N_7041,N_6015,N_6110);
xnor U7042 (N_7042,N_6486,N_6051);
or U7043 (N_7043,N_6628,N_6288);
or U7044 (N_7044,N_6004,N_6555);
nand U7045 (N_7045,N_6494,N_6731);
and U7046 (N_7046,N_6225,N_6183);
nor U7047 (N_7047,N_6239,N_6163);
nand U7048 (N_7048,N_6609,N_6037);
nor U7049 (N_7049,N_6708,N_6487);
and U7050 (N_7050,N_6746,N_6024);
or U7051 (N_7051,N_6441,N_6735);
nand U7052 (N_7052,N_6728,N_6124);
and U7053 (N_7053,N_6286,N_6526);
nor U7054 (N_7054,N_6277,N_6495);
and U7055 (N_7055,N_6653,N_6064);
and U7056 (N_7056,N_6153,N_6472);
nor U7057 (N_7057,N_6134,N_6479);
and U7058 (N_7058,N_6246,N_6097);
nor U7059 (N_7059,N_6172,N_6353);
xor U7060 (N_7060,N_6659,N_6721);
nand U7061 (N_7061,N_6688,N_6201);
nor U7062 (N_7062,N_6531,N_6537);
nand U7063 (N_7063,N_6075,N_6584);
and U7064 (N_7064,N_6333,N_6230);
or U7065 (N_7065,N_6649,N_6268);
nand U7066 (N_7066,N_6100,N_6496);
nand U7067 (N_7067,N_6689,N_6564);
nand U7068 (N_7068,N_6189,N_6427);
nor U7069 (N_7069,N_6565,N_6525);
and U7070 (N_7070,N_6373,N_6624);
nor U7071 (N_7071,N_6722,N_6595);
nor U7072 (N_7072,N_6170,N_6712);
nand U7073 (N_7073,N_6032,N_6387);
nand U7074 (N_7074,N_6195,N_6481);
or U7075 (N_7075,N_6664,N_6676);
nor U7076 (N_7076,N_6672,N_6615);
or U7077 (N_7077,N_6057,N_6133);
nand U7078 (N_7078,N_6503,N_6241);
nor U7079 (N_7079,N_6035,N_6429);
nand U7080 (N_7080,N_6697,N_6572);
nor U7081 (N_7081,N_6216,N_6138);
or U7082 (N_7082,N_6112,N_6351);
nand U7083 (N_7083,N_6273,N_6290);
nand U7084 (N_7084,N_6589,N_6121);
nor U7085 (N_7085,N_6026,N_6518);
or U7086 (N_7086,N_6184,N_6318);
or U7087 (N_7087,N_6366,N_6640);
nand U7088 (N_7088,N_6435,N_6500);
and U7089 (N_7089,N_6690,N_6352);
nor U7090 (N_7090,N_6519,N_6482);
nand U7091 (N_7091,N_6129,N_6425);
and U7092 (N_7092,N_6083,N_6206);
nor U7093 (N_7093,N_6156,N_6695);
xor U7094 (N_7094,N_6292,N_6308);
and U7095 (N_7095,N_6612,N_6167);
xor U7096 (N_7096,N_6604,N_6003);
nor U7097 (N_7097,N_6088,N_6591);
and U7098 (N_7098,N_6577,N_6210);
xnor U7099 (N_7099,N_6686,N_6033);
or U7100 (N_7100,N_6158,N_6742);
and U7101 (N_7101,N_6438,N_6705);
and U7102 (N_7102,N_6458,N_6199);
and U7103 (N_7103,N_6634,N_6080);
nor U7104 (N_7104,N_6008,N_6217);
nand U7105 (N_7105,N_6613,N_6454);
or U7106 (N_7106,N_6011,N_6301);
and U7107 (N_7107,N_6041,N_6548);
xnor U7108 (N_7108,N_6593,N_6497);
or U7109 (N_7109,N_6180,N_6329);
nand U7110 (N_7110,N_6455,N_6581);
nor U7111 (N_7111,N_6528,N_6350);
xor U7112 (N_7112,N_6709,N_6376);
or U7113 (N_7113,N_6707,N_6737);
or U7114 (N_7114,N_6452,N_6724);
or U7115 (N_7115,N_6336,N_6029);
nor U7116 (N_7116,N_6049,N_6111);
and U7117 (N_7117,N_6060,N_6650);
and U7118 (N_7118,N_6418,N_6544);
or U7119 (N_7119,N_6407,N_6606);
and U7120 (N_7120,N_6443,N_6633);
or U7121 (N_7121,N_6231,N_6175);
nor U7122 (N_7122,N_6711,N_6262);
nor U7123 (N_7123,N_6663,N_6623);
and U7124 (N_7124,N_6601,N_6384);
or U7125 (N_7125,N_6118,N_6616);
and U7126 (N_7126,N_6525,N_6478);
and U7127 (N_7127,N_6027,N_6041);
or U7128 (N_7128,N_6186,N_6337);
nor U7129 (N_7129,N_6439,N_6101);
or U7130 (N_7130,N_6654,N_6085);
and U7131 (N_7131,N_6142,N_6138);
nor U7132 (N_7132,N_6442,N_6567);
nand U7133 (N_7133,N_6233,N_6188);
and U7134 (N_7134,N_6447,N_6401);
and U7135 (N_7135,N_6629,N_6001);
or U7136 (N_7136,N_6571,N_6423);
nand U7137 (N_7137,N_6169,N_6402);
nand U7138 (N_7138,N_6327,N_6034);
nor U7139 (N_7139,N_6356,N_6548);
and U7140 (N_7140,N_6275,N_6713);
nand U7141 (N_7141,N_6394,N_6163);
or U7142 (N_7142,N_6546,N_6330);
nor U7143 (N_7143,N_6339,N_6129);
xnor U7144 (N_7144,N_6614,N_6663);
and U7145 (N_7145,N_6254,N_6710);
or U7146 (N_7146,N_6606,N_6245);
or U7147 (N_7147,N_6334,N_6167);
and U7148 (N_7148,N_6371,N_6635);
nand U7149 (N_7149,N_6388,N_6482);
nand U7150 (N_7150,N_6250,N_6635);
or U7151 (N_7151,N_6686,N_6325);
nand U7152 (N_7152,N_6325,N_6684);
and U7153 (N_7153,N_6585,N_6144);
or U7154 (N_7154,N_6211,N_6043);
nor U7155 (N_7155,N_6078,N_6603);
nand U7156 (N_7156,N_6597,N_6513);
or U7157 (N_7157,N_6511,N_6394);
and U7158 (N_7158,N_6076,N_6064);
or U7159 (N_7159,N_6637,N_6506);
nand U7160 (N_7160,N_6716,N_6245);
nor U7161 (N_7161,N_6693,N_6647);
nor U7162 (N_7162,N_6171,N_6396);
nand U7163 (N_7163,N_6206,N_6387);
nor U7164 (N_7164,N_6280,N_6377);
nor U7165 (N_7165,N_6740,N_6364);
nand U7166 (N_7166,N_6057,N_6576);
and U7167 (N_7167,N_6688,N_6650);
and U7168 (N_7168,N_6189,N_6364);
and U7169 (N_7169,N_6397,N_6283);
or U7170 (N_7170,N_6637,N_6600);
and U7171 (N_7171,N_6224,N_6582);
nand U7172 (N_7172,N_6492,N_6030);
nor U7173 (N_7173,N_6707,N_6062);
and U7174 (N_7174,N_6408,N_6171);
and U7175 (N_7175,N_6125,N_6695);
and U7176 (N_7176,N_6110,N_6364);
nand U7177 (N_7177,N_6476,N_6690);
nand U7178 (N_7178,N_6225,N_6721);
and U7179 (N_7179,N_6418,N_6709);
or U7180 (N_7180,N_6108,N_6623);
nor U7181 (N_7181,N_6616,N_6225);
nand U7182 (N_7182,N_6157,N_6271);
xnor U7183 (N_7183,N_6036,N_6621);
nand U7184 (N_7184,N_6668,N_6483);
nand U7185 (N_7185,N_6164,N_6037);
nand U7186 (N_7186,N_6394,N_6134);
nor U7187 (N_7187,N_6340,N_6694);
and U7188 (N_7188,N_6552,N_6419);
and U7189 (N_7189,N_6339,N_6523);
and U7190 (N_7190,N_6622,N_6106);
or U7191 (N_7191,N_6552,N_6537);
and U7192 (N_7192,N_6165,N_6485);
nand U7193 (N_7193,N_6153,N_6474);
and U7194 (N_7194,N_6593,N_6268);
or U7195 (N_7195,N_6399,N_6696);
nand U7196 (N_7196,N_6476,N_6164);
nor U7197 (N_7197,N_6619,N_6268);
or U7198 (N_7198,N_6646,N_6597);
nor U7199 (N_7199,N_6420,N_6153);
or U7200 (N_7200,N_6211,N_6624);
nand U7201 (N_7201,N_6449,N_6282);
nand U7202 (N_7202,N_6557,N_6492);
nor U7203 (N_7203,N_6148,N_6581);
and U7204 (N_7204,N_6140,N_6435);
or U7205 (N_7205,N_6080,N_6387);
nor U7206 (N_7206,N_6655,N_6132);
or U7207 (N_7207,N_6129,N_6052);
nor U7208 (N_7208,N_6186,N_6319);
nand U7209 (N_7209,N_6129,N_6541);
or U7210 (N_7210,N_6493,N_6135);
nor U7211 (N_7211,N_6224,N_6029);
nand U7212 (N_7212,N_6403,N_6658);
and U7213 (N_7213,N_6480,N_6585);
nor U7214 (N_7214,N_6245,N_6200);
and U7215 (N_7215,N_6695,N_6191);
nor U7216 (N_7216,N_6658,N_6054);
nand U7217 (N_7217,N_6577,N_6617);
and U7218 (N_7218,N_6269,N_6225);
and U7219 (N_7219,N_6737,N_6548);
or U7220 (N_7220,N_6247,N_6267);
nor U7221 (N_7221,N_6143,N_6095);
nor U7222 (N_7222,N_6158,N_6427);
or U7223 (N_7223,N_6154,N_6234);
and U7224 (N_7224,N_6427,N_6478);
nand U7225 (N_7225,N_6523,N_6033);
and U7226 (N_7226,N_6149,N_6230);
and U7227 (N_7227,N_6591,N_6124);
nand U7228 (N_7228,N_6457,N_6102);
nor U7229 (N_7229,N_6223,N_6510);
and U7230 (N_7230,N_6554,N_6695);
nor U7231 (N_7231,N_6544,N_6196);
and U7232 (N_7232,N_6299,N_6000);
nand U7233 (N_7233,N_6232,N_6033);
nand U7234 (N_7234,N_6045,N_6497);
or U7235 (N_7235,N_6082,N_6152);
and U7236 (N_7236,N_6564,N_6073);
or U7237 (N_7237,N_6384,N_6294);
nor U7238 (N_7238,N_6521,N_6128);
and U7239 (N_7239,N_6312,N_6642);
nor U7240 (N_7240,N_6077,N_6495);
and U7241 (N_7241,N_6672,N_6612);
nor U7242 (N_7242,N_6030,N_6516);
nand U7243 (N_7243,N_6150,N_6103);
nor U7244 (N_7244,N_6388,N_6543);
nand U7245 (N_7245,N_6274,N_6057);
nand U7246 (N_7246,N_6521,N_6156);
or U7247 (N_7247,N_6009,N_6176);
nor U7248 (N_7248,N_6579,N_6276);
nand U7249 (N_7249,N_6572,N_6737);
or U7250 (N_7250,N_6363,N_6663);
nor U7251 (N_7251,N_6741,N_6165);
nand U7252 (N_7252,N_6288,N_6304);
and U7253 (N_7253,N_6567,N_6383);
or U7254 (N_7254,N_6397,N_6294);
nand U7255 (N_7255,N_6441,N_6716);
nor U7256 (N_7256,N_6530,N_6686);
nand U7257 (N_7257,N_6346,N_6591);
nand U7258 (N_7258,N_6681,N_6047);
or U7259 (N_7259,N_6536,N_6288);
and U7260 (N_7260,N_6227,N_6550);
nand U7261 (N_7261,N_6123,N_6508);
and U7262 (N_7262,N_6514,N_6294);
nand U7263 (N_7263,N_6231,N_6015);
xor U7264 (N_7264,N_6589,N_6741);
nand U7265 (N_7265,N_6212,N_6357);
nand U7266 (N_7266,N_6472,N_6441);
nor U7267 (N_7267,N_6148,N_6469);
nand U7268 (N_7268,N_6563,N_6627);
and U7269 (N_7269,N_6415,N_6193);
or U7270 (N_7270,N_6133,N_6320);
nand U7271 (N_7271,N_6456,N_6701);
nand U7272 (N_7272,N_6432,N_6453);
and U7273 (N_7273,N_6687,N_6290);
or U7274 (N_7274,N_6033,N_6456);
and U7275 (N_7275,N_6672,N_6150);
or U7276 (N_7276,N_6329,N_6702);
and U7277 (N_7277,N_6573,N_6283);
nand U7278 (N_7278,N_6130,N_6129);
and U7279 (N_7279,N_6708,N_6005);
nand U7280 (N_7280,N_6579,N_6527);
nor U7281 (N_7281,N_6735,N_6538);
nor U7282 (N_7282,N_6574,N_6122);
and U7283 (N_7283,N_6229,N_6030);
nand U7284 (N_7284,N_6130,N_6246);
xor U7285 (N_7285,N_6397,N_6158);
or U7286 (N_7286,N_6557,N_6352);
and U7287 (N_7287,N_6203,N_6536);
xor U7288 (N_7288,N_6098,N_6466);
nor U7289 (N_7289,N_6588,N_6464);
and U7290 (N_7290,N_6547,N_6027);
and U7291 (N_7291,N_6436,N_6051);
nand U7292 (N_7292,N_6277,N_6312);
nor U7293 (N_7293,N_6672,N_6010);
nand U7294 (N_7294,N_6680,N_6370);
nand U7295 (N_7295,N_6581,N_6434);
nor U7296 (N_7296,N_6320,N_6581);
nand U7297 (N_7297,N_6067,N_6331);
nand U7298 (N_7298,N_6253,N_6404);
or U7299 (N_7299,N_6075,N_6555);
nand U7300 (N_7300,N_6043,N_6396);
and U7301 (N_7301,N_6028,N_6549);
or U7302 (N_7302,N_6477,N_6348);
nor U7303 (N_7303,N_6598,N_6311);
or U7304 (N_7304,N_6053,N_6271);
or U7305 (N_7305,N_6320,N_6097);
nand U7306 (N_7306,N_6346,N_6040);
nand U7307 (N_7307,N_6307,N_6636);
nand U7308 (N_7308,N_6412,N_6349);
xor U7309 (N_7309,N_6134,N_6027);
nor U7310 (N_7310,N_6193,N_6419);
nand U7311 (N_7311,N_6052,N_6083);
nor U7312 (N_7312,N_6169,N_6262);
nor U7313 (N_7313,N_6627,N_6707);
or U7314 (N_7314,N_6253,N_6324);
and U7315 (N_7315,N_6315,N_6418);
nand U7316 (N_7316,N_6694,N_6537);
xnor U7317 (N_7317,N_6135,N_6697);
nor U7318 (N_7318,N_6442,N_6439);
or U7319 (N_7319,N_6053,N_6323);
nand U7320 (N_7320,N_6037,N_6044);
xor U7321 (N_7321,N_6317,N_6169);
and U7322 (N_7322,N_6011,N_6302);
and U7323 (N_7323,N_6147,N_6153);
or U7324 (N_7324,N_6098,N_6628);
nor U7325 (N_7325,N_6539,N_6310);
nor U7326 (N_7326,N_6706,N_6399);
and U7327 (N_7327,N_6114,N_6351);
and U7328 (N_7328,N_6208,N_6197);
nand U7329 (N_7329,N_6563,N_6723);
or U7330 (N_7330,N_6425,N_6369);
and U7331 (N_7331,N_6073,N_6612);
nor U7332 (N_7332,N_6425,N_6017);
or U7333 (N_7333,N_6107,N_6330);
nand U7334 (N_7334,N_6566,N_6463);
nor U7335 (N_7335,N_6309,N_6581);
or U7336 (N_7336,N_6197,N_6155);
nor U7337 (N_7337,N_6295,N_6467);
nand U7338 (N_7338,N_6404,N_6485);
xor U7339 (N_7339,N_6257,N_6035);
nor U7340 (N_7340,N_6298,N_6255);
or U7341 (N_7341,N_6425,N_6507);
and U7342 (N_7342,N_6084,N_6554);
xor U7343 (N_7343,N_6140,N_6540);
nor U7344 (N_7344,N_6334,N_6554);
and U7345 (N_7345,N_6477,N_6749);
and U7346 (N_7346,N_6582,N_6559);
nand U7347 (N_7347,N_6113,N_6621);
and U7348 (N_7348,N_6106,N_6515);
or U7349 (N_7349,N_6562,N_6579);
and U7350 (N_7350,N_6598,N_6696);
nand U7351 (N_7351,N_6183,N_6066);
nor U7352 (N_7352,N_6171,N_6588);
and U7353 (N_7353,N_6729,N_6302);
nor U7354 (N_7354,N_6746,N_6514);
nand U7355 (N_7355,N_6081,N_6366);
nor U7356 (N_7356,N_6693,N_6319);
nor U7357 (N_7357,N_6629,N_6609);
or U7358 (N_7358,N_6718,N_6625);
nor U7359 (N_7359,N_6704,N_6219);
nor U7360 (N_7360,N_6193,N_6715);
nand U7361 (N_7361,N_6364,N_6527);
nand U7362 (N_7362,N_6048,N_6707);
and U7363 (N_7363,N_6029,N_6615);
and U7364 (N_7364,N_6067,N_6729);
nor U7365 (N_7365,N_6428,N_6125);
nand U7366 (N_7366,N_6288,N_6339);
nor U7367 (N_7367,N_6461,N_6214);
or U7368 (N_7368,N_6221,N_6680);
and U7369 (N_7369,N_6391,N_6107);
and U7370 (N_7370,N_6251,N_6279);
and U7371 (N_7371,N_6393,N_6697);
nor U7372 (N_7372,N_6570,N_6126);
xor U7373 (N_7373,N_6283,N_6725);
nor U7374 (N_7374,N_6411,N_6287);
nor U7375 (N_7375,N_6687,N_6723);
nand U7376 (N_7376,N_6522,N_6104);
nand U7377 (N_7377,N_6479,N_6545);
nand U7378 (N_7378,N_6396,N_6395);
or U7379 (N_7379,N_6667,N_6135);
and U7380 (N_7380,N_6312,N_6327);
and U7381 (N_7381,N_6328,N_6325);
or U7382 (N_7382,N_6443,N_6053);
and U7383 (N_7383,N_6206,N_6332);
nor U7384 (N_7384,N_6357,N_6232);
and U7385 (N_7385,N_6164,N_6571);
or U7386 (N_7386,N_6678,N_6612);
nand U7387 (N_7387,N_6593,N_6010);
or U7388 (N_7388,N_6550,N_6666);
and U7389 (N_7389,N_6688,N_6410);
nand U7390 (N_7390,N_6188,N_6494);
nor U7391 (N_7391,N_6098,N_6151);
and U7392 (N_7392,N_6329,N_6617);
nor U7393 (N_7393,N_6635,N_6316);
nor U7394 (N_7394,N_6476,N_6587);
or U7395 (N_7395,N_6528,N_6223);
nor U7396 (N_7396,N_6280,N_6685);
or U7397 (N_7397,N_6269,N_6623);
and U7398 (N_7398,N_6511,N_6644);
or U7399 (N_7399,N_6410,N_6026);
nor U7400 (N_7400,N_6114,N_6731);
and U7401 (N_7401,N_6071,N_6394);
nor U7402 (N_7402,N_6714,N_6634);
nor U7403 (N_7403,N_6585,N_6111);
xnor U7404 (N_7404,N_6175,N_6551);
nor U7405 (N_7405,N_6363,N_6665);
nand U7406 (N_7406,N_6127,N_6230);
or U7407 (N_7407,N_6625,N_6464);
nor U7408 (N_7408,N_6475,N_6351);
and U7409 (N_7409,N_6718,N_6179);
and U7410 (N_7410,N_6567,N_6267);
nor U7411 (N_7411,N_6711,N_6045);
nor U7412 (N_7412,N_6138,N_6600);
and U7413 (N_7413,N_6141,N_6013);
and U7414 (N_7414,N_6450,N_6567);
nor U7415 (N_7415,N_6204,N_6368);
and U7416 (N_7416,N_6677,N_6190);
nor U7417 (N_7417,N_6171,N_6137);
or U7418 (N_7418,N_6311,N_6323);
nor U7419 (N_7419,N_6538,N_6363);
or U7420 (N_7420,N_6662,N_6738);
and U7421 (N_7421,N_6671,N_6747);
nor U7422 (N_7422,N_6253,N_6452);
xnor U7423 (N_7423,N_6474,N_6452);
nor U7424 (N_7424,N_6581,N_6670);
nand U7425 (N_7425,N_6713,N_6254);
or U7426 (N_7426,N_6311,N_6154);
or U7427 (N_7427,N_6376,N_6483);
xnor U7428 (N_7428,N_6546,N_6632);
and U7429 (N_7429,N_6061,N_6433);
nor U7430 (N_7430,N_6371,N_6391);
nor U7431 (N_7431,N_6283,N_6413);
or U7432 (N_7432,N_6365,N_6656);
nand U7433 (N_7433,N_6551,N_6527);
or U7434 (N_7434,N_6472,N_6525);
nand U7435 (N_7435,N_6074,N_6361);
nor U7436 (N_7436,N_6166,N_6422);
and U7437 (N_7437,N_6593,N_6106);
nor U7438 (N_7438,N_6093,N_6404);
and U7439 (N_7439,N_6223,N_6549);
nor U7440 (N_7440,N_6395,N_6009);
and U7441 (N_7441,N_6465,N_6178);
xnor U7442 (N_7442,N_6599,N_6372);
nor U7443 (N_7443,N_6642,N_6368);
xnor U7444 (N_7444,N_6493,N_6056);
nand U7445 (N_7445,N_6422,N_6694);
and U7446 (N_7446,N_6412,N_6051);
nor U7447 (N_7447,N_6204,N_6481);
or U7448 (N_7448,N_6133,N_6151);
or U7449 (N_7449,N_6580,N_6079);
nor U7450 (N_7450,N_6306,N_6278);
nand U7451 (N_7451,N_6524,N_6062);
nor U7452 (N_7452,N_6110,N_6188);
nor U7453 (N_7453,N_6600,N_6189);
nor U7454 (N_7454,N_6315,N_6554);
or U7455 (N_7455,N_6244,N_6629);
nor U7456 (N_7456,N_6364,N_6709);
or U7457 (N_7457,N_6697,N_6048);
or U7458 (N_7458,N_6424,N_6577);
and U7459 (N_7459,N_6220,N_6343);
or U7460 (N_7460,N_6241,N_6474);
and U7461 (N_7461,N_6277,N_6434);
nand U7462 (N_7462,N_6587,N_6226);
or U7463 (N_7463,N_6212,N_6508);
nand U7464 (N_7464,N_6030,N_6604);
or U7465 (N_7465,N_6611,N_6398);
and U7466 (N_7466,N_6459,N_6569);
nand U7467 (N_7467,N_6622,N_6261);
xnor U7468 (N_7468,N_6574,N_6382);
or U7469 (N_7469,N_6541,N_6683);
xor U7470 (N_7470,N_6356,N_6533);
or U7471 (N_7471,N_6101,N_6096);
nor U7472 (N_7472,N_6007,N_6281);
xor U7473 (N_7473,N_6371,N_6721);
nor U7474 (N_7474,N_6653,N_6256);
or U7475 (N_7475,N_6296,N_6123);
nor U7476 (N_7476,N_6450,N_6316);
nand U7477 (N_7477,N_6547,N_6001);
or U7478 (N_7478,N_6505,N_6086);
nor U7479 (N_7479,N_6712,N_6422);
nor U7480 (N_7480,N_6526,N_6356);
and U7481 (N_7481,N_6291,N_6475);
nor U7482 (N_7482,N_6043,N_6114);
nand U7483 (N_7483,N_6552,N_6422);
nor U7484 (N_7484,N_6520,N_6380);
nand U7485 (N_7485,N_6680,N_6734);
nand U7486 (N_7486,N_6211,N_6190);
or U7487 (N_7487,N_6068,N_6201);
nand U7488 (N_7488,N_6117,N_6353);
or U7489 (N_7489,N_6203,N_6529);
or U7490 (N_7490,N_6618,N_6597);
nand U7491 (N_7491,N_6044,N_6362);
nand U7492 (N_7492,N_6302,N_6165);
xor U7493 (N_7493,N_6501,N_6635);
and U7494 (N_7494,N_6004,N_6343);
or U7495 (N_7495,N_6671,N_6369);
nand U7496 (N_7496,N_6506,N_6232);
or U7497 (N_7497,N_6176,N_6322);
nand U7498 (N_7498,N_6454,N_6719);
or U7499 (N_7499,N_6513,N_6078);
and U7500 (N_7500,N_6908,N_6929);
nand U7501 (N_7501,N_6907,N_7064);
nand U7502 (N_7502,N_7187,N_6925);
nand U7503 (N_7503,N_6864,N_7352);
nor U7504 (N_7504,N_7129,N_7190);
nor U7505 (N_7505,N_6978,N_7109);
nand U7506 (N_7506,N_7106,N_7429);
nand U7507 (N_7507,N_7257,N_6875);
nor U7508 (N_7508,N_6847,N_7354);
nor U7509 (N_7509,N_7313,N_7138);
or U7510 (N_7510,N_7390,N_7164);
or U7511 (N_7511,N_7470,N_7386);
or U7512 (N_7512,N_6848,N_7387);
nor U7513 (N_7513,N_7249,N_7446);
and U7514 (N_7514,N_6899,N_6956);
or U7515 (N_7515,N_7443,N_7020);
and U7516 (N_7516,N_7324,N_6984);
or U7517 (N_7517,N_6814,N_7460);
nand U7518 (N_7518,N_7174,N_7241);
nand U7519 (N_7519,N_7483,N_6770);
or U7520 (N_7520,N_7439,N_7161);
and U7521 (N_7521,N_7225,N_6760);
nor U7522 (N_7522,N_7105,N_7008);
nor U7523 (N_7523,N_7277,N_7240);
or U7524 (N_7524,N_6777,N_6885);
or U7525 (N_7525,N_7166,N_7448);
and U7526 (N_7526,N_7078,N_7034);
or U7527 (N_7527,N_7067,N_7266);
and U7528 (N_7528,N_7260,N_6812);
nor U7529 (N_7529,N_6868,N_7233);
and U7530 (N_7530,N_7217,N_7373);
nand U7531 (N_7531,N_6883,N_7281);
and U7532 (N_7532,N_7419,N_7084);
or U7533 (N_7533,N_7221,N_6850);
nor U7534 (N_7534,N_7424,N_6934);
nand U7535 (N_7535,N_7017,N_7245);
nor U7536 (N_7536,N_7409,N_7335);
and U7537 (N_7537,N_6880,N_6834);
nand U7538 (N_7538,N_7082,N_7079);
or U7539 (N_7539,N_7364,N_6939);
nor U7540 (N_7540,N_7037,N_7388);
nor U7541 (N_7541,N_7278,N_6832);
and U7542 (N_7542,N_6982,N_7425);
nand U7543 (N_7543,N_7003,N_6964);
or U7544 (N_7544,N_6845,N_7494);
or U7545 (N_7545,N_7304,N_7407);
and U7546 (N_7546,N_7087,N_7308);
nand U7547 (N_7547,N_7052,N_7276);
and U7548 (N_7548,N_6961,N_6983);
and U7549 (N_7549,N_7291,N_7381);
nor U7550 (N_7550,N_7211,N_7361);
nand U7551 (N_7551,N_7431,N_7159);
or U7552 (N_7552,N_7420,N_6802);
nand U7553 (N_7553,N_7385,N_7414);
nor U7554 (N_7554,N_6954,N_7176);
nand U7555 (N_7555,N_7123,N_7263);
and U7556 (N_7556,N_6778,N_7392);
and U7557 (N_7557,N_7376,N_7061);
nand U7558 (N_7558,N_7074,N_7382);
and U7559 (N_7559,N_7297,N_7198);
or U7560 (N_7560,N_7498,N_7055);
xnor U7561 (N_7561,N_7347,N_7057);
and U7562 (N_7562,N_7230,N_7092);
xor U7563 (N_7563,N_7449,N_7294);
nor U7564 (N_7564,N_7013,N_6761);
or U7565 (N_7565,N_7345,N_7219);
and U7566 (N_7566,N_6768,N_6863);
and U7567 (N_7567,N_6857,N_7450);
or U7568 (N_7568,N_6931,N_7149);
and U7569 (N_7569,N_6957,N_6785);
nor U7570 (N_7570,N_7377,N_6915);
nor U7571 (N_7571,N_6897,N_7035);
nor U7572 (N_7572,N_7314,N_7328);
nand U7573 (N_7573,N_6909,N_7360);
or U7574 (N_7574,N_6810,N_7333);
and U7575 (N_7575,N_7243,N_7011);
and U7576 (N_7576,N_6902,N_7455);
or U7577 (N_7577,N_6945,N_7036);
or U7578 (N_7578,N_7170,N_7197);
or U7579 (N_7579,N_7027,N_7136);
or U7580 (N_7580,N_6808,N_6855);
nor U7581 (N_7581,N_7332,N_7214);
and U7582 (N_7582,N_6779,N_6865);
and U7583 (N_7583,N_7374,N_7042);
nand U7584 (N_7584,N_6927,N_7380);
and U7585 (N_7585,N_7004,N_7046);
nor U7586 (N_7586,N_7110,N_7412);
and U7587 (N_7587,N_6977,N_7065);
nand U7588 (N_7588,N_7183,N_7395);
nand U7589 (N_7589,N_7496,N_7476);
nand U7590 (N_7590,N_6963,N_7453);
or U7591 (N_7591,N_7442,N_6842);
or U7592 (N_7592,N_6753,N_7461);
and U7593 (N_7593,N_7038,N_7258);
nand U7594 (N_7594,N_7342,N_7089);
and U7595 (N_7595,N_7355,N_6971);
and U7596 (N_7596,N_7045,N_7411);
or U7597 (N_7597,N_7478,N_6936);
nor U7598 (N_7598,N_7338,N_7099);
nor U7599 (N_7599,N_7435,N_7104);
nor U7600 (N_7600,N_7306,N_6960);
nor U7601 (N_7601,N_7349,N_7244);
or U7602 (N_7602,N_6858,N_6991);
and U7603 (N_7603,N_7093,N_7485);
nor U7604 (N_7604,N_6901,N_7206);
nor U7605 (N_7605,N_7299,N_7397);
and U7606 (N_7606,N_6831,N_7154);
or U7607 (N_7607,N_6791,N_7147);
and U7608 (N_7608,N_6773,N_6935);
and U7609 (N_7609,N_6914,N_7053);
or U7610 (N_7610,N_7145,N_7083);
xnor U7611 (N_7611,N_6876,N_6943);
nand U7612 (N_7612,N_7410,N_6951);
and U7613 (N_7613,N_7076,N_6975);
or U7614 (N_7614,N_7125,N_7200);
nand U7615 (N_7615,N_7018,N_7471);
and U7616 (N_7616,N_7317,N_7199);
or U7617 (N_7617,N_7068,N_6952);
nor U7618 (N_7618,N_7408,N_6830);
or U7619 (N_7619,N_7058,N_6843);
nor U7620 (N_7620,N_7438,N_7256);
and U7621 (N_7621,N_7205,N_7457);
and U7622 (N_7622,N_7465,N_6877);
and U7623 (N_7623,N_6998,N_7007);
nand U7624 (N_7624,N_6758,N_7236);
or U7625 (N_7625,N_7116,N_7312);
nor U7626 (N_7626,N_7344,N_7177);
or U7627 (N_7627,N_7127,N_6953);
nor U7628 (N_7628,N_7456,N_7131);
and U7629 (N_7629,N_6829,N_7188);
nor U7630 (N_7630,N_6986,N_6840);
nand U7631 (N_7631,N_7142,N_7040);
or U7632 (N_7632,N_7298,N_7152);
nor U7633 (N_7633,N_7066,N_7340);
and U7634 (N_7634,N_7441,N_6837);
or U7635 (N_7635,N_7030,N_7287);
nand U7636 (N_7636,N_6805,N_6974);
nor U7637 (N_7637,N_7334,N_6890);
nor U7638 (N_7638,N_6759,N_7325);
nor U7639 (N_7639,N_7371,N_7440);
nor U7640 (N_7640,N_6860,N_7091);
and U7641 (N_7641,N_6906,N_7283);
nand U7642 (N_7642,N_6933,N_7097);
or U7643 (N_7643,N_6904,N_6809);
and U7644 (N_7644,N_7095,N_6930);
and U7645 (N_7645,N_7043,N_7228);
nand U7646 (N_7646,N_6979,N_6932);
or U7647 (N_7647,N_7051,N_7454);
nor U7648 (N_7648,N_6985,N_6879);
or U7649 (N_7649,N_6992,N_7146);
nand U7650 (N_7650,N_7015,N_6854);
and U7651 (N_7651,N_7468,N_7293);
nor U7652 (N_7652,N_7265,N_7207);
nor U7653 (N_7653,N_7148,N_7292);
nand U7654 (N_7654,N_7096,N_7447);
nor U7655 (N_7655,N_7296,N_6924);
xnor U7656 (N_7656,N_6870,N_7295);
nor U7657 (N_7657,N_6910,N_6872);
and U7658 (N_7658,N_7075,N_7196);
nand U7659 (N_7659,N_7379,N_6859);
nor U7660 (N_7660,N_7044,N_7389);
or U7661 (N_7661,N_6973,N_7466);
nor U7662 (N_7662,N_6853,N_7032);
nand U7663 (N_7663,N_7418,N_6949);
and U7664 (N_7664,N_7056,N_6962);
xnor U7665 (N_7665,N_6898,N_7318);
nor U7666 (N_7666,N_7238,N_7048);
and U7667 (N_7667,N_7237,N_6946);
nand U7668 (N_7668,N_7216,N_7417);
nand U7669 (N_7669,N_7491,N_7150);
or U7670 (N_7670,N_7289,N_7469);
nor U7671 (N_7671,N_7370,N_7156);
nor U7672 (N_7672,N_7499,N_7253);
nor U7673 (N_7673,N_6800,N_7229);
nor U7674 (N_7674,N_6981,N_7259);
xnor U7675 (N_7675,N_6969,N_7062);
nand U7676 (N_7676,N_7309,N_7002);
or U7677 (N_7677,N_6873,N_7070);
or U7678 (N_7678,N_6941,N_6866);
nand U7679 (N_7679,N_6754,N_7028);
and U7680 (N_7680,N_6839,N_6794);
or U7681 (N_7681,N_7488,N_6756);
and U7682 (N_7682,N_7479,N_7031);
nand U7683 (N_7683,N_7000,N_7366);
and U7684 (N_7684,N_7203,N_6856);
and U7685 (N_7685,N_7246,N_6913);
xnor U7686 (N_7686,N_6895,N_7358);
nand U7687 (N_7687,N_7437,N_7271);
or U7688 (N_7688,N_7365,N_6815);
or U7689 (N_7689,N_7307,N_7115);
and U7690 (N_7690,N_6938,N_6905);
nor U7691 (N_7691,N_7182,N_6900);
and U7692 (N_7692,N_6911,N_7029);
nor U7693 (N_7693,N_6995,N_6921);
and U7694 (N_7694,N_7120,N_6947);
nand U7695 (N_7695,N_7473,N_7351);
nor U7696 (N_7696,N_6793,N_7254);
nand U7697 (N_7697,N_6996,N_6869);
or U7698 (N_7698,N_6757,N_7401);
or U7699 (N_7699,N_7102,N_7047);
nand U7700 (N_7700,N_6783,N_7268);
or U7701 (N_7701,N_7239,N_6867);
nor U7702 (N_7702,N_7300,N_7195);
nor U7703 (N_7703,N_7393,N_6882);
and U7704 (N_7704,N_6811,N_6822);
nand U7705 (N_7705,N_6950,N_7305);
xor U7706 (N_7706,N_7475,N_6804);
or U7707 (N_7707,N_6862,N_6767);
or U7708 (N_7708,N_6958,N_7445);
xor U7709 (N_7709,N_7331,N_6838);
or U7710 (N_7710,N_7022,N_7321);
or U7711 (N_7711,N_7405,N_7033);
or U7712 (N_7712,N_6813,N_7353);
nand U7713 (N_7713,N_7162,N_6878);
nor U7714 (N_7714,N_7081,N_7167);
and U7715 (N_7715,N_7213,N_7073);
nand U7716 (N_7716,N_7232,N_6874);
or U7717 (N_7717,N_6766,N_6780);
nand U7718 (N_7718,N_7326,N_6891);
nor U7719 (N_7719,N_7180,N_7310);
and U7720 (N_7720,N_6942,N_7139);
and U7721 (N_7721,N_7194,N_7322);
nand U7722 (N_7722,N_7172,N_6892);
nor U7723 (N_7723,N_7141,N_6819);
and U7724 (N_7724,N_7169,N_7486);
and U7725 (N_7725,N_7208,N_7158);
nand U7726 (N_7726,N_7416,N_7143);
and U7727 (N_7727,N_7223,N_7215);
and U7728 (N_7728,N_7041,N_7252);
nor U7729 (N_7729,N_7250,N_7059);
nor U7730 (N_7730,N_7133,N_7086);
nor U7731 (N_7731,N_7359,N_6894);
nand U7732 (N_7732,N_7201,N_6786);
nand U7733 (N_7733,N_7262,N_6823);
nand U7734 (N_7734,N_6884,N_7113);
nor U7735 (N_7735,N_7130,N_6918);
or U7736 (N_7736,N_6948,N_7226);
and U7737 (N_7737,N_7436,N_7050);
and U7738 (N_7738,N_6959,N_7121);
xnor U7739 (N_7739,N_7428,N_7480);
and U7740 (N_7740,N_6789,N_6944);
nor U7741 (N_7741,N_6919,N_6955);
nor U7742 (N_7742,N_7406,N_6967);
nand U7743 (N_7743,N_7402,N_7010);
nand U7744 (N_7744,N_6887,N_6751);
and U7745 (N_7745,N_7137,N_7077);
nor U7746 (N_7746,N_6775,N_7090);
and U7747 (N_7747,N_7275,N_6787);
or U7748 (N_7748,N_6903,N_7224);
or U7749 (N_7749,N_7094,N_6806);
and U7750 (N_7750,N_7191,N_7434);
nand U7751 (N_7751,N_7490,N_7462);
and U7752 (N_7752,N_7426,N_6821);
nor U7753 (N_7753,N_7422,N_7383);
nor U7754 (N_7754,N_7181,N_7329);
or U7755 (N_7755,N_6817,N_7012);
nand U7756 (N_7756,N_7384,N_7451);
nand U7757 (N_7757,N_7069,N_7458);
nor U7758 (N_7758,N_6781,N_6797);
or U7759 (N_7759,N_6889,N_7218);
nand U7760 (N_7760,N_6990,N_7452);
and U7761 (N_7761,N_7284,N_6750);
or U7762 (N_7762,N_7220,N_7014);
xor U7763 (N_7763,N_7267,N_7101);
nor U7764 (N_7764,N_7413,N_7122);
nand U7765 (N_7765,N_7155,N_7209);
or U7766 (N_7766,N_7423,N_7492);
nand U7767 (N_7767,N_7489,N_6994);
or U7768 (N_7768,N_7088,N_7134);
and U7769 (N_7769,N_6774,N_7039);
nor U7770 (N_7770,N_7179,N_7311);
nor U7771 (N_7771,N_7135,N_7484);
and U7772 (N_7772,N_7301,N_7153);
or U7773 (N_7773,N_7171,N_7362);
and U7774 (N_7774,N_6835,N_6968);
nor U7775 (N_7775,N_6828,N_7107);
xnor U7776 (N_7776,N_6965,N_7126);
and U7777 (N_7777,N_7280,N_7071);
or U7778 (N_7778,N_7319,N_6966);
nand U7779 (N_7779,N_7339,N_6881);
or U7780 (N_7780,N_6755,N_7330);
xor U7781 (N_7781,N_6916,N_7368);
nor U7782 (N_7782,N_7023,N_7302);
nor U7783 (N_7783,N_6976,N_7118);
or U7784 (N_7784,N_7430,N_7114);
nand U7785 (N_7785,N_6997,N_7021);
nor U7786 (N_7786,N_6776,N_7274);
and U7787 (N_7787,N_6803,N_7157);
or U7788 (N_7788,N_6782,N_7119);
nor U7789 (N_7789,N_7025,N_7255);
nor U7790 (N_7790,N_7290,N_7210);
or U7791 (N_7791,N_7316,N_7320);
nor U7792 (N_7792,N_7444,N_6886);
and U7793 (N_7793,N_7235,N_6764);
nand U7794 (N_7794,N_6849,N_7098);
nor U7795 (N_7795,N_6970,N_6988);
nand U7796 (N_7796,N_7495,N_7103);
or U7797 (N_7797,N_7192,N_7341);
or U7798 (N_7798,N_7006,N_6980);
nor U7799 (N_7799,N_7100,N_7019);
nand U7800 (N_7800,N_7350,N_6861);
and U7801 (N_7801,N_6922,N_6826);
or U7802 (N_7802,N_6920,N_7282);
and U7803 (N_7803,N_6852,N_6846);
nand U7804 (N_7804,N_6771,N_7391);
and U7805 (N_7805,N_7272,N_7189);
nor U7806 (N_7806,N_7270,N_7128);
nor U7807 (N_7807,N_6763,N_6940);
and U7808 (N_7808,N_7227,N_7432);
nor U7809 (N_7809,N_7404,N_6825);
nor U7810 (N_7810,N_7242,N_7111);
nor U7811 (N_7811,N_7394,N_7024);
nand U7812 (N_7812,N_6893,N_7185);
nand U7813 (N_7813,N_6792,N_7343);
nor U7814 (N_7814,N_7348,N_7315);
nand U7815 (N_7815,N_6937,N_7202);
or U7816 (N_7816,N_7193,N_7336);
nor U7817 (N_7817,N_7163,N_7160);
and U7818 (N_7818,N_7108,N_7231);
and U7819 (N_7819,N_7165,N_7009);
nor U7820 (N_7820,N_7144,N_7178);
nor U7821 (N_7821,N_7173,N_6987);
nor U7822 (N_7822,N_7378,N_6795);
or U7823 (N_7823,N_6784,N_7112);
and U7824 (N_7824,N_7464,N_7212);
xnor U7825 (N_7825,N_7474,N_6788);
nor U7826 (N_7826,N_6807,N_7369);
nand U7827 (N_7827,N_7054,N_7399);
nand U7828 (N_7828,N_7168,N_7493);
or U7829 (N_7829,N_6841,N_7140);
and U7830 (N_7830,N_7248,N_6888);
and U7831 (N_7831,N_7049,N_6820);
and U7832 (N_7832,N_6844,N_7286);
or U7833 (N_7833,N_6836,N_7117);
and U7834 (N_7834,N_7175,N_7481);
and U7835 (N_7835,N_7497,N_7467);
nor U7836 (N_7836,N_7288,N_7415);
or U7837 (N_7837,N_6816,N_7337);
or U7838 (N_7838,N_7357,N_6798);
nand U7839 (N_7839,N_7403,N_7398);
or U7840 (N_7840,N_6824,N_7001);
or U7841 (N_7841,N_7234,N_7060);
or U7842 (N_7842,N_6801,N_7026);
or U7843 (N_7843,N_7367,N_7346);
nor U7844 (N_7844,N_6923,N_7372);
or U7845 (N_7845,N_7482,N_7072);
nor U7846 (N_7846,N_7184,N_7247);
and U7847 (N_7847,N_6851,N_7433);
nand U7848 (N_7848,N_7421,N_6818);
nand U7849 (N_7849,N_7251,N_7264);
nor U7850 (N_7850,N_6752,N_6928);
or U7851 (N_7851,N_6762,N_7327);
nor U7852 (N_7852,N_7080,N_7487);
nor U7853 (N_7853,N_7151,N_7279);
nor U7854 (N_7854,N_7222,N_6769);
nor U7855 (N_7855,N_7063,N_6972);
or U7856 (N_7856,N_7303,N_7261);
or U7857 (N_7857,N_7132,N_6772);
nand U7858 (N_7858,N_6827,N_6912);
or U7859 (N_7859,N_6799,N_7427);
nor U7860 (N_7860,N_7472,N_6926);
or U7861 (N_7861,N_6871,N_7204);
or U7862 (N_7862,N_7124,N_6790);
nand U7863 (N_7863,N_7375,N_7363);
nor U7864 (N_7864,N_6765,N_7016);
nor U7865 (N_7865,N_7463,N_6917);
nand U7866 (N_7866,N_7477,N_6993);
and U7867 (N_7867,N_7005,N_7085);
nor U7868 (N_7868,N_7459,N_6796);
and U7869 (N_7869,N_6833,N_6999);
and U7870 (N_7870,N_7285,N_7273);
or U7871 (N_7871,N_6896,N_7269);
nor U7872 (N_7872,N_6989,N_7400);
nand U7873 (N_7873,N_7396,N_7323);
nor U7874 (N_7874,N_7356,N_7186);
nor U7875 (N_7875,N_7011,N_7399);
or U7876 (N_7876,N_7251,N_6905);
nor U7877 (N_7877,N_6936,N_7247);
nand U7878 (N_7878,N_6841,N_7359);
nor U7879 (N_7879,N_7374,N_7021);
nand U7880 (N_7880,N_7046,N_6881);
or U7881 (N_7881,N_7368,N_7180);
nor U7882 (N_7882,N_7263,N_7435);
nand U7883 (N_7883,N_7192,N_6987);
nand U7884 (N_7884,N_7463,N_7124);
or U7885 (N_7885,N_7263,N_6907);
nor U7886 (N_7886,N_7080,N_7351);
and U7887 (N_7887,N_7017,N_7233);
or U7888 (N_7888,N_7007,N_6779);
and U7889 (N_7889,N_7202,N_7154);
and U7890 (N_7890,N_7099,N_7068);
nand U7891 (N_7891,N_6823,N_6866);
and U7892 (N_7892,N_7205,N_7284);
and U7893 (N_7893,N_6805,N_6876);
nor U7894 (N_7894,N_7051,N_6907);
nand U7895 (N_7895,N_7029,N_6781);
or U7896 (N_7896,N_7055,N_6831);
nor U7897 (N_7897,N_6778,N_6759);
nor U7898 (N_7898,N_7256,N_6915);
nand U7899 (N_7899,N_7308,N_7372);
and U7900 (N_7900,N_7252,N_6760);
nand U7901 (N_7901,N_7223,N_7416);
and U7902 (N_7902,N_7153,N_7474);
or U7903 (N_7903,N_6974,N_7194);
and U7904 (N_7904,N_7306,N_6966);
nor U7905 (N_7905,N_7307,N_7303);
and U7906 (N_7906,N_6815,N_7363);
nand U7907 (N_7907,N_7251,N_7480);
nor U7908 (N_7908,N_6979,N_7029);
nor U7909 (N_7909,N_7337,N_7335);
nand U7910 (N_7910,N_7007,N_7006);
nand U7911 (N_7911,N_7465,N_7464);
or U7912 (N_7912,N_7023,N_7405);
nor U7913 (N_7913,N_7212,N_7158);
or U7914 (N_7914,N_6785,N_7176);
or U7915 (N_7915,N_6792,N_6853);
and U7916 (N_7916,N_7107,N_7486);
nor U7917 (N_7917,N_7388,N_6819);
nor U7918 (N_7918,N_7257,N_6845);
nor U7919 (N_7919,N_7238,N_7480);
and U7920 (N_7920,N_7162,N_7163);
nand U7921 (N_7921,N_7087,N_7362);
or U7922 (N_7922,N_6846,N_6939);
nor U7923 (N_7923,N_7390,N_6928);
and U7924 (N_7924,N_7018,N_7380);
nor U7925 (N_7925,N_7484,N_7478);
or U7926 (N_7926,N_6797,N_7369);
nand U7927 (N_7927,N_7166,N_7412);
and U7928 (N_7928,N_7342,N_6911);
and U7929 (N_7929,N_7375,N_6925);
or U7930 (N_7930,N_6897,N_7187);
nor U7931 (N_7931,N_6908,N_7181);
nor U7932 (N_7932,N_7371,N_7332);
nor U7933 (N_7933,N_7489,N_6995);
nand U7934 (N_7934,N_7455,N_7484);
nand U7935 (N_7935,N_6753,N_6899);
or U7936 (N_7936,N_6843,N_7489);
and U7937 (N_7937,N_6890,N_7386);
and U7938 (N_7938,N_6935,N_7322);
nand U7939 (N_7939,N_7188,N_7335);
or U7940 (N_7940,N_7202,N_6949);
or U7941 (N_7941,N_7247,N_7380);
and U7942 (N_7942,N_7213,N_7248);
or U7943 (N_7943,N_7146,N_7405);
and U7944 (N_7944,N_6874,N_7491);
or U7945 (N_7945,N_7112,N_6855);
and U7946 (N_7946,N_7410,N_7158);
and U7947 (N_7947,N_7473,N_7372);
nand U7948 (N_7948,N_7327,N_7361);
and U7949 (N_7949,N_6917,N_7195);
nand U7950 (N_7950,N_6867,N_6937);
nand U7951 (N_7951,N_7153,N_7462);
nand U7952 (N_7952,N_6995,N_7001);
and U7953 (N_7953,N_6969,N_6956);
nand U7954 (N_7954,N_6934,N_7200);
or U7955 (N_7955,N_7303,N_7024);
nand U7956 (N_7956,N_7130,N_6754);
nor U7957 (N_7957,N_6887,N_6944);
and U7958 (N_7958,N_7013,N_7061);
xnor U7959 (N_7959,N_7232,N_7495);
nand U7960 (N_7960,N_7043,N_6892);
nand U7961 (N_7961,N_7140,N_7013);
nor U7962 (N_7962,N_7363,N_7008);
or U7963 (N_7963,N_6858,N_7035);
nand U7964 (N_7964,N_6813,N_7020);
and U7965 (N_7965,N_6784,N_7207);
or U7966 (N_7966,N_6927,N_7123);
and U7967 (N_7967,N_7345,N_7149);
nor U7968 (N_7968,N_7009,N_7369);
nand U7969 (N_7969,N_7278,N_7182);
and U7970 (N_7970,N_6803,N_7439);
nand U7971 (N_7971,N_6978,N_7220);
nor U7972 (N_7972,N_7260,N_7147);
nand U7973 (N_7973,N_7191,N_7246);
nand U7974 (N_7974,N_7119,N_7137);
nor U7975 (N_7975,N_6940,N_6979);
or U7976 (N_7976,N_6943,N_7320);
nand U7977 (N_7977,N_7046,N_7494);
nand U7978 (N_7978,N_6822,N_6926);
nor U7979 (N_7979,N_7242,N_7371);
or U7980 (N_7980,N_7388,N_7077);
nand U7981 (N_7981,N_6928,N_7418);
nor U7982 (N_7982,N_7130,N_6980);
or U7983 (N_7983,N_7224,N_7357);
nand U7984 (N_7984,N_7098,N_6948);
nand U7985 (N_7985,N_7148,N_6926);
xor U7986 (N_7986,N_7357,N_7427);
and U7987 (N_7987,N_7186,N_7387);
and U7988 (N_7988,N_6868,N_7426);
and U7989 (N_7989,N_7168,N_6935);
and U7990 (N_7990,N_7405,N_7202);
nand U7991 (N_7991,N_7059,N_6772);
nand U7992 (N_7992,N_6801,N_7281);
and U7993 (N_7993,N_7158,N_6759);
nand U7994 (N_7994,N_6785,N_7133);
nand U7995 (N_7995,N_7038,N_6760);
nand U7996 (N_7996,N_7170,N_7385);
nand U7997 (N_7997,N_6986,N_6984);
nor U7998 (N_7998,N_7332,N_7020);
and U7999 (N_7999,N_7099,N_7390);
nor U8000 (N_8000,N_7136,N_7126);
nor U8001 (N_8001,N_6839,N_7306);
and U8002 (N_8002,N_6790,N_7363);
or U8003 (N_8003,N_6925,N_7385);
nand U8004 (N_8004,N_7272,N_7375);
and U8005 (N_8005,N_7255,N_7234);
and U8006 (N_8006,N_7429,N_7487);
nor U8007 (N_8007,N_6778,N_7397);
and U8008 (N_8008,N_6842,N_7071);
nor U8009 (N_8009,N_6881,N_6927);
nand U8010 (N_8010,N_7234,N_7351);
nor U8011 (N_8011,N_6905,N_6932);
or U8012 (N_8012,N_6794,N_7432);
nand U8013 (N_8013,N_7290,N_7267);
nor U8014 (N_8014,N_7329,N_7011);
or U8015 (N_8015,N_7292,N_6820);
nand U8016 (N_8016,N_6949,N_6862);
nand U8017 (N_8017,N_6872,N_7390);
nor U8018 (N_8018,N_6935,N_7062);
nor U8019 (N_8019,N_6807,N_7449);
and U8020 (N_8020,N_7092,N_7109);
or U8021 (N_8021,N_7302,N_7270);
or U8022 (N_8022,N_7457,N_7024);
nor U8023 (N_8023,N_7132,N_6961);
and U8024 (N_8024,N_6972,N_6890);
and U8025 (N_8025,N_6776,N_6902);
or U8026 (N_8026,N_7112,N_7265);
nor U8027 (N_8027,N_7010,N_7482);
nor U8028 (N_8028,N_7030,N_6875);
and U8029 (N_8029,N_7157,N_6942);
nand U8030 (N_8030,N_6773,N_7122);
nor U8031 (N_8031,N_7317,N_7404);
or U8032 (N_8032,N_6775,N_7127);
nand U8033 (N_8033,N_7480,N_6754);
nand U8034 (N_8034,N_6814,N_6919);
nand U8035 (N_8035,N_7218,N_7349);
nor U8036 (N_8036,N_7302,N_6949);
nand U8037 (N_8037,N_7105,N_7427);
and U8038 (N_8038,N_7411,N_7126);
or U8039 (N_8039,N_6994,N_7243);
and U8040 (N_8040,N_6816,N_6807);
and U8041 (N_8041,N_7359,N_6851);
or U8042 (N_8042,N_7259,N_7218);
xor U8043 (N_8043,N_7137,N_7461);
nor U8044 (N_8044,N_7101,N_6989);
or U8045 (N_8045,N_7372,N_6890);
nand U8046 (N_8046,N_7296,N_7041);
and U8047 (N_8047,N_7437,N_7401);
nand U8048 (N_8048,N_7075,N_7336);
nand U8049 (N_8049,N_7461,N_6964);
and U8050 (N_8050,N_7433,N_6823);
or U8051 (N_8051,N_6821,N_6946);
nand U8052 (N_8052,N_6986,N_7152);
nor U8053 (N_8053,N_7179,N_7493);
nor U8054 (N_8054,N_6896,N_6988);
and U8055 (N_8055,N_7114,N_7177);
or U8056 (N_8056,N_6752,N_7231);
or U8057 (N_8057,N_7455,N_6763);
or U8058 (N_8058,N_6786,N_6913);
and U8059 (N_8059,N_7297,N_7054);
nand U8060 (N_8060,N_6799,N_7354);
or U8061 (N_8061,N_7347,N_7492);
nand U8062 (N_8062,N_6904,N_6902);
or U8063 (N_8063,N_7410,N_7076);
or U8064 (N_8064,N_7357,N_7082);
or U8065 (N_8065,N_6870,N_7008);
nand U8066 (N_8066,N_6777,N_6902);
nor U8067 (N_8067,N_6970,N_7426);
nor U8068 (N_8068,N_7120,N_6902);
or U8069 (N_8069,N_6833,N_7245);
nor U8070 (N_8070,N_7406,N_7055);
and U8071 (N_8071,N_7383,N_6777);
or U8072 (N_8072,N_7303,N_7374);
nor U8073 (N_8073,N_6781,N_7049);
nand U8074 (N_8074,N_7041,N_6848);
nand U8075 (N_8075,N_7026,N_6930);
nor U8076 (N_8076,N_7327,N_7430);
nand U8077 (N_8077,N_7009,N_7167);
or U8078 (N_8078,N_7284,N_7021);
or U8079 (N_8079,N_6775,N_7312);
nand U8080 (N_8080,N_6956,N_6892);
and U8081 (N_8081,N_6819,N_7206);
and U8082 (N_8082,N_7002,N_6988);
nor U8083 (N_8083,N_7311,N_7267);
nor U8084 (N_8084,N_7388,N_6987);
nand U8085 (N_8085,N_7015,N_7254);
xnor U8086 (N_8086,N_6907,N_7191);
or U8087 (N_8087,N_7206,N_6830);
nand U8088 (N_8088,N_6887,N_7110);
or U8089 (N_8089,N_6911,N_7201);
nor U8090 (N_8090,N_7497,N_7367);
or U8091 (N_8091,N_6786,N_6787);
and U8092 (N_8092,N_6767,N_7353);
and U8093 (N_8093,N_6925,N_7001);
or U8094 (N_8094,N_7090,N_7270);
and U8095 (N_8095,N_6772,N_7261);
nor U8096 (N_8096,N_6861,N_7307);
nor U8097 (N_8097,N_7405,N_7193);
and U8098 (N_8098,N_7358,N_6810);
or U8099 (N_8099,N_6925,N_7329);
nand U8100 (N_8100,N_7227,N_7405);
nand U8101 (N_8101,N_7030,N_7228);
nor U8102 (N_8102,N_7283,N_7039);
xor U8103 (N_8103,N_7003,N_7184);
nand U8104 (N_8104,N_6943,N_6804);
and U8105 (N_8105,N_7014,N_7297);
and U8106 (N_8106,N_7344,N_7205);
or U8107 (N_8107,N_7100,N_6803);
and U8108 (N_8108,N_7424,N_6770);
and U8109 (N_8109,N_7137,N_6983);
xnor U8110 (N_8110,N_6999,N_6995);
xnor U8111 (N_8111,N_6945,N_6774);
or U8112 (N_8112,N_7497,N_7249);
xnor U8113 (N_8113,N_6914,N_7251);
and U8114 (N_8114,N_7371,N_7230);
and U8115 (N_8115,N_7110,N_7028);
nor U8116 (N_8116,N_6862,N_7023);
and U8117 (N_8117,N_7127,N_6959);
or U8118 (N_8118,N_7427,N_7360);
nor U8119 (N_8119,N_7035,N_7258);
nand U8120 (N_8120,N_6786,N_6869);
nor U8121 (N_8121,N_7453,N_6923);
and U8122 (N_8122,N_6967,N_6784);
and U8123 (N_8123,N_7249,N_6780);
nand U8124 (N_8124,N_6979,N_7445);
nand U8125 (N_8125,N_7175,N_6935);
nand U8126 (N_8126,N_7446,N_6783);
and U8127 (N_8127,N_7329,N_7483);
and U8128 (N_8128,N_7180,N_7401);
and U8129 (N_8129,N_7017,N_7039);
nor U8130 (N_8130,N_7487,N_7438);
nand U8131 (N_8131,N_7338,N_7086);
nand U8132 (N_8132,N_7429,N_7100);
nand U8133 (N_8133,N_6911,N_7405);
or U8134 (N_8134,N_7192,N_7497);
and U8135 (N_8135,N_6962,N_7287);
nand U8136 (N_8136,N_7027,N_7451);
and U8137 (N_8137,N_6866,N_7494);
nor U8138 (N_8138,N_7191,N_6920);
nor U8139 (N_8139,N_7476,N_6968);
and U8140 (N_8140,N_6939,N_7367);
and U8141 (N_8141,N_6838,N_7178);
nand U8142 (N_8142,N_7124,N_7245);
and U8143 (N_8143,N_7093,N_7482);
nor U8144 (N_8144,N_7045,N_6926);
nand U8145 (N_8145,N_7334,N_7340);
and U8146 (N_8146,N_7070,N_7259);
nand U8147 (N_8147,N_6909,N_7342);
nand U8148 (N_8148,N_7482,N_6756);
or U8149 (N_8149,N_6966,N_7290);
nor U8150 (N_8150,N_7257,N_6835);
and U8151 (N_8151,N_7116,N_6837);
and U8152 (N_8152,N_7172,N_7374);
and U8153 (N_8153,N_6825,N_7198);
and U8154 (N_8154,N_6831,N_7047);
nand U8155 (N_8155,N_7498,N_6905);
nor U8156 (N_8156,N_6808,N_7115);
nor U8157 (N_8157,N_6848,N_7138);
or U8158 (N_8158,N_7037,N_6847);
and U8159 (N_8159,N_7049,N_7498);
nor U8160 (N_8160,N_7332,N_6874);
and U8161 (N_8161,N_6765,N_6943);
or U8162 (N_8162,N_7295,N_7171);
or U8163 (N_8163,N_7487,N_7267);
and U8164 (N_8164,N_7421,N_7170);
nand U8165 (N_8165,N_7268,N_7497);
nand U8166 (N_8166,N_7231,N_7456);
nor U8167 (N_8167,N_7283,N_6962);
nor U8168 (N_8168,N_7041,N_6964);
or U8169 (N_8169,N_7388,N_7380);
nor U8170 (N_8170,N_6898,N_7150);
nor U8171 (N_8171,N_6852,N_7321);
nand U8172 (N_8172,N_7191,N_6931);
or U8173 (N_8173,N_7308,N_7358);
or U8174 (N_8174,N_7198,N_7410);
nor U8175 (N_8175,N_6907,N_6932);
and U8176 (N_8176,N_7238,N_7214);
xnor U8177 (N_8177,N_6806,N_7410);
nand U8178 (N_8178,N_7043,N_6899);
xnor U8179 (N_8179,N_6928,N_7111);
or U8180 (N_8180,N_7399,N_7003);
or U8181 (N_8181,N_7472,N_7099);
or U8182 (N_8182,N_6858,N_6884);
nand U8183 (N_8183,N_6874,N_6827);
nand U8184 (N_8184,N_7140,N_7475);
nor U8185 (N_8185,N_7160,N_6839);
nor U8186 (N_8186,N_7174,N_7380);
nor U8187 (N_8187,N_7062,N_6831);
or U8188 (N_8188,N_7228,N_7493);
nor U8189 (N_8189,N_6902,N_6790);
and U8190 (N_8190,N_6984,N_6846);
nor U8191 (N_8191,N_7199,N_7127);
or U8192 (N_8192,N_7230,N_7130);
or U8193 (N_8193,N_6765,N_6776);
nor U8194 (N_8194,N_6848,N_6989);
or U8195 (N_8195,N_7328,N_7360);
and U8196 (N_8196,N_7462,N_7424);
or U8197 (N_8197,N_6886,N_7164);
or U8198 (N_8198,N_7196,N_7032);
and U8199 (N_8199,N_7062,N_7374);
and U8200 (N_8200,N_6787,N_7028);
and U8201 (N_8201,N_7263,N_7015);
or U8202 (N_8202,N_6840,N_6978);
or U8203 (N_8203,N_7197,N_7248);
and U8204 (N_8204,N_7380,N_7232);
nand U8205 (N_8205,N_6926,N_7327);
nand U8206 (N_8206,N_7414,N_6869);
or U8207 (N_8207,N_6821,N_7279);
nand U8208 (N_8208,N_6807,N_7478);
nand U8209 (N_8209,N_7406,N_6866);
nand U8210 (N_8210,N_6870,N_7046);
nand U8211 (N_8211,N_7037,N_7254);
or U8212 (N_8212,N_7377,N_6832);
or U8213 (N_8213,N_7108,N_6998);
or U8214 (N_8214,N_6946,N_6863);
nand U8215 (N_8215,N_6755,N_7031);
nand U8216 (N_8216,N_7135,N_7243);
xnor U8217 (N_8217,N_6961,N_6921);
and U8218 (N_8218,N_7452,N_6753);
and U8219 (N_8219,N_7495,N_6926);
nor U8220 (N_8220,N_7401,N_7435);
and U8221 (N_8221,N_6751,N_6775);
or U8222 (N_8222,N_7038,N_7269);
and U8223 (N_8223,N_6764,N_7448);
nor U8224 (N_8224,N_7405,N_7166);
nand U8225 (N_8225,N_7338,N_7163);
nor U8226 (N_8226,N_7420,N_7016);
nand U8227 (N_8227,N_6793,N_7388);
nor U8228 (N_8228,N_6777,N_7360);
nor U8229 (N_8229,N_6907,N_7427);
nor U8230 (N_8230,N_7109,N_7256);
and U8231 (N_8231,N_7098,N_7204);
nor U8232 (N_8232,N_7140,N_7091);
nor U8233 (N_8233,N_6827,N_6775);
nor U8234 (N_8234,N_7284,N_7302);
nor U8235 (N_8235,N_6858,N_7332);
nor U8236 (N_8236,N_7265,N_7485);
nand U8237 (N_8237,N_6776,N_7494);
nor U8238 (N_8238,N_6947,N_7065);
nor U8239 (N_8239,N_7454,N_7357);
or U8240 (N_8240,N_7158,N_6790);
xnor U8241 (N_8241,N_7024,N_7106);
or U8242 (N_8242,N_6968,N_7406);
and U8243 (N_8243,N_6843,N_7403);
and U8244 (N_8244,N_7362,N_7238);
and U8245 (N_8245,N_6924,N_6752);
nor U8246 (N_8246,N_7184,N_6911);
nor U8247 (N_8247,N_7258,N_7051);
nor U8248 (N_8248,N_6942,N_6820);
and U8249 (N_8249,N_7326,N_7155);
nor U8250 (N_8250,N_7893,N_8073);
or U8251 (N_8251,N_7941,N_8190);
and U8252 (N_8252,N_7993,N_7868);
nand U8253 (N_8253,N_7782,N_8072);
nor U8254 (N_8254,N_7953,N_7974);
nand U8255 (N_8255,N_8177,N_8076);
nand U8256 (N_8256,N_8180,N_8226);
nor U8257 (N_8257,N_7535,N_7743);
or U8258 (N_8258,N_8056,N_8128);
nand U8259 (N_8259,N_7942,N_7935);
nand U8260 (N_8260,N_7646,N_7562);
and U8261 (N_8261,N_8044,N_8142);
nand U8262 (N_8262,N_7617,N_7717);
or U8263 (N_8263,N_7614,N_7992);
nor U8264 (N_8264,N_7630,N_8018);
or U8265 (N_8265,N_8011,N_8107);
xnor U8266 (N_8266,N_8178,N_7754);
nor U8267 (N_8267,N_7628,N_7601);
or U8268 (N_8268,N_8003,N_8032);
xor U8269 (N_8269,N_7930,N_7609);
nand U8270 (N_8270,N_7862,N_7874);
nand U8271 (N_8271,N_8160,N_8227);
and U8272 (N_8272,N_8146,N_7708);
nand U8273 (N_8273,N_7904,N_7709);
and U8274 (N_8274,N_7987,N_7653);
or U8275 (N_8275,N_7787,N_8162);
nand U8276 (N_8276,N_8113,N_7737);
nor U8277 (N_8277,N_7813,N_8194);
nand U8278 (N_8278,N_8131,N_8048);
nand U8279 (N_8279,N_7903,N_8191);
and U8280 (N_8280,N_8224,N_7785);
nand U8281 (N_8281,N_7805,N_8125);
nand U8282 (N_8282,N_7781,N_7734);
nand U8283 (N_8283,N_8164,N_7997);
and U8284 (N_8284,N_7691,N_7753);
or U8285 (N_8285,N_7707,N_7553);
nor U8286 (N_8286,N_7970,N_8204);
and U8287 (N_8287,N_7683,N_7674);
or U8288 (N_8288,N_7763,N_7713);
or U8289 (N_8289,N_7612,N_7981);
nand U8290 (N_8290,N_7908,N_7675);
nand U8291 (N_8291,N_7541,N_7777);
or U8292 (N_8292,N_7767,N_8112);
nand U8293 (N_8293,N_7943,N_7559);
nor U8294 (N_8294,N_8139,N_8165);
nor U8295 (N_8295,N_7672,N_7939);
or U8296 (N_8296,N_7976,N_8213);
nor U8297 (N_8297,N_7967,N_8209);
nand U8298 (N_8298,N_7833,N_7568);
and U8299 (N_8299,N_8008,N_8233);
and U8300 (N_8300,N_7772,N_7537);
or U8301 (N_8301,N_7927,N_7622);
and U8302 (N_8302,N_8078,N_8195);
nor U8303 (N_8303,N_7842,N_7725);
nor U8304 (N_8304,N_8031,N_8045);
nor U8305 (N_8305,N_7792,N_8009);
nor U8306 (N_8306,N_8205,N_7996);
or U8307 (N_8307,N_7635,N_7745);
and U8308 (N_8308,N_7984,N_7933);
or U8309 (N_8309,N_7572,N_8055);
nor U8310 (N_8310,N_8021,N_8053);
and U8311 (N_8311,N_8101,N_7826);
nand U8312 (N_8312,N_8109,N_7949);
or U8313 (N_8313,N_7687,N_8066);
or U8314 (N_8314,N_7571,N_8236);
nand U8315 (N_8315,N_7705,N_8099);
nor U8316 (N_8316,N_8102,N_7910);
nor U8317 (N_8317,N_7565,N_7946);
nand U8318 (N_8318,N_8094,N_7944);
nand U8319 (N_8319,N_7850,N_8185);
nand U8320 (N_8320,N_7629,N_7542);
nand U8321 (N_8321,N_7564,N_8183);
nor U8322 (N_8322,N_7593,N_7504);
or U8323 (N_8323,N_8034,N_8010);
and U8324 (N_8324,N_8217,N_7723);
nor U8325 (N_8325,N_8075,N_7727);
and U8326 (N_8326,N_7744,N_7973);
or U8327 (N_8327,N_7776,N_7667);
or U8328 (N_8328,N_7861,N_7902);
or U8329 (N_8329,N_7836,N_7897);
nor U8330 (N_8330,N_7968,N_8087);
xnor U8331 (N_8331,N_7613,N_7872);
nand U8332 (N_8332,N_7748,N_7817);
nor U8333 (N_8333,N_7556,N_7978);
and U8334 (N_8334,N_7647,N_7808);
or U8335 (N_8335,N_7818,N_8141);
nand U8336 (N_8336,N_8081,N_8017);
or U8337 (N_8337,N_7567,N_7681);
nor U8338 (N_8338,N_7979,N_7554);
and U8339 (N_8339,N_7894,N_7584);
and U8340 (N_8340,N_8127,N_8171);
or U8341 (N_8341,N_7631,N_7765);
nand U8342 (N_8342,N_8147,N_7922);
nor U8343 (N_8343,N_7838,N_7769);
and U8344 (N_8344,N_7592,N_7615);
nor U8345 (N_8345,N_7728,N_7561);
nor U8346 (N_8346,N_7654,N_7869);
or U8347 (N_8347,N_7783,N_8214);
nor U8348 (N_8348,N_8098,N_7671);
or U8349 (N_8349,N_7889,N_7719);
and U8350 (N_8350,N_7982,N_7820);
nand U8351 (N_8351,N_8074,N_7914);
and U8352 (N_8352,N_7519,N_7873);
or U8353 (N_8353,N_7505,N_8058);
nor U8354 (N_8354,N_7513,N_7686);
nor U8355 (N_8355,N_7678,N_8135);
or U8356 (N_8356,N_8172,N_8239);
nor U8357 (N_8357,N_7766,N_7742);
nor U8358 (N_8358,N_8245,N_7576);
nor U8359 (N_8359,N_7806,N_8019);
or U8360 (N_8360,N_7954,N_8012);
and U8361 (N_8361,N_8007,N_7814);
nor U8362 (N_8362,N_8004,N_7676);
nor U8363 (N_8363,N_8206,N_7998);
nand U8364 (N_8364,N_7749,N_7652);
and U8365 (N_8365,N_7956,N_7757);
and U8366 (N_8366,N_7530,N_7884);
or U8367 (N_8367,N_8240,N_7768);
and U8368 (N_8368,N_8169,N_7986);
nand U8369 (N_8369,N_7579,N_7896);
nand U8370 (N_8370,N_7701,N_7682);
nand U8371 (N_8371,N_8192,N_7965);
and U8372 (N_8372,N_7828,N_8246);
and U8373 (N_8373,N_8064,N_7695);
or U8374 (N_8374,N_7555,N_7712);
nand U8375 (N_8375,N_7916,N_8089);
nand U8376 (N_8376,N_7692,N_8103);
nand U8377 (N_8377,N_8028,N_7771);
and U8378 (N_8378,N_8049,N_7547);
nand U8379 (N_8379,N_7616,N_7799);
or U8380 (N_8380,N_7878,N_8170);
nand U8381 (N_8381,N_8111,N_8175);
or U8382 (N_8382,N_7520,N_7557);
nor U8383 (N_8383,N_7560,N_7989);
nand U8384 (N_8384,N_7552,N_7661);
or U8385 (N_8385,N_7512,N_7536);
nand U8386 (N_8386,N_7854,N_8063);
or U8387 (N_8387,N_7901,N_7524);
nand U8388 (N_8388,N_7697,N_7926);
and U8389 (N_8389,N_7761,N_7843);
nor U8390 (N_8390,N_7760,N_7634);
nor U8391 (N_8391,N_8030,N_8156);
or U8392 (N_8392,N_7702,N_7639);
or U8393 (N_8393,N_7545,N_8090);
and U8394 (N_8394,N_7955,N_8145);
or U8395 (N_8395,N_7752,N_7837);
nor U8396 (N_8396,N_7740,N_7684);
xnor U8397 (N_8397,N_7971,N_8221);
nor U8398 (N_8398,N_8005,N_8208);
nand U8399 (N_8399,N_7726,N_7807);
xor U8400 (N_8400,N_7762,N_8050);
or U8401 (N_8401,N_7929,N_7583);
nand U8402 (N_8402,N_8243,N_8065);
or U8403 (N_8403,N_7642,N_7506);
and U8404 (N_8404,N_8151,N_7656);
nand U8405 (N_8405,N_8091,N_7832);
or U8406 (N_8406,N_7739,N_8067);
nand U8407 (N_8407,N_8248,N_8013);
or U8408 (N_8408,N_7821,N_7633);
or U8409 (N_8409,N_7881,N_8223);
nor U8410 (N_8410,N_8129,N_7688);
nand U8411 (N_8411,N_7600,N_7599);
nor U8412 (N_8412,N_7580,N_8181);
or U8413 (N_8413,N_8136,N_7509);
and U8414 (N_8414,N_7801,N_8222);
or U8415 (N_8415,N_7680,N_8059);
and U8416 (N_8416,N_7856,N_7879);
and U8417 (N_8417,N_7871,N_8130);
or U8418 (N_8418,N_8144,N_7636);
xor U8419 (N_8419,N_7577,N_8216);
nand U8420 (N_8420,N_7947,N_8054);
xor U8421 (N_8421,N_7747,N_7632);
nor U8422 (N_8422,N_7549,N_7698);
or U8423 (N_8423,N_7511,N_7827);
or U8424 (N_8424,N_8249,N_8202);
nor U8425 (N_8425,N_8092,N_7644);
nand U8426 (N_8426,N_7890,N_7866);
nand U8427 (N_8427,N_7846,N_8158);
nand U8428 (N_8428,N_7528,N_8132);
or U8429 (N_8429,N_7816,N_8197);
nand U8430 (N_8430,N_7885,N_8095);
nor U8431 (N_8431,N_7983,N_7849);
or U8432 (N_8432,N_7962,N_8231);
nand U8433 (N_8433,N_8235,N_7673);
and U8434 (N_8434,N_8122,N_8133);
nand U8435 (N_8435,N_7533,N_7704);
or U8436 (N_8436,N_7733,N_7658);
and U8437 (N_8437,N_8033,N_7508);
nand U8438 (N_8438,N_7711,N_7538);
or U8439 (N_8439,N_8201,N_8186);
nand U8440 (N_8440,N_7751,N_8179);
nand U8441 (N_8441,N_8052,N_8166);
nand U8442 (N_8442,N_7925,N_8163);
nand U8443 (N_8443,N_7840,N_7911);
nand U8444 (N_8444,N_7857,N_7502);
nor U8445 (N_8445,N_7529,N_7764);
nor U8446 (N_8446,N_7811,N_8203);
and U8447 (N_8447,N_7917,N_8211);
nor U8448 (N_8448,N_7887,N_7581);
nand U8449 (N_8449,N_8027,N_7638);
and U8450 (N_8450,N_7664,N_8219);
nor U8451 (N_8451,N_7607,N_7746);
nand U8452 (N_8452,N_7852,N_7665);
nand U8453 (N_8453,N_7755,N_7570);
or U8454 (N_8454,N_7663,N_7810);
and U8455 (N_8455,N_8198,N_7620);
nor U8456 (N_8456,N_7985,N_8006);
nand U8457 (N_8457,N_7829,N_8057);
nor U8458 (N_8458,N_7619,N_7907);
or U8459 (N_8459,N_7500,N_7831);
nor U8460 (N_8460,N_7793,N_8086);
nor U8461 (N_8461,N_7640,N_7608);
and U8462 (N_8462,N_7913,N_7578);
or U8463 (N_8463,N_7899,N_8153);
and U8464 (N_8464,N_8237,N_8016);
nor U8465 (N_8465,N_7657,N_7812);
nor U8466 (N_8466,N_8184,N_7703);
nor U8467 (N_8467,N_7796,N_8174);
nand U8468 (N_8468,N_7527,N_8154);
and U8469 (N_8469,N_8046,N_7980);
and U8470 (N_8470,N_7912,N_7794);
or U8471 (N_8471,N_7550,N_7779);
xor U8472 (N_8472,N_7964,N_8193);
nor U8473 (N_8473,N_7845,N_8143);
xnor U8474 (N_8474,N_8196,N_8134);
and U8475 (N_8475,N_8070,N_7525);
nor U8476 (N_8476,N_8088,N_7741);
nor U8477 (N_8477,N_8026,N_7625);
nor U8478 (N_8478,N_7867,N_7848);
and U8479 (N_8479,N_7778,N_8068);
nor U8480 (N_8480,N_7532,N_7839);
or U8481 (N_8481,N_8085,N_7699);
or U8482 (N_8482,N_8138,N_8061);
nor U8483 (N_8483,N_7940,N_7780);
and U8484 (N_8484,N_7718,N_7855);
and U8485 (N_8485,N_7659,N_7834);
or U8486 (N_8486,N_8152,N_8039);
nor U8487 (N_8487,N_7611,N_7809);
and U8488 (N_8488,N_7602,N_7789);
nor U8489 (N_8489,N_8121,N_7637);
nor U8490 (N_8490,N_7905,N_8150);
or U8491 (N_8491,N_7666,N_7655);
nor U8492 (N_8492,N_8001,N_7750);
xor U8493 (N_8493,N_8029,N_7900);
and U8494 (N_8494,N_7591,N_7724);
and U8495 (N_8495,N_8080,N_7660);
nor U8496 (N_8496,N_7618,N_7870);
and U8497 (N_8497,N_8038,N_7715);
or U8498 (N_8498,N_7626,N_7931);
nand U8499 (N_8499,N_7961,N_8189);
nor U8500 (N_8500,N_7880,N_7918);
xnor U8501 (N_8501,N_8215,N_7966);
xor U8502 (N_8502,N_7875,N_7957);
xor U8503 (N_8503,N_7924,N_7886);
and U8504 (N_8504,N_7994,N_7883);
or U8505 (N_8505,N_7526,N_7604);
and U8506 (N_8506,N_8100,N_8238);
nor U8507 (N_8507,N_7919,N_7898);
or U8508 (N_8508,N_8118,N_7932);
nand U8509 (N_8509,N_7790,N_8104);
and U8510 (N_8510,N_7819,N_8220);
nor U8511 (N_8511,N_7784,N_7795);
or U8512 (N_8512,N_8242,N_8218);
nand U8513 (N_8513,N_8234,N_7507);
xor U8514 (N_8514,N_8037,N_7668);
and U8515 (N_8515,N_7906,N_7860);
xor U8516 (N_8516,N_8043,N_7975);
nor U8517 (N_8517,N_7706,N_7546);
and U8518 (N_8518,N_8071,N_7516);
and U8519 (N_8519,N_8140,N_7669);
or U8520 (N_8520,N_7582,N_8022);
nand U8521 (N_8521,N_7648,N_7877);
nand U8522 (N_8522,N_7830,N_7773);
xnor U8523 (N_8523,N_7685,N_7543);
nor U8524 (N_8524,N_7876,N_8041);
nand U8525 (N_8525,N_7627,N_7595);
nor U8526 (N_8526,N_8230,N_7514);
and U8527 (N_8527,N_7847,N_8002);
or U8528 (N_8528,N_7510,N_7938);
xnor U8529 (N_8529,N_8079,N_7859);
nand U8530 (N_8530,N_8182,N_7523);
nand U8531 (N_8531,N_7920,N_8212);
and U8532 (N_8532,N_7803,N_8168);
nor U8533 (N_8533,N_8159,N_8110);
nor U8534 (N_8534,N_8096,N_8117);
nand U8535 (N_8535,N_8015,N_7714);
or U8536 (N_8536,N_7521,N_8228);
nor U8537 (N_8537,N_7921,N_8225);
or U8538 (N_8538,N_8020,N_8126);
nand U8539 (N_8539,N_8115,N_8083);
nor U8540 (N_8540,N_7522,N_8062);
nand U8541 (N_8541,N_7909,N_7531);
and U8542 (N_8542,N_7597,N_7841);
nand U8543 (N_8543,N_8149,N_8229);
xnor U8544 (N_8544,N_7775,N_7700);
nor U8545 (N_8545,N_8116,N_8036);
and U8546 (N_8546,N_8244,N_7758);
and U8547 (N_8547,N_8167,N_7952);
xnor U8548 (N_8548,N_7735,N_7670);
xor U8549 (N_8549,N_8069,N_7729);
and U8550 (N_8550,N_7732,N_8157);
and U8551 (N_8551,N_7515,N_7650);
and U8552 (N_8552,N_7563,N_8173);
or U8553 (N_8553,N_7936,N_7596);
or U8554 (N_8554,N_7679,N_7645);
nand U8555 (N_8555,N_7590,N_7786);
xor U8556 (N_8556,N_7517,N_7736);
and U8557 (N_8557,N_8023,N_7694);
and U8558 (N_8558,N_7610,N_7689);
nor U8559 (N_8559,N_7853,N_7945);
nor U8560 (N_8560,N_8077,N_7972);
nor U8561 (N_8561,N_8024,N_7937);
and U8562 (N_8562,N_7649,N_7544);
nor U8563 (N_8563,N_7823,N_8105);
or U8564 (N_8564,N_7835,N_7548);
or U8565 (N_8565,N_7603,N_8108);
nand U8566 (N_8566,N_7798,N_8161);
nor U8567 (N_8567,N_7774,N_8014);
xor U8568 (N_8568,N_8051,N_8097);
nand U8569 (N_8569,N_7858,N_7662);
and U8570 (N_8570,N_7540,N_7643);
nor U8571 (N_8571,N_7851,N_7863);
nor U8572 (N_8572,N_8119,N_7791);
nand U8573 (N_8573,N_7958,N_8155);
nor U8574 (N_8574,N_7731,N_7951);
or U8575 (N_8575,N_8093,N_8040);
or U8576 (N_8576,N_7641,N_7677);
or U8577 (N_8577,N_8176,N_7800);
nor U8578 (N_8578,N_7991,N_7503);
or U8579 (N_8579,N_7891,N_7948);
or U8580 (N_8580,N_7759,N_7606);
and U8581 (N_8581,N_7696,N_7534);
nor U8582 (N_8582,N_7501,N_7915);
nor U8583 (N_8583,N_7621,N_7999);
and U8584 (N_8584,N_7605,N_7797);
or U8585 (N_8585,N_7990,N_8148);
or U8586 (N_8586,N_8025,N_7865);
or U8587 (N_8587,N_8199,N_7882);
nand U8588 (N_8588,N_8082,N_7587);
nor U8589 (N_8589,N_7804,N_7815);
or U8590 (N_8590,N_8200,N_7589);
and U8591 (N_8591,N_7574,N_7722);
or U8592 (N_8592,N_7558,N_7825);
nand U8593 (N_8593,N_7738,N_7623);
nor U8594 (N_8594,N_7824,N_8123);
or U8595 (N_8595,N_7988,N_8187);
nor U8596 (N_8596,N_8114,N_8106);
and U8597 (N_8597,N_7569,N_7788);
nor U8598 (N_8598,N_7888,N_7977);
nor U8599 (N_8599,N_8120,N_8047);
and U8600 (N_8600,N_7844,N_7802);
nor U8601 (N_8601,N_7923,N_7959);
or U8602 (N_8602,N_7539,N_7720);
nand U8603 (N_8603,N_7624,N_7995);
and U8604 (N_8604,N_7892,N_7690);
nand U8605 (N_8605,N_8210,N_7960);
nor U8606 (N_8606,N_7716,N_8207);
or U8607 (N_8607,N_7730,N_7950);
nand U8608 (N_8608,N_8137,N_8188);
nor U8609 (N_8609,N_8232,N_7585);
nand U8610 (N_8610,N_7756,N_7551);
nand U8611 (N_8611,N_7575,N_7770);
nand U8612 (N_8612,N_8000,N_7693);
nand U8613 (N_8613,N_7864,N_7969);
and U8614 (N_8614,N_7710,N_7588);
nor U8615 (N_8615,N_8247,N_7963);
and U8616 (N_8616,N_7651,N_8042);
and U8617 (N_8617,N_7822,N_7928);
or U8618 (N_8618,N_7721,N_8035);
and U8619 (N_8619,N_7518,N_7566);
or U8620 (N_8620,N_7586,N_7573);
nand U8621 (N_8621,N_8124,N_8241);
or U8622 (N_8622,N_7598,N_7594);
or U8623 (N_8623,N_8084,N_8060);
nand U8624 (N_8624,N_7934,N_7895);
nor U8625 (N_8625,N_7656,N_8086);
nor U8626 (N_8626,N_8020,N_7841);
xor U8627 (N_8627,N_8167,N_7694);
and U8628 (N_8628,N_7619,N_8209);
nand U8629 (N_8629,N_8064,N_7705);
nor U8630 (N_8630,N_7530,N_8030);
or U8631 (N_8631,N_7911,N_8178);
nor U8632 (N_8632,N_7750,N_8133);
nand U8633 (N_8633,N_7889,N_7581);
or U8634 (N_8634,N_7880,N_8191);
and U8635 (N_8635,N_7527,N_7962);
nand U8636 (N_8636,N_8225,N_7923);
and U8637 (N_8637,N_7805,N_8028);
nor U8638 (N_8638,N_7616,N_7853);
or U8639 (N_8639,N_8153,N_8190);
nand U8640 (N_8640,N_8005,N_7516);
and U8641 (N_8641,N_7604,N_8188);
and U8642 (N_8642,N_8041,N_8062);
or U8643 (N_8643,N_8086,N_8102);
and U8644 (N_8644,N_7845,N_8135);
or U8645 (N_8645,N_7798,N_7692);
and U8646 (N_8646,N_8071,N_7690);
or U8647 (N_8647,N_7943,N_7795);
nand U8648 (N_8648,N_8004,N_8237);
or U8649 (N_8649,N_8129,N_7994);
or U8650 (N_8650,N_8029,N_7688);
nand U8651 (N_8651,N_7619,N_7661);
xor U8652 (N_8652,N_7661,N_8236);
or U8653 (N_8653,N_8229,N_8041);
nand U8654 (N_8654,N_8066,N_7794);
and U8655 (N_8655,N_7836,N_8029);
and U8656 (N_8656,N_7755,N_7978);
and U8657 (N_8657,N_7723,N_7602);
nor U8658 (N_8658,N_7916,N_7521);
and U8659 (N_8659,N_7993,N_7577);
or U8660 (N_8660,N_7552,N_8119);
and U8661 (N_8661,N_7540,N_8227);
and U8662 (N_8662,N_7653,N_8198);
nand U8663 (N_8663,N_7640,N_8106);
nor U8664 (N_8664,N_8031,N_7711);
and U8665 (N_8665,N_7743,N_7715);
nand U8666 (N_8666,N_8198,N_7619);
nand U8667 (N_8667,N_7512,N_7583);
and U8668 (N_8668,N_7598,N_7922);
and U8669 (N_8669,N_7696,N_8054);
nand U8670 (N_8670,N_8232,N_7882);
nor U8671 (N_8671,N_7719,N_8006);
or U8672 (N_8672,N_8066,N_8234);
and U8673 (N_8673,N_7748,N_7592);
or U8674 (N_8674,N_8023,N_7510);
nor U8675 (N_8675,N_7571,N_7500);
or U8676 (N_8676,N_7849,N_8144);
nor U8677 (N_8677,N_7807,N_7745);
or U8678 (N_8678,N_8071,N_7756);
nand U8679 (N_8679,N_7711,N_8192);
and U8680 (N_8680,N_8207,N_7799);
and U8681 (N_8681,N_7729,N_7537);
nand U8682 (N_8682,N_8120,N_8217);
and U8683 (N_8683,N_7567,N_8139);
nand U8684 (N_8684,N_7816,N_7514);
nand U8685 (N_8685,N_8138,N_8022);
and U8686 (N_8686,N_8049,N_7962);
nand U8687 (N_8687,N_7918,N_7964);
nor U8688 (N_8688,N_7787,N_7685);
and U8689 (N_8689,N_7905,N_7833);
or U8690 (N_8690,N_7919,N_7680);
and U8691 (N_8691,N_8076,N_8235);
and U8692 (N_8692,N_7516,N_7633);
and U8693 (N_8693,N_7957,N_8089);
nor U8694 (N_8694,N_7960,N_7771);
nor U8695 (N_8695,N_8232,N_8034);
nor U8696 (N_8696,N_7520,N_7894);
and U8697 (N_8697,N_8058,N_7590);
or U8698 (N_8698,N_7518,N_7805);
nand U8699 (N_8699,N_8204,N_8145);
nor U8700 (N_8700,N_8155,N_7947);
nor U8701 (N_8701,N_8242,N_7633);
or U8702 (N_8702,N_7695,N_7891);
or U8703 (N_8703,N_7697,N_7593);
and U8704 (N_8704,N_7741,N_7955);
nor U8705 (N_8705,N_8042,N_7876);
nand U8706 (N_8706,N_7942,N_7566);
nor U8707 (N_8707,N_8043,N_8119);
or U8708 (N_8708,N_7864,N_8083);
xnor U8709 (N_8709,N_7832,N_7691);
and U8710 (N_8710,N_7531,N_8010);
nand U8711 (N_8711,N_7527,N_8029);
and U8712 (N_8712,N_8016,N_8114);
or U8713 (N_8713,N_7920,N_8141);
or U8714 (N_8714,N_7806,N_7812);
nor U8715 (N_8715,N_8097,N_7730);
nor U8716 (N_8716,N_7785,N_8006);
nand U8717 (N_8717,N_8023,N_7538);
or U8718 (N_8718,N_7902,N_7788);
and U8719 (N_8719,N_8242,N_7747);
nand U8720 (N_8720,N_8174,N_8189);
and U8721 (N_8721,N_7729,N_7705);
nor U8722 (N_8722,N_8236,N_8133);
and U8723 (N_8723,N_7636,N_8074);
nand U8724 (N_8724,N_8102,N_7985);
or U8725 (N_8725,N_7660,N_8006);
and U8726 (N_8726,N_8067,N_7596);
nand U8727 (N_8727,N_7578,N_7561);
nor U8728 (N_8728,N_7982,N_7931);
nor U8729 (N_8729,N_7865,N_7759);
nor U8730 (N_8730,N_7632,N_8006);
and U8731 (N_8731,N_8185,N_7549);
and U8732 (N_8732,N_7691,N_7975);
and U8733 (N_8733,N_8100,N_7521);
nor U8734 (N_8734,N_7968,N_8134);
nor U8735 (N_8735,N_7846,N_7672);
and U8736 (N_8736,N_7873,N_7566);
nor U8737 (N_8737,N_7688,N_7531);
nand U8738 (N_8738,N_8001,N_7790);
and U8739 (N_8739,N_7893,N_7524);
and U8740 (N_8740,N_8119,N_8171);
and U8741 (N_8741,N_8006,N_7695);
and U8742 (N_8742,N_7607,N_7771);
or U8743 (N_8743,N_7967,N_7954);
or U8744 (N_8744,N_7977,N_7617);
or U8745 (N_8745,N_7722,N_8125);
nand U8746 (N_8746,N_7721,N_8163);
nor U8747 (N_8747,N_7870,N_7800);
or U8748 (N_8748,N_7531,N_7597);
or U8749 (N_8749,N_7614,N_8099);
or U8750 (N_8750,N_8159,N_7561);
and U8751 (N_8751,N_7740,N_8101);
or U8752 (N_8752,N_7901,N_7905);
and U8753 (N_8753,N_7929,N_7768);
nand U8754 (N_8754,N_7750,N_7833);
nor U8755 (N_8755,N_8200,N_7889);
nand U8756 (N_8756,N_7572,N_7509);
nor U8757 (N_8757,N_8097,N_7884);
or U8758 (N_8758,N_8132,N_7697);
and U8759 (N_8759,N_8096,N_7718);
and U8760 (N_8760,N_8091,N_7998);
nand U8761 (N_8761,N_7931,N_7780);
nand U8762 (N_8762,N_7786,N_7950);
or U8763 (N_8763,N_7970,N_8199);
or U8764 (N_8764,N_8153,N_8087);
or U8765 (N_8765,N_7753,N_8034);
nand U8766 (N_8766,N_7860,N_7723);
nand U8767 (N_8767,N_7794,N_8186);
or U8768 (N_8768,N_8157,N_7571);
nand U8769 (N_8769,N_7728,N_8206);
nand U8770 (N_8770,N_7869,N_7501);
or U8771 (N_8771,N_8126,N_7987);
xor U8772 (N_8772,N_7817,N_7903);
or U8773 (N_8773,N_8030,N_7776);
nand U8774 (N_8774,N_7941,N_7949);
or U8775 (N_8775,N_7939,N_7606);
nor U8776 (N_8776,N_7569,N_7951);
and U8777 (N_8777,N_7997,N_8197);
or U8778 (N_8778,N_7637,N_8069);
and U8779 (N_8779,N_8229,N_7606);
and U8780 (N_8780,N_7807,N_8010);
or U8781 (N_8781,N_7945,N_7919);
nor U8782 (N_8782,N_7967,N_7972);
and U8783 (N_8783,N_7650,N_8087);
and U8784 (N_8784,N_8101,N_7952);
nor U8785 (N_8785,N_7563,N_8233);
nor U8786 (N_8786,N_7657,N_7703);
and U8787 (N_8787,N_8108,N_8192);
nor U8788 (N_8788,N_7617,N_8142);
or U8789 (N_8789,N_7993,N_8053);
or U8790 (N_8790,N_7718,N_8065);
nand U8791 (N_8791,N_7746,N_7712);
nor U8792 (N_8792,N_8078,N_7934);
or U8793 (N_8793,N_8107,N_7799);
or U8794 (N_8794,N_8024,N_8017);
or U8795 (N_8795,N_7817,N_7845);
and U8796 (N_8796,N_7525,N_7686);
nor U8797 (N_8797,N_7963,N_7634);
or U8798 (N_8798,N_7580,N_7783);
or U8799 (N_8799,N_8239,N_8099);
nand U8800 (N_8800,N_8033,N_7591);
and U8801 (N_8801,N_8085,N_7778);
and U8802 (N_8802,N_7747,N_8243);
nor U8803 (N_8803,N_8034,N_7945);
nor U8804 (N_8804,N_7884,N_7866);
nand U8805 (N_8805,N_7917,N_7548);
and U8806 (N_8806,N_7793,N_7921);
and U8807 (N_8807,N_7817,N_7616);
nand U8808 (N_8808,N_7678,N_7941);
and U8809 (N_8809,N_8103,N_8080);
or U8810 (N_8810,N_7576,N_7698);
nor U8811 (N_8811,N_8020,N_7617);
and U8812 (N_8812,N_8239,N_7509);
nor U8813 (N_8813,N_7706,N_7865);
or U8814 (N_8814,N_8228,N_7819);
or U8815 (N_8815,N_7767,N_7582);
or U8816 (N_8816,N_8016,N_7677);
xor U8817 (N_8817,N_7731,N_8038);
or U8818 (N_8818,N_8089,N_7946);
nand U8819 (N_8819,N_8030,N_8103);
nand U8820 (N_8820,N_7666,N_7928);
and U8821 (N_8821,N_8065,N_7548);
and U8822 (N_8822,N_7625,N_7913);
nand U8823 (N_8823,N_7860,N_8011);
xor U8824 (N_8824,N_7907,N_7608);
nor U8825 (N_8825,N_7951,N_7640);
and U8826 (N_8826,N_7722,N_7706);
nand U8827 (N_8827,N_7742,N_7750);
or U8828 (N_8828,N_7968,N_7625);
and U8829 (N_8829,N_7949,N_8102);
and U8830 (N_8830,N_8145,N_8139);
or U8831 (N_8831,N_7731,N_7773);
nor U8832 (N_8832,N_8147,N_8102);
and U8833 (N_8833,N_8177,N_7866);
or U8834 (N_8834,N_7790,N_7701);
or U8835 (N_8835,N_7811,N_8245);
and U8836 (N_8836,N_7914,N_8041);
or U8837 (N_8837,N_8236,N_8009);
nor U8838 (N_8838,N_7867,N_7523);
nand U8839 (N_8839,N_8095,N_8012);
or U8840 (N_8840,N_7508,N_8198);
nor U8841 (N_8841,N_8133,N_7685);
or U8842 (N_8842,N_8091,N_7646);
nor U8843 (N_8843,N_8172,N_8236);
or U8844 (N_8844,N_7943,N_7987);
xor U8845 (N_8845,N_7877,N_8167);
and U8846 (N_8846,N_7886,N_7738);
or U8847 (N_8847,N_7677,N_8203);
or U8848 (N_8848,N_7831,N_7828);
nand U8849 (N_8849,N_8175,N_7778);
and U8850 (N_8850,N_8082,N_8191);
nand U8851 (N_8851,N_7853,N_7526);
and U8852 (N_8852,N_7620,N_7972);
or U8853 (N_8853,N_7870,N_7822);
and U8854 (N_8854,N_7638,N_8054);
and U8855 (N_8855,N_7994,N_7692);
nand U8856 (N_8856,N_7514,N_7815);
nand U8857 (N_8857,N_7595,N_8155);
nor U8858 (N_8858,N_7995,N_8127);
and U8859 (N_8859,N_7537,N_7946);
or U8860 (N_8860,N_7612,N_7795);
nor U8861 (N_8861,N_7959,N_7843);
nand U8862 (N_8862,N_7647,N_8202);
nor U8863 (N_8863,N_7523,N_7693);
and U8864 (N_8864,N_8116,N_7537);
nand U8865 (N_8865,N_7845,N_7579);
and U8866 (N_8866,N_7938,N_8189);
and U8867 (N_8867,N_7830,N_8173);
nor U8868 (N_8868,N_7888,N_7752);
nand U8869 (N_8869,N_7768,N_8157);
nor U8870 (N_8870,N_7779,N_7690);
or U8871 (N_8871,N_7953,N_8047);
or U8872 (N_8872,N_8141,N_7810);
and U8873 (N_8873,N_7601,N_7643);
nor U8874 (N_8874,N_7522,N_8176);
or U8875 (N_8875,N_7942,N_7537);
or U8876 (N_8876,N_7586,N_7717);
or U8877 (N_8877,N_7692,N_7929);
xor U8878 (N_8878,N_8204,N_8128);
and U8879 (N_8879,N_8213,N_7533);
nor U8880 (N_8880,N_7524,N_8093);
and U8881 (N_8881,N_7685,N_7713);
nand U8882 (N_8882,N_7515,N_7689);
or U8883 (N_8883,N_7940,N_7767);
and U8884 (N_8884,N_7600,N_8085);
nand U8885 (N_8885,N_8009,N_8220);
nand U8886 (N_8886,N_8020,N_7713);
or U8887 (N_8887,N_7695,N_8198);
or U8888 (N_8888,N_7725,N_7779);
nand U8889 (N_8889,N_7719,N_7636);
or U8890 (N_8890,N_7913,N_7869);
and U8891 (N_8891,N_7637,N_8080);
nand U8892 (N_8892,N_7530,N_8241);
nand U8893 (N_8893,N_7792,N_7868);
nor U8894 (N_8894,N_8161,N_7522);
nor U8895 (N_8895,N_7835,N_7503);
nand U8896 (N_8896,N_7770,N_7587);
and U8897 (N_8897,N_8144,N_7615);
xor U8898 (N_8898,N_8237,N_8188);
or U8899 (N_8899,N_7948,N_7860);
and U8900 (N_8900,N_7688,N_8131);
or U8901 (N_8901,N_8075,N_7602);
nand U8902 (N_8902,N_8040,N_8190);
nor U8903 (N_8903,N_8160,N_7550);
nor U8904 (N_8904,N_8029,N_7675);
nand U8905 (N_8905,N_8135,N_7709);
nand U8906 (N_8906,N_7770,N_8249);
or U8907 (N_8907,N_8000,N_7919);
nand U8908 (N_8908,N_7830,N_7607);
nor U8909 (N_8909,N_8039,N_8173);
and U8910 (N_8910,N_7763,N_7975);
and U8911 (N_8911,N_7755,N_8083);
nand U8912 (N_8912,N_7867,N_7701);
nor U8913 (N_8913,N_7554,N_7526);
and U8914 (N_8914,N_7950,N_7981);
nor U8915 (N_8915,N_7833,N_7910);
and U8916 (N_8916,N_7804,N_7930);
xor U8917 (N_8917,N_8208,N_8158);
and U8918 (N_8918,N_7506,N_7725);
and U8919 (N_8919,N_7783,N_7651);
nand U8920 (N_8920,N_7831,N_7634);
or U8921 (N_8921,N_8035,N_7837);
nand U8922 (N_8922,N_7631,N_8192);
and U8923 (N_8923,N_7840,N_7999);
and U8924 (N_8924,N_7712,N_7718);
and U8925 (N_8925,N_7646,N_7791);
or U8926 (N_8926,N_7981,N_7899);
and U8927 (N_8927,N_8224,N_8110);
or U8928 (N_8928,N_7511,N_7906);
and U8929 (N_8929,N_8099,N_8148);
or U8930 (N_8930,N_7999,N_7945);
and U8931 (N_8931,N_7986,N_7625);
nor U8932 (N_8932,N_8017,N_7708);
nor U8933 (N_8933,N_7980,N_8187);
and U8934 (N_8934,N_7713,N_7717);
nor U8935 (N_8935,N_7736,N_8174);
nor U8936 (N_8936,N_7871,N_7800);
nand U8937 (N_8937,N_8199,N_7529);
or U8938 (N_8938,N_7513,N_7667);
nor U8939 (N_8939,N_8173,N_7851);
and U8940 (N_8940,N_7994,N_7632);
nand U8941 (N_8941,N_7813,N_7897);
and U8942 (N_8942,N_7658,N_7889);
nor U8943 (N_8943,N_7619,N_8244);
or U8944 (N_8944,N_7893,N_8156);
or U8945 (N_8945,N_8218,N_8143);
or U8946 (N_8946,N_7747,N_7771);
and U8947 (N_8947,N_7920,N_8103);
and U8948 (N_8948,N_7726,N_7973);
and U8949 (N_8949,N_7885,N_7706);
nor U8950 (N_8950,N_7867,N_7719);
nor U8951 (N_8951,N_7540,N_8107);
nand U8952 (N_8952,N_7910,N_7709);
or U8953 (N_8953,N_7775,N_7926);
and U8954 (N_8954,N_7839,N_8225);
and U8955 (N_8955,N_8085,N_7634);
nor U8956 (N_8956,N_7657,N_8110);
nand U8957 (N_8957,N_7888,N_7518);
or U8958 (N_8958,N_7755,N_7731);
nor U8959 (N_8959,N_8197,N_8140);
or U8960 (N_8960,N_8183,N_7520);
nand U8961 (N_8961,N_8239,N_7980);
and U8962 (N_8962,N_7648,N_7533);
and U8963 (N_8963,N_7569,N_7916);
or U8964 (N_8964,N_8145,N_7720);
or U8965 (N_8965,N_8009,N_8178);
xnor U8966 (N_8966,N_8091,N_7986);
xnor U8967 (N_8967,N_7989,N_7659);
and U8968 (N_8968,N_8140,N_7866);
xnor U8969 (N_8969,N_7812,N_7908);
and U8970 (N_8970,N_7892,N_7750);
nand U8971 (N_8971,N_8095,N_7891);
or U8972 (N_8972,N_8142,N_8170);
or U8973 (N_8973,N_7569,N_7961);
nand U8974 (N_8974,N_7604,N_7993);
and U8975 (N_8975,N_8058,N_7732);
nand U8976 (N_8976,N_7900,N_7993);
or U8977 (N_8977,N_7942,N_8120);
and U8978 (N_8978,N_7757,N_8067);
and U8979 (N_8979,N_7563,N_7784);
nand U8980 (N_8980,N_8216,N_7785);
nor U8981 (N_8981,N_8226,N_7613);
or U8982 (N_8982,N_8170,N_7940);
nand U8983 (N_8983,N_7838,N_7827);
or U8984 (N_8984,N_7773,N_7535);
nor U8985 (N_8985,N_8184,N_8197);
nand U8986 (N_8986,N_7837,N_7911);
nor U8987 (N_8987,N_8143,N_8221);
or U8988 (N_8988,N_7782,N_8068);
nand U8989 (N_8989,N_8142,N_7544);
and U8990 (N_8990,N_7984,N_7803);
nor U8991 (N_8991,N_8099,N_8206);
and U8992 (N_8992,N_7554,N_7778);
and U8993 (N_8993,N_8216,N_7516);
or U8994 (N_8994,N_7627,N_7931);
or U8995 (N_8995,N_7881,N_8248);
nand U8996 (N_8996,N_7987,N_7846);
nor U8997 (N_8997,N_7851,N_7822);
and U8998 (N_8998,N_8145,N_8063);
and U8999 (N_8999,N_7750,N_7845);
and U9000 (N_9000,N_8694,N_8554);
and U9001 (N_9001,N_8276,N_8675);
and U9002 (N_9002,N_8522,N_8772);
and U9003 (N_9003,N_8760,N_8671);
or U9004 (N_9004,N_8487,N_8714);
nand U9005 (N_9005,N_8673,N_8441);
and U9006 (N_9006,N_8503,N_8439);
nor U9007 (N_9007,N_8743,N_8941);
or U9008 (N_9008,N_8952,N_8570);
nor U9009 (N_9009,N_8582,N_8739);
and U9010 (N_9010,N_8676,N_8600);
nand U9011 (N_9011,N_8786,N_8966);
nand U9012 (N_9012,N_8907,N_8720);
nand U9013 (N_9013,N_8428,N_8851);
nand U9014 (N_9014,N_8316,N_8767);
nor U9015 (N_9015,N_8867,N_8454);
and U9016 (N_9016,N_8303,N_8823);
nand U9017 (N_9017,N_8475,N_8365);
nand U9018 (N_9018,N_8822,N_8814);
or U9019 (N_9019,N_8889,N_8343);
and U9020 (N_9020,N_8610,N_8806);
and U9021 (N_9021,N_8840,N_8313);
nand U9022 (N_9022,N_8271,N_8918);
and U9023 (N_9023,N_8565,N_8401);
or U9024 (N_9024,N_8638,N_8521);
nand U9025 (N_9025,N_8652,N_8419);
nor U9026 (N_9026,N_8555,N_8415);
nor U9027 (N_9027,N_8285,N_8452);
nor U9028 (N_9028,N_8580,N_8967);
and U9029 (N_9029,N_8597,N_8985);
or U9030 (N_9030,N_8341,N_8818);
and U9031 (N_9031,N_8911,N_8334);
nand U9032 (N_9032,N_8378,N_8848);
and U9033 (N_9033,N_8844,N_8647);
nor U9034 (N_9034,N_8479,N_8721);
nor U9035 (N_9035,N_8980,N_8595);
and U9036 (N_9036,N_8498,N_8540);
and U9037 (N_9037,N_8813,N_8387);
nand U9038 (N_9038,N_8315,N_8490);
or U9039 (N_9039,N_8320,N_8651);
or U9040 (N_9040,N_8512,N_8527);
nand U9041 (N_9041,N_8278,N_8863);
nand U9042 (N_9042,N_8447,N_8735);
nand U9043 (N_9043,N_8456,N_8978);
or U9044 (N_9044,N_8639,N_8546);
nand U9045 (N_9045,N_8411,N_8658);
nor U9046 (N_9046,N_8504,N_8348);
and U9047 (N_9047,N_8389,N_8587);
or U9048 (N_9048,N_8367,N_8645);
and U9049 (N_9049,N_8843,N_8596);
nor U9050 (N_9050,N_8817,N_8766);
nand U9051 (N_9051,N_8446,N_8514);
nand U9052 (N_9052,N_8869,N_8269);
nor U9053 (N_9053,N_8841,N_8536);
nand U9054 (N_9054,N_8853,N_8268);
nand U9055 (N_9055,N_8513,N_8396);
or U9056 (N_9056,N_8820,N_8888);
nand U9057 (N_9057,N_8252,N_8350);
nand U9058 (N_9058,N_8682,N_8520);
and U9059 (N_9059,N_8277,N_8931);
nand U9060 (N_9060,N_8940,N_8871);
and U9061 (N_9061,N_8724,N_8697);
and U9062 (N_9062,N_8287,N_8924);
or U9063 (N_9063,N_8986,N_8497);
or U9064 (N_9064,N_8898,N_8335);
and U9065 (N_9065,N_8619,N_8649);
nand U9066 (N_9066,N_8391,N_8874);
or U9067 (N_9067,N_8685,N_8865);
or U9068 (N_9068,N_8643,N_8768);
or U9069 (N_9069,N_8662,N_8559);
and U9070 (N_9070,N_8346,N_8255);
nor U9071 (N_9071,N_8880,N_8704);
or U9072 (N_9072,N_8613,N_8405);
or U9073 (N_9073,N_8775,N_8502);
or U9074 (N_9074,N_8796,N_8905);
xor U9075 (N_9075,N_8581,N_8795);
nor U9076 (N_9076,N_8618,N_8584);
or U9077 (N_9077,N_8265,N_8374);
and U9078 (N_9078,N_8921,N_8407);
xor U9079 (N_9079,N_8749,N_8716);
xnor U9080 (N_9080,N_8801,N_8432);
nor U9081 (N_9081,N_8585,N_8528);
or U9082 (N_9082,N_8493,N_8460);
nand U9083 (N_9083,N_8553,N_8511);
nand U9084 (N_9084,N_8572,N_8525);
nor U9085 (N_9085,N_8362,N_8802);
or U9086 (N_9086,N_8949,N_8532);
nor U9087 (N_9087,N_8489,N_8327);
or U9088 (N_9088,N_8609,N_8642);
nor U9089 (N_9089,N_8438,N_8423);
or U9090 (N_9090,N_8925,N_8726);
nor U9091 (N_9091,N_8859,N_8894);
nor U9092 (N_9092,N_8624,N_8462);
nor U9093 (N_9093,N_8424,N_8304);
or U9094 (N_9094,N_8725,N_8288);
nand U9095 (N_9095,N_8355,N_8598);
nor U9096 (N_9096,N_8295,N_8845);
and U9097 (N_9097,N_8302,N_8661);
and U9098 (N_9098,N_8495,N_8975);
or U9099 (N_9099,N_8633,N_8830);
nor U9100 (N_9100,N_8686,N_8896);
or U9101 (N_9101,N_8384,N_8705);
and U9102 (N_9102,N_8308,N_8847);
nand U9103 (N_9103,N_8319,N_8932);
nand U9104 (N_9104,N_8791,N_8640);
or U9105 (N_9105,N_8996,N_8698);
or U9106 (N_9106,N_8336,N_8648);
nor U9107 (N_9107,N_8377,N_8338);
and U9108 (N_9108,N_8782,N_8576);
or U9109 (N_9109,N_8890,N_8435);
or U9110 (N_9110,N_8557,N_8677);
nor U9111 (N_9111,N_8650,N_8608);
nor U9112 (N_9112,N_8449,N_8666);
nor U9113 (N_9113,N_8927,N_8947);
and U9114 (N_9114,N_8551,N_8404);
nor U9115 (N_9115,N_8687,N_8667);
and U9116 (N_9116,N_8885,N_8672);
or U9117 (N_9117,N_8792,N_8264);
or U9118 (N_9118,N_8875,N_8273);
nor U9119 (N_9119,N_8708,N_8761);
or U9120 (N_9120,N_8605,N_8862);
or U9121 (N_9121,N_8937,N_8664);
and U9122 (N_9122,N_8821,N_8852);
or U9123 (N_9123,N_8266,N_8418);
xor U9124 (N_9124,N_8294,N_8606);
nand U9125 (N_9125,N_8534,N_8508);
nand U9126 (N_9126,N_8988,N_8305);
nand U9127 (N_9127,N_8917,N_8524);
nand U9128 (N_9128,N_8310,N_8856);
xor U9129 (N_9129,N_8560,N_8272);
nand U9130 (N_9130,N_8323,N_8542);
nor U9131 (N_9131,N_8437,N_8833);
or U9132 (N_9132,N_8564,N_8933);
nand U9133 (N_9133,N_8466,N_8494);
nor U9134 (N_9134,N_8422,N_8669);
and U9135 (N_9135,N_8627,N_8496);
nand U9136 (N_9136,N_8425,N_8309);
nor U9137 (N_9137,N_8481,N_8701);
and U9138 (N_9138,N_8943,N_8301);
and U9139 (N_9139,N_8733,N_8809);
nor U9140 (N_9140,N_8959,N_8816);
and U9141 (N_9141,N_8413,N_8878);
and U9142 (N_9142,N_8922,N_8939);
nor U9143 (N_9143,N_8530,N_8300);
nor U9144 (N_9144,N_8750,N_8691);
and U9145 (N_9145,N_8457,N_8279);
nor U9146 (N_9146,N_8655,N_8670);
nor U9147 (N_9147,N_8383,N_8262);
nor U9148 (N_9148,N_8854,N_8515);
nand U9149 (N_9149,N_8629,N_8444);
or U9150 (N_9150,N_8261,N_8774);
and U9151 (N_9151,N_8482,N_8469);
nand U9152 (N_9152,N_8797,N_8442);
or U9153 (N_9153,N_8448,N_8681);
and U9154 (N_9154,N_8289,N_8537);
xor U9155 (N_9155,N_8375,N_8403);
nor U9156 (N_9156,N_8882,N_8371);
nand U9157 (N_9157,N_8759,N_8332);
nand U9158 (N_9158,N_8770,N_8286);
nand U9159 (N_9159,N_8891,N_8938);
nor U9160 (N_9160,N_8773,N_8612);
nor U9161 (N_9161,N_8789,N_8794);
nor U9162 (N_9162,N_8951,N_8946);
nor U9163 (N_9163,N_8516,N_8538);
and U9164 (N_9164,N_8634,N_8326);
nor U9165 (N_9165,N_8909,N_8382);
and U9166 (N_9166,N_8824,N_8997);
nand U9167 (N_9167,N_8586,N_8887);
or U9168 (N_9168,N_8656,N_8870);
or U9169 (N_9169,N_8973,N_8736);
nand U9170 (N_9170,N_8290,N_8282);
and U9171 (N_9171,N_8617,N_8588);
and U9172 (N_9172,N_8561,N_8994);
or U9173 (N_9173,N_8730,N_8409);
and U9174 (N_9174,N_8622,N_8602);
or U9175 (N_9175,N_8803,N_8509);
nand U9176 (N_9176,N_8892,N_8427);
nand U9177 (N_9177,N_8765,N_8762);
nand U9178 (N_9178,N_8325,N_8945);
and U9179 (N_9179,N_8529,N_8270);
nor U9180 (N_9180,N_8468,N_8291);
or U9181 (N_9181,N_8747,N_8758);
or U9182 (N_9182,N_8864,N_8583);
and U9183 (N_9183,N_8810,N_8510);
nand U9184 (N_9184,N_8467,N_8707);
and U9185 (N_9185,N_8591,N_8523);
nor U9186 (N_9186,N_8465,N_8410);
or U9187 (N_9187,N_8421,N_8379);
or U9188 (N_9188,N_8683,N_8646);
and U9189 (N_9189,N_8751,N_8636);
nor U9190 (N_9190,N_8397,N_8260);
nand U9191 (N_9191,N_8965,N_8275);
nor U9192 (N_9192,N_8445,N_8877);
nor U9193 (N_9193,N_8936,N_8727);
nor U9194 (N_9194,N_8253,N_8961);
nand U9195 (N_9195,N_8836,N_8414);
and U9196 (N_9196,N_8800,N_8552);
nor U9197 (N_9197,N_8543,N_8307);
and U9198 (N_9198,N_8395,N_8764);
xnor U9199 (N_9199,N_8860,N_8987);
xor U9200 (N_9200,N_8753,N_8531);
or U9201 (N_9201,N_8578,N_8971);
and U9202 (N_9202,N_8904,N_8964);
nor U9203 (N_9203,N_8915,N_8846);
or U9204 (N_9204,N_8989,N_8474);
xor U9205 (N_9205,N_8920,N_8599);
or U9206 (N_9206,N_8855,N_8280);
nor U9207 (N_9207,N_8834,N_8981);
or U9208 (N_9208,N_8778,N_8434);
or U9209 (N_9209,N_8832,N_8977);
xor U9210 (N_9210,N_8416,N_8718);
or U9211 (N_9211,N_8575,N_8505);
or U9212 (N_9212,N_8429,N_8473);
nand U9213 (N_9213,N_8380,N_8501);
and U9214 (N_9214,N_8635,N_8373);
nand U9215 (N_9215,N_8929,N_8630);
nand U9216 (N_9216,N_8982,N_8883);
or U9217 (N_9217,N_8329,N_8254);
or U9218 (N_9218,N_8858,N_8901);
or U9219 (N_9219,N_8393,N_8706);
and U9220 (N_9220,N_8777,N_8665);
or U9221 (N_9221,N_8333,N_8499);
nand U9222 (N_9222,N_8808,N_8680);
and U9223 (N_9223,N_8539,N_8470);
nand U9224 (N_9224,N_8659,N_8954);
and U9225 (N_9225,N_8318,N_8331);
nor U9226 (N_9226,N_8637,N_8363);
nor U9227 (N_9227,N_8620,N_8710);
or U9228 (N_9228,N_8431,N_8563);
and U9229 (N_9229,N_8734,N_8359);
nor U9230 (N_9230,N_8549,N_8259);
and U9231 (N_9231,N_8881,N_8895);
or U9232 (N_9232,N_8284,N_8299);
and U9233 (N_9233,N_8344,N_8547);
nand U9234 (N_9234,N_8893,N_8296);
nor U9235 (N_9235,N_8360,N_8998);
or U9236 (N_9236,N_8577,N_8876);
or U9237 (N_9237,N_8719,N_8740);
nor U9238 (N_9238,N_8616,N_8757);
xor U9239 (N_9239,N_8908,N_8281);
or U9240 (N_9240,N_8558,N_8545);
nand U9241 (N_9241,N_8258,N_8292);
or U9242 (N_9242,N_8314,N_8829);
or U9243 (N_9243,N_8354,N_8679);
and U9244 (N_9244,N_8507,N_8579);
nor U9245 (N_9245,N_8533,N_8400);
and U9246 (N_9246,N_8376,N_8657);
nor U9247 (N_9247,N_8737,N_8283);
xor U9248 (N_9248,N_8914,N_8752);
or U9249 (N_9249,N_8748,N_8611);
or U9250 (N_9250,N_8991,N_8625);
nand U9251 (N_9251,N_8386,N_8461);
nand U9252 (N_9252,N_8715,N_8340);
nand U9253 (N_9253,N_8879,N_8693);
nand U9254 (N_9254,N_8972,N_8594);
or U9255 (N_9255,N_8654,N_8984);
and U9256 (N_9256,N_8607,N_8392);
and U9257 (N_9257,N_8807,N_8787);
or U9258 (N_9258,N_8306,N_8688);
or U9259 (N_9259,N_8717,N_8690);
or U9260 (N_9260,N_8568,N_8500);
or U9261 (N_9261,N_8674,N_8873);
or U9262 (N_9262,N_8983,N_8897);
or U9263 (N_9263,N_8903,N_8556);
nor U9264 (N_9264,N_8783,N_8358);
or U9265 (N_9265,N_8256,N_8886);
nor U9266 (N_9266,N_8408,N_8955);
nand U9267 (N_9267,N_8621,N_8426);
and U9268 (N_9268,N_8593,N_8695);
nand U9269 (N_9269,N_8805,N_8339);
nand U9270 (N_9270,N_8453,N_8250);
nand U9271 (N_9271,N_8369,N_8944);
or U9272 (N_9272,N_8653,N_8571);
nor U9273 (N_9273,N_8484,N_8732);
and U9274 (N_9274,N_8699,N_8398);
nor U9275 (N_9275,N_8324,N_8798);
and U9276 (N_9276,N_8738,N_8550);
and U9277 (N_9277,N_8298,N_8763);
or U9278 (N_9278,N_8488,N_8471);
nand U9279 (N_9279,N_8776,N_8755);
nand U9280 (N_9280,N_8322,N_8696);
nand U9281 (N_9281,N_8267,N_8569);
nand U9282 (N_9282,N_8838,N_8960);
nor U9283 (N_9283,N_8702,N_8990);
or U9284 (N_9284,N_8742,N_8722);
or U9285 (N_9285,N_8970,N_8780);
and U9286 (N_9286,N_8999,N_8388);
nand U9287 (N_9287,N_8979,N_8790);
and U9288 (N_9288,N_8317,N_8900);
and U9289 (N_9289,N_8849,N_8756);
nor U9290 (N_9290,N_8992,N_8463);
or U9291 (N_9291,N_8995,N_8948);
or U9292 (N_9292,N_8562,N_8811);
or U9293 (N_9293,N_8861,N_8349);
and U9294 (N_9294,N_8825,N_8345);
nand U9295 (N_9295,N_8464,N_8517);
nand U9296 (N_9296,N_8480,N_8311);
and U9297 (N_9297,N_8826,N_8574);
or U9298 (N_9298,N_8592,N_8483);
and U9299 (N_9299,N_8935,N_8420);
nand U9300 (N_9300,N_8928,N_8604);
and U9301 (N_9301,N_8785,N_8623);
nor U9302 (N_9302,N_8328,N_8385);
nor U9303 (N_9303,N_8660,N_8899);
and U9304 (N_9304,N_8601,N_8486);
and U9305 (N_9305,N_8402,N_8713);
xor U9306 (N_9306,N_8812,N_8614);
or U9307 (N_9307,N_8417,N_8827);
nor U9308 (N_9308,N_8544,N_8274);
nand U9309 (N_9309,N_8372,N_8950);
nand U9310 (N_9310,N_8731,N_8641);
nand U9311 (N_9311,N_8631,N_8366);
nor U9312 (N_9312,N_8974,N_8626);
or U9313 (N_9313,N_8455,N_8590);
nor U9314 (N_9314,N_8953,N_8919);
or U9315 (N_9315,N_8644,N_8430);
or U9316 (N_9316,N_8526,N_8723);
or U9317 (N_9317,N_8478,N_8458);
nand U9318 (N_9318,N_8728,N_8370);
nor U9319 (N_9319,N_8703,N_8297);
nor U9320 (N_9320,N_8969,N_8835);
or U9321 (N_9321,N_8857,N_8926);
nand U9322 (N_9322,N_8541,N_8963);
or U9323 (N_9323,N_8668,N_8754);
nand U9324 (N_9324,N_8603,N_8263);
nand U9325 (N_9325,N_8729,N_8347);
nand U9326 (N_9326,N_8535,N_8872);
or U9327 (N_9327,N_8912,N_8819);
and U9328 (N_9328,N_8839,N_8485);
and U9329 (N_9329,N_8850,N_8692);
or U9330 (N_9330,N_8968,N_8916);
nand U9331 (N_9331,N_8337,N_8293);
nand U9332 (N_9332,N_8700,N_8842);
or U9333 (N_9333,N_8769,N_8548);
nand U9334 (N_9334,N_8394,N_8684);
and U9335 (N_9335,N_8390,N_8866);
nand U9336 (N_9336,N_8615,N_8815);
nor U9337 (N_9337,N_8788,N_8330);
and U9338 (N_9338,N_8351,N_8257);
and U9339 (N_9339,N_8312,N_8519);
nor U9340 (N_9340,N_8381,N_8712);
or U9341 (N_9341,N_8837,N_8804);
and U9342 (N_9342,N_8746,N_8934);
or U9343 (N_9343,N_8906,N_8433);
nor U9344 (N_9344,N_8744,N_8884);
nand U9345 (N_9345,N_8784,N_8399);
and U9346 (N_9346,N_8406,N_8868);
nand U9347 (N_9347,N_8476,N_8357);
nor U9348 (N_9348,N_8942,N_8976);
or U9349 (N_9349,N_8663,N_8506);
nand U9350 (N_9350,N_8745,N_8793);
and U9351 (N_9351,N_8993,N_8491);
nand U9352 (N_9352,N_8709,N_8910);
and U9353 (N_9353,N_8436,N_8923);
nor U9354 (N_9354,N_8678,N_8251);
and U9355 (N_9355,N_8477,N_8799);
or U9356 (N_9356,N_8828,N_8956);
nor U9357 (N_9357,N_8443,N_8451);
nand U9358 (N_9358,N_8567,N_8472);
nor U9359 (N_9359,N_8632,N_8628);
nor U9360 (N_9360,N_8342,N_8962);
or U9361 (N_9361,N_8779,N_8440);
and U9362 (N_9362,N_8492,N_8364);
nor U9363 (N_9363,N_8321,N_8711);
nor U9364 (N_9364,N_8352,N_8689);
or U9365 (N_9365,N_8913,N_8930);
nand U9366 (N_9366,N_8450,N_8741);
and U9367 (N_9367,N_8459,N_8771);
nor U9368 (N_9368,N_8781,N_8356);
nand U9369 (N_9369,N_8958,N_8831);
nand U9370 (N_9370,N_8353,N_8902);
nor U9371 (N_9371,N_8412,N_8361);
nor U9372 (N_9372,N_8573,N_8518);
or U9373 (N_9373,N_8589,N_8368);
and U9374 (N_9374,N_8566,N_8957);
or U9375 (N_9375,N_8419,N_8587);
nor U9376 (N_9376,N_8869,N_8973);
nor U9377 (N_9377,N_8415,N_8460);
nor U9378 (N_9378,N_8693,N_8920);
nand U9379 (N_9379,N_8882,N_8466);
nand U9380 (N_9380,N_8475,N_8577);
nor U9381 (N_9381,N_8790,N_8491);
and U9382 (N_9382,N_8601,N_8743);
nand U9383 (N_9383,N_8825,N_8886);
or U9384 (N_9384,N_8630,N_8698);
and U9385 (N_9385,N_8751,N_8816);
and U9386 (N_9386,N_8858,N_8747);
nand U9387 (N_9387,N_8933,N_8395);
nand U9388 (N_9388,N_8762,N_8518);
nand U9389 (N_9389,N_8323,N_8447);
xnor U9390 (N_9390,N_8968,N_8653);
or U9391 (N_9391,N_8582,N_8885);
nor U9392 (N_9392,N_8320,N_8865);
nor U9393 (N_9393,N_8813,N_8676);
or U9394 (N_9394,N_8843,N_8303);
and U9395 (N_9395,N_8661,N_8837);
or U9396 (N_9396,N_8976,N_8512);
nand U9397 (N_9397,N_8898,N_8994);
or U9398 (N_9398,N_8990,N_8576);
and U9399 (N_9399,N_8554,N_8640);
nor U9400 (N_9400,N_8636,N_8416);
nand U9401 (N_9401,N_8453,N_8976);
nor U9402 (N_9402,N_8878,N_8885);
or U9403 (N_9403,N_8270,N_8715);
nor U9404 (N_9404,N_8576,N_8410);
nor U9405 (N_9405,N_8720,N_8727);
xor U9406 (N_9406,N_8842,N_8817);
nor U9407 (N_9407,N_8644,N_8402);
and U9408 (N_9408,N_8936,N_8702);
nor U9409 (N_9409,N_8645,N_8661);
nand U9410 (N_9410,N_8734,N_8617);
nor U9411 (N_9411,N_8345,N_8937);
and U9412 (N_9412,N_8969,N_8288);
nor U9413 (N_9413,N_8933,N_8548);
nor U9414 (N_9414,N_8777,N_8950);
or U9415 (N_9415,N_8433,N_8866);
nor U9416 (N_9416,N_8699,N_8722);
nand U9417 (N_9417,N_8629,N_8265);
nor U9418 (N_9418,N_8672,N_8311);
nand U9419 (N_9419,N_8935,N_8741);
or U9420 (N_9420,N_8617,N_8576);
nand U9421 (N_9421,N_8895,N_8803);
or U9422 (N_9422,N_8302,N_8628);
nor U9423 (N_9423,N_8897,N_8740);
nand U9424 (N_9424,N_8818,N_8353);
and U9425 (N_9425,N_8416,N_8926);
nor U9426 (N_9426,N_8558,N_8670);
nor U9427 (N_9427,N_8502,N_8717);
nand U9428 (N_9428,N_8587,N_8414);
xnor U9429 (N_9429,N_8358,N_8719);
nand U9430 (N_9430,N_8935,N_8395);
or U9431 (N_9431,N_8712,N_8973);
nor U9432 (N_9432,N_8444,N_8476);
xor U9433 (N_9433,N_8772,N_8367);
nand U9434 (N_9434,N_8863,N_8640);
and U9435 (N_9435,N_8633,N_8491);
or U9436 (N_9436,N_8951,N_8420);
nand U9437 (N_9437,N_8390,N_8890);
or U9438 (N_9438,N_8930,N_8829);
nand U9439 (N_9439,N_8671,N_8862);
nand U9440 (N_9440,N_8418,N_8414);
xor U9441 (N_9441,N_8829,N_8665);
nand U9442 (N_9442,N_8906,N_8705);
or U9443 (N_9443,N_8643,N_8310);
nor U9444 (N_9444,N_8603,N_8491);
and U9445 (N_9445,N_8548,N_8296);
and U9446 (N_9446,N_8958,N_8785);
nand U9447 (N_9447,N_8709,N_8507);
nand U9448 (N_9448,N_8872,N_8442);
and U9449 (N_9449,N_8678,N_8720);
or U9450 (N_9450,N_8894,N_8305);
nand U9451 (N_9451,N_8822,N_8369);
or U9452 (N_9452,N_8838,N_8852);
nand U9453 (N_9453,N_8935,N_8441);
or U9454 (N_9454,N_8621,N_8917);
or U9455 (N_9455,N_8625,N_8457);
nor U9456 (N_9456,N_8413,N_8661);
nand U9457 (N_9457,N_8980,N_8903);
and U9458 (N_9458,N_8843,N_8565);
nand U9459 (N_9459,N_8303,N_8394);
nand U9460 (N_9460,N_8422,N_8480);
nand U9461 (N_9461,N_8644,N_8631);
and U9462 (N_9462,N_8386,N_8872);
and U9463 (N_9463,N_8850,N_8843);
xnor U9464 (N_9464,N_8984,N_8536);
or U9465 (N_9465,N_8320,N_8699);
nor U9466 (N_9466,N_8877,N_8374);
nand U9467 (N_9467,N_8372,N_8928);
nor U9468 (N_9468,N_8580,N_8491);
nor U9469 (N_9469,N_8876,N_8864);
and U9470 (N_9470,N_8379,N_8448);
nor U9471 (N_9471,N_8791,N_8421);
and U9472 (N_9472,N_8569,N_8311);
nand U9473 (N_9473,N_8256,N_8326);
and U9474 (N_9474,N_8744,N_8600);
nand U9475 (N_9475,N_8896,N_8450);
nor U9476 (N_9476,N_8459,N_8521);
nand U9477 (N_9477,N_8605,N_8873);
nand U9478 (N_9478,N_8518,N_8669);
and U9479 (N_9479,N_8827,N_8493);
nand U9480 (N_9480,N_8699,N_8516);
or U9481 (N_9481,N_8924,N_8795);
nor U9482 (N_9482,N_8603,N_8672);
nor U9483 (N_9483,N_8350,N_8399);
nand U9484 (N_9484,N_8806,N_8346);
nand U9485 (N_9485,N_8298,N_8855);
or U9486 (N_9486,N_8374,N_8561);
nor U9487 (N_9487,N_8276,N_8371);
and U9488 (N_9488,N_8456,N_8466);
nor U9489 (N_9489,N_8631,N_8467);
or U9490 (N_9490,N_8960,N_8280);
and U9491 (N_9491,N_8591,N_8396);
and U9492 (N_9492,N_8952,N_8673);
and U9493 (N_9493,N_8264,N_8405);
and U9494 (N_9494,N_8514,N_8266);
nor U9495 (N_9495,N_8710,N_8459);
nand U9496 (N_9496,N_8612,N_8478);
nand U9497 (N_9497,N_8985,N_8282);
and U9498 (N_9498,N_8856,N_8374);
and U9499 (N_9499,N_8843,N_8993);
or U9500 (N_9500,N_8370,N_8468);
and U9501 (N_9501,N_8965,N_8262);
or U9502 (N_9502,N_8411,N_8946);
nand U9503 (N_9503,N_8306,N_8776);
and U9504 (N_9504,N_8927,N_8545);
nor U9505 (N_9505,N_8863,N_8429);
nand U9506 (N_9506,N_8538,N_8988);
nor U9507 (N_9507,N_8529,N_8474);
nand U9508 (N_9508,N_8461,N_8284);
or U9509 (N_9509,N_8349,N_8310);
nand U9510 (N_9510,N_8599,N_8934);
nor U9511 (N_9511,N_8396,N_8823);
xor U9512 (N_9512,N_8988,N_8261);
xor U9513 (N_9513,N_8468,N_8451);
or U9514 (N_9514,N_8346,N_8302);
and U9515 (N_9515,N_8994,N_8648);
nor U9516 (N_9516,N_8616,N_8658);
nor U9517 (N_9517,N_8382,N_8723);
or U9518 (N_9518,N_8974,N_8509);
nand U9519 (N_9519,N_8717,N_8671);
or U9520 (N_9520,N_8989,N_8836);
nor U9521 (N_9521,N_8354,N_8849);
or U9522 (N_9522,N_8260,N_8438);
nand U9523 (N_9523,N_8258,N_8969);
nor U9524 (N_9524,N_8838,N_8917);
nor U9525 (N_9525,N_8877,N_8829);
nor U9526 (N_9526,N_8614,N_8640);
or U9527 (N_9527,N_8687,N_8495);
nor U9528 (N_9528,N_8647,N_8588);
or U9529 (N_9529,N_8431,N_8419);
nor U9530 (N_9530,N_8568,N_8679);
and U9531 (N_9531,N_8643,N_8850);
and U9532 (N_9532,N_8942,N_8426);
nor U9533 (N_9533,N_8797,N_8826);
xor U9534 (N_9534,N_8440,N_8696);
xor U9535 (N_9535,N_8250,N_8420);
or U9536 (N_9536,N_8855,N_8807);
nor U9537 (N_9537,N_8525,N_8550);
and U9538 (N_9538,N_8753,N_8862);
nand U9539 (N_9539,N_8365,N_8647);
nor U9540 (N_9540,N_8870,N_8977);
and U9541 (N_9541,N_8331,N_8573);
and U9542 (N_9542,N_8937,N_8800);
or U9543 (N_9543,N_8450,N_8283);
or U9544 (N_9544,N_8802,N_8965);
nor U9545 (N_9545,N_8622,N_8254);
nand U9546 (N_9546,N_8489,N_8955);
or U9547 (N_9547,N_8554,N_8803);
and U9548 (N_9548,N_8368,N_8260);
and U9549 (N_9549,N_8309,N_8687);
and U9550 (N_9550,N_8574,N_8614);
nor U9551 (N_9551,N_8652,N_8672);
or U9552 (N_9552,N_8257,N_8719);
nor U9553 (N_9553,N_8343,N_8351);
nand U9554 (N_9554,N_8889,N_8904);
or U9555 (N_9555,N_8940,N_8481);
nor U9556 (N_9556,N_8348,N_8620);
nand U9557 (N_9557,N_8747,N_8634);
or U9558 (N_9558,N_8574,N_8429);
nand U9559 (N_9559,N_8284,N_8336);
nand U9560 (N_9560,N_8472,N_8379);
xnor U9561 (N_9561,N_8534,N_8611);
nor U9562 (N_9562,N_8470,N_8559);
nand U9563 (N_9563,N_8579,N_8924);
or U9564 (N_9564,N_8506,N_8560);
or U9565 (N_9565,N_8603,N_8914);
nor U9566 (N_9566,N_8297,N_8673);
nand U9567 (N_9567,N_8754,N_8419);
nor U9568 (N_9568,N_8253,N_8461);
or U9569 (N_9569,N_8546,N_8664);
and U9570 (N_9570,N_8461,N_8309);
or U9571 (N_9571,N_8283,N_8377);
nor U9572 (N_9572,N_8452,N_8517);
nor U9573 (N_9573,N_8428,N_8612);
nand U9574 (N_9574,N_8706,N_8642);
or U9575 (N_9575,N_8986,N_8755);
nand U9576 (N_9576,N_8697,N_8728);
or U9577 (N_9577,N_8570,N_8582);
or U9578 (N_9578,N_8318,N_8305);
or U9579 (N_9579,N_8984,N_8825);
or U9580 (N_9580,N_8985,N_8299);
nand U9581 (N_9581,N_8649,N_8945);
and U9582 (N_9582,N_8424,N_8335);
nor U9583 (N_9583,N_8267,N_8418);
and U9584 (N_9584,N_8617,N_8571);
nor U9585 (N_9585,N_8697,N_8456);
or U9586 (N_9586,N_8977,N_8555);
or U9587 (N_9587,N_8871,N_8820);
nor U9588 (N_9588,N_8894,N_8667);
nor U9589 (N_9589,N_8691,N_8978);
nand U9590 (N_9590,N_8876,N_8311);
and U9591 (N_9591,N_8338,N_8339);
and U9592 (N_9592,N_8467,N_8684);
nor U9593 (N_9593,N_8991,N_8795);
nor U9594 (N_9594,N_8743,N_8571);
or U9595 (N_9595,N_8576,N_8760);
or U9596 (N_9596,N_8922,N_8949);
nor U9597 (N_9597,N_8705,N_8433);
nand U9598 (N_9598,N_8586,N_8270);
xnor U9599 (N_9599,N_8875,N_8397);
nand U9600 (N_9600,N_8929,N_8476);
nand U9601 (N_9601,N_8706,N_8589);
and U9602 (N_9602,N_8694,N_8971);
or U9603 (N_9603,N_8529,N_8566);
or U9604 (N_9604,N_8614,N_8588);
nor U9605 (N_9605,N_8509,N_8383);
or U9606 (N_9606,N_8674,N_8820);
and U9607 (N_9607,N_8666,N_8788);
or U9608 (N_9608,N_8614,N_8629);
or U9609 (N_9609,N_8410,N_8905);
and U9610 (N_9610,N_8846,N_8740);
nor U9611 (N_9611,N_8457,N_8824);
or U9612 (N_9612,N_8288,N_8683);
nor U9613 (N_9613,N_8852,N_8686);
and U9614 (N_9614,N_8763,N_8656);
nor U9615 (N_9615,N_8693,N_8880);
or U9616 (N_9616,N_8503,N_8352);
and U9617 (N_9617,N_8468,N_8375);
nor U9618 (N_9618,N_8794,N_8688);
and U9619 (N_9619,N_8807,N_8399);
xor U9620 (N_9620,N_8754,N_8600);
xnor U9621 (N_9621,N_8708,N_8798);
or U9622 (N_9622,N_8963,N_8341);
xor U9623 (N_9623,N_8822,N_8930);
nand U9624 (N_9624,N_8887,N_8931);
nand U9625 (N_9625,N_8264,N_8748);
and U9626 (N_9626,N_8758,N_8292);
and U9627 (N_9627,N_8842,N_8981);
or U9628 (N_9628,N_8817,N_8908);
or U9629 (N_9629,N_8393,N_8577);
nor U9630 (N_9630,N_8788,N_8553);
nor U9631 (N_9631,N_8633,N_8658);
nor U9632 (N_9632,N_8779,N_8939);
nand U9633 (N_9633,N_8642,N_8352);
nand U9634 (N_9634,N_8786,N_8294);
or U9635 (N_9635,N_8850,N_8286);
or U9636 (N_9636,N_8567,N_8414);
xnor U9637 (N_9637,N_8745,N_8405);
nor U9638 (N_9638,N_8782,N_8876);
nand U9639 (N_9639,N_8293,N_8396);
nand U9640 (N_9640,N_8912,N_8687);
or U9641 (N_9641,N_8609,N_8277);
nor U9642 (N_9642,N_8486,N_8725);
nor U9643 (N_9643,N_8504,N_8503);
and U9644 (N_9644,N_8428,N_8922);
xnor U9645 (N_9645,N_8714,N_8970);
or U9646 (N_9646,N_8310,N_8597);
or U9647 (N_9647,N_8831,N_8549);
and U9648 (N_9648,N_8654,N_8862);
and U9649 (N_9649,N_8907,N_8882);
nand U9650 (N_9650,N_8827,N_8716);
or U9651 (N_9651,N_8280,N_8478);
or U9652 (N_9652,N_8634,N_8560);
nand U9653 (N_9653,N_8534,N_8750);
or U9654 (N_9654,N_8290,N_8788);
and U9655 (N_9655,N_8839,N_8259);
nand U9656 (N_9656,N_8304,N_8413);
and U9657 (N_9657,N_8757,N_8621);
nor U9658 (N_9658,N_8640,N_8770);
and U9659 (N_9659,N_8616,N_8888);
xor U9660 (N_9660,N_8678,N_8304);
or U9661 (N_9661,N_8365,N_8947);
or U9662 (N_9662,N_8611,N_8552);
nor U9663 (N_9663,N_8308,N_8760);
and U9664 (N_9664,N_8309,N_8768);
nor U9665 (N_9665,N_8885,N_8953);
nand U9666 (N_9666,N_8968,N_8862);
nor U9667 (N_9667,N_8484,N_8989);
nor U9668 (N_9668,N_8712,N_8742);
xnor U9669 (N_9669,N_8976,N_8650);
nand U9670 (N_9670,N_8801,N_8732);
nor U9671 (N_9671,N_8381,N_8535);
and U9672 (N_9672,N_8257,N_8516);
or U9673 (N_9673,N_8929,N_8383);
nand U9674 (N_9674,N_8550,N_8501);
or U9675 (N_9675,N_8638,N_8456);
nor U9676 (N_9676,N_8908,N_8848);
xor U9677 (N_9677,N_8942,N_8439);
or U9678 (N_9678,N_8838,N_8407);
and U9679 (N_9679,N_8471,N_8425);
nand U9680 (N_9680,N_8791,N_8799);
nand U9681 (N_9681,N_8757,N_8359);
nor U9682 (N_9682,N_8750,N_8735);
nand U9683 (N_9683,N_8436,N_8714);
or U9684 (N_9684,N_8292,N_8439);
xor U9685 (N_9685,N_8567,N_8708);
nand U9686 (N_9686,N_8983,N_8503);
or U9687 (N_9687,N_8297,N_8501);
nand U9688 (N_9688,N_8290,N_8878);
nor U9689 (N_9689,N_8411,N_8818);
and U9690 (N_9690,N_8668,N_8354);
nor U9691 (N_9691,N_8367,N_8965);
and U9692 (N_9692,N_8271,N_8433);
nor U9693 (N_9693,N_8376,N_8398);
and U9694 (N_9694,N_8968,N_8902);
nand U9695 (N_9695,N_8311,N_8267);
and U9696 (N_9696,N_8862,N_8394);
nand U9697 (N_9697,N_8693,N_8615);
and U9698 (N_9698,N_8653,N_8951);
or U9699 (N_9699,N_8735,N_8278);
nand U9700 (N_9700,N_8306,N_8730);
nor U9701 (N_9701,N_8914,N_8311);
and U9702 (N_9702,N_8258,N_8687);
nand U9703 (N_9703,N_8692,N_8838);
nand U9704 (N_9704,N_8518,N_8661);
nor U9705 (N_9705,N_8662,N_8710);
and U9706 (N_9706,N_8947,N_8719);
nand U9707 (N_9707,N_8593,N_8806);
nand U9708 (N_9708,N_8650,N_8412);
or U9709 (N_9709,N_8424,N_8647);
or U9710 (N_9710,N_8936,N_8715);
nor U9711 (N_9711,N_8780,N_8805);
nand U9712 (N_9712,N_8338,N_8448);
or U9713 (N_9713,N_8815,N_8281);
nor U9714 (N_9714,N_8255,N_8902);
nor U9715 (N_9715,N_8549,N_8942);
and U9716 (N_9716,N_8772,N_8887);
and U9717 (N_9717,N_8357,N_8301);
nor U9718 (N_9718,N_8718,N_8981);
nor U9719 (N_9719,N_8966,N_8509);
and U9720 (N_9720,N_8667,N_8457);
nor U9721 (N_9721,N_8603,N_8582);
nand U9722 (N_9722,N_8729,N_8563);
nor U9723 (N_9723,N_8927,N_8775);
nor U9724 (N_9724,N_8872,N_8877);
nand U9725 (N_9725,N_8547,N_8306);
nand U9726 (N_9726,N_8472,N_8576);
or U9727 (N_9727,N_8980,N_8509);
or U9728 (N_9728,N_8464,N_8528);
and U9729 (N_9729,N_8470,N_8352);
and U9730 (N_9730,N_8955,N_8353);
nor U9731 (N_9731,N_8806,N_8813);
or U9732 (N_9732,N_8526,N_8366);
nand U9733 (N_9733,N_8368,N_8623);
or U9734 (N_9734,N_8438,N_8993);
or U9735 (N_9735,N_8790,N_8493);
or U9736 (N_9736,N_8413,N_8332);
and U9737 (N_9737,N_8909,N_8582);
and U9738 (N_9738,N_8819,N_8289);
and U9739 (N_9739,N_8713,N_8407);
nand U9740 (N_9740,N_8356,N_8922);
nor U9741 (N_9741,N_8262,N_8416);
nand U9742 (N_9742,N_8628,N_8679);
and U9743 (N_9743,N_8359,N_8314);
or U9744 (N_9744,N_8897,N_8505);
and U9745 (N_9745,N_8279,N_8648);
or U9746 (N_9746,N_8935,N_8925);
and U9747 (N_9747,N_8464,N_8302);
nand U9748 (N_9748,N_8818,N_8797);
nand U9749 (N_9749,N_8840,N_8263);
nor U9750 (N_9750,N_9455,N_9147);
nor U9751 (N_9751,N_9724,N_9504);
or U9752 (N_9752,N_9588,N_9552);
nor U9753 (N_9753,N_9093,N_9076);
nor U9754 (N_9754,N_9451,N_9159);
nand U9755 (N_9755,N_9520,N_9425);
nand U9756 (N_9756,N_9171,N_9363);
or U9757 (N_9757,N_9044,N_9053);
nand U9758 (N_9758,N_9129,N_9556);
nand U9759 (N_9759,N_9305,N_9017);
and U9760 (N_9760,N_9563,N_9679);
nand U9761 (N_9761,N_9394,N_9025);
and U9762 (N_9762,N_9304,N_9105);
nand U9763 (N_9763,N_9663,N_9510);
nor U9764 (N_9764,N_9458,N_9172);
nor U9765 (N_9765,N_9593,N_9306);
nor U9766 (N_9766,N_9100,N_9562);
and U9767 (N_9767,N_9207,N_9448);
nand U9768 (N_9768,N_9364,N_9347);
and U9769 (N_9769,N_9694,N_9617);
xor U9770 (N_9770,N_9126,N_9028);
nand U9771 (N_9771,N_9365,N_9484);
or U9772 (N_9772,N_9567,N_9517);
nor U9773 (N_9773,N_9161,N_9537);
or U9774 (N_9774,N_9378,N_9477);
and U9775 (N_9775,N_9142,N_9439);
nand U9776 (N_9776,N_9581,N_9578);
nand U9777 (N_9777,N_9734,N_9356);
or U9778 (N_9778,N_9672,N_9324);
and U9779 (N_9779,N_9070,N_9460);
or U9780 (N_9780,N_9635,N_9216);
nor U9781 (N_9781,N_9124,N_9587);
or U9782 (N_9782,N_9265,N_9243);
nor U9783 (N_9783,N_9241,N_9113);
nor U9784 (N_9784,N_9175,N_9741);
nor U9785 (N_9785,N_9374,N_9647);
and U9786 (N_9786,N_9162,N_9598);
nand U9787 (N_9787,N_9538,N_9157);
and U9788 (N_9788,N_9329,N_9259);
or U9789 (N_9789,N_9335,N_9426);
nand U9790 (N_9790,N_9287,N_9185);
and U9791 (N_9791,N_9037,N_9186);
nor U9792 (N_9792,N_9453,N_9196);
and U9793 (N_9793,N_9518,N_9383);
or U9794 (N_9794,N_9639,N_9716);
nand U9795 (N_9795,N_9532,N_9302);
nor U9796 (N_9796,N_9678,N_9551);
or U9797 (N_9797,N_9295,N_9720);
and U9798 (N_9798,N_9206,N_9475);
and U9799 (N_9799,N_9388,N_9114);
and U9800 (N_9800,N_9472,N_9368);
xnor U9801 (N_9801,N_9691,N_9208);
or U9802 (N_9802,N_9545,N_9275);
or U9803 (N_9803,N_9205,N_9160);
or U9804 (N_9804,N_9533,N_9336);
or U9805 (N_9805,N_9712,N_9634);
nor U9806 (N_9806,N_9568,N_9345);
nand U9807 (N_9807,N_9688,N_9670);
and U9808 (N_9808,N_9132,N_9586);
nand U9809 (N_9809,N_9673,N_9272);
or U9810 (N_9810,N_9267,N_9310);
and U9811 (N_9811,N_9571,N_9456);
nand U9812 (N_9812,N_9318,N_9121);
or U9813 (N_9813,N_9330,N_9400);
or U9814 (N_9814,N_9402,N_9732);
and U9815 (N_9815,N_9440,N_9137);
nand U9816 (N_9816,N_9506,N_9352);
and U9817 (N_9817,N_9705,N_9300);
or U9818 (N_9818,N_9024,N_9219);
xnor U9819 (N_9819,N_9636,N_9508);
nand U9820 (N_9820,N_9700,N_9513);
and U9821 (N_9821,N_9006,N_9245);
or U9822 (N_9822,N_9393,N_9410);
nor U9823 (N_9823,N_9376,N_9084);
or U9824 (N_9824,N_9155,N_9040);
nor U9825 (N_9825,N_9525,N_9495);
or U9826 (N_9826,N_9441,N_9056);
and U9827 (N_9827,N_9248,N_9689);
xor U9828 (N_9828,N_9746,N_9585);
and U9829 (N_9829,N_9001,N_9215);
and U9830 (N_9830,N_9197,N_9150);
nand U9831 (N_9831,N_9645,N_9022);
nor U9832 (N_9832,N_9686,N_9687);
nand U9833 (N_9833,N_9539,N_9511);
nor U9834 (N_9834,N_9187,N_9156);
nor U9835 (N_9835,N_9291,N_9729);
nor U9836 (N_9836,N_9168,N_9622);
nand U9837 (N_9837,N_9173,N_9303);
nor U9838 (N_9838,N_9608,N_9646);
nand U9839 (N_9839,N_9118,N_9462);
nand U9840 (N_9840,N_9583,N_9199);
nor U9841 (N_9841,N_9260,N_9343);
nor U9842 (N_9842,N_9036,N_9109);
or U9843 (N_9843,N_9500,N_9061);
nor U9844 (N_9844,N_9644,N_9169);
nor U9845 (N_9845,N_9503,N_9619);
xor U9846 (N_9846,N_9375,N_9228);
or U9847 (N_9847,N_9317,N_9222);
nor U9848 (N_9848,N_9650,N_9237);
and U9849 (N_9849,N_9027,N_9722);
nor U9850 (N_9850,N_9195,N_9164);
or U9851 (N_9851,N_9629,N_9014);
and U9852 (N_9852,N_9263,N_9311);
nand U9853 (N_9853,N_9693,N_9086);
and U9854 (N_9854,N_9546,N_9102);
or U9855 (N_9855,N_9602,N_9097);
and U9856 (N_9856,N_9294,N_9348);
and U9857 (N_9857,N_9530,N_9561);
and U9858 (N_9858,N_9083,N_9509);
nor U9859 (N_9859,N_9140,N_9605);
nand U9860 (N_9860,N_9564,N_9019);
and U9861 (N_9861,N_9312,N_9529);
xnor U9862 (N_9862,N_9623,N_9667);
or U9863 (N_9863,N_9062,N_9723);
and U9864 (N_9864,N_9038,N_9218);
nand U9865 (N_9865,N_9049,N_9476);
nor U9866 (N_9866,N_9431,N_9346);
and U9867 (N_9867,N_9337,N_9653);
nor U9868 (N_9868,N_9091,N_9406);
or U9869 (N_9869,N_9103,N_9473);
or U9870 (N_9870,N_9380,N_9013);
and U9871 (N_9871,N_9033,N_9544);
or U9872 (N_9872,N_9603,N_9127);
nand U9873 (N_9873,N_9423,N_9643);
or U9874 (N_9874,N_9180,N_9464);
or U9875 (N_9875,N_9029,N_9236);
nor U9876 (N_9876,N_9744,N_9239);
or U9877 (N_9877,N_9514,N_9242);
nand U9878 (N_9878,N_9106,N_9262);
nor U9879 (N_9879,N_9714,N_9289);
nor U9880 (N_9880,N_9193,N_9201);
and U9881 (N_9881,N_9189,N_9035);
and U9882 (N_9882,N_9077,N_9620);
and U9883 (N_9883,N_9377,N_9471);
nor U9884 (N_9884,N_9493,N_9745);
or U9885 (N_9885,N_9735,N_9069);
and U9886 (N_9886,N_9662,N_9680);
or U9887 (N_9887,N_9665,N_9023);
and U9888 (N_9888,N_9307,N_9313);
and U9889 (N_9889,N_9738,N_9386);
nor U9890 (N_9890,N_9618,N_9284);
and U9891 (N_9891,N_9042,N_9470);
or U9892 (N_9892,N_9727,N_9276);
nor U9893 (N_9893,N_9145,N_9015);
nor U9894 (N_9894,N_9490,N_9261);
nor U9895 (N_9895,N_9521,N_9710);
nor U9896 (N_9896,N_9698,N_9413);
nor U9897 (N_9897,N_9491,N_9685);
nand U9898 (N_9898,N_9749,N_9389);
nor U9899 (N_9899,N_9560,N_9512);
nor U9900 (N_9900,N_9652,N_9020);
or U9901 (N_9901,N_9433,N_9519);
or U9902 (N_9902,N_9535,N_9489);
and U9903 (N_9903,N_9104,N_9391);
or U9904 (N_9904,N_9209,N_9463);
and U9905 (N_9905,N_9592,N_9434);
nor U9906 (N_9906,N_9392,N_9554);
nand U9907 (N_9907,N_9094,N_9234);
and U9908 (N_9908,N_9542,N_9548);
nor U9909 (N_9909,N_9321,N_9485);
nand U9910 (N_9910,N_9674,N_9668);
and U9911 (N_9911,N_9480,N_9213);
or U9912 (N_9912,N_9315,N_9204);
or U9913 (N_9913,N_9338,N_9078);
nand U9914 (N_9914,N_9523,N_9405);
nand U9915 (N_9915,N_9611,N_9696);
nor U9916 (N_9916,N_9153,N_9000);
nand U9917 (N_9917,N_9706,N_9010);
nand U9918 (N_9918,N_9606,N_9254);
or U9919 (N_9919,N_9179,N_9681);
or U9920 (N_9920,N_9395,N_9630);
or U9921 (N_9921,N_9115,N_9297);
and U9922 (N_9922,N_9461,N_9522);
nor U9923 (N_9923,N_9403,N_9609);
or U9924 (N_9924,N_9498,N_9449);
or U9925 (N_9925,N_9507,N_9442);
and U9926 (N_9926,N_9005,N_9730);
nor U9927 (N_9927,N_9158,N_9177);
nand U9928 (N_9928,N_9227,N_9266);
or U9929 (N_9929,N_9255,N_9574);
nand U9930 (N_9930,N_9684,N_9366);
nand U9931 (N_9931,N_9117,N_9429);
nor U9932 (N_9932,N_9057,N_9637);
or U9933 (N_9933,N_9610,N_9045);
nand U9934 (N_9934,N_9041,N_9224);
and U9935 (N_9935,N_9494,N_9584);
or U9936 (N_9936,N_9154,N_9360);
nand U9937 (N_9937,N_9194,N_9279);
and U9938 (N_9938,N_9098,N_9200);
and U9939 (N_9939,N_9247,N_9483);
and U9940 (N_9940,N_9183,N_9709);
or U9941 (N_9941,N_9654,N_9089);
and U9942 (N_9942,N_9296,N_9515);
and U9943 (N_9943,N_9580,N_9092);
or U9944 (N_9944,N_9415,N_9600);
nor U9945 (N_9945,N_9531,N_9387);
or U9946 (N_9946,N_9675,N_9435);
nor U9947 (N_9947,N_9334,N_9528);
and U9948 (N_9948,N_9726,N_9065);
or U9949 (N_9949,N_9055,N_9412);
or U9950 (N_9950,N_9235,N_9399);
nand U9951 (N_9951,N_9594,N_9570);
or U9952 (N_9952,N_9176,N_9074);
nand U9953 (N_9953,N_9323,N_9657);
nor U9954 (N_9954,N_9597,N_9695);
and U9955 (N_9955,N_9407,N_9631);
and U9956 (N_9956,N_9058,N_9221);
nor U9957 (N_9957,N_9314,N_9039);
nor U9958 (N_9958,N_9032,N_9566);
and U9959 (N_9959,N_9099,N_9331);
nor U9960 (N_9960,N_9134,N_9640);
xnor U9961 (N_9961,N_9170,N_9527);
nor U9962 (N_9962,N_9690,N_9664);
and U9963 (N_9963,N_9332,N_9450);
or U9964 (N_9964,N_9719,N_9715);
nor U9965 (N_9965,N_9256,N_9085);
nor U9966 (N_9966,N_9488,N_9613);
and U9967 (N_9967,N_9110,N_9016);
nor U9968 (N_9968,N_9012,N_9181);
nor U9969 (N_9969,N_9601,N_9353);
and U9970 (N_9970,N_9088,N_9344);
or U9971 (N_9971,N_9068,N_9178);
nor U9972 (N_9972,N_9326,N_9656);
nor U9973 (N_9973,N_9649,N_9316);
nor U9974 (N_9974,N_9404,N_9379);
nand U9975 (N_9975,N_9051,N_9550);
or U9976 (N_9976,N_9669,N_9271);
or U9977 (N_9977,N_9184,N_9202);
nor U9978 (N_9978,N_9677,N_9615);
xor U9979 (N_9979,N_9486,N_9298);
nor U9980 (N_9980,N_9210,N_9018);
nand U9981 (N_9981,N_9299,N_9090);
and U9982 (N_9982,N_9082,N_9501);
nand U9983 (N_9983,N_9711,N_9063);
xnor U9984 (N_9984,N_9502,N_9301);
xor U9985 (N_9985,N_9682,N_9370);
nand U9986 (N_9986,N_9572,N_9638);
nand U9987 (N_9987,N_9342,N_9725);
nor U9988 (N_9988,N_9211,N_9340);
and U9989 (N_9989,N_9238,N_9430);
nand U9990 (N_9990,N_9064,N_9273);
and U9991 (N_9991,N_9625,N_9167);
xnor U9992 (N_9992,N_9718,N_9264);
nand U9993 (N_9993,N_9354,N_9658);
and U9994 (N_9994,N_9198,N_9736);
nor U9995 (N_9995,N_9231,N_9174);
nor U9996 (N_9996,N_9748,N_9152);
and U9997 (N_9997,N_9457,N_9474);
or U9998 (N_9998,N_9350,N_9701);
or U9999 (N_9999,N_9432,N_9309);
nand U10000 (N_10000,N_9232,N_9163);
xor U10001 (N_10001,N_9582,N_9130);
nand U10002 (N_10002,N_9226,N_9469);
nand U10003 (N_10003,N_9341,N_9497);
nand U10004 (N_10004,N_9351,N_9229);
nor U10005 (N_10005,N_9595,N_9101);
nand U10006 (N_10006,N_9320,N_9059);
nor U10007 (N_10007,N_9139,N_9050);
and U10008 (N_10008,N_9409,N_9288);
nand U10009 (N_10009,N_9671,N_9553);
and U10010 (N_10010,N_9367,N_9481);
nor U10011 (N_10011,N_9541,N_9743);
and U10012 (N_10012,N_9747,N_9182);
or U10013 (N_10013,N_9191,N_9258);
nor U10014 (N_10014,N_9408,N_9125);
and U10015 (N_10015,N_9459,N_9166);
and U10016 (N_10016,N_9628,N_9146);
nand U10017 (N_10017,N_9257,N_9737);
or U10018 (N_10018,N_9621,N_9339);
and U10019 (N_10019,N_9385,N_9422);
or U10020 (N_10020,N_9359,N_9437);
nand U10021 (N_10021,N_9661,N_9565);
nor U10022 (N_10022,N_9270,N_9398);
nand U10023 (N_10023,N_9703,N_9411);
and U10024 (N_10024,N_9555,N_9225);
nor U10025 (N_10025,N_9283,N_9009);
nor U10026 (N_10026,N_9031,N_9355);
and U10027 (N_10027,N_9655,N_9576);
nor U10028 (N_10028,N_9424,N_9454);
nor U10029 (N_10029,N_9280,N_9641);
nor U10030 (N_10030,N_9604,N_9536);
or U10031 (N_10031,N_9418,N_9203);
nor U10032 (N_10032,N_9417,N_9269);
nand U10033 (N_10033,N_9579,N_9143);
nand U10034 (N_10034,N_9278,N_9419);
nand U10035 (N_10035,N_9190,N_9559);
nor U10036 (N_10036,N_9002,N_9590);
nand U10037 (N_10037,N_9731,N_9361);
nand U10038 (N_10038,N_9692,N_9626);
or U10039 (N_10039,N_9246,N_9624);
and U10040 (N_10040,N_9128,N_9444);
or U10041 (N_10041,N_9438,N_9322);
and U10042 (N_10042,N_9223,N_9072);
nand U10043 (N_10043,N_9148,N_9445);
and U10044 (N_10044,N_9616,N_9697);
and U10045 (N_10045,N_9676,N_9240);
or U10046 (N_10046,N_9487,N_9325);
nor U10047 (N_10047,N_9214,N_9499);
and U10048 (N_10048,N_9372,N_9373);
and U10049 (N_10049,N_9401,N_9707);
or U10050 (N_10050,N_9390,N_9274);
and U10051 (N_10051,N_9591,N_9250);
nand U10052 (N_10052,N_9281,N_9524);
nand U10053 (N_10053,N_9054,N_9446);
or U10054 (N_10054,N_9713,N_9421);
nand U10055 (N_10055,N_9465,N_9052);
or U10056 (N_10056,N_9436,N_9708);
or U10057 (N_10057,N_9575,N_9642);
and U10058 (N_10058,N_9026,N_9285);
or U10059 (N_10059,N_9558,N_9349);
xor U10060 (N_10060,N_9003,N_9358);
nand U10061 (N_10061,N_9122,N_9116);
nand U10062 (N_10062,N_9577,N_9120);
or U10063 (N_10063,N_9443,N_9220);
nor U10064 (N_10064,N_9290,N_9327);
and U10065 (N_10065,N_9381,N_9614);
and U10066 (N_10066,N_9048,N_9149);
nand U10067 (N_10067,N_9420,N_9075);
and U10068 (N_10068,N_9397,N_9478);
or U10069 (N_10069,N_9253,N_9047);
nor U10070 (N_10070,N_9141,N_9466);
and U10071 (N_10071,N_9007,N_9233);
nand U10072 (N_10072,N_9632,N_9308);
nor U10073 (N_10073,N_9540,N_9739);
or U10074 (N_10074,N_9660,N_9268);
nand U10075 (N_10075,N_9721,N_9286);
nand U10076 (N_10076,N_9333,N_9633);
and U10077 (N_10077,N_9212,N_9123);
and U10078 (N_10078,N_9046,N_9319);
nand U10079 (N_10079,N_9557,N_9549);
nand U10080 (N_10080,N_9021,N_9111);
or U10081 (N_10081,N_9071,N_9030);
nand U10082 (N_10082,N_9252,N_9526);
xor U10083 (N_10083,N_9589,N_9496);
and U10084 (N_10084,N_9547,N_9607);
nor U10085 (N_10085,N_9704,N_9627);
nor U10086 (N_10086,N_9188,N_9382);
or U10087 (N_10087,N_9095,N_9596);
and U10088 (N_10088,N_9060,N_9138);
and U10089 (N_10089,N_9096,N_9569);
and U10090 (N_10090,N_9468,N_9144);
nor U10091 (N_10091,N_9293,N_9516);
nand U10092 (N_10092,N_9717,N_9328);
and U10093 (N_10093,N_9011,N_9108);
nand U10094 (N_10094,N_9073,N_9165);
or U10095 (N_10095,N_9357,N_9277);
nand U10096 (N_10096,N_9505,N_9482);
nor U10097 (N_10097,N_9396,N_9230);
nand U10098 (N_10098,N_9131,N_9066);
or U10099 (N_10099,N_9543,N_9384);
or U10100 (N_10100,N_9728,N_9428);
or U10101 (N_10101,N_9251,N_9362);
and U10102 (N_10102,N_9107,N_9416);
nand U10103 (N_10103,N_9244,N_9699);
nor U10104 (N_10104,N_9666,N_9119);
nor U10105 (N_10105,N_9192,N_9651);
and U10106 (N_10106,N_9740,N_9467);
nand U10107 (N_10107,N_9414,N_9135);
and U10108 (N_10108,N_9427,N_9112);
or U10109 (N_10109,N_9599,N_9447);
or U10110 (N_10110,N_9136,N_9008);
and U10111 (N_10111,N_9133,N_9702);
nor U10112 (N_10112,N_9067,N_9659);
nand U10113 (N_10113,N_9151,N_9079);
nor U10114 (N_10114,N_9733,N_9648);
or U10115 (N_10115,N_9217,N_9534);
or U10116 (N_10116,N_9371,N_9249);
nand U10117 (N_10117,N_9612,N_9452);
and U10118 (N_10118,N_9043,N_9292);
and U10119 (N_10119,N_9369,N_9004);
or U10120 (N_10120,N_9492,N_9034);
xnor U10121 (N_10121,N_9087,N_9081);
nand U10122 (N_10122,N_9573,N_9683);
nand U10123 (N_10123,N_9080,N_9742);
nor U10124 (N_10124,N_9282,N_9479);
nand U10125 (N_10125,N_9619,N_9640);
nand U10126 (N_10126,N_9165,N_9110);
nor U10127 (N_10127,N_9415,N_9616);
or U10128 (N_10128,N_9352,N_9523);
and U10129 (N_10129,N_9456,N_9455);
or U10130 (N_10130,N_9328,N_9167);
nand U10131 (N_10131,N_9375,N_9033);
nor U10132 (N_10132,N_9402,N_9129);
and U10133 (N_10133,N_9498,N_9477);
nand U10134 (N_10134,N_9495,N_9592);
and U10135 (N_10135,N_9568,N_9602);
nor U10136 (N_10136,N_9557,N_9742);
and U10137 (N_10137,N_9040,N_9033);
nand U10138 (N_10138,N_9048,N_9125);
nor U10139 (N_10139,N_9568,N_9529);
and U10140 (N_10140,N_9500,N_9070);
and U10141 (N_10141,N_9104,N_9293);
nor U10142 (N_10142,N_9261,N_9185);
and U10143 (N_10143,N_9573,N_9382);
nor U10144 (N_10144,N_9126,N_9734);
nor U10145 (N_10145,N_9396,N_9537);
or U10146 (N_10146,N_9323,N_9339);
and U10147 (N_10147,N_9635,N_9424);
and U10148 (N_10148,N_9196,N_9199);
nor U10149 (N_10149,N_9623,N_9533);
nand U10150 (N_10150,N_9025,N_9499);
and U10151 (N_10151,N_9586,N_9094);
or U10152 (N_10152,N_9381,N_9676);
and U10153 (N_10153,N_9412,N_9406);
or U10154 (N_10154,N_9696,N_9581);
and U10155 (N_10155,N_9165,N_9307);
or U10156 (N_10156,N_9501,N_9160);
nor U10157 (N_10157,N_9438,N_9539);
nor U10158 (N_10158,N_9706,N_9203);
nor U10159 (N_10159,N_9568,N_9037);
and U10160 (N_10160,N_9092,N_9125);
and U10161 (N_10161,N_9040,N_9269);
xnor U10162 (N_10162,N_9208,N_9606);
nor U10163 (N_10163,N_9365,N_9140);
nor U10164 (N_10164,N_9356,N_9451);
or U10165 (N_10165,N_9122,N_9181);
nand U10166 (N_10166,N_9629,N_9049);
nor U10167 (N_10167,N_9032,N_9333);
or U10168 (N_10168,N_9666,N_9185);
and U10169 (N_10169,N_9106,N_9082);
or U10170 (N_10170,N_9519,N_9280);
or U10171 (N_10171,N_9058,N_9486);
nor U10172 (N_10172,N_9514,N_9511);
nand U10173 (N_10173,N_9367,N_9277);
nand U10174 (N_10174,N_9166,N_9746);
and U10175 (N_10175,N_9445,N_9660);
nor U10176 (N_10176,N_9214,N_9220);
or U10177 (N_10177,N_9691,N_9439);
nor U10178 (N_10178,N_9431,N_9282);
xor U10179 (N_10179,N_9241,N_9007);
nand U10180 (N_10180,N_9684,N_9216);
nor U10181 (N_10181,N_9266,N_9509);
nand U10182 (N_10182,N_9306,N_9274);
or U10183 (N_10183,N_9296,N_9319);
and U10184 (N_10184,N_9326,N_9570);
or U10185 (N_10185,N_9398,N_9464);
nor U10186 (N_10186,N_9120,N_9236);
nor U10187 (N_10187,N_9096,N_9514);
and U10188 (N_10188,N_9570,N_9186);
and U10189 (N_10189,N_9201,N_9724);
or U10190 (N_10190,N_9208,N_9615);
and U10191 (N_10191,N_9174,N_9339);
nor U10192 (N_10192,N_9627,N_9258);
or U10193 (N_10193,N_9419,N_9179);
nor U10194 (N_10194,N_9065,N_9323);
xnor U10195 (N_10195,N_9620,N_9207);
nor U10196 (N_10196,N_9332,N_9632);
or U10197 (N_10197,N_9734,N_9060);
and U10198 (N_10198,N_9421,N_9326);
xor U10199 (N_10199,N_9388,N_9302);
nand U10200 (N_10200,N_9393,N_9132);
nor U10201 (N_10201,N_9699,N_9694);
nor U10202 (N_10202,N_9337,N_9628);
and U10203 (N_10203,N_9631,N_9643);
or U10204 (N_10204,N_9712,N_9331);
nor U10205 (N_10205,N_9008,N_9607);
nor U10206 (N_10206,N_9351,N_9325);
nand U10207 (N_10207,N_9243,N_9092);
or U10208 (N_10208,N_9699,N_9107);
nor U10209 (N_10209,N_9256,N_9385);
nand U10210 (N_10210,N_9617,N_9199);
nor U10211 (N_10211,N_9499,N_9100);
or U10212 (N_10212,N_9537,N_9293);
and U10213 (N_10213,N_9184,N_9011);
nor U10214 (N_10214,N_9420,N_9216);
nor U10215 (N_10215,N_9252,N_9381);
and U10216 (N_10216,N_9739,N_9658);
or U10217 (N_10217,N_9276,N_9478);
nor U10218 (N_10218,N_9156,N_9385);
nand U10219 (N_10219,N_9240,N_9678);
nor U10220 (N_10220,N_9327,N_9444);
or U10221 (N_10221,N_9294,N_9115);
and U10222 (N_10222,N_9334,N_9255);
and U10223 (N_10223,N_9674,N_9366);
and U10224 (N_10224,N_9396,N_9472);
nor U10225 (N_10225,N_9477,N_9507);
nor U10226 (N_10226,N_9643,N_9257);
or U10227 (N_10227,N_9526,N_9215);
or U10228 (N_10228,N_9527,N_9533);
nand U10229 (N_10229,N_9231,N_9494);
nand U10230 (N_10230,N_9001,N_9574);
or U10231 (N_10231,N_9749,N_9181);
and U10232 (N_10232,N_9057,N_9427);
xnor U10233 (N_10233,N_9743,N_9441);
nor U10234 (N_10234,N_9091,N_9631);
nand U10235 (N_10235,N_9533,N_9725);
nor U10236 (N_10236,N_9236,N_9411);
nor U10237 (N_10237,N_9526,N_9490);
and U10238 (N_10238,N_9555,N_9070);
or U10239 (N_10239,N_9589,N_9051);
and U10240 (N_10240,N_9264,N_9283);
nand U10241 (N_10241,N_9196,N_9467);
xor U10242 (N_10242,N_9577,N_9314);
nand U10243 (N_10243,N_9293,N_9140);
nand U10244 (N_10244,N_9670,N_9533);
nand U10245 (N_10245,N_9308,N_9362);
nor U10246 (N_10246,N_9150,N_9149);
or U10247 (N_10247,N_9604,N_9134);
nand U10248 (N_10248,N_9222,N_9444);
nor U10249 (N_10249,N_9328,N_9376);
nand U10250 (N_10250,N_9544,N_9489);
and U10251 (N_10251,N_9707,N_9576);
nand U10252 (N_10252,N_9253,N_9570);
nand U10253 (N_10253,N_9031,N_9406);
nor U10254 (N_10254,N_9550,N_9241);
nand U10255 (N_10255,N_9487,N_9091);
nand U10256 (N_10256,N_9054,N_9628);
or U10257 (N_10257,N_9064,N_9155);
nand U10258 (N_10258,N_9494,N_9385);
nand U10259 (N_10259,N_9408,N_9356);
nand U10260 (N_10260,N_9233,N_9191);
and U10261 (N_10261,N_9685,N_9173);
nand U10262 (N_10262,N_9212,N_9420);
and U10263 (N_10263,N_9412,N_9540);
and U10264 (N_10264,N_9586,N_9531);
and U10265 (N_10265,N_9363,N_9653);
and U10266 (N_10266,N_9108,N_9328);
nand U10267 (N_10267,N_9683,N_9475);
or U10268 (N_10268,N_9184,N_9213);
and U10269 (N_10269,N_9621,N_9473);
nand U10270 (N_10270,N_9136,N_9086);
or U10271 (N_10271,N_9660,N_9080);
and U10272 (N_10272,N_9579,N_9667);
nor U10273 (N_10273,N_9277,N_9458);
nand U10274 (N_10274,N_9666,N_9487);
nor U10275 (N_10275,N_9543,N_9195);
and U10276 (N_10276,N_9152,N_9434);
nand U10277 (N_10277,N_9447,N_9100);
and U10278 (N_10278,N_9459,N_9369);
nand U10279 (N_10279,N_9380,N_9157);
and U10280 (N_10280,N_9660,N_9027);
nor U10281 (N_10281,N_9479,N_9263);
and U10282 (N_10282,N_9593,N_9530);
xor U10283 (N_10283,N_9149,N_9494);
nor U10284 (N_10284,N_9658,N_9586);
nor U10285 (N_10285,N_9140,N_9560);
xor U10286 (N_10286,N_9164,N_9694);
or U10287 (N_10287,N_9459,N_9207);
or U10288 (N_10288,N_9376,N_9024);
and U10289 (N_10289,N_9336,N_9032);
nand U10290 (N_10290,N_9669,N_9428);
or U10291 (N_10291,N_9269,N_9458);
or U10292 (N_10292,N_9196,N_9238);
nand U10293 (N_10293,N_9011,N_9042);
and U10294 (N_10294,N_9489,N_9318);
nor U10295 (N_10295,N_9645,N_9576);
nand U10296 (N_10296,N_9307,N_9724);
or U10297 (N_10297,N_9618,N_9653);
nand U10298 (N_10298,N_9111,N_9584);
and U10299 (N_10299,N_9162,N_9712);
or U10300 (N_10300,N_9627,N_9531);
or U10301 (N_10301,N_9201,N_9316);
nor U10302 (N_10302,N_9456,N_9398);
or U10303 (N_10303,N_9701,N_9369);
nor U10304 (N_10304,N_9497,N_9649);
xor U10305 (N_10305,N_9165,N_9707);
xor U10306 (N_10306,N_9167,N_9587);
nand U10307 (N_10307,N_9411,N_9654);
and U10308 (N_10308,N_9287,N_9723);
or U10309 (N_10309,N_9228,N_9520);
nand U10310 (N_10310,N_9328,N_9314);
and U10311 (N_10311,N_9022,N_9407);
nand U10312 (N_10312,N_9393,N_9143);
and U10313 (N_10313,N_9612,N_9466);
nor U10314 (N_10314,N_9192,N_9378);
xor U10315 (N_10315,N_9063,N_9337);
and U10316 (N_10316,N_9258,N_9738);
and U10317 (N_10317,N_9640,N_9546);
or U10318 (N_10318,N_9448,N_9525);
xor U10319 (N_10319,N_9630,N_9293);
or U10320 (N_10320,N_9583,N_9590);
nand U10321 (N_10321,N_9659,N_9090);
or U10322 (N_10322,N_9584,N_9318);
and U10323 (N_10323,N_9726,N_9380);
xor U10324 (N_10324,N_9676,N_9672);
and U10325 (N_10325,N_9474,N_9028);
nand U10326 (N_10326,N_9634,N_9295);
nand U10327 (N_10327,N_9690,N_9233);
nor U10328 (N_10328,N_9735,N_9676);
and U10329 (N_10329,N_9021,N_9084);
nand U10330 (N_10330,N_9170,N_9575);
and U10331 (N_10331,N_9521,N_9749);
and U10332 (N_10332,N_9076,N_9237);
and U10333 (N_10333,N_9446,N_9688);
and U10334 (N_10334,N_9082,N_9682);
and U10335 (N_10335,N_9279,N_9060);
nand U10336 (N_10336,N_9555,N_9619);
or U10337 (N_10337,N_9136,N_9569);
or U10338 (N_10338,N_9432,N_9705);
nor U10339 (N_10339,N_9381,N_9556);
nor U10340 (N_10340,N_9115,N_9320);
nand U10341 (N_10341,N_9048,N_9517);
nor U10342 (N_10342,N_9580,N_9052);
nor U10343 (N_10343,N_9479,N_9130);
nand U10344 (N_10344,N_9020,N_9630);
nor U10345 (N_10345,N_9572,N_9305);
and U10346 (N_10346,N_9024,N_9491);
nand U10347 (N_10347,N_9068,N_9502);
and U10348 (N_10348,N_9262,N_9260);
xnor U10349 (N_10349,N_9405,N_9312);
or U10350 (N_10350,N_9273,N_9636);
or U10351 (N_10351,N_9547,N_9582);
or U10352 (N_10352,N_9205,N_9700);
nand U10353 (N_10353,N_9068,N_9245);
nor U10354 (N_10354,N_9350,N_9074);
nand U10355 (N_10355,N_9669,N_9518);
nand U10356 (N_10356,N_9059,N_9690);
and U10357 (N_10357,N_9196,N_9230);
nor U10358 (N_10358,N_9701,N_9097);
and U10359 (N_10359,N_9072,N_9509);
or U10360 (N_10360,N_9213,N_9072);
and U10361 (N_10361,N_9595,N_9602);
nand U10362 (N_10362,N_9094,N_9743);
and U10363 (N_10363,N_9644,N_9384);
nor U10364 (N_10364,N_9402,N_9122);
xnor U10365 (N_10365,N_9737,N_9701);
nor U10366 (N_10366,N_9290,N_9579);
and U10367 (N_10367,N_9213,N_9294);
and U10368 (N_10368,N_9554,N_9714);
nor U10369 (N_10369,N_9588,N_9745);
nor U10370 (N_10370,N_9504,N_9276);
or U10371 (N_10371,N_9482,N_9120);
and U10372 (N_10372,N_9230,N_9739);
nor U10373 (N_10373,N_9584,N_9696);
and U10374 (N_10374,N_9159,N_9183);
or U10375 (N_10375,N_9389,N_9429);
nor U10376 (N_10376,N_9113,N_9015);
nand U10377 (N_10377,N_9601,N_9153);
and U10378 (N_10378,N_9418,N_9194);
and U10379 (N_10379,N_9587,N_9383);
nand U10380 (N_10380,N_9148,N_9517);
or U10381 (N_10381,N_9645,N_9051);
and U10382 (N_10382,N_9271,N_9524);
nand U10383 (N_10383,N_9487,N_9360);
and U10384 (N_10384,N_9035,N_9678);
nor U10385 (N_10385,N_9416,N_9544);
or U10386 (N_10386,N_9428,N_9296);
or U10387 (N_10387,N_9242,N_9256);
and U10388 (N_10388,N_9196,N_9337);
nor U10389 (N_10389,N_9127,N_9205);
and U10390 (N_10390,N_9698,N_9169);
nand U10391 (N_10391,N_9003,N_9324);
nand U10392 (N_10392,N_9247,N_9704);
or U10393 (N_10393,N_9082,N_9378);
or U10394 (N_10394,N_9262,N_9198);
and U10395 (N_10395,N_9304,N_9053);
or U10396 (N_10396,N_9611,N_9622);
nand U10397 (N_10397,N_9302,N_9320);
and U10398 (N_10398,N_9672,N_9550);
nand U10399 (N_10399,N_9645,N_9471);
nand U10400 (N_10400,N_9734,N_9376);
nand U10401 (N_10401,N_9686,N_9347);
or U10402 (N_10402,N_9091,N_9372);
and U10403 (N_10403,N_9418,N_9060);
or U10404 (N_10404,N_9428,N_9339);
nor U10405 (N_10405,N_9108,N_9053);
nand U10406 (N_10406,N_9528,N_9138);
and U10407 (N_10407,N_9105,N_9370);
nand U10408 (N_10408,N_9035,N_9647);
nor U10409 (N_10409,N_9469,N_9086);
and U10410 (N_10410,N_9633,N_9136);
or U10411 (N_10411,N_9097,N_9343);
and U10412 (N_10412,N_9485,N_9689);
nor U10413 (N_10413,N_9376,N_9112);
and U10414 (N_10414,N_9507,N_9314);
nand U10415 (N_10415,N_9741,N_9444);
nor U10416 (N_10416,N_9732,N_9157);
and U10417 (N_10417,N_9137,N_9080);
nor U10418 (N_10418,N_9558,N_9473);
xnor U10419 (N_10419,N_9473,N_9108);
nand U10420 (N_10420,N_9092,N_9644);
nand U10421 (N_10421,N_9683,N_9449);
or U10422 (N_10422,N_9181,N_9676);
nand U10423 (N_10423,N_9087,N_9328);
nor U10424 (N_10424,N_9558,N_9213);
or U10425 (N_10425,N_9278,N_9359);
nand U10426 (N_10426,N_9652,N_9259);
nor U10427 (N_10427,N_9693,N_9486);
nor U10428 (N_10428,N_9689,N_9281);
nor U10429 (N_10429,N_9165,N_9444);
nand U10430 (N_10430,N_9486,N_9316);
nand U10431 (N_10431,N_9121,N_9049);
nor U10432 (N_10432,N_9329,N_9429);
or U10433 (N_10433,N_9148,N_9170);
nand U10434 (N_10434,N_9547,N_9275);
nor U10435 (N_10435,N_9475,N_9721);
nand U10436 (N_10436,N_9563,N_9056);
nand U10437 (N_10437,N_9073,N_9522);
or U10438 (N_10438,N_9047,N_9114);
nor U10439 (N_10439,N_9076,N_9294);
or U10440 (N_10440,N_9719,N_9223);
or U10441 (N_10441,N_9172,N_9587);
and U10442 (N_10442,N_9449,N_9533);
nand U10443 (N_10443,N_9233,N_9627);
or U10444 (N_10444,N_9594,N_9528);
nand U10445 (N_10445,N_9616,N_9675);
nand U10446 (N_10446,N_9386,N_9497);
nand U10447 (N_10447,N_9479,N_9406);
nand U10448 (N_10448,N_9223,N_9452);
nand U10449 (N_10449,N_9250,N_9496);
or U10450 (N_10450,N_9381,N_9733);
nor U10451 (N_10451,N_9337,N_9542);
nor U10452 (N_10452,N_9474,N_9734);
nand U10453 (N_10453,N_9341,N_9085);
and U10454 (N_10454,N_9653,N_9392);
nor U10455 (N_10455,N_9030,N_9668);
nor U10456 (N_10456,N_9063,N_9143);
nor U10457 (N_10457,N_9699,N_9129);
nand U10458 (N_10458,N_9586,N_9156);
or U10459 (N_10459,N_9247,N_9725);
nand U10460 (N_10460,N_9620,N_9410);
nor U10461 (N_10461,N_9397,N_9539);
or U10462 (N_10462,N_9518,N_9637);
nor U10463 (N_10463,N_9089,N_9309);
and U10464 (N_10464,N_9376,N_9697);
and U10465 (N_10465,N_9011,N_9515);
or U10466 (N_10466,N_9130,N_9138);
and U10467 (N_10467,N_9607,N_9599);
nor U10468 (N_10468,N_9230,N_9619);
nand U10469 (N_10469,N_9425,N_9524);
or U10470 (N_10470,N_9358,N_9532);
nor U10471 (N_10471,N_9264,N_9597);
nor U10472 (N_10472,N_9062,N_9256);
or U10473 (N_10473,N_9252,N_9741);
nor U10474 (N_10474,N_9035,N_9541);
and U10475 (N_10475,N_9412,N_9594);
nor U10476 (N_10476,N_9213,N_9455);
nand U10477 (N_10477,N_9550,N_9381);
nand U10478 (N_10478,N_9492,N_9357);
nor U10479 (N_10479,N_9401,N_9654);
xnor U10480 (N_10480,N_9543,N_9290);
nand U10481 (N_10481,N_9591,N_9409);
or U10482 (N_10482,N_9461,N_9546);
and U10483 (N_10483,N_9236,N_9209);
and U10484 (N_10484,N_9370,N_9319);
nor U10485 (N_10485,N_9279,N_9364);
nand U10486 (N_10486,N_9681,N_9193);
nor U10487 (N_10487,N_9596,N_9249);
nand U10488 (N_10488,N_9706,N_9304);
nand U10489 (N_10489,N_9094,N_9315);
and U10490 (N_10490,N_9574,N_9356);
nand U10491 (N_10491,N_9175,N_9411);
or U10492 (N_10492,N_9567,N_9067);
and U10493 (N_10493,N_9135,N_9225);
or U10494 (N_10494,N_9528,N_9144);
nor U10495 (N_10495,N_9213,N_9134);
nand U10496 (N_10496,N_9720,N_9625);
and U10497 (N_10497,N_9581,N_9515);
and U10498 (N_10498,N_9404,N_9331);
or U10499 (N_10499,N_9017,N_9432);
or U10500 (N_10500,N_10039,N_10233);
or U10501 (N_10501,N_10330,N_9964);
nor U10502 (N_10502,N_10161,N_10055);
or U10503 (N_10503,N_10130,N_10222);
and U10504 (N_10504,N_9775,N_10072);
nor U10505 (N_10505,N_10144,N_10289);
or U10506 (N_10506,N_10250,N_9910);
nand U10507 (N_10507,N_10044,N_10187);
nor U10508 (N_10508,N_10420,N_10362);
nand U10509 (N_10509,N_9876,N_9934);
and U10510 (N_10510,N_10481,N_10297);
and U10511 (N_10511,N_10283,N_10263);
xnor U10512 (N_10512,N_9947,N_10131);
and U10513 (N_10513,N_9965,N_10338);
nor U10514 (N_10514,N_10142,N_10327);
and U10515 (N_10515,N_9782,N_10436);
or U10516 (N_10516,N_10141,N_10412);
nand U10517 (N_10517,N_10337,N_10326);
nor U10518 (N_10518,N_10227,N_10203);
and U10519 (N_10519,N_9764,N_10117);
or U10520 (N_10520,N_10170,N_9878);
nor U10521 (N_10521,N_10288,N_9954);
and U10522 (N_10522,N_10462,N_10185);
or U10523 (N_10523,N_10410,N_10450);
xor U10524 (N_10524,N_9919,N_9872);
and U10525 (N_10525,N_9995,N_9950);
and U10526 (N_10526,N_9756,N_10220);
nand U10527 (N_10527,N_10177,N_9786);
xor U10528 (N_10528,N_10427,N_10439);
nand U10529 (N_10529,N_10484,N_10228);
nor U10530 (N_10530,N_9843,N_10319);
and U10531 (N_10531,N_10242,N_9999);
nand U10532 (N_10532,N_10385,N_10376);
or U10533 (N_10533,N_10490,N_9864);
nor U10534 (N_10534,N_10425,N_10102);
nor U10535 (N_10535,N_10200,N_10322);
and U10536 (N_10536,N_10422,N_10060);
nor U10537 (N_10537,N_9927,N_10247);
and U10538 (N_10538,N_10107,N_9766);
or U10539 (N_10539,N_9821,N_10051);
nor U10540 (N_10540,N_10248,N_10184);
nand U10541 (N_10541,N_9856,N_10007);
nand U10542 (N_10542,N_10380,N_10041);
or U10543 (N_10543,N_10480,N_10014);
nand U10544 (N_10544,N_9789,N_10026);
or U10545 (N_10545,N_10443,N_10042);
and U10546 (N_10546,N_10004,N_10334);
nand U10547 (N_10547,N_10206,N_10295);
nor U10548 (N_10548,N_10179,N_10333);
nand U10549 (N_10549,N_10017,N_10011);
nand U10550 (N_10550,N_10374,N_9905);
nand U10551 (N_10551,N_10080,N_9848);
nand U10552 (N_10552,N_9914,N_10127);
nor U10553 (N_10553,N_9893,N_10448);
and U10554 (N_10554,N_9917,N_9968);
nand U10555 (N_10555,N_9790,N_9819);
and U10556 (N_10556,N_10037,N_9851);
nor U10557 (N_10557,N_10082,N_10109);
nand U10558 (N_10558,N_9904,N_10471);
nand U10559 (N_10559,N_10251,N_10067);
nor U10560 (N_10560,N_10128,N_10482);
and U10561 (N_10561,N_10205,N_10465);
nand U10562 (N_10562,N_9956,N_9976);
nand U10563 (N_10563,N_10252,N_10043);
nand U10564 (N_10564,N_10164,N_10071);
nand U10565 (N_10565,N_9994,N_9831);
or U10566 (N_10566,N_10045,N_9929);
or U10567 (N_10567,N_9804,N_10214);
nand U10568 (N_10568,N_9885,N_10027);
and U10569 (N_10569,N_9977,N_10174);
nand U10570 (N_10570,N_9901,N_9953);
nand U10571 (N_10571,N_10191,N_10488);
or U10572 (N_10572,N_10114,N_9774);
nand U10573 (N_10573,N_10403,N_10497);
and U10574 (N_10574,N_9912,N_9907);
nor U10575 (N_10575,N_9900,N_10413);
or U10576 (N_10576,N_10172,N_10305);
and U10577 (N_10577,N_10238,N_10118);
and U10578 (N_10578,N_10453,N_10303);
or U10579 (N_10579,N_9902,N_10466);
xnor U10580 (N_10580,N_10441,N_10260);
and U10581 (N_10581,N_10301,N_10230);
nor U10582 (N_10582,N_10181,N_10286);
or U10583 (N_10583,N_10396,N_9897);
nor U10584 (N_10584,N_9842,N_10224);
or U10585 (N_10585,N_10212,N_10394);
nand U10586 (N_10586,N_10423,N_10197);
nand U10587 (N_10587,N_10216,N_10239);
and U10588 (N_10588,N_10409,N_10491);
nor U10589 (N_10589,N_9866,N_10078);
and U10590 (N_10590,N_9762,N_10135);
or U10591 (N_10591,N_10133,N_10195);
nand U10592 (N_10592,N_10243,N_9996);
nor U10593 (N_10593,N_10266,N_10094);
and U10594 (N_10594,N_10419,N_10373);
nand U10595 (N_10595,N_9936,N_10321);
nand U10596 (N_10596,N_9845,N_10277);
or U10597 (N_10597,N_9757,N_9779);
xor U10598 (N_10598,N_10032,N_9908);
nand U10599 (N_10599,N_10038,N_10134);
nor U10600 (N_10600,N_10271,N_10324);
xnor U10601 (N_10601,N_9861,N_10311);
or U10602 (N_10602,N_10495,N_10244);
nor U10603 (N_10603,N_10414,N_10132);
nand U10604 (N_10604,N_10178,N_10445);
or U10605 (N_10605,N_10147,N_10265);
nor U10606 (N_10606,N_10235,N_9807);
nand U10607 (N_10607,N_10168,N_9922);
nand U10608 (N_10608,N_10366,N_10281);
or U10609 (N_10609,N_10342,N_10329);
or U10610 (N_10610,N_10034,N_10010);
or U10611 (N_10611,N_10404,N_10282);
xnor U10612 (N_10612,N_9846,N_9990);
nor U10613 (N_10613,N_10309,N_10369);
and U10614 (N_10614,N_10213,N_10189);
or U10615 (N_10615,N_10347,N_10077);
nand U10616 (N_10616,N_10395,N_9798);
nand U10617 (N_10617,N_10461,N_10218);
nand U10618 (N_10618,N_10307,N_9805);
nand U10619 (N_10619,N_10320,N_10318);
and U10620 (N_10620,N_10121,N_10084);
or U10621 (N_10621,N_9773,N_10090);
nand U10622 (N_10622,N_10151,N_9791);
xnor U10623 (N_10623,N_10472,N_10270);
and U10624 (N_10624,N_10036,N_10021);
or U10625 (N_10625,N_10204,N_10440);
or U10626 (N_10626,N_9788,N_10015);
nand U10627 (N_10627,N_9759,N_10175);
or U10628 (N_10628,N_9802,N_9760);
xor U10629 (N_10629,N_10098,N_9752);
nor U10630 (N_10630,N_9800,N_10198);
nand U10631 (N_10631,N_10328,N_10360);
or U10632 (N_10632,N_9827,N_10101);
nor U10633 (N_10633,N_9924,N_10361);
nand U10634 (N_10634,N_10159,N_10381);
or U10635 (N_10635,N_10095,N_10378);
or U10636 (N_10636,N_10382,N_10160);
nand U10637 (N_10637,N_10406,N_9986);
nor U10638 (N_10638,N_9824,N_9911);
nor U10639 (N_10639,N_10207,N_10291);
and U10640 (N_10640,N_10304,N_9808);
nand U10641 (N_10641,N_10083,N_10379);
or U10642 (N_10642,N_10353,N_9892);
nand U10643 (N_10643,N_10188,N_10029);
or U10644 (N_10644,N_10163,N_10140);
nor U10645 (N_10645,N_10389,N_10199);
nand U10646 (N_10646,N_10494,N_10240);
and U10647 (N_10647,N_10006,N_9888);
nor U10648 (N_10648,N_10125,N_10498);
nor U10649 (N_10649,N_10097,N_10371);
xnor U10650 (N_10650,N_9817,N_9873);
nand U10651 (N_10651,N_10398,N_9753);
nand U10652 (N_10652,N_9833,N_10033);
nor U10653 (N_10653,N_9795,N_10193);
or U10654 (N_10654,N_10202,N_10210);
nor U10655 (N_10655,N_10272,N_9896);
or U10656 (N_10656,N_9992,N_9915);
nand U10657 (N_10657,N_10345,N_9889);
or U10658 (N_10658,N_10446,N_10234);
and U10659 (N_10659,N_9942,N_10152);
nand U10660 (N_10660,N_10129,N_9793);
nor U10661 (N_10661,N_10299,N_9899);
nand U10662 (N_10662,N_10390,N_9871);
and U10663 (N_10663,N_10028,N_10232);
or U10664 (N_10664,N_9830,N_9799);
nand U10665 (N_10665,N_10368,N_9792);
nor U10666 (N_10666,N_10183,N_9993);
or U10667 (N_10667,N_10499,N_9933);
nand U10668 (N_10668,N_10259,N_9973);
nand U10669 (N_10669,N_10306,N_10162);
or U10670 (N_10670,N_9928,N_10449);
and U10671 (N_10671,N_10100,N_10110);
and U10672 (N_10672,N_10346,N_9837);
nor U10673 (N_10673,N_9847,N_10377);
or U10674 (N_10674,N_10428,N_10349);
nor U10675 (N_10675,N_10351,N_10287);
nor U10676 (N_10676,N_10386,N_9923);
nand U10677 (N_10677,N_10167,N_9849);
and U10678 (N_10678,N_10253,N_10312);
and U10679 (N_10679,N_10292,N_9988);
or U10680 (N_10680,N_10363,N_10262);
or U10681 (N_10681,N_9980,N_10261);
or U10682 (N_10682,N_10256,N_10106);
or U10683 (N_10683,N_10226,N_9940);
and U10684 (N_10684,N_10217,N_10065);
or U10685 (N_10685,N_10447,N_10056);
nor U10686 (N_10686,N_10241,N_9841);
or U10687 (N_10687,N_10331,N_10358);
nor U10688 (N_10688,N_10444,N_9879);
or U10689 (N_10689,N_10364,N_10057);
nor U10690 (N_10690,N_10076,N_9826);
or U10691 (N_10691,N_10339,N_10470);
or U10692 (N_10692,N_10054,N_10122);
or U10693 (N_10693,N_10171,N_9981);
nor U10694 (N_10694,N_10356,N_10108);
or U10695 (N_10695,N_10387,N_9882);
and U10696 (N_10696,N_10005,N_10008);
nand U10697 (N_10697,N_10023,N_10040);
or U10698 (N_10698,N_10343,N_10479);
and U10699 (N_10699,N_9991,N_10392);
nor U10700 (N_10700,N_10267,N_9772);
nand U10701 (N_10701,N_10116,N_10370);
and U10702 (N_10702,N_10492,N_9967);
nor U10703 (N_10703,N_10279,N_9972);
nor U10704 (N_10704,N_10400,N_10048);
nor U10705 (N_10705,N_9769,N_9906);
nor U10706 (N_10706,N_10158,N_10405);
and U10707 (N_10707,N_10111,N_10437);
nor U10708 (N_10708,N_9877,N_10079);
nor U10709 (N_10709,N_10173,N_10457);
or U10710 (N_10710,N_10201,N_10073);
nand U10711 (N_10711,N_9870,N_9839);
nand U10712 (N_10712,N_9765,N_10464);
nor U10713 (N_10713,N_10085,N_9803);
or U10714 (N_10714,N_10478,N_10146);
and U10715 (N_10715,N_10000,N_10391);
and U10716 (N_10716,N_9894,N_10460);
and U10717 (N_10717,N_10483,N_9858);
or U10718 (N_10718,N_10154,N_9943);
nand U10719 (N_10719,N_10186,N_10407);
nor U10720 (N_10720,N_10225,N_10431);
nor U10721 (N_10721,N_10003,N_10317);
nand U10722 (N_10722,N_10126,N_10138);
and U10723 (N_10723,N_9838,N_10139);
nand U10724 (N_10724,N_9780,N_10426);
nor U10725 (N_10725,N_10310,N_9931);
or U10726 (N_10726,N_10383,N_10325);
nand U10727 (N_10727,N_10352,N_10119);
nand U10728 (N_10728,N_9859,N_10236);
nor U10729 (N_10729,N_10257,N_10009);
nor U10730 (N_10730,N_9771,N_9794);
and U10731 (N_10731,N_9875,N_10416);
nor U10732 (N_10732,N_9758,N_10113);
and U10733 (N_10733,N_10302,N_9835);
and U10734 (N_10734,N_9806,N_9958);
nor U10735 (N_10735,N_10375,N_10344);
nor U10736 (N_10736,N_9913,N_10268);
nand U10737 (N_10737,N_10269,N_10166);
nand U10738 (N_10738,N_10046,N_10081);
and U10739 (N_10739,N_10357,N_10180);
or U10740 (N_10740,N_9939,N_10105);
or U10741 (N_10741,N_9959,N_10053);
nor U10742 (N_10742,N_10208,N_9937);
nor U10743 (N_10743,N_9770,N_10096);
nor U10744 (N_10744,N_10157,N_10255);
nor U10745 (N_10745,N_9969,N_10399);
and U10746 (N_10746,N_10229,N_10274);
nor U10747 (N_10747,N_10355,N_10231);
or U10748 (N_10748,N_10456,N_9853);
and U10749 (N_10749,N_10402,N_10264);
nand U10750 (N_10750,N_9935,N_9857);
and U10751 (N_10751,N_9868,N_9974);
or U10752 (N_10752,N_9829,N_10424);
or U10753 (N_10753,N_10475,N_10074);
nand U10754 (N_10754,N_9865,N_9997);
nand U10755 (N_10755,N_10156,N_9920);
and U10756 (N_10756,N_10052,N_10112);
or U10757 (N_10757,N_9979,N_9984);
and U10758 (N_10758,N_10432,N_10058);
or U10759 (N_10759,N_9815,N_10278);
and U10760 (N_10760,N_10031,N_10417);
nand U10761 (N_10761,N_9822,N_10254);
or U10762 (N_10762,N_10332,N_9989);
or U10763 (N_10763,N_10182,N_9796);
and U10764 (N_10764,N_10245,N_10050);
nand U10765 (N_10765,N_10150,N_10315);
and U10766 (N_10766,N_10223,N_10463);
or U10767 (N_10767,N_9982,N_10314);
nor U10768 (N_10768,N_10165,N_9916);
or U10769 (N_10769,N_9891,N_10438);
nor U10770 (N_10770,N_9895,N_10473);
and U10771 (N_10771,N_10022,N_10468);
xnor U10772 (N_10772,N_10487,N_10384);
xnor U10773 (N_10773,N_9811,N_9962);
and U10774 (N_10774,N_9761,N_10194);
nand U10775 (N_10775,N_10341,N_10421);
and U10776 (N_10776,N_9961,N_10155);
nor U10777 (N_10777,N_9820,N_10249);
nand U10778 (N_10778,N_10469,N_9886);
nor U10779 (N_10779,N_9787,N_10418);
nand U10780 (N_10780,N_9971,N_9925);
nor U10781 (N_10781,N_10354,N_10476);
nand U10782 (N_10782,N_10308,N_9813);
and U10783 (N_10783,N_10365,N_10275);
and U10784 (N_10784,N_10123,N_10002);
or U10785 (N_10785,N_9887,N_9784);
or U10786 (N_10786,N_9755,N_10474);
and U10787 (N_10787,N_10061,N_10024);
and U10788 (N_10788,N_10086,N_10049);
nand U10789 (N_10789,N_9941,N_9785);
and U10790 (N_10790,N_9987,N_10429);
nor U10791 (N_10791,N_9998,N_10196);
nor U10792 (N_10792,N_9754,N_10455);
or U10793 (N_10793,N_10452,N_9921);
or U10794 (N_10794,N_10276,N_10401);
nand U10795 (N_10795,N_10493,N_9855);
nand U10796 (N_10796,N_10093,N_10066);
nand U10797 (N_10797,N_9809,N_10190);
nor U10798 (N_10798,N_10388,N_10246);
nand U10799 (N_10799,N_9944,N_10063);
nor U10800 (N_10800,N_9867,N_9903);
nor U10801 (N_10801,N_9966,N_10068);
or U10802 (N_10802,N_10103,N_10415);
and U10803 (N_10803,N_10298,N_9883);
and U10804 (N_10804,N_10316,N_10408);
and U10805 (N_10805,N_10176,N_10451);
and U10806 (N_10806,N_10300,N_10348);
or U10807 (N_10807,N_10284,N_9862);
nor U10808 (N_10808,N_9960,N_10433);
nand U10809 (N_10809,N_10013,N_10059);
or U10810 (N_10810,N_9975,N_10273);
and U10811 (N_10811,N_9881,N_9832);
and U10812 (N_10812,N_9930,N_10359);
and U10813 (N_10813,N_10153,N_9874);
and U10814 (N_10814,N_10237,N_9834);
nand U10815 (N_10815,N_9777,N_10459);
or U10816 (N_10816,N_10454,N_9863);
nor U10817 (N_10817,N_10221,N_10477);
and U10818 (N_10818,N_10169,N_9970);
and U10819 (N_10819,N_10442,N_10149);
and U10820 (N_10820,N_9840,N_10215);
or U10821 (N_10821,N_9890,N_10104);
nand U10822 (N_10822,N_10335,N_10020);
nor U10823 (N_10823,N_9767,N_10018);
or U10824 (N_10824,N_10016,N_9869);
nor U10825 (N_10825,N_9884,N_9951);
and U10826 (N_10826,N_9778,N_10137);
nor U10827 (N_10827,N_9818,N_10088);
nand U10828 (N_10828,N_10099,N_10496);
nand U10829 (N_10829,N_10489,N_10136);
nand U10830 (N_10830,N_10458,N_10062);
nor U10831 (N_10831,N_10120,N_9825);
nand U10832 (N_10832,N_9781,N_10030);
or U10833 (N_10833,N_9926,N_10296);
and U10834 (N_10834,N_9750,N_10115);
nand U10835 (N_10835,N_10293,N_10285);
and U10836 (N_10836,N_10350,N_9932);
nor U10837 (N_10837,N_10047,N_10075);
or U10838 (N_10838,N_10323,N_10430);
or U10839 (N_10839,N_9955,N_10397);
and U10840 (N_10840,N_10025,N_9836);
nand U10841 (N_10841,N_10294,N_9814);
or U10842 (N_10842,N_9810,N_9823);
or U10843 (N_10843,N_9828,N_10411);
and U10844 (N_10844,N_10435,N_10340);
or U10845 (N_10845,N_9957,N_10209);
or U10846 (N_10846,N_10087,N_9797);
or U10847 (N_10847,N_9948,N_10486);
xnor U10848 (N_10848,N_9898,N_9946);
xnor U10849 (N_10849,N_10393,N_9880);
nor U10850 (N_10850,N_9918,N_9963);
nor U10851 (N_10851,N_10258,N_9776);
or U10852 (N_10852,N_9949,N_10434);
and U10853 (N_10853,N_10001,N_10092);
nand U10854 (N_10854,N_10290,N_10035);
or U10855 (N_10855,N_10485,N_10372);
nand U10856 (N_10856,N_9978,N_9983);
nand U10857 (N_10857,N_9768,N_9909);
and U10858 (N_10858,N_10211,N_9816);
and U10859 (N_10859,N_10012,N_10148);
and U10860 (N_10860,N_9854,N_10336);
and U10861 (N_10861,N_9945,N_9844);
nand U10862 (N_10862,N_9850,N_10467);
xor U10863 (N_10863,N_10143,N_9751);
nand U10864 (N_10864,N_9763,N_9852);
and U10865 (N_10865,N_9783,N_10089);
or U10866 (N_10866,N_10070,N_10069);
and U10867 (N_10867,N_9952,N_10124);
and U10868 (N_10868,N_9860,N_10091);
nand U10869 (N_10869,N_10145,N_10192);
or U10870 (N_10870,N_9985,N_10219);
nand U10871 (N_10871,N_10367,N_9938);
or U10872 (N_10872,N_10313,N_10064);
nand U10873 (N_10873,N_9812,N_10280);
and U10874 (N_10874,N_10019,N_9801);
and U10875 (N_10875,N_9884,N_10481);
xnor U10876 (N_10876,N_10355,N_10396);
nor U10877 (N_10877,N_10088,N_9760);
nor U10878 (N_10878,N_9943,N_10103);
nor U10879 (N_10879,N_10070,N_10169);
nand U10880 (N_10880,N_10098,N_10246);
and U10881 (N_10881,N_10434,N_9775);
nand U10882 (N_10882,N_9967,N_10161);
and U10883 (N_10883,N_10156,N_9786);
nand U10884 (N_10884,N_10382,N_10471);
or U10885 (N_10885,N_10119,N_10045);
and U10886 (N_10886,N_9768,N_10034);
or U10887 (N_10887,N_9926,N_10354);
and U10888 (N_10888,N_10194,N_10311);
or U10889 (N_10889,N_10269,N_9903);
or U10890 (N_10890,N_10195,N_10339);
or U10891 (N_10891,N_10413,N_9981);
and U10892 (N_10892,N_10256,N_10207);
nor U10893 (N_10893,N_10410,N_10115);
nand U10894 (N_10894,N_10385,N_10003);
nand U10895 (N_10895,N_10431,N_10163);
nor U10896 (N_10896,N_10432,N_10001);
nand U10897 (N_10897,N_10000,N_9761);
nor U10898 (N_10898,N_9958,N_10012);
or U10899 (N_10899,N_10479,N_9940);
or U10900 (N_10900,N_10262,N_9798);
or U10901 (N_10901,N_10032,N_10453);
or U10902 (N_10902,N_10332,N_10084);
nor U10903 (N_10903,N_10184,N_10448);
or U10904 (N_10904,N_10269,N_10080);
and U10905 (N_10905,N_10389,N_10236);
nor U10906 (N_10906,N_9816,N_10094);
nor U10907 (N_10907,N_9954,N_10364);
and U10908 (N_10908,N_10022,N_10289);
and U10909 (N_10909,N_10023,N_10082);
nor U10910 (N_10910,N_10439,N_10324);
nand U10911 (N_10911,N_10047,N_10345);
nor U10912 (N_10912,N_10128,N_9861);
and U10913 (N_10913,N_9849,N_9810);
or U10914 (N_10914,N_9796,N_9813);
and U10915 (N_10915,N_10480,N_10108);
nor U10916 (N_10916,N_9839,N_9791);
and U10917 (N_10917,N_10091,N_9993);
nor U10918 (N_10918,N_10461,N_9947);
nor U10919 (N_10919,N_10390,N_10490);
nor U10920 (N_10920,N_10102,N_10139);
nand U10921 (N_10921,N_10032,N_10498);
or U10922 (N_10922,N_9882,N_10307);
nor U10923 (N_10923,N_10011,N_10393);
and U10924 (N_10924,N_10354,N_10376);
or U10925 (N_10925,N_9756,N_10204);
nor U10926 (N_10926,N_10124,N_10178);
or U10927 (N_10927,N_10160,N_10263);
nor U10928 (N_10928,N_10004,N_10101);
nand U10929 (N_10929,N_9869,N_10217);
nand U10930 (N_10930,N_9754,N_10114);
and U10931 (N_10931,N_9777,N_9816);
nor U10932 (N_10932,N_9774,N_9808);
and U10933 (N_10933,N_10123,N_9849);
nor U10934 (N_10934,N_10248,N_9863);
nor U10935 (N_10935,N_9964,N_9827);
nand U10936 (N_10936,N_10085,N_10350);
or U10937 (N_10937,N_10441,N_10408);
xor U10938 (N_10938,N_10472,N_10495);
nor U10939 (N_10939,N_10465,N_10209);
nor U10940 (N_10940,N_10167,N_9926);
and U10941 (N_10941,N_9953,N_9812);
and U10942 (N_10942,N_9751,N_10379);
nor U10943 (N_10943,N_10094,N_10384);
nand U10944 (N_10944,N_10331,N_9797);
nand U10945 (N_10945,N_9799,N_9798);
nand U10946 (N_10946,N_9772,N_10065);
nand U10947 (N_10947,N_10353,N_9849);
nand U10948 (N_10948,N_10121,N_10450);
or U10949 (N_10949,N_10492,N_9848);
or U10950 (N_10950,N_9823,N_9797);
nand U10951 (N_10951,N_9785,N_9767);
nand U10952 (N_10952,N_9929,N_10355);
and U10953 (N_10953,N_10381,N_10499);
or U10954 (N_10954,N_10139,N_10437);
nand U10955 (N_10955,N_10478,N_10411);
or U10956 (N_10956,N_9823,N_10208);
or U10957 (N_10957,N_9765,N_10149);
nor U10958 (N_10958,N_10276,N_10024);
or U10959 (N_10959,N_10129,N_10034);
nand U10960 (N_10960,N_10130,N_10266);
and U10961 (N_10961,N_10181,N_10075);
nand U10962 (N_10962,N_10125,N_10055);
nor U10963 (N_10963,N_10361,N_9838);
nand U10964 (N_10964,N_10273,N_10290);
or U10965 (N_10965,N_10141,N_10205);
xnor U10966 (N_10966,N_10462,N_10452);
or U10967 (N_10967,N_10167,N_10170);
nand U10968 (N_10968,N_9764,N_10499);
nand U10969 (N_10969,N_10124,N_10101);
and U10970 (N_10970,N_10042,N_9965);
and U10971 (N_10971,N_9855,N_10413);
or U10972 (N_10972,N_9777,N_10187);
nand U10973 (N_10973,N_10042,N_10019);
or U10974 (N_10974,N_10335,N_10374);
or U10975 (N_10975,N_10473,N_10181);
and U10976 (N_10976,N_10258,N_9987);
nor U10977 (N_10977,N_10472,N_9828);
nor U10978 (N_10978,N_9983,N_10252);
nand U10979 (N_10979,N_9841,N_9852);
nand U10980 (N_10980,N_10469,N_9829);
and U10981 (N_10981,N_9968,N_10070);
nor U10982 (N_10982,N_10123,N_10290);
nand U10983 (N_10983,N_9909,N_9883);
or U10984 (N_10984,N_10203,N_10109);
and U10985 (N_10985,N_10426,N_9968);
nor U10986 (N_10986,N_10241,N_10109);
nor U10987 (N_10987,N_10193,N_9883);
and U10988 (N_10988,N_9888,N_9787);
nand U10989 (N_10989,N_10125,N_10402);
nor U10990 (N_10990,N_10321,N_10240);
nand U10991 (N_10991,N_9864,N_9842);
nor U10992 (N_10992,N_10085,N_10063);
xnor U10993 (N_10993,N_9828,N_10407);
nand U10994 (N_10994,N_10315,N_10117);
and U10995 (N_10995,N_10236,N_10449);
or U10996 (N_10996,N_9773,N_10072);
or U10997 (N_10997,N_10423,N_10312);
nand U10998 (N_10998,N_9776,N_10192);
nor U10999 (N_10999,N_10193,N_9876);
nor U11000 (N_11000,N_9861,N_10331);
nand U11001 (N_11001,N_10446,N_10353);
or U11002 (N_11002,N_9970,N_9781);
or U11003 (N_11003,N_10270,N_9866);
or U11004 (N_11004,N_10449,N_10440);
nor U11005 (N_11005,N_9872,N_9827);
and U11006 (N_11006,N_9758,N_9813);
nand U11007 (N_11007,N_9860,N_9968);
nor U11008 (N_11008,N_10229,N_10030);
nand U11009 (N_11009,N_9920,N_10229);
nor U11010 (N_11010,N_10381,N_10490);
and U11011 (N_11011,N_10419,N_9915);
or U11012 (N_11012,N_10440,N_10036);
nand U11013 (N_11013,N_10203,N_10202);
and U11014 (N_11014,N_10143,N_10091);
nand U11015 (N_11015,N_10366,N_10018);
and U11016 (N_11016,N_10012,N_9765);
xnor U11017 (N_11017,N_10485,N_10203);
or U11018 (N_11018,N_10090,N_10145);
nor U11019 (N_11019,N_9960,N_9781);
or U11020 (N_11020,N_9792,N_9805);
and U11021 (N_11021,N_10138,N_10311);
nor U11022 (N_11022,N_9884,N_9825);
and U11023 (N_11023,N_9881,N_9782);
and U11024 (N_11024,N_10004,N_10225);
and U11025 (N_11025,N_10258,N_10404);
nor U11026 (N_11026,N_10273,N_10499);
nor U11027 (N_11027,N_9962,N_10321);
and U11028 (N_11028,N_10254,N_10259);
or U11029 (N_11029,N_9943,N_9760);
nand U11030 (N_11030,N_10134,N_9868);
or U11031 (N_11031,N_10473,N_9764);
and U11032 (N_11032,N_10404,N_10154);
nand U11033 (N_11033,N_10089,N_10080);
or U11034 (N_11034,N_10151,N_9777);
nor U11035 (N_11035,N_10362,N_9753);
and U11036 (N_11036,N_10089,N_10024);
or U11037 (N_11037,N_10318,N_10471);
and U11038 (N_11038,N_9926,N_10316);
nor U11039 (N_11039,N_10093,N_10329);
nor U11040 (N_11040,N_10083,N_10322);
nand U11041 (N_11041,N_10490,N_9931);
or U11042 (N_11042,N_9978,N_9998);
or U11043 (N_11043,N_10148,N_10168);
nand U11044 (N_11044,N_10179,N_10287);
nand U11045 (N_11045,N_10232,N_10426);
nand U11046 (N_11046,N_10233,N_10092);
xor U11047 (N_11047,N_10344,N_10430);
or U11048 (N_11048,N_10029,N_10226);
nand U11049 (N_11049,N_10317,N_10400);
nand U11050 (N_11050,N_10306,N_10407);
or U11051 (N_11051,N_10252,N_9955);
or U11052 (N_11052,N_10145,N_9756);
and U11053 (N_11053,N_10246,N_9859);
and U11054 (N_11054,N_9950,N_10295);
or U11055 (N_11055,N_10490,N_9873);
nand U11056 (N_11056,N_10167,N_10047);
xor U11057 (N_11057,N_10075,N_10084);
or U11058 (N_11058,N_10330,N_10411);
or U11059 (N_11059,N_10263,N_9979);
or U11060 (N_11060,N_10410,N_10475);
and U11061 (N_11061,N_10221,N_9976);
and U11062 (N_11062,N_10480,N_9750);
nand U11063 (N_11063,N_9960,N_9993);
nand U11064 (N_11064,N_10358,N_10285);
or U11065 (N_11065,N_10239,N_10463);
nand U11066 (N_11066,N_10016,N_9771);
or U11067 (N_11067,N_10193,N_10361);
nand U11068 (N_11068,N_9807,N_10356);
and U11069 (N_11069,N_10244,N_10257);
nor U11070 (N_11070,N_9772,N_10339);
nand U11071 (N_11071,N_10290,N_10241);
nor U11072 (N_11072,N_10241,N_10161);
nor U11073 (N_11073,N_10001,N_10252);
or U11074 (N_11074,N_10282,N_10197);
or U11075 (N_11075,N_9782,N_10134);
nand U11076 (N_11076,N_10065,N_9993);
and U11077 (N_11077,N_10260,N_10401);
nor U11078 (N_11078,N_10342,N_9780);
nand U11079 (N_11079,N_10004,N_10177);
or U11080 (N_11080,N_9881,N_10132);
nor U11081 (N_11081,N_9915,N_10145);
or U11082 (N_11082,N_10220,N_9752);
xor U11083 (N_11083,N_9851,N_10122);
nand U11084 (N_11084,N_10405,N_10477);
nor U11085 (N_11085,N_10208,N_10252);
nand U11086 (N_11086,N_10006,N_10345);
nand U11087 (N_11087,N_9884,N_10356);
nand U11088 (N_11088,N_10226,N_10319);
and U11089 (N_11089,N_10137,N_10186);
nand U11090 (N_11090,N_10084,N_9969);
or U11091 (N_11091,N_9928,N_10271);
nor U11092 (N_11092,N_9953,N_10171);
and U11093 (N_11093,N_9990,N_9791);
nor U11094 (N_11094,N_10402,N_9903);
or U11095 (N_11095,N_9897,N_10412);
or U11096 (N_11096,N_10443,N_10069);
nand U11097 (N_11097,N_10281,N_9864);
xnor U11098 (N_11098,N_10422,N_10363);
nand U11099 (N_11099,N_10263,N_10421);
nor U11100 (N_11100,N_10133,N_10417);
and U11101 (N_11101,N_10480,N_10195);
and U11102 (N_11102,N_10412,N_9856);
nand U11103 (N_11103,N_10158,N_10482);
nand U11104 (N_11104,N_10455,N_10040);
nor U11105 (N_11105,N_10372,N_10430);
or U11106 (N_11106,N_9957,N_10465);
xor U11107 (N_11107,N_9760,N_9785);
or U11108 (N_11108,N_10488,N_9893);
or U11109 (N_11109,N_10117,N_10062);
nand U11110 (N_11110,N_9750,N_9940);
nand U11111 (N_11111,N_10347,N_10166);
and U11112 (N_11112,N_10216,N_10308);
nor U11113 (N_11113,N_10145,N_9950);
and U11114 (N_11114,N_9992,N_9767);
and U11115 (N_11115,N_10479,N_10252);
or U11116 (N_11116,N_9865,N_10234);
nor U11117 (N_11117,N_9920,N_9923);
nand U11118 (N_11118,N_9959,N_9949);
or U11119 (N_11119,N_10225,N_9814);
nand U11120 (N_11120,N_9758,N_10093);
nand U11121 (N_11121,N_10271,N_10137);
nor U11122 (N_11122,N_10383,N_10154);
or U11123 (N_11123,N_10037,N_10376);
and U11124 (N_11124,N_10313,N_9796);
nor U11125 (N_11125,N_10369,N_9835);
and U11126 (N_11126,N_9802,N_10470);
and U11127 (N_11127,N_10079,N_10153);
and U11128 (N_11128,N_9870,N_10155);
nand U11129 (N_11129,N_10219,N_10323);
xor U11130 (N_11130,N_10499,N_9762);
nor U11131 (N_11131,N_10461,N_10226);
or U11132 (N_11132,N_9815,N_10013);
nand U11133 (N_11133,N_10384,N_10240);
nand U11134 (N_11134,N_9781,N_9770);
and U11135 (N_11135,N_10415,N_10383);
xnor U11136 (N_11136,N_9792,N_9818);
and U11137 (N_11137,N_9751,N_10306);
nand U11138 (N_11138,N_10347,N_9783);
xnor U11139 (N_11139,N_9873,N_10315);
nand U11140 (N_11140,N_10056,N_10022);
xor U11141 (N_11141,N_10121,N_10382);
nand U11142 (N_11142,N_10322,N_10434);
nand U11143 (N_11143,N_10348,N_10043);
xor U11144 (N_11144,N_10373,N_10029);
or U11145 (N_11145,N_9934,N_10451);
and U11146 (N_11146,N_10032,N_10100);
nor U11147 (N_11147,N_9867,N_9945);
and U11148 (N_11148,N_10228,N_9795);
nor U11149 (N_11149,N_10151,N_10281);
nor U11150 (N_11150,N_9777,N_9993);
nand U11151 (N_11151,N_10254,N_10265);
and U11152 (N_11152,N_9809,N_10216);
or U11153 (N_11153,N_10079,N_10445);
nand U11154 (N_11154,N_9786,N_9889);
and U11155 (N_11155,N_10051,N_10164);
or U11156 (N_11156,N_10002,N_10083);
nor U11157 (N_11157,N_10482,N_10266);
nand U11158 (N_11158,N_9954,N_10004);
nor U11159 (N_11159,N_10161,N_10271);
or U11160 (N_11160,N_10328,N_10378);
nand U11161 (N_11161,N_9777,N_9945);
nand U11162 (N_11162,N_10175,N_10375);
nor U11163 (N_11163,N_10442,N_9849);
and U11164 (N_11164,N_9951,N_10088);
and U11165 (N_11165,N_9751,N_10435);
and U11166 (N_11166,N_9905,N_9782);
or U11167 (N_11167,N_10191,N_9764);
nor U11168 (N_11168,N_9862,N_10031);
or U11169 (N_11169,N_10388,N_10320);
nand U11170 (N_11170,N_9920,N_9855);
nor U11171 (N_11171,N_10152,N_9975);
and U11172 (N_11172,N_10486,N_10237);
nor U11173 (N_11173,N_10425,N_10349);
and U11174 (N_11174,N_10148,N_10342);
nand U11175 (N_11175,N_9796,N_10288);
nor U11176 (N_11176,N_10105,N_10243);
or U11177 (N_11177,N_10419,N_9927);
nand U11178 (N_11178,N_10422,N_10058);
nand U11179 (N_11179,N_10391,N_9854);
nor U11180 (N_11180,N_10012,N_10169);
nand U11181 (N_11181,N_10494,N_9792);
or U11182 (N_11182,N_9793,N_10191);
and U11183 (N_11183,N_9913,N_10455);
nand U11184 (N_11184,N_10081,N_10190);
and U11185 (N_11185,N_9886,N_10137);
nor U11186 (N_11186,N_10215,N_10364);
nand U11187 (N_11187,N_10348,N_10299);
or U11188 (N_11188,N_10470,N_10022);
nand U11189 (N_11189,N_9923,N_10267);
and U11190 (N_11190,N_10371,N_9778);
and U11191 (N_11191,N_10388,N_10396);
or U11192 (N_11192,N_10481,N_9927);
xor U11193 (N_11193,N_10038,N_10475);
nor U11194 (N_11194,N_10304,N_9838);
and U11195 (N_11195,N_9892,N_10230);
or U11196 (N_11196,N_9894,N_10478);
or U11197 (N_11197,N_10478,N_10080);
and U11198 (N_11198,N_9814,N_10452);
nand U11199 (N_11199,N_10188,N_10244);
or U11200 (N_11200,N_9935,N_10049);
xnor U11201 (N_11201,N_10275,N_10328);
nor U11202 (N_11202,N_10497,N_10112);
or U11203 (N_11203,N_9843,N_10161);
or U11204 (N_11204,N_10209,N_10062);
nand U11205 (N_11205,N_9982,N_10230);
or U11206 (N_11206,N_10046,N_9783);
nor U11207 (N_11207,N_10429,N_10097);
nand U11208 (N_11208,N_10233,N_9807);
or U11209 (N_11209,N_10298,N_10428);
or U11210 (N_11210,N_10377,N_10260);
and U11211 (N_11211,N_9815,N_10286);
nor U11212 (N_11212,N_10340,N_10288);
nor U11213 (N_11213,N_10317,N_10062);
nor U11214 (N_11214,N_9994,N_9916);
or U11215 (N_11215,N_9836,N_10450);
nor U11216 (N_11216,N_9850,N_10021);
or U11217 (N_11217,N_10023,N_10293);
and U11218 (N_11218,N_10357,N_10201);
nor U11219 (N_11219,N_10061,N_10134);
or U11220 (N_11220,N_10428,N_10202);
or U11221 (N_11221,N_10457,N_10326);
nand U11222 (N_11222,N_10000,N_10475);
nor U11223 (N_11223,N_9786,N_10426);
and U11224 (N_11224,N_10137,N_10121);
and U11225 (N_11225,N_9807,N_9839);
or U11226 (N_11226,N_10065,N_10240);
nor U11227 (N_11227,N_10451,N_10226);
or U11228 (N_11228,N_9816,N_9956);
nor U11229 (N_11229,N_10112,N_10466);
or U11230 (N_11230,N_10440,N_9912);
nand U11231 (N_11231,N_10445,N_10212);
or U11232 (N_11232,N_10344,N_9918);
and U11233 (N_11233,N_10152,N_10091);
nand U11234 (N_11234,N_9967,N_10306);
or U11235 (N_11235,N_10479,N_9788);
nand U11236 (N_11236,N_10302,N_9850);
nor U11237 (N_11237,N_9974,N_9902);
and U11238 (N_11238,N_10204,N_9903);
xnor U11239 (N_11239,N_10027,N_9971);
or U11240 (N_11240,N_9952,N_10246);
nand U11241 (N_11241,N_9979,N_10386);
nand U11242 (N_11242,N_9981,N_9898);
xnor U11243 (N_11243,N_9832,N_9917);
nor U11244 (N_11244,N_10407,N_10361);
and U11245 (N_11245,N_9927,N_10358);
or U11246 (N_11246,N_10195,N_10009);
or U11247 (N_11247,N_10070,N_9751);
or U11248 (N_11248,N_10040,N_10124);
and U11249 (N_11249,N_10345,N_10136);
and U11250 (N_11250,N_11053,N_10991);
and U11251 (N_11251,N_10971,N_11249);
nand U11252 (N_11252,N_11209,N_10836);
and U11253 (N_11253,N_11139,N_11176);
and U11254 (N_11254,N_11124,N_10898);
nor U11255 (N_11255,N_10755,N_10751);
nand U11256 (N_11256,N_10580,N_11152);
or U11257 (N_11257,N_10780,N_10634);
nor U11258 (N_11258,N_11113,N_11031);
nand U11259 (N_11259,N_10949,N_11067);
nand U11260 (N_11260,N_10652,N_11142);
nand U11261 (N_11261,N_10639,N_10960);
nor U11262 (N_11262,N_11170,N_10527);
nand U11263 (N_11263,N_11246,N_10814);
nor U11264 (N_11264,N_11122,N_10940);
nor U11265 (N_11265,N_11131,N_10826);
nor U11266 (N_11266,N_10722,N_11174);
or U11267 (N_11267,N_11038,N_10876);
nand U11268 (N_11268,N_10642,N_10602);
nor U11269 (N_11269,N_10885,N_11068);
nand U11270 (N_11270,N_10516,N_10668);
nand U11271 (N_11271,N_11044,N_11070);
nor U11272 (N_11272,N_10636,N_10804);
and U11273 (N_11273,N_10790,N_11111);
and U11274 (N_11274,N_10700,N_10559);
nand U11275 (N_11275,N_10522,N_10524);
nor U11276 (N_11276,N_11158,N_10909);
or U11277 (N_11277,N_10655,N_10797);
or U11278 (N_11278,N_11042,N_10547);
and U11279 (N_11279,N_10690,N_10881);
and U11280 (N_11280,N_11039,N_10761);
and U11281 (N_11281,N_11030,N_10747);
nand U11282 (N_11282,N_11035,N_11085);
and U11283 (N_11283,N_10604,N_11214);
and U11284 (N_11284,N_10831,N_10593);
or U11285 (N_11285,N_10681,N_10710);
nand U11286 (N_11286,N_11024,N_10573);
nor U11287 (N_11287,N_10846,N_10645);
nand U11288 (N_11288,N_10934,N_10965);
and U11289 (N_11289,N_11164,N_10614);
nand U11290 (N_11290,N_10872,N_10834);
nand U11291 (N_11291,N_11028,N_10801);
and U11292 (N_11292,N_11106,N_10654);
and U11293 (N_11293,N_10674,N_10964);
and U11294 (N_11294,N_10656,N_11102);
nor U11295 (N_11295,N_10558,N_10908);
nand U11296 (N_11296,N_10691,N_10554);
and U11297 (N_11297,N_10629,N_11135);
or U11298 (N_11298,N_10536,N_11133);
nor U11299 (N_11299,N_10776,N_11196);
or U11300 (N_11300,N_10570,N_10754);
and U11301 (N_11301,N_10718,N_11061);
or U11302 (N_11302,N_10810,N_10930);
nand U11303 (N_11303,N_11096,N_10637);
nand U11304 (N_11304,N_11076,N_10677);
nor U11305 (N_11305,N_11224,N_10877);
nand U11306 (N_11306,N_10712,N_10982);
and U11307 (N_11307,N_10640,N_11073);
nor U11308 (N_11308,N_11192,N_10744);
nand U11309 (N_11309,N_11151,N_10842);
or U11310 (N_11310,N_10720,N_10918);
or U11311 (N_11311,N_10886,N_10504);
nor U11312 (N_11312,N_11186,N_10711);
or U11313 (N_11313,N_10592,N_10697);
nand U11314 (N_11314,N_10986,N_10968);
nor U11315 (N_11315,N_11126,N_10596);
or U11316 (N_11316,N_11175,N_11057);
or U11317 (N_11317,N_11244,N_11115);
and U11318 (N_11318,N_11098,N_10803);
or U11319 (N_11319,N_10560,N_10781);
or U11320 (N_11320,N_10648,N_10868);
or U11321 (N_11321,N_11161,N_11237);
or U11322 (N_11322,N_10992,N_10925);
nor U11323 (N_11323,N_10764,N_11091);
and U11324 (N_11324,N_10533,N_10651);
nand U11325 (N_11325,N_10958,N_10505);
nand U11326 (N_11326,N_10721,N_10766);
and U11327 (N_11327,N_11074,N_10724);
nor U11328 (N_11328,N_10920,N_10815);
and U11329 (N_11329,N_10782,N_10743);
nand U11330 (N_11330,N_10963,N_11027);
nor U11331 (N_11331,N_10565,N_10738);
nor U11332 (N_11332,N_10862,N_11206);
or U11333 (N_11333,N_10848,N_11202);
nor U11334 (N_11334,N_11094,N_11146);
or U11335 (N_11335,N_10594,N_11213);
and U11336 (N_11336,N_10546,N_11018);
or U11337 (N_11337,N_11181,N_10799);
nor U11338 (N_11338,N_10715,N_11087);
nand U11339 (N_11339,N_10649,N_11143);
and U11340 (N_11340,N_11183,N_11000);
and U11341 (N_11341,N_10658,N_11032);
nor U11342 (N_11342,N_11112,N_10882);
nor U11343 (N_11343,N_10823,N_10609);
nor U11344 (N_11344,N_10859,N_10897);
nor U11345 (N_11345,N_11145,N_10795);
nand U11346 (N_11346,N_11165,N_10816);
and U11347 (N_11347,N_11166,N_10852);
nor U11348 (N_11348,N_10748,N_10773);
and U11349 (N_11349,N_10980,N_10921);
nor U11350 (N_11350,N_11086,N_10575);
nand U11351 (N_11351,N_10974,N_10551);
and U11352 (N_11352,N_10617,N_10938);
nand U11353 (N_11353,N_11182,N_11003);
and U11354 (N_11354,N_10703,N_11215);
and U11355 (N_11355,N_10684,N_10557);
and U11356 (N_11356,N_10800,N_10664);
or U11357 (N_11357,N_10996,N_10706);
nor U11358 (N_11358,N_11088,N_10623);
nand U11359 (N_11359,N_10981,N_11107);
nand U11360 (N_11360,N_10913,N_10556);
or U11361 (N_11361,N_10895,N_11236);
nand U11362 (N_11362,N_10687,N_10611);
xor U11363 (N_11363,N_11089,N_10583);
nor U11364 (N_11364,N_10979,N_10613);
nor U11365 (N_11365,N_11156,N_11218);
nand U11366 (N_11366,N_11168,N_11242);
and U11367 (N_11367,N_10577,N_10912);
nor U11368 (N_11368,N_10999,N_10535);
nand U11369 (N_11369,N_10817,N_10545);
nand U11370 (N_11370,N_10789,N_11172);
and U11371 (N_11371,N_10669,N_10922);
and U11372 (N_11372,N_10727,N_10796);
or U11373 (N_11373,N_10967,N_10729);
or U11374 (N_11374,N_10973,N_10856);
and U11375 (N_11375,N_10653,N_11138);
and U11376 (N_11376,N_11020,N_11101);
nand U11377 (N_11377,N_10578,N_10830);
or U11378 (N_11378,N_10736,N_10910);
or U11379 (N_11379,N_11178,N_11022);
xor U11380 (N_11380,N_11149,N_11123);
nor U11381 (N_11381,N_10665,N_10605);
xnor U11382 (N_11382,N_10772,N_10569);
nand U11383 (N_11383,N_11210,N_10926);
xnor U11384 (N_11384,N_11048,N_10660);
or U11385 (N_11385,N_10907,N_10869);
or U11386 (N_11386,N_11180,N_10784);
nor U11387 (N_11387,N_10512,N_10673);
and U11388 (N_11388,N_10702,N_10716);
or U11389 (N_11389,N_11064,N_11205);
or U11390 (N_11390,N_11195,N_11216);
nor U11391 (N_11391,N_10879,N_10788);
or U11392 (N_11392,N_10574,N_11239);
nand U11393 (N_11393,N_10820,N_10983);
nand U11394 (N_11394,N_11110,N_10822);
or U11395 (N_11395,N_11160,N_10663);
and U11396 (N_11396,N_10944,N_10819);
nand U11397 (N_11397,N_10765,N_10919);
nand U11398 (N_11398,N_10756,N_11046);
or U11399 (N_11399,N_11014,N_11189);
nor U11400 (N_11400,N_10998,N_10942);
nor U11401 (N_11401,N_11043,N_10825);
or U11402 (N_11402,N_10507,N_10995);
nand U11403 (N_11403,N_10798,N_10643);
nand U11404 (N_11404,N_10576,N_10887);
nand U11405 (N_11405,N_10899,N_11025);
or U11406 (N_11406,N_10923,N_11023);
or U11407 (N_11407,N_11050,N_10564);
and U11408 (N_11408,N_10863,N_11080);
nor U11409 (N_11409,N_10948,N_10883);
and U11410 (N_11410,N_10767,N_10515);
nor U11411 (N_11411,N_10728,N_10933);
or U11412 (N_11412,N_11033,N_10771);
nand U11413 (N_11413,N_10571,N_11203);
or U11414 (N_11414,N_10813,N_10726);
and U11415 (N_11415,N_10977,N_10589);
and U11416 (N_11416,N_10827,N_10845);
nor U11417 (N_11417,N_10851,N_11193);
nor U11418 (N_11418,N_11002,N_11058);
and U11419 (N_11419,N_10550,N_11227);
xnor U11420 (N_11420,N_10915,N_10662);
and U11421 (N_11421,N_10628,N_11201);
and U11422 (N_11422,N_11225,N_10855);
nand U11423 (N_11423,N_11167,N_10840);
and U11424 (N_11424,N_10758,N_10618);
nand U11425 (N_11425,N_10709,N_11200);
or U11426 (N_11426,N_10587,N_10946);
or U11427 (N_11427,N_10952,N_10737);
or U11428 (N_11428,N_10552,N_11051);
nor U11429 (N_11429,N_11054,N_10821);
nor U11430 (N_11430,N_10941,N_10950);
or U11431 (N_11431,N_11127,N_11154);
and U11432 (N_11432,N_10763,N_10770);
and U11433 (N_11433,N_10679,N_11063);
xor U11434 (N_11434,N_10793,N_11229);
nor U11435 (N_11435,N_10695,N_10541);
and U11436 (N_11436,N_10959,N_11134);
nand U11437 (N_11437,N_10905,N_11171);
nand U11438 (N_11438,N_10549,N_10791);
nor U11439 (N_11439,N_10670,N_11093);
nor U11440 (N_11440,N_10633,N_11235);
or U11441 (N_11441,N_10838,N_10947);
or U11442 (N_11442,N_11060,N_10590);
nand U11443 (N_11443,N_10870,N_10532);
or U11444 (N_11444,N_11012,N_10742);
or U11445 (N_11445,N_10599,N_10786);
and U11446 (N_11446,N_11105,N_10635);
or U11447 (N_11447,N_10988,N_11097);
or U11448 (N_11448,N_10752,N_10957);
nor U11449 (N_11449,N_10581,N_11121);
or U11450 (N_11450,N_10762,N_10671);
and U11451 (N_11451,N_10517,N_10719);
and U11452 (N_11452,N_10750,N_11034);
nand U11453 (N_11453,N_10531,N_11036);
nor U11454 (N_11454,N_11011,N_10745);
nand U11455 (N_11455,N_11231,N_11045);
or U11456 (N_11456,N_10875,N_10843);
or U11457 (N_11457,N_11062,N_10794);
or U11458 (N_11458,N_11132,N_10841);
nor U11459 (N_11459,N_10854,N_10625);
and U11460 (N_11460,N_10603,N_10607);
nor U11461 (N_11461,N_10929,N_11245);
or U11462 (N_11462,N_10686,N_11095);
and U11463 (N_11463,N_11117,N_11019);
or U11464 (N_11464,N_11232,N_10543);
nor U11465 (N_11465,N_10503,N_10659);
nand U11466 (N_11466,N_10666,N_11118);
or U11467 (N_11467,N_10867,N_10548);
and U11468 (N_11468,N_10987,N_11148);
nand U11469 (N_11469,N_10866,N_11010);
nor U11470 (N_11470,N_10588,N_10878);
or U11471 (N_11471,N_11004,N_10847);
nor U11472 (N_11472,N_10566,N_10861);
nor U11473 (N_11473,N_10809,N_10530);
or U11474 (N_11474,N_10699,N_10953);
nor U11475 (N_11475,N_10994,N_10509);
nor U11476 (N_11476,N_10534,N_10975);
nand U11477 (N_11477,N_10612,N_10657);
and U11478 (N_11478,N_10627,N_10701);
nand U11479 (N_11479,N_10704,N_11083);
nor U11480 (N_11480,N_10685,N_10966);
and U11481 (N_11481,N_10945,N_10928);
or U11482 (N_11482,N_11072,N_11220);
nand U11483 (N_11483,N_10936,N_10717);
and U11484 (N_11484,N_10993,N_10586);
or U11485 (N_11485,N_11017,N_11177);
or U11486 (N_11486,N_10760,N_11065);
nor U11487 (N_11487,N_11243,N_10775);
nand U11488 (N_11488,N_10582,N_11155);
and U11489 (N_11489,N_10894,N_11015);
and U11490 (N_11490,N_10778,N_10759);
nand U11491 (N_11491,N_10525,N_10740);
or U11492 (N_11492,N_10931,N_10563);
nor U11493 (N_11493,N_10903,N_10807);
nor U11494 (N_11494,N_11191,N_10544);
and U11495 (N_11495,N_10714,N_10880);
and U11496 (N_11496,N_11008,N_11212);
nor U11497 (N_11497,N_10829,N_10777);
or U11498 (N_11498,N_10916,N_10937);
nor U11499 (N_11499,N_11128,N_10984);
and U11500 (N_11500,N_11071,N_10600);
nand U11501 (N_11501,N_10969,N_11056);
nand U11502 (N_11502,N_11233,N_10978);
and U11503 (N_11503,N_10858,N_10610);
and U11504 (N_11504,N_10753,N_10638);
nor U11505 (N_11505,N_10641,N_10956);
nor U11506 (N_11506,N_11234,N_10561);
or U11507 (N_11507,N_10537,N_11219);
and U11508 (N_11508,N_10888,N_10833);
nor U11509 (N_11509,N_10774,N_11040);
and U11510 (N_11510,N_10568,N_10528);
xnor U11511 (N_11511,N_11016,N_11187);
and U11512 (N_11512,N_11190,N_11049);
nor U11513 (N_11513,N_10824,N_10779);
nor U11514 (N_11514,N_10951,N_10874);
or U11515 (N_11515,N_10529,N_11144);
or U11516 (N_11516,N_10631,N_10502);
nand U11517 (N_11517,N_10676,N_10806);
and U11518 (N_11518,N_11184,N_10783);
and U11519 (N_11519,N_11078,N_11079);
and U11520 (N_11520,N_10901,N_11208);
nor U11521 (N_11521,N_10526,N_11137);
nand U11522 (N_11522,N_10990,N_10924);
nand U11523 (N_11523,N_11005,N_10630);
and U11524 (N_11524,N_10723,N_11217);
nand U11525 (N_11525,N_10500,N_10508);
nor U11526 (N_11526,N_10539,N_10802);
nor U11527 (N_11527,N_11082,N_10939);
nand U11528 (N_11528,N_10615,N_10572);
and U11529 (N_11529,N_10914,N_10860);
and U11530 (N_11530,N_10997,N_10540);
nor U11531 (N_11531,N_11006,N_10976);
nand U11532 (N_11532,N_10579,N_10632);
or U11533 (N_11533,N_11084,N_10989);
or U11534 (N_11534,N_11052,N_10889);
and U11535 (N_11535,N_11150,N_11013);
and U11536 (N_11536,N_10917,N_10961);
nand U11537 (N_11537,N_11026,N_10511);
or U11538 (N_11538,N_10890,N_10972);
or U11539 (N_11539,N_11129,N_11136);
nor U11540 (N_11540,N_10892,N_10521);
nor U11541 (N_11541,N_11163,N_10844);
or U11542 (N_11542,N_10601,N_10538);
or U11543 (N_11543,N_10849,N_11081);
and U11544 (N_11544,N_11247,N_10619);
and U11545 (N_11545,N_10884,N_10927);
or U11546 (N_11546,N_11221,N_11204);
nand U11547 (N_11547,N_10891,N_11116);
nor U11548 (N_11548,N_10707,N_10735);
nand U11549 (N_11549,N_10510,N_10585);
or U11550 (N_11550,N_10622,N_10732);
and U11551 (N_11551,N_11092,N_10906);
nand U11552 (N_11552,N_10962,N_10514);
or U11553 (N_11553,N_10692,N_11240);
and U11554 (N_11554,N_11147,N_10713);
nand U11555 (N_11555,N_10620,N_10693);
or U11556 (N_11556,N_11069,N_10694);
nand U11557 (N_11557,N_11179,N_10705);
or U11558 (N_11558,N_11157,N_10562);
and U11559 (N_11559,N_11248,N_11228);
nor U11560 (N_11560,N_10864,N_11047);
and U11561 (N_11561,N_11141,N_11162);
and U11562 (N_11562,N_10698,N_10787);
nor U11563 (N_11563,N_10911,N_10768);
nor U11564 (N_11564,N_10661,N_11238);
or U11565 (N_11565,N_10626,N_10896);
nand U11566 (N_11566,N_10506,N_10857);
nor U11567 (N_11567,N_11109,N_11223);
nand U11568 (N_11568,N_11120,N_10584);
or U11569 (N_11569,N_10902,N_10832);
nor U11570 (N_11570,N_10650,N_11125);
or U11571 (N_11571,N_11103,N_11055);
and U11572 (N_11572,N_10520,N_11199);
and U11573 (N_11573,N_11090,N_11241);
nor U11574 (N_11574,N_10688,N_10850);
or U11575 (N_11575,N_10792,N_10769);
nand U11576 (N_11576,N_10812,N_10893);
nor U11577 (N_11577,N_10621,N_11114);
nand U11578 (N_11578,N_10746,N_10646);
nand U11579 (N_11579,N_11009,N_11226);
and U11580 (N_11580,N_10696,N_10808);
nand U11581 (N_11581,N_10739,N_10553);
and U11582 (N_11582,N_10523,N_10954);
or U11583 (N_11583,N_11222,N_10501);
and U11584 (N_11584,N_11207,N_11104);
or U11585 (N_11585,N_11130,N_10606);
nor U11586 (N_11586,N_11169,N_10598);
or U11587 (N_11587,N_10672,N_11100);
nand U11588 (N_11588,N_10542,N_10595);
nand U11589 (N_11589,N_10865,N_10597);
nand U11590 (N_11590,N_10955,N_10828);
and U11591 (N_11591,N_10608,N_10900);
and U11592 (N_11592,N_11066,N_10734);
xnor U11593 (N_11593,N_10839,N_11119);
nor U11594 (N_11594,N_10749,N_10741);
or U11595 (N_11595,N_11021,N_10811);
and U11596 (N_11596,N_10513,N_10904);
nor U11597 (N_11597,N_10678,N_11159);
or U11598 (N_11598,N_10667,N_11059);
or U11599 (N_11599,N_10555,N_10680);
or U11600 (N_11600,N_10683,N_11198);
nor U11601 (N_11601,N_10932,N_11188);
nor U11602 (N_11602,N_10935,N_10591);
and U11603 (N_11603,N_10818,N_10567);
xor U11604 (N_11604,N_10853,N_11007);
nand U11605 (N_11605,N_10805,N_10682);
nor U11606 (N_11606,N_10731,N_10970);
and U11607 (N_11607,N_10871,N_11173);
nand U11608 (N_11608,N_11029,N_10624);
nand U11609 (N_11609,N_11077,N_10518);
or U11610 (N_11610,N_11041,N_10985);
and U11611 (N_11611,N_10675,N_11037);
or U11612 (N_11612,N_11108,N_10873);
nand U11613 (N_11613,N_10733,N_10708);
nand U11614 (N_11614,N_11099,N_10616);
nand U11615 (N_11615,N_10835,N_11185);
and U11616 (N_11616,N_10730,N_10647);
nor U11617 (N_11617,N_10943,N_11075);
and U11618 (N_11618,N_10519,N_10644);
or U11619 (N_11619,N_11153,N_11211);
nor U11620 (N_11620,N_10837,N_11194);
nand U11621 (N_11621,N_10725,N_11197);
and U11622 (N_11622,N_10689,N_10785);
and U11623 (N_11623,N_10757,N_11140);
or U11624 (N_11624,N_11001,N_11230);
or U11625 (N_11625,N_10939,N_10877);
nor U11626 (N_11626,N_10992,N_11116);
or U11627 (N_11627,N_11031,N_10711);
nand U11628 (N_11628,N_10945,N_10660);
or U11629 (N_11629,N_11160,N_10705);
or U11630 (N_11630,N_10857,N_11244);
and U11631 (N_11631,N_11200,N_10890);
nor U11632 (N_11632,N_10775,N_10896);
or U11633 (N_11633,N_11176,N_11236);
or U11634 (N_11634,N_10985,N_10653);
nand U11635 (N_11635,N_11202,N_11201);
and U11636 (N_11636,N_10920,N_10504);
nand U11637 (N_11637,N_10609,N_10675);
nand U11638 (N_11638,N_10572,N_11227);
and U11639 (N_11639,N_10967,N_11243);
nor U11640 (N_11640,N_10814,N_11239);
nand U11641 (N_11641,N_11124,N_11114);
nor U11642 (N_11642,N_11121,N_10959);
or U11643 (N_11643,N_10898,N_11145);
and U11644 (N_11644,N_10841,N_11041);
xnor U11645 (N_11645,N_10805,N_10794);
and U11646 (N_11646,N_11237,N_11010);
nor U11647 (N_11647,N_10795,N_10659);
nand U11648 (N_11648,N_10649,N_10673);
nor U11649 (N_11649,N_11006,N_10932);
nand U11650 (N_11650,N_10964,N_10575);
or U11651 (N_11651,N_11128,N_10852);
nand U11652 (N_11652,N_11071,N_11180);
nand U11653 (N_11653,N_10988,N_11165);
and U11654 (N_11654,N_10803,N_11070);
nor U11655 (N_11655,N_11047,N_10807);
and U11656 (N_11656,N_10776,N_10916);
and U11657 (N_11657,N_11024,N_11195);
and U11658 (N_11658,N_10570,N_10684);
nor U11659 (N_11659,N_10755,N_11075);
and U11660 (N_11660,N_10885,N_11113);
and U11661 (N_11661,N_10533,N_10741);
and U11662 (N_11662,N_10855,N_10962);
nor U11663 (N_11663,N_11137,N_11018);
and U11664 (N_11664,N_10892,N_11056);
nor U11665 (N_11665,N_10823,N_10826);
and U11666 (N_11666,N_10815,N_10700);
and U11667 (N_11667,N_10993,N_11228);
nor U11668 (N_11668,N_10573,N_11041);
nor U11669 (N_11669,N_11074,N_11030);
xor U11670 (N_11670,N_10626,N_10738);
and U11671 (N_11671,N_10865,N_10568);
or U11672 (N_11672,N_10805,N_10981);
or U11673 (N_11673,N_10635,N_10961);
or U11674 (N_11674,N_10543,N_11066);
nand U11675 (N_11675,N_10543,N_10597);
or U11676 (N_11676,N_11226,N_10528);
nand U11677 (N_11677,N_11158,N_10620);
nand U11678 (N_11678,N_10814,N_10837);
and U11679 (N_11679,N_11142,N_11242);
or U11680 (N_11680,N_10746,N_11177);
nor U11681 (N_11681,N_10804,N_10609);
nor U11682 (N_11682,N_10973,N_11155);
and U11683 (N_11683,N_10607,N_10524);
and U11684 (N_11684,N_10980,N_10780);
or U11685 (N_11685,N_11103,N_10708);
nor U11686 (N_11686,N_11137,N_11087);
or U11687 (N_11687,N_10600,N_10970);
nand U11688 (N_11688,N_10586,N_11154);
xnor U11689 (N_11689,N_11048,N_10686);
nand U11690 (N_11690,N_10662,N_11102);
nor U11691 (N_11691,N_10875,N_11150);
nand U11692 (N_11692,N_10612,N_10995);
nand U11693 (N_11693,N_10869,N_11190);
or U11694 (N_11694,N_10968,N_11206);
nor U11695 (N_11695,N_10706,N_10729);
nor U11696 (N_11696,N_11038,N_10937);
and U11697 (N_11697,N_10661,N_10752);
or U11698 (N_11698,N_10764,N_10846);
or U11699 (N_11699,N_11055,N_10845);
nor U11700 (N_11700,N_11010,N_10557);
or U11701 (N_11701,N_10774,N_11127);
and U11702 (N_11702,N_10865,N_10676);
nor U11703 (N_11703,N_11029,N_11170);
nor U11704 (N_11704,N_10611,N_10762);
nor U11705 (N_11705,N_11112,N_11170);
or U11706 (N_11706,N_10573,N_10646);
or U11707 (N_11707,N_10837,N_10696);
or U11708 (N_11708,N_11069,N_11032);
or U11709 (N_11709,N_10881,N_11246);
xnor U11710 (N_11710,N_10880,N_10748);
and U11711 (N_11711,N_11049,N_10934);
nor U11712 (N_11712,N_11214,N_10572);
nor U11713 (N_11713,N_10718,N_11154);
or U11714 (N_11714,N_11156,N_10903);
and U11715 (N_11715,N_10954,N_10968);
or U11716 (N_11716,N_10574,N_11175);
and U11717 (N_11717,N_10710,N_11127);
or U11718 (N_11718,N_10782,N_10878);
or U11719 (N_11719,N_10666,N_10610);
nor U11720 (N_11720,N_10875,N_10690);
or U11721 (N_11721,N_11038,N_11216);
or U11722 (N_11722,N_10517,N_10644);
nor U11723 (N_11723,N_10631,N_11193);
nand U11724 (N_11724,N_10936,N_10556);
nor U11725 (N_11725,N_10520,N_11126);
nand U11726 (N_11726,N_10892,N_10950);
or U11727 (N_11727,N_10869,N_11223);
and U11728 (N_11728,N_11131,N_11219);
nor U11729 (N_11729,N_11181,N_10822);
nand U11730 (N_11730,N_10672,N_10685);
nor U11731 (N_11731,N_10864,N_10734);
or U11732 (N_11732,N_10512,N_11248);
or U11733 (N_11733,N_10821,N_10575);
nor U11734 (N_11734,N_11233,N_10920);
nor U11735 (N_11735,N_10714,N_11027);
nand U11736 (N_11736,N_10784,N_11124);
nor U11737 (N_11737,N_10683,N_10682);
nand U11738 (N_11738,N_11067,N_11122);
xnor U11739 (N_11739,N_11128,N_10898);
or U11740 (N_11740,N_10865,N_11136);
nor U11741 (N_11741,N_11076,N_10816);
or U11742 (N_11742,N_10903,N_10908);
and U11743 (N_11743,N_11141,N_11073);
and U11744 (N_11744,N_11062,N_11237);
nor U11745 (N_11745,N_11017,N_11010);
or U11746 (N_11746,N_10583,N_11150);
nor U11747 (N_11747,N_11185,N_10767);
or U11748 (N_11748,N_10918,N_11044);
or U11749 (N_11749,N_10580,N_10867);
nor U11750 (N_11750,N_10501,N_10951);
and U11751 (N_11751,N_11020,N_10896);
nand U11752 (N_11752,N_11116,N_11178);
nand U11753 (N_11753,N_10748,N_11148);
nand U11754 (N_11754,N_10520,N_10850);
and U11755 (N_11755,N_10614,N_10512);
nand U11756 (N_11756,N_10866,N_10852);
or U11757 (N_11757,N_10753,N_10889);
xnor U11758 (N_11758,N_11042,N_10552);
nor U11759 (N_11759,N_11110,N_10874);
nor U11760 (N_11760,N_10746,N_11172);
nand U11761 (N_11761,N_10551,N_11079);
and U11762 (N_11762,N_10547,N_11037);
xnor U11763 (N_11763,N_11150,N_10912);
nand U11764 (N_11764,N_10581,N_10687);
nor U11765 (N_11765,N_11187,N_10577);
or U11766 (N_11766,N_11117,N_10646);
nand U11767 (N_11767,N_11171,N_10593);
nand U11768 (N_11768,N_10881,N_10687);
nand U11769 (N_11769,N_10585,N_11243);
nand U11770 (N_11770,N_11083,N_10524);
and U11771 (N_11771,N_10539,N_10855);
nand U11772 (N_11772,N_10702,N_10696);
nand U11773 (N_11773,N_10710,N_11100);
xor U11774 (N_11774,N_10859,N_10551);
nor U11775 (N_11775,N_10968,N_10866);
and U11776 (N_11776,N_11247,N_10992);
nor U11777 (N_11777,N_10772,N_11242);
and U11778 (N_11778,N_11126,N_11015);
or U11779 (N_11779,N_11162,N_10554);
nor U11780 (N_11780,N_10560,N_10523);
and U11781 (N_11781,N_10622,N_10964);
or U11782 (N_11782,N_10717,N_10998);
nand U11783 (N_11783,N_10907,N_10846);
nand U11784 (N_11784,N_10748,N_11002);
and U11785 (N_11785,N_11192,N_10508);
nand U11786 (N_11786,N_11153,N_11201);
or U11787 (N_11787,N_10881,N_10878);
nor U11788 (N_11788,N_10700,N_11229);
nand U11789 (N_11789,N_10750,N_10684);
or U11790 (N_11790,N_11087,N_10920);
and U11791 (N_11791,N_11029,N_10917);
xnor U11792 (N_11792,N_10741,N_11156);
and U11793 (N_11793,N_10849,N_10523);
nor U11794 (N_11794,N_11111,N_10937);
nand U11795 (N_11795,N_11054,N_10923);
and U11796 (N_11796,N_10762,N_10786);
and U11797 (N_11797,N_11204,N_11113);
nand U11798 (N_11798,N_10537,N_11138);
or U11799 (N_11799,N_10953,N_10522);
and U11800 (N_11800,N_10608,N_11196);
or U11801 (N_11801,N_10599,N_10962);
nor U11802 (N_11802,N_11076,N_11216);
or U11803 (N_11803,N_10548,N_10688);
or U11804 (N_11804,N_10996,N_10636);
and U11805 (N_11805,N_11222,N_10574);
nor U11806 (N_11806,N_10951,N_10908);
nor U11807 (N_11807,N_10903,N_10505);
nor U11808 (N_11808,N_10509,N_10656);
or U11809 (N_11809,N_10740,N_11060);
or U11810 (N_11810,N_10813,N_10870);
or U11811 (N_11811,N_10974,N_10722);
or U11812 (N_11812,N_11228,N_10523);
and U11813 (N_11813,N_10570,N_11036);
xnor U11814 (N_11814,N_11047,N_10772);
nand U11815 (N_11815,N_11036,N_10952);
nor U11816 (N_11816,N_10540,N_11030);
nor U11817 (N_11817,N_10506,N_11192);
nor U11818 (N_11818,N_11179,N_11107);
or U11819 (N_11819,N_10554,N_11022);
or U11820 (N_11820,N_10935,N_10618);
nand U11821 (N_11821,N_10641,N_11165);
nand U11822 (N_11822,N_10763,N_10683);
and U11823 (N_11823,N_11017,N_11242);
and U11824 (N_11824,N_11068,N_10712);
nand U11825 (N_11825,N_10717,N_11200);
and U11826 (N_11826,N_11012,N_11074);
nor U11827 (N_11827,N_10895,N_11016);
nor U11828 (N_11828,N_10886,N_10908);
or U11829 (N_11829,N_11125,N_11126);
and U11830 (N_11830,N_10862,N_11126);
nand U11831 (N_11831,N_10856,N_11042);
nor U11832 (N_11832,N_10671,N_10944);
and U11833 (N_11833,N_10798,N_10518);
and U11834 (N_11834,N_11129,N_10618);
and U11835 (N_11835,N_10638,N_11134);
and U11836 (N_11836,N_10571,N_10514);
nor U11837 (N_11837,N_11121,N_11141);
xor U11838 (N_11838,N_10961,N_10773);
nand U11839 (N_11839,N_10679,N_11197);
and U11840 (N_11840,N_11166,N_11001);
nand U11841 (N_11841,N_10963,N_11003);
nor U11842 (N_11842,N_11102,N_10734);
nor U11843 (N_11843,N_10682,N_10834);
or U11844 (N_11844,N_11209,N_10566);
and U11845 (N_11845,N_10606,N_10643);
nand U11846 (N_11846,N_10923,N_10880);
nand U11847 (N_11847,N_10910,N_10513);
or U11848 (N_11848,N_10593,N_11241);
nor U11849 (N_11849,N_10979,N_10554);
nand U11850 (N_11850,N_11194,N_10698);
and U11851 (N_11851,N_10536,N_10538);
or U11852 (N_11852,N_11073,N_10716);
and U11853 (N_11853,N_10887,N_10510);
nand U11854 (N_11854,N_10554,N_11122);
nand U11855 (N_11855,N_10751,N_10662);
or U11856 (N_11856,N_11144,N_10877);
and U11857 (N_11857,N_10518,N_11239);
nor U11858 (N_11858,N_11128,N_11140);
nand U11859 (N_11859,N_10682,N_10842);
or U11860 (N_11860,N_10743,N_10953);
nor U11861 (N_11861,N_10808,N_11229);
or U11862 (N_11862,N_10821,N_10799);
and U11863 (N_11863,N_11125,N_10623);
nand U11864 (N_11864,N_11032,N_10730);
nand U11865 (N_11865,N_11150,N_11085);
nor U11866 (N_11866,N_10911,N_10540);
nand U11867 (N_11867,N_10916,N_11238);
nand U11868 (N_11868,N_10545,N_10727);
nand U11869 (N_11869,N_10628,N_10540);
nor U11870 (N_11870,N_10977,N_11048);
nand U11871 (N_11871,N_10919,N_10722);
or U11872 (N_11872,N_10658,N_10718);
nand U11873 (N_11873,N_10983,N_10673);
and U11874 (N_11874,N_10957,N_10922);
nand U11875 (N_11875,N_10985,N_10535);
nand U11876 (N_11876,N_11018,N_10633);
or U11877 (N_11877,N_10683,N_11004);
nor U11878 (N_11878,N_10661,N_11108);
xor U11879 (N_11879,N_10601,N_10696);
or U11880 (N_11880,N_10745,N_10549);
nand U11881 (N_11881,N_10652,N_10521);
and U11882 (N_11882,N_11114,N_11007);
nand U11883 (N_11883,N_11152,N_10728);
nand U11884 (N_11884,N_10676,N_11063);
nor U11885 (N_11885,N_10731,N_10728);
and U11886 (N_11886,N_11245,N_11106);
and U11887 (N_11887,N_10759,N_11113);
nand U11888 (N_11888,N_10738,N_10641);
and U11889 (N_11889,N_10864,N_10737);
nor U11890 (N_11890,N_10697,N_10910);
nand U11891 (N_11891,N_10889,N_10948);
and U11892 (N_11892,N_10829,N_10801);
and U11893 (N_11893,N_11002,N_10882);
nand U11894 (N_11894,N_10560,N_11071);
nor U11895 (N_11895,N_11133,N_11086);
nor U11896 (N_11896,N_10537,N_11170);
nand U11897 (N_11897,N_10988,N_10780);
and U11898 (N_11898,N_10719,N_11186);
nand U11899 (N_11899,N_10638,N_10760);
and U11900 (N_11900,N_11147,N_10974);
and U11901 (N_11901,N_10704,N_10737);
and U11902 (N_11902,N_10942,N_10720);
or U11903 (N_11903,N_10970,N_11239);
nor U11904 (N_11904,N_11006,N_10633);
or U11905 (N_11905,N_10655,N_10529);
xor U11906 (N_11906,N_10760,N_10580);
nand U11907 (N_11907,N_11235,N_10993);
nor U11908 (N_11908,N_10504,N_11184);
and U11909 (N_11909,N_11011,N_10994);
and U11910 (N_11910,N_11223,N_10962);
nand U11911 (N_11911,N_11194,N_10679);
xor U11912 (N_11912,N_10806,N_10713);
or U11913 (N_11913,N_10611,N_10976);
nand U11914 (N_11914,N_10948,N_11197);
and U11915 (N_11915,N_11031,N_10967);
nand U11916 (N_11916,N_10958,N_10928);
nor U11917 (N_11917,N_10883,N_11241);
nand U11918 (N_11918,N_10787,N_10849);
and U11919 (N_11919,N_10539,N_10987);
nor U11920 (N_11920,N_11135,N_11224);
or U11921 (N_11921,N_10550,N_11063);
or U11922 (N_11922,N_10909,N_10884);
and U11923 (N_11923,N_10747,N_10593);
nand U11924 (N_11924,N_11166,N_10658);
nor U11925 (N_11925,N_10997,N_11208);
nor U11926 (N_11926,N_11035,N_10865);
nor U11927 (N_11927,N_10826,N_11015);
or U11928 (N_11928,N_10893,N_10796);
and U11929 (N_11929,N_11117,N_11110);
or U11930 (N_11930,N_10794,N_11027);
and U11931 (N_11931,N_10580,N_10755);
nand U11932 (N_11932,N_11054,N_11239);
nor U11933 (N_11933,N_10655,N_11235);
nand U11934 (N_11934,N_10583,N_10653);
nor U11935 (N_11935,N_10544,N_11009);
or U11936 (N_11936,N_11070,N_10838);
and U11937 (N_11937,N_11167,N_11001);
xnor U11938 (N_11938,N_11203,N_11035);
and U11939 (N_11939,N_11187,N_10716);
nand U11940 (N_11940,N_11028,N_10789);
nor U11941 (N_11941,N_11124,N_10714);
nand U11942 (N_11942,N_11086,N_10562);
and U11943 (N_11943,N_11018,N_10704);
or U11944 (N_11944,N_10564,N_11008);
or U11945 (N_11945,N_10649,N_10515);
and U11946 (N_11946,N_10783,N_10581);
and U11947 (N_11947,N_10917,N_10746);
nor U11948 (N_11948,N_10704,N_11230);
or U11949 (N_11949,N_11072,N_11237);
nor U11950 (N_11950,N_11222,N_10503);
or U11951 (N_11951,N_10684,N_10679);
or U11952 (N_11952,N_10883,N_10919);
nand U11953 (N_11953,N_11131,N_10810);
nand U11954 (N_11954,N_10675,N_11084);
or U11955 (N_11955,N_10818,N_10580);
and U11956 (N_11956,N_11072,N_10585);
or U11957 (N_11957,N_10739,N_10813);
or U11958 (N_11958,N_11154,N_10990);
nand U11959 (N_11959,N_10893,N_10637);
nor U11960 (N_11960,N_10821,N_10804);
and U11961 (N_11961,N_10812,N_11125);
nand U11962 (N_11962,N_10837,N_10578);
xnor U11963 (N_11963,N_10878,N_10655);
or U11964 (N_11964,N_11043,N_10945);
or U11965 (N_11965,N_10824,N_10665);
nand U11966 (N_11966,N_10678,N_10761);
or U11967 (N_11967,N_10792,N_10708);
or U11968 (N_11968,N_10619,N_11120);
or U11969 (N_11969,N_11110,N_10687);
nor U11970 (N_11970,N_11097,N_10961);
nor U11971 (N_11971,N_11225,N_11150);
nand U11972 (N_11972,N_11009,N_10765);
or U11973 (N_11973,N_10780,N_11111);
nor U11974 (N_11974,N_11061,N_11067);
and U11975 (N_11975,N_11200,N_10598);
or U11976 (N_11976,N_11147,N_11182);
and U11977 (N_11977,N_10521,N_11073);
nor U11978 (N_11978,N_10607,N_10757);
nand U11979 (N_11979,N_10540,N_11141);
and U11980 (N_11980,N_10538,N_10589);
nor U11981 (N_11981,N_11070,N_10788);
and U11982 (N_11982,N_10513,N_11120);
or U11983 (N_11983,N_10872,N_10956);
nor U11984 (N_11984,N_11200,N_11195);
and U11985 (N_11985,N_10565,N_10903);
and U11986 (N_11986,N_10508,N_11087);
nand U11987 (N_11987,N_11049,N_10714);
nand U11988 (N_11988,N_11037,N_11138);
or U11989 (N_11989,N_10668,N_10627);
and U11990 (N_11990,N_10934,N_10659);
and U11991 (N_11991,N_11104,N_10577);
or U11992 (N_11992,N_11003,N_10635);
nand U11993 (N_11993,N_10566,N_11022);
nor U11994 (N_11994,N_11077,N_10976);
and U11995 (N_11995,N_10965,N_10728);
or U11996 (N_11996,N_10975,N_11002);
or U11997 (N_11997,N_10883,N_10501);
nor U11998 (N_11998,N_10751,N_11071);
xor U11999 (N_11999,N_10529,N_10696);
nand U12000 (N_12000,N_11406,N_11742);
or U12001 (N_12001,N_11384,N_11996);
nor U12002 (N_12002,N_11943,N_11734);
nor U12003 (N_12003,N_11444,N_11906);
nand U12004 (N_12004,N_11741,N_11818);
nor U12005 (N_12005,N_11710,N_11763);
and U12006 (N_12006,N_11748,N_11489);
and U12007 (N_12007,N_11524,N_11436);
and U12008 (N_12008,N_11886,N_11671);
or U12009 (N_12009,N_11754,N_11534);
nor U12010 (N_12010,N_11473,N_11761);
or U12011 (N_12011,N_11801,N_11343);
nand U12012 (N_12012,N_11362,N_11861);
or U12013 (N_12013,N_11328,N_11958);
or U12014 (N_12014,N_11461,N_11913);
and U12015 (N_12015,N_11970,N_11568);
and U12016 (N_12016,N_11645,N_11768);
or U12017 (N_12017,N_11796,N_11610);
or U12018 (N_12018,N_11317,N_11577);
and U12019 (N_12019,N_11853,N_11361);
and U12020 (N_12020,N_11306,N_11326);
and U12021 (N_12021,N_11668,N_11371);
nor U12022 (N_12022,N_11498,N_11252);
and U12023 (N_12023,N_11942,N_11960);
nor U12024 (N_12024,N_11916,N_11466);
nand U12025 (N_12025,N_11992,N_11821);
nor U12026 (N_12026,N_11480,N_11695);
nor U12027 (N_12027,N_11562,N_11363);
nor U12028 (N_12028,N_11256,N_11767);
and U12029 (N_12029,N_11526,N_11554);
nor U12030 (N_12030,N_11787,N_11948);
nand U12031 (N_12031,N_11263,N_11520);
or U12032 (N_12032,N_11376,N_11602);
or U12033 (N_12033,N_11826,N_11733);
or U12034 (N_12034,N_11651,N_11907);
nand U12035 (N_12035,N_11389,N_11912);
and U12036 (N_12036,N_11581,N_11936);
nand U12037 (N_12037,N_11421,N_11450);
or U12038 (N_12038,N_11844,N_11267);
nand U12039 (N_12039,N_11337,N_11595);
nand U12040 (N_12040,N_11425,N_11510);
and U12041 (N_12041,N_11762,N_11513);
and U12042 (N_12042,N_11333,N_11437);
or U12043 (N_12043,N_11841,N_11332);
nor U12044 (N_12044,N_11643,N_11751);
nor U12045 (N_12045,N_11653,N_11507);
nor U12046 (N_12046,N_11415,N_11314);
nor U12047 (N_12047,N_11309,N_11257);
nand U12048 (N_12048,N_11722,N_11292);
nor U12049 (N_12049,N_11419,N_11338);
nand U12050 (N_12050,N_11323,N_11740);
or U12051 (N_12051,N_11885,N_11381);
nand U12052 (N_12052,N_11685,N_11692);
nor U12053 (N_12053,N_11542,N_11588);
nor U12054 (N_12054,N_11583,N_11411);
and U12055 (N_12055,N_11879,N_11340);
and U12056 (N_12056,N_11989,N_11817);
nand U12057 (N_12057,N_11730,N_11459);
nor U12058 (N_12058,N_11347,N_11709);
and U12059 (N_12059,N_11639,N_11559);
nand U12060 (N_12060,N_11941,N_11931);
nand U12061 (N_12061,N_11735,N_11327);
nor U12062 (N_12062,N_11616,N_11403);
and U12063 (N_12063,N_11999,N_11860);
or U12064 (N_12064,N_11576,N_11351);
and U12065 (N_12065,N_11802,N_11451);
and U12066 (N_12066,N_11928,N_11873);
nand U12067 (N_12067,N_11519,N_11260);
nor U12068 (N_12068,N_11423,N_11688);
nor U12069 (N_12069,N_11530,N_11500);
and U12070 (N_12070,N_11738,N_11689);
nand U12071 (N_12071,N_11904,N_11478);
and U12072 (N_12072,N_11615,N_11724);
nand U12073 (N_12073,N_11460,N_11587);
or U12074 (N_12074,N_11954,N_11823);
nand U12075 (N_12075,N_11693,N_11798);
nand U12076 (N_12076,N_11998,N_11868);
nand U12077 (N_12077,N_11463,N_11650);
or U12078 (N_12078,N_11882,N_11548);
nand U12079 (N_12079,N_11586,N_11638);
nand U12080 (N_12080,N_11325,N_11287);
and U12081 (N_12081,N_11812,N_11795);
xnor U12082 (N_12082,N_11666,N_11330);
or U12083 (N_12083,N_11825,N_11756);
and U12084 (N_12084,N_11646,N_11346);
nand U12085 (N_12085,N_11273,N_11792);
nor U12086 (N_12086,N_11496,N_11855);
and U12087 (N_12087,N_11870,N_11951);
xor U12088 (N_12088,N_11404,N_11440);
and U12089 (N_12089,N_11301,N_11280);
or U12090 (N_12090,N_11969,N_11591);
nand U12091 (N_12091,N_11471,N_11612);
nor U12092 (N_12092,N_11871,N_11428);
nand U12093 (N_12093,N_11828,N_11558);
nand U12094 (N_12094,N_11445,N_11728);
or U12095 (N_12095,N_11387,N_11431);
nand U12096 (N_12096,N_11791,N_11929);
and U12097 (N_12097,N_11973,N_11902);
nor U12098 (N_12098,N_11848,N_11290);
and U12099 (N_12099,N_11438,N_11567);
and U12100 (N_12100,N_11357,N_11657);
and U12101 (N_12101,N_11769,N_11964);
nor U12102 (N_12102,N_11494,N_11298);
nor U12103 (N_12103,N_11753,N_11383);
nor U12104 (N_12104,N_11749,N_11987);
nor U12105 (N_12105,N_11321,N_11794);
or U12106 (N_12106,N_11770,N_11654);
nor U12107 (N_12107,N_11308,N_11674);
nor U12108 (N_12108,N_11909,N_11479);
nor U12109 (N_12109,N_11565,N_11699);
nand U12110 (N_12110,N_11806,N_11569);
or U12111 (N_12111,N_11963,N_11509);
and U12112 (N_12112,N_11551,N_11433);
nor U12113 (N_12113,N_11726,N_11310);
nand U12114 (N_12114,N_11978,N_11789);
or U12115 (N_12115,N_11599,N_11648);
nand U12116 (N_12116,N_11716,N_11427);
nand U12117 (N_12117,N_11944,N_11621);
nor U12118 (N_12118,N_11329,N_11887);
nand U12119 (N_12119,N_11607,N_11315);
and U12120 (N_12120,N_11635,N_11696);
nor U12121 (N_12121,N_11483,N_11687);
or U12122 (N_12122,N_11430,N_11312);
nor U12123 (N_12123,N_11772,N_11661);
nand U12124 (N_12124,N_11755,N_11446);
or U12125 (N_12125,N_11504,N_11283);
nand U12126 (N_12126,N_11304,N_11596);
nor U12127 (N_12127,N_11401,N_11884);
xor U12128 (N_12128,N_11318,N_11543);
nand U12129 (N_12129,N_11535,N_11555);
and U12130 (N_12130,N_11294,N_11506);
or U12131 (N_12131,N_11593,N_11458);
and U12132 (N_12132,N_11994,N_11972);
nand U12133 (N_12133,N_11660,N_11808);
and U12134 (N_12134,N_11512,N_11549);
nand U12135 (N_12135,N_11609,N_11957);
and U12136 (N_12136,N_11358,N_11541);
or U12137 (N_12137,N_11380,N_11874);
nand U12138 (N_12138,N_11707,N_11307);
nor U12139 (N_12139,N_11842,N_11698);
or U12140 (N_12140,N_11493,N_11764);
and U12141 (N_12141,N_11990,N_11765);
or U12142 (N_12142,N_11903,N_11875);
nor U12143 (N_12143,N_11991,N_11619);
nand U12144 (N_12144,N_11391,N_11293);
xnor U12145 (N_12145,N_11525,N_11484);
nor U12146 (N_12146,N_11590,N_11265);
or U12147 (N_12147,N_11636,N_11774);
and U12148 (N_12148,N_11426,N_11258);
nand U12149 (N_12149,N_11271,N_11827);
nor U12150 (N_12150,N_11529,N_11523);
or U12151 (N_12151,N_11417,N_11608);
nor U12152 (N_12152,N_11331,N_11503);
nand U12153 (N_12153,N_11560,N_11546);
or U12154 (N_12154,N_11659,N_11272);
nand U12155 (N_12155,N_11570,N_11266);
nand U12156 (N_12156,N_11515,N_11898);
or U12157 (N_12157,N_11442,N_11274);
nand U12158 (N_12158,N_11597,N_11594);
and U12159 (N_12159,N_11888,N_11311);
nand U12160 (N_12160,N_11275,N_11930);
nor U12161 (N_12161,N_11382,N_11295);
nand U12162 (N_12162,N_11625,N_11516);
or U12163 (N_12163,N_11713,N_11604);
and U12164 (N_12164,N_11354,N_11335);
nor U12165 (N_12165,N_11322,N_11620);
nand U12166 (N_12166,N_11911,N_11938);
nor U12167 (N_12167,N_11614,N_11447);
nand U12168 (N_12168,N_11270,N_11488);
and U12169 (N_12169,N_11250,N_11708);
or U12170 (N_12170,N_11368,N_11644);
and U12171 (N_12171,N_11965,N_11717);
nor U12172 (N_12172,N_11414,N_11804);
or U12173 (N_12173,N_11353,N_11495);
nor U12174 (N_12174,N_11837,N_11829);
or U12175 (N_12175,N_11302,N_11955);
nor U12176 (N_12176,N_11850,N_11470);
or U12177 (N_12177,N_11719,N_11288);
and U12178 (N_12178,N_11681,N_11505);
and U12179 (N_12179,N_11592,N_11531);
and U12180 (N_12180,N_11396,N_11656);
nor U12181 (N_12181,N_11511,N_11883);
nand U12182 (N_12182,N_11679,N_11824);
nand U12183 (N_12183,N_11703,N_11956);
or U12184 (N_12184,N_11889,N_11634);
and U12185 (N_12185,N_11365,N_11890);
nor U12186 (N_12186,N_11374,N_11405);
xor U12187 (N_12187,N_11908,N_11490);
nor U12188 (N_12188,N_11434,N_11672);
or U12189 (N_12189,N_11851,N_11781);
and U12190 (N_12190,N_11839,N_11527);
and U12191 (N_12191,N_11630,N_11784);
or U12192 (N_12192,N_11891,N_11413);
nor U12193 (N_12193,N_11935,N_11780);
and U12194 (N_12194,N_11550,N_11820);
nand U12195 (N_12195,N_11395,N_11857);
and U12196 (N_12196,N_11350,N_11251);
xnor U12197 (N_12197,N_11962,N_11598);
or U12198 (N_12198,N_11665,N_11945);
and U12199 (N_12199,N_11279,N_11296);
nor U12200 (N_12200,N_11676,N_11746);
and U12201 (N_12201,N_11715,N_11711);
nor U12202 (N_12202,N_11947,N_11453);
or U12203 (N_12203,N_11370,N_11881);
or U12204 (N_12204,N_11601,N_11682);
or U12205 (N_12205,N_11375,N_11876);
or U12206 (N_12206,N_11456,N_11854);
and U12207 (N_12207,N_11959,N_11400);
nand U12208 (N_12208,N_11647,N_11392);
nand U12209 (N_12209,N_11838,N_11297);
nand U12210 (N_12210,N_11552,N_11677);
nand U12211 (N_12211,N_11254,N_11778);
nand U12212 (N_12212,N_11932,N_11632);
and U12213 (N_12213,N_11313,N_11253);
or U12214 (N_12214,N_11984,N_11521);
nor U12215 (N_12215,N_11300,N_11649);
nand U12216 (N_12216,N_11561,N_11918);
nor U12217 (N_12217,N_11939,N_11537);
nor U12218 (N_12218,N_11284,N_11356);
and U12219 (N_12219,N_11725,N_11704);
or U12220 (N_12220,N_11961,N_11575);
or U12221 (N_12221,N_11900,N_11303);
nor U12222 (N_12222,N_11934,N_11914);
nand U12223 (N_12223,N_11544,N_11810);
nor U12224 (N_12224,N_11678,N_11448);
and U12225 (N_12225,N_11536,N_11976);
nor U12226 (N_12226,N_11790,N_11872);
nor U12227 (N_12227,N_11971,N_11831);
nand U12228 (N_12228,N_11631,N_11759);
nand U12229 (N_12229,N_11799,N_11259);
nor U12230 (N_12230,N_11545,N_11336);
or U12231 (N_12231,N_11556,N_11432);
nor U12232 (N_12232,N_11319,N_11443);
xor U12233 (N_12233,N_11547,N_11686);
or U12234 (N_12234,N_11320,N_11901);
and U12235 (N_12235,N_11255,N_11341);
xnor U12236 (N_12236,N_11793,N_11675);
nand U12237 (N_12237,N_11514,N_11452);
and U12238 (N_12238,N_11822,N_11502);
and U12239 (N_12239,N_11986,N_11642);
nor U12240 (N_12240,N_11539,N_11846);
and U12241 (N_12241,N_11833,N_11673);
and U12242 (N_12242,N_11814,N_11830);
and U12243 (N_12243,N_11305,N_11455);
or U12244 (N_12244,N_11540,N_11613);
nor U12245 (N_12245,N_11691,N_11758);
xor U12246 (N_12246,N_11469,N_11757);
or U12247 (N_12247,N_11946,N_11475);
nand U12248 (N_12248,N_11486,N_11464);
and U12249 (N_12249,N_11670,N_11640);
or U12250 (N_12250,N_11979,N_11863);
nor U12251 (N_12251,N_11655,N_11373);
nand U12252 (N_12252,N_11779,N_11264);
and U12253 (N_12253,N_11348,N_11933);
or U12254 (N_12254,N_11416,N_11262);
and U12255 (N_12255,N_11589,N_11840);
nor U12256 (N_12256,N_11269,N_11420);
nand U12257 (N_12257,N_11926,N_11899);
and U12258 (N_12258,N_11624,N_11385);
nor U12259 (N_12259,N_11388,N_11803);
and U12260 (N_12260,N_11892,N_11856);
and U12261 (N_12261,N_11441,N_11983);
nand U12262 (N_12262,N_11422,N_11834);
or U12263 (N_12263,N_11775,N_11584);
and U12264 (N_12264,N_11924,N_11410);
or U12265 (N_12265,N_11532,N_11449);
and U12266 (N_12266,N_11566,N_11574);
nand U12267 (N_12267,N_11334,N_11465);
xnor U12268 (N_12268,N_11866,N_11993);
nand U12269 (N_12269,N_11276,N_11378);
nand U12270 (N_12270,N_11572,N_11797);
nand U12271 (N_12271,N_11750,N_11578);
nor U12272 (N_12272,N_11700,N_11282);
and U12273 (N_12273,N_11342,N_11893);
and U12274 (N_12274,N_11832,N_11807);
nor U12275 (N_12275,N_11760,N_11997);
nand U12276 (N_12276,N_11399,N_11858);
xnor U12277 (N_12277,N_11684,N_11910);
nor U12278 (N_12278,N_11664,N_11501);
and U12279 (N_12279,N_11813,N_11766);
and U12280 (N_12280,N_11582,N_11736);
and U12281 (N_12281,N_11968,N_11737);
nand U12282 (N_12282,N_11980,N_11628);
or U12283 (N_12283,N_11705,N_11905);
nand U12284 (N_12284,N_11407,N_11491);
xor U12285 (N_12285,N_11641,N_11497);
nor U12286 (N_12286,N_11849,N_11720);
or U12287 (N_12287,N_11622,N_11518);
and U12288 (N_12288,N_11988,N_11927);
and U12289 (N_12289,N_11859,N_11667);
or U12290 (N_12290,N_11894,N_11606);
nand U12291 (N_12291,N_11706,N_11811);
nor U12292 (N_12292,N_11472,N_11522);
and U12293 (N_12293,N_11949,N_11268);
nor U12294 (N_12294,N_11285,N_11324);
and U12295 (N_12295,N_11369,N_11771);
nand U12296 (N_12296,N_11937,N_11895);
or U12297 (N_12297,N_11658,N_11950);
nor U12298 (N_12298,N_11800,N_11402);
nor U12299 (N_12299,N_11585,N_11862);
or U12300 (N_12300,N_11739,N_11925);
or U12301 (N_12301,N_11680,N_11835);
nand U12302 (N_12302,N_11915,N_11836);
and U12303 (N_12303,N_11398,N_11605);
nand U12304 (N_12304,N_11424,N_11457);
and U12305 (N_12305,N_11286,N_11517);
and U12306 (N_12306,N_11579,N_11721);
or U12307 (N_12307,N_11880,N_11487);
and U12308 (N_12308,N_11393,N_11474);
xor U12309 (N_12309,N_11299,N_11786);
nand U12310 (N_12310,N_11985,N_11694);
nand U12311 (N_12311,N_11468,N_11669);
nor U12312 (N_12312,N_11919,N_11809);
nor U12313 (N_12313,N_11623,N_11553);
or U12314 (N_12314,N_11953,N_11435);
nor U12315 (N_12315,N_11785,N_11477);
nand U12316 (N_12316,N_11372,N_11409);
nand U12317 (N_12317,N_11379,N_11847);
and U12318 (N_12318,N_11805,N_11611);
and U12319 (N_12319,N_11600,N_11845);
nor U12320 (N_12320,N_11982,N_11974);
nand U12321 (N_12321,N_11701,N_11364);
nand U12322 (N_12322,N_11731,N_11690);
and U12323 (N_12323,N_11788,N_11747);
and U12324 (N_12324,N_11852,N_11439);
or U12325 (N_12325,N_11394,N_11864);
nand U12326 (N_12326,N_11476,N_11714);
nand U12327 (N_12327,N_11896,N_11683);
or U12328 (N_12328,N_11773,N_11627);
nand U12329 (N_12329,N_11481,N_11629);
nor U12330 (N_12330,N_11349,N_11967);
nand U12331 (N_12331,N_11776,N_11727);
nor U12332 (N_12332,N_11777,N_11359);
nor U12333 (N_12333,N_11819,N_11366);
nand U12334 (N_12334,N_11729,N_11580);
or U12335 (N_12335,N_11718,N_11345);
and U12336 (N_12336,N_11744,N_11843);
and U12337 (N_12337,N_11917,N_11386);
xor U12338 (N_12338,N_11662,N_11397);
nor U12339 (N_12339,N_11977,N_11865);
or U12340 (N_12340,N_11557,N_11412);
nand U12341 (N_12341,N_11878,N_11617);
nor U12342 (N_12342,N_11499,N_11816);
nand U12343 (N_12343,N_11723,N_11877);
nand U12344 (N_12344,N_11712,N_11418);
xor U12345 (N_12345,N_11923,N_11360);
nand U12346 (N_12346,N_11277,N_11563);
nand U12347 (N_12347,N_11533,N_11697);
or U12348 (N_12348,N_11940,N_11573);
nor U12349 (N_12349,N_11752,N_11482);
nand U12350 (N_12350,N_11603,N_11377);
or U12351 (N_12351,N_11922,N_11261);
and U12352 (N_12352,N_11339,N_11966);
nand U12353 (N_12353,N_11462,N_11538);
or U12354 (N_12354,N_11637,N_11633);
and U12355 (N_12355,N_11454,N_11408);
and U12356 (N_12356,N_11995,N_11564);
and U12357 (N_12357,N_11352,N_11278);
and U12358 (N_12358,N_11618,N_11815);
or U12359 (N_12359,N_11289,N_11485);
nor U12360 (N_12360,N_11571,N_11745);
nand U12361 (N_12361,N_11467,N_11952);
or U12362 (N_12362,N_11492,N_11981);
and U12363 (N_12363,N_11732,N_11528);
nor U12364 (N_12364,N_11975,N_11783);
and U12365 (N_12365,N_11869,N_11508);
and U12366 (N_12366,N_11390,N_11291);
and U12367 (N_12367,N_11702,N_11367);
and U12368 (N_12368,N_11897,N_11920);
nand U12369 (N_12369,N_11782,N_11429);
or U12370 (N_12370,N_11652,N_11921);
nor U12371 (N_12371,N_11626,N_11281);
or U12372 (N_12372,N_11355,N_11743);
and U12373 (N_12373,N_11867,N_11663);
nand U12374 (N_12374,N_11344,N_11316);
or U12375 (N_12375,N_11998,N_11299);
nor U12376 (N_12376,N_11871,N_11604);
nand U12377 (N_12377,N_11487,N_11977);
nor U12378 (N_12378,N_11985,N_11587);
nand U12379 (N_12379,N_11583,N_11629);
nand U12380 (N_12380,N_11307,N_11889);
nor U12381 (N_12381,N_11582,N_11561);
nor U12382 (N_12382,N_11768,N_11782);
and U12383 (N_12383,N_11621,N_11618);
nor U12384 (N_12384,N_11754,N_11389);
and U12385 (N_12385,N_11312,N_11368);
and U12386 (N_12386,N_11552,N_11984);
nor U12387 (N_12387,N_11769,N_11954);
and U12388 (N_12388,N_11366,N_11316);
nor U12389 (N_12389,N_11264,N_11818);
nand U12390 (N_12390,N_11284,N_11742);
and U12391 (N_12391,N_11716,N_11603);
or U12392 (N_12392,N_11640,N_11368);
or U12393 (N_12393,N_11384,N_11796);
and U12394 (N_12394,N_11536,N_11486);
nor U12395 (N_12395,N_11689,N_11581);
or U12396 (N_12396,N_11309,N_11348);
nand U12397 (N_12397,N_11376,N_11280);
nor U12398 (N_12398,N_11660,N_11781);
and U12399 (N_12399,N_11271,N_11674);
nor U12400 (N_12400,N_11950,N_11387);
nor U12401 (N_12401,N_11559,N_11259);
and U12402 (N_12402,N_11943,N_11724);
or U12403 (N_12403,N_11358,N_11982);
or U12404 (N_12404,N_11744,N_11781);
nor U12405 (N_12405,N_11820,N_11621);
xor U12406 (N_12406,N_11848,N_11279);
nand U12407 (N_12407,N_11832,N_11925);
or U12408 (N_12408,N_11742,N_11967);
and U12409 (N_12409,N_11730,N_11973);
nand U12410 (N_12410,N_11768,N_11764);
or U12411 (N_12411,N_11980,N_11368);
nor U12412 (N_12412,N_11746,N_11682);
and U12413 (N_12413,N_11954,N_11873);
nand U12414 (N_12414,N_11658,N_11616);
nand U12415 (N_12415,N_11334,N_11274);
or U12416 (N_12416,N_11565,N_11376);
or U12417 (N_12417,N_11746,N_11472);
and U12418 (N_12418,N_11911,N_11492);
and U12419 (N_12419,N_11445,N_11311);
or U12420 (N_12420,N_11973,N_11291);
nor U12421 (N_12421,N_11719,N_11360);
nor U12422 (N_12422,N_11430,N_11425);
or U12423 (N_12423,N_11722,N_11475);
xor U12424 (N_12424,N_11953,N_11485);
or U12425 (N_12425,N_11713,N_11950);
nand U12426 (N_12426,N_11342,N_11257);
nand U12427 (N_12427,N_11277,N_11456);
nor U12428 (N_12428,N_11514,N_11714);
and U12429 (N_12429,N_11799,N_11763);
xnor U12430 (N_12430,N_11695,N_11447);
or U12431 (N_12431,N_11964,N_11848);
or U12432 (N_12432,N_11533,N_11880);
nor U12433 (N_12433,N_11458,N_11777);
and U12434 (N_12434,N_11567,N_11914);
nand U12435 (N_12435,N_11945,N_11777);
nand U12436 (N_12436,N_11279,N_11605);
nand U12437 (N_12437,N_11739,N_11620);
and U12438 (N_12438,N_11748,N_11926);
nor U12439 (N_12439,N_11808,N_11874);
nand U12440 (N_12440,N_11800,N_11624);
xor U12441 (N_12441,N_11307,N_11322);
or U12442 (N_12442,N_11637,N_11820);
nand U12443 (N_12443,N_11620,N_11970);
nand U12444 (N_12444,N_11336,N_11260);
and U12445 (N_12445,N_11889,N_11679);
nor U12446 (N_12446,N_11350,N_11549);
or U12447 (N_12447,N_11938,N_11374);
nor U12448 (N_12448,N_11293,N_11797);
and U12449 (N_12449,N_11296,N_11787);
or U12450 (N_12450,N_11797,N_11960);
nand U12451 (N_12451,N_11930,N_11772);
nand U12452 (N_12452,N_11789,N_11517);
or U12453 (N_12453,N_11540,N_11757);
nor U12454 (N_12454,N_11712,N_11572);
and U12455 (N_12455,N_11905,N_11976);
or U12456 (N_12456,N_11844,N_11470);
nand U12457 (N_12457,N_11455,N_11387);
nor U12458 (N_12458,N_11434,N_11633);
and U12459 (N_12459,N_11869,N_11270);
nor U12460 (N_12460,N_11404,N_11268);
or U12461 (N_12461,N_11251,N_11789);
nor U12462 (N_12462,N_11283,N_11986);
nand U12463 (N_12463,N_11407,N_11288);
nand U12464 (N_12464,N_11418,N_11833);
and U12465 (N_12465,N_11262,N_11280);
or U12466 (N_12466,N_11693,N_11302);
and U12467 (N_12467,N_11686,N_11748);
nor U12468 (N_12468,N_11900,N_11872);
and U12469 (N_12469,N_11713,N_11907);
and U12470 (N_12470,N_11878,N_11882);
and U12471 (N_12471,N_11945,N_11954);
nor U12472 (N_12472,N_11293,N_11328);
xnor U12473 (N_12473,N_11589,N_11266);
or U12474 (N_12474,N_11347,N_11977);
nor U12475 (N_12475,N_11327,N_11981);
nor U12476 (N_12476,N_11254,N_11818);
nand U12477 (N_12477,N_11497,N_11575);
nor U12478 (N_12478,N_11958,N_11512);
nor U12479 (N_12479,N_11809,N_11259);
nor U12480 (N_12480,N_11549,N_11913);
nor U12481 (N_12481,N_11296,N_11842);
nor U12482 (N_12482,N_11731,N_11429);
and U12483 (N_12483,N_11873,N_11312);
or U12484 (N_12484,N_11517,N_11757);
or U12485 (N_12485,N_11819,N_11378);
and U12486 (N_12486,N_11578,N_11282);
nand U12487 (N_12487,N_11389,N_11276);
nand U12488 (N_12488,N_11256,N_11318);
nand U12489 (N_12489,N_11489,N_11488);
xor U12490 (N_12490,N_11641,N_11751);
nor U12491 (N_12491,N_11581,N_11576);
nor U12492 (N_12492,N_11467,N_11752);
xnor U12493 (N_12493,N_11352,N_11834);
nor U12494 (N_12494,N_11299,N_11262);
or U12495 (N_12495,N_11603,N_11452);
or U12496 (N_12496,N_11848,N_11859);
nand U12497 (N_12497,N_11841,N_11601);
and U12498 (N_12498,N_11877,N_11805);
and U12499 (N_12499,N_11262,N_11399);
or U12500 (N_12500,N_11295,N_11709);
nor U12501 (N_12501,N_11887,N_11752);
nor U12502 (N_12502,N_11868,N_11833);
nor U12503 (N_12503,N_11968,N_11948);
nand U12504 (N_12504,N_11943,N_11749);
or U12505 (N_12505,N_11739,N_11561);
nor U12506 (N_12506,N_11599,N_11606);
nor U12507 (N_12507,N_11414,N_11413);
nor U12508 (N_12508,N_11696,N_11480);
nor U12509 (N_12509,N_11349,N_11562);
nor U12510 (N_12510,N_11402,N_11796);
and U12511 (N_12511,N_11460,N_11650);
nand U12512 (N_12512,N_11680,N_11845);
nor U12513 (N_12513,N_11792,N_11765);
nor U12514 (N_12514,N_11532,N_11642);
and U12515 (N_12515,N_11979,N_11483);
and U12516 (N_12516,N_11328,N_11815);
nor U12517 (N_12517,N_11955,N_11859);
or U12518 (N_12518,N_11711,N_11527);
nor U12519 (N_12519,N_11250,N_11978);
or U12520 (N_12520,N_11513,N_11662);
nor U12521 (N_12521,N_11712,N_11602);
or U12522 (N_12522,N_11667,N_11942);
xor U12523 (N_12523,N_11809,N_11294);
nor U12524 (N_12524,N_11912,N_11888);
nor U12525 (N_12525,N_11327,N_11831);
or U12526 (N_12526,N_11983,N_11764);
nand U12527 (N_12527,N_11545,N_11414);
nor U12528 (N_12528,N_11913,N_11909);
nor U12529 (N_12529,N_11322,N_11625);
nor U12530 (N_12530,N_11819,N_11386);
and U12531 (N_12531,N_11673,N_11448);
nor U12532 (N_12532,N_11737,N_11903);
nand U12533 (N_12533,N_11525,N_11270);
nand U12534 (N_12534,N_11674,N_11332);
nand U12535 (N_12535,N_11934,N_11619);
nand U12536 (N_12536,N_11783,N_11838);
nand U12537 (N_12537,N_11855,N_11765);
nand U12538 (N_12538,N_11306,N_11957);
or U12539 (N_12539,N_11701,N_11503);
or U12540 (N_12540,N_11399,N_11469);
nand U12541 (N_12541,N_11471,N_11589);
nor U12542 (N_12542,N_11615,N_11625);
nor U12543 (N_12543,N_11610,N_11840);
nor U12544 (N_12544,N_11998,N_11678);
nand U12545 (N_12545,N_11434,N_11334);
xnor U12546 (N_12546,N_11432,N_11254);
or U12547 (N_12547,N_11536,N_11769);
and U12548 (N_12548,N_11888,N_11676);
nor U12549 (N_12549,N_11864,N_11565);
nand U12550 (N_12550,N_11588,N_11418);
or U12551 (N_12551,N_11267,N_11502);
nand U12552 (N_12552,N_11897,N_11554);
and U12553 (N_12553,N_11883,N_11607);
nand U12554 (N_12554,N_11800,N_11981);
or U12555 (N_12555,N_11959,N_11428);
nor U12556 (N_12556,N_11654,N_11823);
nor U12557 (N_12557,N_11926,N_11294);
nor U12558 (N_12558,N_11520,N_11814);
nor U12559 (N_12559,N_11749,N_11935);
nand U12560 (N_12560,N_11665,N_11700);
and U12561 (N_12561,N_11367,N_11729);
nor U12562 (N_12562,N_11576,N_11973);
and U12563 (N_12563,N_11279,N_11471);
or U12564 (N_12564,N_11666,N_11419);
or U12565 (N_12565,N_11487,N_11428);
and U12566 (N_12566,N_11715,N_11906);
or U12567 (N_12567,N_11649,N_11530);
or U12568 (N_12568,N_11565,N_11265);
nand U12569 (N_12569,N_11629,N_11970);
and U12570 (N_12570,N_11691,N_11404);
xor U12571 (N_12571,N_11755,N_11983);
nor U12572 (N_12572,N_11470,N_11799);
xnor U12573 (N_12573,N_11755,N_11811);
nor U12574 (N_12574,N_11363,N_11364);
nand U12575 (N_12575,N_11645,N_11350);
nor U12576 (N_12576,N_11555,N_11253);
or U12577 (N_12577,N_11393,N_11606);
and U12578 (N_12578,N_11709,N_11487);
xor U12579 (N_12579,N_11657,N_11468);
nand U12580 (N_12580,N_11313,N_11550);
nor U12581 (N_12581,N_11353,N_11966);
and U12582 (N_12582,N_11403,N_11617);
nand U12583 (N_12583,N_11490,N_11808);
and U12584 (N_12584,N_11946,N_11459);
nand U12585 (N_12585,N_11444,N_11274);
nor U12586 (N_12586,N_11927,N_11408);
and U12587 (N_12587,N_11911,N_11835);
nor U12588 (N_12588,N_11886,N_11645);
or U12589 (N_12589,N_11376,N_11279);
nor U12590 (N_12590,N_11778,N_11273);
xor U12591 (N_12591,N_11943,N_11362);
xor U12592 (N_12592,N_11256,N_11525);
and U12593 (N_12593,N_11989,N_11753);
or U12594 (N_12594,N_11906,N_11290);
or U12595 (N_12595,N_11368,N_11458);
nand U12596 (N_12596,N_11888,N_11722);
nor U12597 (N_12597,N_11938,N_11565);
and U12598 (N_12598,N_11823,N_11451);
and U12599 (N_12599,N_11555,N_11815);
xnor U12600 (N_12600,N_11400,N_11957);
and U12601 (N_12601,N_11397,N_11711);
nand U12602 (N_12602,N_11260,N_11709);
xnor U12603 (N_12603,N_11364,N_11310);
nand U12604 (N_12604,N_11725,N_11932);
or U12605 (N_12605,N_11967,N_11773);
xnor U12606 (N_12606,N_11619,N_11913);
or U12607 (N_12607,N_11957,N_11668);
nor U12608 (N_12608,N_11555,N_11938);
or U12609 (N_12609,N_11770,N_11652);
and U12610 (N_12610,N_11563,N_11285);
or U12611 (N_12611,N_11892,N_11453);
nand U12612 (N_12612,N_11827,N_11433);
or U12613 (N_12613,N_11444,N_11541);
and U12614 (N_12614,N_11424,N_11599);
nor U12615 (N_12615,N_11894,N_11741);
xor U12616 (N_12616,N_11854,N_11884);
or U12617 (N_12617,N_11544,N_11614);
or U12618 (N_12618,N_11803,N_11927);
nand U12619 (N_12619,N_11683,N_11362);
nor U12620 (N_12620,N_11293,N_11568);
and U12621 (N_12621,N_11966,N_11710);
nor U12622 (N_12622,N_11839,N_11953);
or U12623 (N_12623,N_11950,N_11562);
and U12624 (N_12624,N_11486,N_11874);
and U12625 (N_12625,N_11608,N_11584);
and U12626 (N_12626,N_11887,N_11618);
nor U12627 (N_12627,N_11431,N_11674);
nor U12628 (N_12628,N_11798,N_11673);
and U12629 (N_12629,N_11988,N_11491);
nand U12630 (N_12630,N_11597,N_11286);
xor U12631 (N_12631,N_11585,N_11294);
or U12632 (N_12632,N_11443,N_11418);
and U12633 (N_12633,N_11664,N_11771);
or U12634 (N_12634,N_11519,N_11855);
nor U12635 (N_12635,N_11988,N_11740);
and U12636 (N_12636,N_11654,N_11596);
and U12637 (N_12637,N_11303,N_11395);
and U12638 (N_12638,N_11982,N_11376);
xor U12639 (N_12639,N_11762,N_11511);
or U12640 (N_12640,N_11964,N_11262);
nor U12641 (N_12641,N_11936,N_11423);
or U12642 (N_12642,N_11878,N_11898);
nand U12643 (N_12643,N_11488,N_11294);
and U12644 (N_12644,N_11508,N_11252);
nor U12645 (N_12645,N_11924,N_11678);
nor U12646 (N_12646,N_11647,N_11334);
or U12647 (N_12647,N_11618,N_11486);
or U12648 (N_12648,N_11363,N_11662);
nand U12649 (N_12649,N_11369,N_11300);
nand U12650 (N_12650,N_11254,N_11779);
nor U12651 (N_12651,N_11716,N_11795);
nor U12652 (N_12652,N_11565,N_11324);
or U12653 (N_12653,N_11589,N_11595);
nand U12654 (N_12654,N_11386,N_11959);
nor U12655 (N_12655,N_11425,N_11770);
and U12656 (N_12656,N_11623,N_11562);
and U12657 (N_12657,N_11298,N_11490);
or U12658 (N_12658,N_11781,N_11673);
nand U12659 (N_12659,N_11727,N_11254);
nor U12660 (N_12660,N_11846,N_11348);
nor U12661 (N_12661,N_11987,N_11739);
nand U12662 (N_12662,N_11967,N_11856);
nand U12663 (N_12663,N_11489,N_11648);
nand U12664 (N_12664,N_11656,N_11475);
nand U12665 (N_12665,N_11833,N_11646);
or U12666 (N_12666,N_11274,N_11419);
nand U12667 (N_12667,N_11646,N_11975);
nand U12668 (N_12668,N_11806,N_11585);
nand U12669 (N_12669,N_11795,N_11797);
and U12670 (N_12670,N_11642,N_11667);
or U12671 (N_12671,N_11804,N_11374);
nand U12672 (N_12672,N_11676,N_11310);
and U12673 (N_12673,N_11647,N_11768);
or U12674 (N_12674,N_11283,N_11378);
nor U12675 (N_12675,N_11437,N_11271);
and U12676 (N_12676,N_11514,N_11689);
nand U12677 (N_12677,N_11293,N_11823);
and U12678 (N_12678,N_11733,N_11485);
and U12679 (N_12679,N_11660,N_11399);
or U12680 (N_12680,N_11674,N_11280);
and U12681 (N_12681,N_11876,N_11966);
nor U12682 (N_12682,N_11430,N_11535);
nor U12683 (N_12683,N_11772,N_11337);
nand U12684 (N_12684,N_11318,N_11775);
nor U12685 (N_12685,N_11474,N_11653);
or U12686 (N_12686,N_11360,N_11485);
or U12687 (N_12687,N_11769,N_11411);
nor U12688 (N_12688,N_11667,N_11793);
nor U12689 (N_12689,N_11518,N_11519);
or U12690 (N_12690,N_11988,N_11952);
and U12691 (N_12691,N_11351,N_11779);
and U12692 (N_12692,N_11742,N_11421);
nand U12693 (N_12693,N_11295,N_11303);
nand U12694 (N_12694,N_11989,N_11335);
xor U12695 (N_12695,N_11707,N_11314);
or U12696 (N_12696,N_11333,N_11398);
nor U12697 (N_12697,N_11946,N_11574);
nand U12698 (N_12698,N_11545,N_11848);
or U12699 (N_12699,N_11901,N_11690);
or U12700 (N_12700,N_11731,N_11570);
and U12701 (N_12701,N_11311,N_11467);
nand U12702 (N_12702,N_11855,N_11390);
nand U12703 (N_12703,N_11728,N_11991);
and U12704 (N_12704,N_11569,N_11828);
or U12705 (N_12705,N_11761,N_11804);
nand U12706 (N_12706,N_11264,N_11614);
and U12707 (N_12707,N_11893,N_11971);
nand U12708 (N_12708,N_11796,N_11677);
or U12709 (N_12709,N_11745,N_11673);
nor U12710 (N_12710,N_11559,N_11449);
or U12711 (N_12711,N_11373,N_11311);
and U12712 (N_12712,N_11860,N_11503);
nand U12713 (N_12713,N_11661,N_11458);
nand U12714 (N_12714,N_11285,N_11281);
nand U12715 (N_12715,N_11576,N_11971);
nand U12716 (N_12716,N_11831,N_11793);
or U12717 (N_12717,N_11780,N_11252);
nand U12718 (N_12718,N_11269,N_11329);
and U12719 (N_12719,N_11775,N_11823);
nand U12720 (N_12720,N_11891,N_11521);
or U12721 (N_12721,N_11623,N_11901);
and U12722 (N_12722,N_11784,N_11373);
nand U12723 (N_12723,N_11365,N_11672);
and U12724 (N_12724,N_11534,N_11299);
and U12725 (N_12725,N_11473,N_11287);
nand U12726 (N_12726,N_11955,N_11665);
xor U12727 (N_12727,N_11396,N_11907);
nand U12728 (N_12728,N_11855,N_11717);
nor U12729 (N_12729,N_11973,N_11834);
or U12730 (N_12730,N_11989,N_11960);
nand U12731 (N_12731,N_11399,N_11948);
nor U12732 (N_12732,N_11532,N_11336);
or U12733 (N_12733,N_11599,N_11604);
nand U12734 (N_12734,N_11572,N_11978);
and U12735 (N_12735,N_11771,N_11337);
or U12736 (N_12736,N_11311,N_11790);
nor U12737 (N_12737,N_11276,N_11455);
or U12738 (N_12738,N_11715,N_11330);
and U12739 (N_12739,N_11761,N_11401);
nand U12740 (N_12740,N_11386,N_11491);
and U12741 (N_12741,N_11940,N_11646);
or U12742 (N_12742,N_11395,N_11336);
nor U12743 (N_12743,N_11739,N_11462);
nand U12744 (N_12744,N_11433,N_11555);
nor U12745 (N_12745,N_11697,N_11654);
nor U12746 (N_12746,N_11564,N_11484);
xor U12747 (N_12747,N_11946,N_11263);
or U12748 (N_12748,N_11894,N_11982);
nand U12749 (N_12749,N_11370,N_11571);
or U12750 (N_12750,N_12582,N_12458);
and U12751 (N_12751,N_12669,N_12060);
nand U12752 (N_12752,N_12710,N_12673);
and U12753 (N_12753,N_12742,N_12343);
nor U12754 (N_12754,N_12656,N_12252);
or U12755 (N_12755,N_12520,N_12419);
nand U12756 (N_12756,N_12157,N_12012);
nand U12757 (N_12757,N_12684,N_12098);
or U12758 (N_12758,N_12321,N_12529);
nor U12759 (N_12759,N_12468,N_12709);
or U12760 (N_12760,N_12539,N_12073);
nor U12761 (N_12761,N_12555,N_12714);
or U12762 (N_12762,N_12369,N_12349);
nor U12763 (N_12763,N_12128,N_12659);
xnor U12764 (N_12764,N_12513,N_12324);
or U12765 (N_12765,N_12430,N_12072);
or U12766 (N_12766,N_12246,N_12639);
nor U12767 (N_12767,N_12704,N_12227);
nor U12768 (N_12768,N_12047,N_12233);
or U12769 (N_12769,N_12706,N_12329);
nor U12770 (N_12770,N_12612,N_12033);
or U12771 (N_12771,N_12694,N_12082);
or U12772 (N_12772,N_12665,N_12169);
nand U12773 (N_12773,N_12271,N_12526);
or U12774 (N_12774,N_12168,N_12510);
nor U12775 (N_12775,N_12607,N_12011);
nor U12776 (N_12776,N_12292,N_12002);
or U12777 (N_12777,N_12223,N_12412);
nor U12778 (N_12778,N_12646,N_12186);
and U12779 (N_12779,N_12131,N_12017);
or U12780 (N_12780,N_12117,N_12344);
nand U12781 (N_12781,N_12738,N_12112);
or U12782 (N_12782,N_12103,N_12522);
or U12783 (N_12783,N_12477,N_12148);
nand U12784 (N_12784,N_12456,N_12566);
nor U12785 (N_12785,N_12476,N_12193);
nand U12786 (N_12786,N_12163,N_12201);
or U12787 (N_12787,N_12244,N_12389);
nor U12788 (N_12788,N_12431,N_12268);
nor U12789 (N_12789,N_12417,N_12507);
or U12790 (N_12790,N_12242,N_12400);
xor U12791 (N_12791,N_12494,N_12086);
nand U12792 (N_12792,N_12691,N_12143);
or U12793 (N_12793,N_12726,N_12399);
and U12794 (N_12794,N_12023,N_12018);
and U12795 (N_12795,N_12745,N_12492);
nand U12796 (N_12796,N_12238,N_12631);
nand U12797 (N_12797,N_12040,N_12490);
or U12798 (N_12798,N_12732,N_12303);
nor U12799 (N_12799,N_12683,N_12703);
nand U12800 (N_12800,N_12356,N_12197);
nor U12801 (N_12801,N_12116,N_12693);
xnor U12802 (N_12802,N_12695,N_12099);
nor U12803 (N_12803,N_12453,N_12705);
nor U12804 (N_12804,N_12142,N_12660);
nor U12805 (N_12805,N_12724,N_12104);
nor U12806 (N_12806,N_12406,N_12633);
nor U12807 (N_12807,N_12137,N_12361);
nor U12808 (N_12808,N_12377,N_12000);
or U12809 (N_12809,N_12411,N_12319);
nor U12810 (N_12810,N_12173,N_12578);
or U12811 (N_12811,N_12747,N_12563);
or U12812 (N_12812,N_12110,N_12686);
and U12813 (N_12813,N_12280,N_12249);
nand U12814 (N_12814,N_12382,N_12176);
nand U12815 (N_12815,N_12637,N_12199);
or U12816 (N_12816,N_12122,N_12367);
and U12817 (N_12817,N_12330,N_12003);
and U12818 (N_12818,N_12519,N_12296);
nand U12819 (N_12819,N_12351,N_12636);
or U12820 (N_12820,N_12160,N_12364);
or U12821 (N_12821,N_12149,N_12373);
and U12822 (N_12822,N_12113,N_12467);
nand U12823 (N_12823,N_12595,N_12561);
nand U12824 (N_12824,N_12391,N_12562);
nand U12825 (N_12825,N_12350,N_12679);
nand U12826 (N_12826,N_12415,N_12257);
xnor U12827 (N_12827,N_12312,N_12413);
and U12828 (N_12828,N_12184,N_12346);
or U12829 (N_12829,N_12077,N_12264);
nand U12830 (N_12830,N_12603,N_12090);
nand U12831 (N_12831,N_12590,N_12434);
or U12832 (N_12832,N_12505,N_12056);
nand U12833 (N_12833,N_12697,N_12210);
nor U12834 (N_12834,N_12429,N_12602);
nor U12835 (N_12835,N_12182,N_12470);
or U12836 (N_12836,N_12690,N_12518);
or U12837 (N_12837,N_12301,N_12557);
nand U12838 (N_12838,N_12740,N_12309);
nand U12839 (N_12839,N_12172,N_12304);
and U12840 (N_12840,N_12030,N_12418);
or U12841 (N_12841,N_12258,N_12141);
nor U12842 (N_12842,N_12262,N_12091);
nand U12843 (N_12843,N_12743,N_12071);
nor U12844 (N_12844,N_12611,N_12293);
and U12845 (N_12845,N_12375,N_12632);
nand U12846 (N_12846,N_12594,N_12061);
xnor U12847 (N_12847,N_12010,N_12106);
nand U12848 (N_12848,N_12076,N_12048);
and U12849 (N_12849,N_12069,N_12675);
nor U12850 (N_12850,N_12517,N_12029);
or U12851 (N_12851,N_12663,N_12102);
xnor U12852 (N_12852,N_12386,N_12515);
nor U12853 (N_12853,N_12027,N_12746);
and U12854 (N_12854,N_12081,N_12591);
and U12855 (N_12855,N_12153,N_12674);
or U12856 (N_12856,N_12359,N_12363);
nor U12857 (N_12857,N_12306,N_12063);
xnor U12858 (N_12858,N_12727,N_12008);
nor U12859 (N_12859,N_12536,N_12352);
and U12860 (N_12860,N_12353,N_12028);
or U12861 (N_12861,N_12067,N_12085);
nor U12862 (N_12862,N_12534,N_12336);
nand U12863 (N_12863,N_12692,N_12731);
nand U12864 (N_12864,N_12481,N_12354);
nor U12865 (N_12865,N_12734,N_12243);
nand U12866 (N_12866,N_12652,N_12331);
or U12867 (N_12867,N_12545,N_12339);
or U12868 (N_12868,N_12007,N_12708);
and U12869 (N_12869,N_12298,N_12579);
or U12870 (N_12870,N_12218,N_12613);
nand U12871 (N_12871,N_12118,N_12308);
nand U12872 (N_12872,N_12533,N_12541);
nor U12873 (N_12873,N_12034,N_12586);
or U12874 (N_12874,N_12560,N_12393);
or U12875 (N_12875,N_12164,N_12558);
nand U12876 (N_12876,N_12214,N_12644);
nand U12877 (N_12877,N_12504,N_12688);
or U12878 (N_12878,N_12275,N_12284);
nand U12879 (N_12879,N_12610,N_12715);
and U12880 (N_12880,N_12135,N_12598);
nand U12881 (N_12881,N_12622,N_12383);
or U12882 (N_12882,N_12620,N_12576);
nor U12883 (N_12883,N_12537,N_12402);
nand U12884 (N_12884,N_12256,N_12711);
nor U12885 (N_12885,N_12583,N_12608);
or U12886 (N_12886,N_12667,N_12574);
or U12887 (N_12887,N_12146,N_12315);
nor U12888 (N_12888,N_12016,N_12448);
or U12889 (N_12889,N_12624,N_12449);
and U12890 (N_12890,N_12360,N_12575);
xnor U12891 (N_12891,N_12222,N_12577);
and U12892 (N_12892,N_12295,N_12722);
and U12893 (N_12893,N_12221,N_12682);
or U12894 (N_12894,N_12521,N_12511);
nor U12895 (N_12895,N_12371,N_12634);
nand U12896 (N_12896,N_12328,N_12404);
or U12897 (N_12897,N_12735,N_12443);
nor U12898 (N_12898,N_12119,N_12609);
or U12899 (N_12899,N_12580,N_12635);
or U12900 (N_12900,N_12485,N_12338);
and U12901 (N_12901,N_12744,N_12589);
or U12902 (N_12902,N_12064,N_12604);
and U12903 (N_12903,N_12101,N_12255);
and U12904 (N_12904,N_12203,N_12305);
or U12905 (N_12905,N_12681,N_12089);
nor U12906 (N_12906,N_12035,N_12220);
nand U12907 (N_12907,N_12701,N_12020);
nand U12908 (N_12908,N_12345,N_12668);
nor U12909 (N_12909,N_12124,N_12248);
nand U12910 (N_12910,N_12530,N_12032);
nor U12911 (N_12911,N_12445,N_12551);
and U12912 (N_12912,N_12144,N_12428);
nand U12913 (N_12913,N_12254,N_12538);
or U12914 (N_12914,N_12054,N_12700);
nor U12915 (N_12915,N_12083,N_12278);
nand U12916 (N_12916,N_12230,N_12623);
xor U12917 (N_12917,N_12495,N_12506);
or U12918 (N_12918,N_12341,N_12438);
nand U12919 (N_12919,N_12496,N_12600);
xor U12920 (N_12920,N_12685,N_12488);
and U12921 (N_12921,N_12185,N_12372);
or U12922 (N_12922,N_12599,N_12042);
nor U12923 (N_12923,N_12516,N_12231);
or U12924 (N_12924,N_12190,N_12592);
nor U12925 (N_12925,N_12136,N_12384);
xor U12926 (N_12926,N_12234,N_12297);
or U12927 (N_12927,N_12385,N_12436);
nand U12928 (N_12928,N_12025,N_12721);
nand U12929 (N_12929,N_12707,N_12165);
and U12930 (N_12930,N_12440,N_12426);
nand U12931 (N_12931,N_12676,N_12484);
nor U12932 (N_12932,N_12287,N_12664);
nand U12933 (N_12933,N_12696,N_12217);
nand U12934 (N_12934,N_12272,N_12006);
and U12935 (N_12935,N_12322,N_12314);
nor U12936 (N_12936,N_12626,N_12114);
and U12937 (N_12937,N_12187,N_12627);
nand U12938 (N_12938,N_12074,N_12713);
and U12939 (N_12939,N_12614,N_12587);
and U12940 (N_12940,N_12121,N_12425);
nor U12941 (N_12941,N_12650,N_12410);
or U12942 (N_12942,N_12094,N_12460);
nor U12943 (N_12943,N_12554,N_12045);
and U12944 (N_12944,N_12043,N_12226);
or U12945 (N_12945,N_12605,N_12671);
and U12946 (N_12946,N_12437,N_12191);
nand U12947 (N_12947,N_12316,N_12205);
nor U12948 (N_12948,N_12618,N_12677);
nor U12949 (N_12949,N_12442,N_12568);
nand U12950 (N_12950,N_12617,N_12253);
nand U12951 (N_12951,N_12095,N_12421);
or U12952 (N_12952,N_12347,N_12546);
or U12953 (N_12953,N_12100,N_12718);
nand U12954 (N_12954,N_12125,N_12572);
nor U12955 (N_12955,N_12625,N_12409);
and U12956 (N_12956,N_12672,N_12716);
and U12957 (N_12957,N_12512,N_12235);
nand U12958 (N_12958,N_12161,N_12046);
nand U12959 (N_12959,N_12224,N_12585);
nor U12960 (N_12960,N_12216,N_12736);
nor U12961 (N_12961,N_12208,N_12288);
xnor U12962 (N_12962,N_12155,N_12260);
nor U12963 (N_12963,N_12433,N_12565);
nand U12964 (N_12964,N_12299,N_12240);
and U12965 (N_12965,N_12009,N_12156);
nor U12966 (N_12966,N_12096,N_12283);
nand U12967 (N_12967,N_12263,N_12737);
and U12968 (N_12968,N_12508,N_12597);
nand U12969 (N_12969,N_12424,N_12643);
nand U12970 (N_12970,N_12228,N_12657);
and U12971 (N_12971,N_12648,N_12342);
nand U12972 (N_12972,N_12569,N_12480);
and U12973 (N_12973,N_12024,N_12300);
nor U12974 (N_12974,N_12401,N_12004);
nor U12975 (N_12975,N_12152,N_12088);
and U12976 (N_12976,N_12129,N_12150);
nand U12977 (N_12977,N_12698,N_12212);
nand U12978 (N_12978,N_12318,N_12559);
or U12979 (N_12979,N_12532,N_12446);
nor U12980 (N_12980,N_12188,N_12629);
nor U12981 (N_12981,N_12133,N_12596);
xor U12982 (N_12982,N_12615,N_12464);
nor U12983 (N_12983,N_12049,N_12435);
or U12984 (N_12984,N_12307,N_12621);
nor U12985 (N_12985,N_12057,N_12358);
nor U12986 (N_12986,N_12001,N_12666);
or U12987 (N_12987,N_12368,N_12080);
and U12988 (N_12988,N_12333,N_12134);
and U12989 (N_12989,N_12499,N_12427);
nand U12990 (N_12990,N_12078,N_12447);
nor U12991 (N_12991,N_12289,N_12588);
and U12992 (N_12992,N_12195,N_12570);
and U12993 (N_12993,N_12320,N_12544);
nand U12994 (N_12994,N_12405,N_12274);
and U12995 (N_12995,N_12202,N_12051);
nand U12996 (N_12996,N_12527,N_12092);
or U12997 (N_12997,N_12542,N_12026);
nor U12998 (N_12998,N_12115,N_12337);
nand U12999 (N_12999,N_12403,N_12037);
and U13000 (N_13000,N_12120,N_12500);
or U13001 (N_13001,N_12552,N_12335);
nand U13002 (N_13002,N_12567,N_12107);
or U13003 (N_13003,N_12166,N_12285);
and U13004 (N_13004,N_12712,N_12414);
nor U13005 (N_13005,N_12151,N_12730);
or U13006 (N_13006,N_12466,N_12286);
and U13007 (N_13007,N_12281,N_12454);
or U13008 (N_13008,N_12273,N_12132);
nor U13009 (N_13009,N_12196,N_12439);
nand U13010 (N_13010,N_12649,N_12282);
or U13011 (N_13011,N_12031,N_12105);
nor U13012 (N_13012,N_12139,N_12642);
and U13013 (N_13013,N_12232,N_12111);
and U13014 (N_13014,N_12050,N_12549);
nand U13015 (N_13015,N_12013,N_12325);
nand U13016 (N_13016,N_12501,N_12416);
nand U13017 (N_13017,N_12432,N_12376);
and U13018 (N_13018,N_12179,N_12553);
nor U13019 (N_13019,N_12189,N_12219);
nand U13020 (N_13020,N_12075,N_12702);
nor U13021 (N_13021,N_12465,N_12441);
nor U13022 (N_13022,N_12058,N_12616);
nor U13023 (N_13023,N_12204,N_12066);
and U13024 (N_13024,N_12739,N_12174);
and U13025 (N_13025,N_12245,N_12487);
or U13026 (N_13026,N_12310,N_12229);
and U13027 (N_13027,N_12183,N_12348);
nor U13028 (N_13028,N_12154,N_12159);
and U13029 (N_13029,N_12177,N_12717);
or U13030 (N_13030,N_12525,N_12720);
and U13031 (N_13031,N_12550,N_12327);
and U13032 (N_13032,N_12206,N_12471);
nor U13033 (N_13033,N_12215,N_12236);
nand U13034 (N_13034,N_12138,N_12407);
or U13035 (N_13035,N_12601,N_12455);
nand U13036 (N_13036,N_12171,N_12647);
or U13037 (N_13037,N_12387,N_12162);
nor U13038 (N_13038,N_12323,N_12474);
and U13039 (N_13039,N_12269,N_12019);
or U13040 (N_13040,N_12266,N_12039);
nand U13041 (N_13041,N_12748,N_12317);
or U13042 (N_13042,N_12038,N_12022);
nor U13043 (N_13043,N_12270,N_12564);
nor U13044 (N_13044,N_12380,N_12053);
nand U13045 (N_13045,N_12472,N_12334);
nor U13046 (N_13046,N_12390,N_12654);
and U13047 (N_13047,N_12052,N_12630);
nand U13048 (N_13048,N_12126,N_12420);
or U13049 (N_13049,N_12366,N_12584);
or U13050 (N_13050,N_12689,N_12723);
or U13051 (N_13051,N_12140,N_12398);
or U13052 (N_13052,N_12147,N_12661);
or U13053 (N_13053,N_12491,N_12302);
or U13054 (N_13054,N_12209,N_12370);
nor U13055 (N_13055,N_12241,N_12606);
nand U13056 (N_13056,N_12378,N_12462);
or U13057 (N_13057,N_12524,N_12079);
or U13058 (N_13058,N_12200,N_12540);
and U13059 (N_13059,N_12044,N_12178);
nor U13060 (N_13060,N_12728,N_12408);
or U13061 (N_13061,N_12123,N_12556);
or U13062 (N_13062,N_12489,N_12167);
nor U13063 (N_13063,N_12021,N_12326);
nor U13064 (N_13064,N_12279,N_12379);
and U13065 (N_13065,N_12194,N_12213);
or U13066 (N_13066,N_12547,N_12357);
and U13067 (N_13067,N_12036,N_12482);
or U13068 (N_13068,N_12502,N_12535);
xor U13069 (N_13069,N_12687,N_12145);
xnor U13070 (N_13070,N_12250,N_12093);
nor U13071 (N_13071,N_12493,N_12670);
and U13072 (N_13072,N_12571,N_12514);
and U13073 (N_13073,N_12444,N_12170);
or U13074 (N_13074,N_12207,N_12486);
nor U13075 (N_13075,N_12014,N_12005);
nand U13076 (N_13076,N_12394,N_12459);
and U13077 (N_13077,N_12543,N_12158);
and U13078 (N_13078,N_12503,N_12680);
nand U13079 (N_13079,N_12291,N_12294);
and U13080 (N_13080,N_12059,N_12267);
or U13081 (N_13081,N_12192,N_12619);
nand U13082 (N_13082,N_12340,N_12653);
nand U13083 (N_13083,N_12395,N_12699);
nand U13084 (N_13084,N_12261,N_12641);
nor U13085 (N_13085,N_12108,N_12355);
nor U13086 (N_13086,N_12239,N_12749);
and U13087 (N_13087,N_12397,N_12678);
and U13088 (N_13088,N_12655,N_12311);
nand U13089 (N_13089,N_12109,N_12365);
or U13090 (N_13090,N_12423,N_12247);
nor U13091 (N_13091,N_12548,N_12528);
xor U13092 (N_13092,N_12573,N_12479);
and U13093 (N_13093,N_12725,N_12422);
nor U13094 (N_13094,N_12211,N_12062);
or U13095 (N_13095,N_12070,N_12531);
or U13096 (N_13096,N_12290,N_12180);
xnor U13097 (N_13097,N_12068,N_12084);
and U13098 (N_13098,N_12729,N_12362);
nor U13099 (N_13099,N_12055,N_12175);
or U13100 (N_13100,N_12741,N_12265);
nor U13101 (N_13101,N_12041,N_12225);
or U13102 (N_13102,N_12313,N_12181);
and U13103 (N_13103,N_12593,N_12388);
and U13104 (N_13104,N_12374,N_12015);
nor U13105 (N_13105,N_12087,N_12277);
or U13106 (N_13106,N_12097,N_12478);
xnor U13107 (N_13107,N_12662,N_12198);
or U13108 (N_13108,N_12451,N_12658);
nor U13109 (N_13109,N_12509,N_12450);
and U13110 (N_13110,N_12392,N_12259);
nor U13111 (N_13111,N_12473,N_12645);
or U13112 (N_13112,N_12469,N_12638);
nand U13113 (N_13113,N_12628,N_12640);
nand U13114 (N_13114,N_12719,N_12237);
nor U13115 (N_13115,N_12130,N_12581);
or U13116 (N_13116,N_12251,N_12461);
xnor U13117 (N_13117,N_12498,N_12396);
and U13118 (N_13118,N_12452,N_12483);
nand U13119 (N_13119,N_12332,N_12463);
nand U13120 (N_13120,N_12065,N_12651);
or U13121 (N_13121,N_12523,N_12276);
xnor U13122 (N_13122,N_12381,N_12457);
or U13123 (N_13123,N_12497,N_12475);
or U13124 (N_13124,N_12127,N_12733);
nand U13125 (N_13125,N_12306,N_12637);
or U13126 (N_13126,N_12639,N_12275);
and U13127 (N_13127,N_12419,N_12010);
or U13128 (N_13128,N_12460,N_12281);
nand U13129 (N_13129,N_12238,N_12225);
and U13130 (N_13130,N_12072,N_12283);
nand U13131 (N_13131,N_12635,N_12213);
nand U13132 (N_13132,N_12513,N_12040);
or U13133 (N_13133,N_12579,N_12069);
or U13134 (N_13134,N_12034,N_12434);
or U13135 (N_13135,N_12600,N_12077);
nand U13136 (N_13136,N_12343,N_12686);
or U13137 (N_13137,N_12406,N_12124);
nor U13138 (N_13138,N_12344,N_12220);
and U13139 (N_13139,N_12442,N_12112);
and U13140 (N_13140,N_12239,N_12643);
or U13141 (N_13141,N_12449,N_12303);
nor U13142 (N_13142,N_12591,N_12108);
and U13143 (N_13143,N_12154,N_12246);
or U13144 (N_13144,N_12684,N_12394);
nand U13145 (N_13145,N_12256,N_12636);
nor U13146 (N_13146,N_12748,N_12381);
nand U13147 (N_13147,N_12732,N_12424);
nand U13148 (N_13148,N_12555,N_12557);
nand U13149 (N_13149,N_12265,N_12627);
nand U13150 (N_13150,N_12406,N_12099);
or U13151 (N_13151,N_12459,N_12540);
nand U13152 (N_13152,N_12070,N_12373);
or U13153 (N_13153,N_12354,N_12313);
nand U13154 (N_13154,N_12587,N_12383);
nand U13155 (N_13155,N_12223,N_12406);
and U13156 (N_13156,N_12363,N_12445);
nand U13157 (N_13157,N_12365,N_12396);
nor U13158 (N_13158,N_12587,N_12486);
and U13159 (N_13159,N_12457,N_12586);
and U13160 (N_13160,N_12302,N_12109);
and U13161 (N_13161,N_12683,N_12028);
or U13162 (N_13162,N_12530,N_12648);
or U13163 (N_13163,N_12589,N_12534);
nor U13164 (N_13164,N_12227,N_12613);
or U13165 (N_13165,N_12688,N_12065);
or U13166 (N_13166,N_12598,N_12675);
or U13167 (N_13167,N_12485,N_12167);
and U13168 (N_13168,N_12676,N_12659);
and U13169 (N_13169,N_12212,N_12547);
nand U13170 (N_13170,N_12321,N_12562);
or U13171 (N_13171,N_12125,N_12731);
and U13172 (N_13172,N_12087,N_12076);
xnor U13173 (N_13173,N_12554,N_12363);
nor U13174 (N_13174,N_12499,N_12664);
and U13175 (N_13175,N_12351,N_12321);
nor U13176 (N_13176,N_12191,N_12568);
and U13177 (N_13177,N_12555,N_12722);
nor U13178 (N_13178,N_12587,N_12237);
or U13179 (N_13179,N_12212,N_12570);
or U13180 (N_13180,N_12616,N_12665);
and U13181 (N_13181,N_12108,N_12312);
nand U13182 (N_13182,N_12550,N_12017);
nor U13183 (N_13183,N_12681,N_12709);
or U13184 (N_13184,N_12123,N_12672);
or U13185 (N_13185,N_12648,N_12054);
nand U13186 (N_13186,N_12579,N_12594);
or U13187 (N_13187,N_12117,N_12653);
and U13188 (N_13188,N_12509,N_12543);
nor U13189 (N_13189,N_12720,N_12572);
and U13190 (N_13190,N_12730,N_12492);
nand U13191 (N_13191,N_12566,N_12593);
and U13192 (N_13192,N_12273,N_12062);
or U13193 (N_13193,N_12116,N_12709);
and U13194 (N_13194,N_12574,N_12630);
or U13195 (N_13195,N_12022,N_12337);
nor U13196 (N_13196,N_12222,N_12747);
or U13197 (N_13197,N_12279,N_12037);
nor U13198 (N_13198,N_12553,N_12450);
and U13199 (N_13199,N_12039,N_12551);
nor U13200 (N_13200,N_12282,N_12210);
nand U13201 (N_13201,N_12486,N_12362);
nor U13202 (N_13202,N_12221,N_12354);
nand U13203 (N_13203,N_12381,N_12280);
nand U13204 (N_13204,N_12018,N_12633);
and U13205 (N_13205,N_12651,N_12455);
nor U13206 (N_13206,N_12631,N_12622);
and U13207 (N_13207,N_12284,N_12552);
or U13208 (N_13208,N_12061,N_12190);
or U13209 (N_13209,N_12514,N_12719);
nand U13210 (N_13210,N_12208,N_12188);
nor U13211 (N_13211,N_12295,N_12746);
nand U13212 (N_13212,N_12347,N_12604);
and U13213 (N_13213,N_12578,N_12197);
nand U13214 (N_13214,N_12036,N_12406);
or U13215 (N_13215,N_12464,N_12185);
and U13216 (N_13216,N_12118,N_12366);
nor U13217 (N_13217,N_12651,N_12273);
nor U13218 (N_13218,N_12240,N_12059);
and U13219 (N_13219,N_12311,N_12409);
or U13220 (N_13220,N_12245,N_12691);
xor U13221 (N_13221,N_12370,N_12624);
nand U13222 (N_13222,N_12155,N_12643);
and U13223 (N_13223,N_12169,N_12417);
nor U13224 (N_13224,N_12548,N_12080);
nor U13225 (N_13225,N_12149,N_12111);
and U13226 (N_13226,N_12190,N_12488);
nor U13227 (N_13227,N_12334,N_12560);
xnor U13228 (N_13228,N_12658,N_12606);
nand U13229 (N_13229,N_12347,N_12067);
nand U13230 (N_13230,N_12640,N_12214);
nand U13231 (N_13231,N_12345,N_12492);
and U13232 (N_13232,N_12588,N_12099);
and U13233 (N_13233,N_12683,N_12213);
and U13234 (N_13234,N_12738,N_12687);
and U13235 (N_13235,N_12134,N_12190);
and U13236 (N_13236,N_12581,N_12136);
and U13237 (N_13237,N_12292,N_12253);
or U13238 (N_13238,N_12399,N_12289);
or U13239 (N_13239,N_12440,N_12234);
and U13240 (N_13240,N_12309,N_12673);
nor U13241 (N_13241,N_12694,N_12328);
nor U13242 (N_13242,N_12138,N_12403);
nor U13243 (N_13243,N_12739,N_12263);
or U13244 (N_13244,N_12711,N_12117);
and U13245 (N_13245,N_12420,N_12081);
nand U13246 (N_13246,N_12084,N_12112);
nand U13247 (N_13247,N_12202,N_12561);
and U13248 (N_13248,N_12199,N_12641);
and U13249 (N_13249,N_12120,N_12520);
or U13250 (N_13250,N_12533,N_12233);
nor U13251 (N_13251,N_12239,N_12613);
nor U13252 (N_13252,N_12041,N_12194);
and U13253 (N_13253,N_12032,N_12301);
nand U13254 (N_13254,N_12088,N_12450);
or U13255 (N_13255,N_12423,N_12656);
or U13256 (N_13256,N_12654,N_12381);
nor U13257 (N_13257,N_12246,N_12469);
nor U13258 (N_13258,N_12535,N_12590);
nor U13259 (N_13259,N_12223,N_12452);
and U13260 (N_13260,N_12107,N_12042);
nand U13261 (N_13261,N_12518,N_12198);
nor U13262 (N_13262,N_12508,N_12519);
xnor U13263 (N_13263,N_12694,N_12594);
or U13264 (N_13264,N_12072,N_12205);
nand U13265 (N_13265,N_12562,N_12117);
and U13266 (N_13266,N_12415,N_12607);
and U13267 (N_13267,N_12092,N_12727);
nor U13268 (N_13268,N_12197,N_12036);
and U13269 (N_13269,N_12111,N_12344);
or U13270 (N_13270,N_12535,N_12681);
or U13271 (N_13271,N_12127,N_12626);
nand U13272 (N_13272,N_12125,N_12274);
nand U13273 (N_13273,N_12209,N_12461);
nand U13274 (N_13274,N_12002,N_12462);
and U13275 (N_13275,N_12215,N_12450);
and U13276 (N_13276,N_12644,N_12663);
and U13277 (N_13277,N_12486,N_12161);
nor U13278 (N_13278,N_12641,N_12458);
and U13279 (N_13279,N_12501,N_12585);
nor U13280 (N_13280,N_12362,N_12391);
nand U13281 (N_13281,N_12352,N_12563);
nor U13282 (N_13282,N_12718,N_12407);
nor U13283 (N_13283,N_12101,N_12699);
and U13284 (N_13284,N_12635,N_12486);
or U13285 (N_13285,N_12711,N_12126);
or U13286 (N_13286,N_12465,N_12406);
nor U13287 (N_13287,N_12027,N_12302);
and U13288 (N_13288,N_12171,N_12163);
or U13289 (N_13289,N_12490,N_12683);
or U13290 (N_13290,N_12199,N_12152);
nor U13291 (N_13291,N_12714,N_12526);
or U13292 (N_13292,N_12705,N_12367);
nor U13293 (N_13293,N_12190,N_12644);
xor U13294 (N_13294,N_12160,N_12266);
nand U13295 (N_13295,N_12559,N_12680);
and U13296 (N_13296,N_12153,N_12425);
xnor U13297 (N_13297,N_12561,N_12260);
or U13298 (N_13298,N_12593,N_12502);
and U13299 (N_13299,N_12057,N_12687);
nor U13300 (N_13300,N_12409,N_12330);
nand U13301 (N_13301,N_12235,N_12084);
nand U13302 (N_13302,N_12411,N_12470);
nand U13303 (N_13303,N_12739,N_12324);
nand U13304 (N_13304,N_12320,N_12678);
xor U13305 (N_13305,N_12331,N_12063);
nand U13306 (N_13306,N_12332,N_12622);
and U13307 (N_13307,N_12440,N_12473);
nor U13308 (N_13308,N_12290,N_12507);
nor U13309 (N_13309,N_12395,N_12348);
and U13310 (N_13310,N_12514,N_12532);
or U13311 (N_13311,N_12187,N_12250);
and U13312 (N_13312,N_12352,N_12077);
nand U13313 (N_13313,N_12303,N_12724);
and U13314 (N_13314,N_12533,N_12084);
nor U13315 (N_13315,N_12597,N_12561);
nor U13316 (N_13316,N_12654,N_12194);
and U13317 (N_13317,N_12292,N_12645);
nand U13318 (N_13318,N_12239,N_12599);
nor U13319 (N_13319,N_12281,N_12720);
nor U13320 (N_13320,N_12478,N_12231);
nand U13321 (N_13321,N_12181,N_12613);
nor U13322 (N_13322,N_12493,N_12312);
nor U13323 (N_13323,N_12548,N_12652);
nor U13324 (N_13324,N_12287,N_12622);
nor U13325 (N_13325,N_12189,N_12603);
or U13326 (N_13326,N_12093,N_12226);
and U13327 (N_13327,N_12523,N_12018);
or U13328 (N_13328,N_12091,N_12637);
nand U13329 (N_13329,N_12384,N_12076);
and U13330 (N_13330,N_12284,N_12248);
or U13331 (N_13331,N_12657,N_12635);
nand U13332 (N_13332,N_12695,N_12290);
or U13333 (N_13333,N_12480,N_12492);
nand U13334 (N_13334,N_12033,N_12118);
nor U13335 (N_13335,N_12719,N_12466);
nand U13336 (N_13336,N_12155,N_12641);
nand U13337 (N_13337,N_12684,N_12312);
nand U13338 (N_13338,N_12277,N_12343);
and U13339 (N_13339,N_12456,N_12637);
nor U13340 (N_13340,N_12154,N_12452);
and U13341 (N_13341,N_12388,N_12304);
nand U13342 (N_13342,N_12706,N_12305);
and U13343 (N_13343,N_12483,N_12562);
or U13344 (N_13344,N_12354,N_12515);
nor U13345 (N_13345,N_12048,N_12538);
or U13346 (N_13346,N_12629,N_12380);
or U13347 (N_13347,N_12724,N_12169);
or U13348 (N_13348,N_12561,N_12453);
xor U13349 (N_13349,N_12226,N_12727);
nor U13350 (N_13350,N_12631,N_12399);
or U13351 (N_13351,N_12183,N_12551);
or U13352 (N_13352,N_12626,N_12261);
and U13353 (N_13353,N_12217,N_12288);
xnor U13354 (N_13354,N_12393,N_12652);
or U13355 (N_13355,N_12501,N_12710);
or U13356 (N_13356,N_12382,N_12183);
or U13357 (N_13357,N_12530,N_12014);
and U13358 (N_13358,N_12359,N_12095);
or U13359 (N_13359,N_12534,N_12525);
nor U13360 (N_13360,N_12637,N_12737);
nand U13361 (N_13361,N_12663,N_12631);
or U13362 (N_13362,N_12202,N_12073);
and U13363 (N_13363,N_12440,N_12384);
and U13364 (N_13364,N_12448,N_12698);
nor U13365 (N_13365,N_12454,N_12246);
and U13366 (N_13366,N_12430,N_12015);
or U13367 (N_13367,N_12575,N_12493);
or U13368 (N_13368,N_12090,N_12270);
nor U13369 (N_13369,N_12138,N_12185);
xnor U13370 (N_13370,N_12672,N_12038);
nor U13371 (N_13371,N_12250,N_12284);
nor U13372 (N_13372,N_12133,N_12104);
or U13373 (N_13373,N_12414,N_12158);
or U13374 (N_13374,N_12516,N_12403);
and U13375 (N_13375,N_12343,N_12581);
or U13376 (N_13376,N_12189,N_12740);
or U13377 (N_13377,N_12228,N_12467);
nor U13378 (N_13378,N_12095,N_12686);
and U13379 (N_13379,N_12096,N_12229);
nor U13380 (N_13380,N_12553,N_12106);
or U13381 (N_13381,N_12472,N_12694);
and U13382 (N_13382,N_12594,N_12017);
or U13383 (N_13383,N_12045,N_12365);
nor U13384 (N_13384,N_12111,N_12078);
nor U13385 (N_13385,N_12380,N_12005);
nand U13386 (N_13386,N_12064,N_12042);
nand U13387 (N_13387,N_12725,N_12191);
and U13388 (N_13388,N_12047,N_12721);
and U13389 (N_13389,N_12367,N_12550);
and U13390 (N_13390,N_12379,N_12456);
nand U13391 (N_13391,N_12532,N_12604);
nand U13392 (N_13392,N_12596,N_12667);
and U13393 (N_13393,N_12418,N_12703);
nor U13394 (N_13394,N_12748,N_12287);
or U13395 (N_13395,N_12487,N_12361);
nand U13396 (N_13396,N_12604,N_12618);
or U13397 (N_13397,N_12395,N_12109);
nand U13398 (N_13398,N_12201,N_12022);
or U13399 (N_13399,N_12103,N_12571);
nor U13400 (N_13400,N_12237,N_12572);
nor U13401 (N_13401,N_12645,N_12516);
nor U13402 (N_13402,N_12341,N_12649);
and U13403 (N_13403,N_12490,N_12545);
and U13404 (N_13404,N_12340,N_12588);
and U13405 (N_13405,N_12108,N_12262);
nor U13406 (N_13406,N_12224,N_12487);
and U13407 (N_13407,N_12352,N_12572);
or U13408 (N_13408,N_12075,N_12475);
nor U13409 (N_13409,N_12008,N_12744);
nor U13410 (N_13410,N_12594,N_12657);
nor U13411 (N_13411,N_12598,N_12431);
nand U13412 (N_13412,N_12455,N_12584);
nand U13413 (N_13413,N_12527,N_12269);
nand U13414 (N_13414,N_12495,N_12368);
xnor U13415 (N_13415,N_12111,N_12353);
nand U13416 (N_13416,N_12457,N_12564);
nor U13417 (N_13417,N_12094,N_12165);
or U13418 (N_13418,N_12472,N_12006);
and U13419 (N_13419,N_12553,N_12311);
nor U13420 (N_13420,N_12471,N_12158);
and U13421 (N_13421,N_12293,N_12233);
or U13422 (N_13422,N_12417,N_12495);
nand U13423 (N_13423,N_12694,N_12334);
or U13424 (N_13424,N_12511,N_12271);
or U13425 (N_13425,N_12511,N_12678);
and U13426 (N_13426,N_12005,N_12619);
or U13427 (N_13427,N_12649,N_12553);
nand U13428 (N_13428,N_12289,N_12463);
nor U13429 (N_13429,N_12635,N_12412);
nor U13430 (N_13430,N_12749,N_12109);
nand U13431 (N_13431,N_12642,N_12309);
and U13432 (N_13432,N_12291,N_12739);
or U13433 (N_13433,N_12262,N_12285);
nand U13434 (N_13434,N_12498,N_12603);
and U13435 (N_13435,N_12403,N_12632);
and U13436 (N_13436,N_12617,N_12207);
nand U13437 (N_13437,N_12050,N_12245);
and U13438 (N_13438,N_12514,N_12236);
nand U13439 (N_13439,N_12038,N_12336);
and U13440 (N_13440,N_12538,N_12731);
nor U13441 (N_13441,N_12400,N_12357);
or U13442 (N_13442,N_12082,N_12076);
nand U13443 (N_13443,N_12663,N_12345);
nor U13444 (N_13444,N_12036,N_12183);
nand U13445 (N_13445,N_12224,N_12172);
nor U13446 (N_13446,N_12657,N_12176);
and U13447 (N_13447,N_12565,N_12319);
nor U13448 (N_13448,N_12020,N_12700);
nand U13449 (N_13449,N_12171,N_12273);
or U13450 (N_13450,N_12292,N_12045);
nand U13451 (N_13451,N_12722,N_12160);
or U13452 (N_13452,N_12352,N_12156);
nand U13453 (N_13453,N_12452,N_12096);
nand U13454 (N_13454,N_12064,N_12695);
and U13455 (N_13455,N_12035,N_12609);
or U13456 (N_13456,N_12107,N_12483);
and U13457 (N_13457,N_12267,N_12611);
and U13458 (N_13458,N_12535,N_12127);
nor U13459 (N_13459,N_12697,N_12524);
or U13460 (N_13460,N_12316,N_12543);
nor U13461 (N_13461,N_12621,N_12324);
nand U13462 (N_13462,N_12485,N_12407);
or U13463 (N_13463,N_12168,N_12583);
or U13464 (N_13464,N_12650,N_12614);
nor U13465 (N_13465,N_12708,N_12376);
nand U13466 (N_13466,N_12360,N_12218);
and U13467 (N_13467,N_12046,N_12268);
nand U13468 (N_13468,N_12221,N_12288);
nor U13469 (N_13469,N_12390,N_12502);
and U13470 (N_13470,N_12183,N_12368);
nor U13471 (N_13471,N_12257,N_12572);
or U13472 (N_13472,N_12477,N_12547);
nor U13473 (N_13473,N_12594,N_12575);
and U13474 (N_13474,N_12523,N_12407);
and U13475 (N_13475,N_12718,N_12344);
nand U13476 (N_13476,N_12430,N_12054);
and U13477 (N_13477,N_12015,N_12573);
nand U13478 (N_13478,N_12620,N_12120);
nor U13479 (N_13479,N_12602,N_12044);
nand U13480 (N_13480,N_12498,N_12326);
and U13481 (N_13481,N_12207,N_12341);
nand U13482 (N_13482,N_12366,N_12245);
and U13483 (N_13483,N_12549,N_12338);
or U13484 (N_13484,N_12037,N_12449);
nand U13485 (N_13485,N_12110,N_12711);
nand U13486 (N_13486,N_12674,N_12378);
xnor U13487 (N_13487,N_12368,N_12325);
nor U13488 (N_13488,N_12459,N_12535);
and U13489 (N_13489,N_12580,N_12148);
and U13490 (N_13490,N_12488,N_12198);
nor U13491 (N_13491,N_12227,N_12289);
nor U13492 (N_13492,N_12682,N_12563);
nor U13493 (N_13493,N_12049,N_12521);
nand U13494 (N_13494,N_12301,N_12064);
or U13495 (N_13495,N_12398,N_12556);
nand U13496 (N_13496,N_12167,N_12404);
nand U13497 (N_13497,N_12183,N_12673);
and U13498 (N_13498,N_12192,N_12231);
and U13499 (N_13499,N_12012,N_12081);
nor U13500 (N_13500,N_13494,N_12995);
or U13501 (N_13501,N_13388,N_12966);
or U13502 (N_13502,N_12996,N_13176);
nand U13503 (N_13503,N_13138,N_13367);
and U13504 (N_13504,N_13072,N_13129);
or U13505 (N_13505,N_12949,N_12972);
nand U13506 (N_13506,N_12921,N_13147);
and U13507 (N_13507,N_12950,N_12779);
nor U13508 (N_13508,N_13317,N_13050);
nand U13509 (N_13509,N_12960,N_13068);
and U13510 (N_13510,N_13361,N_12870);
xor U13511 (N_13511,N_12862,N_13464);
or U13512 (N_13512,N_13121,N_12797);
nor U13513 (N_13513,N_13160,N_12982);
nor U13514 (N_13514,N_13302,N_13360);
and U13515 (N_13515,N_12992,N_13233);
nor U13516 (N_13516,N_13287,N_13220);
or U13517 (N_13517,N_13093,N_13470);
and U13518 (N_13518,N_13208,N_13135);
nor U13519 (N_13519,N_12787,N_13276);
or U13520 (N_13520,N_12910,N_12917);
and U13521 (N_13521,N_13019,N_13338);
or U13522 (N_13522,N_13458,N_13422);
nand U13523 (N_13523,N_12984,N_13178);
and U13524 (N_13524,N_12845,N_13217);
and U13525 (N_13525,N_13001,N_12867);
or U13526 (N_13526,N_13474,N_12963);
nor U13527 (N_13527,N_12844,N_13359);
nor U13528 (N_13528,N_13188,N_13164);
xnor U13529 (N_13529,N_13061,N_13415);
or U13530 (N_13530,N_13163,N_13099);
nand U13531 (N_13531,N_13023,N_13230);
nor U13532 (N_13532,N_12881,N_13288);
nor U13533 (N_13533,N_12926,N_13394);
nand U13534 (N_13534,N_13169,N_13312);
or U13535 (N_13535,N_12800,N_13268);
nand U13536 (N_13536,N_13213,N_13381);
or U13537 (N_13537,N_13095,N_12761);
nand U13538 (N_13538,N_13335,N_12752);
and U13539 (N_13539,N_13366,N_13244);
and U13540 (N_13540,N_12836,N_13401);
nand U13541 (N_13541,N_13145,N_13227);
nor U13542 (N_13542,N_13106,N_12994);
or U13543 (N_13543,N_13278,N_13232);
xnor U13544 (N_13544,N_12915,N_13175);
nor U13545 (N_13545,N_13140,N_12932);
nor U13546 (N_13546,N_12876,N_13168);
or U13547 (N_13547,N_12883,N_13329);
xor U13548 (N_13548,N_13075,N_12802);
or U13549 (N_13549,N_13300,N_13431);
and U13550 (N_13550,N_13081,N_13310);
and U13551 (N_13551,N_13391,N_12942);
or U13552 (N_13552,N_13284,N_13141);
or U13553 (N_13553,N_12891,N_13030);
nor U13554 (N_13554,N_12771,N_12773);
nand U13555 (N_13555,N_13127,N_13405);
nor U13556 (N_13556,N_12998,N_13286);
nor U13557 (N_13557,N_13441,N_13451);
nor U13558 (N_13558,N_12894,N_12803);
nand U13559 (N_13559,N_13013,N_13454);
nand U13560 (N_13560,N_12853,N_12916);
or U13561 (N_13561,N_13117,N_12945);
and U13562 (N_13562,N_12871,N_13444);
nor U13563 (N_13563,N_13457,N_13209);
or U13564 (N_13564,N_12946,N_13442);
nor U13565 (N_13565,N_13222,N_12880);
and U13566 (N_13566,N_12959,N_13488);
and U13567 (N_13567,N_13231,N_12772);
or U13568 (N_13568,N_13341,N_13396);
or U13569 (N_13569,N_12987,N_12830);
and U13570 (N_13570,N_13150,N_12792);
and U13571 (N_13571,N_12937,N_13468);
nand U13572 (N_13572,N_12850,N_13151);
or U13573 (N_13573,N_13314,N_13449);
and U13574 (N_13574,N_13346,N_13065);
nand U13575 (N_13575,N_13301,N_13035);
and U13576 (N_13576,N_13193,N_12923);
nor U13577 (N_13577,N_13331,N_13434);
nand U13578 (N_13578,N_13161,N_12939);
and U13579 (N_13579,N_13012,N_12912);
and U13580 (N_13580,N_13290,N_13328);
nor U13581 (N_13581,N_13408,N_13097);
nor U13582 (N_13582,N_13192,N_13320);
and U13583 (N_13583,N_13461,N_12753);
nor U13584 (N_13584,N_12885,N_13111);
nor U13585 (N_13585,N_12927,N_12914);
nor U13586 (N_13586,N_12857,N_13271);
and U13587 (N_13587,N_12825,N_13297);
nand U13588 (N_13588,N_13223,N_13282);
nor U13589 (N_13589,N_13045,N_13113);
nor U13590 (N_13590,N_13028,N_13060);
and U13591 (N_13591,N_12962,N_12813);
or U13592 (N_13592,N_13390,N_13191);
and U13593 (N_13593,N_13294,N_13203);
nor U13594 (N_13594,N_13197,N_12934);
nor U13595 (N_13595,N_13033,N_13283);
and U13596 (N_13596,N_13275,N_13265);
nor U13597 (N_13597,N_12971,N_13246);
nand U13598 (N_13598,N_13462,N_13272);
nor U13599 (N_13599,N_12888,N_13003);
nand U13600 (N_13600,N_13376,N_13166);
nor U13601 (N_13601,N_12837,N_13085);
and U13602 (N_13602,N_13477,N_13206);
nor U13603 (N_13603,N_13031,N_13254);
or U13604 (N_13604,N_12865,N_13108);
nor U13605 (N_13605,N_12806,N_12955);
and U13606 (N_13606,N_13309,N_13103);
or U13607 (N_13607,N_13256,N_12847);
nor U13608 (N_13608,N_13148,N_13403);
and U13609 (N_13609,N_13435,N_13353);
xnor U13610 (N_13610,N_13295,N_13006);
and U13611 (N_13611,N_12933,N_13364);
nor U13612 (N_13612,N_12755,N_13267);
and U13613 (N_13613,N_12819,N_12811);
and U13614 (N_13614,N_13427,N_13445);
nand U13615 (N_13615,N_13032,N_13443);
or U13616 (N_13616,N_12775,N_12935);
nor U13617 (N_13617,N_13305,N_13102);
and U13618 (N_13618,N_13260,N_12849);
nor U13619 (N_13619,N_12970,N_12941);
nand U13620 (N_13620,N_12790,N_13333);
and U13621 (N_13621,N_13262,N_13101);
and U13622 (N_13622,N_12983,N_13096);
xnor U13623 (N_13623,N_13253,N_13411);
nor U13624 (N_13624,N_13429,N_13195);
or U13625 (N_13625,N_12873,N_13387);
nor U13626 (N_13626,N_13397,N_13071);
nor U13627 (N_13627,N_13481,N_13414);
nand U13628 (N_13628,N_13067,N_13484);
nand U13629 (N_13629,N_13123,N_12986);
nand U13630 (N_13630,N_13077,N_13257);
and U13631 (N_13631,N_13418,N_13384);
and U13632 (N_13632,N_12879,N_13053);
nor U13633 (N_13633,N_12897,N_13172);
nand U13634 (N_13634,N_12760,N_12788);
nor U13635 (N_13635,N_13303,N_12777);
nand U13636 (N_13636,N_13412,N_12889);
nor U13637 (N_13637,N_12785,N_12979);
and U13638 (N_13638,N_12877,N_13018);
or U13639 (N_13639,N_13348,N_12791);
or U13640 (N_13640,N_12991,N_13363);
and U13641 (N_13641,N_13465,N_13498);
nand U13642 (N_13642,N_12750,N_13337);
or U13643 (N_13643,N_13450,N_13466);
nand U13644 (N_13644,N_13350,N_13090);
or U13645 (N_13645,N_13002,N_13351);
and U13646 (N_13646,N_12816,N_13385);
or U13647 (N_13647,N_12776,N_13142);
nor U13648 (N_13648,N_12913,N_12833);
nand U13649 (N_13649,N_13467,N_13460);
or U13650 (N_13650,N_13110,N_13228);
and U13651 (N_13651,N_13034,N_13428);
nand U13652 (N_13652,N_13130,N_13298);
and U13653 (N_13653,N_13378,N_13089);
nand U13654 (N_13654,N_12920,N_12809);
or U13655 (N_13655,N_13119,N_13311);
nand U13656 (N_13656,N_12938,N_12922);
nand U13657 (N_13657,N_13196,N_12956);
nand U13658 (N_13658,N_12975,N_12969);
and U13659 (N_13659,N_13029,N_13218);
or U13660 (N_13660,N_13436,N_12804);
nand U13661 (N_13661,N_12884,N_12954);
or U13662 (N_13662,N_13291,N_13400);
and U13663 (N_13663,N_12909,N_12848);
nand U13664 (N_13664,N_13373,N_13125);
or U13665 (N_13665,N_12856,N_12821);
and U13666 (N_13666,N_13183,N_13432);
nand U13667 (N_13667,N_12842,N_13389);
and U13668 (N_13668,N_13149,N_13369);
nand U13669 (N_13669,N_13368,N_13371);
nor U13670 (N_13670,N_13440,N_13332);
nor U13671 (N_13671,N_13027,N_13413);
xnor U13672 (N_13672,N_13010,N_13330);
and U13673 (N_13673,N_12908,N_13198);
nand U13674 (N_13674,N_12965,N_12762);
nand U13675 (N_13675,N_12798,N_13008);
or U13676 (N_13676,N_12823,N_13046);
xor U13677 (N_13677,N_13308,N_13316);
nand U13678 (N_13678,N_13358,N_12808);
or U13679 (N_13679,N_12858,N_13062);
nor U13680 (N_13680,N_13041,N_12756);
or U13681 (N_13681,N_12905,N_12812);
or U13682 (N_13682,N_13181,N_13370);
nor U13683 (N_13683,N_12895,N_13237);
or U13684 (N_13684,N_13025,N_12989);
nand U13685 (N_13685,N_13423,N_13327);
nand U13686 (N_13686,N_13162,N_13105);
nand U13687 (N_13687,N_13069,N_12831);
nor U13688 (N_13688,N_13115,N_13490);
and U13689 (N_13689,N_13448,N_13107);
nand U13690 (N_13690,N_12974,N_13251);
nor U13691 (N_13691,N_13352,N_13374);
nor U13692 (N_13692,N_13021,N_13236);
or U13693 (N_13693,N_13354,N_13070);
or U13694 (N_13694,N_13334,N_12943);
nor U13695 (N_13695,N_13205,N_13165);
nor U13696 (N_13696,N_13094,N_12826);
nand U13697 (N_13697,N_13372,N_13009);
or U13698 (N_13698,N_13489,N_13049);
or U13699 (N_13699,N_13395,N_13005);
nand U13700 (N_13700,N_12968,N_13190);
nor U13701 (N_13701,N_13098,N_12861);
and U13702 (N_13702,N_13215,N_13024);
and U13703 (N_13703,N_12952,N_13000);
nor U13704 (N_13704,N_13425,N_13296);
and U13705 (N_13705,N_13120,N_12774);
or U13706 (N_13706,N_13132,N_12864);
nand U13707 (N_13707,N_13247,N_13078);
or U13708 (N_13708,N_13326,N_13088);
nand U13709 (N_13709,N_13473,N_13037);
or U13710 (N_13710,N_12841,N_13185);
or U13711 (N_13711,N_13083,N_13076);
nand U13712 (N_13712,N_13420,N_13261);
or U13713 (N_13713,N_13020,N_13365);
and U13714 (N_13714,N_13289,N_12789);
or U13715 (N_13715,N_13048,N_12782);
or U13716 (N_13716,N_12948,N_13017);
nor U13717 (N_13717,N_13134,N_12817);
and U13718 (N_13718,N_13421,N_12754);
nor U13719 (N_13719,N_12928,N_12758);
nor U13720 (N_13720,N_13323,N_12786);
or U13721 (N_13721,N_12799,N_13402);
and U13722 (N_13722,N_13259,N_12824);
nand U13723 (N_13723,N_13211,N_13056);
or U13724 (N_13724,N_13124,N_12957);
or U13725 (N_13725,N_13340,N_13398);
nand U13726 (N_13726,N_12770,N_12818);
and U13727 (N_13727,N_12796,N_13495);
nand U13728 (N_13728,N_13399,N_12902);
or U13729 (N_13729,N_13362,N_13249);
or U13730 (N_13730,N_13144,N_12784);
nor U13731 (N_13731,N_13128,N_13255);
and U13732 (N_13732,N_13199,N_12794);
or U13733 (N_13733,N_12924,N_13375);
or U13734 (N_13734,N_13281,N_13383);
or U13735 (N_13735,N_13382,N_12985);
or U13736 (N_13736,N_13040,N_12906);
nor U13737 (N_13737,N_13344,N_13492);
nor U13738 (N_13738,N_13409,N_13219);
or U13739 (N_13739,N_13379,N_13476);
nand U13740 (N_13740,N_13136,N_13258);
and U13741 (N_13741,N_13216,N_13349);
or U13742 (N_13742,N_13059,N_12901);
nand U13743 (N_13743,N_13245,N_12820);
and U13744 (N_13744,N_13240,N_13453);
and U13745 (N_13745,N_13250,N_13235);
xor U13746 (N_13746,N_12840,N_12827);
nand U13747 (N_13747,N_12993,N_13226);
or U13748 (N_13748,N_13055,N_13437);
nand U13749 (N_13749,N_12835,N_13064);
xor U13750 (N_13750,N_12999,N_13377);
or U13751 (N_13751,N_12810,N_13225);
nor U13752 (N_13752,N_13118,N_13480);
nor U13753 (N_13753,N_13043,N_12887);
and U13754 (N_13754,N_12757,N_13022);
nor U13755 (N_13755,N_12838,N_13322);
nor U13756 (N_13756,N_13154,N_13343);
nand U13757 (N_13757,N_13086,N_12763);
and U13758 (N_13758,N_12832,N_13357);
xor U13759 (N_13759,N_12859,N_13189);
nor U13760 (N_13760,N_13447,N_13293);
and U13761 (N_13761,N_13347,N_13184);
or U13762 (N_13762,N_13285,N_13011);
xnor U13763 (N_13763,N_13242,N_13221);
nor U13764 (N_13764,N_13380,N_13496);
or U13765 (N_13765,N_13292,N_13194);
nand U13766 (N_13766,N_13252,N_13100);
nor U13767 (N_13767,N_13084,N_13167);
nand U13768 (N_13768,N_13336,N_12919);
nand U13769 (N_13769,N_13455,N_13015);
or U13770 (N_13770,N_13315,N_12815);
or U13771 (N_13771,N_13073,N_12843);
or U13772 (N_13772,N_13277,N_13407);
and U13773 (N_13773,N_13430,N_13321);
and U13774 (N_13774,N_12769,N_12958);
nand U13775 (N_13775,N_13171,N_12766);
nor U13776 (N_13776,N_13463,N_13116);
nand U13777 (N_13777,N_13087,N_13438);
or U13778 (N_13778,N_12767,N_13109);
nor U13779 (N_13779,N_12860,N_12961);
nand U13780 (N_13780,N_13174,N_13016);
xnor U13781 (N_13781,N_12869,N_13180);
nor U13782 (N_13782,N_12855,N_12977);
nand U13783 (N_13783,N_12997,N_12973);
or U13784 (N_13784,N_13306,N_13146);
nor U13785 (N_13785,N_13269,N_12793);
nand U13786 (N_13786,N_13497,N_13241);
and U13787 (N_13787,N_12990,N_13325);
or U13788 (N_13788,N_13313,N_13419);
or U13789 (N_13789,N_13133,N_13047);
nor U13790 (N_13790,N_13186,N_13273);
nand U13791 (N_13791,N_12846,N_12911);
and U13792 (N_13792,N_12768,N_13386);
xor U13793 (N_13793,N_13092,N_13339);
nand U13794 (N_13794,N_13263,N_12978);
nor U13795 (N_13795,N_13446,N_13173);
nand U13796 (N_13796,N_13479,N_13342);
nor U13797 (N_13797,N_12900,N_13157);
or U13798 (N_13798,N_13091,N_12903);
nand U13799 (N_13799,N_13248,N_13299);
nand U13800 (N_13800,N_12801,N_12807);
and U13801 (N_13801,N_12783,N_12890);
and U13802 (N_13802,N_13318,N_13439);
nand U13803 (N_13803,N_13239,N_13424);
nor U13804 (N_13804,N_12765,N_13036);
nand U13805 (N_13805,N_13417,N_13229);
nand U13806 (N_13806,N_13044,N_13304);
or U13807 (N_13807,N_13074,N_13014);
and U13808 (N_13808,N_13319,N_13416);
and U13809 (N_13809,N_13426,N_13042);
or U13810 (N_13810,N_13122,N_13404);
nor U13811 (N_13811,N_13212,N_13410);
or U13812 (N_13812,N_13210,N_12834);
or U13813 (N_13813,N_12872,N_13112);
and U13814 (N_13814,N_13038,N_13406);
nor U13815 (N_13815,N_13224,N_13079);
nor U13816 (N_13816,N_12795,N_12878);
or U13817 (N_13817,N_13131,N_12851);
and U13818 (N_13818,N_13052,N_12947);
nor U13819 (N_13819,N_12780,N_12866);
and U13820 (N_13820,N_13039,N_12918);
nor U13821 (N_13821,N_13080,N_13007);
and U13822 (N_13822,N_12898,N_13177);
or U13823 (N_13823,N_13472,N_12967);
nand U13824 (N_13824,N_13307,N_13114);
or U13825 (N_13825,N_12863,N_13170);
nor U13826 (N_13826,N_13475,N_13026);
and U13827 (N_13827,N_12781,N_13202);
nand U13828 (N_13828,N_13187,N_13280);
nor U13829 (N_13829,N_12829,N_13126);
nand U13830 (N_13830,N_13485,N_13139);
nor U13831 (N_13831,N_12778,N_13469);
nor U13832 (N_13832,N_12852,N_12976);
nand U13833 (N_13833,N_12764,N_13264);
and U13834 (N_13834,N_13324,N_13471);
nand U13835 (N_13835,N_12981,N_12899);
and U13836 (N_13836,N_12875,N_13058);
xor U13837 (N_13837,N_13478,N_13156);
and U13838 (N_13838,N_13355,N_13159);
and U13839 (N_13839,N_12839,N_13456);
or U13840 (N_13840,N_13207,N_13392);
nand U13841 (N_13841,N_13345,N_13243);
nand U13842 (N_13842,N_13158,N_12980);
or U13843 (N_13843,N_13066,N_13499);
or U13844 (N_13844,N_13486,N_12882);
and U13845 (N_13845,N_13054,N_13266);
nand U13846 (N_13846,N_13491,N_13459);
or U13847 (N_13847,N_13487,N_13057);
or U13848 (N_13848,N_12893,N_12944);
nor U13849 (N_13849,N_13051,N_12751);
or U13850 (N_13850,N_13153,N_12904);
xor U13851 (N_13851,N_13063,N_13274);
nand U13852 (N_13852,N_12925,N_13152);
or U13853 (N_13853,N_13482,N_13433);
or U13854 (N_13854,N_13356,N_13234);
nor U13855 (N_13855,N_12886,N_12929);
or U13856 (N_13856,N_13155,N_13179);
and U13857 (N_13857,N_12854,N_12951);
and U13858 (N_13858,N_13204,N_12828);
nand U13859 (N_13859,N_13270,N_13279);
xnor U13860 (N_13860,N_12822,N_12759);
xnor U13861 (N_13861,N_12964,N_13393);
nor U13862 (N_13862,N_12896,N_12892);
nor U13863 (N_13863,N_13200,N_13182);
and U13864 (N_13864,N_12931,N_12953);
nor U13865 (N_13865,N_13214,N_13493);
and U13866 (N_13866,N_13238,N_13082);
or U13867 (N_13867,N_13143,N_12988);
nand U13868 (N_13868,N_13452,N_13004);
and U13869 (N_13869,N_12874,N_12930);
nor U13870 (N_13870,N_12907,N_13104);
or U13871 (N_13871,N_13137,N_12868);
nor U13872 (N_13872,N_13201,N_13483);
nor U13873 (N_13873,N_12814,N_12940);
and U13874 (N_13874,N_12805,N_12936);
nand U13875 (N_13875,N_12857,N_13138);
nand U13876 (N_13876,N_13017,N_13295);
nand U13877 (N_13877,N_12763,N_12828);
nor U13878 (N_13878,N_12986,N_12772);
nand U13879 (N_13879,N_13360,N_13316);
and U13880 (N_13880,N_13162,N_13138);
and U13881 (N_13881,N_13291,N_12823);
and U13882 (N_13882,N_13010,N_12932);
or U13883 (N_13883,N_13216,N_13259);
xnor U13884 (N_13884,N_13306,N_12904);
nand U13885 (N_13885,N_13016,N_13366);
xnor U13886 (N_13886,N_13422,N_13086);
nor U13887 (N_13887,N_13492,N_12828);
nor U13888 (N_13888,N_13132,N_13217);
nor U13889 (N_13889,N_13364,N_13224);
and U13890 (N_13890,N_13169,N_12828);
nor U13891 (N_13891,N_13422,N_12981);
nand U13892 (N_13892,N_13274,N_12827);
nand U13893 (N_13893,N_12795,N_12903);
nor U13894 (N_13894,N_13212,N_13181);
nand U13895 (N_13895,N_13207,N_13256);
or U13896 (N_13896,N_12984,N_13094);
and U13897 (N_13897,N_13394,N_13319);
nor U13898 (N_13898,N_13232,N_12846);
or U13899 (N_13899,N_13445,N_13022);
or U13900 (N_13900,N_12761,N_13171);
nand U13901 (N_13901,N_12918,N_12799);
or U13902 (N_13902,N_12852,N_13371);
or U13903 (N_13903,N_13133,N_13166);
and U13904 (N_13904,N_12783,N_13228);
or U13905 (N_13905,N_12849,N_12880);
nand U13906 (N_13906,N_12918,N_12854);
or U13907 (N_13907,N_13077,N_12901);
and U13908 (N_13908,N_12832,N_12845);
and U13909 (N_13909,N_13079,N_13294);
nand U13910 (N_13910,N_13296,N_13082);
nand U13911 (N_13911,N_12786,N_13402);
nand U13912 (N_13912,N_13366,N_13175);
or U13913 (N_13913,N_12779,N_12963);
and U13914 (N_13914,N_13351,N_13302);
and U13915 (N_13915,N_13216,N_13245);
or U13916 (N_13916,N_13338,N_13288);
nor U13917 (N_13917,N_13367,N_13389);
nor U13918 (N_13918,N_13013,N_13378);
and U13919 (N_13919,N_13395,N_13317);
or U13920 (N_13920,N_12934,N_13489);
nor U13921 (N_13921,N_12819,N_12929);
or U13922 (N_13922,N_13446,N_13221);
and U13923 (N_13923,N_12978,N_12823);
and U13924 (N_13924,N_13364,N_12951);
or U13925 (N_13925,N_13410,N_12999);
nand U13926 (N_13926,N_12917,N_12948);
and U13927 (N_13927,N_13494,N_13498);
or U13928 (N_13928,N_13299,N_13100);
or U13929 (N_13929,N_13146,N_13427);
nand U13930 (N_13930,N_13447,N_13263);
and U13931 (N_13931,N_13028,N_12883);
nor U13932 (N_13932,N_13253,N_13073);
nand U13933 (N_13933,N_13212,N_13032);
or U13934 (N_13934,N_13169,N_12881);
nor U13935 (N_13935,N_13259,N_12902);
or U13936 (N_13936,N_12926,N_13408);
nand U13937 (N_13937,N_13432,N_13202);
or U13938 (N_13938,N_13242,N_13012);
nor U13939 (N_13939,N_12962,N_13100);
or U13940 (N_13940,N_12968,N_13351);
nor U13941 (N_13941,N_13335,N_13299);
and U13942 (N_13942,N_12909,N_13096);
or U13943 (N_13943,N_13151,N_13079);
nor U13944 (N_13944,N_13044,N_13192);
xnor U13945 (N_13945,N_12905,N_12917);
nand U13946 (N_13946,N_12849,N_13467);
and U13947 (N_13947,N_13006,N_13300);
or U13948 (N_13948,N_13438,N_12770);
or U13949 (N_13949,N_13295,N_13388);
or U13950 (N_13950,N_12923,N_13024);
nor U13951 (N_13951,N_13050,N_13238);
or U13952 (N_13952,N_13341,N_12970);
or U13953 (N_13953,N_13035,N_12824);
and U13954 (N_13954,N_13285,N_13274);
nand U13955 (N_13955,N_13134,N_13243);
nand U13956 (N_13956,N_13465,N_13101);
and U13957 (N_13957,N_13188,N_12830);
nor U13958 (N_13958,N_13161,N_12973);
or U13959 (N_13959,N_12830,N_13352);
and U13960 (N_13960,N_13301,N_13432);
nor U13961 (N_13961,N_13246,N_13187);
and U13962 (N_13962,N_13028,N_13042);
and U13963 (N_13963,N_13497,N_13426);
and U13964 (N_13964,N_13475,N_13104);
and U13965 (N_13965,N_12877,N_12932);
and U13966 (N_13966,N_13418,N_12861);
nand U13967 (N_13967,N_13091,N_13023);
and U13968 (N_13968,N_13345,N_12982);
and U13969 (N_13969,N_13024,N_13095);
nor U13970 (N_13970,N_13079,N_13278);
and U13971 (N_13971,N_13224,N_12967);
or U13972 (N_13972,N_13050,N_13192);
or U13973 (N_13973,N_13467,N_13423);
and U13974 (N_13974,N_13329,N_12852);
or U13975 (N_13975,N_13022,N_13441);
or U13976 (N_13976,N_13232,N_13335);
or U13977 (N_13977,N_12812,N_13464);
nor U13978 (N_13978,N_12832,N_12771);
or U13979 (N_13979,N_13134,N_12965);
nor U13980 (N_13980,N_13052,N_13120);
and U13981 (N_13981,N_12940,N_13164);
nand U13982 (N_13982,N_12991,N_12891);
nor U13983 (N_13983,N_13234,N_12791);
or U13984 (N_13984,N_13491,N_13476);
nand U13985 (N_13985,N_13467,N_12832);
nor U13986 (N_13986,N_12813,N_13113);
and U13987 (N_13987,N_13175,N_12993);
nand U13988 (N_13988,N_13282,N_13499);
nand U13989 (N_13989,N_13134,N_13152);
xnor U13990 (N_13990,N_12934,N_13256);
nor U13991 (N_13991,N_13067,N_13066);
or U13992 (N_13992,N_13118,N_13001);
and U13993 (N_13993,N_13135,N_13233);
or U13994 (N_13994,N_13474,N_12990);
and U13995 (N_13995,N_13358,N_13360);
or U13996 (N_13996,N_13309,N_12853);
and U13997 (N_13997,N_13374,N_13345);
and U13998 (N_13998,N_12929,N_13147);
nand U13999 (N_13999,N_13412,N_13491);
nor U14000 (N_14000,N_13261,N_13342);
or U14001 (N_14001,N_13268,N_12867);
nor U14002 (N_14002,N_12854,N_13083);
and U14003 (N_14003,N_12891,N_13211);
nor U14004 (N_14004,N_13144,N_13274);
and U14005 (N_14005,N_13060,N_12905);
and U14006 (N_14006,N_13321,N_12859);
nand U14007 (N_14007,N_13129,N_13268);
or U14008 (N_14008,N_13193,N_13020);
or U14009 (N_14009,N_13496,N_12935);
or U14010 (N_14010,N_13415,N_13224);
nand U14011 (N_14011,N_12845,N_13000);
nor U14012 (N_14012,N_12777,N_12926);
nand U14013 (N_14013,N_12813,N_13123);
or U14014 (N_14014,N_12766,N_13335);
nand U14015 (N_14015,N_13329,N_13323);
nor U14016 (N_14016,N_12982,N_13346);
nand U14017 (N_14017,N_13226,N_12884);
or U14018 (N_14018,N_13244,N_13254);
nor U14019 (N_14019,N_13242,N_12915);
nand U14020 (N_14020,N_12900,N_12838);
and U14021 (N_14021,N_13468,N_13143);
and U14022 (N_14022,N_13289,N_12754);
or U14023 (N_14023,N_12841,N_12958);
nand U14024 (N_14024,N_13024,N_13088);
and U14025 (N_14025,N_13409,N_13066);
and U14026 (N_14026,N_12841,N_13087);
or U14027 (N_14027,N_13320,N_12859);
or U14028 (N_14028,N_13085,N_13037);
nand U14029 (N_14029,N_12826,N_13022);
nor U14030 (N_14030,N_13031,N_12834);
nand U14031 (N_14031,N_13085,N_13341);
or U14032 (N_14032,N_13095,N_13424);
nor U14033 (N_14033,N_13100,N_13006);
nand U14034 (N_14034,N_13156,N_13498);
and U14035 (N_14035,N_13359,N_12884);
nand U14036 (N_14036,N_13478,N_12880);
nor U14037 (N_14037,N_12801,N_13120);
or U14038 (N_14038,N_13126,N_13358);
nor U14039 (N_14039,N_13180,N_13311);
nor U14040 (N_14040,N_13215,N_13201);
and U14041 (N_14041,N_12940,N_13201);
nand U14042 (N_14042,N_12947,N_13455);
nand U14043 (N_14043,N_13460,N_13447);
or U14044 (N_14044,N_13393,N_12865);
or U14045 (N_14045,N_13172,N_13232);
nor U14046 (N_14046,N_13078,N_12856);
nand U14047 (N_14047,N_13293,N_13028);
nand U14048 (N_14048,N_13085,N_13300);
or U14049 (N_14049,N_13294,N_13069);
or U14050 (N_14050,N_13266,N_13308);
nand U14051 (N_14051,N_12846,N_13479);
nand U14052 (N_14052,N_12899,N_12971);
and U14053 (N_14053,N_13264,N_13349);
nor U14054 (N_14054,N_13263,N_13383);
nor U14055 (N_14055,N_13132,N_13403);
nor U14056 (N_14056,N_12909,N_13109);
or U14057 (N_14057,N_12939,N_13497);
xor U14058 (N_14058,N_13402,N_13358);
nand U14059 (N_14059,N_13311,N_12817);
or U14060 (N_14060,N_13289,N_13174);
or U14061 (N_14061,N_13247,N_13108);
nand U14062 (N_14062,N_12828,N_13167);
nor U14063 (N_14063,N_13179,N_13008);
nand U14064 (N_14064,N_13318,N_12850);
nor U14065 (N_14065,N_13417,N_13032);
xor U14066 (N_14066,N_12981,N_13147);
and U14067 (N_14067,N_13289,N_12797);
and U14068 (N_14068,N_13114,N_13392);
and U14069 (N_14069,N_13302,N_12893);
and U14070 (N_14070,N_13216,N_13398);
nand U14071 (N_14071,N_13005,N_13150);
nor U14072 (N_14072,N_12954,N_12893);
nand U14073 (N_14073,N_12962,N_13229);
nand U14074 (N_14074,N_13391,N_13349);
nor U14075 (N_14075,N_12806,N_12799);
or U14076 (N_14076,N_13092,N_13444);
nand U14077 (N_14077,N_12829,N_13129);
or U14078 (N_14078,N_13430,N_12771);
or U14079 (N_14079,N_12768,N_13277);
nor U14080 (N_14080,N_13192,N_13181);
or U14081 (N_14081,N_12940,N_12795);
and U14082 (N_14082,N_12839,N_13335);
nand U14083 (N_14083,N_12954,N_13139);
and U14084 (N_14084,N_13233,N_12938);
and U14085 (N_14085,N_13042,N_13379);
nor U14086 (N_14086,N_13245,N_12854);
nor U14087 (N_14087,N_13207,N_13467);
or U14088 (N_14088,N_13045,N_12845);
nor U14089 (N_14089,N_13148,N_12841);
and U14090 (N_14090,N_13019,N_13092);
nand U14091 (N_14091,N_12866,N_13197);
nand U14092 (N_14092,N_13085,N_12816);
nand U14093 (N_14093,N_13098,N_13158);
nand U14094 (N_14094,N_12876,N_12954);
or U14095 (N_14095,N_12777,N_12804);
or U14096 (N_14096,N_13435,N_12938);
nor U14097 (N_14097,N_13235,N_13315);
nand U14098 (N_14098,N_13227,N_13412);
nor U14099 (N_14099,N_12762,N_12955);
nor U14100 (N_14100,N_13287,N_13203);
or U14101 (N_14101,N_13457,N_13424);
nand U14102 (N_14102,N_13342,N_13280);
and U14103 (N_14103,N_12837,N_12776);
and U14104 (N_14104,N_13438,N_12989);
nor U14105 (N_14105,N_13360,N_13010);
nor U14106 (N_14106,N_12777,N_13389);
nand U14107 (N_14107,N_13070,N_13306);
or U14108 (N_14108,N_12990,N_13446);
nor U14109 (N_14109,N_13040,N_13427);
nand U14110 (N_14110,N_12940,N_13321);
or U14111 (N_14111,N_13318,N_13486);
and U14112 (N_14112,N_13488,N_13456);
nand U14113 (N_14113,N_12877,N_12977);
xor U14114 (N_14114,N_13447,N_13440);
or U14115 (N_14115,N_13107,N_12855);
nor U14116 (N_14116,N_13449,N_13481);
nand U14117 (N_14117,N_13283,N_13157);
nand U14118 (N_14118,N_12956,N_12871);
nand U14119 (N_14119,N_12763,N_13345);
xnor U14120 (N_14120,N_12870,N_13243);
and U14121 (N_14121,N_13161,N_12985);
and U14122 (N_14122,N_13471,N_13142);
and U14123 (N_14123,N_12820,N_13422);
or U14124 (N_14124,N_13120,N_12928);
and U14125 (N_14125,N_13197,N_13115);
nand U14126 (N_14126,N_13151,N_13242);
nor U14127 (N_14127,N_13414,N_13231);
nand U14128 (N_14128,N_12783,N_12958);
and U14129 (N_14129,N_13446,N_12994);
nor U14130 (N_14130,N_13266,N_12878);
nand U14131 (N_14131,N_13230,N_12934);
nand U14132 (N_14132,N_13202,N_12888);
or U14133 (N_14133,N_12933,N_12878);
nor U14134 (N_14134,N_13018,N_13308);
nor U14135 (N_14135,N_13376,N_13467);
or U14136 (N_14136,N_12952,N_13362);
or U14137 (N_14137,N_13392,N_13337);
nand U14138 (N_14138,N_12786,N_12761);
xor U14139 (N_14139,N_12845,N_13067);
nand U14140 (N_14140,N_13145,N_13264);
and U14141 (N_14141,N_12921,N_13069);
nand U14142 (N_14142,N_13405,N_13178);
and U14143 (N_14143,N_13451,N_13252);
nor U14144 (N_14144,N_12826,N_13364);
and U14145 (N_14145,N_13210,N_13207);
or U14146 (N_14146,N_12821,N_13376);
nand U14147 (N_14147,N_12903,N_13416);
nor U14148 (N_14148,N_13230,N_13279);
nor U14149 (N_14149,N_13184,N_13091);
nand U14150 (N_14150,N_12812,N_13321);
nor U14151 (N_14151,N_13340,N_13232);
or U14152 (N_14152,N_13178,N_13461);
and U14153 (N_14153,N_12943,N_12780);
nand U14154 (N_14154,N_12907,N_13396);
xor U14155 (N_14155,N_13333,N_13410);
nor U14156 (N_14156,N_12828,N_13399);
or U14157 (N_14157,N_13474,N_12855);
or U14158 (N_14158,N_12965,N_13137);
nor U14159 (N_14159,N_13320,N_12780);
nor U14160 (N_14160,N_12945,N_13193);
nand U14161 (N_14161,N_12960,N_12814);
and U14162 (N_14162,N_13300,N_13398);
and U14163 (N_14163,N_13264,N_13366);
nor U14164 (N_14164,N_13152,N_13250);
and U14165 (N_14165,N_13448,N_13034);
or U14166 (N_14166,N_13039,N_13298);
and U14167 (N_14167,N_12826,N_13498);
nand U14168 (N_14168,N_13279,N_13252);
nand U14169 (N_14169,N_13167,N_13250);
nor U14170 (N_14170,N_13284,N_13266);
nand U14171 (N_14171,N_13494,N_12993);
or U14172 (N_14172,N_13422,N_13243);
and U14173 (N_14173,N_12915,N_13262);
or U14174 (N_14174,N_12768,N_13171);
or U14175 (N_14175,N_13497,N_12783);
and U14176 (N_14176,N_13307,N_12789);
nand U14177 (N_14177,N_13256,N_13028);
or U14178 (N_14178,N_13140,N_13196);
nand U14179 (N_14179,N_12755,N_13055);
nand U14180 (N_14180,N_12925,N_12804);
and U14181 (N_14181,N_13036,N_13206);
nand U14182 (N_14182,N_13204,N_13122);
nor U14183 (N_14183,N_13055,N_13142);
or U14184 (N_14184,N_13206,N_13081);
or U14185 (N_14185,N_13047,N_12921);
nor U14186 (N_14186,N_12942,N_13063);
nor U14187 (N_14187,N_13212,N_12896);
or U14188 (N_14188,N_13308,N_12799);
nand U14189 (N_14189,N_12812,N_13059);
and U14190 (N_14190,N_13427,N_13274);
nand U14191 (N_14191,N_13024,N_12863);
nor U14192 (N_14192,N_13450,N_13257);
or U14193 (N_14193,N_13439,N_13401);
and U14194 (N_14194,N_13073,N_12894);
or U14195 (N_14195,N_12902,N_13280);
and U14196 (N_14196,N_13451,N_13048);
or U14197 (N_14197,N_13233,N_13438);
nor U14198 (N_14198,N_13319,N_13257);
nand U14199 (N_14199,N_13498,N_13283);
and U14200 (N_14200,N_13405,N_13134);
nor U14201 (N_14201,N_13061,N_12989);
and U14202 (N_14202,N_12857,N_13460);
and U14203 (N_14203,N_13425,N_12971);
nor U14204 (N_14204,N_13386,N_13253);
nand U14205 (N_14205,N_13367,N_13324);
nand U14206 (N_14206,N_13099,N_13471);
nor U14207 (N_14207,N_13276,N_13227);
nand U14208 (N_14208,N_12848,N_13434);
nand U14209 (N_14209,N_12851,N_13293);
nand U14210 (N_14210,N_12828,N_13318);
nor U14211 (N_14211,N_12847,N_13159);
and U14212 (N_14212,N_13332,N_12754);
nand U14213 (N_14213,N_12833,N_13482);
nor U14214 (N_14214,N_12935,N_12846);
and U14215 (N_14215,N_12832,N_13228);
and U14216 (N_14216,N_12826,N_12869);
nor U14217 (N_14217,N_13026,N_12798);
nor U14218 (N_14218,N_12976,N_13027);
or U14219 (N_14219,N_13169,N_12853);
nor U14220 (N_14220,N_13321,N_12874);
nand U14221 (N_14221,N_12914,N_13096);
nand U14222 (N_14222,N_12922,N_13030);
and U14223 (N_14223,N_13083,N_12835);
or U14224 (N_14224,N_13215,N_12812);
xor U14225 (N_14225,N_12928,N_13076);
nor U14226 (N_14226,N_12956,N_13342);
and U14227 (N_14227,N_13298,N_12765);
nor U14228 (N_14228,N_13264,N_13190);
nand U14229 (N_14229,N_13249,N_13111);
nand U14230 (N_14230,N_12891,N_13327);
nand U14231 (N_14231,N_13029,N_13322);
or U14232 (N_14232,N_13171,N_12762);
nand U14233 (N_14233,N_12854,N_12979);
nor U14234 (N_14234,N_12936,N_12751);
nor U14235 (N_14235,N_13081,N_13482);
and U14236 (N_14236,N_13464,N_12760);
nand U14237 (N_14237,N_12929,N_12762);
nand U14238 (N_14238,N_13420,N_13095);
xor U14239 (N_14239,N_13033,N_12864);
or U14240 (N_14240,N_12840,N_12845);
nor U14241 (N_14241,N_13013,N_12829);
nor U14242 (N_14242,N_13129,N_13350);
or U14243 (N_14243,N_13094,N_13126);
or U14244 (N_14244,N_12843,N_13221);
nand U14245 (N_14245,N_13310,N_13251);
and U14246 (N_14246,N_13066,N_13044);
xnor U14247 (N_14247,N_13199,N_12856);
or U14248 (N_14248,N_13210,N_13243);
nand U14249 (N_14249,N_13478,N_12928);
nand U14250 (N_14250,N_13643,N_13984);
nand U14251 (N_14251,N_13696,N_13741);
nand U14252 (N_14252,N_13665,N_13860);
or U14253 (N_14253,N_14230,N_13944);
nor U14254 (N_14254,N_13865,N_14132);
and U14255 (N_14255,N_13770,N_13928);
and U14256 (N_14256,N_14039,N_13875);
nor U14257 (N_14257,N_13676,N_13743);
nand U14258 (N_14258,N_14136,N_13744);
or U14259 (N_14259,N_13710,N_14143);
nor U14260 (N_14260,N_13756,N_14072);
nand U14261 (N_14261,N_13653,N_13949);
xnor U14262 (N_14262,N_14111,N_13524);
nand U14263 (N_14263,N_13712,N_13622);
nor U14264 (N_14264,N_13648,N_13686);
and U14265 (N_14265,N_13742,N_14134);
nor U14266 (N_14266,N_13651,N_13593);
or U14267 (N_14267,N_13790,N_13571);
or U14268 (N_14268,N_14018,N_13572);
or U14269 (N_14269,N_13609,N_14188);
and U14270 (N_14270,N_13697,N_14218);
nor U14271 (N_14271,N_13706,N_14228);
nand U14272 (N_14272,N_14145,N_13924);
or U14273 (N_14273,N_13728,N_14179);
and U14274 (N_14274,N_13867,N_13847);
nor U14275 (N_14275,N_13632,N_13916);
and U14276 (N_14276,N_14138,N_14240);
nand U14277 (N_14277,N_13739,N_14144);
and U14278 (N_14278,N_14060,N_13723);
or U14279 (N_14279,N_13608,N_14006);
nor U14280 (N_14280,N_13635,N_14189);
nor U14281 (N_14281,N_13624,N_13797);
and U14282 (N_14282,N_14090,N_13887);
nand U14283 (N_14283,N_14055,N_14159);
and U14284 (N_14284,N_13817,N_14244);
nand U14285 (N_14285,N_13920,N_14000);
xor U14286 (N_14286,N_13563,N_13904);
and U14287 (N_14287,N_13729,N_13844);
nand U14288 (N_14288,N_13833,N_14012);
nand U14289 (N_14289,N_13557,N_14243);
and U14290 (N_14290,N_13985,N_13546);
or U14291 (N_14291,N_14223,N_13559);
nor U14292 (N_14292,N_13783,N_14029);
or U14293 (N_14293,N_13955,N_13718);
nand U14294 (N_14294,N_13664,N_14104);
nand U14295 (N_14295,N_13510,N_13699);
nand U14296 (N_14296,N_14091,N_13879);
or U14297 (N_14297,N_13597,N_13972);
or U14298 (N_14298,N_13599,N_14222);
nor U14299 (N_14299,N_13550,N_13780);
nand U14300 (N_14300,N_13650,N_14085);
nor U14301 (N_14301,N_13895,N_13812);
nand U14302 (N_14302,N_13787,N_14219);
or U14303 (N_14303,N_13607,N_14140);
and U14304 (N_14304,N_13900,N_14096);
nand U14305 (N_14305,N_13574,N_14206);
nand U14306 (N_14306,N_13842,N_14028);
or U14307 (N_14307,N_14120,N_13583);
xor U14308 (N_14308,N_13766,N_13529);
nor U14309 (N_14309,N_13601,N_14087);
nand U14310 (N_14310,N_13631,N_13936);
xor U14311 (N_14311,N_14214,N_13694);
nor U14312 (N_14312,N_14142,N_13575);
nor U14313 (N_14313,N_13621,N_13685);
or U14314 (N_14314,N_13737,N_13657);
nand U14315 (N_14315,N_14036,N_14125);
nand U14316 (N_14316,N_13745,N_14075);
nor U14317 (N_14317,N_13692,N_13771);
xor U14318 (N_14318,N_14050,N_13813);
nor U14319 (N_14319,N_13795,N_13940);
and U14320 (N_14320,N_13625,N_13809);
nor U14321 (N_14321,N_13827,N_13682);
and U14322 (N_14322,N_14108,N_14068);
or U14323 (N_14323,N_13990,N_14157);
nor U14324 (N_14324,N_14112,N_13560);
xnor U14325 (N_14325,N_13604,N_13616);
and U14326 (N_14326,N_13722,N_14187);
nand U14327 (N_14327,N_13644,N_13979);
or U14328 (N_14328,N_13964,N_14163);
xor U14329 (N_14329,N_14242,N_14161);
or U14330 (N_14330,N_13957,N_13781);
or U14331 (N_14331,N_13590,N_13514);
nand U14332 (N_14332,N_13769,N_13782);
or U14333 (N_14333,N_14046,N_14180);
nand U14334 (N_14334,N_14025,N_13548);
or U14335 (N_14335,N_14040,N_13760);
and U14336 (N_14336,N_13731,N_13610);
or U14337 (N_14337,N_13912,N_13713);
nor U14338 (N_14338,N_14093,N_13855);
nor U14339 (N_14339,N_14007,N_14098);
or U14340 (N_14340,N_13589,N_13568);
nor U14341 (N_14341,N_13939,N_14213);
or U14342 (N_14342,N_13603,N_14131);
or U14343 (N_14343,N_14146,N_14209);
and U14344 (N_14344,N_13901,N_14081);
or U14345 (N_14345,N_14182,N_13824);
or U14346 (N_14346,N_13750,N_13998);
nand U14347 (N_14347,N_13947,N_14186);
or U14348 (N_14348,N_14066,N_13974);
nand U14349 (N_14349,N_14153,N_13841);
nand U14350 (N_14350,N_14114,N_14015);
nor U14351 (N_14351,N_14003,N_13700);
or U14352 (N_14352,N_13522,N_14162);
and U14353 (N_14353,N_13945,N_14231);
or U14354 (N_14354,N_13826,N_14211);
nor U14355 (N_14355,N_14249,N_13871);
nand U14356 (N_14356,N_14118,N_14070);
and U14357 (N_14357,N_13831,N_13558);
or U14358 (N_14358,N_14048,N_14172);
and U14359 (N_14359,N_14129,N_13882);
nor U14360 (N_14360,N_14052,N_13630);
nor U14361 (N_14361,N_14024,N_14110);
and U14362 (N_14362,N_13537,N_13883);
nor U14363 (N_14363,N_13645,N_14170);
and U14364 (N_14364,N_14234,N_13776);
and U14365 (N_14365,N_14079,N_14109);
and U14366 (N_14366,N_13956,N_13897);
or U14367 (N_14367,N_13561,N_13997);
or U14368 (N_14368,N_13500,N_14019);
or U14369 (N_14369,N_14002,N_14225);
and U14370 (N_14370,N_14247,N_14226);
and U14371 (N_14371,N_13840,N_13677);
nand U14372 (N_14372,N_13881,N_14205);
xnor U14373 (N_14373,N_13646,N_13751);
or U14374 (N_14374,N_13820,N_13856);
and U14375 (N_14375,N_14196,N_13633);
or U14376 (N_14376,N_13950,N_14013);
nor U14377 (N_14377,N_13768,N_13556);
nand U14378 (N_14378,N_13672,N_13838);
and U14379 (N_14379,N_14154,N_14042);
nand U14380 (N_14380,N_13687,N_14216);
nor U14381 (N_14381,N_13815,N_14097);
nand U14382 (N_14382,N_13937,N_13963);
nor U14383 (N_14383,N_13970,N_13701);
nand U14384 (N_14384,N_13836,N_14168);
or U14385 (N_14385,N_13932,N_13849);
or U14386 (N_14386,N_13618,N_14232);
and U14387 (N_14387,N_13654,N_13663);
and U14388 (N_14388,N_13927,N_14160);
nand U14389 (N_14389,N_13905,N_13872);
nor U14390 (N_14390,N_13878,N_13503);
or U14391 (N_14391,N_13688,N_13555);
nor U14392 (N_14392,N_13906,N_13767);
xnor U14393 (N_14393,N_14178,N_14167);
and U14394 (N_14394,N_13716,N_13702);
nor U14395 (N_14395,N_13647,N_13890);
nor U14396 (N_14396,N_13715,N_13981);
nor U14397 (N_14397,N_14126,N_13885);
nor U14398 (N_14398,N_13851,N_14026);
nor U14399 (N_14399,N_13938,N_13825);
nor U14400 (N_14400,N_13542,N_14043);
or U14401 (N_14401,N_14010,N_13794);
nor U14402 (N_14402,N_13775,N_13764);
and U14403 (N_14403,N_13868,N_14238);
nand U14404 (N_14404,N_14008,N_14204);
and U14405 (N_14405,N_14175,N_13870);
nor U14406 (N_14406,N_13530,N_13948);
nand U14407 (N_14407,N_13965,N_14217);
nor U14408 (N_14408,N_13693,N_13791);
nor U14409 (N_14409,N_13547,N_13993);
nor U14410 (N_14410,N_13951,N_14047);
nand U14411 (N_14411,N_14235,N_14014);
xnor U14412 (N_14412,N_13536,N_14094);
xnor U14413 (N_14413,N_14053,N_13892);
nand U14414 (N_14414,N_13942,N_13977);
nand U14415 (N_14415,N_13914,N_13858);
xnor U14416 (N_14416,N_14001,N_13578);
nand U14417 (N_14417,N_14128,N_13954);
nor U14418 (N_14418,N_13501,N_13786);
or U14419 (N_14419,N_14033,N_13995);
or U14420 (N_14420,N_13511,N_13545);
and U14421 (N_14421,N_13789,N_13926);
or U14422 (N_14422,N_13620,N_14076);
or U14423 (N_14423,N_13573,N_13921);
and U14424 (N_14424,N_13839,N_14022);
and U14425 (N_14425,N_14005,N_14184);
nor U14426 (N_14426,N_13543,N_13991);
nand U14427 (N_14427,N_14173,N_13999);
and U14428 (N_14428,N_13758,N_13505);
or U14429 (N_14429,N_13988,N_13658);
nand U14430 (N_14430,N_14199,N_14084);
nor U14431 (N_14431,N_13866,N_13735);
or U14432 (N_14432,N_14246,N_13891);
nand U14433 (N_14433,N_13757,N_14065);
nor U14434 (N_14434,N_13869,N_14032);
nand U14435 (N_14435,N_13535,N_13580);
and U14436 (N_14436,N_13896,N_13551);
nand U14437 (N_14437,N_13639,N_14041);
nand U14438 (N_14438,N_13818,N_13553);
or U14439 (N_14439,N_13661,N_14017);
nand U14440 (N_14440,N_14020,N_13520);
nand U14441 (N_14441,N_13835,N_13711);
nor U14442 (N_14442,N_13864,N_13634);
nand U14443 (N_14443,N_13538,N_13637);
or U14444 (N_14444,N_13541,N_14045);
or U14445 (N_14445,N_13534,N_14082);
nor U14446 (N_14446,N_14044,N_13843);
nor U14447 (N_14447,N_13698,N_13502);
xor U14448 (N_14448,N_13755,N_13800);
or U14449 (N_14449,N_13606,N_13525);
nand U14450 (N_14450,N_13832,N_14183);
nand U14451 (N_14451,N_13982,N_14038);
or U14452 (N_14452,N_14004,N_13674);
or U14453 (N_14453,N_13941,N_14095);
or U14454 (N_14454,N_13747,N_14124);
and U14455 (N_14455,N_13959,N_13953);
nor U14456 (N_14456,N_13935,N_13933);
and U14457 (N_14457,N_14139,N_14227);
nor U14458 (N_14458,N_14220,N_14195);
nor U14459 (N_14459,N_14049,N_14059);
nor U14460 (N_14460,N_14191,N_14245);
nor U14461 (N_14461,N_13913,N_14203);
nor U14462 (N_14462,N_13627,N_13512);
or U14463 (N_14463,N_13778,N_13798);
nor U14464 (N_14464,N_13684,N_13504);
nand U14465 (N_14465,N_13893,N_13822);
or U14466 (N_14466,N_13642,N_13554);
nand U14467 (N_14467,N_14063,N_13805);
or U14468 (N_14468,N_14171,N_13752);
nand U14469 (N_14469,N_14021,N_13670);
and U14470 (N_14470,N_14086,N_14210);
or U14471 (N_14471,N_13703,N_14080);
and U14472 (N_14472,N_14116,N_14207);
nor U14473 (N_14473,N_13989,N_14169);
and U14474 (N_14474,N_13585,N_13588);
or U14475 (N_14475,N_13929,N_14229);
nor U14476 (N_14476,N_13669,N_13626);
and U14477 (N_14477,N_13969,N_13814);
and U14478 (N_14478,N_13721,N_13763);
and U14479 (N_14479,N_14034,N_13733);
nor U14480 (N_14480,N_14155,N_13788);
nand U14481 (N_14481,N_14176,N_14174);
nand U14482 (N_14482,N_13638,N_14099);
xor U14483 (N_14483,N_13777,N_13876);
nor U14484 (N_14484,N_13811,N_13980);
nor U14485 (N_14485,N_13726,N_14239);
or U14486 (N_14486,N_13943,N_14233);
or U14487 (N_14487,N_13884,N_14202);
nor U14488 (N_14488,N_13615,N_13738);
or U14489 (N_14489,N_13544,N_13848);
or U14490 (N_14490,N_13894,N_14101);
or U14491 (N_14491,N_13886,N_14221);
nor U14492 (N_14492,N_13819,N_13837);
nor U14493 (N_14493,N_13584,N_13857);
nand U14494 (N_14494,N_14089,N_13908);
nor U14495 (N_14495,N_13666,N_13911);
or U14496 (N_14496,N_14057,N_14127);
nor U14497 (N_14497,N_13803,N_13614);
or U14498 (N_14498,N_13598,N_13804);
and U14499 (N_14499,N_13660,N_14148);
and U14500 (N_14500,N_14088,N_14105);
xor U14501 (N_14501,N_13834,N_13528);
nand U14502 (N_14502,N_13679,N_13532);
and U14503 (N_14503,N_13533,N_14192);
or U14504 (N_14504,N_13976,N_13829);
or U14505 (N_14505,N_13996,N_14241);
nand U14506 (N_14506,N_13673,N_13730);
or U14507 (N_14507,N_13569,N_13952);
nor U14508 (N_14508,N_13570,N_13774);
or U14509 (N_14509,N_13968,N_14137);
or U14510 (N_14510,N_13992,N_13652);
or U14511 (N_14511,N_13695,N_14119);
nor U14512 (N_14512,N_13678,N_13612);
or U14513 (N_14513,N_13531,N_14151);
or U14514 (N_14514,N_13773,N_13507);
nand U14515 (N_14515,N_13772,N_13523);
and U14516 (N_14516,N_13845,N_13960);
and U14517 (N_14517,N_13641,N_14166);
or U14518 (N_14518,N_13792,N_13539);
or U14519 (N_14519,N_13807,N_13907);
or U14520 (N_14520,N_13705,N_14100);
and U14521 (N_14521,N_13724,N_14147);
and U14522 (N_14522,N_13978,N_13823);
nor U14523 (N_14523,N_14117,N_13962);
and U14524 (N_14524,N_14011,N_14193);
or U14525 (N_14525,N_13662,N_13517);
xor U14526 (N_14526,N_13566,N_13748);
and U14527 (N_14527,N_13521,N_13828);
nand U14528 (N_14528,N_14200,N_14164);
nor U14529 (N_14529,N_14133,N_13581);
and U14530 (N_14530,N_14054,N_13975);
nor U14531 (N_14531,N_13902,N_14236);
nand U14532 (N_14532,N_13785,N_13873);
nand U14533 (N_14533,N_13753,N_13613);
and U14534 (N_14534,N_13810,N_13675);
or U14535 (N_14535,N_14073,N_13898);
nand U14536 (N_14536,N_13602,N_13565);
xnor U14537 (N_14537,N_13889,N_13727);
nand U14538 (N_14538,N_13714,N_14078);
xnor U14539 (N_14539,N_13587,N_13987);
nand U14540 (N_14540,N_13564,N_13910);
xor U14541 (N_14541,N_13600,N_13617);
and U14542 (N_14542,N_13717,N_14141);
or U14543 (N_14543,N_13934,N_13506);
and U14544 (N_14544,N_14115,N_13863);
nand U14545 (N_14545,N_14009,N_14083);
or U14546 (N_14546,N_14061,N_14135);
or U14547 (N_14547,N_13946,N_13862);
xor U14548 (N_14548,N_14092,N_13594);
nand U14549 (N_14549,N_13909,N_13779);
nor U14550 (N_14550,N_13793,N_13983);
nand U14551 (N_14551,N_13704,N_13667);
or U14552 (N_14552,N_13552,N_13899);
nor U14553 (N_14553,N_13853,N_14023);
or U14554 (N_14554,N_14102,N_14149);
and U14555 (N_14555,N_13680,N_14031);
or U14556 (N_14556,N_14067,N_13888);
nor U14557 (N_14557,N_14121,N_13852);
and U14558 (N_14558,N_14030,N_13799);
and U14559 (N_14559,N_13736,N_13515);
or U14560 (N_14560,N_13579,N_13519);
and U14561 (N_14561,N_13966,N_13725);
xnor U14562 (N_14562,N_14150,N_14113);
or U14563 (N_14563,N_14190,N_13567);
or U14564 (N_14564,N_14208,N_14123);
nand U14565 (N_14565,N_13821,N_13762);
nor U14566 (N_14566,N_13986,N_13659);
nand U14567 (N_14567,N_13709,N_13683);
nand U14568 (N_14568,N_13761,N_13967);
xor U14569 (N_14569,N_14185,N_14107);
and U14570 (N_14570,N_13880,N_14077);
or U14571 (N_14571,N_13918,N_13754);
or U14572 (N_14572,N_13759,N_13619);
xor U14573 (N_14573,N_13690,N_13516);
nand U14574 (N_14574,N_14056,N_13877);
nor U14575 (N_14575,N_13527,N_13861);
or U14576 (N_14576,N_13508,N_13586);
and U14577 (N_14577,N_13719,N_13595);
nor U14578 (N_14578,N_13816,N_13846);
and U14579 (N_14579,N_13720,N_13919);
nor U14580 (N_14580,N_13784,N_14103);
and U14581 (N_14581,N_14074,N_13973);
and U14582 (N_14582,N_14156,N_13796);
nand U14583 (N_14583,N_14122,N_13509);
nor U14584 (N_14584,N_13596,N_13922);
nand U14585 (N_14585,N_13749,N_13915);
nand U14586 (N_14586,N_13874,N_13806);
xnor U14587 (N_14587,N_14198,N_13576);
nor U14588 (N_14588,N_14177,N_13689);
xor U14589 (N_14589,N_13931,N_14152);
nand U14590 (N_14590,N_14035,N_13923);
nor U14591 (N_14591,N_14106,N_13707);
or U14592 (N_14592,N_13801,N_13540);
nor U14593 (N_14593,N_13961,N_13802);
nor U14594 (N_14594,N_13591,N_14181);
nor U14595 (N_14595,N_14224,N_14062);
and U14596 (N_14596,N_14212,N_13746);
nand U14597 (N_14597,N_13925,N_13605);
and U14598 (N_14598,N_14201,N_13958);
xnor U14599 (N_14599,N_13611,N_13734);
and U14600 (N_14600,N_13930,N_14194);
and U14601 (N_14601,N_13592,N_13518);
and U14602 (N_14602,N_14069,N_13668);
nor U14603 (N_14603,N_13917,N_13740);
and U14604 (N_14604,N_14158,N_13577);
nand U14605 (N_14605,N_14237,N_14058);
nor U14606 (N_14606,N_13549,N_14037);
and U14607 (N_14607,N_13708,N_13765);
or U14608 (N_14608,N_13562,N_13994);
nand U14609 (N_14609,N_14071,N_13671);
nand U14610 (N_14610,N_13850,N_13903);
or U14611 (N_14611,N_13649,N_13854);
or U14612 (N_14612,N_13526,N_14248);
xnor U14613 (N_14613,N_14215,N_13513);
or U14614 (N_14614,N_13629,N_14165);
nand U14615 (N_14615,N_14016,N_14197);
nand U14616 (N_14616,N_13691,N_13640);
nand U14617 (N_14617,N_13732,N_13808);
and U14618 (N_14618,N_13636,N_13859);
or U14619 (N_14619,N_13623,N_14027);
and U14620 (N_14620,N_14064,N_14051);
nor U14621 (N_14621,N_13656,N_13971);
nand U14622 (N_14622,N_14130,N_13655);
nor U14623 (N_14623,N_13582,N_13628);
and U14624 (N_14624,N_13681,N_13830);
nand U14625 (N_14625,N_14149,N_13567);
nor U14626 (N_14626,N_13890,N_14143);
and U14627 (N_14627,N_14023,N_14025);
or U14628 (N_14628,N_13633,N_13646);
nand U14629 (N_14629,N_13958,N_14038);
xor U14630 (N_14630,N_13651,N_13559);
and U14631 (N_14631,N_13578,N_13853);
or U14632 (N_14632,N_13913,N_13635);
nor U14633 (N_14633,N_13751,N_13870);
nor U14634 (N_14634,N_14111,N_13742);
and U14635 (N_14635,N_13634,N_13890);
nand U14636 (N_14636,N_13834,N_14153);
nor U14637 (N_14637,N_13642,N_14019);
nand U14638 (N_14638,N_14141,N_14083);
nand U14639 (N_14639,N_14081,N_13685);
nor U14640 (N_14640,N_14218,N_13514);
or U14641 (N_14641,N_13622,N_13931);
and U14642 (N_14642,N_13699,N_14058);
and U14643 (N_14643,N_13719,N_13968);
nand U14644 (N_14644,N_13934,N_13566);
nor U14645 (N_14645,N_14115,N_13997);
xnor U14646 (N_14646,N_14243,N_13787);
or U14647 (N_14647,N_13780,N_13740);
and U14648 (N_14648,N_13894,N_13748);
and U14649 (N_14649,N_14249,N_13708);
or U14650 (N_14650,N_13857,N_13813);
nand U14651 (N_14651,N_13520,N_13927);
or U14652 (N_14652,N_13537,N_14188);
or U14653 (N_14653,N_14036,N_13960);
nand U14654 (N_14654,N_14128,N_13891);
nand U14655 (N_14655,N_14229,N_14101);
and U14656 (N_14656,N_13675,N_13607);
and U14657 (N_14657,N_13944,N_13709);
nand U14658 (N_14658,N_14211,N_14033);
or U14659 (N_14659,N_13543,N_13930);
and U14660 (N_14660,N_14017,N_14230);
and U14661 (N_14661,N_13939,N_14177);
and U14662 (N_14662,N_14097,N_14075);
nor U14663 (N_14663,N_13772,N_14120);
nand U14664 (N_14664,N_13755,N_13543);
nor U14665 (N_14665,N_13632,N_13593);
nand U14666 (N_14666,N_14225,N_14006);
or U14667 (N_14667,N_14004,N_13961);
or U14668 (N_14668,N_13723,N_14105);
nor U14669 (N_14669,N_13881,N_13804);
or U14670 (N_14670,N_13637,N_14195);
nand U14671 (N_14671,N_14240,N_14084);
nand U14672 (N_14672,N_13792,N_14175);
or U14673 (N_14673,N_13563,N_13623);
nor U14674 (N_14674,N_13781,N_14112);
xor U14675 (N_14675,N_13838,N_13894);
nand U14676 (N_14676,N_14235,N_13592);
and U14677 (N_14677,N_13564,N_13990);
and U14678 (N_14678,N_13874,N_13970);
nand U14679 (N_14679,N_13799,N_13559);
nand U14680 (N_14680,N_13526,N_13574);
and U14681 (N_14681,N_13786,N_13526);
nand U14682 (N_14682,N_13863,N_13826);
nor U14683 (N_14683,N_14110,N_13623);
nor U14684 (N_14684,N_13815,N_13988);
nand U14685 (N_14685,N_13553,N_13860);
nor U14686 (N_14686,N_13965,N_13895);
or U14687 (N_14687,N_13965,N_14161);
and U14688 (N_14688,N_13566,N_14112);
and U14689 (N_14689,N_14004,N_14122);
or U14690 (N_14690,N_14150,N_13802);
nor U14691 (N_14691,N_14167,N_13718);
or U14692 (N_14692,N_14122,N_13834);
and U14693 (N_14693,N_13579,N_14089);
or U14694 (N_14694,N_13734,N_13665);
nor U14695 (N_14695,N_13885,N_13855);
nor U14696 (N_14696,N_13748,N_13927);
and U14697 (N_14697,N_14018,N_14090);
nor U14698 (N_14698,N_14186,N_13913);
and U14699 (N_14699,N_14023,N_14134);
and U14700 (N_14700,N_14140,N_14082);
xnor U14701 (N_14701,N_13917,N_14086);
and U14702 (N_14702,N_13524,N_13596);
or U14703 (N_14703,N_13769,N_13718);
nor U14704 (N_14704,N_14188,N_13628);
nand U14705 (N_14705,N_13987,N_14151);
nor U14706 (N_14706,N_13924,N_13742);
and U14707 (N_14707,N_14154,N_13771);
nand U14708 (N_14708,N_13633,N_14004);
or U14709 (N_14709,N_13697,N_14154);
nor U14710 (N_14710,N_13603,N_13718);
nor U14711 (N_14711,N_13976,N_13730);
and U14712 (N_14712,N_14102,N_13608);
or U14713 (N_14713,N_13619,N_13569);
nand U14714 (N_14714,N_13627,N_13651);
and U14715 (N_14715,N_13850,N_14031);
nor U14716 (N_14716,N_13786,N_14027);
nand U14717 (N_14717,N_13824,N_13857);
nor U14718 (N_14718,N_13507,N_14248);
or U14719 (N_14719,N_14224,N_13907);
nor U14720 (N_14720,N_13732,N_14204);
and U14721 (N_14721,N_14242,N_14118);
and U14722 (N_14722,N_13802,N_13513);
or U14723 (N_14723,N_13789,N_13961);
nor U14724 (N_14724,N_13703,N_13770);
nor U14725 (N_14725,N_14234,N_13786);
and U14726 (N_14726,N_14030,N_13925);
nor U14727 (N_14727,N_14234,N_13729);
or U14728 (N_14728,N_14051,N_13717);
and U14729 (N_14729,N_13549,N_14102);
and U14730 (N_14730,N_13866,N_13789);
and U14731 (N_14731,N_13531,N_13644);
nand U14732 (N_14732,N_13929,N_14016);
and U14733 (N_14733,N_13853,N_13665);
or U14734 (N_14734,N_13997,N_13935);
nand U14735 (N_14735,N_13633,N_14022);
or U14736 (N_14736,N_14183,N_13622);
or U14737 (N_14737,N_13729,N_13706);
xnor U14738 (N_14738,N_13929,N_13557);
nand U14739 (N_14739,N_13677,N_13539);
nor U14740 (N_14740,N_14210,N_13590);
nand U14741 (N_14741,N_13619,N_13618);
and U14742 (N_14742,N_13628,N_13612);
nor U14743 (N_14743,N_13972,N_13701);
nand U14744 (N_14744,N_13756,N_14228);
nand U14745 (N_14745,N_14023,N_13560);
nor U14746 (N_14746,N_13647,N_13930);
or U14747 (N_14747,N_13976,N_13875);
or U14748 (N_14748,N_14121,N_13662);
or U14749 (N_14749,N_13786,N_13916);
and U14750 (N_14750,N_14091,N_13615);
or U14751 (N_14751,N_13936,N_14226);
and U14752 (N_14752,N_14207,N_14027);
nand U14753 (N_14753,N_13811,N_13758);
and U14754 (N_14754,N_14022,N_13572);
and U14755 (N_14755,N_13584,N_14212);
nand U14756 (N_14756,N_14177,N_13904);
nand U14757 (N_14757,N_13696,N_14029);
nor U14758 (N_14758,N_13688,N_14095);
nor U14759 (N_14759,N_14003,N_13893);
nand U14760 (N_14760,N_13613,N_13736);
nand U14761 (N_14761,N_13705,N_13701);
nor U14762 (N_14762,N_13694,N_13622);
nand U14763 (N_14763,N_13789,N_14052);
nand U14764 (N_14764,N_14231,N_13674);
and U14765 (N_14765,N_13870,N_13637);
and U14766 (N_14766,N_13754,N_13837);
nand U14767 (N_14767,N_14205,N_13869);
and U14768 (N_14768,N_14071,N_13733);
or U14769 (N_14769,N_13556,N_13918);
or U14770 (N_14770,N_13946,N_14135);
and U14771 (N_14771,N_13660,N_13727);
or U14772 (N_14772,N_14025,N_14189);
nor U14773 (N_14773,N_14122,N_13725);
and U14774 (N_14774,N_14182,N_13730);
xnor U14775 (N_14775,N_13922,N_13883);
xor U14776 (N_14776,N_14188,N_14012);
or U14777 (N_14777,N_14207,N_13827);
nor U14778 (N_14778,N_13769,N_13693);
nor U14779 (N_14779,N_13772,N_13663);
nor U14780 (N_14780,N_13553,N_13755);
nor U14781 (N_14781,N_14172,N_13705);
nor U14782 (N_14782,N_13780,N_14244);
or U14783 (N_14783,N_13563,N_13529);
xnor U14784 (N_14784,N_13538,N_14016);
or U14785 (N_14785,N_14127,N_14107);
and U14786 (N_14786,N_14081,N_13564);
nor U14787 (N_14787,N_14239,N_13626);
or U14788 (N_14788,N_14220,N_14140);
nand U14789 (N_14789,N_13694,N_13912);
nor U14790 (N_14790,N_13844,N_14157);
xor U14791 (N_14791,N_14028,N_13692);
nand U14792 (N_14792,N_14037,N_13971);
or U14793 (N_14793,N_13878,N_13581);
nand U14794 (N_14794,N_13912,N_13889);
nand U14795 (N_14795,N_13902,N_13980);
and U14796 (N_14796,N_14086,N_13961);
and U14797 (N_14797,N_14215,N_13958);
nor U14798 (N_14798,N_14131,N_13635);
nor U14799 (N_14799,N_14003,N_13760);
or U14800 (N_14800,N_13592,N_13522);
nand U14801 (N_14801,N_13708,N_14109);
and U14802 (N_14802,N_13899,N_13502);
nand U14803 (N_14803,N_13610,N_13515);
or U14804 (N_14804,N_13642,N_14214);
nand U14805 (N_14805,N_13779,N_13845);
nor U14806 (N_14806,N_13765,N_13682);
nand U14807 (N_14807,N_13952,N_13531);
nor U14808 (N_14808,N_13889,N_13645);
nand U14809 (N_14809,N_14100,N_13939);
and U14810 (N_14810,N_13679,N_14115);
and U14811 (N_14811,N_14219,N_13970);
nand U14812 (N_14812,N_14145,N_13669);
nand U14813 (N_14813,N_13997,N_13796);
and U14814 (N_14814,N_14167,N_13781);
nand U14815 (N_14815,N_13844,N_13651);
and U14816 (N_14816,N_14123,N_14207);
and U14817 (N_14817,N_14010,N_14016);
or U14818 (N_14818,N_13868,N_14169);
xor U14819 (N_14819,N_14035,N_14040);
nand U14820 (N_14820,N_14060,N_13664);
and U14821 (N_14821,N_13579,N_14173);
nand U14822 (N_14822,N_13564,N_14136);
and U14823 (N_14823,N_13522,N_13911);
and U14824 (N_14824,N_14039,N_13815);
and U14825 (N_14825,N_13964,N_13649);
and U14826 (N_14826,N_13814,N_13520);
nand U14827 (N_14827,N_14119,N_13517);
nand U14828 (N_14828,N_13667,N_13833);
nor U14829 (N_14829,N_13614,N_14100);
nand U14830 (N_14830,N_14198,N_13885);
and U14831 (N_14831,N_13884,N_14207);
nand U14832 (N_14832,N_13720,N_13562);
nor U14833 (N_14833,N_13544,N_13655);
nand U14834 (N_14834,N_13936,N_13677);
or U14835 (N_14835,N_13836,N_14191);
and U14836 (N_14836,N_13596,N_13706);
and U14837 (N_14837,N_13978,N_14207);
xor U14838 (N_14838,N_14149,N_14047);
nand U14839 (N_14839,N_14160,N_14014);
and U14840 (N_14840,N_14087,N_13646);
nand U14841 (N_14841,N_13831,N_14193);
nand U14842 (N_14842,N_14193,N_13741);
nor U14843 (N_14843,N_14045,N_13751);
and U14844 (N_14844,N_13947,N_13538);
nor U14845 (N_14845,N_13510,N_13928);
and U14846 (N_14846,N_14196,N_13911);
xor U14847 (N_14847,N_13761,N_14039);
nand U14848 (N_14848,N_13650,N_13845);
or U14849 (N_14849,N_13994,N_13527);
or U14850 (N_14850,N_13653,N_13784);
or U14851 (N_14851,N_14162,N_13683);
and U14852 (N_14852,N_14163,N_14124);
and U14853 (N_14853,N_13572,N_14056);
or U14854 (N_14854,N_13656,N_13977);
or U14855 (N_14855,N_13585,N_13982);
nand U14856 (N_14856,N_13627,N_14150);
nand U14857 (N_14857,N_13670,N_13907);
nand U14858 (N_14858,N_13744,N_14039);
and U14859 (N_14859,N_14234,N_14078);
nor U14860 (N_14860,N_14128,N_14085);
nand U14861 (N_14861,N_13569,N_14150);
and U14862 (N_14862,N_13919,N_14192);
or U14863 (N_14863,N_14233,N_13575);
nor U14864 (N_14864,N_13687,N_13861);
and U14865 (N_14865,N_14140,N_13809);
and U14866 (N_14866,N_13513,N_14111);
nor U14867 (N_14867,N_14238,N_13795);
and U14868 (N_14868,N_13585,N_13933);
and U14869 (N_14869,N_13887,N_14125);
nand U14870 (N_14870,N_14162,N_14103);
or U14871 (N_14871,N_13963,N_14216);
nand U14872 (N_14872,N_13612,N_13795);
and U14873 (N_14873,N_13572,N_13881);
nand U14874 (N_14874,N_13767,N_13619);
nand U14875 (N_14875,N_13611,N_13779);
nand U14876 (N_14876,N_14131,N_13686);
or U14877 (N_14877,N_14174,N_13646);
nor U14878 (N_14878,N_13665,N_13532);
nor U14879 (N_14879,N_13744,N_13784);
nor U14880 (N_14880,N_13920,N_13775);
and U14881 (N_14881,N_13996,N_13666);
or U14882 (N_14882,N_14085,N_14139);
nand U14883 (N_14883,N_13632,N_13855);
and U14884 (N_14884,N_13662,N_14116);
xor U14885 (N_14885,N_13832,N_13590);
nand U14886 (N_14886,N_13543,N_13604);
or U14887 (N_14887,N_14200,N_14143);
and U14888 (N_14888,N_14127,N_13715);
or U14889 (N_14889,N_13766,N_13884);
or U14890 (N_14890,N_14125,N_14099);
and U14891 (N_14891,N_14009,N_14156);
and U14892 (N_14892,N_13942,N_13764);
or U14893 (N_14893,N_14113,N_14009);
nand U14894 (N_14894,N_13620,N_13866);
nor U14895 (N_14895,N_13876,N_14230);
nand U14896 (N_14896,N_13571,N_14224);
or U14897 (N_14897,N_13882,N_13613);
nor U14898 (N_14898,N_14213,N_13644);
xnor U14899 (N_14899,N_13844,N_13984);
nor U14900 (N_14900,N_13897,N_14153);
and U14901 (N_14901,N_13524,N_13808);
nor U14902 (N_14902,N_13959,N_13823);
xnor U14903 (N_14903,N_13796,N_13504);
nor U14904 (N_14904,N_14001,N_13856);
or U14905 (N_14905,N_14227,N_14100);
or U14906 (N_14906,N_14147,N_13662);
nand U14907 (N_14907,N_14128,N_13603);
and U14908 (N_14908,N_13651,N_13793);
or U14909 (N_14909,N_13892,N_13763);
or U14910 (N_14910,N_13514,N_13604);
and U14911 (N_14911,N_13626,N_13625);
nor U14912 (N_14912,N_14024,N_14146);
or U14913 (N_14913,N_13978,N_13963);
xor U14914 (N_14914,N_13611,N_14188);
nand U14915 (N_14915,N_14182,N_14179);
nor U14916 (N_14916,N_13645,N_13752);
nand U14917 (N_14917,N_13685,N_13725);
nand U14918 (N_14918,N_14168,N_13923);
nand U14919 (N_14919,N_13621,N_13963);
nor U14920 (N_14920,N_13715,N_13593);
nor U14921 (N_14921,N_14015,N_13880);
nor U14922 (N_14922,N_13567,N_14015);
nand U14923 (N_14923,N_14135,N_14181);
nor U14924 (N_14924,N_14239,N_14163);
nand U14925 (N_14925,N_13678,N_14173);
and U14926 (N_14926,N_13918,N_13589);
nand U14927 (N_14927,N_14121,N_14114);
nand U14928 (N_14928,N_14004,N_13574);
and U14929 (N_14929,N_14249,N_14148);
or U14930 (N_14930,N_13919,N_13542);
or U14931 (N_14931,N_14173,N_13664);
nor U14932 (N_14932,N_13833,N_13739);
or U14933 (N_14933,N_13823,N_14191);
or U14934 (N_14934,N_14079,N_13749);
nor U14935 (N_14935,N_14190,N_13543);
nor U14936 (N_14936,N_14065,N_14010);
nor U14937 (N_14937,N_13781,N_14141);
nand U14938 (N_14938,N_13617,N_14114);
and U14939 (N_14939,N_14110,N_14243);
nor U14940 (N_14940,N_13800,N_13770);
nand U14941 (N_14941,N_13574,N_13589);
nand U14942 (N_14942,N_13655,N_13691);
nand U14943 (N_14943,N_14088,N_13912);
nand U14944 (N_14944,N_14242,N_14218);
nand U14945 (N_14945,N_13729,N_13894);
nor U14946 (N_14946,N_14033,N_13924);
or U14947 (N_14947,N_13776,N_13646);
or U14948 (N_14948,N_13623,N_13546);
and U14949 (N_14949,N_13712,N_14003);
nand U14950 (N_14950,N_14042,N_14125);
nor U14951 (N_14951,N_13691,N_13630);
nand U14952 (N_14952,N_14157,N_13850);
or U14953 (N_14953,N_13719,N_13982);
or U14954 (N_14954,N_13793,N_13857);
and U14955 (N_14955,N_13556,N_13513);
nor U14956 (N_14956,N_13702,N_13984);
nor U14957 (N_14957,N_13873,N_14157);
and U14958 (N_14958,N_14073,N_13658);
nor U14959 (N_14959,N_13919,N_14222);
nor U14960 (N_14960,N_13738,N_14105);
or U14961 (N_14961,N_14065,N_13755);
and U14962 (N_14962,N_14110,N_14233);
nor U14963 (N_14963,N_13907,N_13728);
and U14964 (N_14964,N_13994,N_13745);
nor U14965 (N_14965,N_13579,N_13814);
or U14966 (N_14966,N_13929,N_13595);
xor U14967 (N_14967,N_14057,N_13586);
nor U14968 (N_14968,N_13835,N_13819);
nor U14969 (N_14969,N_13862,N_14150);
nor U14970 (N_14970,N_14226,N_13707);
and U14971 (N_14971,N_14146,N_14003);
nor U14972 (N_14972,N_13616,N_14018);
or U14973 (N_14973,N_13599,N_13712);
nor U14974 (N_14974,N_14217,N_14219);
nor U14975 (N_14975,N_13646,N_14213);
nor U14976 (N_14976,N_13549,N_13537);
nand U14977 (N_14977,N_14154,N_13999);
nand U14978 (N_14978,N_14168,N_14064);
nor U14979 (N_14979,N_13960,N_14120);
and U14980 (N_14980,N_14151,N_13974);
nor U14981 (N_14981,N_13510,N_13734);
xor U14982 (N_14982,N_14188,N_13639);
or U14983 (N_14983,N_13948,N_14158);
and U14984 (N_14984,N_13661,N_13819);
and U14985 (N_14985,N_14073,N_14126);
nand U14986 (N_14986,N_14055,N_13763);
and U14987 (N_14987,N_14161,N_13622);
or U14988 (N_14988,N_14191,N_13579);
nand U14989 (N_14989,N_13882,N_13541);
and U14990 (N_14990,N_13956,N_14153);
or U14991 (N_14991,N_13961,N_13600);
or U14992 (N_14992,N_14132,N_13902);
or U14993 (N_14993,N_13856,N_13818);
nand U14994 (N_14994,N_14244,N_14073);
and U14995 (N_14995,N_13885,N_14217);
and U14996 (N_14996,N_13721,N_13865);
nand U14997 (N_14997,N_13628,N_13991);
and U14998 (N_14998,N_13820,N_14233);
or U14999 (N_14999,N_14160,N_13932);
or UO_0 (O_0,N_14790,N_14851);
nor UO_1 (O_1,N_14413,N_14883);
nand UO_2 (O_2,N_14256,N_14973);
and UO_3 (O_3,N_14745,N_14711);
nor UO_4 (O_4,N_14374,N_14697);
nor UO_5 (O_5,N_14926,N_14674);
xor UO_6 (O_6,N_14512,N_14972);
and UO_7 (O_7,N_14966,N_14971);
or UO_8 (O_8,N_14623,N_14569);
nor UO_9 (O_9,N_14500,N_14733);
and UO_10 (O_10,N_14616,N_14730);
nand UO_11 (O_11,N_14476,N_14905);
nor UO_12 (O_12,N_14408,N_14902);
or UO_13 (O_13,N_14968,N_14490);
nand UO_14 (O_14,N_14660,N_14329);
nor UO_15 (O_15,N_14554,N_14387);
or UO_16 (O_16,N_14867,N_14295);
nand UO_17 (O_17,N_14786,N_14946);
and UO_18 (O_18,N_14738,N_14301);
nand UO_19 (O_19,N_14510,N_14687);
nor UO_20 (O_20,N_14911,N_14705);
nand UO_21 (O_21,N_14322,N_14441);
and UO_22 (O_22,N_14662,N_14725);
or UO_23 (O_23,N_14773,N_14798);
nand UO_24 (O_24,N_14758,N_14896);
or UO_25 (O_25,N_14255,N_14586);
xnor UO_26 (O_26,N_14317,N_14970);
nor UO_27 (O_27,N_14346,N_14690);
and UO_28 (O_28,N_14478,N_14370);
and UO_29 (O_29,N_14986,N_14800);
and UO_30 (O_30,N_14678,N_14344);
or UO_31 (O_31,N_14348,N_14732);
nand UO_32 (O_32,N_14991,N_14382);
nor UO_33 (O_33,N_14856,N_14827);
nor UO_34 (O_34,N_14275,N_14866);
nor UO_35 (O_35,N_14661,N_14708);
or UO_36 (O_36,N_14843,N_14960);
or UO_37 (O_37,N_14753,N_14313);
or UO_38 (O_38,N_14840,N_14283);
nor UO_39 (O_39,N_14962,N_14625);
and UO_40 (O_40,N_14273,N_14629);
nor UO_41 (O_41,N_14521,N_14395);
nand UO_42 (O_42,N_14304,N_14760);
nand UO_43 (O_43,N_14543,N_14761);
nand UO_44 (O_44,N_14749,N_14872);
and UO_45 (O_45,N_14795,N_14701);
and UO_46 (O_46,N_14812,N_14292);
nor UO_47 (O_47,N_14784,N_14974);
nor UO_48 (O_48,N_14850,N_14864);
and UO_49 (O_49,N_14757,N_14855);
or UO_50 (O_50,N_14639,N_14552);
or UO_51 (O_51,N_14355,N_14405);
and UO_52 (O_52,N_14755,N_14744);
and UO_53 (O_53,N_14578,N_14963);
nor UO_54 (O_54,N_14652,N_14797);
nand UO_55 (O_55,N_14527,N_14734);
or UO_56 (O_56,N_14637,N_14858);
nor UO_57 (O_57,N_14445,N_14540);
or UO_58 (O_58,N_14716,N_14307);
or UO_59 (O_59,N_14516,N_14647);
nand UO_60 (O_60,N_14293,N_14710);
and UO_61 (O_61,N_14547,N_14923);
nor UO_62 (O_62,N_14717,N_14581);
and UO_63 (O_63,N_14965,N_14912);
nand UO_64 (O_64,N_14494,N_14465);
and UO_65 (O_65,N_14916,N_14781);
nor UO_66 (O_66,N_14859,N_14961);
nand UO_67 (O_67,N_14453,N_14567);
and UO_68 (O_68,N_14604,N_14615);
or UO_69 (O_69,N_14895,N_14650);
nand UO_70 (O_70,N_14993,N_14544);
nor UO_71 (O_71,N_14303,N_14684);
or UO_72 (O_72,N_14836,N_14828);
nand UO_73 (O_73,N_14357,N_14680);
nand UO_74 (O_74,N_14549,N_14546);
nor UO_75 (O_75,N_14854,N_14466);
nand UO_76 (O_76,N_14253,N_14898);
or UO_77 (O_77,N_14954,N_14979);
and UO_78 (O_78,N_14443,N_14940);
and UO_79 (O_79,N_14311,N_14664);
and UO_80 (O_80,N_14978,N_14523);
nor UO_81 (O_81,N_14642,N_14358);
nand UO_82 (O_82,N_14285,N_14340);
nor UO_83 (O_83,N_14553,N_14673);
xor UO_84 (O_84,N_14702,N_14967);
and UO_85 (O_85,N_14868,N_14341);
nor UO_86 (O_86,N_14485,N_14522);
and UO_87 (O_87,N_14372,N_14832);
xor UO_88 (O_88,N_14474,N_14666);
or UO_89 (O_89,N_14506,N_14281);
and UO_90 (O_90,N_14752,N_14998);
nand UO_91 (O_91,N_14767,N_14406);
nor UO_92 (O_92,N_14556,N_14955);
nor UO_93 (O_93,N_14751,N_14486);
and UO_94 (O_94,N_14918,N_14507);
and UO_95 (O_95,N_14397,N_14645);
and UO_96 (O_96,N_14739,N_14729);
or UO_97 (O_97,N_14468,N_14719);
and UO_98 (O_98,N_14877,N_14462);
and UO_99 (O_99,N_14876,N_14457);
or UO_100 (O_100,N_14252,N_14721);
nor UO_101 (O_101,N_14422,N_14391);
or UO_102 (O_102,N_14538,N_14614);
nor UO_103 (O_103,N_14658,N_14446);
nand UO_104 (O_104,N_14309,N_14934);
xnor UO_105 (O_105,N_14885,N_14349);
or UO_106 (O_106,N_14712,N_14321);
or UO_107 (O_107,N_14250,N_14557);
and UO_108 (O_108,N_14780,N_14617);
xnor UO_109 (O_109,N_14822,N_14805);
and UO_110 (O_110,N_14342,N_14499);
or UO_111 (O_111,N_14359,N_14682);
or UO_112 (O_112,N_14772,N_14897);
or UO_113 (O_113,N_14597,N_14601);
nand UO_114 (O_114,N_14891,N_14371);
or UO_115 (O_115,N_14437,N_14939);
nor UO_116 (O_116,N_14996,N_14699);
nand UO_117 (O_117,N_14904,N_14361);
nand UO_118 (O_118,N_14400,N_14802);
or UO_119 (O_119,N_14381,N_14770);
or UO_120 (O_120,N_14644,N_14439);
and UO_121 (O_121,N_14456,N_14913);
nor UO_122 (O_122,N_14718,N_14525);
xor UO_123 (O_123,N_14427,N_14548);
and UO_124 (O_124,N_14769,N_14299);
nor UO_125 (O_125,N_14590,N_14407);
or UO_126 (O_126,N_14768,N_14574);
nand UO_127 (O_127,N_14881,N_14793);
nor UO_128 (O_128,N_14670,N_14871);
nand UO_129 (O_129,N_14845,N_14630);
nand UO_130 (O_130,N_14448,N_14353);
and UO_131 (O_131,N_14583,N_14611);
and UO_132 (O_132,N_14539,N_14620);
nor UO_133 (O_133,N_14860,N_14917);
or UO_134 (O_134,N_14847,N_14906);
nand UO_135 (O_135,N_14584,N_14260);
or UO_136 (O_136,N_14354,N_14862);
nor UO_137 (O_137,N_14811,N_14541);
and UO_138 (O_138,N_14915,N_14338);
or UO_139 (O_139,N_14640,N_14975);
or UO_140 (O_140,N_14345,N_14312);
nor UO_141 (O_141,N_14766,N_14818);
xor UO_142 (O_142,N_14560,N_14429);
or UO_143 (O_143,N_14782,N_14376);
nand UO_144 (O_144,N_14264,N_14930);
and UO_145 (O_145,N_14924,N_14835);
xor UO_146 (O_146,N_14430,N_14715);
nand UO_147 (O_147,N_14631,N_14933);
nor UO_148 (O_148,N_14756,N_14657);
nor UO_149 (O_149,N_14424,N_14839);
and UO_150 (O_150,N_14771,N_14692);
and UO_151 (O_151,N_14691,N_14450);
nand UO_152 (O_152,N_14816,N_14663);
nor UO_153 (O_153,N_14505,N_14580);
or UO_154 (O_154,N_14689,N_14438);
nor UO_155 (O_155,N_14774,N_14696);
and UO_156 (O_156,N_14988,N_14792);
and UO_157 (O_157,N_14368,N_14587);
or UO_158 (O_158,N_14987,N_14762);
nand UO_159 (O_159,N_14727,N_14641);
xor UO_160 (O_160,N_14347,N_14783);
nor UO_161 (O_161,N_14598,N_14633);
and UO_162 (O_162,N_14364,N_14314);
nand UO_163 (O_163,N_14722,N_14935);
or UO_164 (O_164,N_14621,N_14509);
nor UO_165 (O_165,N_14679,N_14706);
or UO_166 (O_166,N_14251,N_14296);
nand UO_167 (O_167,N_14903,N_14573);
and UO_168 (O_168,N_14852,N_14334);
xor UO_169 (O_169,N_14272,N_14740);
nand UO_170 (O_170,N_14654,N_14263);
and UO_171 (O_171,N_14414,N_14817);
nor UO_172 (O_172,N_14579,N_14681);
or UO_173 (O_173,N_14600,N_14735);
nand UO_174 (O_174,N_14534,N_14473);
and UO_175 (O_175,N_14984,N_14393);
or UO_176 (O_176,N_14571,N_14801);
nor UO_177 (O_177,N_14724,N_14919);
nand UO_178 (O_178,N_14981,N_14291);
and UO_179 (O_179,N_14594,N_14305);
and UO_180 (O_180,N_14375,N_14269);
nor UO_181 (O_181,N_14532,N_14791);
and UO_182 (O_182,N_14308,N_14677);
nand UO_183 (O_183,N_14373,N_14969);
and UO_184 (O_184,N_14964,N_14636);
nor UO_185 (O_185,N_14700,N_14537);
xor UO_186 (O_186,N_14565,N_14433);
nor UO_187 (O_187,N_14297,N_14831);
and UO_188 (O_188,N_14432,N_14813);
nor UO_189 (O_189,N_14412,N_14488);
nand UO_190 (O_190,N_14524,N_14363);
xor UO_191 (O_191,N_14563,N_14316);
nand UO_192 (O_192,N_14794,N_14695);
or UO_193 (O_193,N_14280,N_14460);
nand UO_194 (O_194,N_14815,N_14775);
or UO_195 (O_195,N_14997,N_14992);
and UO_196 (O_196,N_14814,N_14779);
nor UO_197 (O_197,N_14288,N_14282);
or UO_198 (O_198,N_14515,N_14471);
or UO_199 (O_199,N_14356,N_14315);
nor UO_200 (O_200,N_14572,N_14907);
and UO_201 (O_201,N_14953,N_14990);
and UO_202 (O_202,N_14884,N_14807);
nor UO_203 (O_203,N_14958,N_14931);
nand UO_204 (O_204,N_14665,N_14886);
or UO_205 (O_205,N_14746,N_14469);
or UO_206 (O_206,N_14632,N_14577);
nand UO_207 (O_207,N_14276,N_14526);
nand UO_208 (O_208,N_14319,N_14480);
xor UO_209 (O_209,N_14452,N_14863);
and UO_210 (O_210,N_14849,N_14945);
or UO_211 (O_211,N_14952,N_14893);
nor UO_212 (O_212,N_14592,N_14809);
and UO_213 (O_213,N_14846,N_14367);
nor UO_214 (O_214,N_14325,N_14726);
nor UO_215 (O_215,N_14634,N_14378);
nand UO_216 (O_216,N_14651,N_14489);
nand UO_217 (O_217,N_14709,N_14390);
xnor UO_218 (O_218,N_14351,N_14550);
nor UO_219 (O_219,N_14459,N_14418);
and UO_220 (O_220,N_14423,N_14901);
or UO_221 (O_221,N_14582,N_14741);
or UO_222 (O_222,N_14808,N_14983);
nor UO_223 (O_223,N_14834,N_14461);
nand UO_224 (O_224,N_14910,N_14938);
nor UO_225 (O_225,N_14564,N_14360);
and UO_226 (O_226,N_14982,N_14638);
nor UO_227 (O_227,N_14530,N_14747);
nor UO_228 (O_228,N_14607,N_14880);
and UO_229 (O_229,N_14326,N_14323);
or UO_230 (O_230,N_14415,N_14501);
and UO_231 (O_231,N_14261,N_14384);
nor UO_232 (O_232,N_14514,N_14482);
and UO_233 (O_233,N_14622,N_14610);
or UO_234 (O_234,N_14436,N_14873);
and UO_235 (O_235,N_14558,N_14300);
nor UO_236 (O_236,N_14442,N_14754);
and UO_237 (O_237,N_14824,N_14704);
nor UO_238 (O_238,N_14908,N_14421);
or UO_239 (O_239,N_14268,N_14287);
nor UO_240 (O_240,N_14612,N_14402);
nand UO_241 (O_241,N_14551,N_14948);
nand UO_242 (O_242,N_14343,N_14942);
and UO_243 (O_243,N_14936,N_14330);
nor UO_244 (O_244,N_14520,N_14545);
or UO_245 (O_245,N_14528,N_14737);
or UO_246 (O_246,N_14324,N_14602);
or UO_247 (O_247,N_14417,N_14892);
nor UO_248 (O_248,N_14535,N_14675);
or UO_249 (O_249,N_14366,N_14404);
and UO_250 (O_250,N_14869,N_14799);
nand UO_251 (O_251,N_14603,N_14561);
nand UO_252 (O_252,N_14497,N_14492);
or UO_253 (O_253,N_14266,N_14267);
nand UO_254 (O_254,N_14686,N_14257);
xnor UO_255 (O_255,N_14643,N_14508);
nor UO_256 (O_256,N_14830,N_14380);
and UO_257 (O_257,N_14444,N_14927);
nand UO_258 (O_258,N_14826,N_14454);
nand UO_259 (O_259,N_14882,N_14591);
nand UO_260 (O_260,N_14742,N_14925);
or UO_261 (O_261,N_14626,N_14498);
nor UO_262 (O_262,N_14608,N_14928);
nor UO_263 (O_263,N_14589,N_14467);
nand UO_264 (O_264,N_14995,N_14890);
and UO_265 (O_265,N_14286,N_14483);
and UO_266 (O_266,N_14861,N_14331);
or UO_267 (O_267,N_14932,N_14947);
nor UO_268 (O_268,N_14878,N_14401);
nand UO_269 (O_269,N_14796,N_14416);
and UO_270 (O_270,N_14409,N_14504);
or UO_271 (O_271,N_14676,N_14750);
and UO_272 (O_272,N_14669,N_14555);
nor UO_273 (O_273,N_14277,N_14875);
or UO_274 (O_274,N_14328,N_14479);
nand UO_275 (O_275,N_14688,N_14865);
and UO_276 (O_276,N_14278,N_14369);
or UO_277 (O_277,N_14458,N_14956);
nor UO_278 (O_278,N_14672,N_14656);
nor UO_279 (O_279,N_14698,N_14804);
nand UO_280 (O_280,N_14274,N_14435);
and UO_281 (O_281,N_14655,N_14398);
nand UO_282 (O_282,N_14542,N_14477);
nand UO_283 (O_283,N_14517,N_14491);
nand UO_284 (O_284,N_14713,N_14562);
nor UO_285 (O_285,N_14909,N_14289);
or UO_286 (O_286,N_14844,N_14270);
or UO_287 (O_287,N_14627,N_14985);
nor UO_288 (O_288,N_14659,N_14759);
xor UO_289 (O_289,N_14671,N_14944);
nor UO_290 (O_290,N_14821,N_14887);
and UO_291 (O_291,N_14743,N_14352);
nand UO_292 (O_292,N_14829,N_14874);
nand UO_293 (O_293,N_14624,N_14254);
nor UO_294 (O_294,N_14857,N_14994);
nand UO_295 (O_295,N_14842,N_14529);
nor UO_296 (O_296,N_14399,N_14487);
nor UO_297 (O_297,N_14628,N_14989);
and UO_298 (O_298,N_14394,N_14320);
nor UO_299 (O_299,N_14837,N_14502);
or UO_300 (O_300,N_14833,N_14588);
nand UO_301 (O_301,N_14720,N_14332);
nand UO_302 (O_302,N_14685,N_14511);
or UO_303 (O_303,N_14362,N_14447);
or UO_304 (O_304,N_14888,N_14379);
and UO_305 (O_305,N_14464,N_14568);
nand UO_306 (O_306,N_14976,N_14449);
and UO_307 (O_307,N_14959,N_14787);
or UO_308 (O_308,N_14957,N_14294);
nor UO_309 (O_309,N_14765,N_14570);
nor UO_310 (O_310,N_14694,N_14778);
or UO_311 (O_311,N_14853,N_14425);
nand UO_312 (O_312,N_14302,N_14619);
or UO_313 (O_313,N_14377,N_14870);
nor UO_314 (O_314,N_14518,N_14820);
and UO_315 (O_315,N_14493,N_14403);
or UO_316 (O_316,N_14823,N_14599);
nor UO_317 (O_317,N_14575,N_14764);
nor UO_318 (O_318,N_14419,N_14503);
or UO_319 (O_319,N_14365,N_14475);
or UO_320 (O_320,N_14980,N_14310);
or UO_321 (O_321,N_14949,N_14595);
and UO_322 (O_322,N_14290,N_14977);
and UO_323 (O_323,N_14336,N_14396);
nor UO_324 (O_324,N_14566,N_14484);
nor UO_325 (O_325,N_14848,N_14776);
nand UO_326 (O_326,N_14819,N_14728);
nor UO_327 (O_327,N_14585,N_14736);
and UO_328 (O_328,N_14879,N_14922);
and UO_329 (O_329,N_14411,N_14386);
or UO_330 (O_330,N_14618,N_14388);
or UO_331 (O_331,N_14606,N_14306);
nand UO_332 (O_332,N_14941,N_14455);
nand UO_333 (O_333,N_14279,N_14649);
nand UO_334 (O_334,N_14383,N_14810);
xnor UO_335 (O_335,N_14259,N_14788);
and UO_336 (O_336,N_14533,N_14265);
and UO_337 (O_337,N_14648,N_14333);
nand UO_338 (O_338,N_14668,N_14519);
and UO_339 (O_339,N_14667,N_14803);
nand UO_340 (O_340,N_14298,N_14440);
nor UO_341 (O_341,N_14481,N_14596);
or UO_342 (O_342,N_14613,N_14899);
nand UO_343 (O_343,N_14937,N_14763);
nand UO_344 (O_344,N_14536,N_14531);
nor UO_345 (O_345,N_14463,N_14605);
nand UO_346 (O_346,N_14339,N_14841);
nand UO_347 (O_347,N_14559,N_14693);
nand UO_348 (O_348,N_14789,N_14825);
nand UO_349 (O_349,N_14284,N_14426);
nor UO_350 (O_350,N_14495,N_14496);
and UO_351 (O_351,N_14723,N_14950);
nor UO_352 (O_352,N_14806,N_14335);
and UO_353 (O_353,N_14318,N_14748);
nor UO_354 (O_354,N_14894,N_14777);
and UO_355 (O_355,N_14434,N_14327);
or UO_356 (O_356,N_14576,N_14350);
nand UO_357 (O_357,N_14707,N_14714);
and UO_358 (O_358,N_14943,N_14785);
nand UO_359 (O_359,N_14431,N_14258);
and UO_360 (O_360,N_14472,N_14900);
or UO_361 (O_361,N_14731,N_14635);
nand UO_362 (O_362,N_14921,N_14420);
or UO_363 (O_363,N_14914,N_14951);
nand UO_364 (O_364,N_14410,N_14889);
nand UO_365 (O_365,N_14470,N_14385);
and UO_366 (O_366,N_14262,N_14929);
or UO_367 (O_367,N_14451,N_14609);
nor UO_368 (O_368,N_14392,N_14703);
nor UO_369 (O_369,N_14428,N_14920);
nand UO_370 (O_370,N_14513,N_14389);
nand UO_371 (O_371,N_14271,N_14838);
nor UO_372 (O_372,N_14593,N_14683);
nor UO_373 (O_373,N_14999,N_14646);
nand UO_374 (O_374,N_14653,N_14337);
and UO_375 (O_375,N_14380,N_14326);
nor UO_376 (O_376,N_14623,N_14486);
or UO_377 (O_377,N_14387,N_14676);
nor UO_378 (O_378,N_14684,N_14933);
xor UO_379 (O_379,N_14819,N_14668);
or UO_380 (O_380,N_14755,N_14399);
nor UO_381 (O_381,N_14441,N_14679);
nand UO_382 (O_382,N_14559,N_14251);
nor UO_383 (O_383,N_14903,N_14531);
nor UO_384 (O_384,N_14697,N_14653);
or UO_385 (O_385,N_14255,N_14652);
or UO_386 (O_386,N_14808,N_14698);
or UO_387 (O_387,N_14307,N_14729);
or UO_388 (O_388,N_14845,N_14867);
or UO_389 (O_389,N_14257,N_14864);
nor UO_390 (O_390,N_14835,N_14512);
and UO_391 (O_391,N_14911,N_14268);
nand UO_392 (O_392,N_14559,N_14910);
nand UO_393 (O_393,N_14515,N_14801);
nor UO_394 (O_394,N_14912,N_14469);
nand UO_395 (O_395,N_14819,N_14857);
or UO_396 (O_396,N_14586,N_14641);
or UO_397 (O_397,N_14444,N_14610);
nor UO_398 (O_398,N_14803,N_14793);
nor UO_399 (O_399,N_14898,N_14874);
nor UO_400 (O_400,N_14632,N_14826);
xnor UO_401 (O_401,N_14711,N_14719);
nor UO_402 (O_402,N_14276,N_14454);
or UO_403 (O_403,N_14390,N_14266);
nor UO_404 (O_404,N_14558,N_14666);
or UO_405 (O_405,N_14339,N_14745);
nor UO_406 (O_406,N_14638,N_14408);
nor UO_407 (O_407,N_14723,N_14319);
nor UO_408 (O_408,N_14637,N_14873);
and UO_409 (O_409,N_14838,N_14456);
nand UO_410 (O_410,N_14568,N_14701);
and UO_411 (O_411,N_14977,N_14914);
and UO_412 (O_412,N_14420,N_14894);
and UO_413 (O_413,N_14623,N_14911);
and UO_414 (O_414,N_14308,N_14688);
and UO_415 (O_415,N_14841,N_14762);
or UO_416 (O_416,N_14536,N_14339);
nor UO_417 (O_417,N_14443,N_14777);
nor UO_418 (O_418,N_14624,N_14960);
nand UO_419 (O_419,N_14555,N_14861);
nor UO_420 (O_420,N_14827,N_14364);
nor UO_421 (O_421,N_14976,N_14309);
nor UO_422 (O_422,N_14268,N_14611);
nor UO_423 (O_423,N_14302,N_14553);
nand UO_424 (O_424,N_14550,N_14934);
nand UO_425 (O_425,N_14759,N_14332);
and UO_426 (O_426,N_14413,N_14919);
nor UO_427 (O_427,N_14335,N_14452);
and UO_428 (O_428,N_14417,N_14535);
or UO_429 (O_429,N_14944,N_14512);
nand UO_430 (O_430,N_14914,N_14955);
or UO_431 (O_431,N_14763,N_14469);
and UO_432 (O_432,N_14482,N_14887);
and UO_433 (O_433,N_14372,N_14350);
nor UO_434 (O_434,N_14825,N_14958);
or UO_435 (O_435,N_14929,N_14443);
or UO_436 (O_436,N_14943,N_14869);
or UO_437 (O_437,N_14725,N_14688);
nand UO_438 (O_438,N_14908,N_14783);
nor UO_439 (O_439,N_14744,N_14957);
nor UO_440 (O_440,N_14615,N_14333);
or UO_441 (O_441,N_14387,N_14738);
and UO_442 (O_442,N_14885,N_14931);
nand UO_443 (O_443,N_14455,N_14755);
nand UO_444 (O_444,N_14821,N_14320);
and UO_445 (O_445,N_14910,N_14422);
and UO_446 (O_446,N_14374,N_14716);
or UO_447 (O_447,N_14932,N_14503);
nor UO_448 (O_448,N_14368,N_14990);
or UO_449 (O_449,N_14792,N_14251);
or UO_450 (O_450,N_14269,N_14405);
or UO_451 (O_451,N_14263,N_14450);
or UO_452 (O_452,N_14772,N_14371);
nand UO_453 (O_453,N_14800,N_14675);
nor UO_454 (O_454,N_14708,N_14691);
nand UO_455 (O_455,N_14515,N_14844);
nand UO_456 (O_456,N_14951,N_14625);
nor UO_457 (O_457,N_14400,N_14427);
or UO_458 (O_458,N_14691,N_14564);
and UO_459 (O_459,N_14950,N_14697);
nand UO_460 (O_460,N_14859,N_14343);
nor UO_461 (O_461,N_14444,N_14675);
nor UO_462 (O_462,N_14595,N_14777);
or UO_463 (O_463,N_14417,N_14826);
or UO_464 (O_464,N_14741,N_14419);
or UO_465 (O_465,N_14556,N_14392);
nand UO_466 (O_466,N_14382,N_14533);
and UO_467 (O_467,N_14817,N_14990);
nor UO_468 (O_468,N_14571,N_14553);
nor UO_469 (O_469,N_14979,N_14469);
and UO_470 (O_470,N_14933,N_14355);
and UO_471 (O_471,N_14372,N_14336);
and UO_472 (O_472,N_14300,N_14613);
or UO_473 (O_473,N_14465,N_14418);
nor UO_474 (O_474,N_14577,N_14739);
or UO_475 (O_475,N_14337,N_14972);
nor UO_476 (O_476,N_14544,N_14506);
and UO_477 (O_477,N_14676,N_14748);
and UO_478 (O_478,N_14635,N_14602);
or UO_479 (O_479,N_14991,N_14348);
or UO_480 (O_480,N_14837,N_14739);
nand UO_481 (O_481,N_14335,N_14920);
and UO_482 (O_482,N_14547,N_14366);
nand UO_483 (O_483,N_14780,N_14599);
or UO_484 (O_484,N_14788,N_14985);
or UO_485 (O_485,N_14301,N_14811);
nor UO_486 (O_486,N_14927,N_14806);
and UO_487 (O_487,N_14458,N_14943);
nand UO_488 (O_488,N_14594,N_14663);
nor UO_489 (O_489,N_14686,N_14611);
nor UO_490 (O_490,N_14760,N_14295);
and UO_491 (O_491,N_14401,N_14810);
nor UO_492 (O_492,N_14429,N_14398);
and UO_493 (O_493,N_14629,N_14760);
nand UO_494 (O_494,N_14975,N_14904);
and UO_495 (O_495,N_14631,N_14476);
xor UO_496 (O_496,N_14466,N_14430);
or UO_497 (O_497,N_14770,N_14796);
nand UO_498 (O_498,N_14554,N_14823);
nor UO_499 (O_499,N_14251,N_14885);
nor UO_500 (O_500,N_14596,N_14741);
or UO_501 (O_501,N_14749,N_14408);
or UO_502 (O_502,N_14251,N_14723);
and UO_503 (O_503,N_14751,N_14262);
nor UO_504 (O_504,N_14855,N_14717);
nor UO_505 (O_505,N_14516,N_14876);
or UO_506 (O_506,N_14264,N_14294);
or UO_507 (O_507,N_14386,N_14456);
nor UO_508 (O_508,N_14834,N_14320);
nor UO_509 (O_509,N_14626,N_14743);
nand UO_510 (O_510,N_14588,N_14882);
nand UO_511 (O_511,N_14652,N_14727);
nor UO_512 (O_512,N_14366,N_14768);
nand UO_513 (O_513,N_14845,N_14403);
and UO_514 (O_514,N_14919,N_14847);
and UO_515 (O_515,N_14276,N_14257);
nor UO_516 (O_516,N_14252,N_14868);
or UO_517 (O_517,N_14716,N_14880);
or UO_518 (O_518,N_14572,N_14322);
or UO_519 (O_519,N_14622,N_14351);
and UO_520 (O_520,N_14296,N_14813);
nor UO_521 (O_521,N_14584,N_14442);
nor UO_522 (O_522,N_14303,N_14345);
nor UO_523 (O_523,N_14552,N_14841);
nor UO_524 (O_524,N_14499,N_14374);
or UO_525 (O_525,N_14489,N_14323);
and UO_526 (O_526,N_14931,N_14814);
and UO_527 (O_527,N_14634,N_14254);
nand UO_528 (O_528,N_14315,N_14413);
nor UO_529 (O_529,N_14439,N_14807);
nor UO_530 (O_530,N_14870,N_14469);
and UO_531 (O_531,N_14924,N_14257);
nor UO_532 (O_532,N_14643,N_14604);
or UO_533 (O_533,N_14770,N_14919);
nor UO_534 (O_534,N_14351,N_14648);
nand UO_535 (O_535,N_14939,N_14403);
or UO_536 (O_536,N_14900,N_14709);
nand UO_537 (O_537,N_14650,N_14576);
and UO_538 (O_538,N_14438,N_14668);
and UO_539 (O_539,N_14386,N_14881);
nand UO_540 (O_540,N_14371,N_14829);
or UO_541 (O_541,N_14522,N_14649);
or UO_542 (O_542,N_14715,N_14469);
nor UO_543 (O_543,N_14610,N_14419);
xnor UO_544 (O_544,N_14331,N_14788);
nor UO_545 (O_545,N_14666,N_14885);
or UO_546 (O_546,N_14787,N_14347);
nand UO_547 (O_547,N_14728,N_14603);
and UO_548 (O_548,N_14300,N_14504);
nand UO_549 (O_549,N_14265,N_14302);
nand UO_550 (O_550,N_14335,N_14608);
nand UO_551 (O_551,N_14513,N_14309);
nor UO_552 (O_552,N_14328,N_14911);
nor UO_553 (O_553,N_14976,N_14633);
nand UO_554 (O_554,N_14605,N_14716);
xor UO_555 (O_555,N_14274,N_14343);
or UO_556 (O_556,N_14915,N_14696);
nand UO_557 (O_557,N_14621,N_14976);
nand UO_558 (O_558,N_14935,N_14919);
or UO_559 (O_559,N_14774,N_14326);
nor UO_560 (O_560,N_14280,N_14521);
or UO_561 (O_561,N_14498,N_14917);
nand UO_562 (O_562,N_14953,N_14550);
and UO_563 (O_563,N_14350,N_14575);
nand UO_564 (O_564,N_14610,N_14817);
and UO_565 (O_565,N_14442,N_14992);
nand UO_566 (O_566,N_14933,N_14922);
and UO_567 (O_567,N_14332,N_14985);
nand UO_568 (O_568,N_14315,N_14285);
nor UO_569 (O_569,N_14424,N_14767);
nand UO_570 (O_570,N_14731,N_14780);
nand UO_571 (O_571,N_14497,N_14596);
or UO_572 (O_572,N_14266,N_14523);
nand UO_573 (O_573,N_14321,N_14425);
and UO_574 (O_574,N_14948,N_14552);
and UO_575 (O_575,N_14418,N_14735);
nand UO_576 (O_576,N_14768,N_14808);
nand UO_577 (O_577,N_14882,N_14957);
and UO_578 (O_578,N_14374,N_14641);
nor UO_579 (O_579,N_14306,N_14665);
and UO_580 (O_580,N_14319,N_14293);
nor UO_581 (O_581,N_14327,N_14906);
and UO_582 (O_582,N_14811,N_14929);
or UO_583 (O_583,N_14255,N_14977);
and UO_584 (O_584,N_14407,N_14526);
xnor UO_585 (O_585,N_14435,N_14781);
nor UO_586 (O_586,N_14423,N_14751);
and UO_587 (O_587,N_14332,N_14304);
nor UO_588 (O_588,N_14982,N_14761);
nor UO_589 (O_589,N_14669,N_14642);
or UO_590 (O_590,N_14364,N_14700);
or UO_591 (O_591,N_14772,N_14713);
nor UO_592 (O_592,N_14507,N_14294);
and UO_593 (O_593,N_14434,N_14772);
and UO_594 (O_594,N_14436,N_14341);
or UO_595 (O_595,N_14834,N_14289);
or UO_596 (O_596,N_14451,N_14926);
or UO_597 (O_597,N_14597,N_14887);
or UO_598 (O_598,N_14765,N_14256);
or UO_599 (O_599,N_14460,N_14952);
nor UO_600 (O_600,N_14450,N_14744);
nand UO_601 (O_601,N_14399,N_14886);
nand UO_602 (O_602,N_14364,N_14633);
or UO_603 (O_603,N_14307,N_14864);
and UO_604 (O_604,N_14542,N_14373);
nand UO_605 (O_605,N_14530,N_14743);
nor UO_606 (O_606,N_14471,N_14665);
nor UO_607 (O_607,N_14912,N_14466);
and UO_608 (O_608,N_14709,N_14579);
nor UO_609 (O_609,N_14839,N_14440);
and UO_610 (O_610,N_14707,N_14516);
nand UO_611 (O_611,N_14549,N_14494);
and UO_612 (O_612,N_14493,N_14325);
or UO_613 (O_613,N_14723,N_14810);
nor UO_614 (O_614,N_14634,N_14684);
and UO_615 (O_615,N_14301,N_14963);
nand UO_616 (O_616,N_14604,N_14454);
or UO_617 (O_617,N_14969,N_14983);
and UO_618 (O_618,N_14987,N_14807);
or UO_619 (O_619,N_14892,N_14459);
and UO_620 (O_620,N_14472,N_14657);
nor UO_621 (O_621,N_14324,N_14842);
and UO_622 (O_622,N_14508,N_14921);
and UO_623 (O_623,N_14388,N_14515);
nand UO_624 (O_624,N_14812,N_14608);
nor UO_625 (O_625,N_14383,N_14377);
or UO_626 (O_626,N_14491,N_14881);
or UO_627 (O_627,N_14389,N_14809);
nand UO_628 (O_628,N_14520,N_14549);
and UO_629 (O_629,N_14693,N_14744);
nor UO_630 (O_630,N_14856,N_14336);
or UO_631 (O_631,N_14374,N_14831);
nor UO_632 (O_632,N_14600,N_14597);
or UO_633 (O_633,N_14946,N_14353);
nand UO_634 (O_634,N_14983,N_14270);
nand UO_635 (O_635,N_14862,N_14694);
or UO_636 (O_636,N_14594,N_14791);
nor UO_637 (O_637,N_14344,N_14302);
nor UO_638 (O_638,N_14542,N_14605);
or UO_639 (O_639,N_14555,N_14989);
nand UO_640 (O_640,N_14706,N_14648);
and UO_641 (O_641,N_14854,N_14331);
nand UO_642 (O_642,N_14721,N_14504);
xor UO_643 (O_643,N_14494,N_14688);
nor UO_644 (O_644,N_14838,N_14713);
nand UO_645 (O_645,N_14641,N_14366);
xnor UO_646 (O_646,N_14457,N_14330);
and UO_647 (O_647,N_14293,N_14639);
nor UO_648 (O_648,N_14446,N_14400);
nand UO_649 (O_649,N_14768,N_14478);
nor UO_650 (O_650,N_14959,N_14681);
or UO_651 (O_651,N_14782,N_14771);
nand UO_652 (O_652,N_14418,N_14766);
nor UO_653 (O_653,N_14272,N_14577);
or UO_654 (O_654,N_14505,N_14256);
and UO_655 (O_655,N_14314,N_14390);
and UO_656 (O_656,N_14971,N_14572);
or UO_657 (O_657,N_14876,N_14892);
and UO_658 (O_658,N_14359,N_14523);
and UO_659 (O_659,N_14433,N_14956);
or UO_660 (O_660,N_14680,N_14454);
nor UO_661 (O_661,N_14789,N_14605);
nor UO_662 (O_662,N_14282,N_14571);
nand UO_663 (O_663,N_14514,N_14447);
and UO_664 (O_664,N_14589,N_14949);
nand UO_665 (O_665,N_14494,N_14359);
nor UO_666 (O_666,N_14368,N_14767);
nor UO_667 (O_667,N_14425,N_14459);
and UO_668 (O_668,N_14984,N_14369);
and UO_669 (O_669,N_14941,N_14785);
nor UO_670 (O_670,N_14971,N_14657);
nor UO_671 (O_671,N_14676,N_14502);
or UO_672 (O_672,N_14520,N_14634);
nor UO_673 (O_673,N_14386,N_14590);
or UO_674 (O_674,N_14978,N_14298);
nand UO_675 (O_675,N_14335,N_14514);
nor UO_676 (O_676,N_14655,N_14631);
nor UO_677 (O_677,N_14325,N_14954);
and UO_678 (O_678,N_14494,N_14351);
or UO_679 (O_679,N_14991,N_14900);
nand UO_680 (O_680,N_14751,N_14719);
and UO_681 (O_681,N_14962,N_14690);
nand UO_682 (O_682,N_14581,N_14821);
or UO_683 (O_683,N_14923,N_14886);
nor UO_684 (O_684,N_14535,N_14747);
and UO_685 (O_685,N_14302,N_14251);
nand UO_686 (O_686,N_14900,N_14426);
and UO_687 (O_687,N_14806,N_14965);
and UO_688 (O_688,N_14602,N_14791);
nor UO_689 (O_689,N_14775,N_14842);
nor UO_690 (O_690,N_14294,N_14870);
or UO_691 (O_691,N_14471,N_14925);
nand UO_692 (O_692,N_14536,N_14469);
nor UO_693 (O_693,N_14825,N_14281);
nand UO_694 (O_694,N_14707,N_14431);
nor UO_695 (O_695,N_14252,N_14750);
or UO_696 (O_696,N_14574,N_14868);
nor UO_697 (O_697,N_14739,N_14473);
or UO_698 (O_698,N_14557,N_14758);
xnor UO_699 (O_699,N_14484,N_14561);
nand UO_700 (O_700,N_14324,N_14274);
nand UO_701 (O_701,N_14810,N_14819);
or UO_702 (O_702,N_14688,N_14624);
nand UO_703 (O_703,N_14679,N_14558);
and UO_704 (O_704,N_14455,N_14724);
or UO_705 (O_705,N_14892,N_14954);
and UO_706 (O_706,N_14368,N_14981);
or UO_707 (O_707,N_14499,N_14603);
nor UO_708 (O_708,N_14919,N_14260);
or UO_709 (O_709,N_14839,N_14253);
or UO_710 (O_710,N_14282,N_14354);
nand UO_711 (O_711,N_14788,N_14438);
or UO_712 (O_712,N_14560,N_14505);
nand UO_713 (O_713,N_14859,N_14393);
and UO_714 (O_714,N_14583,N_14322);
or UO_715 (O_715,N_14720,N_14830);
or UO_716 (O_716,N_14453,N_14446);
or UO_717 (O_717,N_14965,N_14930);
and UO_718 (O_718,N_14550,N_14594);
or UO_719 (O_719,N_14497,N_14264);
and UO_720 (O_720,N_14320,N_14779);
nand UO_721 (O_721,N_14622,N_14536);
nor UO_722 (O_722,N_14257,N_14645);
or UO_723 (O_723,N_14353,N_14920);
or UO_724 (O_724,N_14838,N_14625);
nor UO_725 (O_725,N_14565,N_14813);
and UO_726 (O_726,N_14705,N_14893);
nor UO_727 (O_727,N_14830,N_14786);
nand UO_728 (O_728,N_14362,N_14590);
nor UO_729 (O_729,N_14953,N_14621);
and UO_730 (O_730,N_14614,N_14610);
or UO_731 (O_731,N_14731,N_14537);
xnor UO_732 (O_732,N_14421,N_14699);
and UO_733 (O_733,N_14982,N_14272);
nand UO_734 (O_734,N_14772,N_14601);
or UO_735 (O_735,N_14622,N_14448);
and UO_736 (O_736,N_14876,N_14643);
and UO_737 (O_737,N_14746,N_14733);
or UO_738 (O_738,N_14481,N_14343);
or UO_739 (O_739,N_14655,N_14983);
and UO_740 (O_740,N_14258,N_14675);
nor UO_741 (O_741,N_14715,N_14306);
or UO_742 (O_742,N_14327,N_14522);
or UO_743 (O_743,N_14691,N_14928);
and UO_744 (O_744,N_14362,N_14805);
or UO_745 (O_745,N_14983,N_14620);
or UO_746 (O_746,N_14454,N_14402);
and UO_747 (O_747,N_14285,N_14942);
and UO_748 (O_748,N_14915,N_14381);
nor UO_749 (O_749,N_14992,N_14712);
nand UO_750 (O_750,N_14767,N_14275);
nand UO_751 (O_751,N_14859,N_14877);
or UO_752 (O_752,N_14470,N_14913);
nor UO_753 (O_753,N_14669,N_14398);
nor UO_754 (O_754,N_14349,N_14263);
or UO_755 (O_755,N_14915,N_14801);
nand UO_756 (O_756,N_14439,N_14805);
or UO_757 (O_757,N_14621,N_14868);
or UO_758 (O_758,N_14547,N_14781);
nor UO_759 (O_759,N_14657,N_14965);
and UO_760 (O_760,N_14415,N_14998);
nor UO_761 (O_761,N_14586,N_14793);
and UO_762 (O_762,N_14572,N_14595);
nand UO_763 (O_763,N_14421,N_14587);
nand UO_764 (O_764,N_14321,N_14831);
nand UO_765 (O_765,N_14708,N_14705);
nand UO_766 (O_766,N_14531,N_14803);
or UO_767 (O_767,N_14487,N_14432);
nor UO_768 (O_768,N_14863,N_14690);
or UO_769 (O_769,N_14438,N_14981);
or UO_770 (O_770,N_14696,N_14677);
nand UO_771 (O_771,N_14322,N_14473);
and UO_772 (O_772,N_14833,N_14464);
xor UO_773 (O_773,N_14822,N_14694);
and UO_774 (O_774,N_14671,N_14454);
or UO_775 (O_775,N_14696,N_14803);
nor UO_776 (O_776,N_14585,N_14315);
xnor UO_777 (O_777,N_14729,N_14289);
nand UO_778 (O_778,N_14583,N_14700);
and UO_779 (O_779,N_14868,N_14305);
or UO_780 (O_780,N_14849,N_14798);
and UO_781 (O_781,N_14309,N_14812);
or UO_782 (O_782,N_14933,N_14472);
or UO_783 (O_783,N_14387,N_14372);
nand UO_784 (O_784,N_14422,N_14746);
nor UO_785 (O_785,N_14704,N_14689);
nand UO_786 (O_786,N_14496,N_14430);
or UO_787 (O_787,N_14392,N_14428);
and UO_788 (O_788,N_14554,N_14370);
nor UO_789 (O_789,N_14757,N_14946);
or UO_790 (O_790,N_14862,N_14438);
nor UO_791 (O_791,N_14271,N_14679);
and UO_792 (O_792,N_14395,N_14491);
nand UO_793 (O_793,N_14567,N_14776);
nor UO_794 (O_794,N_14638,N_14969);
or UO_795 (O_795,N_14968,N_14657);
nor UO_796 (O_796,N_14329,N_14517);
or UO_797 (O_797,N_14905,N_14977);
or UO_798 (O_798,N_14331,N_14439);
or UO_799 (O_799,N_14653,N_14952);
and UO_800 (O_800,N_14979,N_14403);
and UO_801 (O_801,N_14996,N_14607);
and UO_802 (O_802,N_14675,N_14377);
or UO_803 (O_803,N_14623,N_14573);
and UO_804 (O_804,N_14629,N_14944);
nand UO_805 (O_805,N_14621,N_14654);
or UO_806 (O_806,N_14388,N_14552);
and UO_807 (O_807,N_14333,N_14989);
nor UO_808 (O_808,N_14824,N_14754);
nand UO_809 (O_809,N_14410,N_14524);
nor UO_810 (O_810,N_14452,N_14638);
or UO_811 (O_811,N_14975,N_14616);
nand UO_812 (O_812,N_14552,N_14532);
and UO_813 (O_813,N_14505,N_14597);
nand UO_814 (O_814,N_14280,N_14262);
nor UO_815 (O_815,N_14936,N_14418);
or UO_816 (O_816,N_14721,N_14679);
and UO_817 (O_817,N_14397,N_14371);
and UO_818 (O_818,N_14830,N_14286);
nor UO_819 (O_819,N_14645,N_14376);
or UO_820 (O_820,N_14816,N_14755);
and UO_821 (O_821,N_14448,N_14667);
nor UO_822 (O_822,N_14627,N_14809);
nor UO_823 (O_823,N_14554,N_14550);
nor UO_824 (O_824,N_14953,N_14688);
nand UO_825 (O_825,N_14731,N_14589);
or UO_826 (O_826,N_14772,N_14919);
and UO_827 (O_827,N_14819,N_14350);
nand UO_828 (O_828,N_14705,N_14487);
and UO_829 (O_829,N_14487,N_14607);
nand UO_830 (O_830,N_14800,N_14389);
nor UO_831 (O_831,N_14933,N_14794);
nand UO_832 (O_832,N_14497,N_14395);
and UO_833 (O_833,N_14626,N_14837);
nor UO_834 (O_834,N_14970,N_14336);
nand UO_835 (O_835,N_14606,N_14574);
nand UO_836 (O_836,N_14831,N_14599);
or UO_837 (O_837,N_14840,N_14699);
and UO_838 (O_838,N_14704,N_14959);
or UO_839 (O_839,N_14465,N_14750);
nand UO_840 (O_840,N_14360,N_14751);
or UO_841 (O_841,N_14892,N_14872);
or UO_842 (O_842,N_14495,N_14599);
nand UO_843 (O_843,N_14756,N_14940);
xnor UO_844 (O_844,N_14670,N_14904);
and UO_845 (O_845,N_14777,N_14307);
xnor UO_846 (O_846,N_14610,N_14853);
nor UO_847 (O_847,N_14295,N_14347);
or UO_848 (O_848,N_14801,N_14572);
and UO_849 (O_849,N_14705,N_14449);
or UO_850 (O_850,N_14837,N_14912);
xnor UO_851 (O_851,N_14500,N_14806);
or UO_852 (O_852,N_14660,N_14781);
and UO_853 (O_853,N_14321,N_14250);
nor UO_854 (O_854,N_14476,N_14849);
or UO_855 (O_855,N_14715,N_14256);
nand UO_856 (O_856,N_14305,N_14272);
and UO_857 (O_857,N_14632,N_14680);
nor UO_858 (O_858,N_14382,N_14685);
or UO_859 (O_859,N_14506,N_14758);
or UO_860 (O_860,N_14259,N_14331);
and UO_861 (O_861,N_14846,N_14744);
or UO_862 (O_862,N_14902,N_14752);
nor UO_863 (O_863,N_14323,N_14677);
nand UO_864 (O_864,N_14701,N_14912);
nand UO_865 (O_865,N_14527,N_14892);
nand UO_866 (O_866,N_14324,N_14861);
nand UO_867 (O_867,N_14428,N_14945);
nor UO_868 (O_868,N_14794,N_14752);
and UO_869 (O_869,N_14513,N_14895);
and UO_870 (O_870,N_14615,N_14984);
nor UO_871 (O_871,N_14474,N_14453);
or UO_872 (O_872,N_14438,N_14759);
or UO_873 (O_873,N_14250,N_14500);
nor UO_874 (O_874,N_14292,N_14545);
and UO_875 (O_875,N_14508,N_14427);
nand UO_876 (O_876,N_14306,N_14478);
xor UO_877 (O_877,N_14668,N_14262);
nand UO_878 (O_878,N_14820,N_14940);
nand UO_879 (O_879,N_14834,N_14563);
xor UO_880 (O_880,N_14730,N_14756);
nand UO_881 (O_881,N_14982,N_14444);
and UO_882 (O_882,N_14391,N_14949);
and UO_883 (O_883,N_14581,N_14957);
or UO_884 (O_884,N_14595,N_14995);
and UO_885 (O_885,N_14924,N_14272);
or UO_886 (O_886,N_14328,N_14966);
and UO_887 (O_887,N_14611,N_14810);
nor UO_888 (O_888,N_14496,N_14735);
nor UO_889 (O_889,N_14295,N_14378);
and UO_890 (O_890,N_14707,N_14445);
or UO_891 (O_891,N_14432,N_14435);
and UO_892 (O_892,N_14490,N_14882);
nand UO_893 (O_893,N_14639,N_14859);
and UO_894 (O_894,N_14834,N_14466);
nor UO_895 (O_895,N_14714,N_14411);
nand UO_896 (O_896,N_14337,N_14365);
or UO_897 (O_897,N_14677,N_14830);
nor UO_898 (O_898,N_14566,N_14659);
and UO_899 (O_899,N_14524,N_14610);
nor UO_900 (O_900,N_14336,N_14922);
nand UO_901 (O_901,N_14585,N_14276);
nand UO_902 (O_902,N_14590,N_14573);
or UO_903 (O_903,N_14628,N_14851);
xor UO_904 (O_904,N_14661,N_14358);
nand UO_905 (O_905,N_14563,N_14754);
nand UO_906 (O_906,N_14516,N_14302);
and UO_907 (O_907,N_14615,N_14437);
or UO_908 (O_908,N_14603,N_14402);
nand UO_909 (O_909,N_14836,N_14998);
nor UO_910 (O_910,N_14656,N_14868);
nor UO_911 (O_911,N_14895,N_14558);
nor UO_912 (O_912,N_14385,N_14508);
nor UO_913 (O_913,N_14665,N_14386);
and UO_914 (O_914,N_14294,N_14829);
or UO_915 (O_915,N_14995,N_14310);
and UO_916 (O_916,N_14431,N_14789);
or UO_917 (O_917,N_14879,N_14823);
nor UO_918 (O_918,N_14739,N_14802);
nand UO_919 (O_919,N_14833,N_14367);
and UO_920 (O_920,N_14760,N_14331);
nor UO_921 (O_921,N_14867,N_14860);
nand UO_922 (O_922,N_14334,N_14923);
and UO_923 (O_923,N_14287,N_14790);
and UO_924 (O_924,N_14321,N_14952);
nand UO_925 (O_925,N_14395,N_14768);
nand UO_926 (O_926,N_14827,N_14368);
and UO_927 (O_927,N_14328,N_14389);
and UO_928 (O_928,N_14674,N_14586);
nand UO_929 (O_929,N_14459,N_14291);
and UO_930 (O_930,N_14731,N_14758);
nand UO_931 (O_931,N_14787,N_14814);
nor UO_932 (O_932,N_14950,N_14680);
and UO_933 (O_933,N_14301,N_14360);
nand UO_934 (O_934,N_14528,N_14775);
xnor UO_935 (O_935,N_14704,N_14491);
nor UO_936 (O_936,N_14628,N_14900);
nor UO_937 (O_937,N_14665,N_14427);
nand UO_938 (O_938,N_14539,N_14698);
and UO_939 (O_939,N_14273,N_14743);
nand UO_940 (O_940,N_14336,N_14363);
nor UO_941 (O_941,N_14603,N_14955);
nor UO_942 (O_942,N_14597,N_14760);
and UO_943 (O_943,N_14497,N_14498);
nand UO_944 (O_944,N_14288,N_14398);
and UO_945 (O_945,N_14555,N_14349);
and UO_946 (O_946,N_14729,N_14662);
or UO_947 (O_947,N_14283,N_14279);
nor UO_948 (O_948,N_14984,N_14551);
or UO_949 (O_949,N_14726,N_14800);
nor UO_950 (O_950,N_14271,N_14866);
nand UO_951 (O_951,N_14773,N_14546);
nor UO_952 (O_952,N_14454,N_14783);
nor UO_953 (O_953,N_14449,N_14568);
nand UO_954 (O_954,N_14477,N_14911);
nor UO_955 (O_955,N_14906,N_14314);
nand UO_956 (O_956,N_14668,N_14317);
or UO_957 (O_957,N_14259,N_14856);
or UO_958 (O_958,N_14481,N_14550);
nor UO_959 (O_959,N_14758,N_14722);
nor UO_960 (O_960,N_14837,N_14573);
and UO_961 (O_961,N_14668,N_14602);
nor UO_962 (O_962,N_14422,N_14774);
or UO_963 (O_963,N_14424,N_14359);
nor UO_964 (O_964,N_14622,N_14276);
nor UO_965 (O_965,N_14393,N_14441);
nand UO_966 (O_966,N_14528,N_14932);
nor UO_967 (O_967,N_14623,N_14795);
nor UO_968 (O_968,N_14838,N_14571);
or UO_969 (O_969,N_14882,N_14896);
or UO_970 (O_970,N_14532,N_14255);
nand UO_971 (O_971,N_14266,N_14420);
and UO_972 (O_972,N_14864,N_14780);
or UO_973 (O_973,N_14528,N_14736);
and UO_974 (O_974,N_14456,N_14540);
xor UO_975 (O_975,N_14921,N_14475);
nand UO_976 (O_976,N_14943,N_14619);
or UO_977 (O_977,N_14578,N_14765);
nor UO_978 (O_978,N_14799,N_14856);
xor UO_979 (O_979,N_14511,N_14566);
nor UO_980 (O_980,N_14741,N_14561);
nand UO_981 (O_981,N_14594,N_14767);
and UO_982 (O_982,N_14552,N_14310);
nand UO_983 (O_983,N_14278,N_14517);
or UO_984 (O_984,N_14838,N_14617);
and UO_985 (O_985,N_14956,N_14827);
or UO_986 (O_986,N_14517,N_14445);
nand UO_987 (O_987,N_14977,N_14297);
nand UO_988 (O_988,N_14515,N_14853);
or UO_989 (O_989,N_14426,N_14309);
or UO_990 (O_990,N_14297,N_14414);
nand UO_991 (O_991,N_14588,N_14268);
nand UO_992 (O_992,N_14747,N_14353);
nor UO_993 (O_993,N_14908,N_14757);
or UO_994 (O_994,N_14511,N_14714);
nand UO_995 (O_995,N_14917,N_14428);
and UO_996 (O_996,N_14513,N_14538);
nand UO_997 (O_997,N_14779,N_14751);
nor UO_998 (O_998,N_14936,N_14781);
and UO_999 (O_999,N_14993,N_14538);
nand UO_1000 (O_1000,N_14991,N_14580);
and UO_1001 (O_1001,N_14661,N_14260);
nand UO_1002 (O_1002,N_14699,N_14338);
nand UO_1003 (O_1003,N_14439,N_14641);
nand UO_1004 (O_1004,N_14526,N_14855);
nor UO_1005 (O_1005,N_14880,N_14311);
and UO_1006 (O_1006,N_14933,N_14427);
or UO_1007 (O_1007,N_14502,N_14681);
and UO_1008 (O_1008,N_14379,N_14787);
nor UO_1009 (O_1009,N_14974,N_14628);
and UO_1010 (O_1010,N_14428,N_14482);
nand UO_1011 (O_1011,N_14762,N_14593);
nand UO_1012 (O_1012,N_14603,N_14838);
nand UO_1013 (O_1013,N_14577,N_14760);
nor UO_1014 (O_1014,N_14958,N_14582);
and UO_1015 (O_1015,N_14555,N_14326);
nor UO_1016 (O_1016,N_14910,N_14325);
or UO_1017 (O_1017,N_14263,N_14720);
nand UO_1018 (O_1018,N_14329,N_14582);
nor UO_1019 (O_1019,N_14472,N_14732);
nand UO_1020 (O_1020,N_14709,N_14379);
or UO_1021 (O_1021,N_14438,N_14368);
and UO_1022 (O_1022,N_14594,N_14826);
nor UO_1023 (O_1023,N_14768,N_14259);
and UO_1024 (O_1024,N_14262,N_14857);
nand UO_1025 (O_1025,N_14611,N_14494);
or UO_1026 (O_1026,N_14945,N_14715);
and UO_1027 (O_1027,N_14620,N_14602);
nand UO_1028 (O_1028,N_14493,N_14412);
or UO_1029 (O_1029,N_14823,N_14710);
nor UO_1030 (O_1030,N_14624,N_14899);
nand UO_1031 (O_1031,N_14654,N_14613);
nand UO_1032 (O_1032,N_14919,N_14805);
or UO_1033 (O_1033,N_14496,N_14684);
or UO_1034 (O_1034,N_14695,N_14399);
nor UO_1035 (O_1035,N_14806,N_14663);
nand UO_1036 (O_1036,N_14796,N_14383);
nor UO_1037 (O_1037,N_14686,N_14765);
nor UO_1038 (O_1038,N_14631,N_14640);
nand UO_1039 (O_1039,N_14547,N_14409);
nor UO_1040 (O_1040,N_14376,N_14816);
or UO_1041 (O_1041,N_14319,N_14296);
nand UO_1042 (O_1042,N_14493,N_14979);
nand UO_1043 (O_1043,N_14669,N_14337);
and UO_1044 (O_1044,N_14655,N_14408);
nand UO_1045 (O_1045,N_14340,N_14471);
nor UO_1046 (O_1046,N_14372,N_14814);
and UO_1047 (O_1047,N_14946,N_14267);
and UO_1048 (O_1048,N_14414,N_14351);
nand UO_1049 (O_1049,N_14984,N_14828);
or UO_1050 (O_1050,N_14659,N_14269);
nand UO_1051 (O_1051,N_14809,N_14718);
or UO_1052 (O_1052,N_14789,N_14864);
and UO_1053 (O_1053,N_14725,N_14970);
and UO_1054 (O_1054,N_14544,N_14730);
nor UO_1055 (O_1055,N_14892,N_14713);
nor UO_1056 (O_1056,N_14724,N_14665);
nor UO_1057 (O_1057,N_14705,N_14776);
and UO_1058 (O_1058,N_14471,N_14476);
nor UO_1059 (O_1059,N_14312,N_14976);
or UO_1060 (O_1060,N_14578,N_14764);
nor UO_1061 (O_1061,N_14820,N_14931);
and UO_1062 (O_1062,N_14605,N_14585);
nand UO_1063 (O_1063,N_14554,N_14945);
nand UO_1064 (O_1064,N_14520,N_14361);
nor UO_1065 (O_1065,N_14447,N_14941);
and UO_1066 (O_1066,N_14460,N_14939);
nand UO_1067 (O_1067,N_14805,N_14303);
nor UO_1068 (O_1068,N_14874,N_14767);
or UO_1069 (O_1069,N_14375,N_14503);
or UO_1070 (O_1070,N_14657,N_14954);
and UO_1071 (O_1071,N_14871,N_14418);
or UO_1072 (O_1072,N_14330,N_14868);
and UO_1073 (O_1073,N_14740,N_14963);
and UO_1074 (O_1074,N_14276,N_14464);
or UO_1075 (O_1075,N_14400,N_14998);
or UO_1076 (O_1076,N_14272,N_14735);
or UO_1077 (O_1077,N_14735,N_14358);
or UO_1078 (O_1078,N_14409,N_14371);
nand UO_1079 (O_1079,N_14740,N_14741);
and UO_1080 (O_1080,N_14333,N_14824);
nor UO_1081 (O_1081,N_14463,N_14737);
or UO_1082 (O_1082,N_14874,N_14541);
and UO_1083 (O_1083,N_14826,N_14683);
or UO_1084 (O_1084,N_14959,N_14841);
and UO_1085 (O_1085,N_14800,N_14893);
and UO_1086 (O_1086,N_14990,N_14457);
or UO_1087 (O_1087,N_14900,N_14921);
and UO_1088 (O_1088,N_14419,N_14890);
nor UO_1089 (O_1089,N_14775,N_14967);
and UO_1090 (O_1090,N_14553,N_14518);
nand UO_1091 (O_1091,N_14262,N_14484);
or UO_1092 (O_1092,N_14765,N_14853);
or UO_1093 (O_1093,N_14980,N_14964);
and UO_1094 (O_1094,N_14328,N_14533);
nor UO_1095 (O_1095,N_14927,N_14461);
nor UO_1096 (O_1096,N_14390,N_14594);
nand UO_1097 (O_1097,N_14820,N_14324);
and UO_1098 (O_1098,N_14603,N_14431);
nor UO_1099 (O_1099,N_14842,N_14836);
and UO_1100 (O_1100,N_14878,N_14554);
and UO_1101 (O_1101,N_14747,N_14660);
nand UO_1102 (O_1102,N_14439,N_14840);
nor UO_1103 (O_1103,N_14789,N_14368);
nand UO_1104 (O_1104,N_14397,N_14950);
nor UO_1105 (O_1105,N_14894,N_14432);
nor UO_1106 (O_1106,N_14508,N_14340);
and UO_1107 (O_1107,N_14289,N_14898);
or UO_1108 (O_1108,N_14480,N_14757);
and UO_1109 (O_1109,N_14669,N_14379);
and UO_1110 (O_1110,N_14542,N_14867);
nand UO_1111 (O_1111,N_14851,N_14332);
or UO_1112 (O_1112,N_14589,N_14509);
or UO_1113 (O_1113,N_14822,N_14902);
nor UO_1114 (O_1114,N_14627,N_14344);
nand UO_1115 (O_1115,N_14450,N_14594);
or UO_1116 (O_1116,N_14870,N_14609);
and UO_1117 (O_1117,N_14821,N_14911);
nor UO_1118 (O_1118,N_14684,N_14685);
nand UO_1119 (O_1119,N_14850,N_14319);
nand UO_1120 (O_1120,N_14763,N_14863);
and UO_1121 (O_1121,N_14729,N_14908);
nand UO_1122 (O_1122,N_14812,N_14274);
or UO_1123 (O_1123,N_14614,N_14625);
nand UO_1124 (O_1124,N_14528,N_14843);
nand UO_1125 (O_1125,N_14489,N_14457);
and UO_1126 (O_1126,N_14649,N_14548);
nor UO_1127 (O_1127,N_14912,N_14765);
and UO_1128 (O_1128,N_14509,N_14768);
or UO_1129 (O_1129,N_14406,N_14903);
nand UO_1130 (O_1130,N_14442,N_14406);
and UO_1131 (O_1131,N_14525,N_14604);
nor UO_1132 (O_1132,N_14654,N_14909);
or UO_1133 (O_1133,N_14862,N_14387);
or UO_1134 (O_1134,N_14492,N_14419);
nor UO_1135 (O_1135,N_14328,N_14473);
nand UO_1136 (O_1136,N_14979,N_14953);
nor UO_1137 (O_1137,N_14974,N_14650);
nand UO_1138 (O_1138,N_14857,N_14651);
or UO_1139 (O_1139,N_14361,N_14772);
or UO_1140 (O_1140,N_14420,N_14934);
and UO_1141 (O_1141,N_14818,N_14357);
nand UO_1142 (O_1142,N_14808,N_14777);
and UO_1143 (O_1143,N_14895,N_14556);
nor UO_1144 (O_1144,N_14839,N_14673);
nand UO_1145 (O_1145,N_14650,N_14994);
nand UO_1146 (O_1146,N_14450,N_14906);
or UO_1147 (O_1147,N_14749,N_14768);
nor UO_1148 (O_1148,N_14826,N_14483);
nand UO_1149 (O_1149,N_14592,N_14961);
or UO_1150 (O_1150,N_14270,N_14286);
nor UO_1151 (O_1151,N_14644,N_14871);
or UO_1152 (O_1152,N_14822,N_14670);
and UO_1153 (O_1153,N_14924,N_14253);
nand UO_1154 (O_1154,N_14855,N_14869);
nand UO_1155 (O_1155,N_14408,N_14425);
xnor UO_1156 (O_1156,N_14942,N_14939);
or UO_1157 (O_1157,N_14630,N_14909);
nand UO_1158 (O_1158,N_14251,N_14444);
or UO_1159 (O_1159,N_14535,N_14483);
nor UO_1160 (O_1160,N_14688,N_14372);
xnor UO_1161 (O_1161,N_14461,N_14960);
and UO_1162 (O_1162,N_14373,N_14342);
and UO_1163 (O_1163,N_14393,N_14339);
nor UO_1164 (O_1164,N_14849,N_14559);
and UO_1165 (O_1165,N_14269,N_14530);
nor UO_1166 (O_1166,N_14887,N_14779);
or UO_1167 (O_1167,N_14992,N_14778);
or UO_1168 (O_1168,N_14373,N_14487);
and UO_1169 (O_1169,N_14533,N_14275);
nand UO_1170 (O_1170,N_14361,N_14348);
nand UO_1171 (O_1171,N_14308,N_14955);
nor UO_1172 (O_1172,N_14750,N_14758);
nand UO_1173 (O_1173,N_14349,N_14863);
nand UO_1174 (O_1174,N_14670,N_14693);
nand UO_1175 (O_1175,N_14604,N_14575);
nand UO_1176 (O_1176,N_14780,N_14373);
nand UO_1177 (O_1177,N_14740,N_14593);
nor UO_1178 (O_1178,N_14317,N_14413);
nand UO_1179 (O_1179,N_14930,N_14642);
nand UO_1180 (O_1180,N_14746,N_14740);
and UO_1181 (O_1181,N_14502,N_14584);
and UO_1182 (O_1182,N_14333,N_14560);
or UO_1183 (O_1183,N_14966,N_14774);
nand UO_1184 (O_1184,N_14251,N_14729);
and UO_1185 (O_1185,N_14988,N_14810);
and UO_1186 (O_1186,N_14745,N_14484);
and UO_1187 (O_1187,N_14557,N_14662);
nand UO_1188 (O_1188,N_14975,N_14510);
nor UO_1189 (O_1189,N_14576,N_14375);
and UO_1190 (O_1190,N_14978,N_14985);
or UO_1191 (O_1191,N_14468,N_14620);
nor UO_1192 (O_1192,N_14834,N_14428);
or UO_1193 (O_1193,N_14418,N_14381);
nand UO_1194 (O_1194,N_14732,N_14573);
and UO_1195 (O_1195,N_14829,N_14783);
nor UO_1196 (O_1196,N_14770,N_14350);
or UO_1197 (O_1197,N_14561,N_14883);
nor UO_1198 (O_1198,N_14633,N_14603);
nand UO_1199 (O_1199,N_14372,N_14490);
and UO_1200 (O_1200,N_14378,N_14558);
or UO_1201 (O_1201,N_14506,N_14967);
nand UO_1202 (O_1202,N_14547,N_14707);
or UO_1203 (O_1203,N_14616,N_14561);
and UO_1204 (O_1204,N_14963,N_14924);
nor UO_1205 (O_1205,N_14282,N_14351);
or UO_1206 (O_1206,N_14953,N_14422);
nand UO_1207 (O_1207,N_14701,N_14371);
and UO_1208 (O_1208,N_14631,N_14856);
nand UO_1209 (O_1209,N_14504,N_14785);
and UO_1210 (O_1210,N_14775,N_14961);
nand UO_1211 (O_1211,N_14531,N_14599);
or UO_1212 (O_1212,N_14685,N_14492);
xnor UO_1213 (O_1213,N_14988,N_14801);
and UO_1214 (O_1214,N_14910,N_14424);
nor UO_1215 (O_1215,N_14701,N_14659);
nor UO_1216 (O_1216,N_14905,N_14737);
or UO_1217 (O_1217,N_14355,N_14464);
nor UO_1218 (O_1218,N_14388,N_14608);
nor UO_1219 (O_1219,N_14656,N_14314);
or UO_1220 (O_1220,N_14278,N_14570);
and UO_1221 (O_1221,N_14494,N_14878);
or UO_1222 (O_1222,N_14513,N_14541);
nor UO_1223 (O_1223,N_14569,N_14321);
nor UO_1224 (O_1224,N_14749,N_14960);
nor UO_1225 (O_1225,N_14974,N_14630);
and UO_1226 (O_1226,N_14846,N_14617);
or UO_1227 (O_1227,N_14691,N_14523);
nand UO_1228 (O_1228,N_14932,N_14752);
nor UO_1229 (O_1229,N_14711,N_14910);
or UO_1230 (O_1230,N_14562,N_14776);
nand UO_1231 (O_1231,N_14357,N_14698);
nand UO_1232 (O_1232,N_14859,N_14615);
and UO_1233 (O_1233,N_14258,N_14594);
nand UO_1234 (O_1234,N_14286,N_14698);
and UO_1235 (O_1235,N_14620,N_14357);
nor UO_1236 (O_1236,N_14942,N_14316);
and UO_1237 (O_1237,N_14323,N_14722);
nand UO_1238 (O_1238,N_14770,N_14340);
or UO_1239 (O_1239,N_14997,N_14708);
xor UO_1240 (O_1240,N_14801,N_14588);
and UO_1241 (O_1241,N_14957,N_14567);
nand UO_1242 (O_1242,N_14621,N_14451);
nor UO_1243 (O_1243,N_14581,N_14873);
or UO_1244 (O_1244,N_14343,N_14720);
and UO_1245 (O_1245,N_14380,N_14537);
nor UO_1246 (O_1246,N_14463,N_14623);
nand UO_1247 (O_1247,N_14940,N_14932);
and UO_1248 (O_1248,N_14924,N_14582);
nand UO_1249 (O_1249,N_14526,N_14743);
or UO_1250 (O_1250,N_14502,N_14921);
and UO_1251 (O_1251,N_14422,N_14567);
nand UO_1252 (O_1252,N_14369,N_14898);
nor UO_1253 (O_1253,N_14574,N_14429);
and UO_1254 (O_1254,N_14740,N_14250);
and UO_1255 (O_1255,N_14462,N_14831);
or UO_1256 (O_1256,N_14722,N_14525);
and UO_1257 (O_1257,N_14853,N_14881);
and UO_1258 (O_1258,N_14733,N_14664);
nand UO_1259 (O_1259,N_14855,N_14387);
or UO_1260 (O_1260,N_14429,N_14342);
and UO_1261 (O_1261,N_14975,N_14739);
or UO_1262 (O_1262,N_14288,N_14763);
or UO_1263 (O_1263,N_14479,N_14733);
nor UO_1264 (O_1264,N_14998,N_14722);
or UO_1265 (O_1265,N_14802,N_14454);
xor UO_1266 (O_1266,N_14415,N_14682);
nand UO_1267 (O_1267,N_14623,N_14625);
nor UO_1268 (O_1268,N_14488,N_14991);
or UO_1269 (O_1269,N_14743,N_14795);
and UO_1270 (O_1270,N_14579,N_14305);
nor UO_1271 (O_1271,N_14847,N_14870);
nand UO_1272 (O_1272,N_14694,N_14644);
xor UO_1273 (O_1273,N_14648,N_14804);
or UO_1274 (O_1274,N_14881,N_14327);
xnor UO_1275 (O_1275,N_14368,N_14718);
nand UO_1276 (O_1276,N_14423,N_14923);
or UO_1277 (O_1277,N_14945,N_14953);
nand UO_1278 (O_1278,N_14875,N_14570);
nand UO_1279 (O_1279,N_14825,N_14450);
nand UO_1280 (O_1280,N_14963,N_14368);
nor UO_1281 (O_1281,N_14292,N_14326);
nor UO_1282 (O_1282,N_14880,N_14363);
and UO_1283 (O_1283,N_14949,N_14833);
or UO_1284 (O_1284,N_14781,N_14885);
or UO_1285 (O_1285,N_14566,N_14536);
and UO_1286 (O_1286,N_14909,N_14475);
nor UO_1287 (O_1287,N_14371,N_14394);
and UO_1288 (O_1288,N_14836,N_14476);
nand UO_1289 (O_1289,N_14270,N_14770);
nand UO_1290 (O_1290,N_14840,N_14304);
nand UO_1291 (O_1291,N_14957,N_14326);
nor UO_1292 (O_1292,N_14416,N_14441);
or UO_1293 (O_1293,N_14748,N_14263);
or UO_1294 (O_1294,N_14315,N_14277);
nand UO_1295 (O_1295,N_14684,N_14794);
and UO_1296 (O_1296,N_14623,N_14745);
or UO_1297 (O_1297,N_14988,N_14261);
or UO_1298 (O_1298,N_14784,N_14624);
nand UO_1299 (O_1299,N_14383,N_14603);
nand UO_1300 (O_1300,N_14683,N_14946);
nand UO_1301 (O_1301,N_14788,N_14908);
nor UO_1302 (O_1302,N_14360,N_14550);
nand UO_1303 (O_1303,N_14908,N_14968);
nand UO_1304 (O_1304,N_14523,N_14345);
nand UO_1305 (O_1305,N_14942,N_14752);
xnor UO_1306 (O_1306,N_14463,N_14524);
nand UO_1307 (O_1307,N_14761,N_14620);
and UO_1308 (O_1308,N_14463,N_14279);
nor UO_1309 (O_1309,N_14677,N_14518);
nand UO_1310 (O_1310,N_14731,N_14307);
and UO_1311 (O_1311,N_14663,N_14863);
nor UO_1312 (O_1312,N_14918,N_14981);
or UO_1313 (O_1313,N_14266,N_14401);
nand UO_1314 (O_1314,N_14476,N_14652);
nand UO_1315 (O_1315,N_14700,N_14434);
and UO_1316 (O_1316,N_14788,N_14653);
nor UO_1317 (O_1317,N_14854,N_14690);
nand UO_1318 (O_1318,N_14292,N_14818);
and UO_1319 (O_1319,N_14936,N_14286);
nand UO_1320 (O_1320,N_14908,N_14474);
nor UO_1321 (O_1321,N_14339,N_14326);
nand UO_1322 (O_1322,N_14471,N_14263);
nand UO_1323 (O_1323,N_14993,N_14348);
nor UO_1324 (O_1324,N_14732,N_14586);
nand UO_1325 (O_1325,N_14573,N_14796);
or UO_1326 (O_1326,N_14819,N_14622);
and UO_1327 (O_1327,N_14315,N_14917);
nand UO_1328 (O_1328,N_14771,N_14806);
nor UO_1329 (O_1329,N_14734,N_14365);
or UO_1330 (O_1330,N_14695,N_14722);
and UO_1331 (O_1331,N_14706,N_14453);
or UO_1332 (O_1332,N_14424,N_14445);
and UO_1333 (O_1333,N_14902,N_14681);
nand UO_1334 (O_1334,N_14356,N_14617);
nand UO_1335 (O_1335,N_14541,N_14621);
or UO_1336 (O_1336,N_14680,N_14433);
or UO_1337 (O_1337,N_14399,N_14488);
or UO_1338 (O_1338,N_14925,N_14277);
or UO_1339 (O_1339,N_14315,N_14345);
nand UO_1340 (O_1340,N_14568,N_14741);
nor UO_1341 (O_1341,N_14299,N_14917);
nand UO_1342 (O_1342,N_14789,N_14514);
and UO_1343 (O_1343,N_14859,N_14871);
nor UO_1344 (O_1344,N_14381,N_14400);
or UO_1345 (O_1345,N_14436,N_14913);
nand UO_1346 (O_1346,N_14395,N_14945);
nand UO_1347 (O_1347,N_14925,N_14432);
nand UO_1348 (O_1348,N_14761,N_14303);
and UO_1349 (O_1349,N_14613,N_14354);
nand UO_1350 (O_1350,N_14758,N_14416);
or UO_1351 (O_1351,N_14715,N_14602);
nand UO_1352 (O_1352,N_14493,N_14837);
nand UO_1353 (O_1353,N_14598,N_14323);
nand UO_1354 (O_1354,N_14299,N_14923);
nand UO_1355 (O_1355,N_14508,N_14313);
or UO_1356 (O_1356,N_14564,N_14787);
or UO_1357 (O_1357,N_14501,N_14635);
nand UO_1358 (O_1358,N_14780,N_14614);
or UO_1359 (O_1359,N_14455,N_14800);
and UO_1360 (O_1360,N_14576,N_14626);
nand UO_1361 (O_1361,N_14975,N_14995);
and UO_1362 (O_1362,N_14462,N_14397);
nor UO_1363 (O_1363,N_14968,N_14323);
nor UO_1364 (O_1364,N_14749,N_14894);
nor UO_1365 (O_1365,N_14388,N_14544);
nor UO_1366 (O_1366,N_14642,N_14594);
nor UO_1367 (O_1367,N_14578,N_14833);
nand UO_1368 (O_1368,N_14707,N_14526);
and UO_1369 (O_1369,N_14466,N_14360);
or UO_1370 (O_1370,N_14875,N_14776);
or UO_1371 (O_1371,N_14580,N_14287);
and UO_1372 (O_1372,N_14668,N_14664);
or UO_1373 (O_1373,N_14381,N_14679);
nand UO_1374 (O_1374,N_14680,N_14986);
and UO_1375 (O_1375,N_14350,N_14883);
and UO_1376 (O_1376,N_14548,N_14956);
or UO_1377 (O_1377,N_14687,N_14279);
or UO_1378 (O_1378,N_14672,N_14589);
nand UO_1379 (O_1379,N_14611,N_14889);
or UO_1380 (O_1380,N_14842,N_14263);
or UO_1381 (O_1381,N_14712,N_14401);
and UO_1382 (O_1382,N_14833,N_14820);
or UO_1383 (O_1383,N_14530,N_14668);
nand UO_1384 (O_1384,N_14408,N_14514);
nand UO_1385 (O_1385,N_14414,N_14876);
nor UO_1386 (O_1386,N_14890,N_14718);
and UO_1387 (O_1387,N_14523,N_14812);
nor UO_1388 (O_1388,N_14991,N_14640);
nor UO_1389 (O_1389,N_14697,N_14917);
nand UO_1390 (O_1390,N_14894,N_14447);
or UO_1391 (O_1391,N_14366,N_14574);
nand UO_1392 (O_1392,N_14982,N_14683);
nand UO_1393 (O_1393,N_14699,N_14277);
and UO_1394 (O_1394,N_14342,N_14812);
or UO_1395 (O_1395,N_14673,N_14682);
and UO_1396 (O_1396,N_14665,N_14547);
or UO_1397 (O_1397,N_14579,N_14768);
nand UO_1398 (O_1398,N_14383,N_14860);
nor UO_1399 (O_1399,N_14813,N_14289);
or UO_1400 (O_1400,N_14727,N_14474);
nand UO_1401 (O_1401,N_14517,N_14954);
xnor UO_1402 (O_1402,N_14357,N_14828);
nand UO_1403 (O_1403,N_14621,N_14990);
or UO_1404 (O_1404,N_14792,N_14617);
or UO_1405 (O_1405,N_14258,N_14981);
nor UO_1406 (O_1406,N_14689,N_14901);
nor UO_1407 (O_1407,N_14871,N_14659);
or UO_1408 (O_1408,N_14578,N_14277);
nand UO_1409 (O_1409,N_14580,N_14409);
nor UO_1410 (O_1410,N_14549,N_14318);
nor UO_1411 (O_1411,N_14780,N_14435);
nor UO_1412 (O_1412,N_14894,N_14824);
nor UO_1413 (O_1413,N_14777,N_14611);
nor UO_1414 (O_1414,N_14711,N_14480);
nand UO_1415 (O_1415,N_14916,N_14665);
or UO_1416 (O_1416,N_14372,N_14602);
and UO_1417 (O_1417,N_14481,N_14438);
nor UO_1418 (O_1418,N_14406,N_14334);
nor UO_1419 (O_1419,N_14825,N_14509);
nand UO_1420 (O_1420,N_14859,N_14554);
and UO_1421 (O_1421,N_14743,N_14828);
xor UO_1422 (O_1422,N_14297,N_14772);
nor UO_1423 (O_1423,N_14481,N_14279);
nor UO_1424 (O_1424,N_14689,N_14769);
nand UO_1425 (O_1425,N_14875,N_14965);
xnor UO_1426 (O_1426,N_14612,N_14391);
xnor UO_1427 (O_1427,N_14755,N_14711);
nor UO_1428 (O_1428,N_14502,N_14304);
and UO_1429 (O_1429,N_14260,N_14856);
nor UO_1430 (O_1430,N_14864,N_14264);
nand UO_1431 (O_1431,N_14842,N_14488);
xnor UO_1432 (O_1432,N_14986,N_14897);
nand UO_1433 (O_1433,N_14934,N_14316);
nor UO_1434 (O_1434,N_14708,N_14770);
nand UO_1435 (O_1435,N_14326,N_14583);
and UO_1436 (O_1436,N_14323,N_14631);
xor UO_1437 (O_1437,N_14528,N_14910);
nor UO_1438 (O_1438,N_14364,N_14524);
and UO_1439 (O_1439,N_14823,N_14756);
nor UO_1440 (O_1440,N_14944,N_14459);
nand UO_1441 (O_1441,N_14538,N_14556);
and UO_1442 (O_1442,N_14847,N_14813);
nor UO_1443 (O_1443,N_14511,N_14913);
nand UO_1444 (O_1444,N_14328,N_14923);
xnor UO_1445 (O_1445,N_14844,N_14906);
nand UO_1446 (O_1446,N_14824,N_14867);
nor UO_1447 (O_1447,N_14455,N_14798);
nand UO_1448 (O_1448,N_14758,N_14373);
or UO_1449 (O_1449,N_14709,N_14471);
or UO_1450 (O_1450,N_14715,N_14338);
or UO_1451 (O_1451,N_14599,N_14486);
and UO_1452 (O_1452,N_14330,N_14394);
nand UO_1453 (O_1453,N_14398,N_14796);
and UO_1454 (O_1454,N_14315,N_14817);
and UO_1455 (O_1455,N_14536,N_14935);
nand UO_1456 (O_1456,N_14720,N_14957);
nand UO_1457 (O_1457,N_14613,N_14640);
and UO_1458 (O_1458,N_14674,N_14962);
and UO_1459 (O_1459,N_14748,N_14775);
and UO_1460 (O_1460,N_14620,N_14972);
or UO_1461 (O_1461,N_14411,N_14496);
or UO_1462 (O_1462,N_14557,N_14800);
nand UO_1463 (O_1463,N_14414,N_14677);
nor UO_1464 (O_1464,N_14320,N_14838);
and UO_1465 (O_1465,N_14430,N_14837);
nor UO_1466 (O_1466,N_14366,N_14879);
nand UO_1467 (O_1467,N_14956,N_14390);
nor UO_1468 (O_1468,N_14397,N_14986);
nor UO_1469 (O_1469,N_14667,N_14918);
or UO_1470 (O_1470,N_14417,N_14314);
nor UO_1471 (O_1471,N_14493,N_14429);
nand UO_1472 (O_1472,N_14702,N_14870);
nand UO_1473 (O_1473,N_14935,N_14773);
nor UO_1474 (O_1474,N_14512,N_14823);
nor UO_1475 (O_1475,N_14533,N_14773);
nor UO_1476 (O_1476,N_14875,N_14256);
and UO_1477 (O_1477,N_14614,N_14511);
nand UO_1478 (O_1478,N_14711,N_14419);
and UO_1479 (O_1479,N_14932,N_14476);
or UO_1480 (O_1480,N_14309,N_14654);
or UO_1481 (O_1481,N_14507,N_14864);
nor UO_1482 (O_1482,N_14933,N_14309);
and UO_1483 (O_1483,N_14486,N_14806);
nand UO_1484 (O_1484,N_14904,N_14284);
nand UO_1485 (O_1485,N_14355,N_14861);
and UO_1486 (O_1486,N_14425,N_14331);
or UO_1487 (O_1487,N_14861,N_14373);
nand UO_1488 (O_1488,N_14614,N_14909);
nand UO_1489 (O_1489,N_14624,N_14611);
nand UO_1490 (O_1490,N_14881,N_14627);
nand UO_1491 (O_1491,N_14791,N_14865);
and UO_1492 (O_1492,N_14697,N_14402);
nand UO_1493 (O_1493,N_14395,N_14743);
or UO_1494 (O_1494,N_14490,N_14904);
and UO_1495 (O_1495,N_14668,N_14393);
nor UO_1496 (O_1496,N_14715,N_14355);
nor UO_1497 (O_1497,N_14344,N_14894);
or UO_1498 (O_1498,N_14396,N_14686);
or UO_1499 (O_1499,N_14932,N_14766);
and UO_1500 (O_1500,N_14478,N_14941);
and UO_1501 (O_1501,N_14733,N_14619);
nand UO_1502 (O_1502,N_14880,N_14283);
and UO_1503 (O_1503,N_14385,N_14530);
and UO_1504 (O_1504,N_14708,N_14782);
nor UO_1505 (O_1505,N_14326,N_14305);
nand UO_1506 (O_1506,N_14355,N_14432);
or UO_1507 (O_1507,N_14396,N_14661);
xnor UO_1508 (O_1508,N_14754,N_14630);
nor UO_1509 (O_1509,N_14911,N_14654);
or UO_1510 (O_1510,N_14647,N_14810);
and UO_1511 (O_1511,N_14378,N_14562);
xor UO_1512 (O_1512,N_14668,N_14696);
nand UO_1513 (O_1513,N_14872,N_14549);
and UO_1514 (O_1514,N_14820,N_14426);
nor UO_1515 (O_1515,N_14446,N_14367);
nor UO_1516 (O_1516,N_14579,N_14915);
nor UO_1517 (O_1517,N_14349,N_14348);
nand UO_1518 (O_1518,N_14455,N_14769);
nor UO_1519 (O_1519,N_14739,N_14458);
or UO_1520 (O_1520,N_14273,N_14657);
or UO_1521 (O_1521,N_14402,N_14370);
or UO_1522 (O_1522,N_14497,N_14374);
and UO_1523 (O_1523,N_14823,N_14698);
and UO_1524 (O_1524,N_14656,N_14559);
or UO_1525 (O_1525,N_14914,N_14657);
nor UO_1526 (O_1526,N_14254,N_14267);
and UO_1527 (O_1527,N_14637,N_14963);
or UO_1528 (O_1528,N_14893,N_14942);
or UO_1529 (O_1529,N_14652,N_14753);
and UO_1530 (O_1530,N_14394,N_14512);
and UO_1531 (O_1531,N_14343,N_14510);
and UO_1532 (O_1532,N_14370,N_14307);
nand UO_1533 (O_1533,N_14658,N_14400);
or UO_1534 (O_1534,N_14400,N_14631);
nor UO_1535 (O_1535,N_14994,N_14803);
or UO_1536 (O_1536,N_14285,N_14789);
or UO_1537 (O_1537,N_14464,N_14433);
and UO_1538 (O_1538,N_14294,N_14809);
xor UO_1539 (O_1539,N_14982,N_14958);
or UO_1540 (O_1540,N_14696,N_14650);
or UO_1541 (O_1541,N_14927,N_14696);
nand UO_1542 (O_1542,N_14775,N_14374);
and UO_1543 (O_1543,N_14860,N_14812);
and UO_1544 (O_1544,N_14343,N_14881);
nand UO_1545 (O_1545,N_14589,N_14340);
nor UO_1546 (O_1546,N_14332,N_14751);
nor UO_1547 (O_1547,N_14868,N_14419);
or UO_1548 (O_1548,N_14492,N_14280);
or UO_1549 (O_1549,N_14976,N_14632);
and UO_1550 (O_1550,N_14465,N_14334);
and UO_1551 (O_1551,N_14334,N_14905);
or UO_1552 (O_1552,N_14588,N_14817);
and UO_1553 (O_1553,N_14800,N_14870);
nand UO_1554 (O_1554,N_14997,N_14467);
nor UO_1555 (O_1555,N_14288,N_14903);
nor UO_1556 (O_1556,N_14473,N_14692);
nor UO_1557 (O_1557,N_14293,N_14339);
nand UO_1558 (O_1558,N_14508,N_14586);
and UO_1559 (O_1559,N_14952,N_14592);
or UO_1560 (O_1560,N_14265,N_14935);
or UO_1561 (O_1561,N_14528,N_14895);
and UO_1562 (O_1562,N_14876,N_14542);
nor UO_1563 (O_1563,N_14440,N_14525);
and UO_1564 (O_1564,N_14612,N_14933);
and UO_1565 (O_1565,N_14461,N_14691);
xnor UO_1566 (O_1566,N_14355,N_14261);
nor UO_1567 (O_1567,N_14582,N_14936);
nor UO_1568 (O_1568,N_14581,N_14900);
and UO_1569 (O_1569,N_14839,N_14983);
xor UO_1570 (O_1570,N_14400,N_14553);
nor UO_1571 (O_1571,N_14661,N_14457);
nor UO_1572 (O_1572,N_14957,N_14624);
and UO_1573 (O_1573,N_14776,N_14796);
and UO_1574 (O_1574,N_14897,N_14800);
nor UO_1575 (O_1575,N_14495,N_14494);
nand UO_1576 (O_1576,N_14284,N_14864);
or UO_1577 (O_1577,N_14395,N_14341);
nor UO_1578 (O_1578,N_14552,N_14919);
and UO_1579 (O_1579,N_14376,N_14336);
or UO_1580 (O_1580,N_14743,N_14393);
xor UO_1581 (O_1581,N_14337,N_14392);
or UO_1582 (O_1582,N_14570,N_14442);
and UO_1583 (O_1583,N_14844,N_14516);
or UO_1584 (O_1584,N_14849,N_14901);
nand UO_1585 (O_1585,N_14269,N_14703);
nand UO_1586 (O_1586,N_14832,N_14675);
nand UO_1587 (O_1587,N_14750,N_14495);
nand UO_1588 (O_1588,N_14902,N_14688);
or UO_1589 (O_1589,N_14866,N_14520);
nor UO_1590 (O_1590,N_14251,N_14592);
nor UO_1591 (O_1591,N_14559,N_14418);
xnor UO_1592 (O_1592,N_14970,N_14856);
nor UO_1593 (O_1593,N_14531,N_14353);
nor UO_1594 (O_1594,N_14748,N_14888);
and UO_1595 (O_1595,N_14890,N_14568);
or UO_1596 (O_1596,N_14687,N_14732);
and UO_1597 (O_1597,N_14882,N_14416);
or UO_1598 (O_1598,N_14594,N_14703);
and UO_1599 (O_1599,N_14801,N_14325);
nand UO_1600 (O_1600,N_14831,N_14512);
nand UO_1601 (O_1601,N_14743,N_14638);
nand UO_1602 (O_1602,N_14842,N_14736);
nor UO_1603 (O_1603,N_14814,N_14675);
or UO_1604 (O_1604,N_14449,N_14473);
nand UO_1605 (O_1605,N_14939,N_14409);
and UO_1606 (O_1606,N_14931,N_14969);
nor UO_1607 (O_1607,N_14859,N_14566);
nand UO_1608 (O_1608,N_14498,N_14529);
or UO_1609 (O_1609,N_14939,N_14662);
nand UO_1610 (O_1610,N_14914,N_14738);
and UO_1611 (O_1611,N_14806,N_14906);
nand UO_1612 (O_1612,N_14945,N_14925);
or UO_1613 (O_1613,N_14563,N_14945);
or UO_1614 (O_1614,N_14899,N_14538);
nand UO_1615 (O_1615,N_14797,N_14955);
or UO_1616 (O_1616,N_14371,N_14688);
or UO_1617 (O_1617,N_14785,N_14266);
nor UO_1618 (O_1618,N_14385,N_14568);
nand UO_1619 (O_1619,N_14657,N_14731);
nand UO_1620 (O_1620,N_14868,N_14824);
or UO_1621 (O_1621,N_14942,N_14655);
nand UO_1622 (O_1622,N_14612,N_14261);
or UO_1623 (O_1623,N_14337,N_14553);
and UO_1624 (O_1624,N_14468,N_14538);
nand UO_1625 (O_1625,N_14490,N_14819);
nand UO_1626 (O_1626,N_14364,N_14609);
or UO_1627 (O_1627,N_14352,N_14631);
nand UO_1628 (O_1628,N_14636,N_14572);
and UO_1629 (O_1629,N_14415,N_14914);
nor UO_1630 (O_1630,N_14645,N_14293);
nand UO_1631 (O_1631,N_14965,N_14629);
nor UO_1632 (O_1632,N_14389,N_14946);
nor UO_1633 (O_1633,N_14613,N_14293);
and UO_1634 (O_1634,N_14512,N_14796);
nand UO_1635 (O_1635,N_14972,N_14452);
or UO_1636 (O_1636,N_14255,N_14956);
nand UO_1637 (O_1637,N_14746,N_14315);
or UO_1638 (O_1638,N_14669,N_14782);
nand UO_1639 (O_1639,N_14815,N_14275);
or UO_1640 (O_1640,N_14366,N_14340);
nor UO_1641 (O_1641,N_14668,N_14285);
or UO_1642 (O_1642,N_14382,N_14863);
nor UO_1643 (O_1643,N_14740,N_14332);
or UO_1644 (O_1644,N_14873,N_14686);
and UO_1645 (O_1645,N_14854,N_14469);
nor UO_1646 (O_1646,N_14951,N_14423);
and UO_1647 (O_1647,N_14946,N_14553);
nor UO_1648 (O_1648,N_14910,N_14419);
or UO_1649 (O_1649,N_14252,N_14948);
and UO_1650 (O_1650,N_14403,N_14982);
and UO_1651 (O_1651,N_14643,N_14788);
and UO_1652 (O_1652,N_14876,N_14466);
and UO_1653 (O_1653,N_14319,N_14898);
nor UO_1654 (O_1654,N_14645,N_14818);
nor UO_1655 (O_1655,N_14263,N_14932);
nor UO_1656 (O_1656,N_14717,N_14531);
or UO_1657 (O_1657,N_14629,N_14773);
and UO_1658 (O_1658,N_14285,N_14803);
nand UO_1659 (O_1659,N_14767,N_14446);
and UO_1660 (O_1660,N_14851,N_14856);
nand UO_1661 (O_1661,N_14496,N_14394);
or UO_1662 (O_1662,N_14811,N_14615);
nand UO_1663 (O_1663,N_14321,N_14878);
nand UO_1664 (O_1664,N_14272,N_14487);
or UO_1665 (O_1665,N_14778,N_14981);
or UO_1666 (O_1666,N_14928,N_14350);
nor UO_1667 (O_1667,N_14257,N_14538);
xor UO_1668 (O_1668,N_14640,N_14525);
nor UO_1669 (O_1669,N_14411,N_14852);
or UO_1670 (O_1670,N_14793,N_14859);
and UO_1671 (O_1671,N_14344,N_14547);
nand UO_1672 (O_1672,N_14510,N_14659);
or UO_1673 (O_1673,N_14599,N_14692);
nand UO_1674 (O_1674,N_14749,N_14612);
nand UO_1675 (O_1675,N_14583,N_14462);
or UO_1676 (O_1676,N_14259,N_14815);
or UO_1677 (O_1677,N_14458,N_14592);
or UO_1678 (O_1678,N_14999,N_14815);
or UO_1679 (O_1679,N_14692,N_14427);
or UO_1680 (O_1680,N_14784,N_14817);
xnor UO_1681 (O_1681,N_14959,N_14817);
or UO_1682 (O_1682,N_14513,N_14377);
and UO_1683 (O_1683,N_14816,N_14300);
nand UO_1684 (O_1684,N_14921,N_14415);
or UO_1685 (O_1685,N_14615,N_14465);
or UO_1686 (O_1686,N_14484,N_14294);
or UO_1687 (O_1687,N_14351,N_14346);
nor UO_1688 (O_1688,N_14552,N_14275);
or UO_1689 (O_1689,N_14915,N_14700);
nor UO_1690 (O_1690,N_14895,N_14759);
and UO_1691 (O_1691,N_14725,N_14998);
nor UO_1692 (O_1692,N_14523,N_14640);
nor UO_1693 (O_1693,N_14435,N_14774);
nand UO_1694 (O_1694,N_14608,N_14660);
and UO_1695 (O_1695,N_14525,N_14952);
xnor UO_1696 (O_1696,N_14970,N_14984);
nand UO_1697 (O_1697,N_14824,N_14748);
nor UO_1698 (O_1698,N_14838,N_14697);
nand UO_1699 (O_1699,N_14573,N_14861);
nor UO_1700 (O_1700,N_14766,N_14596);
or UO_1701 (O_1701,N_14783,N_14383);
nand UO_1702 (O_1702,N_14902,N_14578);
or UO_1703 (O_1703,N_14319,N_14250);
and UO_1704 (O_1704,N_14853,N_14567);
xor UO_1705 (O_1705,N_14568,N_14782);
nand UO_1706 (O_1706,N_14600,N_14343);
nand UO_1707 (O_1707,N_14389,N_14961);
or UO_1708 (O_1708,N_14292,N_14357);
nor UO_1709 (O_1709,N_14524,N_14518);
nand UO_1710 (O_1710,N_14489,N_14987);
and UO_1711 (O_1711,N_14640,N_14624);
or UO_1712 (O_1712,N_14855,N_14390);
or UO_1713 (O_1713,N_14954,N_14898);
nor UO_1714 (O_1714,N_14404,N_14398);
nand UO_1715 (O_1715,N_14684,N_14923);
and UO_1716 (O_1716,N_14534,N_14373);
and UO_1717 (O_1717,N_14344,N_14481);
or UO_1718 (O_1718,N_14346,N_14784);
or UO_1719 (O_1719,N_14397,N_14992);
nand UO_1720 (O_1720,N_14845,N_14917);
nor UO_1721 (O_1721,N_14335,N_14363);
nand UO_1722 (O_1722,N_14640,N_14406);
and UO_1723 (O_1723,N_14810,N_14549);
nor UO_1724 (O_1724,N_14765,N_14745);
and UO_1725 (O_1725,N_14509,N_14859);
or UO_1726 (O_1726,N_14691,N_14503);
or UO_1727 (O_1727,N_14623,N_14379);
nand UO_1728 (O_1728,N_14903,N_14656);
nor UO_1729 (O_1729,N_14953,N_14866);
xor UO_1730 (O_1730,N_14975,N_14466);
or UO_1731 (O_1731,N_14598,N_14513);
nand UO_1732 (O_1732,N_14479,N_14608);
or UO_1733 (O_1733,N_14776,N_14785);
or UO_1734 (O_1734,N_14963,N_14449);
nor UO_1735 (O_1735,N_14669,N_14586);
or UO_1736 (O_1736,N_14862,N_14589);
nor UO_1737 (O_1737,N_14356,N_14998);
nand UO_1738 (O_1738,N_14680,N_14817);
nand UO_1739 (O_1739,N_14747,N_14828);
nand UO_1740 (O_1740,N_14578,N_14463);
nand UO_1741 (O_1741,N_14697,N_14773);
or UO_1742 (O_1742,N_14972,N_14755);
nor UO_1743 (O_1743,N_14450,N_14703);
nand UO_1744 (O_1744,N_14725,N_14958);
xnor UO_1745 (O_1745,N_14954,N_14844);
xnor UO_1746 (O_1746,N_14525,N_14435);
xnor UO_1747 (O_1747,N_14429,N_14649);
nor UO_1748 (O_1748,N_14432,N_14696);
xnor UO_1749 (O_1749,N_14616,N_14879);
and UO_1750 (O_1750,N_14505,N_14762);
nand UO_1751 (O_1751,N_14993,N_14712);
xnor UO_1752 (O_1752,N_14621,N_14339);
or UO_1753 (O_1753,N_14656,N_14342);
and UO_1754 (O_1754,N_14798,N_14572);
and UO_1755 (O_1755,N_14562,N_14704);
and UO_1756 (O_1756,N_14893,N_14397);
and UO_1757 (O_1757,N_14423,N_14339);
or UO_1758 (O_1758,N_14939,N_14475);
nand UO_1759 (O_1759,N_14635,N_14367);
nor UO_1760 (O_1760,N_14912,N_14286);
and UO_1761 (O_1761,N_14941,N_14277);
or UO_1762 (O_1762,N_14659,N_14454);
nor UO_1763 (O_1763,N_14636,N_14656);
and UO_1764 (O_1764,N_14432,N_14838);
or UO_1765 (O_1765,N_14348,N_14292);
or UO_1766 (O_1766,N_14827,N_14557);
and UO_1767 (O_1767,N_14888,N_14450);
nor UO_1768 (O_1768,N_14908,N_14938);
nor UO_1769 (O_1769,N_14607,N_14618);
nor UO_1770 (O_1770,N_14404,N_14575);
and UO_1771 (O_1771,N_14870,N_14644);
nor UO_1772 (O_1772,N_14294,N_14330);
or UO_1773 (O_1773,N_14990,N_14504);
and UO_1774 (O_1774,N_14406,N_14550);
nand UO_1775 (O_1775,N_14676,N_14675);
and UO_1776 (O_1776,N_14711,N_14886);
nand UO_1777 (O_1777,N_14412,N_14782);
or UO_1778 (O_1778,N_14782,N_14587);
xor UO_1779 (O_1779,N_14743,N_14824);
nor UO_1780 (O_1780,N_14457,N_14984);
or UO_1781 (O_1781,N_14530,N_14866);
and UO_1782 (O_1782,N_14363,N_14276);
nand UO_1783 (O_1783,N_14374,N_14449);
nor UO_1784 (O_1784,N_14296,N_14904);
or UO_1785 (O_1785,N_14637,N_14649);
nor UO_1786 (O_1786,N_14276,N_14989);
and UO_1787 (O_1787,N_14439,N_14426);
nand UO_1788 (O_1788,N_14885,N_14568);
or UO_1789 (O_1789,N_14770,N_14789);
and UO_1790 (O_1790,N_14760,N_14350);
and UO_1791 (O_1791,N_14820,N_14550);
or UO_1792 (O_1792,N_14322,N_14744);
nor UO_1793 (O_1793,N_14795,N_14495);
nand UO_1794 (O_1794,N_14437,N_14266);
nor UO_1795 (O_1795,N_14984,N_14823);
or UO_1796 (O_1796,N_14454,N_14631);
nand UO_1797 (O_1797,N_14575,N_14418);
or UO_1798 (O_1798,N_14406,N_14712);
xor UO_1799 (O_1799,N_14890,N_14311);
nand UO_1800 (O_1800,N_14316,N_14396);
nand UO_1801 (O_1801,N_14514,N_14300);
xnor UO_1802 (O_1802,N_14769,N_14530);
or UO_1803 (O_1803,N_14590,N_14784);
and UO_1804 (O_1804,N_14840,N_14274);
and UO_1805 (O_1805,N_14295,N_14539);
and UO_1806 (O_1806,N_14598,N_14349);
nor UO_1807 (O_1807,N_14324,N_14459);
nor UO_1808 (O_1808,N_14784,N_14501);
nor UO_1809 (O_1809,N_14571,N_14613);
or UO_1810 (O_1810,N_14290,N_14767);
nor UO_1811 (O_1811,N_14643,N_14404);
and UO_1812 (O_1812,N_14691,N_14900);
or UO_1813 (O_1813,N_14668,N_14284);
or UO_1814 (O_1814,N_14523,N_14768);
and UO_1815 (O_1815,N_14930,N_14473);
or UO_1816 (O_1816,N_14749,N_14939);
nor UO_1817 (O_1817,N_14378,N_14330);
and UO_1818 (O_1818,N_14355,N_14699);
nor UO_1819 (O_1819,N_14476,N_14296);
nand UO_1820 (O_1820,N_14786,N_14847);
nor UO_1821 (O_1821,N_14910,N_14830);
xor UO_1822 (O_1822,N_14580,N_14707);
and UO_1823 (O_1823,N_14594,N_14729);
or UO_1824 (O_1824,N_14376,N_14682);
or UO_1825 (O_1825,N_14622,N_14965);
and UO_1826 (O_1826,N_14763,N_14283);
and UO_1827 (O_1827,N_14742,N_14896);
nor UO_1828 (O_1828,N_14532,N_14768);
nand UO_1829 (O_1829,N_14362,N_14269);
nor UO_1830 (O_1830,N_14680,N_14589);
nand UO_1831 (O_1831,N_14467,N_14637);
or UO_1832 (O_1832,N_14816,N_14353);
nand UO_1833 (O_1833,N_14522,N_14909);
nor UO_1834 (O_1834,N_14874,N_14914);
and UO_1835 (O_1835,N_14501,N_14827);
nand UO_1836 (O_1836,N_14776,N_14788);
and UO_1837 (O_1837,N_14486,N_14658);
or UO_1838 (O_1838,N_14304,N_14635);
nor UO_1839 (O_1839,N_14620,N_14301);
and UO_1840 (O_1840,N_14929,N_14523);
and UO_1841 (O_1841,N_14395,N_14988);
or UO_1842 (O_1842,N_14457,N_14912);
nand UO_1843 (O_1843,N_14793,N_14515);
or UO_1844 (O_1844,N_14316,N_14452);
nand UO_1845 (O_1845,N_14902,N_14560);
nor UO_1846 (O_1846,N_14889,N_14488);
nand UO_1847 (O_1847,N_14772,N_14405);
or UO_1848 (O_1848,N_14440,N_14534);
nor UO_1849 (O_1849,N_14667,N_14305);
nand UO_1850 (O_1850,N_14808,N_14410);
or UO_1851 (O_1851,N_14559,N_14868);
or UO_1852 (O_1852,N_14937,N_14957);
or UO_1853 (O_1853,N_14724,N_14402);
nand UO_1854 (O_1854,N_14534,N_14730);
and UO_1855 (O_1855,N_14987,N_14545);
nand UO_1856 (O_1856,N_14366,N_14359);
nand UO_1857 (O_1857,N_14888,N_14352);
and UO_1858 (O_1858,N_14398,N_14823);
or UO_1859 (O_1859,N_14364,N_14269);
nor UO_1860 (O_1860,N_14853,N_14667);
nor UO_1861 (O_1861,N_14844,N_14418);
and UO_1862 (O_1862,N_14487,N_14641);
or UO_1863 (O_1863,N_14315,N_14587);
or UO_1864 (O_1864,N_14637,N_14937);
and UO_1865 (O_1865,N_14763,N_14544);
nor UO_1866 (O_1866,N_14500,N_14551);
nor UO_1867 (O_1867,N_14730,N_14741);
and UO_1868 (O_1868,N_14607,N_14579);
or UO_1869 (O_1869,N_14933,N_14460);
and UO_1870 (O_1870,N_14505,N_14786);
and UO_1871 (O_1871,N_14337,N_14837);
and UO_1872 (O_1872,N_14568,N_14398);
and UO_1873 (O_1873,N_14333,N_14931);
or UO_1874 (O_1874,N_14488,N_14403);
or UO_1875 (O_1875,N_14693,N_14608);
and UO_1876 (O_1876,N_14608,N_14521);
nand UO_1877 (O_1877,N_14767,N_14307);
nor UO_1878 (O_1878,N_14491,N_14296);
and UO_1879 (O_1879,N_14547,N_14505);
and UO_1880 (O_1880,N_14827,N_14615);
nor UO_1881 (O_1881,N_14329,N_14720);
or UO_1882 (O_1882,N_14516,N_14495);
nor UO_1883 (O_1883,N_14512,N_14839);
nor UO_1884 (O_1884,N_14911,N_14349);
or UO_1885 (O_1885,N_14373,N_14886);
nor UO_1886 (O_1886,N_14288,N_14930);
and UO_1887 (O_1887,N_14956,N_14891);
and UO_1888 (O_1888,N_14818,N_14610);
and UO_1889 (O_1889,N_14583,N_14345);
nor UO_1890 (O_1890,N_14854,N_14882);
or UO_1891 (O_1891,N_14354,N_14957);
nand UO_1892 (O_1892,N_14869,N_14639);
or UO_1893 (O_1893,N_14816,N_14886);
and UO_1894 (O_1894,N_14999,N_14561);
nand UO_1895 (O_1895,N_14792,N_14539);
nor UO_1896 (O_1896,N_14822,N_14769);
nor UO_1897 (O_1897,N_14914,N_14506);
nor UO_1898 (O_1898,N_14892,N_14645);
nor UO_1899 (O_1899,N_14564,N_14614);
nand UO_1900 (O_1900,N_14379,N_14468);
xnor UO_1901 (O_1901,N_14758,N_14507);
nor UO_1902 (O_1902,N_14550,N_14935);
and UO_1903 (O_1903,N_14752,N_14586);
or UO_1904 (O_1904,N_14676,N_14755);
nand UO_1905 (O_1905,N_14891,N_14464);
nand UO_1906 (O_1906,N_14984,N_14618);
or UO_1907 (O_1907,N_14958,N_14573);
nand UO_1908 (O_1908,N_14515,N_14702);
and UO_1909 (O_1909,N_14483,N_14706);
nor UO_1910 (O_1910,N_14536,N_14605);
or UO_1911 (O_1911,N_14301,N_14798);
nand UO_1912 (O_1912,N_14341,N_14672);
nand UO_1913 (O_1913,N_14320,N_14509);
nor UO_1914 (O_1914,N_14304,N_14521);
nand UO_1915 (O_1915,N_14848,N_14459);
nand UO_1916 (O_1916,N_14784,N_14396);
nor UO_1917 (O_1917,N_14282,N_14718);
or UO_1918 (O_1918,N_14755,N_14595);
nand UO_1919 (O_1919,N_14843,N_14424);
xnor UO_1920 (O_1920,N_14322,N_14638);
and UO_1921 (O_1921,N_14566,N_14449);
or UO_1922 (O_1922,N_14792,N_14392);
nand UO_1923 (O_1923,N_14974,N_14729);
xor UO_1924 (O_1924,N_14674,N_14483);
or UO_1925 (O_1925,N_14641,N_14708);
or UO_1926 (O_1926,N_14809,N_14804);
or UO_1927 (O_1927,N_14743,N_14544);
and UO_1928 (O_1928,N_14905,N_14979);
and UO_1929 (O_1929,N_14787,N_14789);
nand UO_1930 (O_1930,N_14446,N_14996);
nand UO_1931 (O_1931,N_14570,N_14561);
nand UO_1932 (O_1932,N_14672,N_14983);
nor UO_1933 (O_1933,N_14473,N_14517);
or UO_1934 (O_1934,N_14514,N_14720);
or UO_1935 (O_1935,N_14981,N_14839);
or UO_1936 (O_1936,N_14769,N_14913);
and UO_1937 (O_1937,N_14504,N_14577);
and UO_1938 (O_1938,N_14892,N_14514);
nand UO_1939 (O_1939,N_14827,N_14969);
or UO_1940 (O_1940,N_14305,N_14855);
nand UO_1941 (O_1941,N_14457,N_14873);
or UO_1942 (O_1942,N_14490,N_14283);
nand UO_1943 (O_1943,N_14777,N_14905);
or UO_1944 (O_1944,N_14550,N_14723);
or UO_1945 (O_1945,N_14630,N_14806);
xnor UO_1946 (O_1946,N_14872,N_14507);
nor UO_1947 (O_1947,N_14389,N_14552);
xor UO_1948 (O_1948,N_14302,N_14671);
nand UO_1949 (O_1949,N_14330,N_14354);
and UO_1950 (O_1950,N_14996,N_14345);
or UO_1951 (O_1951,N_14812,N_14500);
nand UO_1952 (O_1952,N_14504,N_14749);
or UO_1953 (O_1953,N_14490,N_14575);
or UO_1954 (O_1954,N_14509,N_14372);
nor UO_1955 (O_1955,N_14431,N_14992);
nand UO_1956 (O_1956,N_14324,N_14506);
or UO_1957 (O_1957,N_14744,N_14746);
and UO_1958 (O_1958,N_14552,N_14604);
nand UO_1959 (O_1959,N_14957,N_14644);
and UO_1960 (O_1960,N_14439,N_14812);
xor UO_1961 (O_1961,N_14395,N_14796);
nand UO_1962 (O_1962,N_14904,N_14739);
nor UO_1963 (O_1963,N_14315,N_14263);
nor UO_1964 (O_1964,N_14438,N_14756);
nor UO_1965 (O_1965,N_14770,N_14805);
nor UO_1966 (O_1966,N_14941,N_14521);
nor UO_1967 (O_1967,N_14569,N_14312);
and UO_1968 (O_1968,N_14950,N_14617);
or UO_1969 (O_1969,N_14946,N_14901);
nand UO_1970 (O_1970,N_14604,N_14567);
or UO_1971 (O_1971,N_14273,N_14971);
or UO_1972 (O_1972,N_14814,N_14420);
nor UO_1973 (O_1973,N_14775,N_14973);
nand UO_1974 (O_1974,N_14718,N_14994);
nor UO_1975 (O_1975,N_14491,N_14574);
nor UO_1976 (O_1976,N_14715,N_14557);
or UO_1977 (O_1977,N_14569,N_14334);
or UO_1978 (O_1978,N_14981,N_14547);
nor UO_1979 (O_1979,N_14359,N_14508);
nor UO_1980 (O_1980,N_14779,N_14763);
and UO_1981 (O_1981,N_14710,N_14676);
and UO_1982 (O_1982,N_14433,N_14880);
nor UO_1983 (O_1983,N_14455,N_14411);
or UO_1984 (O_1984,N_14930,N_14912);
nand UO_1985 (O_1985,N_14793,N_14905);
and UO_1986 (O_1986,N_14973,N_14592);
nor UO_1987 (O_1987,N_14292,N_14498);
nor UO_1988 (O_1988,N_14577,N_14669);
nor UO_1989 (O_1989,N_14730,N_14919);
nand UO_1990 (O_1990,N_14326,N_14743);
or UO_1991 (O_1991,N_14372,N_14566);
and UO_1992 (O_1992,N_14362,N_14974);
or UO_1993 (O_1993,N_14779,N_14343);
nor UO_1994 (O_1994,N_14817,N_14434);
and UO_1995 (O_1995,N_14986,N_14412);
and UO_1996 (O_1996,N_14405,N_14950);
or UO_1997 (O_1997,N_14639,N_14854);
and UO_1998 (O_1998,N_14425,N_14284);
nand UO_1999 (O_1999,N_14730,N_14823);
endmodule