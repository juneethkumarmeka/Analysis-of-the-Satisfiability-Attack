module basic_1500_15000_2000_5_levels_10xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
or U0 (N_0,In_994,In_463);
or U1 (N_1,In_1186,In_377);
or U2 (N_2,In_1148,In_584);
xnor U3 (N_3,In_105,In_870);
nor U4 (N_4,In_1291,In_383);
or U5 (N_5,In_77,In_1457);
xnor U6 (N_6,In_173,In_20);
or U7 (N_7,In_973,In_165);
xor U8 (N_8,In_408,In_1007);
or U9 (N_9,In_739,In_495);
nor U10 (N_10,In_1162,In_258);
xnor U11 (N_11,In_751,In_1089);
xor U12 (N_12,In_796,In_915);
nor U13 (N_13,In_1355,In_855);
nand U14 (N_14,In_129,In_1410);
nand U15 (N_15,In_656,In_638);
or U16 (N_16,In_1102,In_347);
and U17 (N_17,In_271,In_445);
or U18 (N_18,In_810,In_1404);
xor U19 (N_19,In_1121,In_1100);
nand U20 (N_20,In_1422,In_7);
xnor U21 (N_21,In_1199,In_1456);
nor U22 (N_22,In_261,In_663);
nand U23 (N_23,In_373,In_916);
xnor U24 (N_24,In_322,In_812);
and U25 (N_25,In_324,In_1172);
and U26 (N_26,In_543,In_542);
xnor U27 (N_27,In_1015,In_795);
nand U28 (N_28,In_1223,In_244);
nand U29 (N_29,In_110,In_597);
and U30 (N_30,In_717,In_200);
nor U31 (N_31,In_1224,In_306);
or U32 (N_32,In_1308,In_1282);
xor U33 (N_33,In_867,In_699);
nor U34 (N_34,In_202,In_166);
nand U35 (N_35,In_201,In_1117);
nand U36 (N_36,In_1154,In_520);
xor U37 (N_37,In_159,In_706);
nand U38 (N_38,In_1055,In_102);
xnor U39 (N_39,In_1363,In_466);
nor U40 (N_40,In_884,In_1019);
nand U41 (N_41,In_1315,In_1240);
nor U42 (N_42,In_1392,In_483);
and U43 (N_43,In_797,In_1150);
and U44 (N_44,In_835,In_344);
and U45 (N_45,In_1462,In_1129);
or U46 (N_46,In_553,In_960);
nor U47 (N_47,In_632,In_1083);
xor U48 (N_48,In_147,In_1396);
xnor U49 (N_49,In_1384,In_729);
nand U50 (N_50,In_397,In_1445);
and U51 (N_51,In_1173,In_1274);
xor U52 (N_52,In_414,In_177);
xor U53 (N_53,In_277,In_1378);
xnor U54 (N_54,In_137,In_1185);
nand U55 (N_55,In_66,In_395);
xnor U56 (N_56,In_1249,In_907);
and U57 (N_57,In_874,In_227);
nand U58 (N_58,In_711,In_278);
nand U59 (N_59,In_279,In_1234);
xor U60 (N_60,In_684,In_472);
nor U61 (N_61,In_903,In_1080);
nand U62 (N_62,In_438,In_672);
xor U63 (N_63,In_898,In_492);
and U64 (N_64,In_1218,In_1229);
and U65 (N_65,In_253,In_231);
nor U66 (N_66,In_1027,In_1081);
nor U67 (N_67,In_735,In_1372);
nand U68 (N_68,In_963,In_1295);
and U69 (N_69,In_561,In_134);
nand U70 (N_70,In_753,In_1245);
and U71 (N_71,In_103,In_1072);
and U72 (N_72,In_409,In_404);
xnor U73 (N_73,In_303,In_1478);
or U74 (N_74,In_1464,In_1495);
nand U75 (N_75,In_539,In_487);
nand U76 (N_76,In_60,In_1443);
nor U77 (N_77,In_815,In_698);
or U78 (N_78,In_1092,In_386);
nand U79 (N_79,In_384,In_170);
xnor U80 (N_80,In_872,In_741);
xnor U81 (N_81,In_862,In_673);
nand U82 (N_82,In_164,In_1426);
and U83 (N_83,In_1126,In_636);
and U84 (N_84,In_692,In_136);
nand U85 (N_85,In_1451,In_908);
nand U86 (N_86,In_484,In_1269);
or U87 (N_87,In_1198,In_285);
or U88 (N_88,In_1023,In_993);
nor U89 (N_89,In_28,In_189);
or U90 (N_90,In_219,In_1119);
nand U91 (N_91,In_167,In_1267);
and U92 (N_92,In_233,In_922);
nand U93 (N_93,In_1020,In_410);
xnor U94 (N_94,In_1242,In_175);
xnor U95 (N_95,In_1319,In_49);
xnor U96 (N_96,In_462,In_932);
nand U97 (N_97,In_881,In_834);
and U98 (N_98,In_567,In_947);
nand U99 (N_99,In_1367,In_390);
and U100 (N_100,In_118,In_930);
or U101 (N_101,In_1140,In_215);
xor U102 (N_102,In_1303,In_3);
xor U103 (N_103,In_599,In_1491);
or U104 (N_104,In_1048,In_1111);
and U105 (N_105,In_419,In_671);
and U106 (N_106,In_512,In_995);
and U107 (N_107,In_1460,In_1429);
and U108 (N_108,In_133,In_1196);
and U109 (N_109,In_548,In_989);
xor U110 (N_110,In_1473,In_582);
nand U111 (N_111,In_239,In_267);
xnor U112 (N_112,In_935,In_157);
nand U113 (N_113,In_878,In_1062);
xor U114 (N_114,In_1005,In_55);
and U115 (N_115,In_73,In_1311);
and U116 (N_116,In_427,In_356);
and U117 (N_117,In_762,In_986);
nand U118 (N_118,In_961,In_1304);
and U119 (N_119,In_65,In_413);
nand U120 (N_120,In_1342,In_1492);
and U121 (N_121,In_152,In_603);
and U122 (N_122,In_1217,In_1123);
and U123 (N_123,In_148,In_689);
nand U124 (N_124,In_1003,In_422);
xor U125 (N_125,In_1167,In_280);
nor U126 (N_126,In_199,In_1400);
nand U127 (N_127,In_194,In_1493);
and U128 (N_128,In_593,In_92);
or U129 (N_129,In_1268,In_926);
or U130 (N_130,In_153,In_400);
or U131 (N_131,In_155,In_1037);
xor U132 (N_132,In_658,In_1250);
nor U133 (N_133,In_868,In_300);
or U134 (N_134,In_311,In_851);
xnor U135 (N_135,In_772,In_140);
and U136 (N_136,In_666,In_744);
xor U137 (N_137,In_1133,In_708);
and U138 (N_138,In_398,In_1323);
xor U139 (N_139,In_1135,In_578);
nand U140 (N_140,In_1236,In_508);
xnor U141 (N_141,In_992,In_864);
and U142 (N_142,In_1307,In_837);
and U143 (N_143,In_363,In_1439);
nand U144 (N_144,In_909,In_1216);
or U145 (N_145,In_1090,In_1278);
nor U146 (N_146,In_904,In_591);
and U147 (N_147,In_1043,In_1352);
or U148 (N_148,In_920,In_1051);
or U149 (N_149,In_720,In_357);
nor U150 (N_150,In_873,In_798);
nor U151 (N_151,In_607,In_212);
and U152 (N_152,In_968,In_610);
nor U153 (N_153,In_1130,In_559);
xnor U154 (N_154,In_1275,In_1064);
xor U155 (N_155,In_13,In_293);
xnor U156 (N_156,In_1298,In_132);
and U157 (N_157,In_565,In_1287);
or U158 (N_158,In_1309,In_191);
and U159 (N_159,In_645,In_382);
or U160 (N_160,In_43,In_417);
and U161 (N_161,In_830,In_564);
nor U162 (N_162,In_845,In_1115);
and U163 (N_163,In_576,In_707);
and U164 (N_164,In_563,In_1440);
nand U165 (N_165,In_475,In_63);
or U166 (N_166,In_1138,In_447);
or U167 (N_167,In_1073,In_195);
nand U168 (N_168,In_635,In_45);
xor U169 (N_169,In_710,In_1207);
xnor U170 (N_170,In_31,In_583);
and U171 (N_171,In_81,In_1000);
and U172 (N_172,In_977,In_911);
and U173 (N_173,In_449,In_641);
or U174 (N_174,In_613,In_323);
nor U175 (N_175,In_499,In_1262);
nor U176 (N_176,In_946,In_704);
nor U177 (N_177,In_524,In_53);
nand U178 (N_178,In_1095,In_282);
or U179 (N_179,In_522,In_469);
nor U180 (N_180,In_976,In_198);
or U181 (N_181,In_683,In_1159);
nor U182 (N_182,In_1455,In_997);
and U183 (N_183,In_1347,In_560);
xnor U184 (N_184,In_885,In_262);
nand U185 (N_185,In_1403,In_566);
xnor U186 (N_186,In_1407,In_33);
xnor U187 (N_187,In_75,In_677);
and U188 (N_188,In_1345,In_824);
and U189 (N_189,In_573,In_1335);
or U190 (N_190,In_435,In_256);
and U191 (N_191,In_1132,In_819);
and U192 (N_192,In_631,In_661);
nor U193 (N_193,In_954,In_1255);
and U194 (N_194,In_161,In_245);
xor U195 (N_195,In_62,In_1034);
xor U196 (N_196,In_1299,In_85);
or U197 (N_197,In_1060,In_72);
xor U198 (N_198,In_305,In_432);
nor U199 (N_199,In_728,In_1099);
or U200 (N_200,In_1297,In_1428);
or U201 (N_201,In_442,In_491);
nand U202 (N_202,In_959,In_1074);
xnor U203 (N_203,In_1373,In_682);
or U204 (N_204,In_655,In_1344);
and U205 (N_205,In_93,In_80);
nor U206 (N_206,In_817,In_336);
nand U207 (N_207,In_224,In_1273);
xor U208 (N_208,In_241,In_82);
or U209 (N_209,In_604,In_204);
or U210 (N_210,In_957,In_730);
nand U211 (N_211,In_326,In_1178);
nand U212 (N_212,In_828,In_42);
nand U213 (N_213,In_117,In_1340);
xor U214 (N_214,In_289,In_138);
and U215 (N_215,In_562,In_1014);
xnor U216 (N_216,In_467,In_489);
nor U217 (N_217,In_251,In_1409);
nand U218 (N_218,In_10,In_470);
nor U219 (N_219,In_1179,In_374);
nand U220 (N_220,In_446,In_154);
or U221 (N_221,In_1243,In_473);
xnor U222 (N_222,In_813,In_1393);
nand U223 (N_223,In_998,In_83);
nand U224 (N_224,In_1017,In_1168);
or U225 (N_225,In_1305,In_1353);
nand U226 (N_226,In_1024,In_950);
and U227 (N_227,In_95,In_625);
xnor U228 (N_228,In_1324,In_1227);
and U229 (N_229,In_338,In_1124);
xor U230 (N_230,In_951,In_1477);
nand U231 (N_231,In_925,In_19);
nor U232 (N_232,In_126,In_601);
nor U233 (N_233,In_1012,In_853);
nand U234 (N_234,In_1244,In_498);
nand U235 (N_235,In_768,In_273);
or U236 (N_236,In_1200,In_1164);
or U237 (N_237,In_1257,In_1106);
and U238 (N_238,In_517,In_1076);
and U239 (N_239,In_274,In_431);
nand U240 (N_240,In_927,In_931);
nand U241 (N_241,In_680,In_1412);
and U242 (N_242,In_169,In_142);
or U243 (N_243,In_35,In_365);
xnor U244 (N_244,In_307,In_1052);
xnor U245 (N_245,In_220,In_379);
and U246 (N_246,In_1221,In_724);
xor U247 (N_247,In_691,In_1112);
and U248 (N_248,In_718,In_600);
nand U249 (N_249,In_1075,In_809);
or U250 (N_250,In_296,In_1388);
nor U251 (N_251,In_1487,In_1417);
or U252 (N_252,In_1433,In_1086);
or U253 (N_253,In_24,In_1390);
or U254 (N_254,In_1,In_807);
and U255 (N_255,In_1375,In_1424);
or U256 (N_256,In_1071,In_1006);
nor U257 (N_257,In_702,In_918);
nand U258 (N_258,In_1193,In_521);
nand U259 (N_259,In_722,In_353);
and U260 (N_260,In_1341,In_1039);
and U261 (N_261,In_263,In_98);
xor U262 (N_262,In_971,In_331);
or U263 (N_263,In_847,In_1110);
nor U264 (N_264,In_709,In_569);
nand U265 (N_265,In_1206,In_122);
and U266 (N_266,In_90,In_1471);
xnor U267 (N_267,In_1016,In_767);
xor U268 (N_268,In_1430,In_1098);
nor U269 (N_269,In_1449,In_747);
or U270 (N_270,In_380,In_1021);
or U271 (N_271,In_1266,In_158);
nor U272 (N_272,In_388,In_477);
nand U273 (N_273,In_1067,In_705);
nand U274 (N_274,In_1408,In_940);
or U275 (N_275,In_1056,In_291);
or U276 (N_276,In_308,In_1225);
and U277 (N_277,In_877,In_779);
xnor U278 (N_278,In_39,In_283);
nor U279 (N_279,In_1070,In_646);
or U280 (N_280,In_433,In_1452);
nor U281 (N_281,In_1170,In_823);
or U282 (N_282,In_1038,In_953);
xor U283 (N_283,In_1033,In_89);
nand U284 (N_284,In_1141,In_642);
nand U285 (N_285,In_459,In_314);
nor U286 (N_286,In_574,In_76);
and U287 (N_287,In_733,In_162);
and U288 (N_288,In_1143,In_1108);
xor U289 (N_289,In_69,In_203);
nand U290 (N_290,In_1368,In_1394);
xor U291 (N_291,In_242,In_660);
nand U292 (N_292,In_890,In_782);
and U293 (N_293,In_501,In_125);
nor U294 (N_294,In_448,In_549);
nor U295 (N_295,In_701,In_135);
nor U296 (N_296,In_1204,In_1316);
or U297 (N_297,In_1416,In_319);
xnor U298 (N_298,In_1087,In_939);
xnor U299 (N_299,In_455,In_123);
nand U300 (N_300,In_690,In_52);
or U301 (N_301,In_131,In_630);
and U302 (N_302,In_956,In_727);
nor U303 (N_303,In_965,In_313);
xnor U304 (N_304,In_674,In_493);
nor U305 (N_305,In_206,In_974);
nor U306 (N_306,In_115,In_770);
nand U307 (N_307,In_30,In_511);
xor U308 (N_308,In_1018,In_1151);
nor U309 (N_309,In_1238,In_286);
nand U310 (N_310,In_1271,In_91);
or U311 (N_311,In_179,In_468);
or U312 (N_312,In_236,In_776);
or U313 (N_313,In_647,In_50);
xnor U314 (N_314,In_309,In_248);
and U315 (N_315,In_1166,In_514);
and U316 (N_316,In_988,In_765);
or U317 (N_317,In_737,In_889);
or U318 (N_318,In_1283,In_742);
xor U319 (N_319,In_1157,In_943);
nor U320 (N_320,In_376,In_844);
xnor U321 (N_321,In_1128,In_608);
and U322 (N_322,In_958,In_478);
nand U323 (N_323,In_128,In_633);
xor U324 (N_324,In_1049,In_1369);
or U325 (N_325,In_420,In_1435);
xor U326 (N_326,In_355,In_385);
or U327 (N_327,In_1374,In_500);
or U328 (N_328,In_425,In_228);
and U329 (N_329,In_457,In_1284);
nand U330 (N_330,In_1009,In_387);
nor U331 (N_331,In_1091,In_465);
xnor U332 (N_332,In_151,In_577);
and U333 (N_333,In_537,In_726);
and U334 (N_334,In_910,In_688);
or U335 (N_335,In_952,In_679);
or U336 (N_336,In_1187,In_1097);
nor U337 (N_337,In_453,In_1125);
nor U338 (N_338,In_1285,In_1254);
xnor U339 (N_339,In_1028,In_96);
nand U340 (N_340,In_987,In_972);
nand U341 (N_341,In_748,In_1155);
nor U342 (N_342,In_145,In_32);
nor U343 (N_343,In_866,In_174);
xnor U344 (N_344,In_854,In_528);
and U345 (N_345,In_840,In_257);
and U346 (N_346,In_415,In_111);
and U347 (N_347,In_523,In_452);
nor U348 (N_348,In_361,In_757);
nor U349 (N_349,In_801,In_1175);
xor U350 (N_350,In_675,In_615);
xnor U351 (N_351,In_1068,In_299);
or U352 (N_352,In_1183,In_1362);
nand U353 (N_353,In_394,In_21);
or U354 (N_354,In_571,In_57);
nor U355 (N_355,In_980,In_1177);
or U356 (N_356,In_1475,In_1398);
nor U357 (N_357,In_1136,In_247);
and U358 (N_358,In_1431,In_964);
or U359 (N_359,In_506,In_79);
nor U360 (N_360,In_222,In_846);
nor U361 (N_361,In_476,In_766);
nor U362 (N_362,In_1359,In_121);
xnor U363 (N_363,In_101,In_1358);
nand U364 (N_364,In_962,In_693);
xor U365 (N_365,In_156,In_1251);
xnor U366 (N_366,In_315,In_749);
nor U367 (N_367,In_1467,In_301);
nor U368 (N_368,In_586,In_1153);
xor U369 (N_369,In_61,In_1114);
nand U370 (N_370,In_1182,In_350);
and U371 (N_371,In_769,In_783);
nor U372 (N_372,In_970,In_186);
nand U373 (N_373,In_474,In_1010);
or U374 (N_374,In_1171,In_1330);
or U375 (N_375,In_507,In_1228);
xor U376 (N_376,In_1453,In_1397);
and U377 (N_377,In_1226,In_536);
nand U378 (N_378,In_1025,In_1399);
or U379 (N_379,In_1231,In_1146);
or U380 (N_380,In_525,In_270);
xor U381 (N_381,In_1263,In_1061);
or U382 (N_382,In_502,In_503);
nor U383 (N_383,In_1205,In_981);
nor U384 (N_384,In_1041,In_183);
or U385 (N_385,In_771,In_160);
nand U386 (N_386,In_1265,In_401);
and U387 (N_387,In_168,In_781);
or U388 (N_388,In_1279,In_287);
xnor U389 (N_389,In_1122,In_345);
nor U390 (N_390,In_71,In_668);
nor U391 (N_391,In_141,In_354);
or U392 (N_392,In_371,In_942);
or U393 (N_393,In_1022,In_624);
and U394 (N_394,In_1192,In_1239);
xnor U395 (N_395,In_1063,In_1446);
nor U396 (N_396,In_295,In_598);
xor U397 (N_397,In_23,In_255);
or U398 (N_398,In_617,In_649);
and U399 (N_399,In_450,In_1026);
nand U400 (N_400,In_1360,In_1292);
nor U401 (N_401,In_1137,In_1450);
and U402 (N_402,In_780,In_288);
xor U403 (N_403,In_436,In_1253);
nor U404 (N_404,In_1296,In_205);
nand U405 (N_405,In_1474,In_70);
or U406 (N_406,In_1461,In_1211);
or U407 (N_407,In_944,In_541);
or U408 (N_408,In_1486,In_1120);
or U409 (N_409,In_1194,In_696);
or U410 (N_410,In_1142,In_1105);
or U411 (N_411,In_831,In_622);
nor U412 (N_412,In_513,In_572);
and U413 (N_413,In_94,In_213);
xor U414 (N_414,In_1413,In_334);
and U415 (N_415,In_15,In_454);
and U416 (N_416,In_1322,In_421);
xor U417 (N_417,In_1259,In_1351);
nand U418 (N_418,In_529,In_1288);
nand U419 (N_419,In_694,In_58);
and U420 (N_420,In_510,In_490);
and U421 (N_421,In_917,In_1332);
nor U422 (N_422,In_1482,In_480);
or U423 (N_423,In_34,In_290);
xor U424 (N_424,In_556,In_806);
and U425 (N_425,In_609,In_1195);
and U426 (N_426,In_188,In_1107);
nand U427 (N_427,In_197,In_746);
or U428 (N_428,In_518,In_1383);
nor U429 (N_429,In_337,In_298);
or U430 (N_430,In_12,In_1047);
nand U431 (N_431,In_822,In_1045);
nand U432 (N_432,In_1405,In_805);
nor U433 (N_433,In_914,In_1277);
or U434 (N_434,In_265,In_629);
nor U435 (N_435,In_996,In_399);
xnor U436 (N_436,In_731,In_1468);
nand U437 (N_437,In_378,In_1432);
and U438 (N_438,In_1290,In_217);
nor U439 (N_439,In_1088,In_348);
nand U440 (N_440,In_403,In_1069);
or U441 (N_441,In_312,In_619);
and U442 (N_442,In_848,In_897);
or U443 (N_443,In_1312,In_859);
xor U444 (N_444,In_112,In_602);
nor U445 (N_445,In_934,In_392);
nand U446 (N_446,In_1203,In_1260);
or U447 (N_447,In_310,In_1050);
xnor U448 (N_448,In_342,In_614);
xnor U449 (N_449,In_424,In_193);
xnor U450 (N_450,In_1113,In_1215);
or U451 (N_451,In_46,In_339);
and U452 (N_452,In_1078,In_437);
nor U453 (N_453,In_1427,In_941);
or U454 (N_454,In_650,In_856);
nand U455 (N_455,In_1310,In_329);
and U456 (N_456,In_370,In_252);
and U457 (N_457,In_393,In_955);
or U458 (N_458,In_734,In_181);
nor U459 (N_459,In_341,In_1233);
or U460 (N_460,In_725,In_626);
xor U461 (N_461,In_999,In_893);
nor U462 (N_462,In_1160,In_349);
nor U463 (N_463,In_1036,In_428);
and U464 (N_464,In_552,In_533);
or U465 (N_465,In_736,In_1145);
xor U466 (N_466,In_761,In_802);
or U467 (N_467,In_544,In_929);
nor U468 (N_468,In_557,In_1189);
nor U469 (N_469,In_829,In_894);
and U470 (N_470,In_527,In_555);
or U471 (N_471,In_1371,In_1096);
nand U472 (N_472,In_665,In_1382);
nor U473 (N_473,In_892,In_87);
xnor U474 (N_474,In_1219,In_16);
or U475 (N_475,In_1356,In_444);
xnor U476 (N_476,In_1437,In_1414);
and U477 (N_477,In_333,In_358);
or U478 (N_478,In_494,In_697);
and U479 (N_479,In_1326,In_1208);
or U480 (N_480,In_1389,In_25);
or U481 (N_481,In_237,In_1476);
and U482 (N_482,In_643,In_818);
nor U483 (N_483,In_461,In_715);
or U484 (N_484,In_865,In_654);
xnor U485 (N_485,In_302,In_1436);
nor U486 (N_486,In_686,In_1008);
nand U487 (N_487,In_209,In_732);
nor U488 (N_488,In_621,In_1498);
nand U489 (N_489,In_1101,In_86);
nand U490 (N_490,In_1011,In_412);
and U491 (N_491,In_804,In_416);
xor U492 (N_492,In_575,In_225);
xnor U493 (N_493,In_1386,In_1261);
or U494 (N_494,In_841,In_616);
and U495 (N_495,In_1441,In_40);
nand U496 (N_496,In_924,In_1480);
or U497 (N_497,In_628,In_1118);
nand U498 (N_498,In_238,In_667);
xor U499 (N_499,In_990,In_451);
and U500 (N_500,In_568,In_871);
or U501 (N_501,In_1210,In_208);
and U502 (N_502,In_1066,In_481);
xor U503 (N_503,In_116,In_187);
or U504 (N_504,In_443,In_406);
xnor U505 (N_505,In_1059,In_249);
nor U506 (N_506,In_367,In_662);
or U507 (N_507,In_664,In_836);
or U508 (N_508,In_594,In_1448);
nand U509 (N_509,In_1329,In_687);
and U510 (N_510,In_790,In_721);
xor U511 (N_511,In_1201,In_785);
xnor U512 (N_512,In_670,In_1212);
or U513 (N_513,In_429,In_1246);
nor U514 (N_514,In_1419,In_1302);
nor U515 (N_515,In_1222,In_814);
nand U516 (N_516,In_1376,In_226);
xor U517 (N_517,In_411,In_928);
and U518 (N_518,In_1489,In_18);
nand U519 (N_519,In_6,In_588);
nor U520 (N_520,In_786,In_106);
or U521 (N_521,In_254,In_328);
nand U522 (N_522,In_669,In_886);
nand U523 (N_523,In_1381,In_945);
nor U524 (N_524,In_832,In_281);
and U525 (N_525,In_214,In_869);
nor U526 (N_526,In_109,In_1169);
and U527 (N_527,In_1272,In_612);
nand U528 (N_528,In_74,In_763);
xor U529 (N_529,In_838,In_1191);
nor U530 (N_530,In_975,In_434);
xor U531 (N_531,In_857,In_794);
or U532 (N_532,In_485,In_1209);
nor U533 (N_533,In_139,In_891);
nor U534 (N_534,In_774,In_888);
xnor U535 (N_535,In_861,In_1454);
or U536 (N_536,In_405,In_1001);
xnor U537 (N_537,In_863,In_146);
and U538 (N_538,In_816,In_531);
nand U539 (N_539,In_1044,In_933);
xnor U540 (N_540,In_372,In_723);
nand U541 (N_541,In_912,In_784);
xnor U542 (N_542,In_496,In_519);
nand U543 (N_543,In_1002,In_1214);
xnor U544 (N_544,In_464,In_368);
nand U545 (N_545,In_232,In_1156);
or U546 (N_546,In_9,In_713);
and U547 (N_547,In_595,In_243);
xnor U548 (N_548,In_876,In_259);
nor U549 (N_549,In_700,In_740);
nand U550 (N_550,In_107,In_1472);
nor U551 (N_551,In_852,In_1029);
xnor U552 (N_552,In_27,In_811);
nor U553 (N_553,In_130,In_5);
nor U554 (N_554,In_1294,In_800);
and U555 (N_555,In_983,In_1377);
or U556 (N_556,In_570,In_360);
and U557 (N_557,In_266,In_879);
nor U558 (N_558,In_1438,In_272);
xor U559 (N_559,In_540,In_407);
and U560 (N_560,In_104,In_606);
or U561 (N_561,In_64,In_396);
and U562 (N_562,In_221,In_919);
xor U563 (N_563,In_547,In_1289);
or U564 (N_564,In_332,In_1385);
and U565 (N_565,In_51,In_11);
or U566 (N_566,In_1354,In_505);
nor U567 (N_567,In_991,In_1174);
nor U568 (N_568,In_596,In_1395);
nand U569 (N_569,In_778,In_850);
nor U570 (N_570,In_26,In_216);
nor U571 (N_571,In_842,In_14);
or U572 (N_572,In_755,In_471);
and U573 (N_573,In_1077,In_1084);
xnor U574 (N_574,In_1313,In_627);
nand U575 (N_575,In_230,In_937);
xnor U576 (N_576,In_1364,In_178);
or U577 (N_577,In_587,In_275);
or U578 (N_578,In_1337,In_789);
nor U579 (N_579,In_906,In_1248);
or U580 (N_580,In_497,In_48);
nand U581 (N_581,In_0,In_192);
and U582 (N_582,In_426,In_967);
nor U583 (N_583,In_88,In_882);
and U584 (N_584,In_144,In_590);
nor U585 (N_585,In_1336,In_196);
xor U586 (N_586,In_589,In_234);
or U587 (N_587,In_1349,In_317);
nand U588 (N_588,In_1065,In_678);
or U589 (N_589,In_1458,In_44);
nand U590 (N_590,In_1152,In_532);
and U591 (N_591,In_546,In_1479);
xor U592 (N_592,In_580,In_1483);
or U593 (N_593,In_37,In_764);
xor U594 (N_594,In_346,In_681);
nand U595 (N_595,In_659,In_826);
or U596 (N_596,In_223,In_1365);
xnor U597 (N_597,In_1004,In_738);
and U598 (N_598,In_1402,In_1237);
xor U599 (N_599,In_1109,In_369);
nor U600 (N_600,In_509,In_685);
nand U601 (N_601,In_551,In_895);
nor U602 (N_602,In_535,In_1366);
and U603 (N_603,In_843,In_381);
or U604 (N_604,In_1258,In_359);
and U605 (N_605,In_558,In_1497);
and U606 (N_606,In_849,In_340);
xnor U607 (N_607,In_440,In_1116);
nand U608 (N_608,In_488,In_54);
nand U609 (N_609,In_325,In_808);
nor U610 (N_610,In_1465,In_773);
nand U611 (N_611,In_210,In_949);
and U612 (N_612,In_1202,In_418);
or U613 (N_613,In_460,In_1180);
or U614 (N_614,In_150,In_240);
and U615 (N_615,In_1147,In_754);
or U616 (N_616,In_833,In_343);
or U617 (N_617,In_1348,In_352);
xor U618 (N_618,In_441,In_1481);
xor U619 (N_619,In_1357,In_585);
nand U620 (N_620,In_29,In_639);
nor U621 (N_621,In_1447,In_184);
and U622 (N_622,In_127,In_880);
xnor U623 (N_623,In_775,In_1387);
xor U624 (N_624,In_791,In_896);
and U625 (N_625,In_1276,In_482);
and U626 (N_626,In_56,In_297);
or U627 (N_627,In_839,In_182);
nand U628 (N_628,In_858,In_1470);
xor U629 (N_629,In_318,In_366);
nand U630 (N_630,In_1380,In_479);
nor U631 (N_631,In_1339,In_550);
or U632 (N_632,In_172,In_276);
nand U633 (N_633,In_375,In_268);
nand U634 (N_634,In_1082,In_391);
xnor U635 (N_635,In_579,In_1361);
or U636 (N_636,In_1176,In_1411);
and U637 (N_637,In_113,In_1197);
xnor U638 (N_638,In_788,In_269);
xor U639 (N_639,In_777,In_8);
xnor U640 (N_640,In_1434,In_486);
and U641 (N_641,In_1343,In_1032);
xor U642 (N_642,In_260,In_84);
or U643 (N_643,In_207,In_1163);
xor U644 (N_644,In_41,In_149);
xor U645 (N_645,In_456,In_623);
nand U646 (N_646,In_1421,In_787);
nor U647 (N_647,In_1318,In_821);
nand U648 (N_648,In_1494,In_703);
and U649 (N_649,In_554,In_1134);
or U650 (N_650,In_1103,In_321);
and U651 (N_651,In_294,In_1252);
or U652 (N_652,In_1490,In_1230);
nand U653 (N_653,In_905,In_923);
and U654 (N_654,In_676,In_250);
xor U655 (N_655,In_180,In_657);
xnor U656 (N_656,In_99,In_190);
and U657 (N_657,In_163,In_538);
or U658 (N_658,In_284,In_351);
or U659 (N_659,In_1415,In_1320);
xnor U660 (N_660,In_651,In_439);
xor U661 (N_661,In_1281,In_1423);
nand U662 (N_662,In_100,In_978);
or U663 (N_663,In_745,In_304);
and U664 (N_664,In_1093,In_108);
and U665 (N_665,In_185,In_330);
xnor U666 (N_666,In_1331,In_38);
nand U667 (N_667,In_860,In_1190);
nand U668 (N_668,In_752,In_712);
and U669 (N_669,In_1232,In_1264);
and U670 (N_670,In_2,In_875);
xnor U671 (N_671,In_1139,In_1256);
nand U672 (N_672,In_900,In_913);
xor U673 (N_673,In_1420,In_1328);
xnor U674 (N_674,In_1484,In_362);
nand U675 (N_675,In_652,In_68);
nand U676 (N_676,In_966,In_47);
nor U677 (N_677,In_1144,In_618);
nor U678 (N_678,In_936,In_1442);
or U679 (N_679,In_1499,In_264);
nand U680 (N_680,In_1333,In_1425);
and U681 (N_681,In_1321,In_1030);
and U682 (N_682,In_1235,In_1270);
xor U683 (N_683,In_1220,In_1042);
or U684 (N_684,In_176,In_1325);
and U685 (N_685,In_979,In_327);
xnor U686 (N_686,In_504,In_292);
nand U687 (N_687,In_534,In_526);
or U688 (N_688,In_124,In_423);
nor U689 (N_689,In_1293,In_1301);
xor U690 (N_690,In_1314,In_1040);
xnor U691 (N_691,In_793,In_760);
nand U692 (N_692,In_1188,In_1327);
nor U693 (N_693,In_1300,In_458);
xor U694 (N_694,In_634,In_887);
nor U695 (N_695,In_1161,In_756);
or U696 (N_696,In_901,In_581);
nand U697 (N_697,In_984,In_1418);
nand U698 (N_698,In_316,In_67);
and U699 (N_699,In_235,In_218);
nor U700 (N_700,In_1053,In_921);
and U701 (N_701,In_1131,In_750);
nor U702 (N_702,In_1469,In_1149);
or U703 (N_703,In_899,In_611);
and U704 (N_704,In_1338,In_1350);
and U705 (N_705,In_743,In_143);
nand U706 (N_706,In_36,In_78);
and U707 (N_707,In_4,In_1379);
nor U708 (N_708,In_1184,In_1444);
xnor U709 (N_709,In_389,In_22);
and U710 (N_710,In_653,In_1334);
xor U711 (N_711,In_902,In_1158);
and U712 (N_712,In_1046,In_640);
nor U713 (N_713,In_515,In_799);
xnor U714 (N_714,In_120,In_246);
and U715 (N_715,In_171,In_402);
or U716 (N_716,In_648,In_825);
and U717 (N_717,In_1391,In_1213);
nand U718 (N_718,In_620,In_827);
or U719 (N_719,In_17,In_516);
nor U720 (N_720,In_1401,In_1058);
nand U721 (N_721,In_1079,In_1165);
nand U722 (N_722,In_1485,In_1247);
or U723 (N_723,In_119,In_982);
and U724 (N_724,In_792,In_97);
xnor U725 (N_725,In_1085,In_1181);
or U726 (N_726,In_716,In_758);
or U727 (N_727,In_1035,In_1306);
nand U728 (N_728,In_1094,In_948);
xor U729 (N_729,In_320,In_545);
or U730 (N_730,In_1463,In_1054);
nor U731 (N_731,In_1346,In_229);
or U732 (N_732,In_1013,In_1459);
or U733 (N_733,In_335,In_883);
nor U734 (N_734,In_592,In_644);
nor U735 (N_735,In_759,In_530);
nor U736 (N_736,In_1317,In_1406);
nand U737 (N_737,In_59,In_211);
nand U738 (N_738,In_695,In_1496);
and U739 (N_739,In_1466,In_969);
nor U740 (N_740,In_637,In_714);
and U741 (N_741,In_938,In_1286);
xor U742 (N_742,In_1241,In_364);
nand U743 (N_743,In_1127,In_1488);
xor U744 (N_744,In_1280,In_985);
xnor U745 (N_745,In_1031,In_114);
xnor U746 (N_746,In_820,In_803);
nor U747 (N_747,In_1370,In_1057);
and U748 (N_748,In_1104,In_430);
nor U749 (N_749,In_605,In_719);
and U750 (N_750,In_1311,In_1017);
nor U751 (N_751,In_599,In_1412);
nand U752 (N_752,In_1069,In_462);
nor U753 (N_753,In_274,In_164);
and U754 (N_754,In_471,In_70);
xnor U755 (N_755,In_1481,In_160);
or U756 (N_756,In_76,In_1023);
and U757 (N_757,In_952,In_761);
or U758 (N_758,In_196,In_1316);
nand U759 (N_759,In_1070,In_1413);
or U760 (N_760,In_764,In_525);
xor U761 (N_761,In_660,In_1289);
nor U762 (N_762,In_52,In_357);
nor U763 (N_763,In_852,In_252);
and U764 (N_764,In_902,In_439);
nor U765 (N_765,In_681,In_379);
and U766 (N_766,In_781,In_829);
xor U767 (N_767,In_1459,In_1269);
xor U768 (N_768,In_610,In_1172);
nor U769 (N_769,In_463,In_1164);
xor U770 (N_770,In_1140,In_381);
or U771 (N_771,In_749,In_269);
nor U772 (N_772,In_366,In_1335);
or U773 (N_773,In_32,In_708);
nor U774 (N_774,In_332,In_110);
and U775 (N_775,In_521,In_1223);
and U776 (N_776,In_1443,In_1068);
xor U777 (N_777,In_1371,In_1013);
nand U778 (N_778,In_266,In_65);
or U779 (N_779,In_1379,In_1073);
or U780 (N_780,In_602,In_35);
nand U781 (N_781,In_1010,In_665);
xor U782 (N_782,In_1278,In_1332);
nor U783 (N_783,In_7,In_168);
and U784 (N_784,In_172,In_796);
and U785 (N_785,In_1059,In_664);
nand U786 (N_786,In_1042,In_660);
or U787 (N_787,In_649,In_1413);
xnor U788 (N_788,In_987,In_1129);
and U789 (N_789,In_1138,In_234);
xnor U790 (N_790,In_1257,In_933);
nand U791 (N_791,In_248,In_365);
or U792 (N_792,In_67,In_1008);
nor U793 (N_793,In_9,In_1251);
or U794 (N_794,In_1463,In_129);
xnor U795 (N_795,In_1392,In_3);
xor U796 (N_796,In_232,In_988);
or U797 (N_797,In_1169,In_48);
nor U798 (N_798,In_333,In_685);
and U799 (N_799,In_607,In_926);
xnor U800 (N_800,In_921,In_143);
nor U801 (N_801,In_745,In_1180);
nor U802 (N_802,In_219,In_781);
nand U803 (N_803,In_780,In_1428);
nor U804 (N_804,In_992,In_1364);
or U805 (N_805,In_979,In_342);
and U806 (N_806,In_1362,In_910);
nand U807 (N_807,In_817,In_570);
and U808 (N_808,In_1434,In_657);
nand U809 (N_809,In_1183,In_305);
nor U810 (N_810,In_1076,In_241);
and U811 (N_811,In_409,In_471);
and U812 (N_812,In_1137,In_1215);
and U813 (N_813,In_1279,In_970);
and U814 (N_814,In_401,In_595);
nor U815 (N_815,In_394,In_1057);
and U816 (N_816,In_1134,In_1375);
and U817 (N_817,In_239,In_362);
nor U818 (N_818,In_1448,In_853);
nor U819 (N_819,In_985,In_1140);
nand U820 (N_820,In_27,In_366);
and U821 (N_821,In_1030,In_1081);
nor U822 (N_822,In_873,In_1353);
nand U823 (N_823,In_1431,In_148);
nand U824 (N_824,In_1016,In_591);
nand U825 (N_825,In_793,In_936);
and U826 (N_826,In_1064,In_465);
xnor U827 (N_827,In_537,In_702);
and U828 (N_828,In_1388,In_1124);
and U829 (N_829,In_1249,In_498);
nor U830 (N_830,In_946,In_61);
xor U831 (N_831,In_47,In_812);
and U832 (N_832,In_1039,In_25);
or U833 (N_833,In_62,In_640);
or U834 (N_834,In_1477,In_738);
nor U835 (N_835,In_226,In_340);
nand U836 (N_836,In_125,In_386);
or U837 (N_837,In_116,In_1010);
xor U838 (N_838,In_910,In_1119);
xnor U839 (N_839,In_1360,In_555);
and U840 (N_840,In_340,In_189);
and U841 (N_841,In_661,In_543);
xnor U842 (N_842,In_633,In_104);
or U843 (N_843,In_22,In_114);
and U844 (N_844,In_503,In_29);
nand U845 (N_845,In_1246,In_457);
xor U846 (N_846,In_570,In_1308);
nand U847 (N_847,In_807,In_271);
nand U848 (N_848,In_965,In_681);
nor U849 (N_849,In_1082,In_1114);
and U850 (N_850,In_122,In_309);
nor U851 (N_851,In_871,In_792);
xor U852 (N_852,In_1211,In_184);
nand U853 (N_853,In_1102,In_263);
and U854 (N_854,In_357,In_386);
or U855 (N_855,In_1378,In_47);
xnor U856 (N_856,In_960,In_1237);
and U857 (N_857,In_167,In_215);
nor U858 (N_858,In_444,In_660);
nand U859 (N_859,In_1353,In_373);
nand U860 (N_860,In_482,In_159);
nand U861 (N_861,In_1366,In_950);
nor U862 (N_862,In_967,In_1404);
and U863 (N_863,In_338,In_9);
or U864 (N_864,In_784,In_1175);
nand U865 (N_865,In_1370,In_1284);
and U866 (N_866,In_308,In_475);
or U867 (N_867,In_353,In_685);
xor U868 (N_868,In_707,In_991);
and U869 (N_869,In_297,In_228);
nor U870 (N_870,In_215,In_589);
or U871 (N_871,In_126,In_567);
nor U872 (N_872,In_75,In_505);
xnor U873 (N_873,In_752,In_763);
and U874 (N_874,In_461,In_56);
nor U875 (N_875,In_1359,In_34);
nand U876 (N_876,In_9,In_1481);
nor U877 (N_877,In_721,In_101);
xnor U878 (N_878,In_661,In_1021);
nand U879 (N_879,In_1172,In_628);
xnor U880 (N_880,In_1137,In_103);
and U881 (N_881,In_611,In_562);
and U882 (N_882,In_882,In_831);
xor U883 (N_883,In_921,In_137);
and U884 (N_884,In_1243,In_1296);
nor U885 (N_885,In_740,In_837);
or U886 (N_886,In_754,In_729);
xnor U887 (N_887,In_646,In_148);
or U888 (N_888,In_1390,In_1469);
and U889 (N_889,In_350,In_921);
and U890 (N_890,In_1383,In_765);
nor U891 (N_891,In_1458,In_861);
nor U892 (N_892,In_1250,In_122);
and U893 (N_893,In_431,In_1437);
xnor U894 (N_894,In_1176,In_151);
nor U895 (N_895,In_1238,In_201);
xor U896 (N_896,In_906,In_1298);
nor U897 (N_897,In_985,In_66);
xor U898 (N_898,In_100,In_510);
nand U899 (N_899,In_409,In_141);
nor U900 (N_900,In_176,In_807);
or U901 (N_901,In_501,In_246);
or U902 (N_902,In_567,In_1184);
nor U903 (N_903,In_532,In_807);
nor U904 (N_904,In_1443,In_1241);
nor U905 (N_905,In_1362,In_740);
and U906 (N_906,In_1088,In_191);
nand U907 (N_907,In_132,In_482);
nand U908 (N_908,In_1138,In_101);
nor U909 (N_909,In_861,In_1141);
xor U910 (N_910,In_1309,In_480);
xnor U911 (N_911,In_322,In_734);
nor U912 (N_912,In_723,In_626);
nand U913 (N_913,In_687,In_926);
or U914 (N_914,In_1338,In_802);
xnor U915 (N_915,In_1253,In_618);
nor U916 (N_916,In_395,In_251);
or U917 (N_917,In_1322,In_698);
nand U918 (N_918,In_1145,In_337);
and U919 (N_919,In_842,In_787);
nor U920 (N_920,In_876,In_601);
or U921 (N_921,In_1241,In_313);
and U922 (N_922,In_380,In_1010);
nor U923 (N_923,In_738,In_841);
or U924 (N_924,In_1174,In_1097);
nand U925 (N_925,In_1405,In_1280);
or U926 (N_926,In_20,In_826);
nand U927 (N_927,In_912,In_1339);
and U928 (N_928,In_709,In_545);
nand U929 (N_929,In_1116,In_1379);
nand U930 (N_930,In_992,In_644);
nor U931 (N_931,In_122,In_998);
and U932 (N_932,In_924,In_625);
nand U933 (N_933,In_311,In_907);
xnor U934 (N_934,In_367,In_387);
and U935 (N_935,In_1202,In_563);
nor U936 (N_936,In_992,In_1008);
xor U937 (N_937,In_1389,In_404);
or U938 (N_938,In_1057,In_513);
xnor U939 (N_939,In_722,In_250);
and U940 (N_940,In_32,In_1470);
or U941 (N_941,In_976,In_512);
or U942 (N_942,In_1141,In_1225);
and U943 (N_943,In_219,In_914);
nand U944 (N_944,In_58,In_998);
nor U945 (N_945,In_940,In_1466);
nand U946 (N_946,In_836,In_1322);
or U947 (N_947,In_416,In_706);
and U948 (N_948,In_600,In_809);
nand U949 (N_949,In_969,In_740);
or U950 (N_950,In_361,In_155);
nand U951 (N_951,In_1308,In_559);
xnor U952 (N_952,In_546,In_709);
nor U953 (N_953,In_1156,In_650);
or U954 (N_954,In_262,In_747);
nor U955 (N_955,In_581,In_1397);
xor U956 (N_956,In_1028,In_816);
or U957 (N_957,In_1474,In_673);
or U958 (N_958,In_126,In_1197);
nor U959 (N_959,In_1136,In_332);
nor U960 (N_960,In_889,In_356);
nor U961 (N_961,In_448,In_137);
xnor U962 (N_962,In_890,In_1252);
nor U963 (N_963,In_1437,In_442);
and U964 (N_964,In_515,In_429);
and U965 (N_965,In_45,In_940);
and U966 (N_966,In_611,In_84);
or U967 (N_967,In_720,In_1077);
or U968 (N_968,In_336,In_1170);
and U969 (N_969,In_1341,In_31);
xor U970 (N_970,In_923,In_85);
and U971 (N_971,In_578,In_933);
or U972 (N_972,In_1136,In_1088);
or U973 (N_973,In_1181,In_1007);
nand U974 (N_974,In_1182,In_455);
xnor U975 (N_975,In_853,In_1460);
or U976 (N_976,In_1169,In_1324);
or U977 (N_977,In_910,In_796);
nand U978 (N_978,In_819,In_859);
and U979 (N_979,In_844,In_1119);
nand U980 (N_980,In_1436,In_236);
nor U981 (N_981,In_1374,In_442);
or U982 (N_982,In_985,In_967);
nor U983 (N_983,In_47,In_475);
xor U984 (N_984,In_395,In_796);
nor U985 (N_985,In_623,In_86);
and U986 (N_986,In_977,In_713);
nand U987 (N_987,In_463,In_960);
or U988 (N_988,In_772,In_661);
nand U989 (N_989,In_47,In_159);
xnor U990 (N_990,In_755,In_673);
nand U991 (N_991,In_1289,In_645);
nor U992 (N_992,In_603,In_113);
xnor U993 (N_993,In_1094,In_445);
or U994 (N_994,In_1434,In_1339);
xor U995 (N_995,In_1460,In_801);
nand U996 (N_996,In_1332,In_198);
nand U997 (N_997,In_202,In_1313);
nand U998 (N_998,In_85,In_269);
and U999 (N_999,In_217,In_914);
xor U1000 (N_1000,In_706,In_868);
and U1001 (N_1001,In_892,In_528);
nand U1002 (N_1002,In_1421,In_504);
or U1003 (N_1003,In_1263,In_128);
nor U1004 (N_1004,In_124,In_110);
nor U1005 (N_1005,In_950,In_534);
xnor U1006 (N_1006,In_234,In_1010);
nor U1007 (N_1007,In_1058,In_720);
and U1008 (N_1008,In_1001,In_1350);
nor U1009 (N_1009,In_1484,In_83);
nor U1010 (N_1010,In_809,In_1447);
xnor U1011 (N_1011,In_953,In_1294);
xor U1012 (N_1012,In_465,In_977);
nand U1013 (N_1013,In_1065,In_763);
xor U1014 (N_1014,In_1120,In_321);
nor U1015 (N_1015,In_1203,In_635);
xnor U1016 (N_1016,In_1245,In_295);
xor U1017 (N_1017,In_628,In_303);
nand U1018 (N_1018,In_1023,In_1131);
nand U1019 (N_1019,In_1067,In_217);
or U1020 (N_1020,In_489,In_1256);
xnor U1021 (N_1021,In_987,In_1023);
and U1022 (N_1022,In_1367,In_143);
nand U1023 (N_1023,In_535,In_81);
and U1024 (N_1024,In_135,In_1199);
nand U1025 (N_1025,In_1288,In_1205);
xnor U1026 (N_1026,In_369,In_443);
and U1027 (N_1027,In_301,In_677);
nor U1028 (N_1028,In_1044,In_88);
and U1029 (N_1029,In_1454,In_307);
or U1030 (N_1030,In_511,In_142);
nand U1031 (N_1031,In_725,In_783);
or U1032 (N_1032,In_410,In_292);
nor U1033 (N_1033,In_1084,In_548);
or U1034 (N_1034,In_499,In_996);
or U1035 (N_1035,In_534,In_1414);
or U1036 (N_1036,In_1329,In_767);
nand U1037 (N_1037,In_562,In_205);
nand U1038 (N_1038,In_281,In_483);
nand U1039 (N_1039,In_1411,In_505);
or U1040 (N_1040,In_1225,In_229);
xor U1041 (N_1041,In_789,In_983);
and U1042 (N_1042,In_258,In_1476);
and U1043 (N_1043,In_582,In_568);
xor U1044 (N_1044,In_984,In_357);
nand U1045 (N_1045,In_806,In_1173);
nand U1046 (N_1046,In_1490,In_1043);
or U1047 (N_1047,In_389,In_496);
or U1048 (N_1048,In_257,In_1237);
or U1049 (N_1049,In_936,In_1022);
nand U1050 (N_1050,In_130,In_972);
nor U1051 (N_1051,In_1167,In_401);
and U1052 (N_1052,In_290,In_650);
nor U1053 (N_1053,In_1123,In_1170);
nand U1054 (N_1054,In_421,In_716);
nor U1055 (N_1055,In_534,In_1128);
and U1056 (N_1056,In_975,In_1042);
nor U1057 (N_1057,In_67,In_1461);
or U1058 (N_1058,In_1286,In_1243);
and U1059 (N_1059,In_253,In_522);
nor U1060 (N_1060,In_1172,In_182);
and U1061 (N_1061,In_940,In_1389);
and U1062 (N_1062,In_978,In_915);
or U1063 (N_1063,In_1459,In_1249);
nand U1064 (N_1064,In_172,In_268);
or U1065 (N_1065,In_248,In_1091);
xnor U1066 (N_1066,In_1035,In_835);
nor U1067 (N_1067,In_1232,In_576);
nor U1068 (N_1068,In_518,In_636);
nand U1069 (N_1069,In_1363,In_863);
xnor U1070 (N_1070,In_412,In_789);
nand U1071 (N_1071,In_190,In_759);
nor U1072 (N_1072,In_1224,In_492);
or U1073 (N_1073,In_379,In_664);
xnor U1074 (N_1074,In_980,In_1275);
nor U1075 (N_1075,In_420,In_564);
xor U1076 (N_1076,In_114,In_1172);
nor U1077 (N_1077,In_1411,In_1360);
nand U1078 (N_1078,In_1193,In_486);
nor U1079 (N_1079,In_244,In_1474);
nand U1080 (N_1080,In_140,In_933);
nand U1081 (N_1081,In_272,In_590);
or U1082 (N_1082,In_1418,In_386);
xnor U1083 (N_1083,In_396,In_518);
and U1084 (N_1084,In_261,In_270);
xor U1085 (N_1085,In_1031,In_67);
xnor U1086 (N_1086,In_1001,In_277);
or U1087 (N_1087,In_45,In_1037);
and U1088 (N_1088,In_1446,In_651);
xnor U1089 (N_1089,In_413,In_341);
nand U1090 (N_1090,In_533,In_1434);
xor U1091 (N_1091,In_885,In_776);
or U1092 (N_1092,In_1432,In_629);
nor U1093 (N_1093,In_141,In_1267);
nand U1094 (N_1094,In_1274,In_411);
and U1095 (N_1095,In_71,In_284);
nor U1096 (N_1096,In_883,In_478);
or U1097 (N_1097,In_475,In_745);
and U1098 (N_1098,In_1305,In_1378);
nand U1099 (N_1099,In_860,In_1264);
xnor U1100 (N_1100,In_801,In_689);
nor U1101 (N_1101,In_853,In_58);
and U1102 (N_1102,In_821,In_344);
xor U1103 (N_1103,In_639,In_120);
or U1104 (N_1104,In_1413,In_1293);
nand U1105 (N_1105,In_959,In_1025);
nor U1106 (N_1106,In_461,In_495);
or U1107 (N_1107,In_1166,In_313);
nand U1108 (N_1108,In_833,In_498);
nand U1109 (N_1109,In_1441,In_1101);
or U1110 (N_1110,In_1221,In_1488);
nor U1111 (N_1111,In_988,In_886);
nor U1112 (N_1112,In_1112,In_895);
and U1113 (N_1113,In_1019,In_494);
or U1114 (N_1114,In_246,In_1307);
and U1115 (N_1115,In_946,In_51);
nor U1116 (N_1116,In_777,In_89);
nor U1117 (N_1117,In_309,In_799);
nand U1118 (N_1118,In_1074,In_239);
nand U1119 (N_1119,In_464,In_1308);
nand U1120 (N_1120,In_618,In_270);
and U1121 (N_1121,In_585,In_830);
and U1122 (N_1122,In_279,In_965);
and U1123 (N_1123,In_691,In_1138);
nand U1124 (N_1124,In_938,In_110);
xor U1125 (N_1125,In_1015,In_944);
or U1126 (N_1126,In_641,In_1362);
nor U1127 (N_1127,In_228,In_224);
nor U1128 (N_1128,In_1181,In_365);
nor U1129 (N_1129,In_1335,In_1062);
nor U1130 (N_1130,In_144,In_1190);
and U1131 (N_1131,In_1242,In_402);
and U1132 (N_1132,In_645,In_997);
and U1133 (N_1133,In_240,In_847);
xor U1134 (N_1134,In_1392,In_1195);
or U1135 (N_1135,In_63,In_599);
xor U1136 (N_1136,In_1416,In_84);
nand U1137 (N_1137,In_1147,In_592);
or U1138 (N_1138,In_902,In_1145);
or U1139 (N_1139,In_1421,In_291);
nand U1140 (N_1140,In_1376,In_105);
and U1141 (N_1141,In_64,In_1214);
and U1142 (N_1142,In_233,In_293);
nor U1143 (N_1143,In_733,In_1432);
nand U1144 (N_1144,In_1279,In_253);
xnor U1145 (N_1145,In_1421,In_1488);
nor U1146 (N_1146,In_635,In_1384);
xnor U1147 (N_1147,In_22,In_215);
nor U1148 (N_1148,In_48,In_399);
nand U1149 (N_1149,In_1462,In_1066);
xor U1150 (N_1150,In_850,In_897);
and U1151 (N_1151,In_246,In_1038);
and U1152 (N_1152,In_643,In_1181);
nand U1153 (N_1153,In_481,In_545);
and U1154 (N_1154,In_829,In_100);
nand U1155 (N_1155,In_896,In_319);
or U1156 (N_1156,In_1138,In_813);
xor U1157 (N_1157,In_1218,In_278);
or U1158 (N_1158,In_460,In_1325);
or U1159 (N_1159,In_117,In_1023);
and U1160 (N_1160,In_688,In_887);
and U1161 (N_1161,In_737,In_905);
and U1162 (N_1162,In_980,In_444);
nand U1163 (N_1163,In_1342,In_1333);
nor U1164 (N_1164,In_724,In_1467);
nand U1165 (N_1165,In_1039,In_910);
xor U1166 (N_1166,In_836,In_893);
or U1167 (N_1167,In_646,In_540);
and U1168 (N_1168,In_1306,In_372);
xnor U1169 (N_1169,In_41,In_715);
and U1170 (N_1170,In_768,In_1160);
or U1171 (N_1171,In_851,In_1011);
xnor U1172 (N_1172,In_833,In_296);
or U1173 (N_1173,In_1076,In_544);
xnor U1174 (N_1174,In_1051,In_807);
or U1175 (N_1175,In_55,In_529);
nor U1176 (N_1176,In_1010,In_564);
and U1177 (N_1177,In_486,In_438);
nand U1178 (N_1178,In_696,In_10);
or U1179 (N_1179,In_452,In_870);
nor U1180 (N_1180,In_821,In_589);
and U1181 (N_1181,In_1096,In_35);
xnor U1182 (N_1182,In_1008,In_910);
or U1183 (N_1183,In_208,In_946);
xor U1184 (N_1184,In_1285,In_543);
or U1185 (N_1185,In_346,In_129);
and U1186 (N_1186,In_391,In_511);
and U1187 (N_1187,In_1304,In_1374);
nand U1188 (N_1188,In_579,In_857);
xnor U1189 (N_1189,In_1171,In_788);
xor U1190 (N_1190,In_1108,In_241);
or U1191 (N_1191,In_628,In_519);
and U1192 (N_1192,In_759,In_309);
xor U1193 (N_1193,In_811,In_1440);
nand U1194 (N_1194,In_678,In_707);
or U1195 (N_1195,In_825,In_752);
or U1196 (N_1196,In_343,In_1050);
and U1197 (N_1197,In_665,In_691);
nor U1198 (N_1198,In_886,In_1327);
nor U1199 (N_1199,In_28,In_1098);
nand U1200 (N_1200,In_1326,In_588);
xnor U1201 (N_1201,In_270,In_1277);
nand U1202 (N_1202,In_238,In_456);
and U1203 (N_1203,In_559,In_1158);
nor U1204 (N_1204,In_883,In_533);
and U1205 (N_1205,In_731,In_310);
nor U1206 (N_1206,In_75,In_915);
nand U1207 (N_1207,In_1165,In_864);
xnor U1208 (N_1208,In_93,In_168);
xor U1209 (N_1209,In_1322,In_62);
or U1210 (N_1210,In_331,In_339);
nor U1211 (N_1211,In_1442,In_504);
nor U1212 (N_1212,In_1136,In_19);
or U1213 (N_1213,In_90,In_714);
nor U1214 (N_1214,In_950,In_1142);
xnor U1215 (N_1215,In_502,In_1469);
nor U1216 (N_1216,In_1236,In_1355);
or U1217 (N_1217,In_1216,In_530);
and U1218 (N_1218,In_121,In_1072);
nor U1219 (N_1219,In_1045,In_536);
nor U1220 (N_1220,In_41,In_349);
xor U1221 (N_1221,In_116,In_1293);
xor U1222 (N_1222,In_784,In_1485);
or U1223 (N_1223,In_1470,In_480);
or U1224 (N_1224,In_689,In_979);
nor U1225 (N_1225,In_345,In_928);
or U1226 (N_1226,In_173,In_680);
nand U1227 (N_1227,In_1192,In_8);
nand U1228 (N_1228,In_725,In_134);
and U1229 (N_1229,In_1001,In_132);
xor U1230 (N_1230,In_7,In_476);
or U1231 (N_1231,In_394,In_356);
xnor U1232 (N_1232,In_1271,In_608);
nand U1233 (N_1233,In_644,In_1070);
nand U1234 (N_1234,In_1110,In_866);
xnor U1235 (N_1235,In_1329,In_783);
nor U1236 (N_1236,In_90,In_458);
or U1237 (N_1237,In_1419,In_1174);
and U1238 (N_1238,In_1221,In_1317);
xnor U1239 (N_1239,In_148,In_852);
nand U1240 (N_1240,In_20,In_985);
and U1241 (N_1241,In_1127,In_325);
nor U1242 (N_1242,In_522,In_1056);
or U1243 (N_1243,In_1457,In_993);
nor U1244 (N_1244,In_1029,In_1179);
nand U1245 (N_1245,In_226,In_30);
xor U1246 (N_1246,In_472,In_43);
nor U1247 (N_1247,In_633,In_852);
xnor U1248 (N_1248,In_624,In_1229);
or U1249 (N_1249,In_1280,In_476);
or U1250 (N_1250,In_145,In_858);
or U1251 (N_1251,In_824,In_1055);
and U1252 (N_1252,In_659,In_284);
nor U1253 (N_1253,In_315,In_1037);
or U1254 (N_1254,In_228,In_954);
and U1255 (N_1255,In_1499,In_770);
and U1256 (N_1256,In_882,In_249);
xor U1257 (N_1257,In_655,In_814);
and U1258 (N_1258,In_643,In_98);
nand U1259 (N_1259,In_1301,In_67);
xnor U1260 (N_1260,In_502,In_547);
nor U1261 (N_1261,In_1260,In_674);
xnor U1262 (N_1262,In_303,In_376);
nand U1263 (N_1263,In_828,In_879);
and U1264 (N_1264,In_331,In_1437);
or U1265 (N_1265,In_486,In_224);
and U1266 (N_1266,In_1455,In_598);
nor U1267 (N_1267,In_561,In_1238);
nor U1268 (N_1268,In_912,In_758);
xor U1269 (N_1269,In_987,In_1337);
and U1270 (N_1270,In_914,In_166);
and U1271 (N_1271,In_723,In_1012);
nand U1272 (N_1272,In_911,In_1182);
and U1273 (N_1273,In_1122,In_1454);
nand U1274 (N_1274,In_396,In_322);
nand U1275 (N_1275,In_513,In_1480);
nand U1276 (N_1276,In_1487,In_1252);
xor U1277 (N_1277,In_307,In_916);
and U1278 (N_1278,In_692,In_66);
or U1279 (N_1279,In_1350,In_845);
or U1280 (N_1280,In_450,In_1358);
xor U1281 (N_1281,In_59,In_1272);
nor U1282 (N_1282,In_946,In_598);
and U1283 (N_1283,In_911,In_349);
and U1284 (N_1284,In_423,In_597);
nand U1285 (N_1285,In_418,In_989);
and U1286 (N_1286,In_372,In_943);
xnor U1287 (N_1287,In_609,In_454);
and U1288 (N_1288,In_1103,In_603);
or U1289 (N_1289,In_61,In_995);
nor U1290 (N_1290,In_808,In_1038);
xor U1291 (N_1291,In_76,In_499);
xnor U1292 (N_1292,In_1369,In_917);
and U1293 (N_1293,In_1012,In_1104);
nor U1294 (N_1294,In_374,In_452);
xnor U1295 (N_1295,In_1048,In_511);
nor U1296 (N_1296,In_1340,In_1277);
and U1297 (N_1297,In_134,In_990);
nand U1298 (N_1298,In_256,In_795);
and U1299 (N_1299,In_1226,In_733);
and U1300 (N_1300,In_729,In_2);
xnor U1301 (N_1301,In_1383,In_236);
nor U1302 (N_1302,In_740,In_993);
xnor U1303 (N_1303,In_845,In_626);
xor U1304 (N_1304,In_1486,In_874);
nor U1305 (N_1305,In_1186,In_434);
nand U1306 (N_1306,In_1272,In_1033);
xnor U1307 (N_1307,In_1487,In_597);
nand U1308 (N_1308,In_1193,In_339);
nand U1309 (N_1309,In_117,In_176);
or U1310 (N_1310,In_1310,In_1349);
nor U1311 (N_1311,In_836,In_765);
nor U1312 (N_1312,In_1193,In_284);
xor U1313 (N_1313,In_691,In_303);
xnor U1314 (N_1314,In_1116,In_81);
xnor U1315 (N_1315,In_250,In_304);
nor U1316 (N_1316,In_1018,In_378);
and U1317 (N_1317,In_879,In_1231);
nor U1318 (N_1318,In_1435,In_80);
nor U1319 (N_1319,In_759,In_1105);
or U1320 (N_1320,In_628,In_1200);
xnor U1321 (N_1321,In_1193,In_357);
nand U1322 (N_1322,In_475,In_229);
or U1323 (N_1323,In_13,In_890);
xor U1324 (N_1324,In_237,In_1405);
and U1325 (N_1325,In_1298,In_1362);
nor U1326 (N_1326,In_276,In_1358);
xor U1327 (N_1327,In_588,In_142);
or U1328 (N_1328,In_1209,In_1085);
and U1329 (N_1329,In_595,In_1018);
nand U1330 (N_1330,In_5,In_95);
xor U1331 (N_1331,In_530,In_1075);
xor U1332 (N_1332,In_1244,In_12);
nand U1333 (N_1333,In_674,In_444);
nand U1334 (N_1334,In_857,In_1);
nor U1335 (N_1335,In_838,In_1066);
or U1336 (N_1336,In_652,In_736);
xnor U1337 (N_1337,In_1019,In_1136);
nor U1338 (N_1338,In_45,In_661);
or U1339 (N_1339,In_582,In_1078);
xnor U1340 (N_1340,In_242,In_1448);
or U1341 (N_1341,In_472,In_1298);
and U1342 (N_1342,In_189,In_1216);
and U1343 (N_1343,In_856,In_917);
or U1344 (N_1344,In_1293,In_60);
nor U1345 (N_1345,In_903,In_40);
nor U1346 (N_1346,In_105,In_78);
or U1347 (N_1347,In_597,In_885);
nand U1348 (N_1348,In_849,In_439);
and U1349 (N_1349,In_1027,In_2);
or U1350 (N_1350,In_394,In_1103);
nand U1351 (N_1351,In_1252,In_1306);
nor U1352 (N_1352,In_381,In_979);
nor U1353 (N_1353,In_42,In_1095);
xnor U1354 (N_1354,In_728,In_1391);
nand U1355 (N_1355,In_342,In_42);
nand U1356 (N_1356,In_1238,In_519);
or U1357 (N_1357,In_85,In_1166);
nor U1358 (N_1358,In_896,In_631);
xor U1359 (N_1359,In_782,In_417);
and U1360 (N_1360,In_58,In_651);
and U1361 (N_1361,In_411,In_254);
and U1362 (N_1362,In_142,In_230);
or U1363 (N_1363,In_595,In_844);
and U1364 (N_1364,In_988,In_557);
and U1365 (N_1365,In_832,In_1100);
nor U1366 (N_1366,In_420,In_932);
nand U1367 (N_1367,In_1366,In_846);
nand U1368 (N_1368,In_1273,In_1479);
xnor U1369 (N_1369,In_574,In_669);
and U1370 (N_1370,In_253,In_425);
nor U1371 (N_1371,In_949,In_1179);
nor U1372 (N_1372,In_265,In_159);
or U1373 (N_1373,In_82,In_1334);
and U1374 (N_1374,In_910,In_1113);
xor U1375 (N_1375,In_1208,In_266);
nor U1376 (N_1376,In_91,In_1121);
xnor U1377 (N_1377,In_990,In_427);
xnor U1378 (N_1378,In_281,In_562);
xor U1379 (N_1379,In_420,In_1180);
or U1380 (N_1380,In_1169,In_1484);
nand U1381 (N_1381,In_415,In_723);
and U1382 (N_1382,In_246,In_732);
nand U1383 (N_1383,In_1086,In_188);
xnor U1384 (N_1384,In_415,In_497);
and U1385 (N_1385,In_358,In_864);
nand U1386 (N_1386,In_797,In_987);
or U1387 (N_1387,In_458,In_841);
and U1388 (N_1388,In_891,In_885);
or U1389 (N_1389,In_606,In_239);
and U1390 (N_1390,In_1372,In_1326);
or U1391 (N_1391,In_1169,In_1420);
nor U1392 (N_1392,In_718,In_914);
nor U1393 (N_1393,In_416,In_200);
and U1394 (N_1394,In_285,In_1326);
and U1395 (N_1395,In_856,In_274);
xnor U1396 (N_1396,In_706,In_71);
xor U1397 (N_1397,In_1392,In_1371);
xor U1398 (N_1398,In_719,In_1407);
nor U1399 (N_1399,In_246,In_58);
or U1400 (N_1400,In_1345,In_672);
xnor U1401 (N_1401,In_861,In_1131);
xnor U1402 (N_1402,In_624,In_1023);
xnor U1403 (N_1403,In_444,In_765);
nand U1404 (N_1404,In_988,In_828);
nor U1405 (N_1405,In_685,In_938);
and U1406 (N_1406,In_61,In_1275);
nand U1407 (N_1407,In_1160,In_1374);
nand U1408 (N_1408,In_402,In_278);
or U1409 (N_1409,In_1157,In_1468);
nand U1410 (N_1410,In_261,In_1066);
xnor U1411 (N_1411,In_818,In_552);
nand U1412 (N_1412,In_22,In_1201);
nor U1413 (N_1413,In_341,In_1499);
nor U1414 (N_1414,In_810,In_1121);
xor U1415 (N_1415,In_325,In_337);
or U1416 (N_1416,In_758,In_173);
or U1417 (N_1417,In_821,In_1253);
or U1418 (N_1418,In_739,In_86);
and U1419 (N_1419,In_357,In_681);
or U1420 (N_1420,In_199,In_845);
and U1421 (N_1421,In_1069,In_1020);
and U1422 (N_1422,In_1207,In_928);
or U1423 (N_1423,In_846,In_653);
nand U1424 (N_1424,In_1207,In_1094);
nand U1425 (N_1425,In_459,In_358);
and U1426 (N_1426,In_22,In_827);
nand U1427 (N_1427,In_1229,In_898);
nand U1428 (N_1428,In_1170,In_109);
nor U1429 (N_1429,In_1167,In_1139);
nand U1430 (N_1430,In_1393,In_532);
nand U1431 (N_1431,In_1337,In_434);
and U1432 (N_1432,In_786,In_519);
and U1433 (N_1433,In_1375,In_133);
and U1434 (N_1434,In_315,In_1242);
nand U1435 (N_1435,In_626,In_608);
nor U1436 (N_1436,In_470,In_72);
nor U1437 (N_1437,In_1257,In_1013);
xnor U1438 (N_1438,In_1024,In_445);
nor U1439 (N_1439,In_1044,In_1273);
or U1440 (N_1440,In_982,In_70);
nand U1441 (N_1441,In_1010,In_569);
nor U1442 (N_1442,In_772,In_431);
and U1443 (N_1443,In_1138,In_977);
or U1444 (N_1444,In_68,In_1310);
xor U1445 (N_1445,In_182,In_61);
and U1446 (N_1446,In_376,In_664);
and U1447 (N_1447,In_229,In_892);
and U1448 (N_1448,In_435,In_1018);
nand U1449 (N_1449,In_181,In_893);
and U1450 (N_1450,In_336,In_872);
or U1451 (N_1451,In_947,In_1142);
or U1452 (N_1452,In_1197,In_1062);
nand U1453 (N_1453,In_452,In_397);
nand U1454 (N_1454,In_1486,In_953);
xor U1455 (N_1455,In_393,In_725);
or U1456 (N_1456,In_952,In_615);
nand U1457 (N_1457,In_626,In_1194);
xor U1458 (N_1458,In_481,In_646);
nand U1459 (N_1459,In_1453,In_249);
nor U1460 (N_1460,In_1490,In_137);
and U1461 (N_1461,In_878,In_674);
or U1462 (N_1462,In_544,In_1482);
or U1463 (N_1463,In_1032,In_651);
nor U1464 (N_1464,In_776,In_1367);
xor U1465 (N_1465,In_525,In_861);
xor U1466 (N_1466,In_574,In_1464);
or U1467 (N_1467,In_198,In_1092);
or U1468 (N_1468,In_208,In_532);
or U1469 (N_1469,In_400,In_183);
or U1470 (N_1470,In_1264,In_340);
nor U1471 (N_1471,In_502,In_902);
nand U1472 (N_1472,In_707,In_398);
xnor U1473 (N_1473,In_1209,In_228);
nor U1474 (N_1474,In_161,In_283);
and U1475 (N_1475,In_364,In_902);
nor U1476 (N_1476,In_688,In_752);
or U1477 (N_1477,In_1259,In_713);
and U1478 (N_1478,In_1474,In_1250);
and U1479 (N_1479,In_1410,In_647);
nor U1480 (N_1480,In_1358,In_1216);
or U1481 (N_1481,In_556,In_191);
xor U1482 (N_1482,In_288,In_1051);
nand U1483 (N_1483,In_1144,In_561);
and U1484 (N_1484,In_1365,In_176);
nor U1485 (N_1485,In_469,In_1133);
nand U1486 (N_1486,In_1301,In_62);
xor U1487 (N_1487,In_1120,In_278);
and U1488 (N_1488,In_894,In_504);
and U1489 (N_1489,In_848,In_589);
nand U1490 (N_1490,In_1130,In_1379);
nor U1491 (N_1491,In_420,In_1303);
xor U1492 (N_1492,In_1167,In_371);
nor U1493 (N_1493,In_255,In_606);
nand U1494 (N_1494,In_334,In_955);
nand U1495 (N_1495,In_326,In_828);
or U1496 (N_1496,In_87,In_1352);
nand U1497 (N_1497,In_928,In_1209);
or U1498 (N_1498,In_1078,In_1399);
xor U1499 (N_1499,In_326,In_867);
or U1500 (N_1500,In_1295,In_1005);
and U1501 (N_1501,In_852,In_6);
xor U1502 (N_1502,In_578,In_832);
xor U1503 (N_1503,In_927,In_320);
nand U1504 (N_1504,In_657,In_128);
and U1505 (N_1505,In_1476,In_900);
xor U1506 (N_1506,In_693,In_612);
xnor U1507 (N_1507,In_822,In_67);
xnor U1508 (N_1508,In_399,In_1231);
nand U1509 (N_1509,In_1441,In_262);
and U1510 (N_1510,In_1490,In_141);
xor U1511 (N_1511,In_610,In_402);
and U1512 (N_1512,In_445,In_1058);
nor U1513 (N_1513,In_1198,In_75);
nand U1514 (N_1514,In_820,In_1424);
nand U1515 (N_1515,In_168,In_338);
and U1516 (N_1516,In_982,In_849);
and U1517 (N_1517,In_511,In_1063);
xor U1518 (N_1518,In_736,In_646);
or U1519 (N_1519,In_270,In_1065);
and U1520 (N_1520,In_1167,In_380);
nor U1521 (N_1521,In_1112,In_320);
nor U1522 (N_1522,In_759,In_323);
nand U1523 (N_1523,In_983,In_1324);
nor U1524 (N_1524,In_583,In_711);
nand U1525 (N_1525,In_202,In_1302);
nand U1526 (N_1526,In_638,In_898);
nand U1527 (N_1527,In_130,In_272);
xnor U1528 (N_1528,In_84,In_832);
and U1529 (N_1529,In_134,In_595);
nor U1530 (N_1530,In_1119,In_1250);
xnor U1531 (N_1531,In_1108,In_504);
or U1532 (N_1532,In_452,In_935);
xor U1533 (N_1533,In_142,In_240);
xor U1534 (N_1534,In_971,In_1015);
nand U1535 (N_1535,In_1206,In_396);
nor U1536 (N_1536,In_217,In_1224);
and U1537 (N_1537,In_578,In_1388);
nor U1538 (N_1538,In_795,In_164);
nand U1539 (N_1539,In_1044,In_794);
nor U1540 (N_1540,In_2,In_285);
nand U1541 (N_1541,In_222,In_1361);
nor U1542 (N_1542,In_632,In_432);
or U1543 (N_1543,In_1006,In_814);
or U1544 (N_1544,In_809,In_6);
and U1545 (N_1545,In_1258,In_933);
and U1546 (N_1546,In_891,In_526);
xnor U1547 (N_1547,In_1263,In_844);
xnor U1548 (N_1548,In_1035,In_393);
and U1549 (N_1549,In_593,In_792);
xor U1550 (N_1550,In_358,In_365);
nand U1551 (N_1551,In_675,In_461);
or U1552 (N_1552,In_988,In_613);
xor U1553 (N_1553,In_19,In_460);
xnor U1554 (N_1554,In_870,In_961);
nor U1555 (N_1555,In_1306,In_1352);
nand U1556 (N_1556,In_146,In_718);
and U1557 (N_1557,In_188,In_480);
nand U1558 (N_1558,In_732,In_548);
or U1559 (N_1559,In_1259,In_1312);
or U1560 (N_1560,In_254,In_442);
xor U1561 (N_1561,In_604,In_299);
or U1562 (N_1562,In_862,In_154);
nor U1563 (N_1563,In_1353,In_964);
xor U1564 (N_1564,In_858,In_1352);
or U1565 (N_1565,In_729,In_1447);
nand U1566 (N_1566,In_1454,In_1377);
or U1567 (N_1567,In_1408,In_116);
xnor U1568 (N_1568,In_1087,In_55);
nor U1569 (N_1569,In_1293,In_703);
xnor U1570 (N_1570,In_1305,In_1254);
and U1571 (N_1571,In_1215,In_953);
xor U1572 (N_1572,In_1135,In_699);
nand U1573 (N_1573,In_629,In_970);
xor U1574 (N_1574,In_719,In_1113);
nand U1575 (N_1575,In_897,In_857);
or U1576 (N_1576,In_791,In_1274);
nor U1577 (N_1577,In_202,In_839);
or U1578 (N_1578,In_1266,In_191);
xnor U1579 (N_1579,In_195,In_621);
nor U1580 (N_1580,In_1095,In_179);
xor U1581 (N_1581,In_156,In_1225);
xnor U1582 (N_1582,In_1402,In_1008);
and U1583 (N_1583,In_772,In_924);
or U1584 (N_1584,In_1195,In_1046);
nor U1585 (N_1585,In_228,In_629);
or U1586 (N_1586,In_262,In_23);
nor U1587 (N_1587,In_328,In_688);
and U1588 (N_1588,In_1200,In_1221);
nor U1589 (N_1589,In_1206,In_928);
nand U1590 (N_1590,In_313,In_149);
xnor U1591 (N_1591,In_1437,In_946);
or U1592 (N_1592,In_423,In_881);
nor U1593 (N_1593,In_584,In_728);
or U1594 (N_1594,In_192,In_967);
and U1595 (N_1595,In_925,In_1427);
xor U1596 (N_1596,In_1264,In_37);
xnor U1597 (N_1597,In_267,In_399);
xnor U1598 (N_1598,In_747,In_953);
or U1599 (N_1599,In_1053,In_5);
or U1600 (N_1600,In_61,In_177);
nand U1601 (N_1601,In_1082,In_68);
and U1602 (N_1602,In_873,In_400);
and U1603 (N_1603,In_76,In_1441);
and U1604 (N_1604,In_673,In_15);
nor U1605 (N_1605,In_281,In_1266);
nand U1606 (N_1606,In_828,In_186);
nor U1607 (N_1607,In_882,In_1154);
xnor U1608 (N_1608,In_380,In_1250);
nor U1609 (N_1609,In_96,In_1386);
nor U1610 (N_1610,In_881,In_135);
nor U1611 (N_1611,In_589,In_2);
nor U1612 (N_1612,In_1285,In_1420);
nand U1613 (N_1613,In_1333,In_1011);
nor U1614 (N_1614,In_1029,In_1409);
xnor U1615 (N_1615,In_1154,In_741);
xnor U1616 (N_1616,In_260,In_1239);
xor U1617 (N_1617,In_323,In_1277);
nor U1618 (N_1618,In_919,In_721);
nor U1619 (N_1619,In_721,In_281);
nor U1620 (N_1620,In_784,In_1257);
and U1621 (N_1621,In_79,In_965);
nand U1622 (N_1622,In_579,In_743);
and U1623 (N_1623,In_1079,In_821);
nor U1624 (N_1624,In_197,In_948);
xnor U1625 (N_1625,In_451,In_17);
or U1626 (N_1626,In_495,In_126);
xnor U1627 (N_1627,In_669,In_290);
xnor U1628 (N_1628,In_1119,In_412);
nand U1629 (N_1629,In_715,In_1297);
nor U1630 (N_1630,In_611,In_1002);
or U1631 (N_1631,In_900,In_1172);
nor U1632 (N_1632,In_885,In_224);
xnor U1633 (N_1633,In_145,In_560);
nand U1634 (N_1634,In_222,In_687);
nand U1635 (N_1635,In_318,In_1365);
xnor U1636 (N_1636,In_1369,In_499);
and U1637 (N_1637,In_1376,In_758);
nand U1638 (N_1638,In_208,In_1388);
or U1639 (N_1639,In_1179,In_0);
nand U1640 (N_1640,In_1013,In_232);
or U1641 (N_1641,In_1326,In_1082);
nor U1642 (N_1642,In_887,In_44);
or U1643 (N_1643,In_432,In_1494);
or U1644 (N_1644,In_1181,In_559);
and U1645 (N_1645,In_261,In_75);
or U1646 (N_1646,In_442,In_1089);
nor U1647 (N_1647,In_864,In_610);
or U1648 (N_1648,In_1024,In_653);
xor U1649 (N_1649,In_1167,In_822);
nand U1650 (N_1650,In_1457,In_27);
or U1651 (N_1651,In_852,In_1218);
nand U1652 (N_1652,In_1252,In_765);
or U1653 (N_1653,In_1044,In_857);
nand U1654 (N_1654,In_436,In_1092);
nor U1655 (N_1655,In_889,In_121);
xnor U1656 (N_1656,In_1088,In_1023);
nor U1657 (N_1657,In_648,In_286);
xor U1658 (N_1658,In_802,In_1168);
or U1659 (N_1659,In_659,In_519);
nor U1660 (N_1660,In_1040,In_71);
and U1661 (N_1661,In_744,In_659);
xnor U1662 (N_1662,In_1011,In_528);
xor U1663 (N_1663,In_856,In_72);
nand U1664 (N_1664,In_1050,In_156);
or U1665 (N_1665,In_707,In_937);
or U1666 (N_1666,In_76,In_347);
nor U1667 (N_1667,In_37,In_1135);
or U1668 (N_1668,In_831,In_1152);
nor U1669 (N_1669,In_736,In_397);
and U1670 (N_1670,In_376,In_874);
and U1671 (N_1671,In_409,In_134);
nand U1672 (N_1672,In_747,In_1354);
or U1673 (N_1673,In_1333,In_1465);
nand U1674 (N_1674,In_693,In_1141);
and U1675 (N_1675,In_740,In_1015);
xnor U1676 (N_1676,In_979,In_880);
and U1677 (N_1677,In_150,In_767);
nor U1678 (N_1678,In_181,In_33);
xnor U1679 (N_1679,In_307,In_801);
nand U1680 (N_1680,In_1196,In_991);
and U1681 (N_1681,In_994,In_607);
nor U1682 (N_1682,In_338,In_659);
nor U1683 (N_1683,In_1204,In_849);
and U1684 (N_1684,In_1074,In_1012);
xor U1685 (N_1685,In_1064,In_1355);
or U1686 (N_1686,In_1204,In_1249);
nand U1687 (N_1687,In_551,In_1420);
xnor U1688 (N_1688,In_1113,In_1206);
xnor U1689 (N_1689,In_1370,In_612);
or U1690 (N_1690,In_624,In_1084);
and U1691 (N_1691,In_511,In_363);
nor U1692 (N_1692,In_711,In_1116);
and U1693 (N_1693,In_796,In_196);
and U1694 (N_1694,In_271,In_89);
nand U1695 (N_1695,In_57,In_432);
nor U1696 (N_1696,In_589,In_931);
and U1697 (N_1697,In_93,In_1277);
xor U1698 (N_1698,In_255,In_404);
nand U1699 (N_1699,In_1400,In_243);
nand U1700 (N_1700,In_966,In_1365);
or U1701 (N_1701,In_444,In_403);
xor U1702 (N_1702,In_981,In_570);
or U1703 (N_1703,In_1060,In_288);
or U1704 (N_1704,In_276,In_95);
xnor U1705 (N_1705,In_930,In_444);
nor U1706 (N_1706,In_427,In_172);
xnor U1707 (N_1707,In_1480,In_1487);
nand U1708 (N_1708,In_744,In_537);
or U1709 (N_1709,In_810,In_444);
nor U1710 (N_1710,In_1456,In_569);
nand U1711 (N_1711,In_1133,In_1393);
nand U1712 (N_1712,In_663,In_386);
or U1713 (N_1713,In_27,In_1406);
nand U1714 (N_1714,In_96,In_702);
and U1715 (N_1715,In_915,In_1010);
nor U1716 (N_1716,In_873,In_906);
xor U1717 (N_1717,In_289,In_376);
xor U1718 (N_1718,In_1493,In_767);
xor U1719 (N_1719,In_999,In_526);
nor U1720 (N_1720,In_366,In_545);
or U1721 (N_1721,In_1438,In_2);
or U1722 (N_1722,In_1423,In_1326);
or U1723 (N_1723,In_968,In_1145);
nor U1724 (N_1724,In_969,In_1053);
xnor U1725 (N_1725,In_104,In_982);
or U1726 (N_1726,In_1301,In_13);
or U1727 (N_1727,In_253,In_1175);
xnor U1728 (N_1728,In_1250,In_719);
nand U1729 (N_1729,In_1435,In_268);
nand U1730 (N_1730,In_514,In_421);
nand U1731 (N_1731,In_1388,In_308);
and U1732 (N_1732,In_1192,In_598);
or U1733 (N_1733,In_279,In_356);
nor U1734 (N_1734,In_572,In_919);
xnor U1735 (N_1735,In_1017,In_1137);
and U1736 (N_1736,In_817,In_1354);
or U1737 (N_1737,In_964,In_1134);
nor U1738 (N_1738,In_934,In_982);
and U1739 (N_1739,In_74,In_754);
xor U1740 (N_1740,In_57,In_713);
and U1741 (N_1741,In_360,In_842);
and U1742 (N_1742,In_57,In_419);
xnor U1743 (N_1743,In_735,In_782);
xor U1744 (N_1744,In_578,In_1461);
and U1745 (N_1745,In_1041,In_307);
and U1746 (N_1746,In_815,In_373);
or U1747 (N_1747,In_58,In_804);
or U1748 (N_1748,In_1049,In_1045);
or U1749 (N_1749,In_589,In_1011);
nor U1750 (N_1750,In_362,In_999);
xor U1751 (N_1751,In_626,In_520);
nor U1752 (N_1752,In_113,In_776);
or U1753 (N_1753,In_1024,In_906);
and U1754 (N_1754,In_1364,In_1449);
nand U1755 (N_1755,In_704,In_623);
or U1756 (N_1756,In_909,In_918);
and U1757 (N_1757,In_1098,In_130);
nor U1758 (N_1758,In_488,In_426);
xnor U1759 (N_1759,In_319,In_1369);
or U1760 (N_1760,In_1131,In_1220);
or U1761 (N_1761,In_1434,In_725);
and U1762 (N_1762,In_635,In_536);
nand U1763 (N_1763,In_1097,In_1085);
xnor U1764 (N_1764,In_573,In_840);
xor U1765 (N_1765,In_1048,In_1409);
nand U1766 (N_1766,In_92,In_364);
and U1767 (N_1767,In_161,In_21);
nand U1768 (N_1768,In_523,In_1133);
or U1769 (N_1769,In_727,In_109);
xnor U1770 (N_1770,In_421,In_1170);
xnor U1771 (N_1771,In_361,In_437);
and U1772 (N_1772,In_572,In_151);
or U1773 (N_1773,In_1086,In_814);
nor U1774 (N_1774,In_222,In_674);
and U1775 (N_1775,In_7,In_573);
nand U1776 (N_1776,In_1394,In_896);
nand U1777 (N_1777,In_376,In_91);
and U1778 (N_1778,In_963,In_1194);
nor U1779 (N_1779,In_675,In_1311);
or U1780 (N_1780,In_1072,In_1176);
nand U1781 (N_1781,In_220,In_1107);
nand U1782 (N_1782,In_523,In_423);
or U1783 (N_1783,In_568,In_1478);
or U1784 (N_1784,In_1478,In_1463);
nand U1785 (N_1785,In_410,In_97);
xor U1786 (N_1786,In_1202,In_153);
or U1787 (N_1787,In_229,In_305);
and U1788 (N_1788,In_885,In_986);
xor U1789 (N_1789,In_975,In_1333);
or U1790 (N_1790,In_33,In_1039);
nand U1791 (N_1791,In_458,In_693);
or U1792 (N_1792,In_1377,In_263);
nor U1793 (N_1793,In_673,In_937);
and U1794 (N_1794,In_1244,In_906);
xor U1795 (N_1795,In_1244,In_1128);
or U1796 (N_1796,In_548,In_586);
nor U1797 (N_1797,In_962,In_464);
and U1798 (N_1798,In_224,In_192);
nand U1799 (N_1799,In_966,In_1318);
and U1800 (N_1800,In_580,In_184);
nand U1801 (N_1801,In_954,In_1487);
and U1802 (N_1802,In_25,In_142);
nand U1803 (N_1803,In_1092,In_534);
or U1804 (N_1804,In_1265,In_888);
xor U1805 (N_1805,In_840,In_1274);
or U1806 (N_1806,In_424,In_1264);
nor U1807 (N_1807,In_328,In_1304);
xor U1808 (N_1808,In_460,In_1032);
and U1809 (N_1809,In_335,In_1157);
and U1810 (N_1810,In_1285,In_391);
and U1811 (N_1811,In_517,In_1009);
nor U1812 (N_1812,In_1221,In_391);
and U1813 (N_1813,In_183,In_506);
or U1814 (N_1814,In_1147,In_904);
or U1815 (N_1815,In_418,In_325);
nor U1816 (N_1816,In_1389,In_1443);
and U1817 (N_1817,In_533,In_921);
nand U1818 (N_1818,In_370,In_841);
or U1819 (N_1819,In_918,In_1031);
xnor U1820 (N_1820,In_591,In_12);
nand U1821 (N_1821,In_269,In_909);
nor U1822 (N_1822,In_504,In_297);
xnor U1823 (N_1823,In_1210,In_615);
nand U1824 (N_1824,In_278,In_437);
nand U1825 (N_1825,In_377,In_399);
nor U1826 (N_1826,In_289,In_1048);
and U1827 (N_1827,In_565,In_562);
or U1828 (N_1828,In_500,In_113);
or U1829 (N_1829,In_910,In_1061);
and U1830 (N_1830,In_1255,In_432);
xnor U1831 (N_1831,In_428,In_1421);
xor U1832 (N_1832,In_464,In_228);
nor U1833 (N_1833,In_134,In_1319);
xor U1834 (N_1834,In_1351,In_368);
xor U1835 (N_1835,In_792,In_126);
xor U1836 (N_1836,In_919,In_1281);
and U1837 (N_1837,In_611,In_1414);
and U1838 (N_1838,In_1337,In_120);
and U1839 (N_1839,In_8,In_247);
nor U1840 (N_1840,In_1062,In_839);
and U1841 (N_1841,In_880,In_1380);
and U1842 (N_1842,In_250,In_1326);
xor U1843 (N_1843,In_11,In_197);
nand U1844 (N_1844,In_1212,In_211);
and U1845 (N_1845,In_545,In_1195);
or U1846 (N_1846,In_1266,In_239);
or U1847 (N_1847,In_341,In_1180);
xnor U1848 (N_1848,In_1489,In_1434);
nor U1849 (N_1849,In_923,In_1497);
xnor U1850 (N_1850,In_1156,In_75);
xnor U1851 (N_1851,In_377,In_1449);
nand U1852 (N_1852,In_1402,In_104);
or U1853 (N_1853,In_222,In_1496);
xnor U1854 (N_1854,In_1020,In_839);
nand U1855 (N_1855,In_504,In_610);
and U1856 (N_1856,In_899,In_962);
and U1857 (N_1857,In_359,In_130);
nand U1858 (N_1858,In_834,In_547);
and U1859 (N_1859,In_1160,In_105);
nor U1860 (N_1860,In_1136,In_1311);
and U1861 (N_1861,In_795,In_852);
nand U1862 (N_1862,In_1457,In_285);
xor U1863 (N_1863,In_54,In_725);
or U1864 (N_1864,In_1378,In_1442);
or U1865 (N_1865,In_783,In_750);
or U1866 (N_1866,In_484,In_553);
and U1867 (N_1867,In_623,In_1027);
and U1868 (N_1868,In_698,In_314);
or U1869 (N_1869,In_1283,In_595);
nor U1870 (N_1870,In_1221,In_997);
and U1871 (N_1871,In_294,In_139);
and U1872 (N_1872,In_597,In_1121);
nor U1873 (N_1873,In_735,In_246);
xnor U1874 (N_1874,In_174,In_905);
nand U1875 (N_1875,In_1255,In_147);
nor U1876 (N_1876,In_586,In_420);
or U1877 (N_1877,In_1348,In_1245);
nand U1878 (N_1878,In_239,In_1101);
or U1879 (N_1879,In_118,In_470);
nor U1880 (N_1880,In_810,In_874);
or U1881 (N_1881,In_168,In_584);
nand U1882 (N_1882,In_1204,In_982);
xnor U1883 (N_1883,In_146,In_607);
nand U1884 (N_1884,In_665,In_870);
nand U1885 (N_1885,In_920,In_1104);
nor U1886 (N_1886,In_517,In_126);
and U1887 (N_1887,In_1167,In_971);
nor U1888 (N_1888,In_950,In_25);
or U1889 (N_1889,In_383,In_484);
nor U1890 (N_1890,In_850,In_1076);
and U1891 (N_1891,In_536,In_1390);
nand U1892 (N_1892,In_443,In_483);
xor U1893 (N_1893,In_1158,In_1497);
xor U1894 (N_1894,In_85,In_966);
nor U1895 (N_1895,In_171,In_925);
or U1896 (N_1896,In_984,In_445);
nor U1897 (N_1897,In_224,In_702);
or U1898 (N_1898,In_405,In_230);
nand U1899 (N_1899,In_661,In_857);
or U1900 (N_1900,In_1250,In_1235);
nand U1901 (N_1901,In_859,In_293);
xor U1902 (N_1902,In_82,In_166);
nor U1903 (N_1903,In_998,In_929);
xor U1904 (N_1904,In_530,In_766);
xnor U1905 (N_1905,In_614,In_250);
nor U1906 (N_1906,In_1364,In_1083);
nor U1907 (N_1907,In_370,In_1046);
or U1908 (N_1908,In_1438,In_990);
nor U1909 (N_1909,In_407,In_1492);
nor U1910 (N_1910,In_1244,In_565);
xnor U1911 (N_1911,In_238,In_857);
or U1912 (N_1912,In_493,In_57);
or U1913 (N_1913,In_883,In_432);
and U1914 (N_1914,In_844,In_1424);
or U1915 (N_1915,In_1226,In_473);
nor U1916 (N_1916,In_35,In_430);
and U1917 (N_1917,In_1116,In_1136);
nor U1918 (N_1918,In_1102,In_1022);
or U1919 (N_1919,In_57,In_538);
nand U1920 (N_1920,In_460,In_314);
nand U1921 (N_1921,In_174,In_1042);
or U1922 (N_1922,In_844,In_342);
and U1923 (N_1923,In_387,In_1258);
xor U1924 (N_1924,In_557,In_533);
and U1925 (N_1925,In_1351,In_1336);
nand U1926 (N_1926,In_266,In_795);
nand U1927 (N_1927,In_1482,In_682);
and U1928 (N_1928,In_379,In_43);
nor U1929 (N_1929,In_786,In_911);
or U1930 (N_1930,In_127,In_1098);
nand U1931 (N_1931,In_805,In_212);
or U1932 (N_1932,In_1056,In_597);
and U1933 (N_1933,In_99,In_863);
or U1934 (N_1934,In_1417,In_1219);
or U1935 (N_1935,In_376,In_436);
or U1936 (N_1936,In_993,In_94);
nand U1937 (N_1937,In_432,In_112);
xor U1938 (N_1938,In_208,In_587);
nand U1939 (N_1939,In_553,In_1171);
xnor U1940 (N_1940,In_262,In_1012);
and U1941 (N_1941,In_489,In_658);
nand U1942 (N_1942,In_67,In_236);
nor U1943 (N_1943,In_992,In_476);
or U1944 (N_1944,In_48,In_793);
nand U1945 (N_1945,In_559,In_334);
nand U1946 (N_1946,In_1459,In_273);
xnor U1947 (N_1947,In_554,In_41);
nor U1948 (N_1948,In_728,In_464);
and U1949 (N_1949,In_1281,In_350);
and U1950 (N_1950,In_621,In_1466);
nor U1951 (N_1951,In_922,In_158);
nand U1952 (N_1952,In_1365,In_392);
xnor U1953 (N_1953,In_1379,In_1444);
xor U1954 (N_1954,In_355,In_646);
nand U1955 (N_1955,In_727,In_36);
nand U1956 (N_1956,In_109,In_1005);
nand U1957 (N_1957,In_1143,In_0);
or U1958 (N_1958,In_1223,In_235);
nand U1959 (N_1959,In_69,In_1154);
or U1960 (N_1960,In_776,In_159);
or U1961 (N_1961,In_1448,In_1483);
xor U1962 (N_1962,In_1266,In_829);
and U1963 (N_1963,In_1295,In_1383);
and U1964 (N_1964,In_175,In_1199);
nor U1965 (N_1965,In_907,In_792);
xor U1966 (N_1966,In_1140,In_976);
nand U1967 (N_1967,In_439,In_943);
and U1968 (N_1968,In_876,In_66);
and U1969 (N_1969,In_401,In_1089);
nand U1970 (N_1970,In_1131,In_1206);
nor U1971 (N_1971,In_1163,In_1173);
or U1972 (N_1972,In_1138,In_1250);
xnor U1973 (N_1973,In_71,In_992);
xnor U1974 (N_1974,In_994,In_977);
nand U1975 (N_1975,In_1224,In_649);
and U1976 (N_1976,In_546,In_638);
nand U1977 (N_1977,In_679,In_1451);
xor U1978 (N_1978,In_244,In_290);
or U1979 (N_1979,In_180,In_453);
and U1980 (N_1980,In_1033,In_909);
and U1981 (N_1981,In_687,In_33);
and U1982 (N_1982,In_530,In_239);
nor U1983 (N_1983,In_80,In_861);
nand U1984 (N_1984,In_990,In_255);
xnor U1985 (N_1985,In_1034,In_953);
nand U1986 (N_1986,In_772,In_420);
or U1987 (N_1987,In_1379,In_256);
nand U1988 (N_1988,In_1449,In_1036);
xor U1989 (N_1989,In_1309,In_819);
xor U1990 (N_1990,In_454,In_1320);
or U1991 (N_1991,In_174,In_1339);
nor U1992 (N_1992,In_82,In_1447);
or U1993 (N_1993,In_154,In_1273);
nand U1994 (N_1994,In_1100,In_497);
and U1995 (N_1995,In_1106,In_83);
xnor U1996 (N_1996,In_231,In_421);
nor U1997 (N_1997,In_261,In_1438);
nor U1998 (N_1998,In_52,In_925);
or U1999 (N_1999,In_873,In_697);
or U2000 (N_2000,In_88,In_1083);
nor U2001 (N_2001,In_1297,In_926);
xnor U2002 (N_2002,In_612,In_1081);
nand U2003 (N_2003,In_772,In_999);
nor U2004 (N_2004,In_193,In_544);
nor U2005 (N_2005,In_44,In_612);
xor U2006 (N_2006,In_1015,In_1177);
nand U2007 (N_2007,In_545,In_1399);
xnor U2008 (N_2008,In_958,In_346);
nand U2009 (N_2009,In_1043,In_1365);
nand U2010 (N_2010,In_783,In_737);
xnor U2011 (N_2011,In_466,In_897);
or U2012 (N_2012,In_1187,In_14);
and U2013 (N_2013,In_1241,In_1165);
nor U2014 (N_2014,In_739,In_965);
and U2015 (N_2015,In_533,In_1120);
or U2016 (N_2016,In_922,In_1337);
and U2017 (N_2017,In_1082,In_916);
nor U2018 (N_2018,In_1372,In_1194);
nand U2019 (N_2019,In_784,In_175);
xor U2020 (N_2020,In_456,In_575);
xor U2021 (N_2021,In_1133,In_418);
nand U2022 (N_2022,In_734,In_1128);
and U2023 (N_2023,In_1005,In_111);
nand U2024 (N_2024,In_1351,In_559);
nand U2025 (N_2025,In_333,In_1163);
nand U2026 (N_2026,In_1115,In_999);
nor U2027 (N_2027,In_667,In_229);
and U2028 (N_2028,In_1168,In_708);
and U2029 (N_2029,In_430,In_597);
xor U2030 (N_2030,In_1461,In_942);
or U2031 (N_2031,In_1141,In_276);
xnor U2032 (N_2032,In_394,In_1499);
and U2033 (N_2033,In_801,In_35);
or U2034 (N_2034,In_381,In_893);
and U2035 (N_2035,In_537,In_644);
xnor U2036 (N_2036,In_384,In_956);
xnor U2037 (N_2037,In_1314,In_410);
or U2038 (N_2038,In_83,In_1176);
xor U2039 (N_2039,In_1149,In_112);
nor U2040 (N_2040,In_953,In_104);
nand U2041 (N_2041,In_32,In_508);
nand U2042 (N_2042,In_1158,In_1001);
nor U2043 (N_2043,In_75,In_809);
and U2044 (N_2044,In_971,In_257);
xnor U2045 (N_2045,In_1479,In_754);
nor U2046 (N_2046,In_316,In_120);
xor U2047 (N_2047,In_656,In_513);
or U2048 (N_2048,In_286,In_941);
nor U2049 (N_2049,In_1368,In_1302);
xor U2050 (N_2050,In_401,In_259);
or U2051 (N_2051,In_608,In_363);
or U2052 (N_2052,In_1293,In_1195);
xor U2053 (N_2053,In_1373,In_604);
nand U2054 (N_2054,In_821,In_441);
nand U2055 (N_2055,In_370,In_830);
or U2056 (N_2056,In_11,In_318);
nand U2057 (N_2057,In_1075,In_938);
or U2058 (N_2058,In_1352,In_437);
nor U2059 (N_2059,In_835,In_65);
and U2060 (N_2060,In_31,In_1196);
nor U2061 (N_2061,In_951,In_16);
xnor U2062 (N_2062,In_1003,In_960);
nor U2063 (N_2063,In_568,In_1365);
xnor U2064 (N_2064,In_292,In_395);
and U2065 (N_2065,In_649,In_963);
nor U2066 (N_2066,In_1033,In_223);
nand U2067 (N_2067,In_793,In_652);
or U2068 (N_2068,In_606,In_176);
xor U2069 (N_2069,In_783,In_1079);
nand U2070 (N_2070,In_1110,In_407);
and U2071 (N_2071,In_195,In_772);
nand U2072 (N_2072,In_1078,In_166);
and U2073 (N_2073,In_1002,In_658);
nor U2074 (N_2074,In_264,In_501);
nand U2075 (N_2075,In_1061,In_775);
xnor U2076 (N_2076,In_666,In_59);
nand U2077 (N_2077,In_1201,In_1159);
or U2078 (N_2078,In_746,In_288);
nand U2079 (N_2079,In_1424,In_856);
and U2080 (N_2080,In_648,In_297);
and U2081 (N_2081,In_464,In_150);
and U2082 (N_2082,In_566,In_346);
xnor U2083 (N_2083,In_683,In_50);
or U2084 (N_2084,In_568,In_969);
xnor U2085 (N_2085,In_566,In_1196);
or U2086 (N_2086,In_110,In_200);
and U2087 (N_2087,In_341,In_221);
or U2088 (N_2088,In_381,In_1112);
and U2089 (N_2089,In_190,In_1006);
xnor U2090 (N_2090,In_584,In_773);
or U2091 (N_2091,In_1107,In_1262);
xnor U2092 (N_2092,In_707,In_42);
or U2093 (N_2093,In_521,In_121);
xnor U2094 (N_2094,In_1267,In_926);
xor U2095 (N_2095,In_1379,In_159);
nand U2096 (N_2096,In_1024,In_884);
nor U2097 (N_2097,In_473,In_877);
nand U2098 (N_2098,In_419,In_349);
and U2099 (N_2099,In_1273,In_1406);
nor U2100 (N_2100,In_704,In_406);
or U2101 (N_2101,In_244,In_745);
or U2102 (N_2102,In_256,In_325);
and U2103 (N_2103,In_1169,In_874);
or U2104 (N_2104,In_975,In_126);
nand U2105 (N_2105,In_871,In_888);
and U2106 (N_2106,In_418,In_144);
nor U2107 (N_2107,In_1434,In_299);
or U2108 (N_2108,In_379,In_710);
xor U2109 (N_2109,In_1228,In_1484);
nand U2110 (N_2110,In_541,In_774);
nor U2111 (N_2111,In_1071,In_270);
nand U2112 (N_2112,In_1239,In_1188);
xnor U2113 (N_2113,In_1396,In_203);
xor U2114 (N_2114,In_766,In_1088);
nor U2115 (N_2115,In_1425,In_783);
nand U2116 (N_2116,In_528,In_819);
and U2117 (N_2117,In_1018,In_927);
nor U2118 (N_2118,In_657,In_751);
xnor U2119 (N_2119,In_207,In_439);
or U2120 (N_2120,In_844,In_1389);
nand U2121 (N_2121,In_1499,In_969);
nor U2122 (N_2122,In_574,In_386);
nor U2123 (N_2123,In_299,In_888);
or U2124 (N_2124,In_671,In_229);
nand U2125 (N_2125,In_246,In_1113);
xnor U2126 (N_2126,In_645,In_69);
and U2127 (N_2127,In_825,In_592);
nor U2128 (N_2128,In_1140,In_1269);
or U2129 (N_2129,In_782,In_314);
or U2130 (N_2130,In_1021,In_986);
nand U2131 (N_2131,In_1235,In_99);
xor U2132 (N_2132,In_1396,In_1153);
nand U2133 (N_2133,In_1169,In_1104);
or U2134 (N_2134,In_903,In_146);
or U2135 (N_2135,In_42,In_860);
or U2136 (N_2136,In_243,In_980);
xor U2137 (N_2137,In_416,In_683);
or U2138 (N_2138,In_192,In_574);
and U2139 (N_2139,In_1362,In_128);
xor U2140 (N_2140,In_1225,In_482);
nand U2141 (N_2141,In_560,In_1290);
and U2142 (N_2142,In_463,In_1296);
nand U2143 (N_2143,In_1380,In_102);
or U2144 (N_2144,In_97,In_814);
nor U2145 (N_2145,In_131,In_438);
or U2146 (N_2146,In_308,In_1193);
nand U2147 (N_2147,In_1326,In_308);
and U2148 (N_2148,In_188,In_1241);
and U2149 (N_2149,In_488,In_337);
and U2150 (N_2150,In_193,In_970);
and U2151 (N_2151,In_246,In_1425);
or U2152 (N_2152,In_746,In_1348);
xor U2153 (N_2153,In_874,In_439);
or U2154 (N_2154,In_932,In_1029);
or U2155 (N_2155,In_1167,In_433);
and U2156 (N_2156,In_884,In_131);
xnor U2157 (N_2157,In_776,In_523);
nand U2158 (N_2158,In_1418,In_906);
nand U2159 (N_2159,In_1221,In_436);
and U2160 (N_2160,In_540,In_935);
or U2161 (N_2161,In_1388,In_144);
and U2162 (N_2162,In_265,In_389);
or U2163 (N_2163,In_1033,In_360);
nand U2164 (N_2164,In_670,In_1457);
or U2165 (N_2165,In_496,In_410);
nor U2166 (N_2166,In_980,In_1138);
xor U2167 (N_2167,In_590,In_433);
nand U2168 (N_2168,In_1093,In_446);
nor U2169 (N_2169,In_1060,In_27);
xor U2170 (N_2170,In_304,In_582);
nand U2171 (N_2171,In_828,In_1034);
nor U2172 (N_2172,In_430,In_977);
or U2173 (N_2173,In_282,In_1101);
or U2174 (N_2174,In_895,In_307);
or U2175 (N_2175,In_1116,In_1292);
nor U2176 (N_2176,In_203,In_785);
nand U2177 (N_2177,In_77,In_409);
nor U2178 (N_2178,In_154,In_1478);
or U2179 (N_2179,In_1225,In_1072);
nor U2180 (N_2180,In_506,In_1307);
or U2181 (N_2181,In_540,In_136);
nand U2182 (N_2182,In_1324,In_915);
or U2183 (N_2183,In_726,In_1214);
or U2184 (N_2184,In_448,In_1298);
xnor U2185 (N_2185,In_997,In_873);
nor U2186 (N_2186,In_234,In_1428);
nor U2187 (N_2187,In_244,In_5);
or U2188 (N_2188,In_1417,In_489);
and U2189 (N_2189,In_1011,In_1154);
nor U2190 (N_2190,In_1471,In_1147);
xor U2191 (N_2191,In_588,In_903);
or U2192 (N_2192,In_445,In_550);
or U2193 (N_2193,In_259,In_996);
and U2194 (N_2194,In_939,In_1402);
nor U2195 (N_2195,In_1080,In_571);
nor U2196 (N_2196,In_471,In_419);
and U2197 (N_2197,In_1395,In_912);
nand U2198 (N_2198,In_82,In_1112);
or U2199 (N_2199,In_953,In_1042);
nand U2200 (N_2200,In_434,In_1154);
nor U2201 (N_2201,In_1283,In_510);
nor U2202 (N_2202,In_65,In_1293);
nor U2203 (N_2203,In_108,In_394);
nand U2204 (N_2204,In_184,In_629);
nand U2205 (N_2205,In_132,In_250);
and U2206 (N_2206,In_1387,In_1333);
and U2207 (N_2207,In_677,In_1104);
nor U2208 (N_2208,In_853,In_138);
and U2209 (N_2209,In_424,In_342);
and U2210 (N_2210,In_832,In_271);
and U2211 (N_2211,In_491,In_361);
nand U2212 (N_2212,In_463,In_1209);
xor U2213 (N_2213,In_541,In_1461);
nand U2214 (N_2214,In_417,In_614);
or U2215 (N_2215,In_355,In_671);
nor U2216 (N_2216,In_622,In_598);
and U2217 (N_2217,In_387,In_454);
xnor U2218 (N_2218,In_454,In_544);
nand U2219 (N_2219,In_28,In_1445);
or U2220 (N_2220,In_1106,In_290);
xnor U2221 (N_2221,In_1148,In_743);
nand U2222 (N_2222,In_922,In_55);
or U2223 (N_2223,In_1169,In_1268);
or U2224 (N_2224,In_1279,In_1255);
or U2225 (N_2225,In_921,In_577);
nor U2226 (N_2226,In_525,In_1050);
xnor U2227 (N_2227,In_1212,In_652);
or U2228 (N_2228,In_260,In_1462);
and U2229 (N_2229,In_675,In_421);
and U2230 (N_2230,In_181,In_1332);
and U2231 (N_2231,In_1293,In_320);
nand U2232 (N_2232,In_1383,In_423);
nand U2233 (N_2233,In_247,In_202);
nand U2234 (N_2234,In_1067,In_86);
xnor U2235 (N_2235,In_1033,In_961);
nand U2236 (N_2236,In_816,In_79);
or U2237 (N_2237,In_562,In_883);
and U2238 (N_2238,In_635,In_189);
nor U2239 (N_2239,In_373,In_200);
nand U2240 (N_2240,In_288,In_796);
and U2241 (N_2241,In_242,In_532);
and U2242 (N_2242,In_107,In_1408);
and U2243 (N_2243,In_812,In_770);
nor U2244 (N_2244,In_1418,In_615);
nor U2245 (N_2245,In_369,In_612);
nand U2246 (N_2246,In_284,In_880);
or U2247 (N_2247,In_547,In_678);
nor U2248 (N_2248,In_1213,In_877);
nor U2249 (N_2249,In_727,In_1030);
xnor U2250 (N_2250,In_45,In_510);
nor U2251 (N_2251,In_247,In_452);
nor U2252 (N_2252,In_605,In_1070);
xor U2253 (N_2253,In_369,In_666);
xor U2254 (N_2254,In_1327,In_431);
and U2255 (N_2255,In_1133,In_1288);
nand U2256 (N_2256,In_167,In_84);
xor U2257 (N_2257,In_1280,In_521);
xnor U2258 (N_2258,In_489,In_611);
or U2259 (N_2259,In_611,In_898);
nor U2260 (N_2260,In_86,In_127);
nand U2261 (N_2261,In_587,In_917);
nand U2262 (N_2262,In_1227,In_718);
nand U2263 (N_2263,In_1209,In_703);
nand U2264 (N_2264,In_250,In_222);
and U2265 (N_2265,In_163,In_1390);
nor U2266 (N_2266,In_530,In_1483);
or U2267 (N_2267,In_1126,In_668);
xor U2268 (N_2268,In_1202,In_979);
or U2269 (N_2269,In_1044,In_322);
xnor U2270 (N_2270,In_83,In_963);
nor U2271 (N_2271,In_1024,In_971);
or U2272 (N_2272,In_314,In_308);
nand U2273 (N_2273,In_15,In_1095);
nand U2274 (N_2274,In_773,In_1314);
nor U2275 (N_2275,In_466,In_1285);
nor U2276 (N_2276,In_961,In_188);
or U2277 (N_2277,In_1086,In_898);
nand U2278 (N_2278,In_1397,In_683);
or U2279 (N_2279,In_1002,In_373);
xnor U2280 (N_2280,In_1175,In_297);
nand U2281 (N_2281,In_749,In_16);
nor U2282 (N_2282,In_1178,In_620);
nor U2283 (N_2283,In_762,In_1026);
xnor U2284 (N_2284,In_271,In_1206);
nor U2285 (N_2285,In_495,In_949);
nor U2286 (N_2286,In_1086,In_1391);
nor U2287 (N_2287,In_1352,In_1004);
nor U2288 (N_2288,In_299,In_177);
xnor U2289 (N_2289,In_330,In_231);
nor U2290 (N_2290,In_1185,In_945);
nand U2291 (N_2291,In_1203,In_1074);
and U2292 (N_2292,In_138,In_1224);
and U2293 (N_2293,In_364,In_460);
nand U2294 (N_2294,In_1104,In_1413);
or U2295 (N_2295,In_248,In_732);
or U2296 (N_2296,In_1416,In_1167);
and U2297 (N_2297,In_1386,In_1112);
nand U2298 (N_2298,In_1100,In_930);
and U2299 (N_2299,In_870,In_505);
and U2300 (N_2300,In_578,In_1288);
nor U2301 (N_2301,In_507,In_1143);
nand U2302 (N_2302,In_1289,In_1427);
nand U2303 (N_2303,In_766,In_208);
nand U2304 (N_2304,In_1213,In_548);
nand U2305 (N_2305,In_1239,In_1087);
nand U2306 (N_2306,In_1091,In_1110);
or U2307 (N_2307,In_478,In_912);
or U2308 (N_2308,In_168,In_617);
nand U2309 (N_2309,In_1431,In_1452);
nor U2310 (N_2310,In_286,In_1336);
nand U2311 (N_2311,In_770,In_683);
nor U2312 (N_2312,In_161,In_997);
nand U2313 (N_2313,In_962,In_750);
xnor U2314 (N_2314,In_547,In_925);
or U2315 (N_2315,In_1026,In_370);
or U2316 (N_2316,In_1453,In_1127);
and U2317 (N_2317,In_767,In_248);
nand U2318 (N_2318,In_1332,In_341);
nand U2319 (N_2319,In_1273,In_1216);
nand U2320 (N_2320,In_1237,In_339);
or U2321 (N_2321,In_753,In_1247);
nor U2322 (N_2322,In_523,In_753);
or U2323 (N_2323,In_1021,In_266);
nor U2324 (N_2324,In_1076,In_292);
or U2325 (N_2325,In_558,In_274);
xor U2326 (N_2326,In_932,In_1108);
xnor U2327 (N_2327,In_378,In_1236);
and U2328 (N_2328,In_956,In_1214);
or U2329 (N_2329,In_885,In_1386);
or U2330 (N_2330,In_1092,In_411);
and U2331 (N_2331,In_43,In_946);
or U2332 (N_2332,In_31,In_1250);
nand U2333 (N_2333,In_79,In_669);
or U2334 (N_2334,In_1027,In_480);
nand U2335 (N_2335,In_822,In_1176);
nand U2336 (N_2336,In_601,In_898);
and U2337 (N_2337,In_529,In_140);
and U2338 (N_2338,In_184,In_1413);
and U2339 (N_2339,In_786,In_185);
and U2340 (N_2340,In_61,In_419);
nor U2341 (N_2341,In_4,In_1243);
or U2342 (N_2342,In_1165,In_1261);
xor U2343 (N_2343,In_1007,In_316);
nand U2344 (N_2344,In_604,In_223);
and U2345 (N_2345,In_591,In_955);
xor U2346 (N_2346,In_336,In_1002);
or U2347 (N_2347,In_97,In_1386);
xnor U2348 (N_2348,In_157,In_1071);
xor U2349 (N_2349,In_1038,In_1464);
nand U2350 (N_2350,In_230,In_1176);
or U2351 (N_2351,In_13,In_1025);
xnor U2352 (N_2352,In_583,In_1093);
nand U2353 (N_2353,In_873,In_1170);
or U2354 (N_2354,In_580,In_788);
xnor U2355 (N_2355,In_253,In_506);
nor U2356 (N_2356,In_146,In_603);
nor U2357 (N_2357,In_40,In_1484);
nor U2358 (N_2358,In_1185,In_126);
nor U2359 (N_2359,In_872,In_198);
xor U2360 (N_2360,In_1266,In_758);
xor U2361 (N_2361,In_347,In_390);
or U2362 (N_2362,In_353,In_1022);
or U2363 (N_2363,In_1053,In_699);
nor U2364 (N_2364,In_1322,In_711);
or U2365 (N_2365,In_1048,In_1291);
nor U2366 (N_2366,In_100,In_1490);
nor U2367 (N_2367,In_821,In_1037);
nor U2368 (N_2368,In_1300,In_229);
xnor U2369 (N_2369,In_682,In_315);
or U2370 (N_2370,In_1025,In_41);
or U2371 (N_2371,In_1141,In_1444);
nor U2372 (N_2372,In_1020,In_665);
xor U2373 (N_2373,In_236,In_53);
or U2374 (N_2374,In_238,In_1051);
nor U2375 (N_2375,In_932,In_276);
xor U2376 (N_2376,In_155,In_459);
nor U2377 (N_2377,In_374,In_1463);
or U2378 (N_2378,In_429,In_295);
nand U2379 (N_2379,In_1256,In_38);
or U2380 (N_2380,In_1325,In_1219);
nor U2381 (N_2381,In_261,In_415);
and U2382 (N_2382,In_1317,In_108);
and U2383 (N_2383,In_1040,In_670);
and U2384 (N_2384,In_334,In_1250);
nand U2385 (N_2385,In_116,In_150);
and U2386 (N_2386,In_360,In_199);
nand U2387 (N_2387,In_1449,In_724);
nand U2388 (N_2388,In_461,In_1466);
nor U2389 (N_2389,In_397,In_1394);
or U2390 (N_2390,In_423,In_220);
nor U2391 (N_2391,In_1292,In_74);
nor U2392 (N_2392,In_10,In_1171);
nand U2393 (N_2393,In_1071,In_208);
or U2394 (N_2394,In_396,In_143);
xnor U2395 (N_2395,In_904,In_1291);
and U2396 (N_2396,In_1394,In_997);
nor U2397 (N_2397,In_882,In_515);
nand U2398 (N_2398,In_493,In_534);
nor U2399 (N_2399,In_917,In_660);
xor U2400 (N_2400,In_448,In_240);
and U2401 (N_2401,In_573,In_738);
or U2402 (N_2402,In_675,In_1308);
or U2403 (N_2403,In_569,In_772);
xor U2404 (N_2404,In_482,In_823);
xor U2405 (N_2405,In_374,In_579);
nor U2406 (N_2406,In_996,In_638);
or U2407 (N_2407,In_217,In_721);
and U2408 (N_2408,In_1268,In_528);
nor U2409 (N_2409,In_638,In_670);
or U2410 (N_2410,In_1378,In_770);
nor U2411 (N_2411,In_1100,In_502);
xnor U2412 (N_2412,In_669,In_1239);
nand U2413 (N_2413,In_688,In_1405);
and U2414 (N_2414,In_882,In_668);
nor U2415 (N_2415,In_856,In_156);
nand U2416 (N_2416,In_1303,In_665);
nor U2417 (N_2417,In_1007,In_1376);
nand U2418 (N_2418,In_136,In_101);
nor U2419 (N_2419,In_1188,In_1317);
nand U2420 (N_2420,In_406,In_919);
and U2421 (N_2421,In_1234,In_94);
and U2422 (N_2422,In_1028,In_45);
or U2423 (N_2423,In_295,In_374);
or U2424 (N_2424,In_1412,In_266);
nand U2425 (N_2425,In_412,In_829);
nor U2426 (N_2426,In_1362,In_1409);
or U2427 (N_2427,In_1312,In_1020);
xor U2428 (N_2428,In_1427,In_1026);
nand U2429 (N_2429,In_722,In_1468);
nor U2430 (N_2430,In_762,In_1157);
nor U2431 (N_2431,In_762,In_1473);
xnor U2432 (N_2432,In_973,In_473);
nor U2433 (N_2433,In_1258,In_813);
or U2434 (N_2434,In_1464,In_549);
xnor U2435 (N_2435,In_890,In_498);
nor U2436 (N_2436,In_107,In_780);
xnor U2437 (N_2437,In_1325,In_967);
xor U2438 (N_2438,In_1089,In_813);
xor U2439 (N_2439,In_1402,In_1110);
nor U2440 (N_2440,In_448,In_232);
nor U2441 (N_2441,In_780,In_351);
nor U2442 (N_2442,In_875,In_1326);
nand U2443 (N_2443,In_1491,In_210);
or U2444 (N_2444,In_1167,In_926);
nand U2445 (N_2445,In_907,In_496);
xor U2446 (N_2446,In_737,In_24);
nor U2447 (N_2447,In_1187,In_770);
and U2448 (N_2448,In_698,In_78);
xnor U2449 (N_2449,In_496,In_351);
and U2450 (N_2450,In_1189,In_1256);
xor U2451 (N_2451,In_95,In_844);
or U2452 (N_2452,In_107,In_98);
and U2453 (N_2453,In_1362,In_1344);
and U2454 (N_2454,In_599,In_823);
and U2455 (N_2455,In_66,In_1084);
nand U2456 (N_2456,In_129,In_1322);
nor U2457 (N_2457,In_152,In_51);
or U2458 (N_2458,In_310,In_580);
or U2459 (N_2459,In_78,In_1337);
or U2460 (N_2460,In_70,In_913);
nor U2461 (N_2461,In_1071,In_827);
or U2462 (N_2462,In_1415,In_926);
and U2463 (N_2463,In_5,In_678);
and U2464 (N_2464,In_1232,In_1000);
or U2465 (N_2465,In_1077,In_947);
nor U2466 (N_2466,In_440,In_846);
or U2467 (N_2467,In_1039,In_58);
nor U2468 (N_2468,In_96,In_1029);
nor U2469 (N_2469,In_925,In_1222);
xnor U2470 (N_2470,In_790,In_620);
nor U2471 (N_2471,In_1122,In_1325);
or U2472 (N_2472,In_341,In_504);
xor U2473 (N_2473,In_1345,In_1213);
nand U2474 (N_2474,In_31,In_990);
xnor U2475 (N_2475,In_23,In_1126);
nor U2476 (N_2476,In_1168,In_1313);
nand U2477 (N_2477,In_212,In_82);
nor U2478 (N_2478,In_335,In_298);
and U2479 (N_2479,In_592,In_103);
nand U2480 (N_2480,In_847,In_1130);
nor U2481 (N_2481,In_923,In_1435);
or U2482 (N_2482,In_1417,In_835);
nand U2483 (N_2483,In_1211,In_745);
nand U2484 (N_2484,In_919,In_418);
nand U2485 (N_2485,In_530,In_1155);
and U2486 (N_2486,In_487,In_439);
xnor U2487 (N_2487,In_1056,In_347);
or U2488 (N_2488,In_1212,In_1066);
or U2489 (N_2489,In_1282,In_147);
or U2490 (N_2490,In_291,In_739);
or U2491 (N_2491,In_646,In_694);
nor U2492 (N_2492,In_1009,In_1409);
xor U2493 (N_2493,In_1117,In_1353);
nand U2494 (N_2494,In_846,In_226);
xnor U2495 (N_2495,In_962,In_146);
nor U2496 (N_2496,In_430,In_1048);
or U2497 (N_2497,In_1111,In_283);
and U2498 (N_2498,In_337,In_1023);
and U2499 (N_2499,In_280,In_1301);
nand U2500 (N_2500,In_1190,In_1154);
or U2501 (N_2501,In_1185,In_1435);
nand U2502 (N_2502,In_1275,In_290);
nor U2503 (N_2503,In_326,In_710);
and U2504 (N_2504,In_38,In_788);
or U2505 (N_2505,In_902,In_1115);
and U2506 (N_2506,In_784,In_1354);
and U2507 (N_2507,In_795,In_1204);
xnor U2508 (N_2508,In_1310,In_362);
and U2509 (N_2509,In_199,In_108);
nand U2510 (N_2510,In_1103,In_285);
xor U2511 (N_2511,In_1356,In_1360);
and U2512 (N_2512,In_433,In_266);
nand U2513 (N_2513,In_1348,In_800);
nor U2514 (N_2514,In_192,In_373);
and U2515 (N_2515,In_1174,In_1277);
xnor U2516 (N_2516,In_408,In_538);
and U2517 (N_2517,In_851,In_1190);
or U2518 (N_2518,In_1368,In_1451);
or U2519 (N_2519,In_148,In_1475);
and U2520 (N_2520,In_682,In_252);
nor U2521 (N_2521,In_223,In_1123);
nand U2522 (N_2522,In_443,In_1224);
xnor U2523 (N_2523,In_791,In_773);
xnor U2524 (N_2524,In_540,In_178);
and U2525 (N_2525,In_842,In_97);
xnor U2526 (N_2526,In_258,In_942);
or U2527 (N_2527,In_161,In_1062);
and U2528 (N_2528,In_51,In_0);
and U2529 (N_2529,In_1360,In_381);
xnor U2530 (N_2530,In_257,In_8);
xnor U2531 (N_2531,In_1034,In_160);
nor U2532 (N_2532,In_353,In_583);
or U2533 (N_2533,In_836,In_569);
nand U2534 (N_2534,In_1331,In_1178);
xnor U2535 (N_2535,In_1213,In_1136);
xor U2536 (N_2536,In_1229,In_442);
and U2537 (N_2537,In_534,In_78);
and U2538 (N_2538,In_669,In_62);
and U2539 (N_2539,In_1489,In_1273);
nor U2540 (N_2540,In_210,In_5);
nand U2541 (N_2541,In_360,In_475);
xnor U2542 (N_2542,In_1470,In_71);
nand U2543 (N_2543,In_1198,In_369);
xnor U2544 (N_2544,In_1289,In_371);
and U2545 (N_2545,In_1110,In_295);
nand U2546 (N_2546,In_963,In_416);
nand U2547 (N_2547,In_29,In_828);
nor U2548 (N_2548,In_1280,In_1030);
nand U2549 (N_2549,In_86,In_608);
nor U2550 (N_2550,In_514,In_836);
xor U2551 (N_2551,In_1417,In_761);
xnor U2552 (N_2552,In_25,In_211);
nand U2553 (N_2553,In_734,In_551);
and U2554 (N_2554,In_578,In_1316);
nand U2555 (N_2555,In_1498,In_246);
nand U2556 (N_2556,In_1462,In_823);
and U2557 (N_2557,In_253,In_1260);
and U2558 (N_2558,In_257,In_1282);
nor U2559 (N_2559,In_1003,In_596);
xnor U2560 (N_2560,In_1183,In_451);
and U2561 (N_2561,In_1272,In_867);
nor U2562 (N_2562,In_326,In_102);
nor U2563 (N_2563,In_1152,In_1053);
xnor U2564 (N_2564,In_394,In_1245);
and U2565 (N_2565,In_1398,In_786);
nand U2566 (N_2566,In_806,In_845);
xor U2567 (N_2567,In_1443,In_649);
nor U2568 (N_2568,In_1474,In_826);
xor U2569 (N_2569,In_1328,In_666);
and U2570 (N_2570,In_1065,In_1164);
and U2571 (N_2571,In_1214,In_466);
nor U2572 (N_2572,In_137,In_823);
and U2573 (N_2573,In_1247,In_860);
and U2574 (N_2574,In_1393,In_1207);
nand U2575 (N_2575,In_950,In_670);
or U2576 (N_2576,In_1036,In_188);
xnor U2577 (N_2577,In_986,In_603);
or U2578 (N_2578,In_806,In_838);
xnor U2579 (N_2579,In_457,In_42);
and U2580 (N_2580,In_477,In_352);
xor U2581 (N_2581,In_194,In_790);
and U2582 (N_2582,In_247,In_820);
and U2583 (N_2583,In_194,In_1405);
and U2584 (N_2584,In_599,In_603);
nor U2585 (N_2585,In_415,In_264);
xnor U2586 (N_2586,In_132,In_668);
xor U2587 (N_2587,In_387,In_79);
and U2588 (N_2588,In_292,In_1129);
or U2589 (N_2589,In_132,In_922);
or U2590 (N_2590,In_1275,In_86);
nand U2591 (N_2591,In_1249,In_1048);
xor U2592 (N_2592,In_1151,In_351);
or U2593 (N_2593,In_1017,In_1229);
and U2594 (N_2594,In_493,In_351);
nand U2595 (N_2595,In_561,In_403);
nand U2596 (N_2596,In_1167,In_184);
or U2597 (N_2597,In_993,In_549);
and U2598 (N_2598,In_1326,In_46);
or U2599 (N_2599,In_235,In_403);
nor U2600 (N_2600,In_60,In_896);
and U2601 (N_2601,In_591,In_1164);
nand U2602 (N_2602,In_7,In_1444);
nor U2603 (N_2603,In_120,In_1379);
or U2604 (N_2604,In_645,In_1352);
and U2605 (N_2605,In_827,In_284);
xnor U2606 (N_2606,In_620,In_1295);
or U2607 (N_2607,In_28,In_671);
nor U2608 (N_2608,In_998,In_532);
and U2609 (N_2609,In_327,In_904);
nand U2610 (N_2610,In_586,In_761);
or U2611 (N_2611,In_102,In_202);
nand U2612 (N_2612,In_1220,In_1432);
xor U2613 (N_2613,In_918,In_1115);
and U2614 (N_2614,In_79,In_937);
nand U2615 (N_2615,In_1314,In_313);
and U2616 (N_2616,In_1275,In_931);
nand U2617 (N_2617,In_232,In_637);
nor U2618 (N_2618,In_436,In_773);
or U2619 (N_2619,In_215,In_95);
or U2620 (N_2620,In_220,In_411);
xnor U2621 (N_2621,In_1332,In_201);
and U2622 (N_2622,In_267,In_570);
nor U2623 (N_2623,In_637,In_1192);
and U2624 (N_2624,In_619,In_983);
xnor U2625 (N_2625,In_905,In_1482);
and U2626 (N_2626,In_673,In_1354);
and U2627 (N_2627,In_632,In_592);
nor U2628 (N_2628,In_1046,In_647);
and U2629 (N_2629,In_876,In_1371);
nor U2630 (N_2630,In_316,In_1468);
nand U2631 (N_2631,In_429,In_953);
and U2632 (N_2632,In_28,In_475);
or U2633 (N_2633,In_662,In_537);
xnor U2634 (N_2634,In_1313,In_1268);
nor U2635 (N_2635,In_903,In_1469);
nor U2636 (N_2636,In_4,In_463);
nor U2637 (N_2637,In_1281,In_916);
or U2638 (N_2638,In_1446,In_1449);
nor U2639 (N_2639,In_1110,In_665);
or U2640 (N_2640,In_1215,In_133);
nor U2641 (N_2641,In_1260,In_1004);
xnor U2642 (N_2642,In_1162,In_784);
xor U2643 (N_2643,In_375,In_1085);
nor U2644 (N_2644,In_979,In_216);
or U2645 (N_2645,In_1240,In_1332);
nor U2646 (N_2646,In_103,In_1469);
nand U2647 (N_2647,In_1321,In_425);
nand U2648 (N_2648,In_349,In_182);
or U2649 (N_2649,In_1162,In_30);
xnor U2650 (N_2650,In_1308,In_56);
or U2651 (N_2651,In_676,In_652);
nor U2652 (N_2652,In_68,In_526);
nand U2653 (N_2653,In_470,In_140);
xnor U2654 (N_2654,In_392,In_908);
nand U2655 (N_2655,In_93,In_1173);
xor U2656 (N_2656,In_212,In_792);
xnor U2657 (N_2657,In_1396,In_387);
nand U2658 (N_2658,In_1220,In_1214);
or U2659 (N_2659,In_1465,In_438);
or U2660 (N_2660,In_988,In_112);
nor U2661 (N_2661,In_930,In_1490);
and U2662 (N_2662,In_841,In_782);
xor U2663 (N_2663,In_597,In_385);
nor U2664 (N_2664,In_1043,In_235);
or U2665 (N_2665,In_221,In_965);
nand U2666 (N_2666,In_231,In_1036);
nand U2667 (N_2667,In_718,In_1404);
or U2668 (N_2668,In_935,In_160);
nor U2669 (N_2669,In_1367,In_308);
nor U2670 (N_2670,In_387,In_626);
xor U2671 (N_2671,In_387,In_464);
nor U2672 (N_2672,In_775,In_40);
nand U2673 (N_2673,In_634,In_349);
and U2674 (N_2674,In_735,In_602);
xor U2675 (N_2675,In_522,In_42);
nor U2676 (N_2676,In_33,In_705);
nand U2677 (N_2677,In_1082,In_733);
nor U2678 (N_2678,In_823,In_1004);
or U2679 (N_2679,In_74,In_329);
nor U2680 (N_2680,In_976,In_536);
or U2681 (N_2681,In_1007,In_1303);
xnor U2682 (N_2682,In_1276,In_1327);
xor U2683 (N_2683,In_63,In_412);
or U2684 (N_2684,In_950,In_574);
nor U2685 (N_2685,In_1003,In_1469);
and U2686 (N_2686,In_106,In_1467);
nor U2687 (N_2687,In_621,In_1184);
nor U2688 (N_2688,In_1172,In_365);
xor U2689 (N_2689,In_295,In_386);
nor U2690 (N_2690,In_227,In_885);
and U2691 (N_2691,In_42,In_637);
and U2692 (N_2692,In_997,In_523);
or U2693 (N_2693,In_846,In_323);
nand U2694 (N_2694,In_699,In_1395);
xnor U2695 (N_2695,In_1075,In_1456);
and U2696 (N_2696,In_289,In_1100);
xnor U2697 (N_2697,In_1134,In_830);
nand U2698 (N_2698,In_645,In_156);
xnor U2699 (N_2699,In_301,In_1257);
xnor U2700 (N_2700,In_1413,In_1283);
nor U2701 (N_2701,In_815,In_926);
nor U2702 (N_2702,In_765,In_771);
xor U2703 (N_2703,In_1269,In_770);
or U2704 (N_2704,In_1460,In_812);
or U2705 (N_2705,In_405,In_383);
xnor U2706 (N_2706,In_753,In_1338);
and U2707 (N_2707,In_507,In_50);
nor U2708 (N_2708,In_481,In_558);
xor U2709 (N_2709,In_1067,In_965);
nor U2710 (N_2710,In_815,In_527);
xnor U2711 (N_2711,In_291,In_702);
nand U2712 (N_2712,In_53,In_658);
nor U2713 (N_2713,In_1456,In_332);
xnor U2714 (N_2714,In_604,In_583);
and U2715 (N_2715,In_1181,In_14);
nand U2716 (N_2716,In_162,In_1277);
and U2717 (N_2717,In_1269,In_147);
and U2718 (N_2718,In_1367,In_792);
and U2719 (N_2719,In_1128,In_535);
nand U2720 (N_2720,In_217,In_396);
and U2721 (N_2721,In_809,In_843);
xnor U2722 (N_2722,In_1101,In_254);
xor U2723 (N_2723,In_285,In_1372);
nand U2724 (N_2724,In_516,In_1130);
and U2725 (N_2725,In_1465,In_590);
and U2726 (N_2726,In_419,In_1417);
nor U2727 (N_2727,In_1366,In_376);
nor U2728 (N_2728,In_673,In_995);
xnor U2729 (N_2729,In_611,In_584);
nor U2730 (N_2730,In_959,In_1027);
or U2731 (N_2731,In_1036,In_191);
and U2732 (N_2732,In_1443,In_0);
or U2733 (N_2733,In_1381,In_368);
nand U2734 (N_2734,In_1286,In_1168);
and U2735 (N_2735,In_1190,In_946);
nand U2736 (N_2736,In_1331,In_999);
xor U2737 (N_2737,In_580,In_531);
and U2738 (N_2738,In_672,In_611);
nand U2739 (N_2739,In_208,In_23);
and U2740 (N_2740,In_294,In_698);
and U2741 (N_2741,In_1081,In_1147);
or U2742 (N_2742,In_729,In_751);
nor U2743 (N_2743,In_682,In_442);
nand U2744 (N_2744,In_1495,In_638);
nand U2745 (N_2745,In_953,In_1282);
and U2746 (N_2746,In_474,In_1431);
and U2747 (N_2747,In_233,In_1119);
xor U2748 (N_2748,In_916,In_651);
xor U2749 (N_2749,In_1119,In_241);
nand U2750 (N_2750,In_1219,In_831);
nor U2751 (N_2751,In_1495,In_816);
or U2752 (N_2752,In_472,In_439);
nor U2753 (N_2753,In_700,In_790);
nor U2754 (N_2754,In_1298,In_324);
or U2755 (N_2755,In_1072,In_583);
nand U2756 (N_2756,In_1494,In_41);
or U2757 (N_2757,In_629,In_1051);
or U2758 (N_2758,In_643,In_953);
and U2759 (N_2759,In_1238,In_458);
nor U2760 (N_2760,In_983,In_691);
nand U2761 (N_2761,In_1106,In_1490);
or U2762 (N_2762,In_165,In_1254);
nor U2763 (N_2763,In_361,In_672);
xnor U2764 (N_2764,In_1386,In_10);
xnor U2765 (N_2765,In_132,In_94);
and U2766 (N_2766,In_944,In_169);
nor U2767 (N_2767,In_726,In_430);
nor U2768 (N_2768,In_185,In_378);
nand U2769 (N_2769,In_477,In_1490);
xnor U2770 (N_2770,In_1432,In_510);
or U2771 (N_2771,In_862,In_716);
nor U2772 (N_2772,In_847,In_854);
or U2773 (N_2773,In_1213,In_1298);
nand U2774 (N_2774,In_873,In_1205);
or U2775 (N_2775,In_1,In_345);
and U2776 (N_2776,In_391,In_235);
nor U2777 (N_2777,In_968,In_1465);
nor U2778 (N_2778,In_236,In_1157);
xnor U2779 (N_2779,In_648,In_653);
or U2780 (N_2780,In_865,In_106);
or U2781 (N_2781,In_261,In_174);
and U2782 (N_2782,In_1054,In_50);
or U2783 (N_2783,In_630,In_818);
and U2784 (N_2784,In_118,In_1386);
and U2785 (N_2785,In_834,In_557);
nand U2786 (N_2786,In_386,In_1108);
or U2787 (N_2787,In_521,In_914);
xor U2788 (N_2788,In_903,In_523);
nor U2789 (N_2789,In_1431,In_61);
and U2790 (N_2790,In_478,In_1103);
or U2791 (N_2791,In_138,In_1407);
nand U2792 (N_2792,In_496,In_361);
xor U2793 (N_2793,In_897,In_49);
xor U2794 (N_2794,In_1002,In_1039);
and U2795 (N_2795,In_1392,In_1118);
or U2796 (N_2796,In_9,In_1433);
nor U2797 (N_2797,In_892,In_611);
nand U2798 (N_2798,In_114,In_1497);
nor U2799 (N_2799,In_1478,In_812);
and U2800 (N_2800,In_765,In_690);
or U2801 (N_2801,In_974,In_1013);
and U2802 (N_2802,In_667,In_1473);
nor U2803 (N_2803,In_1227,In_421);
nand U2804 (N_2804,In_1239,In_337);
xor U2805 (N_2805,In_314,In_649);
nand U2806 (N_2806,In_1046,In_559);
nand U2807 (N_2807,In_467,In_284);
xor U2808 (N_2808,In_1262,In_1010);
and U2809 (N_2809,In_543,In_1247);
nor U2810 (N_2810,In_1496,In_1157);
or U2811 (N_2811,In_138,In_1300);
nor U2812 (N_2812,In_1448,In_162);
or U2813 (N_2813,In_823,In_91);
xor U2814 (N_2814,In_319,In_295);
or U2815 (N_2815,In_1109,In_889);
xor U2816 (N_2816,In_1008,In_461);
xor U2817 (N_2817,In_991,In_1416);
nor U2818 (N_2818,In_798,In_444);
nand U2819 (N_2819,In_896,In_207);
xor U2820 (N_2820,In_1144,In_143);
or U2821 (N_2821,In_1306,In_971);
and U2822 (N_2822,In_969,In_738);
nor U2823 (N_2823,In_652,In_894);
xor U2824 (N_2824,In_444,In_583);
xnor U2825 (N_2825,In_454,In_929);
xnor U2826 (N_2826,In_37,In_623);
nor U2827 (N_2827,In_1223,In_167);
xnor U2828 (N_2828,In_910,In_132);
nor U2829 (N_2829,In_1202,In_924);
and U2830 (N_2830,In_355,In_899);
xnor U2831 (N_2831,In_1470,In_1050);
or U2832 (N_2832,In_264,In_616);
nor U2833 (N_2833,In_352,In_353);
nand U2834 (N_2834,In_524,In_358);
or U2835 (N_2835,In_208,In_480);
xor U2836 (N_2836,In_960,In_417);
and U2837 (N_2837,In_714,In_984);
or U2838 (N_2838,In_1075,In_931);
nand U2839 (N_2839,In_172,In_1347);
nor U2840 (N_2840,In_26,In_96);
and U2841 (N_2841,In_473,In_678);
xor U2842 (N_2842,In_19,In_264);
nand U2843 (N_2843,In_365,In_670);
nor U2844 (N_2844,In_400,In_478);
or U2845 (N_2845,In_184,In_1239);
or U2846 (N_2846,In_160,In_410);
nand U2847 (N_2847,In_265,In_919);
nand U2848 (N_2848,In_711,In_676);
and U2849 (N_2849,In_1365,In_334);
and U2850 (N_2850,In_246,In_515);
and U2851 (N_2851,In_1253,In_609);
nand U2852 (N_2852,In_186,In_742);
xnor U2853 (N_2853,In_999,In_290);
or U2854 (N_2854,In_1097,In_1077);
xor U2855 (N_2855,In_214,In_995);
nand U2856 (N_2856,In_1163,In_709);
or U2857 (N_2857,In_186,In_0);
nand U2858 (N_2858,In_173,In_987);
nor U2859 (N_2859,In_717,In_1043);
nor U2860 (N_2860,In_990,In_795);
nand U2861 (N_2861,In_533,In_663);
and U2862 (N_2862,In_675,In_151);
nand U2863 (N_2863,In_1438,In_1352);
xor U2864 (N_2864,In_71,In_1423);
and U2865 (N_2865,In_845,In_1083);
nor U2866 (N_2866,In_1236,In_1198);
and U2867 (N_2867,In_1409,In_958);
nand U2868 (N_2868,In_1195,In_96);
or U2869 (N_2869,In_925,In_1274);
nor U2870 (N_2870,In_291,In_864);
nand U2871 (N_2871,In_53,In_850);
nand U2872 (N_2872,In_339,In_556);
nand U2873 (N_2873,In_566,In_1357);
nand U2874 (N_2874,In_81,In_855);
or U2875 (N_2875,In_637,In_797);
and U2876 (N_2876,In_1308,In_51);
nand U2877 (N_2877,In_905,In_1117);
xor U2878 (N_2878,In_540,In_680);
and U2879 (N_2879,In_930,In_1225);
or U2880 (N_2880,In_1027,In_1332);
or U2881 (N_2881,In_1207,In_543);
xor U2882 (N_2882,In_1116,In_1413);
and U2883 (N_2883,In_611,In_953);
nand U2884 (N_2884,In_1228,In_1460);
xnor U2885 (N_2885,In_815,In_746);
or U2886 (N_2886,In_360,In_1474);
or U2887 (N_2887,In_137,In_735);
xnor U2888 (N_2888,In_72,In_467);
xnor U2889 (N_2889,In_534,In_686);
nor U2890 (N_2890,In_854,In_1424);
and U2891 (N_2891,In_1282,In_800);
nand U2892 (N_2892,In_154,In_475);
and U2893 (N_2893,In_558,In_847);
nor U2894 (N_2894,In_997,In_1047);
or U2895 (N_2895,In_1151,In_1327);
or U2896 (N_2896,In_1036,In_1293);
or U2897 (N_2897,In_48,In_159);
xnor U2898 (N_2898,In_666,In_1389);
nor U2899 (N_2899,In_754,In_68);
xnor U2900 (N_2900,In_1278,In_576);
and U2901 (N_2901,In_229,In_84);
nand U2902 (N_2902,In_543,In_934);
nand U2903 (N_2903,In_301,In_511);
nor U2904 (N_2904,In_526,In_729);
nand U2905 (N_2905,In_1153,In_919);
xor U2906 (N_2906,In_835,In_7);
and U2907 (N_2907,In_900,In_1024);
nand U2908 (N_2908,In_373,In_1217);
nand U2909 (N_2909,In_880,In_845);
nand U2910 (N_2910,In_1121,In_1329);
and U2911 (N_2911,In_1239,In_1496);
and U2912 (N_2912,In_1366,In_1442);
nor U2913 (N_2913,In_709,In_473);
xor U2914 (N_2914,In_240,In_1202);
nor U2915 (N_2915,In_1472,In_1329);
nand U2916 (N_2916,In_547,In_979);
or U2917 (N_2917,In_122,In_338);
or U2918 (N_2918,In_746,In_1311);
nand U2919 (N_2919,In_899,In_1107);
or U2920 (N_2920,In_1014,In_1142);
or U2921 (N_2921,In_399,In_610);
xnor U2922 (N_2922,In_391,In_561);
nand U2923 (N_2923,In_158,In_1032);
or U2924 (N_2924,In_951,In_237);
and U2925 (N_2925,In_655,In_52);
or U2926 (N_2926,In_1182,In_1128);
nand U2927 (N_2927,In_540,In_856);
nor U2928 (N_2928,In_825,In_1039);
nand U2929 (N_2929,In_137,In_1082);
or U2930 (N_2930,In_686,In_130);
or U2931 (N_2931,In_1341,In_1292);
or U2932 (N_2932,In_703,In_1120);
xnor U2933 (N_2933,In_686,In_1179);
nor U2934 (N_2934,In_519,In_76);
nand U2935 (N_2935,In_1097,In_347);
xnor U2936 (N_2936,In_129,In_353);
and U2937 (N_2937,In_1408,In_281);
and U2938 (N_2938,In_859,In_227);
and U2939 (N_2939,In_1369,In_211);
nand U2940 (N_2940,In_1405,In_722);
nand U2941 (N_2941,In_1013,In_956);
xnor U2942 (N_2942,In_1023,In_920);
nand U2943 (N_2943,In_230,In_1012);
nor U2944 (N_2944,In_680,In_513);
nand U2945 (N_2945,In_842,In_105);
nand U2946 (N_2946,In_757,In_373);
nand U2947 (N_2947,In_1118,In_1138);
xnor U2948 (N_2948,In_585,In_278);
and U2949 (N_2949,In_1260,In_888);
nor U2950 (N_2950,In_1154,In_109);
xnor U2951 (N_2951,In_212,In_859);
xnor U2952 (N_2952,In_236,In_1466);
and U2953 (N_2953,In_1026,In_20);
nand U2954 (N_2954,In_1395,In_953);
nand U2955 (N_2955,In_526,In_1131);
xor U2956 (N_2956,In_990,In_1209);
xor U2957 (N_2957,In_667,In_1192);
nand U2958 (N_2958,In_579,In_1069);
or U2959 (N_2959,In_1262,In_1191);
or U2960 (N_2960,In_1297,In_178);
or U2961 (N_2961,In_1224,In_580);
nand U2962 (N_2962,In_1318,In_1226);
nand U2963 (N_2963,In_1362,In_554);
or U2964 (N_2964,In_1246,In_922);
xnor U2965 (N_2965,In_1422,In_1333);
nor U2966 (N_2966,In_989,In_1131);
xor U2967 (N_2967,In_1372,In_1409);
and U2968 (N_2968,In_45,In_709);
nand U2969 (N_2969,In_206,In_621);
nand U2970 (N_2970,In_368,In_134);
nand U2971 (N_2971,In_731,In_1028);
or U2972 (N_2972,In_1068,In_1455);
nor U2973 (N_2973,In_87,In_159);
and U2974 (N_2974,In_776,In_1193);
nand U2975 (N_2975,In_554,In_1049);
nor U2976 (N_2976,In_1019,In_1362);
nand U2977 (N_2977,In_572,In_210);
and U2978 (N_2978,In_394,In_638);
and U2979 (N_2979,In_337,In_566);
xor U2980 (N_2980,In_1300,In_206);
or U2981 (N_2981,In_310,In_38);
nand U2982 (N_2982,In_939,In_964);
nand U2983 (N_2983,In_1285,In_312);
and U2984 (N_2984,In_1404,In_542);
xnor U2985 (N_2985,In_551,In_1122);
xnor U2986 (N_2986,In_642,In_1437);
or U2987 (N_2987,In_383,In_825);
xor U2988 (N_2988,In_241,In_847);
nand U2989 (N_2989,In_405,In_896);
and U2990 (N_2990,In_643,In_183);
and U2991 (N_2991,In_1083,In_1424);
nor U2992 (N_2992,In_99,In_1499);
and U2993 (N_2993,In_926,In_1285);
nor U2994 (N_2994,In_417,In_361);
nand U2995 (N_2995,In_82,In_383);
xnor U2996 (N_2996,In_959,In_1451);
and U2997 (N_2997,In_907,In_222);
nor U2998 (N_2998,In_796,In_1248);
nor U2999 (N_2999,In_512,In_1484);
xnor U3000 (N_3000,N_1470,N_928);
nand U3001 (N_3001,N_1501,N_2593);
xor U3002 (N_3002,N_1107,N_854);
or U3003 (N_3003,N_1607,N_2494);
and U3004 (N_3004,N_896,N_186);
and U3005 (N_3005,N_1329,N_2290);
nand U3006 (N_3006,N_1478,N_1512);
nand U3007 (N_3007,N_339,N_2533);
nor U3008 (N_3008,N_465,N_1833);
and U3009 (N_3009,N_894,N_1580);
xnor U3010 (N_3010,N_2824,N_964);
and U3011 (N_3011,N_1727,N_2259);
nand U3012 (N_3012,N_114,N_772);
nor U3013 (N_3013,N_2847,N_1691);
and U3014 (N_3014,N_2811,N_788);
and U3015 (N_3015,N_192,N_1369);
or U3016 (N_3016,N_1779,N_2237);
or U3017 (N_3017,N_1586,N_1170);
nand U3018 (N_3018,N_2115,N_1150);
nand U3019 (N_3019,N_1790,N_481);
and U3020 (N_3020,N_1886,N_2429);
and U3021 (N_3021,N_2686,N_793);
nor U3022 (N_3022,N_2222,N_127);
nand U3023 (N_3023,N_2634,N_920);
nand U3024 (N_3024,N_2372,N_1022);
nor U3025 (N_3025,N_2940,N_446);
or U3026 (N_3026,N_852,N_1915);
nand U3027 (N_3027,N_2487,N_662);
xnor U3028 (N_3028,N_2488,N_840);
and U3029 (N_3029,N_2955,N_2101);
or U3030 (N_3030,N_2961,N_783);
xnor U3031 (N_3031,N_1422,N_439);
or U3032 (N_3032,N_1386,N_2774);
nand U3033 (N_3033,N_194,N_727);
xnor U3034 (N_3034,N_2716,N_1489);
or U3035 (N_3035,N_8,N_2854);
xnor U3036 (N_3036,N_257,N_137);
nand U3037 (N_3037,N_283,N_1967);
nor U3038 (N_3038,N_1947,N_2310);
xnor U3039 (N_3039,N_897,N_2345);
nand U3040 (N_3040,N_2951,N_364);
nor U3041 (N_3041,N_1785,N_131);
xor U3042 (N_3042,N_2668,N_2631);
xor U3043 (N_3043,N_948,N_1709);
or U3044 (N_3044,N_246,N_2515);
nor U3045 (N_3045,N_1866,N_1415);
nand U3046 (N_3046,N_1941,N_13);
xnor U3047 (N_3047,N_2540,N_2053);
xnor U3048 (N_3048,N_1961,N_2689);
nor U3049 (N_3049,N_1867,N_904);
nor U3050 (N_3050,N_559,N_2097);
nor U3051 (N_3051,N_2519,N_975);
xnor U3052 (N_3052,N_1364,N_2470);
xor U3053 (N_3053,N_682,N_1603);
and U3054 (N_3054,N_678,N_1495);
nor U3055 (N_3055,N_947,N_1493);
or U3056 (N_3056,N_1793,N_926);
and U3057 (N_3057,N_537,N_667);
xor U3058 (N_3058,N_2830,N_202);
xor U3059 (N_3059,N_2085,N_832);
nand U3060 (N_3060,N_2428,N_277);
or U3061 (N_3061,N_2850,N_1417);
or U3062 (N_3062,N_1815,N_891);
and U3063 (N_3063,N_1678,N_542);
xnor U3064 (N_3064,N_1176,N_1774);
and U3065 (N_3065,N_2625,N_800);
nand U3066 (N_3066,N_1046,N_493);
xnor U3067 (N_3067,N_2321,N_280);
and U3068 (N_3068,N_2495,N_2232);
and U3069 (N_3069,N_549,N_2814);
xor U3070 (N_3070,N_922,N_1572);
nand U3071 (N_3071,N_744,N_2558);
or U3072 (N_3072,N_1756,N_2045);
nand U3073 (N_3073,N_1058,N_961);
or U3074 (N_3074,N_1716,N_2245);
nor U3075 (N_3075,N_2159,N_63);
or U3076 (N_3076,N_2818,N_1073);
nand U3077 (N_3077,N_478,N_1085);
xor U3078 (N_3078,N_750,N_123);
xor U3079 (N_3079,N_607,N_1304);
xor U3080 (N_3080,N_847,N_1506);
and U3081 (N_3081,N_201,N_801);
nor U3082 (N_3082,N_1248,N_2144);
xnor U3083 (N_3083,N_1281,N_1735);
nand U3084 (N_3084,N_1582,N_2160);
and U3085 (N_3085,N_142,N_468);
xor U3086 (N_3086,N_1570,N_424);
nand U3087 (N_3087,N_291,N_2279);
and U3088 (N_3088,N_370,N_554);
xnor U3089 (N_3089,N_2147,N_1340);
nor U3090 (N_3090,N_398,N_511);
and U3091 (N_3091,N_787,N_634);
or U3092 (N_3092,N_2369,N_1623);
xnor U3093 (N_3093,N_1261,N_1410);
nor U3094 (N_3094,N_2141,N_617);
nand U3095 (N_3095,N_2435,N_1724);
nand U3096 (N_3096,N_668,N_2441);
and U3097 (N_3097,N_2808,N_303);
and U3098 (N_3098,N_2229,N_818);
or U3099 (N_3099,N_1347,N_409);
xor U3100 (N_3100,N_2535,N_2082);
nand U3101 (N_3101,N_2303,N_1646);
xnor U3102 (N_3102,N_1579,N_2354);
and U3103 (N_3103,N_1097,N_2623);
or U3104 (N_3104,N_1042,N_2296);
or U3105 (N_3105,N_2035,N_73);
and U3106 (N_3106,N_19,N_1481);
xor U3107 (N_3107,N_1882,N_2282);
xnor U3108 (N_3108,N_2554,N_82);
nor U3109 (N_3109,N_1492,N_2556);
xor U3110 (N_3110,N_701,N_1523);
xnor U3111 (N_3111,N_376,N_2460);
or U3112 (N_3112,N_429,N_2718);
nor U3113 (N_3113,N_1153,N_168);
and U3114 (N_3114,N_1426,N_1794);
and U3115 (N_3115,N_2327,N_2105);
nor U3116 (N_3116,N_785,N_1970);
nor U3117 (N_3117,N_1801,N_2944);
and U3118 (N_3118,N_1126,N_1302);
and U3119 (N_3119,N_1745,N_942);
nor U3120 (N_3120,N_1662,N_1462);
and U3121 (N_3121,N_1902,N_2498);
nand U3122 (N_3122,N_2373,N_2083);
or U3123 (N_3123,N_2236,N_2063);
or U3124 (N_3124,N_2520,N_2061);
nand U3125 (N_3125,N_872,N_1036);
and U3126 (N_3126,N_2760,N_2189);
nor U3127 (N_3127,N_2763,N_2611);
nor U3128 (N_3128,N_1389,N_2953);
and U3129 (N_3129,N_455,N_599);
nand U3130 (N_3130,N_284,N_865);
nand U3131 (N_3131,N_1697,N_2306);
nor U3132 (N_3132,N_641,N_766);
xor U3133 (N_3133,N_1013,N_1968);
xnor U3134 (N_3134,N_2761,N_765);
xnor U3135 (N_3135,N_1002,N_1577);
nand U3136 (N_3136,N_2234,N_987);
nor U3137 (N_3137,N_2564,N_677);
xor U3138 (N_3138,N_1513,N_1247);
and U3139 (N_3139,N_1676,N_2071);
or U3140 (N_3140,N_2208,N_1589);
nor U3141 (N_3141,N_2162,N_1154);
nand U3142 (N_3142,N_2813,N_2375);
nor U3143 (N_3143,N_1445,N_2052);
or U3144 (N_3144,N_2870,N_479);
nor U3145 (N_3145,N_1590,N_68);
nor U3146 (N_3146,N_2251,N_2644);
nor U3147 (N_3147,N_999,N_1475);
nor U3148 (N_3148,N_1411,N_2243);
xor U3149 (N_3149,N_567,N_2902);
nand U3150 (N_3150,N_2295,N_2650);
or U3151 (N_3151,N_1904,N_2202);
or U3152 (N_3152,N_1711,N_440);
xor U3153 (N_3153,N_1357,N_2181);
nor U3154 (N_3154,N_445,N_2945);
xnor U3155 (N_3155,N_2527,N_585);
or U3156 (N_3156,N_2575,N_1230);
nand U3157 (N_3157,N_531,N_2578);
nand U3158 (N_3158,N_2649,N_2696);
or U3159 (N_3159,N_1224,N_2618);
or U3160 (N_3160,N_2167,N_1219);
or U3161 (N_3161,N_2797,N_1373);
and U3162 (N_3162,N_1504,N_130);
nand U3163 (N_3163,N_1124,N_688);
nor U3164 (N_3164,N_2472,N_331);
nand U3165 (N_3165,N_1121,N_2285);
xnor U3166 (N_3166,N_1100,N_2415);
nand U3167 (N_3167,N_2842,N_1522);
and U3168 (N_3168,N_2687,N_372);
nand U3169 (N_3169,N_1959,N_1356);
nand U3170 (N_3170,N_516,N_2614);
and U3171 (N_3171,N_1976,N_839);
or U3172 (N_3172,N_2276,N_1909);
nand U3173 (N_3173,N_2709,N_2802);
or U3174 (N_3174,N_1051,N_391);
or U3175 (N_3175,N_1682,N_288);
and U3176 (N_3176,N_1378,N_1510);
nor U3177 (N_3177,N_1893,N_914);
xnor U3178 (N_3178,N_855,N_1898);
nor U3179 (N_3179,N_1458,N_2198);
nor U3180 (N_3180,N_1050,N_721);
and U3181 (N_3181,N_2499,N_714);
nand U3182 (N_3182,N_2673,N_2371);
or U3183 (N_3183,N_33,N_2021);
nor U3184 (N_3184,N_1116,N_673);
or U3185 (N_3185,N_204,N_230);
nor U3186 (N_3186,N_2133,N_2806);
and U3187 (N_3187,N_1158,N_2734);
and U3188 (N_3188,N_2901,N_960);
nand U3189 (N_3189,N_2672,N_2065);
and U3190 (N_3190,N_93,N_48);
xnor U3191 (N_3191,N_2466,N_720);
xor U3192 (N_3192,N_2148,N_1529);
xnor U3193 (N_3193,N_1675,N_2597);
and U3194 (N_3194,N_527,N_2359);
nor U3195 (N_3195,N_2778,N_1640);
xor U3196 (N_3196,N_2370,N_2586);
or U3197 (N_3197,N_1317,N_2240);
and U3198 (N_3198,N_135,N_1811);
and U3199 (N_3199,N_1459,N_2989);
nor U3200 (N_3200,N_162,N_546);
nand U3201 (N_3201,N_2538,N_133);
xnor U3202 (N_3202,N_1279,N_524);
or U3203 (N_3203,N_2723,N_2308);
nand U3204 (N_3204,N_1943,N_301);
xor U3205 (N_3205,N_341,N_562);
nor U3206 (N_3206,N_2403,N_1206);
xnor U3207 (N_3207,N_826,N_1635);
nor U3208 (N_3208,N_84,N_1249);
and U3209 (N_3209,N_706,N_320);
xnor U3210 (N_3210,N_2815,N_597);
nand U3211 (N_3211,N_1535,N_275);
or U3212 (N_3212,N_660,N_2084);
nand U3213 (N_3213,N_260,N_332);
nor U3214 (N_3214,N_1914,N_2023);
and U3215 (N_3215,N_2984,N_2637);
nor U3216 (N_3216,N_919,N_1533);
or U3217 (N_3217,N_53,N_1738);
nand U3218 (N_3218,N_2302,N_215);
nor U3219 (N_3219,N_427,N_1721);
xor U3220 (N_3220,N_2798,N_1026);
or U3221 (N_3221,N_1131,N_472);
nand U3222 (N_3222,N_1074,N_492);
xnor U3223 (N_3223,N_642,N_1268);
and U3224 (N_3224,N_2380,N_646);
or U3225 (N_3225,N_2246,N_880);
nor U3226 (N_3226,N_1986,N_1092);
nor U3227 (N_3227,N_984,N_694);
xnor U3228 (N_3228,N_1323,N_2338);
and U3229 (N_3229,N_1796,N_1425);
and U3230 (N_3230,N_1087,N_2534);
nor U3231 (N_3231,N_349,N_1578);
nand U3232 (N_3232,N_629,N_187);
nand U3233 (N_3233,N_1555,N_2343);
nor U3234 (N_3234,N_497,N_62);
nand U3235 (N_3235,N_595,N_2863);
xnor U3236 (N_3236,N_2486,N_217);
xnor U3237 (N_3237,N_778,N_1642);
xnor U3238 (N_3238,N_2217,N_944);
xnor U3239 (N_3239,N_2173,N_1521);
and U3240 (N_3240,N_1981,N_1985);
and U3241 (N_3241,N_1413,N_1692);
nand U3242 (N_3242,N_469,N_1838);
or U3243 (N_3243,N_739,N_868);
or U3244 (N_3244,N_1265,N_2081);
or U3245 (N_3245,N_271,N_823);
nand U3246 (N_3246,N_200,N_1044);
or U3247 (N_3247,N_146,N_2913);
nor U3248 (N_3248,N_181,N_536);
or U3249 (N_3249,N_154,N_1138);
nand U3250 (N_3250,N_659,N_611);
or U3251 (N_3251,N_2209,N_2925);
nor U3252 (N_3252,N_1146,N_2078);
or U3253 (N_3253,N_620,N_1250);
nand U3254 (N_3254,N_2465,N_2627);
or U3255 (N_3255,N_541,N_2670);
and U3256 (N_3256,N_1576,N_2393);
nor U3257 (N_3257,N_2107,N_2985);
nor U3258 (N_3258,N_2932,N_881);
nand U3259 (N_3259,N_767,N_875);
nand U3260 (N_3260,N_2005,N_2439);
and U3261 (N_3261,N_2665,N_426);
nor U3262 (N_3262,N_1343,N_2213);
or U3263 (N_3263,N_451,N_1958);
or U3264 (N_3264,N_2029,N_1220);
nor U3265 (N_3265,N_2032,N_2457);
or U3266 (N_3266,N_1924,N_2075);
xor U3267 (N_3267,N_965,N_582);
nor U3268 (N_3268,N_1132,N_1136);
and U3269 (N_3269,N_1665,N_794);
and U3270 (N_3270,N_1208,N_1229);
and U3271 (N_3271,N_2201,N_2312);
and U3272 (N_3272,N_705,N_980);
nand U3273 (N_3273,N_702,N_365);
nor U3274 (N_3274,N_864,N_38);
nor U3275 (N_3275,N_1012,N_25);
or U3276 (N_3276,N_2873,N_2390);
and U3277 (N_3277,N_1974,N_761);
or U3278 (N_3278,N_2292,N_1218);
nor U3279 (N_3279,N_300,N_1710);
nor U3280 (N_3280,N_2787,N_1911);
or U3281 (N_3281,N_1518,N_2469);
nor U3282 (N_3282,N_109,N_917);
nor U3283 (N_3283,N_1851,N_2579);
nor U3284 (N_3284,N_1753,N_1830);
nand U3285 (N_3285,N_2166,N_1877);
and U3286 (N_3286,N_1626,N_2658);
nor U3287 (N_3287,N_716,N_265);
nor U3288 (N_3288,N_722,N_1718);
xor U3289 (N_3289,N_1179,N_333);
nand U3290 (N_3290,N_105,N_1502);
nand U3291 (N_3291,N_2894,N_2377);
or U3292 (N_3292,N_625,N_462);
and U3293 (N_3293,N_2652,N_268);
nor U3294 (N_3294,N_2752,N_1729);
nand U3295 (N_3295,N_35,N_467);
or U3296 (N_3296,N_58,N_2777);
or U3297 (N_3297,N_657,N_2956);
nor U3298 (N_3298,N_1379,N_2108);
and U3299 (N_3299,N_976,N_278);
nand U3300 (N_3300,N_1029,N_2915);
xor U3301 (N_3301,N_1260,N_2361);
or U3302 (N_3302,N_1544,N_2746);
and U3303 (N_3303,N_46,N_247);
xnor U3304 (N_3304,N_1566,N_1883);
or U3305 (N_3305,N_2526,N_2930);
and U3306 (N_3306,N_1634,N_645);
xor U3307 (N_3307,N_1918,N_2230);
or U3308 (N_3308,N_590,N_790);
or U3309 (N_3309,N_208,N_406);
nand U3310 (N_3310,N_2187,N_1547);
xor U3311 (N_3311,N_2622,N_652);
and U3312 (N_3312,N_488,N_809);
xnor U3313 (N_3313,N_2699,N_1734);
or U3314 (N_3314,N_1203,N_547);
or U3315 (N_3315,N_2987,N_2514);
nand U3316 (N_3316,N_1172,N_1957);
xnor U3317 (N_3317,N_1795,N_2445);
or U3318 (N_3318,N_806,N_2911);
and U3319 (N_3319,N_1056,N_2907);
and U3320 (N_3320,N_2130,N_2799);
nor U3321 (N_3321,N_1617,N_2626);
and U3322 (N_3322,N_1420,N_2333);
xor U3323 (N_3323,N_464,N_2512);
and U3324 (N_3324,N_2730,N_2682);
or U3325 (N_3325,N_74,N_2205);
xnor U3326 (N_3326,N_182,N_423);
xor U3327 (N_3327,N_1820,N_780);
and U3328 (N_3328,N_1668,N_2161);
xnor U3329 (N_3329,N_1400,N_1066);
nor U3330 (N_3330,N_2381,N_2999);
nand U3331 (N_3331,N_1490,N_1856);
or U3332 (N_3332,N_1723,N_2825);
nand U3333 (N_3333,N_1631,N_2212);
nand U3334 (N_3334,N_1342,N_1696);
nand U3335 (N_3335,N_1977,N_2134);
nor U3336 (N_3336,N_656,N_1719);
nand U3337 (N_3337,N_2800,N_889);
nand U3338 (N_3338,N_2522,N_350);
or U3339 (N_3339,N_971,N_1892);
nand U3340 (N_3340,N_2153,N_458);
and U3341 (N_3341,N_405,N_1895);
nand U3342 (N_3342,N_1054,N_2753);
xor U3343 (N_3343,N_1949,N_2139);
xnor U3344 (N_3344,N_1139,N_1240);
or U3345 (N_3345,N_2566,N_388);
or U3346 (N_3346,N_1083,N_2386);
and U3347 (N_3347,N_1093,N_2553);
xnor U3348 (N_3348,N_2991,N_2829);
xnor U3349 (N_3349,N_615,N_1003);
or U3350 (N_3350,N_2170,N_1669);
nor U3351 (N_3351,N_658,N_1822);
nor U3352 (N_3352,N_2335,N_1848);
xnor U3353 (N_3353,N_250,N_266);
nor U3354 (N_3354,N_2507,N_2484);
and U3355 (N_3355,N_340,N_1464);
or U3356 (N_3356,N_1316,N_67);
or U3357 (N_3357,N_573,N_1468);
and U3358 (N_3358,N_401,N_2450);
xnor U3359 (N_3359,N_1060,N_2412);
xnor U3360 (N_3360,N_2104,N_1767);
and U3361 (N_3361,N_2404,N_1847);
nor U3362 (N_3362,N_251,N_893);
nor U3363 (N_3363,N_600,N_185);
nor U3364 (N_3364,N_59,N_962);
nor U3365 (N_3365,N_2549,N_1216);
xor U3366 (N_3366,N_1094,N_648);
xor U3367 (N_3367,N_444,N_95);
nand U3368 (N_3368,N_2031,N_403);
nor U3369 (N_3369,N_1466,N_1252);
nor U3370 (N_3370,N_2924,N_2529);
xor U3371 (N_3371,N_17,N_795);
nand U3372 (N_3372,N_1207,N_1587);
or U3373 (N_3373,N_680,N_2418);
and U3374 (N_3374,N_1913,N_1287);
xor U3375 (N_3375,N_2376,N_2118);
nor U3376 (N_3376,N_1430,N_2009);
and U3377 (N_3377,N_2272,N_2176);
and U3378 (N_3378,N_286,N_1780);
xnor U3379 (N_3379,N_1200,N_2040);
and U3380 (N_3380,N_1483,N_2794);
nor U3381 (N_3381,N_1602,N_501);
or U3382 (N_3382,N_1267,N_1887);
xor U3383 (N_3383,N_96,N_2643);
xnor U3384 (N_3384,N_2669,N_1749);
and U3385 (N_3385,N_2909,N_1402);
xnor U3386 (N_3386,N_1558,N_1648);
xor U3387 (N_3387,N_1568,N_639);
or U3388 (N_3388,N_2957,N_1188);
nand U3389 (N_3389,N_650,N_1407);
or U3390 (N_3390,N_718,N_1151);
nand U3391 (N_3391,N_1177,N_2655);
nand U3392 (N_3392,N_1872,N_326);
and U3393 (N_3393,N_1608,N_526);
and U3394 (N_3394,N_2250,N_129);
or U3395 (N_3395,N_2789,N_2890);
or U3396 (N_3396,N_1541,N_2523);
and U3397 (N_3397,N_1312,N_2536);
xor U3398 (N_3398,N_2452,N_1862);
xor U3399 (N_3399,N_2449,N_579);
xnor U3400 (N_3400,N_1186,N_770);
and U3401 (N_3401,N_1775,N_1409);
xnor U3402 (N_3402,N_2918,N_2776);
xnor U3403 (N_3403,N_564,N_776);
and U3404 (N_3404,N_282,N_2318);
nand U3405 (N_3405,N_294,N_2524);
nor U3406 (N_3406,N_2796,N_2378);
and U3407 (N_3407,N_972,N_2837);
nor U3408 (N_3408,N_654,N_2131);
nand U3409 (N_3409,N_1827,N_2066);
nand U3410 (N_3410,N_1078,N_2255);
nor U3411 (N_3411,N_1463,N_1601);
or U3412 (N_3412,N_2978,N_1987);
or U3413 (N_3413,N_671,N_1077);
nor U3414 (N_3414,N_1398,N_2966);
xor U3415 (N_3415,N_2064,N_784);
or U3416 (N_3416,N_1596,N_1108);
or U3417 (N_3417,N_2455,N_989);
nor U3418 (N_3418,N_2177,N_1556);
or U3419 (N_3419,N_489,N_1989);
or U3420 (N_3420,N_2417,N_2585);
nand U3421 (N_3421,N_2750,N_233);
or U3422 (N_3422,N_709,N_1182);
nand U3423 (N_3423,N_731,N_934);
nor U3424 (N_3424,N_329,N_2698);
and U3425 (N_3425,N_2152,N_65);
nor U3426 (N_3426,N_2478,N_1034);
nand U3427 (N_3427,N_2993,N_2490);
and U3428 (N_3428,N_1440,N_636);
xor U3429 (N_3429,N_2917,N_1931);
nor U3430 (N_3430,N_2633,N_2908);
nand U3431 (N_3431,N_1027,N_311);
and U3432 (N_3432,N_1704,N_2054);
xnor U3433 (N_3433,N_2897,N_1404);
nand U3434 (N_3434,N_463,N_1781);
and U3435 (N_3435,N_2119,N_2963);
xor U3436 (N_3436,N_64,N_2542);
nor U3437 (N_3437,N_955,N_12);
nand U3438 (N_3438,N_762,N_2392);
nor U3439 (N_3439,N_2283,N_1419);
or U3440 (N_3440,N_433,N_85);
or U3441 (N_3441,N_115,N_2352);
nand U3442 (N_3442,N_1303,N_2543);
nor U3443 (N_3443,N_1401,N_2977);
nand U3444 (N_3444,N_2431,N_245);
nor U3445 (N_3445,N_2679,N_1109);
nand U3446 (N_3446,N_1447,N_1246);
or U3447 (N_3447,N_846,N_1204);
nor U3448 (N_3448,N_155,N_1254);
or U3449 (N_3449,N_1000,N_2719);
or U3450 (N_3450,N_2659,N_385);
nor U3451 (N_3451,N_1543,N_2560);
nor U3452 (N_3452,N_106,N_1853);
and U3453 (N_3453,N_2812,N_2663);
nand U3454 (N_3454,N_1688,N_2122);
nor U3455 (N_3455,N_2297,N_1903);
and U3456 (N_3456,N_2459,N_44);
and U3457 (N_3457,N_2434,N_1198);
xnor U3458 (N_3458,N_726,N_907);
xnor U3459 (N_3459,N_1731,N_2771);
nor U3460 (N_3460,N_2326,N_1846);
nand U3461 (N_3461,N_102,N_2258);
nand U3462 (N_3462,N_995,N_1102);
or U3463 (N_3463,N_2442,N_1052);
xnor U3464 (N_3464,N_1612,N_2573);
xor U3465 (N_3465,N_2408,N_1751);
or U3466 (N_3466,N_2188,N_1199);
nand U3467 (N_3467,N_1449,N_1628);
or U3468 (N_3468,N_2155,N_1318);
or U3469 (N_3469,N_211,N_935);
xor U3470 (N_3470,N_1284,N_2934);
nand U3471 (N_3471,N_2299,N_812);
nor U3472 (N_3472,N_510,N_1406);
and U3473 (N_3473,N_2210,N_2142);
or U3474 (N_3474,N_363,N_1859);
or U3475 (N_3475,N_2982,N_2006);
xnor U3476 (N_3476,N_2454,N_1752);
or U3477 (N_3477,N_2601,N_36);
xnor U3478 (N_3478,N_2826,N_1212);
or U3479 (N_3479,N_378,N_1476);
nor U3480 (N_3480,N_2906,N_1591);
nor U3481 (N_3481,N_664,N_1333);
nand U3482 (N_3482,N_1484,N_1921);
and U3483 (N_3483,N_1414,N_570);
and U3484 (N_3484,N_2544,N_1714);
or U3485 (N_3485,N_2356,N_939);
nand U3486 (N_3486,N_2003,N_313);
and U3487 (N_3487,N_1004,N_111);
and U3488 (N_3488,N_814,N_475);
nand U3489 (N_3489,N_2595,N_2976);
or U3490 (N_3490,N_878,N_491);
or U3491 (N_3491,N_2904,N_1861);
and U3492 (N_3492,N_884,N_47);
and U3493 (N_3493,N_1485,N_2946);
nor U3494 (N_3494,N_2163,N_2015);
or U3495 (N_3495,N_343,N_849);
nand U3496 (N_3496,N_2717,N_687);
or U3497 (N_3497,N_1797,N_2583);
nand U3498 (N_3498,N_441,N_256);
and U3499 (N_3499,N_1538,N_2509);
and U3500 (N_3500,N_2671,N_906);
and U3501 (N_3501,N_2517,N_1906);
and U3502 (N_3502,N_2630,N_1605);
nand U3503 (N_3503,N_1244,N_1105);
xor U3504 (N_3504,N_2334,N_2056);
and U3505 (N_3505,N_993,N_2301);
xor U3506 (N_3506,N_1952,N_170);
nor U3507 (N_3507,N_2211,N_923);
xor U3508 (N_3508,N_1019,N_2729);
nand U3509 (N_3509,N_2143,N_151);
and U3510 (N_3510,N_627,N_165);
nor U3511 (N_3511,N_663,N_221);
or U3512 (N_3512,N_950,N_1649);
xor U3513 (N_3513,N_308,N_60);
xor U3514 (N_3514,N_239,N_248);
nand U3515 (N_3515,N_2233,N_1944);
nor U3516 (N_3516,N_945,N_2349);
and U3517 (N_3517,N_1359,N_755);
or U3518 (N_3518,N_474,N_2775);
xnor U3519 (N_3519,N_2025,N_2784);
and U3520 (N_3520,N_1446,N_1891);
nor U3521 (N_3521,N_1670,N_1299);
or U3522 (N_3522,N_1071,N_1890);
xor U3523 (N_3523,N_1194,N_504);
nor U3524 (N_3524,N_1270,N_695);
xnor U3525 (N_3525,N_399,N_863);
nor U3526 (N_3526,N_1005,N_2430);
nor U3527 (N_3527,N_258,N_1600);
and U3528 (N_3528,N_1355,N_24);
xor U3529 (N_3529,N_2008,N_1832);
and U3530 (N_3530,N_2489,N_1122);
or U3531 (N_3531,N_2998,N_2964);
and U3532 (N_3532,N_1599,N_2759);
nand U3533 (N_3533,N_1597,N_374);
nand U3534 (N_3534,N_2346,N_2843);
and U3535 (N_3535,N_43,N_436);
nand U3536 (N_3536,N_545,N_548);
nand U3537 (N_3537,N_610,N_310);
or U3538 (N_3538,N_532,N_1174);
or U3539 (N_3539,N_315,N_1344);
and U3540 (N_3540,N_1349,N_669);
nor U3541 (N_3541,N_226,N_2810);
and U3542 (N_3542,N_833,N_1500);
nand U3543 (N_3543,N_1162,N_707);
nand U3544 (N_3544,N_742,N_1687);
nor U3545 (N_3545,N_1875,N_149);
or U3546 (N_3546,N_1370,N_1037);
or U3547 (N_3547,N_2766,N_1842);
nor U3548 (N_3548,N_1345,N_899);
and U3549 (N_3549,N_1024,N_2204);
nor U3550 (N_3550,N_1982,N_262);
and U3551 (N_3551,N_591,N_2280);
nor U3552 (N_3552,N_1115,N_1280);
or U3553 (N_3553,N_612,N_2223);
xor U3554 (N_3554,N_2785,N_2463);
and U3555 (N_3555,N_1629,N_2026);
and U3556 (N_3556,N_408,N_1840);
or U3557 (N_3557,N_1120,N_1868);
and U3558 (N_3558,N_306,N_348);
nand U3559 (N_3559,N_2972,N_2440);
nand U3560 (N_3560,N_1062,N_55);
nand U3561 (N_3561,N_1454,N_2660);
nor U3562 (N_3562,N_434,N_2547);
xnor U3563 (N_3563,N_1730,N_1095);
or U3564 (N_3564,N_1016,N_2313);
nand U3565 (N_3565,N_2616,N_608);
and U3566 (N_3566,N_1955,N_1091);
or U3567 (N_3567,N_281,N_1325);
nor U3568 (N_3568,N_270,N_23);
nor U3569 (N_3569,N_392,N_1652);
or U3570 (N_3570,N_1155,N_815);
and U3571 (N_3571,N_2183,N_2508);
nor U3572 (N_3572,N_126,N_87);
nand U3573 (N_3573,N_1185,N_1610);
nand U3574 (N_3574,N_2281,N_2744);
or U3575 (N_3575,N_1217,N_252);
nor U3576 (N_3576,N_2410,N_1908);
nand U3577 (N_3577,N_605,N_2893);
or U3578 (N_3578,N_2949,N_1292);
nand U3579 (N_3579,N_224,N_2116);
or U3580 (N_3580,N_973,N_1881);
or U3581 (N_3581,N_622,N_666);
nand U3582 (N_3582,N_2421,N_1283);
xor U3583 (N_3583,N_1722,N_101);
xor U3584 (N_3584,N_2974,N_2036);
or U3585 (N_3585,N_1432,N_753);
nor U3586 (N_3586,N_988,N_1561);
nand U3587 (N_3587,N_2200,N_538);
xor U3588 (N_3588,N_834,N_843);
nand U3589 (N_3589,N_1098,N_2220);
xor U3590 (N_3590,N_813,N_2094);
and U3591 (N_3591,N_1588,N_2185);
nor U3592 (N_3592,N_2001,N_1905);
or U3593 (N_3593,N_1408,N_209);
and U3594 (N_3594,N_435,N_2612);
or U3595 (N_3595,N_2596,N_991);
nor U3596 (N_3596,N_2941,N_1684);
nand U3597 (N_3597,N_684,N_2444);
xnor U3598 (N_3598,N_1831,N_1808);
nand U3599 (N_3599,N_2007,N_184);
or U3600 (N_3600,N_2022,N_696);
nor U3601 (N_3601,N_1341,N_2511);
xnor U3602 (N_3602,N_2278,N_166);
and U3603 (N_3603,N_1945,N_366);
xnor U3604 (N_3604,N_1826,N_249);
nand U3605 (N_3605,N_1812,N_1685);
nand U3606 (N_3606,N_887,N_487);
nor U3607 (N_3607,N_2548,N_2033);
nor U3608 (N_3608,N_2598,N_1679);
nor U3609 (N_3609,N_473,N_2565);
nand U3610 (N_3610,N_1683,N_2462);
nor U3611 (N_3611,N_951,N_1762);
and U3612 (N_3612,N_2876,N_2706);
nor U3613 (N_3613,N_799,N_1701);
xor U3614 (N_3614,N_2831,N_956);
nand U3615 (N_3615,N_2357,N_691);
nor U3616 (N_3616,N_592,N_598);
and U3617 (N_3617,N_147,N_2958);
nand U3618 (N_3618,N_2340,N_1467);
nand U3619 (N_3619,N_1593,N_136);
and U3620 (N_3620,N_1508,N_901);
xor U3621 (N_3621,N_992,N_2051);
nand U3622 (N_3622,N_104,N_870);
and U3623 (N_3623,N_1375,N_482);
nand U3624 (N_3624,N_5,N_1559);
nor U3625 (N_3625,N_2887,N_456);
and U3626 (N_3626,N_285,N_749);
nor U3627 (N_3627,N_777,N_231);
and U3628 (N_3628,N_996,N_1145);
and U3629 (N_3629,N_119,N_494);
nand U3630 (N_3630,N_2725,N_1114);
xor U3631 (N_3631,N_2922,N_633);
or U3632 (N_3632,N_1392,N_2703);
or U3633 (N_3633,N_819,N_791);
nor U3634 (N_3634,N_2747,N_728);
and U3635 (N_3635,N_797,N_1);
nor U3636 (N_3636,N_572,N_1653);
nand U3637 (N_3637,N_2179,N_2059);
xnor U3638 (N_3638,N_1849,N_2331);
xnor U3639 (N_3639,N_851,N_1874);
nand U3640 (N_3640,N_2034,N_1766);
xnor U3641 (N_3641,N_1423,N_1234);
or U3642 (N_3642,N_601,N_1382);
nor U3643 (N_3643,N_2867,N_460);
and U3644 (N_3644,N_1358,N_2261);
nand U3645 (N_3645,N_342,N_2145);
and U3646 (N_3646,N_1166,N_1137);
or U3647 (N_3647,N_2394,N_1860);
or U3648 (N_3648,N_2014,N_2479);
nor U3649 (N_3649,N_982,N_741);
and U3650 (N_3650,N_2467,N_34);
and U3651 (N_3651,N_2124,N_866);
xnor U3652 (N_3652,N_49,N_2865);
or U3653 (N_3653,N_2362,N_1023);
xor U3654 (N_3654,N_410,N_1011);
xor U3655 (N_3655,N_2353,N_651);
or U3656 (N_3656,N_227,N_2674);
xor U3657 (N_3657,N_1695,N_596);
or U3658 (N_3658,N_824,N_1157);
nor U3659 (N_3659,N_2398,N_1937);
nor U3660 (N_3660,N_1604,N_2845);
nor U3661 (N_3661,N_1390,N_1479);
nor U3662 (N_3662,N_52,N_1017);
and U3663 (N_3663,N_1549,N_2662);
or U3664 (N_3664,N_1789,N_2624);
nand U3665 (N_3665,N_1063,N_518);
xor U3666 (N_3666,N_1067,N_2792);
or U3667 (N_3667,N_2273,N_2587);
nand U3668 (N_3668,N_1272,N_621);
and U3669 (N_3669,N_1225,N_3);
or U3670 (N_3670,N_1387,N_2342);
or U3671 (N_3671,N_1773,N_882);
xnor U3672 (N_3672,N_1030,N_2242);
nor U3673 (N_3673,N_2726,N_683);
or U3674 (N_3674,N_2602,N_1778);
or U3675 (N_3675,N_2309,N_2606);
xor U3676 (N_3676,N_2728,N_2923);
or U3677 (N_3677,N_2809,N_415);
nor U3678 (N_3678,N_1850,N_1705);
nor U3679 (N_3679,N_1658,N_1118);
xnor U3680 (N_3680,N_860,N_1584);
and U3681 (N_3681,N_952,N_1350);
or U3682 (N_3682,N_2214,N_2137);
nor U3683 (N_3683,N_203,N_853);
nor U3684 (N_3684,N_1433,N_2742);
and U3685 (N_3685,N_626,N_1326);
and U3686 (N_3686,N_2090,N_477);
nor U3687 (N_3687,N_1972,N_1076);
nor U3688 (N_3688,N_1332,N_2895);
or U3689 (N_3689,N_1650,N_1839);
nor U3690 (N_3690,N_842,N_1178);
xnor U3691 (N_3691,N_2504,N_936);
xor U3692 (N_3692,N_565,N_2068);
or U3693 (N_3693,N_1759,N_1858);
or U3694 (N_3694,N_318,N_1231);
nand U3695 (N_3695,N_1187,N_737);
or U3696 (N_3696,N_2990,N_2482);
nand U3697 (N_3697,N_2314,N_977);
nand U3698 (N_3698,N_2041,N_2086);
nor U3699 (N_3699,N_1010,N_2379);
or U3700 (N_3700,N_116,N_1737);
or U3701 (N_3701,N_1618,N_1035);
xor U3702 (N_3702,N_232,N_1450);
and U3703 (N_3703,N_983,N_628);
nand U3704 (N_3704,N_76,N_898);
nand U3705 (N_3705,N_1845,N_312);
or U3706 (N_3706,N_2690,N_1025);
and U3707 (N_3707,N_2438,N_1551);
nand U3708 (N_3708,N_2146,N_51);
or U3709 (N_3709,N_1213,N_2106);
nor U3710 (N_3710,N_2114,N_351);
xnor U3711 (N_3711,N_2748,N_2653);
nor U3712 (N_3712,N_890,N_1726);
nand U3713 (N_3713,N_2095,N_2715);
and U3714 (N_3714,N_2835,N_1798);
xnor U3715 (N_3715,N_1130,N_1542);
or U3716 (N_3716,N_925,N_1288);
xor U3717 (N_3717,N_1674,N_2400);
and U3718 (N_3718,N_327,N_1993);
nand U3719 (N_3719,N_876,N_425);
nor U3720 (N_3720,N_2833,N_387);
nand U3721 (N_3721,N_693,N_2275);
nand U3722 (N_3722,N_1371,N_1743);
and U3723 (N_3723,N_2165,N_2607);
nor U3724 (N_3724,N_2402,N_1487);
and U3725 (N_3725,N_1196,N_1884);
or U3726 (N_3726,N_1259,N_873);
nor U3727 (N_3727,N_134,N_1301);
and U3728 (N_3728,N_1660,N_644);
and U3729 (N_3729,N_2678,N_1509);
nand U3730 (N_3730,N_337,N_437);
and U3731 (N_3731,N_1616,N_1048);
and U3732 (N_3732,N_183,N_2580);
xnor U3733 (N_3733,N_1140,N_754);
nand U3734 (N_3734,N_1156,N_199);
nor U3735 (N_3735,N_1061,N_4);
nand U3736 (N_3736,N_1910,N_1611);
or U3737 (N_3737,N_1519,N_1671);
nand U3738 (N_3738,N_2399,N_2140);
and U3739 (N_3739,N_932,N_2171);
or U3740 (N_3740,N_2293,N_2174);
and U3741 (N_3741,N_302,N_223);
nor U3742 (N_3742,N_828,N_124);
nor U3743 (N_3743,N_1971,N_2286);
or U3744 (N_3744,N_2804,N_1659);
xnor U3745 (N_3745,N_2136,N_588);
nand U3746 (N_3746,N_1368,N_1656);
nor U3747 (N_3747,N_1143,N_2099);
or U3748 (N_3748,N_1245,N_2683);
and U3749 (N_3749,N_299,N_2582);
nand U3750 (N_3750,N_869,N_2019);
or U3751 (N_3751,N_422,N_1306);
and U3752 (N_3752,N_2667,N_1376);
and U3753 (N_3753,N_91,N_676);
nand U3754 (N_3754,N_1009,N_2782);
xnor U3755 (N_3755,N_1750,N_1015);
or U3756 (N_3756,N_2239,N_2407);
or U3757 (N_3757,N_328,N_1256);
nand U3758 (N_3758,N_1285,N_1293);
or U3759 (N_3759,N_1442,N_1363);
or U3760 (N_3760,N_2164,N_1885);
or U3761 (N_3761,N_1817,N_1045);
or U3762 (N_3762,N_2270,N_1021);
nor U3763 (N_3763,N_2948,N_927);
or U3764 (N_3764,N_1197,N_1262);
and U3765 (N_3765,N_272,N_1428);
or U3766 (N_3766,N_1516,N_2632);
xor U3767 (N_3767,N_2884,N_2433);
and U3768 (N_3768,N_733,N_835);
xor U3769 (N_3769,N_140,N_1777);
or U3770 (N_3770,N_139,N_164);
or U3771 (N_3771,N_1257,N_1829);
xnor U3772 (N_3772,N_2695,N_1388);
nand U3773 (N_3773,N_2685,N_879);
or U3774 (N_3774,N_1765,N_1263);
nor U3775 (N_3775,N_1804,N_1253);
nor U3776 (N_3776,N_15,N_2323);
or U3777 (N_3777,N_2089,N_2013);
and U3778 (N_3778,N_2330,N_2491);
nor U3779 (N_3779,N_2363,N_1128);
and U3780 (N_3780,N_725,N_512);
or U3781 (N_3781,N_2193,N_2531);
or U3782 (N_3782,N_20,N_2749);
or U3783 (N_3783,N_1702,N_99);
or U3784 (N_3784,N_1814,N_994);
nand U3785 (N_3785,N_1135,N_1698);
xor U3786 (N_3786,N_316,N_395);
xnor U3787 (N_3787,N_163,N_580);
nor U3788 (N_3788,N_2608,N_530);
xnor U3789 (N_3789,N_1546,N_2707);
and U3790 (N_3790,N_1337,N_1258);
nand U3791 (N_3791,N_428,N_471);
nand U3792 (N_3792,N_11,N_756);
and U3793 (N_3793,N_416,N_829);
and U3794 (N_3794,N_389,N_1837);
xnor U3795 (N_3795,N_2852,N_2939);
xnor U3796 (N_3796,N_1835,N_966);
or U3797 (N_3797,N_632,N_381);
or U3798 (N_3798,N_2839,N_1028);
or U3799 (N_3799,N_918,N_933);
and U3800 (N_3800,N_2360,N_297);
nand U3801 (N_3801,N_2620,N_1746);
and U3802 (N_3802,N_2959,N_1296);
nand U3803 (N_3803,N_2389,N_1499);
and U3804 (N_3804,N_2737,N_1160);
nand U3805 (N_3805,N_2260,N_2391);
and U3806 (N_3806,N_2588,N_1936);
and U3807 (N_3807,N_796,N_346);
or U3808 (N_3808,N_2882,N_1006);
or U3809 (N_3809,N_236,N_1032);
or U3810 (N_3810,N_1437,N_675);
nand U3811 (N_3811,N_2599,N_1548);
nor U3812 (N_3812,N_2426,N_647);
nor U3813 (N_3813,N_2823,N_393);
xor U3814 (N_3814,N_1787,N_1557);
or U3815 (N_3815,N_2938,N_2092);
and U3816 (N_3816,N_2332,N_78);
nor U3817 (N_3817,N_1290,N_1324);
xnor U3818 (N_3818,N_1563,N_2795);
or U3819 (N_3819,N_1482,N_2860);
nor U3820 (N_3820,N_1664,N_2395);
and U3821 (N_3821,N_2899,N_118);
nand U3822 (N_3822,N_1096,N_1540);
xor U3823 (N_3823,N_1585,N_1190);
or U3824 (N_3824,N_2539,N_2840);
nand U3825 (N_3825,N_2180,N_2641);
or U3826 (N_3826,N_2781,N_1351);
or U3827 (N_3827,N_2047,N_290);
xnor U3828 (N_3828,N_990,N_2738);
and U3829 (N_3829,N_1996,N_2049);
or U3830 (N_3830,N_2866,N_421);
and U3831 (N_3831,N_125,N_2758);
nand U3832 (N_3832,N_1142,N_1520);
nand U3833 (N_3833,N_1888,N_2740);
or U3834 (N_3834,N_2864,N_1537);
nand U3835 (N_3835,N_2117,N_336);
xor U3836 (N_3836,N_2448,N_1497);
nor U3837 (N_3837,N_1223,N_841);
or U3838 (N_3838,N_2425,N_27);
nor U3839 (N_3839,N_2832,N_836);
and U3840 (N_3840,N_1979,N_2567);
or U3841 (N_3841,N_1825,N_1643);
nand U3842 (N_3842,N_466,N_1079);
and U3843 (N_3843,N_273,N_2186);
xor U3844 (N_3844,N_150,N_782);
nor U3845 (N_3845,N_1725,N_757);
nor U3846 (N_3846,N_1486,N_1149);
nand U3847 (N_3847,N_781,N_1090);
nor U3848 (N_3848,N_858,N_916);
xnor U3849 (N_3849,N_2688,N_1622);
and U3850 (N_3850,N_2704,N_41);
nor U3851 (N_3851,N_845,N_902);
and U3852 (N_3852,N_912,N_1031);
nand U3853 (N_3853,N_1531,N_1070);
nor U3854 (N_3854,N_2768,N_334);
nor U3855 (N_3855,N_1620,N_1739);
xnor U3856 (N_3856,N_2960,N_529);
xor U3857 (N_3857,N_407,N_1661);
nor U3858 (N_3858,N_1007,N_1141);
and U3859 (N_3859,N_2048,N_2190);
xor U3860 (N_3860,N_2537,N_1530);
nand U3861 (N_3861,N_969,N_692);
and U3862 (N_3862,N_1939,N_486);
nand U3863 (N_3863,N_2705,N_1241);
and U3864 (N_3864,N_1308,N_2510);
nor U3865 (N_3865,N_1637,N_2341);
or U3866 (N_3866,N_2248,N_1214);
nand U3867 (N_3867,N_22,N_2559);
or U3868 (N_3868,N_2385,N_1421);
nor U3869 (N_3869,N_205,N_724);
nor U3870 (N_3870,N_2844,N_177);
nor U3871 (N_3871,N_2476,N_514);
xnor U3872 (N_3872,N_803,N_2413);
xnor U3873 (N_3873,N_2287,N_430);
and U3874 (N_3874,N_242,N_1181);
nand U3875 (N_3875,N_2770,N_943);
nand U3876 (N_3876,N_1498,N_225);
xnor U3877 (N_3877,N_775,N_40);
and U3878 (N_3878,N_1416,N_2856);
nand U3879 (N_3879,N_442,N_1038);
nor U3880 (N_3880,N_490,N_1960);
nand U3881 (N_3881,N_1039,N_190);
nor U3882 (N_3882,N_1277,N_1033);
nand U3883 (N_3883,N_1946,N_1167);
nand U3884 (N_3884,N_2700,N_525);
or U3885 (N_3885,N_1163,N_2121);
or U3886 (N_3886,N_2883,N_1923);
nor U3887 (N_3887,N_1334,N_2432);
and U3888 (N_3888,N_1954,N_1715);
nor U3889 (N_3889,N_2184,N_2307);
or U3890 (N_3890,N_1841,N_276);
and U3891 (N_3891,N_394,N_2322);
nand U3892 (N_3892,N_1980,N_1381);
nor U3893 (N_3893,N_2570,N_734);
or U3894 (N_3894,N_121,N_1418);
and U3895 (N_3895,N_2500,N_2584);
xnor U3896 (N_3896,N_1152,N_637);
nor U3897 (N_3897,N_2401,N_238);
and U3898 (N_3898,N_1638,N_1168);
nand U3899 (N_3899,N_175,N_189);
nor U3900 (N_3900,N_2574,N_2819);
nand U3901 (N_3901,N_2492,N_635);
nand U3902 (N_3902,N_1348,N_2151);
and U3903 (N_3903,N_908,N_1770);
xor U3904 (N_3904,N_2447,N_1171);
nor U3905 (N_3905,N_2091,N_2241);
nand U3906 (N_3906,N_1330,N_689);
or U3907 (N_3907,N_2983,N_1064);
nand U3908 (N_3908,N_2358,N_937);
and U3909 (N_3909,N_1984,N_1942);
or U3910 (N_3910,N_2267,N_2027);
and U3911 (N_3911,N_2979,N_1236);
nor U3912 (N_3912,N_2110,N_1819);
nand U3913 (N_3913,N_1235,N_2409);
nor U3914 (N_3914,N_2736,N_1123);
nor U3915 (N_3915,N_1894,N_1889);
or U3916 (N_3916,N_2645,N_83);
xor U3917 (N_3917,N_2150,N_173);
and U3918 (N_3918,N_1657,N_924);
or U3919 (N_3919,N_1782,N_2569);
xnor U3920 (N_3920,N_2727,N_566);
and U3921 (N_3921,N_2123,N_2997);
nor U3922 (N_3922,N_347,N_359);
xnor U3923 (N_3923,N_419,N_2967);
xnor U3924 (N_3924,N_2720,N_1314);
or U3925 (N_3925,N_255,N_1119);
nor U3926 (N_3926,N_369,N_1125);
and U3927 (N_3927,N_322,N_2821);
xnor U3928 (N_3928,N_877,N_2779);
nand U3929 (N_3929,N_98,N_1873);
and U3930 (N_3930,N_2249,N_1001);
nor U3931 (N_3931,N_1677,N_2518);
or U3932 (N_3932,N_289,N_1496);
or U3933 (N_3933,N_2262,N_1309);
and U3934 (N_3934,N_602,N_900);
nor U3935 (N_3935,N_2900,N_2820);
nand U3936 (N_3936,N_296,N_2892);
nand U3937 (N_3937,N_499,N_2677);
and U3938 (N_3938,N_2291,N_2080);
nor U3939 (N_3939,N_515,N_2468);
xor U3940 (N_3940,N_26,N_2581);
nor U3941 (N_3941,N_561,N_2862);
nor U3942 (N_3942,N_1477,N_1365);
xnor U3943 (N_3943,N_122,N_2067);
nor U3944 (N_3944,N_2714,N_1338);
nand U3945 (N_3945,N_1080,N_1769);
nor U3946 (N_3946,N_88,N_2786);
or U3947 (N_3947,N_307,N_2355);
and U3948 (N_3948,N_2836,N_1768);
nand U3949 (N_3949,N_1792,N_1636);
or U3950 (N_3950,N_1880,N_2914);
nand U3951 (N_3951,N_1818,N_2228);
xnor U3952 (N_3952,N_2096,N_979);
nand U3953 (N_3953,N_584,N_2793);
xnor U3954 (N_3954,N_752,N_2192);
or U3955 (N_3955,N_1869,N_198);
nand U3956 (N_3956,N_402,N_1879);
nor U3957 (N_3957,N_1367,N_2437);
nor U3958 (N_3958,N_949,N_2002);
and U3959 (N_3959,N_2996,N_1165);
nand U3960 (N_3960,N_54,N_1014);
and U3961 (N_3961,N_1282,N_411);
and U3962 (N_3962,N_145,N_1925);
nor U3963 (N_3963,N_2073,N_2339);
nand U3964 (N_3964,N_32,N_2732);
xnor U3965 (N_3965,N_480,N_2783);
nor U3966 (N_3966,N_1975,N_2206);
nand U3967 (N_3967,N_1465,N_352);
nand U3968 (N_3968,N_21,N_2069);
xor U3969 (N_3969,N_2271,N_2100);
nor U3970 (N_3970,N_1964,N_485);
xor U3971 (N_3971,N_2218,N_1361);
and U3972 (N_3972,N_723,N_848);
or U3973 (N_3973,N_986,N_643);
nand U3974 (N_3974,N_2988,N_1057);
nor U3975 (N_3975,N_1471,N_1242);
xor U3976 (N_3976,N_2405,N_1366);
xnor U3977 (N_3977,N_1474,N_2871);
nor U3978 (N_3978,N_2571,N_1791);
and U3979 (N_3979,N_1346,N_1900);
and U3980 (N_3980,N_2879,N_1699);
nor U3981 (N_3981,N_1226,N_2880);
nand U3982 (N_3982,N_220,N_2493);
xnor U3983 (N_3983,N_2288,N_981);
and U3984 (N_3984,N_2263,N_253);
and U3985 (N_3985,N_1239,N_2039);
nand U3986 (N_3986,N_2231,N_670);
nor U3987 (N_3987,N_2387,N_219);
and U3988 (N_3988,N_2886,N_431);
or U3989 (N_3989,N_382,N_1438);
nand U3990 (N_3990,N_1755,N_708);
or U3991 (N_3991,N_71,N_2000);
or U3992 (N_3992,N_1928,N_2102);
xor U3993 (N_3993,N_1965,N_520);
nand U3994 (N_3994,N_1184,N_2743);
or U3995 (N_3995,N_1805,N_2219);
or U3996 (N_3996,N_1741,N_1673);
nor U3997 (N_3997,N_2112,N_1075);
and U3998 (N_3998,N_1221,N_218);
and U3999 (N_3999,N_152,N_1238);
xor U4000 (N_4000,N_16,N_1472);
nand U4001 (N_4001,N_568,N_167);
or U4002 (N_4002,N_143,N_2530);
xor U4003 (N_4003,N_2898,N_2817);
nor U4004 (N_4004,N_913,N_2724);
xor U4005 (N_4005,N_1439,N_30);
and U4006 (N_4006,N_2577,N_2541);
and U4007 (N_4007,N_2848,N_2238);
nor U4008 (N_4008,N_56,N_2968);
and U4009 (N_4009,N_1809,N_589);
xor U4010 (N_4010,N_713,N_362);
xor U4011 (N_4011,N_1550,N_2603);
nor U4012 (N_4012,N_892,N_70);
or U4013 (N_4013,N_859,N_604);
nor U4014 (N_4014,N_506,N_1159);
xnor U4015 (N_4015,N_2277,N_2367);
nand U4016 (N_4016,N_528,N_555);
nand U4017 (N_4017,N_747,N_2903);
nand U4018 (N_4018,N_1973,N_805);
nand U4019 (N_4019,N_1211,N_2994);
or U4020 (N_4020,N_476,N_459);
and U4021 (N_4021,N_138,N_1227);
and U4022 (N_4022,N_97,N_1295);
nand U4023 (N_4023,N_293,N_1651);
nor U4024 (N_4024,N_2680,N_1362);
nand U4025 (N_4025,N_2675,N_420);
nand U4026 (N_4026,N_1243,N_172);
xor U4027 (N_4027,N_940,N_1956);
and U4028 (N_4028,N_2182,N_2416);
nand U4029 (N_4029,N_1040,N_867);
nor U4030 (N_4030,N_1539,N_2849);
xor U4031 (N_4031,N_321,N_1494);
and U4032 (N_4032,N_1863,N_2803);
nand U4033 (N_4033,N_557,N_740);
or U4034 (N_4034,N_2456,N_2697);
and U4035 (N_4035,N_2965,N_1630);
nor U4036 (N_4036,N_2629,N_1427);
or U4037 (N_4037,N_2483,N_1854);
nand U4038 (N_4038,N_509,N_521);
or U4039 (N_4039,N_191,N_50);
and U4040 (N_4040,N_2319,N_1321);
nand U4041 (N_4041,N_2024,N_1581);
nor U4042 (N_4042,N_1926,N_319);
xnor U4043 (N_4043,N_1747,N_1396);
and U4044 (N_4044,N_2648,N_543);
xnor U4045 (N_4045,N_66,N_2191);
nand U4046 (N_4046,N_1728,N_586);
or U4047 (N_4047,N_237,N_874);
xnor U4048 (N_4048,N_2550,N_2935);
xor U4049 (N_4049,N_2702,N_228);
or U4050 (N_4050,N_2816,N_1999);
xor U4051 (N_4051,N_2244,N_2169);
nor U4052 (N_4052,N_368,N_1532);
or U4053 (N_4053,N_1460,N_502);
xor U4054 (N_4054,N_1803,N_1291);
nand U4055 (N_4055,N_2942,N_1491);
xor U4056 (N_4056,N_1717,N_2927);
or U4057 (N_4057,N_117,N_1953);
or U4058 (N_4058,N_1978,N_210);
nor U4059 (N_4059,N_2446,N_2364);
nor U4060 (N_4060,N_108,N_2197);
and U4061 (N_4061,N_2528,N_325);
nand U4062 (N_4062,N_2551,N_69);
nand U4063 (N_4063,N_1456,N_89);
xnor U4064 (N_4064,N_379,N_2087);
nor U4065 (N_4065,N_1621,N_2791);
xor U4066 (N_4066,N_1639,N_206);
nor U4067 (N_4067,N_2221,N_2872);
xnor U4068 (N_4068,N_1049,N_1082);
nand U4069 (N_4069,N_857,N_1072);
xnor U4070 (N_4070,N_2154,N_1255);
or U4071 (N_4071,N_1391,N_2420);
xnor U4072 (N_4072,N_1339,N_2868);
or U4073 (N_4073,N_2928,N_517);
or U4074 (N_4074,N_759,N_1784);
nand U4075 (N_4075,N_263,N_2555);
nand U4076 (N_4076,N_743,N_1384);
nor U4077 (N_4077,N_1276,N_697);
or U4078 (N_4078,N_1865,N_2857);
nor U4079 (N_4079,N_2028,N_715);
or U4080 (N_4080,N_42,N_539);
nor U4081 (N_4081,N_229,N_345);
xor U4082 (N_4082,N_2168,N_2336);
xnor U4083 (N_4083,N_769,N_2933);
xnor U4084 (N_4084,N_176,N_1515);
or U4085 (N_4085,N_1655,N_2017);
xor U4086 (N_4086,N_2070,N_2639);
or U4087 (N_4087,N_413,N_2875);
or U4088 (N_4088,N_1113,N_386);
and U4089 (N_4089,N_533,N_1320);
and U4090 (N_4090,N_1560,N_2298);
and U4091 (N_4091,N_86,N_2919);
nand U4092 (N_4092,N_1810,N_412);
nand U4093 (N_4093,N_1271,N_1776);
xnor U4094 (N_4094,N_120,N_274);
nor U4095 (N_4095,N_804,N_75);
nand U4096 (N_4096,N_540,N_1008);
nand U4097 (N_4097,N_1663,N_861);
xnor U4098 (N_4098,N_638,N_1666);
or U4099 (N_4099,N_593,N_496);
nor U4100 (N_4100,N_1681,N_1545);
nand U4101 (N_4101,N_2374,N_1645);
and U4102 (N_4102,N_2337,N_2411);
and U4103 (N_4103,N_2305,N_712);
xnor U4104 (N_4104,N_371,N_244);
xor U4105 (N_4105,N_156,N_1429);
or U4106 (N_4106,N_1632,N_811);
or U4107 (N_4107,N_2962,N_2711);
xnor U4108 (N_4108,N_2461,N_470);
xor U4109 (N_4109,N_193,N_1736);
xnor U4110 (N_4110,N_1733,N_2621);
xnor U4111 (N_4111,N_771,N_1127);
and U4112 (N_4112,N_2224,N_1686);
or U4113 (N_4113,N_2647,N_2525);
and U4114 (N_4114,N_1619,N_2149);
nor U4115 (N_4115,N_1598,N_1328);
xor U4116 (N_4116,N_1594,N_438);
xnor U4117 (N_4117,N_871,N_72);
nor U4118 (N_4118,N_2613,N_90);
or U4119 (N_4119,N_798,N_1101);
nor U4120 (N_4120,N_2419,N_2497);
and U4121 (N_4121,N_844,N_1700);
or U4122 (N_4122,N_196,N_614);
or U4123 (N_4123,N_1834,N_2954);
nor U4124 (N_4124,N_2505,N_1595);
nor U4125 (N_4125,N_686,N_2838);
xor U4126 (N_4126,N_2388,N_779);
nand U4127 (N_4127,N_295,N_2769);
and U4128 (N_4128,N_2256,N_1930);
xor U4129 (N_4129,N_817,N_1436);
and U4130 (N_4130,N_2657,N_888);
nor U4131 (N_4131,N_1189,N_1708);
xnor U4132 (N_4132,N_1081,N_2739);
nand U4133 (N_4133,N_1099,N_2172);
xor U4134 (N_4134,N_1286,N_2453);
or U4135 (N_4135,N_1553,N_1319);
nand U4136 (N_4136,N_553,N_2735);
or U4137 (N_4137,N_1053,N_484);
or U4138 (N_4138,N_2252,N_2266);
or U4139 (N_4139,N_2253,N_830);
or U4140 (N_4140,N_367,N_77);
xor U4141 (N_4141,N_344,N_856);
and U4142 (N_4142,N_309,N_2320);
xor U4143 (N_4143,N_746,N_1654);
nor U4144 (N_4144,N_2733,N_235);
and U4145 (N_4145,N_1431,N_2600);
or U4146 (N_4146,N_314,N_2368);
or U4147 (N_4147,N_959,N_304);
or U4148 (N_4148,N_2681,N_404);
nor U4149 (N_4149,N_1457,N_623);
and U4150 (N_4150,N_1763,N_1374);
xnor U4151 (N_4151,N_1222,N_2636);
xor U4152 (N_4152,N_1966,N_158);
xnor U4153 (N_4153,N_1988,N_2109);
and U4154 (N_4154,N_1372,N_169);
xnor U4155 (N_4155,N_1201,N_732);
nor U4156 (N_4156,N_1473,N_2656);
nor U4157 (N_4157,N_452,N_1644);
nor U4158 (N_4158,N_1133,N_1933);
or U4159 (N_4159,N_377,N_1251);
or U4160 (N_4160,N_1435,N_786);
nand U4161 (N_4161,N_2628,N_2128);
nor U4162 (N_4162,N_1278,N_2822);
and U4163 (N_4163,N_953,N_132);
nand U4164 (N_4164,N_240,N_1806);
and U4165 (N_4165,N_1647,N_1274);
and U4166 (N_4166,N_417,N_2397);
nand U4167 (N_4167,N_1112,N_361);
or U4168 (N_4168,N_910,N_1055);
or U4169 (N_4169,N_2382,N_1824);
and U4170 (N_4170,N_383,N_2615);
or U4171 (N_4171,N_862,N_613);
nor U4172 (N_4172,N_1760,N_1899);
nand U4173 (N_4173,N_1294,N_1173);
and U4174 (N_4174,N_717,N_2175);
xnor U4175 (N_4175,N_384,N_2590);
nand U4176 (N_4176,N_1424,N_1209);
nand U4177 (N_4177,N_764,N_2227);
nor U4178 (N_4178,N_2111,N_2772);
nand U4179 (N_4179,N_213,N_1451);
or U4180 (N_4180,N_1574,N_2098);
nand U4181 (N_4181,N_2891,N_1627);
or U4182 (N_4182,N_1997,N_1311);
nand U4183 (N_4183,N_269,N_330);
or U4184 (N_4184,N_1237,N_1707);
nand U4185 (N_4185,N_2103,N_418);
and U4186 (N_4186,N_2125,N_1693);
and U4187 (N_4187,N_2610,N_1788);
nor U4188 (N_4188,N_1571,N_160);
or U4189 (N_4189,N_1524,N_513);
and U4190 (N_4190,N_2926,N_763);
and U4191 (N_4191,N_2986,N_838);
and U4192 (N_4192,N_970,N_552);
or U4193 (N_4193,N_1232,N_681);
nand U4194 (N_4194,N_1453,N_1480);
nand U4195 (N_4195,N_1305,N_1855);
xnor U4196 (N_4196,N_2315,N_2496);
or U4197 (N_4197,N_690,N_2317);
or U4198 (N_4198,N_672,N_80);
and U4199 (N_4199,N_1935,N_2853);
xor U4200 (N_4200,N_958,N_2869);
xor U4201 (N_4201,N_1689,N_1289);
nor U4202 (N_4202,N_1641,N_558);
nor U4203 (N_4203,N_1761,N_1994);
nand U4204 (N_4204,N_2257,N_1110);
and U4205 (N_4205,N_1744,N_2423);
or U4206 (N_4206,N_483,N_1191);
nand U4207 (N_4207,N_2561,N_606);
nand U4208 (N_4208,N_0,N_1503);
nor U4209 (N_4209,N_2195,N_214);
or U4210 (N_4210,N_730,N_2501);
nor U4211 (N_4211,N_45,N_2194);
and U4212 (N_4212,N_2436,N_2878);
nand U4213 (N_4213,N_2135,N_2617);
nand U4214 (N_4214,N_2199,N_2888);
or U4215 (N_4215,N_905,N_264);
nand U4216 (N_4216,N_100,N_1948);
xor U4217 (N_4217,N_216,N_2348);
xnor U4218 (N_4218,N_2516,N_2350);
nand U4219 (N_4219,N_9,N_503);
nand U4220 (N_4220,N_850,N_7);
xor U4221 (N_4221,N_1443,N_2037);
xor U4222 (N_4222,N_820,N_2443);
and U4223 (N_4223,N_1534,N_1086);
nor U4224 (N_4224,N_2851,N_335);
and U4225 (N_4225,N_2563,N_1383);
and U4226 (N_4226,N_2422,N_2694);
nand U4227 (N_4227,N_2471,N_1394);
and U4228 (N_4228,N_534,N_2889);
and U4229 (N_4229,N_79,N_148);
xnor U4230 (N_4230,N_1385,N_954);
xnor U4231 (N_4231,N_397,N_141);
and U4232 (N_4232,N_2328,N_1298);
or U4233 (N_4233,N_2093,N_1799);
xnor U4234 (N_4234,N_2651,N_2594);
nor U4235 (N_4235,N_1907,N_1917);
or U4236 (N_4236,N_2576,N_375);
and U4237 (N_4237,N_61,N_603);
or U4238 (N_4238,N_2157,N_373);
or U4239 (N_4239,N_1526,N_1871);
xnor U4240 (N_4240,N_2178,N_2552);
nor U4241 (N_4241,N_432,N_2474);
xnor U4242 (N_4242,N_2502,N_449);
nand U4243 (N_4243,N_1772,N_1089);
nor U4244 (N_4244,N_569,N_1901);
xor U4245 (N_4245,N_254,N_508);
nor U4246 (N_4246,N_323,N_2931);
and U4247 (N_4247,N_447,N_1169);
and U4248 (N_4248,N_631,N_207);
or U4249 (N_4249,N_2254,N_1983);
nor U4250 (N_4250,N_2731,N_2545);
nand U4251 (N_4251,N_2207,N_551);
or U4252 (N_4252,N_578,N_2304);
nand U4253 (N_4253,N_2088,N_2912);
or U4254 (N_4254,N_700,N_2921);
and U4255 (N_4255,N_2654,N_563);
xor U4256 (N_4256,N_1104,N_259);
and U4257 (N_4257,N_2316,N_1448);
nor U4258 (N_4258,N_1331,N_1452);
xor U4259 (N_4259,N_29,N_1469);
nor U4260 (N_4260,N_885,N_1963);
nand U4261 (N_4261,N_808,N_2589);
nor U4262 (N_4262,N_2755,N_1313);
and U4263 (N_4263,N_1018,N_792);
and U4264 (N_4264,N_453,N_1511);
and U4265 (N_4265,N_39,N_179);
or U4266 (N_4266,N_886,N_1583);
nor U4267 (N_4267,N_1322,N_2030);
nor U4268 (N_4268,N_1821,N_448);
nor U4269 (N_4269,N_1395,N_1399);
or U4270 (N_4270,N_234,N_738);
and U4271 (N_4271,N_1919,N_2344);
xnor U4272 (N_4272,N_338,N_1043);
nor U4273 (N_4273,N_1625,N_1403);
or U4274 (N_4274,N_1041,N_1706);
and U4275 (N_4275,N_2269,N_774);
nand U4276 (N_4276,N_1210,N_2692);
xnor U4277 (N_4277,N_2969,N_1934);
xnor U4278 (N_4278,N_1843,N_1275);
and U4279 (N_4279,N_2841,N_2661);
nand U4280 (N_4280,N_2756,N_1614);
xor U4281 (N_4281,N_930,N_2767);
or U4282 (N_4282,N_665,N_1352);
or U4283 (N_4283,N_998,N_2562);
or U4284 (N_4284,N_816,N_522);
nand U4285 (N_4285,N_1297,N_1615);
and U4286 (N_4286,N_2635,N_1507);
nor U4287 (N_4287,N_968,N_2203);
nand U4288 (N_4288,N_2708,N_2129);
nand U4289 (N_4289,N_1148,N_2881);
nand U4290 (N_4290,N_457,N_1059);
or U4291 (N_4291,N_2712,N_2764);
xor U4292 (N_4292,N_2805,N_2347);
xnor U4293 (N_4293,N_903,N_1106);
nand U4294 (N_4294,N_1505,N_1183);
or U4295 (N_4295,N_2427,N_2042);
and U4296 (N_4296,N_450,N_576);
nand U4297 (N_4297,N_2722,N_535);
or U4298 (N_4298,N_180,N_1800);
xnor U4299 (N_4299,N_2012,N_2300);
nand U4300 (N_4300,N_748,N_2062);
and U4301 (N_4301,N_1488,N_2666);
or U4302 (N_4302,N_1667,N_18);
and U4303 (N_4303,N_1527,N_685);
and U4304 (N_4304,N_2043,N_1927);
nand U4305 (N_4305,N_1393,N_1273);
xnor U4306 (N_4306,N_2351,N_356);
nor U4307 (N_4307,N_357,N_768);
nand U4308 (N_4308,N_2807,N_1269);
nand U4309 (N_4309,N_1742,N_2950);
or U4310 (N_4310,N_1703,N_2885);
nand U4311 (N_4311,N_1266,N_1300);
and U4312 (N_4312,N_1732,N_1969);
nand U4313 (N_4313,N_2264,N_2827);
nor U4314 (N_4314,N_594,N_112);
and U4315 (N_4315,N_1405,N_2055);
nand U4316 (N_4316,N_2751,N_2225);
nand U4317 (N_4317,N_1912,N_2937);
nor U4318 (N_4318,N_1380,N_195);
and U4319 (N_4319,N_822,N_1517);
and U4320 (N_4320,N_1932,N_1573);
nor U4321 (N_4321,N_2018,N_2646);
nor U4322 (N_4322,N_640,N_2311);
and U4323 (N_4323,N_2120,N_630);
nor U4324 (N_4324,N_2074,N_2046);
xnor U4325 (N_4325,N_661,N_2294);
and U4326 (N_4326,N_360,N_2406);
and U4327 (N_4327,N_355,N_2970);
nor U4328 (N_4328,N_305,N_2664);
and U4329 (N_4329,N_2325,N_2485);
nor U4330 (N_4330,N_1129,N_2591);
nand U4331 (N_4331,N_911,N_2506);
and U4332 (N_4332,N_1461,N_1147);
and U4333 (N_4333,N_128,N_2846);
nand U4334 (N_4334,N_2980,N_2324);
xnor U4335 (N_4335,N_461,N_2480);
or U4336 (N_4336,N_1068,N_1215);
or U4337 (N_4337,N_581,N_2684);
and U4338 (N_4338,N_1047,N_2773);
nor U4339 (N_4339,N_2572,N_1536);
nand U4340 (N_4340,N_174,N_358);
xor U4341 (N_4341,N_2995,N_2952);
xor U4342 (N_4342,N_1353,N_380);
nand U4343 (N_4343,N_292,N_2127);
nor U4344 (N_4344,N_241,N_400);
or U4345 (N_4345,N_1065,N_1307);
xor U4346 (N_4346,N_2710,N_1444);
nand U4347 (N_4347,N_1564,N_110);
nor U4348 (N_4348,N_1852,N_1202);
nor U4349 (N_4349,N_500,N_2289);
xor U4350 (N_4350,N_2284,N_915);
or U4351 (N_4351,N_616,N_1069);
xnor U4352 (N_4352,N_1134,N_1828);
nand U4353 (N_4353,N_1712,N_495);
xor U4354 (N_4354,N_2473,N_31);
nor U4355 (N_4355,N_1327,N_703);
nand U4356 (N_4356,N_719,N_704);
and U4357 (N_4357,N_575,N_414);
nand U4358 (N_4358,N_1816,N_1990);
xnor U4359 (N_4359,N_619,N_571);
and U4360 (N_4360,N_729,N_2713);
nand U4361 (N_4361,N_178,N_895);
and U4362 (N_4362,N_2226,N_1592);
and U4363 (N_4363,N_1088,N_941);
nand U4364 (N_4364,N_94,N_505);
nand U4365 (N_4365,N_1609,N_2691);
and U4366 (N_4366,N_2077,N_2640);
xor U4367 (N_4367,N_938,N_1455);
and U4368 (N_4368,N_745,N_1844);
or U4369 (N_4369,N_2058,N_1554);
or U4370 (N_4370,N_2050,N_107);
xor U4371 (N_4371,N_2414,N_1916);
nand U4372 (N_4372,N_1929,N_574);
and U4373 (N_4373,N_1233,N_10);
nand U4374 (N_4374,N_2079,N_2329);
and U4375 (N_4375,N_583,N_831);
or U4376 (N_4376,N_1613,N_1020);
nand U4377 (N_4377,N_2464,N_188);
or U4378 (N_4378,N_1377,N_997);
and U4379 (N_4379,N_1680,N_2010);
and U4380 (N_4380,N_2521,N_2992);
or U4381 (N_4381,N_2947,N_978);
and U4382 (N_4382,N_2874,N_649);
and U4383 (N_4383,N_103,N_1672);
nor U4384 (N_4384,N_2855,N_2072);
or U4385 (N_4385,N_2757,N_153);
xnor U4386 (N_4386,N_2604,N_1748);
nand U4387 (N_4387,N_1565,N_2196);
or U4388 (N_4388,N_1962,N_931);
nand U4389 (N_4389,N_1084,N_2532);
or U4390 (N_4390,N_2126,N_655);
nor U4391 (N_4391,N_2701,N_909);
nand U4392 (N_4392,N_609,N_2916);
nor U4393 (N_4393,N_1786,N_1771);
nor U4394 (N_4394,N_2060,N_507);
nand U4395 (N_4395,N_1857,N_1441);
and U4396 (N_4396,N_1412,N_2016);
nor U4397 (N_4397,N_2020,N_2642);
nor U4398 (N_4398,N_2568,N_261);
nand U4399 (N_4399,N_1896,N_2834);
nand U4400 (N_4400,N_1161,N_2481);
nor U4401 (N_4401,N_498,N_2619);
nor U4402 (N_4402,N_2780,N_2366);
nand U4403 (N_4403,N_698,N_279);
nor U4404 (N_4404,N_2113,N_921);
or U4405 (N_4405,N_2801,N_2896);
and U4406 (N_4406,N_758,N_519);
and U4407 (N_4407,N_710,N_92);
and U4408 (N_4408,N_883,N_821);
nand U4409 (N_4409,N_2605,N_2044);
and U4410 (N_4410,N_2216,N_1569);
and U4411 (N_4411,N_1192,N_1264);
and U4412 (N_4412,N_550,N_2274);
xor U4413 (N_4413,N_711,N_171);
nor U4414 (N_4414,N_2475,N_1995);
nor U4415 (N_4415,N_1740,N_2754);
xor U4416 (N_4416,N_2557,N_2790);
nand U4417 (N_4417,N_2609,N_2235);
nand U4418 (N_4418,N_679,N_789);
and U4419 (N_4419,N_161,N_2546);
or U4420 (N_4420,N_1180,N_802);
nor U4421 (N_4421,N_1998,N_1525);
or U4422 (N_4422,N_1195,N_653);
or U4423 (N_4423,N_6,N_2076);
nor U4424 (N_4424,N_577,N_1950);
nor U4425 (N_4425,N_587,N_736);
xor U4426 (N_4426,N_2910,N_354);
and U4427 (N_4427,N_556,N_1783);
or U4428 (N_4428,N_2158,N_1836);
nor U4429 (N_4429,N_1992,N_2451);
or U4430 (N_4430,N_1757,N_2424);
nor U4431 (N_4431,N_1802,N_946);
nor U4432 (N_4432,N_1514,N_760);
nand U4433 (N_4433,N_1567,N_113);
and U4434 (N_4434,N_1694,N_1315);
nor U4435 (N_4435,N_2638,N_523);
and U4436 (N_4436,N_2132,N_2);
xnor U4437 (N_4437,N_2503,N_2268);
xor U4438 (N_4438,N_2458,N_454);
or U4439 (N_4439,N_2011,N_1111);
nand U4440 (N_4440,N_1690,N_1360);
xor U4441 (N_4441,N_2057,N_2828);
xnor U4442 (N_4442,N_1624,N_2513);
nand U4443 (N_4443,N_2383,N_28);
nor U4444 (N_4444,N_2038,N_1335);
nand U4445 (N_4445,N_1807,N_810);
xor U4446 (N_4446,N_1897,N_243);
or U4447 (N_4447,N_2861,N_37);
or U4448 (N_4448,N_2973,N_287);
nor U4449 (N_4449,N_2004,N_2247);
nor U4450 (N_4450,N_773,N_396);
nor U4451 (N_4451,N_2215,N_674);
xnor U4452 (N_4452,N_157,N_1434);
and U4453 (N_4453,N_317,N_267);
nor U4454 (N_4454,N_624,N_2981);
nor U4455 (N_4455,N_1228,N_2365);
or U4456 (N_4456,N_1606,N_2693);
or U4457 (N_4457,N_1864,N_1878);
xor U4458 (N_4458,N_1175,N_618);
xnor U4459 (N_4459,N_699,N_2762);
xor U4460 (N_4460,N_1205,N_1552);
and U4461 (N_4461,N_1575,N_735);
nor U4462 (N_4462,N_1310,N_1951);
and U4463 (N_4463,N_2396,N_1528);
xnor U4464 (N_4464,N_2721,N_837);
nand U4465 (N_4465,N_57,N_2745);
nand U4466 (N_4466,N_1354,N_957);
xnor U4467 (N_4467,N_2936,N_2592);
xor U4468 (N_4468,N_353,N_751);
nor U4469 (N_4469,N_2788,N_1164);
xor U4470 (N_4470,N_2676,N_1758);
nor U4471 (N_4471,N_967,N_560);
nand U4472 (N_4472,N_929,N_974);
or U4473 (N_4473,N_1938,N_544);
nand U4474 (N_4474,N_1144,N_1991);
or U4475 (N_4475,N_2858,N_1920);
and U4476 (N_4476,N_197,N_1336);
xnor U4477 (N_4477,N_2920,N_2877);
nor U4478 (N_4478,N_2765,N_443);
or U4479 (N_4479,N_985,N_1103);
or U4480 (N_4480,N_1813,N_81);
nand U4481 (N_4481,N_1764,N_212);
or U4482 (N_4482,N_1922,N_1940);
and U4483 (N_4483,N_2138,N_1870);
or U4484 (N_4484,N_2905,N_2971);
nor U4485 (N_4485,N_298,N_1633);
and U4486 (N_4486,N_2384,N_2859);
xor U4487 (N_4487,N_1713,N_390);
nand U4488 (N_4488,N_2975,N_963);
xor U4489 (N_4489,N_1754,N_1193);
and U4490 (N_4490,N_807,N_1823);
nand U4491 (N_4491,N_144,N_324);
xnor U4492 (N_4492,N_2477,N_825);
nand U4493 (N_4493,N_2943,N_1876);
or U4494 (N_4494,N_159,N_2265);
nor U4495 (N_4495,N_1720,N_1562);
and U4496 (N_4496,N_2156,N_222);
and U4497 (N_4497,N_2929,N_827);
nand U4498 (N_4498,N_14,N_1117);
nor U4499 (N_4499,N_2741,N_1397);
nand U4500 (N_4500,N_282,N_1171);
nand U4501 (N_4501,N_46,N_2336);
and U4502 (N_4502,N_2075,N_1584);
and U4503 (N_4503,N_984,N_136);
or U4504 (N_4504,N_1376,N_2733);
nor U4505 (N_4505,N_1605,N_1686);
nor U4506 (N_4506,N_29,N_2056);
and U4507 (N_4507,N_56,N_959);
nand U4508 (N_4508,N_1389,N_629);
nand U4509 (N_4509,N_1109,N_1316);
nand U4510 (N_4510,N_2396,N_1450);
nand U4511 (N_4511,N_921,N_2814);
nand U4512 (N_4512,N_319,N_95);
nand U4513 (N_4513,N_1661,N_1142);
nand U4514 (N_4514,N_2305,N_1928);
nand U4515 (N_4515,N_812,N_2137);
or U4516 (N_4516,N_2680,N_1879);
and U4517 (N_4517,N_2758,N_373);
xnor U4518 (N_4518,N_200,N_1186);
nand U4519 (N_4519,N_1018,N_1775);
or U4520 (N_4520,N_1935,N_2633);
xnor U4521 (N_4521,N_2629,N_874);
nand U4522 (N_4522,N_967,N_2609);
xor U4523 (N_4523,N_1093,N_1163);
and U4524 (N_4524,N_1488,N_179);
or U4525 (N_4525,N_139,N_2976);
or U4526 (N_4526,N_765,N_2577);
nor U4527 (N_4527,N_2119,N_2034);
and U4528 (N_4528,N_2180,N_801);
nand U4529 (N_4529,N_1847,N_1244);
nor U4530 (N_4530,N_2818,N_1540);
xor U4531 (N_4531,N_1044,N_1174);
and U4532 (N_4532,N_1195,N_2959);
or U4533 (N_4533,N_69,N_2249);
and U4534 (N_4534,N_65,N_2444);
xor U4535 (N_4535,N_321,N_2525);
xnor U4536 (N_4536,N_1085,N_2132);
xor U4537 (N_4537,N_2973,N_1504);
nand U4538 (N_4538,N_2059,N_1252);
or U4539 (N_4539,N_1167,N_2787);
or U4540 (N_4540,N_2002,N_14);
nor U4541 (N_4541,N_82,N_2186);
xnor U4542 (N_4542,N_2808,N_2147);
xor U4543 (N_4543,N_2678,N_1063);
and U4544 (N_4544,N_1613,N_493);
nor U4545 (N_4545,N_582,N_1048);
xnor U4546 (N_4546,N_527,N_1827);
xor U4547 (N_4547,N_1795,N_568);
nand U4548 (N_4548,N_423,N_893);
or U4549 (N_4549,N_821,N_1064);
and U4550 (N_4550,N_1328,N_300);
or U4551 (N_4551,N_2968,N_712);
or U4552 (N_4552,N_1673,N_2702);
and U4553 (N_4553,N_1786,N_2321);
nor U4554 (N_4554,N_2463,N_2256);
nand U4555 (N_4555,N_1327,N_1791);
nand U4556 (N_4556,N_1323,N_2683);
nand U4557 (N_4557,N_2261,N_2311);
and U4558 (N_4558,N_392,N_819);
nor U4559 (N_4559,N_275,N_1986);
nor U4560 (N_4560,N_1652,N_1598);
nor U4561 (N_4561,N_2719,N_607);
and U4562 (N_4562,N_1245,N_238);
nand U4563 (N_4563,N_2524,N_2759);
nand U4564 (N_4564,N_221,N_430);
nor U4565 (N_4565,N_2299,N_1661);
and U4566 (N_4566,N_2496,N_805);
and U4567 (N_4567,N_888,N_320);
or U4568 (N_4568,N_416,N_276);
and U4569 (N_4569,N_2429,N_2110);
nand U4570 (N_4570,N_1100,N_1161);
nor U4571 (N_4571,N_458,N_2018);
nor U4572 (N_4572,N_1986,N_2049);
and U4573 (N_4573,N_993,N_1439);
xor U4574 (N_4574,N_1156,N_891);
nand U4575 (N_4575,N_794,N_2793);
or U4576 (N_4576,N_1512,N_788);
nor U4577 (N_4577,N_2779,N_2089);
and U4578 (N_4578,N_400,N_1878);
nor U4579 (N_4579,N_889,N_821);
or U4580 (N_4580,N_72,N_1735);
or U4581 (N_4581,N_2225,N_2019);
xor U4582 (N_4582,N_360,N_1114);
xnor U4583 (N_4583,N_1477,N_2581);
or U4584 (N_4584,N_313,N_264);
nand U4585 (N_4585,N_2856,N_426);
and U4586 (N_4586,N_2385,N_2777);
nor U4587 (N_4587,N_834,N_429);
xor U4588 (N_4588,N_1447,N_2308);
and U4589 (N_4589,N_83,N_2503);
xnor U4590 (N_4590,N_565,N_2536);
or U4591 (N_4591,N_616,N_1143);
nand U4592 (N_4592,N_2478,N_2523);
nor U4593 (N_4593,N_1106,N_2293);
nand U4594 (N_4594,N_1299,N_2909);
nand U4595 (N_4595,N_1840,N_1337);
xor U4596 (N_4596,N_71,N_645);
and U4597 (N_4597,N_2028,N_621);
nor U4598 (N_4598,N_2409,N_1758);
nor U4599 (N_4599,N_2500,N_2029);
or U4600 (N_4600,N_2194,N_815);
nor U4601 (N_4601,N_274,N_934);
and U4602 (N_4602,N_1210,N_2762);
or U4603 (N_4603,N_1012,N_2172);
and U4604 (N_4604,N_1851,N_1805);
xor U4605 (N_4605,N_1208,N_994);
and U4606 (N_4606,N_2081,N_291);
nand U4607 (N_4607,N_2213,N_2210);
nor U4608 (N_4608,N_797,N_1370);
xor U4609 (N_4609,N_203,N_957);
and U4610 (N_4610,N_542,N_2052);
or U4611 (N_4611,N_197,N_1102);
nor U4612 (N_4612,N_1757,N_2521);
nor U4613 (N_4613,N_1821,N_1163);
or U4614 (N_4614,N_2804,N_376);
or U4615 (N_4615,N_113,N_615);
xnor U4616 (N_4616,N_1977,N_1283);
nor U4617 (N_4617,N_755,N_1426);
nand U4618 (N_4618,N_1605,N_2437);
nand U4619 (N_4619,N_1403,N_113);
and U4620 (N_4620,N_2078,N_1269);
nand U4621 (N_4621,N_2580,N_656);
nand U4622 (N_4622,N_1541,N_2638);
xnor U4623 (N_4623,N_1456,N_156);
and U4624 (N_4624,N_1995,N_324);
nand U4625 (N_4625,N_1559,N_2219);
nor U4626 (N_4626,N_1255,N_2014);
nor U4627 (N_4627,N_385,N_585);
xor U4628 (N_4628,N_741,N_2941);
or U4629 (N_4629,N_2468,N_1601);
nand U4630 (N_4630,N_2969,N_2869);
and U4631 (N_4631,N_2222,N_2395);
or U4632 (N_4632,N_2170,N_401);
and U4633 (N_4633,N_1506,N_2666);
and U4634 (N_4634,N_1850,N_782);
and U4635 (N_4635,N_204,N_494);
nor U4636 (N_4636,N_2683,N_1020);
and U4637 (N_4637,N_203,N_681);
xor U4638 (N_4638,N_1949,N_2272);
nand U4639 (N_4639,N_2968,N_2863);
nand U4640 (N_4640,N_1454,N_1048);
or U4641 (N_4641,N_698,N_2013);
nor U4642 (N_4642,N_2367,N_2701);
nor U4643 (N_4643,N_2845,N_1127);
nor U4644 (N_4644,N_2963,N_2011);
or U4645 (N_4645,N_550,N_842);
xnor U4646 (N_4646,N_1609,N_1463);
or U4647 (N_4647,N_398,N_687);
and U4648 (N_4648,N_2538,N_2065);
nand U4649 (N_4649,N_1560,N_276);
nand U4650 (N_4650,N_2945,N_2549);
or U4651 (N_4651,N_2935,N_2388);
nor U4652 (N_4652,N_11,N_359);
and U4653 (N_4653,N_2352,N_193);
xor U4654 (N_4654,N_1514,N_307);
nor U4655 (N_4655,N_1890,N_1378);
and U4656 (N_4656,N_625,N_1177);
nand U4657 (N_4657,N_1375,N_2148);
nor U4658 (N_4658,N_1500,N_449);
nor U4659 (N_4659,N_1169,N_201);
or U4660 (N_4660,N_1427,N_434);
nor U4661 (N_4661,N_2127,N_2406);
and U4662 (N_4662,N_691,N_1985);
xnor U4663 (N_4663,N_1742,N_1573);
nor U4664 (N_4664,N_2756,N_266);
nand U4665 (N_4665,N_751,N_2207);
and U4666 (N_4666,N_2791,N_1838);
and U4667 (N_4667,N_1420,N_616);
nor U4668 (N_4668,N_796,N_40);
nand U4669 (N_4669,N_1102,N_1133);
xnor U4670 (N_4670,N_474,N_910);
and U4671 (N_4671,N_2751,N_1617);
nand U4672 (N_4672,N_2788,N_562);
nand U4673 (N_4673,N_565,N_1473);
xnor U4674 (N_4674,N_2013,N_94);
nand U4675 (N_4675,N_1526,N_914);
nand U4676 (N_4676,N_1215,N_1351);
xnor U4677 (N_4677,N_2512,N_1468);
nand U4678 (N_4678,N_1671,N_1855);
and U4679 (N_4679,N_1102,N_132);
xnor U4680 (N_4680,N_2214,N_1829);
xor U4681 (N_4681,N_836,N_1268);
or U4682 (N_4682,N_1215,N_55);
and U4683 (N_4683,N_20,N_1279);
nand U4684 (N_4684,N_2317,N_504);
nor U4685 (N_4685,N_377,N_2705);
xor U4686 (N_4686,N_1068,N_1805);
or U4687 (N_4687,N_1559,N_4);
or U4688 (N_4688,N_2443,N_2033);
and U4689 (N_4689,N_1508,N_381);
nand U4690 (N_4690,N_1123,N_2346);
and U4691 (N_4691,N_593,N_663);
nand U4692 (N_4692,N_1908,N_127);
or U4693 (N_4693,N_1635,N_2953);
or U4694 (N_4694,N_2206,N_611);
nand U4695 (N_4695,N_813,N_1525);
and U4696 (N_4696,N_1927,N_1862);
xnor U4697 (N_4697,N_896,N_185);
and U4698 (N_4698,N_1919,N_1904);
xor U4699 (N_4699,N_2383,N_2064);
or U4700 (N_4700,N_2473,N_2812);
nor U4701 (N_4701,N_1317,N_2470);
nor U4702 (N_4702,N_2025,N_2838);
nand U4703 (N_4703,N_1122,N_536);
nor U4704 (N_4704,N_2198,N_706);
and U4705 (N_4705,N_625,N_2048);
nand U4706 (N_4706,N_769,N_1401);
nand U4707 (N_4707,N_2293,N_2647);
nand U4708 (N_4708,N_930,N_1592);
xnor U4709 (N_4709,N_33,N_1159);
and U4710 (N_4710,N_1061,N_2641);
nand U4711 (N_4711,N_1760,N_518);
xor U4712 (N_4712,N_2643,N_1980);
nand U4713 (N_4713,N_673,N_1325);
or U4714 (N_4714,N_127,N_128);
xnor U4715 (N_4715,N_946,N_2385);
and U4716 (N_4716,N_2674,N_2689);
nand U4717 (N_4717,N_2169,N_1521);
xor U4718 (N_4718,N_1982,N_1720);
nor U4719 (N_4719,N_759,N_2370);
nand U4720 (N_4720,N_58,N_2492);
nand U4721 (N_4721,N_651,N_1331);
nor U4722 (N_4722,N_1896,N_262);
nand U4723 (N_4723,N_2813,N_2245);
xor U4724 (N_4724,N_992,N_2084);
xnor U4725 (N_4725,N_1280,N_1220);
xor U4726 (N_4726,N_1674,N_1732);
xnor U4727 (N_4727,N_2819,N_2309);
or U4728 (N_4728,N_2259,N_1997);
nand U4729 (N_4729,N_280,N_2811);
or U4730 (N_4730,N_2842,N_962);
or U4731 (N_4731,N_837,N_1996);
nor U4732 (N_4732,N_1110,N_1191);
nand U4733 (N_4733,N_970,N_1852);
nor U4734 (N_4734,N_2536,N_913);
nand U4735 (N_4735,N_543,N_950);
nor U4736 (N_4736,N_2104,N_88);
or U4737 (N_4737,N_380,N_1583);
and U4738 (N_4738,N_2804,N_1649);
or U4739 (N_4739,N_488,N_2129);
or U4740 (N_4740,N_829,N_1381);
nand U4741 (N_4741,N_176,N_698);
nand U4742 (N_4742,N_2250,N_2316);
nand U4743 (N_4743,N_1541,N_331);
nand U4744 (N_4744,N_2349,N_2265);
xnor U4745 (N_4745,N_1106,N_2135);
nand U4746 (N_4746,N_1220,N_931);
and U4747 (N_4747,N_1,N_1744);
nand U4748 (N_4748,N_2014,N_183);
and U4749 (N_4749,N_631,N_2467);
nor U4750 (N_4750,N_202,N_1590);
nor U4751 (N_4751,N_1467,N_2783);
or U4752 (N_4752,N_94,N_2876);
or U4753 (N_4753,N_292,N_2602);
nand U4754 (N_4754,N_413,N_640);
or U4755 (N_4755,N_1556,N_2);
and U4756 (N_4756,N_2363,N_1884);
nand U4757 (N_4757,N_2478,N_1201);
nor U4758 (N_4758,N_23,N_1020);
or U4759 (N_4759,N_1810,N_2362);
nor U4760 (N_4760,N_2345,N_2971);
xnor U4761 (N_4761,N_714,N_561);
nor U4762 (N_4762,N_1534,N_1604);
or U4763 (N_4763,N_2546,N_651);
nor U4764 (N_4764,N_1663,N_1890);
nand U4765 (N_4765,N_1379,N_1565);
or U4766 (N_4766,N_605,N_2488);
nor U4767 (N_4767,N_237,N_2164);
nor U4768 (N_4768,N_1808,N_1412);
nor U4769 (N_4769,N_681,N_2069);
or U4770 (N_4770,N_2392,N_724);
or U4771 (N_4771,N_2884,N_2950);
nor U4772 (N_4772,N_81,N_766);
and U4773 (N_4773,N_1485,N_288);
xor U4774 (N_4774,N_759,N_1421);
and U4775 (N_4775,N_26,N_1633);
xnor U4776 (N_4776,N_1869,N_737);
or U4777 (N_4777,N_2644,N_406);
nor U4778 (N_4778,N_1809,N_738);
or U4779 (N_4779,N_1744,N_2592);
and U4780 (N_4780,N_2019,N_431);
xor U4781 (N_4781,N_2514,N_917);
or U4782 (N_4782,N_1436,N_2804);
or U4783 (N_4783,N_2080,N_1343);
nor U4784 (N_4784,N_380,N_1620);
xor U4785 (N_4785,N_543,N_743);
nor U4786 (N_4786,N_731,N_1552);
or U4787 (N_4787,N_1480,N_986);
or U4788 (N_4788,N_2567,N_625);
nor U4789 (N_4789,N_1667,N_47);
and U4790 (N_4790,N_1252,N_2764);
nand U4791 (N_4791,N_2554,N_2261);
or U4792 (N_4792,N_2488,N_1994);
and U4793 (N_4793,N_2836,N_1285);
xnor U4794 (N_4794,N_2666,N_611);
xor U4795 (N_4795,N_98,N_1269);
xor U4796 (N_4796,N_826,N_450);
and U4797 (N_4797,N_1383,N_1514);
and U4798 (N_4798,N_1711,N_2327);
nor U4799 (N_4799,N_2205,N_625);
nor U4800 (N_4800,N_2474,N_1475);
xnor U4801 (N_4801,N_485,N_2482);
and U4802 (N_4802,N_2598,N_75);
and U4803 (N_4803,N_644,N_2732);
or U4804 (N_4804,N_1851,N_94);
nand U4805 (N_4805,N_2861,N_127);
nor U4806 (N_4806,N_2116,N_2420);
or U4807 (N_4807,N_980,N_2771);
xor U4808 (N_4808,N_1724,N_2734);
xnor U4809 (N_4809,N_15,N_1003);
nand U4810 (N_4810,N_219,N_90);
xnor U4811 (N_4811,N_1942,N_2667);
xor U4812 (N_4812,N_809,N_747);
nand U4813 (N_4813,N_825,N_475);
nand U4814 (N_4814,N_570,N_1376);
or U4815 (N_4815,N_491,N_519);
or U4816 (N_4816,N_1989,N_1854);
nor U4817 (N_4817,N_1407,N_2800);
nand U4818 (N_4818,N_1034,N_2694);
and U4819 (N_4819,N_2649,N_2142);
and U4820 (N_4820,N_961,N_2686);
and U4821 (N_4821,N_2626,N_141);
xnor U4822 (N_4822,N_18,N_554);
xnor U4823 (N_4823,N_2560,N_2135);
or U4824 (N_4824,N_2219,N_212);
or U4825 (N_4825,N_1000,N_242);
nand U4826 (N_4826,N_1902,N_978);
nor U4827 (N_4827,N_531,N_2586);
nor U4828 (N_4828,N_2754,N_2315);
or U4829 (N_4829,N_1886,N_1858);
and U4830 (N_4830,N_2169,N_2362);
and U4831 (N_4831,N_2699,N_2104);
nor U4832 (N_4832,N_294,N_1396);
xnor U4833 (N_4833,N_368,N_432);
xnor U4834 (N_4834,N_336,N_960);
nor U4835 (N_4835,N_976,N_485);
and U4836 (N_4836,N_2195,N_261);
or U4837 (N_4837,N_2766,N_1746);
nand U4838 (N_4838,N_1304,N_782);
or U4839 (N_4839,N_1773,N_2217);
and U4840 (N_4840,N_444,N_837);
nand U4841 (N_4841,N_705,N_887);
nand U4842 (N_4842,N_973,N_2512);
and U4843 (N_4843,N_2461,N_601);
or U4844 (N_4844,N_847,N_501);
and U4845 (N_4845,N_2037,N_1162);
nand U4846 (N_4846,N_765,N_2877);
and U4847 (N_4847,N_2672,N_886);
or U4848 (N_4848,N_1991,N_367);
and U4849 (N_4849,N_2666,N_622);
and U4850 (N_4850,N_1921,N_1079);
xor U4851 (N_4851,N_231,N_2908);
xor U4852 (N_4852,N_22,N_1595);
and U4853 (N_4853,N_896,N_2428);
or U4854 (N_4854,N_1078,N_2490);
nand U4855 (N_4855,N_2467,N_2239);
nor U4856 (N_4856,N_1580,N_1702);
nor U4857 (N_4857,N_53,N_2880);
nand U4858 (N_4858,N_2128,N_734);
and U4859 (N_4859,N_190,N_278);
nor U4860 (N_4860,N_1770,N_356);
and U4861 (N_4861,N_1969,N_2042);
xor U4862 (N_4862,N_1052,N_986);
and U4863 (N_4863,N_573,N_1713);
nand U4864 (N_4864,N_1621,N_1301);
nor U4865 (N_4865,N_1550,N_806);
xor U4866 (N_4866,N_1773,N_1932);
nor U4867 (N_4867,N_1529,N_2104);
nand U4868 (N_4868,N_933,N_1870);
or U4869 (N_4869,N_998,N_2257);
nand U4870 (N_4870,N_2331,N_2241);
nand U4871 (N_4871,N_703,N_286);
or U4872 (N_4872,N_2181,N_40);
xnor U4873 (N_4873,N_2354,N_409);
nand U4874 (N_4874,N_2755,N_2862);
nand U4875 (N_4875,N_1109,N_960);
nor U4876 (N_4876,N_1337,N_2516);
nand U4877 (N_4877,N_2006,N_585);
or U4878 (N_4878,N_1903,N_2255);
or U4879 (N_4879,N_2367,N_553);
and U4880 (N_4880,N_2655,N_19);
or U4881 (N_4881,N_1002,N_452);
nor U4882 (N_4882,N_1757,N_1199);
and U4883 (N_4883,N_901,N_2566);
or U4884 (N_4884,N_681,N_108);
nor U4885 (N_4885,N_2654,N_2317);
and U4886 (N_4886,N_179,N_1659);
nor U4887 (N_4887,N_129,N_2277);
nand U4888 (N_4888,N_1780,N_1464);
nor U4889 (N_4889,N_1846,N_584);
nor U4890 (N_4890,N_2482,N_101);
or U4891 (N_4891,N_1233,N_1584);
nand U4892 (N_4892,N_1106,N_700);
nor U4893 (N_4893,N_441,N_1823);
xnor U4894 (N_4894,N_2104,N_1005);
or U4895 (N_4895,N_935,N_1201);
xor U4896 (N_4896,N_2277,N_2084);
nor U4897 (N_4897,N_1797,N_530);
and U4898 (N_4898,N_1445,N_1348);
and U4899 (N_4899,N_648,N_1466);
nand U4900 (N_4900,N_222,N_2800);
or U4901 (N_4901,N_1006,N_209);
nand U4902 (N_4902,N_927,N_946);
and U4903 (N_4903,N_348,N_1837);
xor U4904 (N_4904,N_941,N_2825);
nand U4905 (N_4905,N_1297,N_446);
xor U4906 (N_4906,N_945,N_1201);
xor U4907 (N_4907,N_240,N_1430);
xnor U4908 (N_4908,N_526,N_1015);
or U4909 (N_4909,N_2116,N_388);
or U4910 (N_4910,N_1427,N_2154);
or U4911 (N_4911,N_1478,N_2930);
nand U4912 (N_4912,N_312,N_2804);
xnor U4913 (N_4913,N_1895,N_1487);
and U4914 (N_4914,N_70,N_741);
nand U4915 (N_4915,N_1686,N_1851);
nand U4916 (N_4916,N_1947,N_2085);
xor U4917 (N_4917,N_2466,N_2128);
and U4918 (N_4918,N_1800,N_1482);
or U4919 (N_4919,N_2987,N_436);
nor U4920 (N_4920,N_46,N_2101);
nand U4921 (N_4921,N_1720,N_26);
nand U4922 (N_4922,N_597,N_257);
nor U4923 (N_4923,N_662,N_1539);
nor U4924 (N_4924,N_800,N_772);
nand U4925 (N_4925,N_858,N_2130);
nor U4926 (N_4926,N_1276,N_1151);
or U4927 (N_4927,N_2028,N_111);
nand U4928 (N_4928,N_21,N_2182);
nand U4929 (N_4929,N_2424,N_179);
and U4930 (N_4930,N_2452,N_1237);
and U4931 (N_4931,N_1858,N_44);
or U4932 (N_4932,N_803,N_2340);
nor U4933 (N_4933,N_327,N_1087);
nand U4934 (N_4934,N_2953,N_438);
nand U4935 (N_4935,N_2378,N_321);
xor U4936 (N_4936,N_667,N_899);
nor U4937 (N_4937,N_735,N_322);
or U4938 (N_4938,N_1894,N_790);
and U4939 (N_4939,N_2287,N_1674);
nor U4940 (N_4940,N_492,N_1725);
or U4941 (N_4941,N_676,N_135);
and U4942 (N_4942,N_900,N_10);
and U4943 (N_4943,N_1259,N_2427);
and U4944 (N_4944,N_2148,N_1963);
nor U4945 (N_4945,N_2222,N_1147);
nand U4946 (N_4946,N_478,N_1690);
nand U4947 (N_4947,N_624,N_2116);
xnor U4948 (N_4948,N_702,N_1776);
xor U4949 (N_4949,N_2112,N_489);
nor U4950 (N_4950,N_2102,N_174);
nand U4951 (N_4951,N_1770,N_2256);
or U4952 (N_4952,N_1551,N_1797);
and U4953 (N_4953,N_2893,N_2655);
nor U4954 (N_4954,N_106,N_455);
xnor U4955 (N_4955,N_1233,N_1587);
xnor U4956 (N_4956,N_1043,N_2407);
or U4957 (N_4957,N_729,N_502);
or U4958 (N_4958,N_1182,N_1705);
and U4959 (N_4959,N_798,N_1076);
and U4960 (N_4960,N_796,N_518);
and U4961 (N_4961,N_175,N_672);
nand U4962 (N_4962,N_1760,N_1402);
nand U4963 (N_4963,N_2687,N_2879);
and U4964 (N_4964,N_2499,N_1701);
or U4965 (N_4965,N_2459,N_1538);
or U4966 (N_4966,N_1505,N_2684);
nor U4967 (N_4967,N_545,N_1761);
xor U4968 (N_4968,N_2309,N_2120);
xor U4969 (N_4969,N_786,N_2575);
nor U4970 (N_4970,N_2741,N_849);
or U4971 (N_4971,N_958,N_2567);
and U4972 (N_4972,N_224,N_2725);
xnor U4973 (N_4973,N_1715,N_1935);
or U4974 (N_4974,N_1279,N_896);
or U4975 (N_4975,N_1500,N_335);
and U4976 (N_4976,N_238,N_1718);
nor U4977 (N_4977,N_74,N_2255);
and U4978 (N_4978,N_2667,N_2473);
nand U4979 (N_4979,N_2257,N_842);
or U4980 (N_4980,N_1992,N_221);
and U4981 (N_4981,N_4,N_371);
and U4982 (N_4982,N_2516,N_2409);
and U4983 (N_4983,N_1980,N_712);
or U4984 (N_4984,N_1211,N_1154);
xnor U4985 (N_4985,N_1123,N_1224);
or U4986 (N_4986,N_748,N_11);
and U4987 (N_4987,N_1523,N_2577);
nand U4988 (N_4988,N_1652,N_1836);
xor U4989 (N_4989,N_1102,N_2317);
or U4990 (N_4990,N_1646,N_1720);
nor U4991 (N_4991,N_2487,N_949);
nand U4992 (N_4992,N_1697,N_2397);
or U4993 (N_4993,N_2249,N_866);
nand U4994 (N_4994,N_2377,N_816);
or U4995 (N_4995,N_1411,N_1226);
nand U4996 (N_4996,N_1531,N_929);
and U4997 (N_4997,N_161,N_2020);
nor U4998 (N_4998,N_2245,N_1303);
nor U4999 (N_4999,N_338,N_2458);
nor U5000 (N_5000,N_2511,N_2626);
xnor U5001 (N_5001,N_2859,N_2017);
and U5002 (N_5002,N_152,N_697);
and U5003 (N_5003,N_1477,N_1138);
and U5004 (N_5004,N_544,N_2473);
xor U5005 (N_5005,N_759,N_2738);
xnor U5006 (N_5006,N_2916,N_117);
nand U5007 (N_5007,N_208,N_2423);
or U5008 (N_5008,N_3,N_895);
nor U5009 (N_5009,N_343,N_813);
xnor U5010 (N_5010,N_2997,N_1001);
nor U5011 (N_5011,N_2068,N_531);
or U5012 (N_5012,N_2982,N_1693);
nand U5013 (N_5013,N_1913,N_544);
xnor U5014 (N_5014,N_1509,N_1355);
and U5015 (N_5015,N_1875,N_2641);
nor U5016 (N_5016,N_2950,N_1344);
and U5017 (N_5017,N_958,N_251);
nor U5018 (N_5018,N_32,N_2022);
nand U5019 (N_5019,N_2557,N_1312);
xnor U5020 (N_5020,N_1154,N_457);
and U5021 (N_5021,N_1344,N_1123);
nand U5022 (N_5022,N_293,N_2011);
or U5023 (N_5023,N_657,N_1834);
xnor U5024 (N_5024,N_2325,N_355);
nor U5025 (N_5025,N_2193,N_2941);
nor U5026 (N_5026,N_1417,N_2477);
xor U5027 (N_5027,N_1589,N_186);
or U5028 (N_5028,N_1380,N_1318);
or U5029 (N_5029,N_504,N_952);
nor U5030 (N_5030,N_780,N_2828);
nand U5031 (N_5031,N_2083,N_967);
nand U5032 (N_5032,N_692,N_2074);
and U5033 (N_5033,N_703,N_1473);
or U5034 (N_5034,N_260,N_1665);
nand U5035 (N_5035,N_1446,N_777);
and U5036 (N_5036,N_2209,N_2980);
or U5037 (N_5037,N_2453,N_137);
and U5038 (N_5038,N_2771,N_2545);
nand U5039 (N_5039,N_45,N_85);
nand U5040 (N_5040,N_2948,N_1152);
nor U5041 (N_5041,N_997,N_1288);
or U5042 (N_5042,N_1756,N_753);
nand U5043 (N_5043,N_946,N_1708);
nand U5044 (N_5044,N_502,N_2683);
or U5045 (N_5045,N_2656,N_2264);
or U5046 (N_5046,N_230,N_2507);
nand U5047 (N_5047,N_2956,N_2831);
and U5048 (N_5048,N_664,N_2659);
nand U5049 (N_5049,N_1467,N_2618);
nor U5050 (N_5050,N_49,N_537);
or U5051 (N_5051,N_2908,N_2815);
or U5052 (N_5052,N_426,N_1069);
xor U5053 (N_5053,N_2208,N_1218);
or U5054 (N_5054,N_1867,N_912);
nand U5055 (N_5055,N_198,N_2555);
and U5056 (N_5056,N_628,N_974);
nor U5057 (N_5057,N_2928,N_102);
and U5058 (N_5058,N_2950,N_2202);
xor U5059 (N_5059,N_1762,N_2459);
xor U5060 (N_5060,N_2982,N_208);
and U5061 (N_5061,N_2230,N_2559);
xnor U5062 (N_5062,N_2679,N_1137);
xor U5063 (N_5063,N_1083,N_1878);
xor U5064 (N_5064,N_2914,N_1723);
xnor U5065 (N_5065,N_1749,N_2889);
and U5066 (N_5066,N_1844,N_243);
nand U5067 (N_5067,N_997,N_2976);
or U5068 (N_5068,N_611,N_2283);
xnor U5069 (N_5069,N_617,N_879);
xnor U5070 (N_5070,N_588,N_2463);
or U5071 (N_5071,N_2454,N_2444);
xor U5072 (N_5072,N_1186,N_1542);
nor U5073 (N_5073,N_2883,N_2146);
xor U5074 (N_5074,N_2256,N_1906);
or U5075 (N_5075,N_1736,N_1947);
nand U5076 (N_5076,N_2588,N_2521);
nand U5077 (N_5077,N_2662,N_51);
nand U5078 (N_5078,N_2936,N_87);
and U5079 (N_5079,N_1252,N_992);
nor U5080 (N_5080,N_2605,N_2661);
nand U5081 (N_5081,N_2325,N_780);
nor U5082 (N_5082,N_2812,N_1908);
nor U5083 (N_5083,N_2461,N_2171);
nand U5084 (N_5084,N_427,N_1506);
nand U5085 (N_5085,N_804,N_1321);
and U5086 (N_5086,N_2955,N_1426);
xnor U5087 (N_5087,N_2356,N_2366);
xnor U5088 (N_5088,N_2873,N_294);
xor U5089 (N_5089,N_2721,N_281);
xor U5090 (N_5090,N_766,N_1870);
xnor U5091 (N_5091,N_1404,N_2404);
or U5092 (N_5092,N_65,N_169);
nor U5093 (N_5093,N_2195,N_2063);
or U5094 (N_5094,N_12,N_1517);
nand U5095 (N_5095,N_1701,N_1829);
or U5096 (N_5096,N_1811,N_2519);
xor U5097 (N_5097,N_2043,N_2450);
nand U5098 (N_5098,N_1362,N_102);
and U5099 (N_5099,N_971,N_1468);
nor U5100 (N_5100,N_2150,N_1327);
or U5101 (N_5101,N_1922,N_2881);
nor U5102 (N_5102,N_2261,N_2672);
nor U5103 (N_5103,N_712,N_1623);
and U5104 (N_5104,N_1654,N_236);
and U5105 (N_5105,N_1638,N_939);
and U5106 (N_5106,N_383,N_502);
or U5107 (N_5107,N_377,N_2207);
or U5108 (N_5108,N_978,N_2282);
and U5109 (N_5109,N_587,N_2701);
nor U5110 (N_5110,N_1292,N_2242);
and U5111 (N_5111,N_778,N_2583);
nand U5112 (N_5112,N_1201,N_2609);
and U5113 (N_5113,N_621,N_2807);
or U5114 (N_5114,N_2092,N_2832);
nand U5115 (N_5115,N_2510,N_538);
xnor U5116 (N_5116,N_734,N_2718);
xor U5117 (N_5117,N_389,N_2102);
nor U5118 (N_5118,N_2634,N_1630);
nand U5119 (N_5119,N_202,N_1978);
and U5120 (N_5120,N_908,N_2631);
xnor U5121 (N_5121,N_2124,N_1008);
nor U5122 (N_5122,N_2389,N_823);
nor U5123 (N_5123,N_908,N_2842);
nor U5124 (N_5124,N_845,N_2147);
nand U5125 (N_5125,N_2703,N_936);
nor U5126 (N_5126,N_2417,N_2221);
nor U5127 (N_5127,N_1578,N_1487);
nor U5128 (N_5128,N_1170,N_1047);
nor U5129 (N_5129,N_1828,N_2656);
xnor U5130 (N_5130,N_29,N_2535);
nor U5131 (N_5131,N_2572,N_1612);
nor U5132 (N_5132,N_2783,N_2774);
nand U5133 (N_5133,N_1407,N_1124);
or U5134 (N_5134,N_2352,N_212);
xor U5135 (N_5135,N_2112,N_2660);
nor U5136 (N_5136,N_925,N_5);
nand U5137 (N_5137,N_1794,N_1230);
nor U5138 (N_5138,N_1605,N_259);
xnor U5139 (N_5139,N_2131,N_1847);
xnor U5140 (N_5140,N_2710,N_1628);
or U5141 (N_5141,N_2075,N_723);
nand U5142 (N_5142,N_1116,N_2832);
and U5143 (N_5143,N_2385,N_1826);
or U5144 (N_5144,N_502,N_458);
nand U5145 (N_5145,N_1792,N_2892);
nand U5146 (N_5146,N_614,N_535);
nor U5147 (N_5147,N_1463,N_2314);
or U5148 (N_5148,N_668,N_1828);
nand U5149 (N_5149,N_24,N_1812);
xnor U5150 (N_5150,N_1050,N_736);
nor U5151 (N_5151,N_435,N_2507);
nand U5152 (N_5152,N_863,N_2418);
nand U5153 (N_5153,N_2017,N_2554);
or U5154 (N_5154,N_2227,N_2872);
nand U5155 (N_5155,N_366,N_2730);
xor U5156 (N_5156,N_2963,N_2169);
and U5157 (N_5157,N_1527,N_400);
xor U5158 (N_5158,N_921,N_1379);
and U5159 (N_5159,N_1123,N_255);
or U5160 (N_5160,N_445,N_919);
nand U5161 (N_5161,N_1306,N_2244);
or U5162 (N_5162,N_2048,N_1998);
or U5163 (N_5163,N_2645,N_1691);
nand U5164 (N_5164,N_627,N_1678);
nand U5165 (N_5165,N_957,N_300);
or U5166 (N_5166,N_1272,N_1298);
nand U5167 (N_5167,N_1923,N_1177);
nand U5168 (N_5168,N_2704,N_2995);
xor U5169 (N_5169,N_2118,N_1540);
nand U5170 (N_5170,N_2494,N_1353);
or U5171 (N_5171,N_816,N_1055);
nand U5172 (N_5172,N_986,N_1976);
and U5173 (N_5173,N_854,N_381);
nand U5174 (N_5174,N_576,N_2481);
or U5175 (N_5175,N_1124,N_2523);
xnor U5176 (N_5176,N_2848,N_1994);
nand U5177 (N_5177,N_583,N_1720);
nand U5178 (N_5178,N_1638,N_1384);
nor U5179 (N_5179,N_1857,N_1673);
nand U5180 (N_5180,N_2012,N_2101);
and U5181 (N_5181,N_1176,N_922);
and U5182 (N_5182,N_153,N_1826);
nor U5183 (N_5183,N_39,N_1410);
nor U5184 (N_5184,N_74,N_2752);
or U5185 (N_5185,N_1955,N_1252);
and U5186 (N_5186,N_506,N_2321);
or U5187 (N_5187,N_14,N_2738);
and U5188 (N_5188,N_1318,N_1835);
or U5189 (N_5189,N_1407,N_142);
and U5190 (N_5190,N_1738,N_2610);
or U5191 (N_5191,N_1757,N_2651);
nand U5192 (N_5192,N_2813,N_2068);
xor U5193 (N_5193,N_1732,N_2803);
or U5194 (N_5194,N_1854,N_1028);
nor U5195 (N_5195,N_2847,N_2057);
and U5196 (N_5196,N_175,N_2549);
and U5197 (N_5197,N_2058,N_2884);
and U5198 (N_5198,N_1854,N_2779);
nor U5199 (N_5199,N_2122,N_1916);
nor U5200 (N_5200,N_1818,N_372);
xor U5201 (N_5201,N_2054,N_1959);
or U5202 (N_5202,N_173,N_882);
xor U5203 (N_5203,N_1664,N_1499);
and U5204 (N_5204,N_1307,N_1039);
nor U5205 (N_5205,N_2519,N_143);
and U5206 (N_5206,N_2892,N_1248);
or U5207 (N_5207,N_2673,N_578);
nand U5208 (N_5208,N_6,N_2011);
nor U5209 (N_5209,N_1255,N_1231);
xnor U5210 (N_5210,N_682,N_2460);
xnor U5211 (N_5211,N_44,N_2291);
xnor U5212 (N_5212,N_1147,N_1619);
xnor U5213 (N_5213,N_80,N_2527);
or U5214 (N_5214,N_1497,N_1059);
or U5215 (N_5215,N_1460,N_2904);
and U5216 (N_5216,N_762,N_1673);
nand U5217 (N_5217,N_1778,N_1627);
and U5218 (N_5218,N_1082,N_2317);
and U5219 (N_5219,N_2029,N_2196);
xor U5220 (N_5220,N_2524,N_627);
or U5221 (N_5221,N_1952,N_1327);
nor U5222 (N_5222,N_1013,N_158);
nand U5223 (N_5223,N_293,N_1769);
or U5224 (N_5224,N_554,N_1900);
and U5225 (N_5225,N_323,N_482);
and U5226 (N_5226,N_2378,N_2636);
nor U5227 (N_5227,N_702,N_1599);
nand U5228 (N_5228,N_1836,N_1474);
nand U5229 (N_5229,N_1167,N_2485);
nand U5230 (N_5230,N_1362,N_827);
and U5231 (N_5231,N_1868,N_1559);
and U5232 (N_5232,N_2639,N_2924);
xnor U5233 (N_5233,N_2846,N_2835);
nor U5234 (N_5234,N_808,N_158);
or U5235 (N_5235,N_2285,N_2826);
nand U5236 (N_5236,N_1454,N_2182);
or U5237 (N_5237,N_262,N_677);
xnor U5238 (N_5238,N_338,N_2585);
xnor U5239 (N_5239,N_1141,N_2263);
nor U5240 (N_5240,N_197,N_1201);
and U5241 (N_5241,N_2448,N_370);
xor U5242 (N_5242,N_82,N_2047);
xor U5243 (N_5243,N_2475,N_768);
xnor U5244 (N_5244,N_2138,N_2748);
or U5245 (N_5245,N_1028,N_1073);
or U5246 (N_5246,N_1654,N_816);
xor U5247 (N_5247,N_1634,N_2162);
or U5248 (N_5248,N_2729,N_2656);
and U5249 (N_5249,N_45,N_1276);
nand U5250 (N_5250,N_2272,N_960);
xor U5251 (N_5251,N_1654,N_1658);
and U5252 (N_5252,N_1870,N_255);
xor U5253 (N_5253,N_2359,N_274);
or U5254 (N_5254,N_1359,N_2419);
nor U5255 (N_5255,N_2199,N_2840);
or U5256 (N_5256,N_832,N_622);
nand U5257 (N_5257,N_148,N_2339);
nor U5258 (N_5258,N_2622,N_1781);
and U5259 (N_5259,N_573,N_2390);
xor U5260 (N_5260,N_838,N_2693);
nor U5261 (N_5261,N_607,N_1110);
nor U5262 (N_5262,N_2023,N_2478);
and U5263 (N_5263,N_1170,N_291);
and U5264 (N_5264,N_2022,N_187);
nor U5265 (N_5265,N_606,N_2217);
nor U5266 (N_5266,N_2469,N_1845);
xnor U5267 (N_5267,N_2405,N_2632);
or U5268 (N_5268,N_467,N_2739);
nor U5269 (N_5269,N_1409,N_2794);
nor U5270 (N_5270,N_204,N_125);
nand U5271 (N_5271,N_210,N_1931);
xor U5272 (N_5272,N_1315,N_1037);
nand U5273 (N_5273,N_2268,N_675);
nand U5274 (N_5274,N_1796,N_1652);
and U5275 (N_5275,N_2714,N_477);
or U5276 (N_5276,N_779,N_375);
xnor U5277 (N_5277,N_1380,N_1427);
nand U5278 (N_5278,N_1743,N_2904);
nor U5279 (N_5279,N_1760,N_1185);
nand U5280 (N_5280,N_2758,N_2307);
and U5281 (N_5281,N_1067,N_820);
nor U5282 (N_5282,N_517,N_1483);
nand U5283 (N_5283,N_1896,N_2120);
nor U5284 (N_5284,N_1081,N_2623);
nor U5285 (N_5285,N_866,N_2340);
nor U5286 (N_5286,N_2999,N_2184);
and U5287 (N_5287,N_359,N_1637);
or U5288 (N_5288,N_357,N_1256);
or U5289 (N_5289,N_2925,N_2951);
and U5290 (N_5290,N_2542,N_1169);
xnor U5291 (N_5291,N_2990,N_2484);
or U5292 (N_5292,N_581,N_2394);
and U5293 (N_5293,N_1766,N_678);
nand U5294 (N_5294,N_1458,N_2061);
and U5295 (N_5295,N_1748,N_1481);
and U5296 (N_5296,N_2839,N_1987);
xor U5297 (N_5297,N_1892,N_2905);
nor U5298 (N_5298,N_588,N_2898);
or U5299 (N_5299,N_915,N_2772);
and U5300 (N_5300,N_2661,N_687);
and U5301 (N_5301,N_939,N_742);
or U5302 (N_5302,N_787,N_745);
nor U5303 (N_5303,N_578,N_2055);
xnor U5304 (N_5304,N_1037,N_784);
nor U5305 (N_5305,N_597,N_1800);
xnor U5306 (N_5306,N_1896,N_426);
nand U5307 (N_5307,N_2590,N_259);
nor U5308 (N_5308,N_81,N_964);
or U5309 (N_5309,N_1308,N_173);
nor U5310 (N_5310,N_125,N_2938);
and U5311 (N_5311,N_278,N_900);
nand U5312 (N_5312,N_1831,N_2427);
xnor U5313 (N_5313,N_802,N_599);
nor U5314 (N_5314,N_1164,N_2558);
or U5315 (N_5315,N_442,N_525);
nand U5316 (N_5316,N_811,N_158);
nor U5317 (N_5317,N_1503,N_839);
or U5318 (N_5318,N_2021,N_1181);
nand U5319 (N_5319,N_1287,N_961);
nand U5320 (N_5320,N_1763,N_1442);
or U5321 (N_5321,N_384,N_215);
and U5322 (N_5322,N_2195,N_1067);
nand U5323 (N_5323,N_328,N_340);
xor U5324 (N_5324,N_1431,N_207);
or U5325 (N_5325,N_399,N_2161);
and U5326 (N_5326,N_464,N_1805);
and U5327 (N_5327,N_386,N_1908);
xor U5328 (N_5328,N_1351,N_451);
nor U5329 (N_5329,N_1317,N_2819);
nand U5330 (N_5330,N_375,N_1736);
and U5331 (N_5331,N_1241,N_2809);
nor U5332 (N_5332,N_1032,N_773);
nor U5333 (N_5333,N_1232,N_1624);
or U5334 (N_5334,N_321,N_960);
xor U5335 (N_5335,N_2867,N_573);
xor U5336 (N_5336,N_2470,N_319);
nand U5337 (N_5337,N_2556,N_2843);
xor U5338 (N_5338,N_325,N_2038);
and U5339 (N_5339,N_1906,N_517);
xnor U5340 (N_5340,N_1706,N_470);
nor U5341 (N_5341,N_2060,N_371);
nor U5342 (N_5342,N_89,N_540);
and U5343 (N_5343,N_1827,N_2658);
and U5344 (N_5344,N_1616,N_351);
xor U5345 (N_5345,N_1068,N_1793);
xnor U5346 (N_5346,N_144,N_545);
or U5347 (N_5347,N_2318,N_870);
xnor U5348 (N_5348,N_2865,N_752);
nor U5349 (N_5349,N_1112,N_1040);
nand U5350 (N_5350,N_2332,N_2839);
xor U5351 (N_5351,N_1869,N_2621);
or U5352 (N_5352,N_805,N_2335);
nand U5353 (N_5353,N_1254,N_2635);
nand U5354 (N_5354,N_1960,N_2819);
and U5355 (N_5355,N_2295,N_2359);
nand U5356 (N_5356,N_708,N_1070);
xor U5357 (N_5357,N_1313,N_450);
or U5358 (N_5358,N_378,N_2178);
and U5359 (N_5359,N_1346,N_2127);
nor U5360 (N_5360,N_1959,N_505);
nor U5361 (N_5361,N_2972,N_1318);
xnor U5362 (N_5362,N_2881,N_124);
nor U5363 (N_5363,N_474,N_2881);
nor U5364 (N_5364,N_2091,N_1324);
nand U5365 (N_5365,N_958,N_356);
and U5366 (N_5366,N_1615,N_2063);
nand U5367 (N_5367,N_801,N_1472);
nor U5368 (N_5368,N_824,N_603);
xnor U5369 (N_5369,N_231,N_177);
or U5370 (N_5370,N_278,N_1960);
and U5371 (N_5371,N_2198,N_1657);
or U5372 (N_5372,N_793,N_1433);
nand U5373 (N_5373,N_666,N_2389);
and U5374 (N_5374,N_62,N_2009);
and U5375 (N_5375,N_1533,N_1731);
nand U5376 (N_5376,N_1334,N_157);
xnor U5377 (N_5377,N_474,N_167);
and U5378 (N_5378,N_2860,N_990);
and U5379 (N_5379,N_27,N_1091);
xnor U5380 (N_5380,N_1778,N_442);
or U5381 (N_5381,N_2368,N_440);
xnor U5382 (N_5382,N_1685,N_2564);
xor U5383 (N_5383,N_2269,N_469);
nor U5384 (N_5384,N_1378,N_1092);
nor U5385 (N_5385,N_128,N_2731);
nand U5386 (N_5386,N_420,N_831);
and U5387 (N_5387,N_2627,N_2662);
nand U5388 (N_5388,N_2419,N_2086);
xnor U5389 (N_5389,N_2038,N_2438);
and U5390 (N_5390,N_1493,N_2413);
nand U5391 (N_5391,N_897,N_2752);
and U5392 (N_5392,N_900,N_728);
xnor U5393 (N_5393,N_1524,N_1006);
and U5394 (N_5394,N_1476,N_2825);
and U5395 (N_5395,N_460,N_2453);
nand U5396 (N_5396,N_2097,N_1683);
or U5397 (N_5397,N_2003,N_2013);
xnor U5398 (N_5398,N_1203,N_809);
xor U5399 (N_5399,N_2104,N_526);
and U5400 (N_5400,N_974,N_2774);
nor U5401 (N_5401,N_1810,N_2041);
and U5402 (N_5402,N_826,N_365);
nand U5403 (N_5403,N_2257,N_1353);
nor U5404 (N_5404,N_695,N_2872);
xnor U5405 (N_5405,N_2676,N_858);
nor U5406 (N_5406,N_2433,N_1518);
and U5407 (N_5407,N_1283,N_1021);
nor U5408 (N_5408,N_329,N_2263);
nand U5409 (N_5409,N_220,N_1720);
and U5410 (N_5410,N_2004,N_2528);
or U5411 (N_5411,N_1011,N_849);
xnor U5412 (N_5412,N_711,N_1186);
and U5413 (N_5413,N_1720,N_1478);
nand U5414 (N_5414,N_2104,N_1969);
nand U5415 (N_5415,N_2383,N_2048);
nand U5416 (N_5416,N_1148,N_176);
nor U5417 (N_5417,N_1571,N_916);
nand U5418 (N_5418,N_1194,N_2456);
nor U5419 (N_5419,N_2598,N_1856);
and U5420 (N_5420,N_184,N_2588);
and U5421 (N_5421,N_1940,N_1336);
or U5422 (N_5422,N_1641,N_2524);
xor U5423 (N_5423,N_793,N_1517);
nor U5424 (N_5424,N_2976,N_998);
xnor U5425 (N_5425,N_450,N_1058);
nand U5426 (N_5426,N_2045,N_1245);
and U5427 (N_5427,N_1330,N_15);
and U5428 (N_5428,N_1478,N_1667);
or U5429 (N_5429,N_541,N_1304);
nor U5430 (N_5430,N_460,N_1876);
nand U5431 (N_5431,N_1114,N_1949);
or U5432 (N_5432,N_2671,N_1694);
nor U5433 (N_5433,N_116,N_2008);
or U5434 (N_5434,N_961,N_118);
nor U5435 (N_5435,N_2090,N_1068);
and U5436 (N_5436,N_2796,N_1265);
xor U5437 (N_5437,N_2562,N_2091);
and U5438 (N_5438,N_1442,N_1144);
xor U5439 (N_5439,N_2267,N_1373);
or U5440 (N_5440,N_1947,N_2942);
nand U5441 (N_5441,N_2353,N_1171);
and U5442 (N_5442,N_618,N_2495);
or U5443 (N_5443,N_1593,N_634);
and U5444 (N_5444,N_2675,N_680);
xor U5445 (N_5445,N_1463,N_179);
or U5446 (N_5446,N_1093,N_1654);
nor U5447 (N_5447,N_1320,N_1746);
and U5448 (N_5448,N_883,N_2676);
or U5449 (N_5449,N_2717,N_2726);
nor U5450 (N_5450,N_1426,N_619);
nand U5451 (N_5451,N_2084,N_62);
and U5452 (N_5452,N_2292,N_859);
nand U5453 (N_5453,N_2518,N_1088);
or U5454 (N_5454,N_2840,N_1474);
and U5455 (N_5455,N_1539,N_1244);
nor U5456 (N_5456,N_1526,N_873);
xnor U5457 (N_5457,N_2157,N_1911);
nor U5458 (N_5458,N_2196,N_184);
xor U5459 (N_5459,N_1427,N_2433);
or U5460 (N_5460,N_2165,N_2841);
xor U5461 (N_5461,N_283,N_988);
nand U5462 (N_5462,N_1408,N_2281);
nand U5463 (N_5463,N_2889,N_2001);
nand U5464 (N_5464,N_1416,N_2403);
nor U5465 (N_5465,N_428,N_1823);
nor U5466 (N_5466,N_60,N_1901);
and U5467 (N_5467,N_698,N_1741);
and U5468 (N_5468,N_90,N_677);
nand U5469 (N_5469,N_1309,N_614);
and U5470 (N_5470,N_158,N_2177);
and U5471 (N_5471,N_1081,N_1211);
and U5472 (N_5472,N_1213,N_1243);
or U5473 (N_5473,N_300,N_233);
nor U5474 (N_5474,N_557,N_2165);
xor U5475 (N_5475,N_1059,N_2244);
or U5476 (N_5476,N_150,N_176);
nor U5477 (N_5477,N_1132,N_1355);
nand U5478 (N_5478,N_559,N_1158);
and U5479 (N_5479,N_2724,N_1582);
nor U5480 (N_5480,N_1882,N_1664);
or U5481 (N_5481,N_492,N_2663);
or U5482 (N_5482,N_2116,N_2738);
xnor U5483 (N_5483,N_2361,N_1981);
and U5484 (N_5484,N_1017,N_2324);
and U5485 (N_5485,N_2015,N_1565);
and U5486 (N_5486,N_693,N_589);
or U5487 (N_5487,N_253,N_2446);
nor U5488 (N_5488,N_2527,N_2231);
nand U5489 (N_5489,N_1256,N_813);
xor U5490 (N_5490,N_595,N_2152);
xor U5491 (N_5491,N_2434,N_1838);
nor U5492 (N_5492,N_1265,N_2775);
nor U5493 (N_5493,N_980,N_537);
xor U5494 (N_5494,N_1187,N_2916);
xor U5495 (N_5495,N_1019,N_1222);
nand U5496 (N_5496,N_753,N_78);
or U5497 (N_5497,N_1889,N_604);
nand U5498 (N_5498,N_198,N_2955);
nor U5499 (N_5499,N_2418,N_221);
and U5500 (N_5500,N_1946,N_2259);
or U5501 (N_5501,N_1509,N_257);
and U5502 (N_5502,N_2935,N_45);
xor U5503 (N_5503,N_2641,N_2882);
xor U5504 (N_5504,N_2520,N_346);
xor U5505 (N_5505,N_1423,N_2553);
and U5506 (N_5506,N_186,N_244);
nor U5507 (N_5507,N_1178,N_2058);
and U5508 (N_5508,N_1597,N_967);
nand U5509 (N_5509,N_1278,N_762);
nor U5510 (N_5510,N_814,N_659);
and U5511 (N_5511,N_677,N_2370);
or U5512 (N_5512,N_2549,N_631);
and U5513 (N_5513,N_725,N_42);
nand U5514 (N_5514,N_1371,N_409);
nor U5515 (N_5515,N_2158,N_1136);
xnor U5516 (N_5516,N_2158,N_2773);
xnor U5517 (N_5517,N_555,N_300);
and U5518 (N_5518,N_2863,N_1278);
or U5519 (N_5519,N_1743,N_2528);
nand U5520 (N_5520,N_992,N_1599);
nor U5521 (N_5521,N_2985,N_2588);
xor U5522 (N_5522,N_2291,N_2949);
and U5523 (N_5523,N_1492,N_1317);
and U5524 (N_5524,N_319,N_662);
xnor U5525 (N_5525,N_2665,N_1508);
nor U5526 (N_5526,N_66,N_303);
nor U5527 (N_5527,N_2133,N_2192);
or U5528 (N_5528,N_337,N_688);
or U5529 (N_5529,N_1332,N_2246);
xnor U5530 (N_5530,N_808,N_814);
nor U5531 (N_5531,N_813,N_1657);
and U5532 (N_5532,N_2370,N_315);
nor U5533 (N_5533,N_1615,N_2405);
or U5534 (N_5534,N_1634,N_162);
xor U5535 (N_5535,N_2926,N_1742);
nor U5536 (N_5536,N_485,N_2562);
and U5537 (N_5537,N_1659,N_2267);
nand U5538 (N_5538,N_490,N_20);
or U5539 (N_5539,N_833,N_2403);
nand U5540 (N_5540,N_639,N_661);
nand U5541 (N_5541,N_2979,N_2698);
nand U5542 (N_5542,N_216,N_1815);
nand U5543 (N_5543,N_1695,N_2819);
nand U5544 (N_5544,N_1280,N_491);
and U5545 (N_5545,N_1844,N_989);
or U5546 (N_5546,N_2750,N_2335);
nand U5547 (N_5547,N_2308,N_2005);
nand U5548 (N_5548,N_1399,N_1605);
and U5549 (N_5549,N_1295,N_988);
nand U5550 (N_5550,N_2323,N_1244);
xor U5551 (N_5551,N_754,N_558);
nand U5552 (N_5552,N_81,N_1659);
or U5553 (N_5553,N_2125,N_496);
or U5554 (N_5554,N_1883,N_887);
xnor U5555 (N_5555,N_188,N_1153);
xor U5556 (N_5556,N_578,N_2931);
or U5557 (N_5557,N_2162,N_2408);
xnor U5558 (N_5558,N_890,N_2815);
xor U5559 (N_5559,N_656,N_1258);
and U5560 (N_5560,N_2361,N_181);
nor U5561 (N_5561,N_2001,N_480);
and U5562 (N_5562,N_1045,N_481);
nor U5563 (N_5563,N_2253,N_351);
nor U5564 (N_5564,N_2584,N_16);
nor U5565 (N_5565,N_1927,N_108);
and U5566 (N_5566,N_2726,N_493);
nand U5567 (N_5567,N_2632,N_623);
and U5568 (N_5568,N_1379,N_1124);
and U5569 (N_5569,N_2771,N_412);
nand U5570 (N_5570,N_859,N_2760);
nand U5571 (N_5571,N_1285,N_279);
nand U5572 (N_5572,N_2975,N_2949);
nand U5573 (N_5573,N_583,N_643);
or U5574 (N_5574,N_2906,N_2903);
or U5575 (N_5575,N_124,N_2400);
nor U5576 (N_5576,N_2332,N_1540);
and U5577 (N_5577,N_1224,N_481);
and U5578 (N_5578,N_296,N_2527);
or U5579 (N_5579,N_418,N_2676);
xnor U5580 (N_5580,N_2372,N_2811);
and U5581 (N_5581,N_721,N_2230);
xnor U5582 (N_5582,N_1234,N_1365);
or U5583 (N_5583,N_1485,N_418);
xnor U5584 (N_5584,N_1533,N_2360);
xnor U5585 (N_5585,N_36,N_1727);
nand U5586 (N_5586,N_401,N_2787);
xnor U5587 (N_5587,N_1632,N_584);
nor U5588 (N_5588,N_1371,N_50);
nand U5589 (N_5589,N_2403,N_95);
nand U5590 (N_5590,N_1908,N_1370);
nand U5591 (N_5591,N_599,N_1603);
xor U5592 (N_5592,N_1998,N_1426);
nand U5593 (N_5593,N_2171,N_1603);
or U5594 (N_5594,N_2067,N_2242);
nand U5595 (N_5595,N_1746,N_613);
nor U5596 (N_5596,N_2925,N_1761);
nand U5597 (N_5597,N_425,N_1973);
nor U5598 (N_5598,N_2224,N_2809);
nand U5599 (N_5599,N_2562,N_1201);
or U5600 (N_5600,N_1261,N_1968);
nor U5601 (N_5601,N_2255,N_948);
or U5602 (N_5602,N_729,N_1233);
and U5603 (N_5603,N_2786,N_563);
or U5604 (N_5604,N_2537,N_2850);
nand U5605 (N_5605,N_2504,N_2506);
and U5606 (N_5606,N_2571,N_1759);
nand U5607 (N_5607,N_2857,N_2407);
nor U5608 (N_5608,N_653,N_2366);
and U5609 (N_5609,N_1189,N_1621);
or U5610 (N_5610,N_537,N_1614);
or U5611 (N_5611,N_1628,N_392);
xor U5612 (N_5612,N_15,N_2987);
or U5613 (N_5613,N_1843,N_1174);
nor U5614 (N_5614,N_2838,N_512);
or U5615 (N_5615,N_838,N_1912);
and U5616 (N_5616,N_841,N_2822);
nor U5617 (N_5617,N_1490,N_2068);
or U5618 (N_5618,N_258,N_2392);
xnor U5619 (N_5619,N_1321,N_941);
or U5620 (N_5620,N_1397,N_1972);
nor U5621 (N_5621,N_1988,N_2775);
xnor U5622 (N_5622,N_151,N_2100);
nand U5623 (N_5623,N_468,N_1990);
nand U5624 (N_5624,N_2036,N_2007);
or U5625 (N_5625,N_267,N_2200);
or U5626 (N_5626,N_150,N_1027);
nand U5627 (N_5627,N_2072,N_106);
and U5628 (N_5628,N_2710,N_1601);
and U5629 (N_5629,N_2143,N_1365);
and U5630 (N_5630,N_687,N_2650);
nand U5631 (N_5631,N_38,N_1882);
or U5632 (N_5632,N_2825,N_2395);
nand U5633 (N_5633,N_2075,N_1362);
nand U5634 (N_5634,N_2982,N_1214);
nor U5635 (N_5635,N_612,N_978);
and U5636 (N_5636,N_1220,N_1807);
or U5637 (N_5637,N_991,N_2635);
and U5638 (N_5638,N_1153,N_1463);
or U5639 (N_5639,N_342,N_2642);
and U5640 (N_5640,N_2501,N_64);
nand U5641 (N_5641,N_206,N_1324);
xor U5642 (N_5642,N_960,N_1076);
or U5643 (N_5643,N_797,N_560);
or U5644 (N_5644,N_2570,N_333);
xnor U5645 (N_5645,N_2256,N_1103);
and U5646 (N_5646,N_2962,N_1680);
and U5647 (N_5647,N_1240,N_211);
and U5648 (N_5648,N_2715,N_560);
or U5649 (N_5649,N_2025,N_104);
or U5650 (N_5650,N_1081,N_2661);
nor U5651 (N_5651,N_2711,N_1759);
xor U5652 (N_5652,N_384,N_2530);
nor U5653 (N_5653,N_2181,N_2044);
nand U5654 (N_5654,N_811,N_2432);
or U5655 (N_5655,N_2054,N_2355);
nor U5656 (N_5656,N_2925,N_703);
and U5657 (N_5657,N_1712,N_2357);
or U5658 (N_5658,N_262,N_1761);
and U5659 (N_5659,N_1069,N_2045);
and U5660 (N_5660,N_1748,N_1523);
nand U5661 (N_5661,N_1280,N_1272);
nor U5662 (N_5662,N_1848,N_332);
nor U5663 (N_5663,N_288,N_2190);
xnor U5664 (N_5664,N_1864,N_1682);
nor U5665 (N_5665,N_1833,N_1790);
or U5666 (N_5666,N_0,N_1102);
or U5667 (N_5667,N_2074,N_2464);
xnor U5668 (N_5668,N_909,N_2174);
and U5669 (N_5669,N_1523,N_1924);
nand U5670 (N_5670,N_1536,N_1704);
xor U5671 (N_5671,N_2859,N_1865);
xor U5672 (N_5672,N_2902,N_2461);
xnor U5673 (N_5673,N_2204,N_2949);
xnor U5674 (N_5674,N_1889,N_1111);
nand U5675 (N_5675,N_2219,N_2091);
xor U5676 (N_5676,N_241,N_964);
nor U5677 (N_5677,N_599,N_2814);
nor U5678 (N_5678,N_1054,N_2528);
or U5679 (N_5679,N_1923,N_1086);
nand U5680 (N_5680,N_1105,N_1764);
or U5681 (N_5681,N_2274,N_78);
nor U5682 (N_5682,N_296,N_1356);
xor U5683 (N_5683,N_1104,N_1796);
xor U5684 (N_5684,N_504,N_692);
nor U5685 (N_5685,N_4,N_822);
nand U5686 (N_5686,N_2226,N_738);
nor U5687 (N_5687,N_2281,N_2074);
xnor U5688 (N_5688,N_477,N_25);
nor U5689 (N_5689,N_2560,N_2760);
and U5690 (N_5690,N_2582,N_440);
and U5691 (N_5691,N_1396,N_926);
and U5692 (N_5692,N_594,N_2223);
nand U5693 (N_5693,N_2635,N_1146);
and U5694 (N_5694,N_948,N_483);
nor U5695 (N_5695,N_1310,N_294);
nor U5696 (N_5696,N_1572,N_522);
or U5697 (N_5697,N_1715,N_1296);
or U5698 (N_5698,N_2895,N_2883);
or U5699 (N_5699,N_545,N_2518);
xor U5700 (N_5700,N_600,N_1769);
or U5701 (N_5701,N_1210,N_2028);
and U5702 (N_5702,N_1493,N_1627);
or U5703 (N_5703,N_1411,N_2710);
nand U5704 (N_5704,N_856,N_933);
or U5705 (N_5705,N_2036,N_1835);
or U5706 (N_5706,N_207,N_1011);
nor U5707 (N_5707,N_703,N_2760);
or U5708 (N_5708,N_1858,N_2140);
xor U5709 (N_5709,N_2077,N_440);
or U5710 (N_5710,N_2175,N_1255);
xnor U5711 (N_5711,N_128,N_2180);
and U5712 (N_5712,N_747,N_1334);
nor U5713 (N_5713,N_658,N_2917);
nand U5714 (N_5714,N_1991,N_2479);
nor U5715 (N_5715,N_657,N_2258);
and U5716 (N_5716,N_2971,N_2882);
nand U5717 (N_5717,N_27,N_2197);
or U5718 (N_5718,N_1271,N_331);
nor U5719 (N_5719,N_2818,N_1414);
xnor U5720 (N_5720,N_2698,N_1592);
nor U5721 (N_5721,N_373,N_2353);
nor U5722 (N_5722,N_768,N_2853);
nand U5723 (N_5723,N_2531,N_2990);
xnor U5724 (N_5724,N_1594,N_1746);
xor U5725 (N_5725,N_1706,N_588);
or U5726 (N_5726,N_739,N_2873);
nand U5727 (N_5727,N_239,N_18);
and U5728 (N_5728,N_1674,N_410);
nor U5729 (N_5729,N_1012,N_1134);
xor U5730 (N_5730,N_539,N_818);
nand U5731 (N_5731,N_2350,N_792);
and U5732 (N_5732,N_1849,N_292);
nand U5733 (N_5733,N_2047,N_2076);
or U5734 (N_5734,N_1897,N_2918);
and U5735 (N_5735,N_1637,N_1418);
nor U5736 (N_5736,N_3,N_2445);
and U5737 (N_5737,N_1599,N_2342);
xnor U5738 (N_5738,N_2494,N_1105);
nand U5739 (N_5739,N_511,N_655);
nor U5740 (N_5740,N_1301,N_1265);
xor U5741 (N_5741,N_1053,N_1745);
nand U5742 (N_5742,N_1337,N_1036);
xor U5743 (N_5743,N_2288,N_304);
or U5744 (N_5744,N_1862,N_974);
nand U5745 (N_5745,N_811,N_1618);
nand U5746 (N_5746,N_453,N_2845);
nand U5747 (N_5747,N_2337,N_1988);
or U5748 (N_5748,N_1434,N_2839);
nor U5749 (N_5749,N_2409,N_1570);
or U5750 (N_5750,N_211,N_132);
or U5751 (N_5751,N_634,N_2499);
nor U5752 (N_5752,N_2604,N_2614);
or U5753 (N_5753,N_2329,N_1712);
and U5754 (N_5754,N_2847,N_2291);
or U5755 (N_5755,N_1411,N_1092);
and U5756 (N_5756,N_1331,N_2810);
and U5757 (N_5757,N_2148,N_773);
nor U5758 (N_5758,N_1919,N_1211);
or U5759 (N_5759,N_1745,N_1425);
and U5760 (N_5760,N_537,N_1139);
nor U5761 (N_5761,N_325,N_1845);
nand U5762 (N_5762,N_449,N_155);
and U5763 (N_5763,N_2547,N_2989);
or U5764 (N_5764,N_2238,N_356);
and U5765 (N_5765,N_1190,N_423);
and U5766 (N_5766,N_862,N_2306);
xor U5767 (N_5767,N_2826,N_2921);
xor U5768 (N_5768,N_1390,N_324);
and U5769 (N_5769,N_481,N_2891);
xor U5770 (N_5770,N_168,N_656);
nand U5771 (N_5771,N_2954,N_197);
nor U5772 (N_5772,N_1210,N_1242);
and U5773 (N_5773,N_2509,N_2627);
and U5774 (N_5774,N_518,N_2803);
xnor U5775 (N_5775,N_2636,N_2773);
xnor U5776 (N_5776,N_1338,N_966);
xnor U5777 (N_5777,N_345,N_252);
nor U5778 (N_5778,N_2114,N_416);
nor U5779 (N_5779,N_206,N_2305);
and U5780 (N_5780,N_363,N_2142);
nor U5781 (N_5781,N_2843,N_1942);
and U5782 (N_5782,N_758,N_340);
or U5783 (N_5783,N_222,N_1484);
nand U5784 (N_5784,N_2319,N_452);
xnor U5785 (N_5785,N_2879,N_213);
nor U5786 (N_5786,N_328,N_1310);
nand U5787 (N_5787,N_266,N_569);
nand U5788 (N_5788,N_201,N_24);
nand U5789 (N_5789,N_1975,N_1211);
xor U5790 (N_5790,N_1231,N_1780);
and U5791 (N_5791,N_902,N_178);
xor U5792 (N_5792,N_2166,N_2069);
xnor U5793 (N_5793,N_687,N_1804);
xnor U5794 (N_5794,N_1695,N_2545);
xor U5795 (N_5795,N_2817,N_2508);
nor U5796 (N_5796,N_1427,N_788);
nand U5797 (N_5797,N_2488,N_462);
nor U5798 (N_5798,N_1418,N_2443);
nor U5799 (N_5799,N_2218,N_1116);
nor U5800 (N_5800,N_347,N_2562);
or U5801 (N_5801,N_159,N_485);
or U5802 (N_5802,N_2704,N_2237);
nand U5803 (N_5803,N_1816,N_2726);
and U5804 (N_5804,N_499,N_536);
nand U5805 (N_5805,N_1585,N_2332);
and U5806 (N_5806,N_2626,N_2153);
xnor U5807 (N_5807,N_1024,N_1113);
xor U5808 (N_5808,N_1173,N_2817);
nor U5809 (N_5809,N_711,N_670);
nand U5810 (N_5810,N_1472,N_2846);
nand U5811 (N_5811,N_97,N_2294);
and U5812 (N_5812,N_247,N_897);
xor U5813 (N_5813,N_1682,N_2165);
and U5814 (N_5814,N_2471,N_2780);
xnor U5815 (N_5815,N_936,N_2301);
or U5816 (N_5816,N_2371,N_2441);
xor U5817 (N_5817,N_1738,N_834);
nor U5818 (N_5818,N_650,N_1781);
xor U5819 (N_5819,N_2043,N_2352);
and U5820 (N_5820,N_438,N_787);
xnor U5821 (N_5821,N_2575,N_97);
nor U5822 (N_5822,N_1137,N_1827);
and U5823 (N_5823,N_2185,N_802);
nor U5824 (N_5824,N_1277,N_2940);
nand U5825 (N_5825,N_1237,N_1189);
and U5826 (N_5826,N_1694,N_1222);
or U5827 (N_5827,N_2806,N_2942);
or U5828 (N_5828,N_640,N_1507);
xor U5829 (N_5829,N_2967,N_1671);
nor U5830 (N_5830,N_2539,N_928);
or U5831 (N_5831,N_1484,N_5);
nand U5832 (N_5832,N_1354,N_1629);
and U5833 (N_5833,N_408,N_1997);
nand U5834 (N_5834,N_134,N_1453);
or U5835 (N_5835,N_808,N_1954);
or U5836 (N_5836,N_1796,N_1114);
or U5837 (N_5837,N_332,N_531);
and U5838 (N_5838,N_2124,N_1359);
nand U5839 (N_5839,N_808,N_2766);
nor U5840 (N_5840,N_1897,N_1724);
xor U5841 (N_5841,N_1116,N_556);
nor U5842 (N_5842,N_1761,N_1036);
or U5843 (N_5843,N_2444,N_2601);
xnor U5844 (N_5844,N_1957,N_1255);
nor U5845 (N_5845,N_196,N_863);
nor U5846 (N_5846,N_72,N_349);
or U5847 (N_5847,N_2645,N_2354);
xor U5848 (N_5848,N_2231,N_1402);
and U5849 (N_5849,N_1784,N_1519);
nand U5850 (N_5850,N_540,N_0);
nand U5851 (N_5851,N_239,N_1376);
or U5852 (N_5852,N_1940,N_253);
and U5853 (N_5853,N_928,N_2589);
or U5854 (N_5854,N_2178,N_546);
nor U5855 (N_5855,N_16,N_372);
or U5856 (N_5856,N_1392,N_1523);
nand U5857 (N_5857,N_2784,N_175);
nor U5858 (N_5858,N_1993,N_989);
nor U5859 (N_5859,N_927,N_1591);
or U5860 (N_5860,N_1023,N_2675);
or U5861 (N_5861,N_1043,N_1787);
nand U5862 (N_5862,N_2547,N_1445);
nand U5863 (N_5863,N_102,N_2770);
or U5864 (N_5864,N_1619,N_1681);
or U5865 (N_5865,N_2074,N_2444);
or U5866 (N_5866,N_540,N_983);
xnor U5867 (N_5867,N_1349,N_567);
and U5868 (N_5868,N_2597,N_1201);
xor U5869 (N_5869,N_1041,N_2604);
and U5870 (N_5870,N_2919,N_2291);
or U5871 (N_5871,N_1405,N_2812);
xor U5872 (N_5872,N_1109,N_1645);
nand U5873 (N_5873,N_1236,N_784);
xnor U5874 (N_5874,N_1836,N_558);
nor U5875 (N_5875,N_2819,N_2082);
nor U5876 (N_5876,N_2869,N_521);
nor U5877 (N_5877,N_2989,N_2304);
nand U5878 (N_5878,N_456,N_1198);
and U5879 (N_5879,N_36,N_1921);
or U5880 (N_5880,N_1594,N_1015);
or U5881 (N_5881,N_2222,N_1366);
nand U5882 (N_5882,N_1091,N_465);
or U5883 (N_5883,N_1111,N_592);
nand U5884 (N_5884,N_1865,N_1220);
nand U5885 (N_5885,N_1035,N_1511);
or U5886 (N_5886,N_1970,N_2669);
nor U5887 (N_5887,N_453,N_118);
xor U5888 (N_5888,N_615,N_2775);
and U5889 (N_5889,N_1350,N_1291);
or U5890 (N_5890,N_441,N_1856);
xnor U5891 (N_5891,N_2497,N_2380);
nor U5892 (N_5892,N_1797,N_72);
or U5893 (N_5893,N_934,N_1867);
nand U5894 (N_5894,N_1327,N_2218);
and U5895 (N_5895,N_2448,N_2690);
nand U5896 (N_5896,N_2089,N_646);
or U5897 (N_5897,N_1084,N_1002);
xnor U5898 (N_5898,N_761,N_1213);
nand U5899 (N_5899,N_1414,N_446);
nor U5900 (N_5900,N_362,N_2516);
xnor U5901 (N_5901,N_108,N_642);
xor U5902 (N_5902,N_988,N_2973);
nand U5903 (N_5903,N_2102,N_1700);
nand U5904 (N_5904,N_1054,N_2904);
xnor U5905 (N_5905,N_1318,N_2820);
or U5906 (N_5906,N_2388,N_459);
or U5907 (N_5907,N_1384,N_656);
nand U5908 (N_5908,N_2747,N_1923);
or U5909 (N_5909,N_2250,N_979);
nand U5910 (N_5910,N_1049,N_275);
nor U5911 (N_5911,N_278,N_2472);
and U5912 (N_5912,N_570,N_2799);
nand U5913 (N_5913,N_1872,N_16);
nand U5914 (N_5914,N_2746,N_707);
and U5915 (N_5915,N_1548,N_1923);
or U5916 (N_5916,N_1521,N_2503);
nor U5917 (N_5917,N_2117,N_389);
or U5918 (N_5918,N_711,N_2206);
nor U5919 (N_5919,N_1183,N_2559);
xnor U5920 (N_5920,N_1126,N_709);
or U5921 (N_5921,N_2745,N_2325);
nand U5922 (N_5922,N_1197,N_164);
or U5923 (N_5923,N_145,N_1811);
or U5924 (N_5924,N_70,N_1836);
xnor U5925 (N_5925,N_1285,N_1564);
and U5926 (N_5926,N_2454,N_1705);
and U5927 (N_5927,N_603,N_2508);
or U5928 (N_5928,N_2311,N_274);
nand U5929 (N_5929,N_226,N_664);
nor U5930 (N_5930,N_2291,N_2262);
nand U5931 (N_5931,N_2437,N_295);
and U5932 (N_5932,N_1097,N_2930);
xnor U5933 (N_5933,N_2375,N_411);
nand U5934 (N_5934,N_1709,N_496);
and U5935 (N_5935,N_2156,N_2613);
and U5936 (N_5936,N_2198,N_2710);
xnor U5937 (N_5937,N_2503,N_1445);
xnor U5938 (N_5938,N_623,N_54);
and U5939 (N_5939,N_2661,N_1027);
and U5940 (N_5940,N_1932,N_237);
and U5941 (N_5941,N_1857,N_1347);
nand U5942 (N_5942,N_133,N_93);
xor U5943 (N_5943,N_2875,N_865);
and U5944 (N_5944,N_466,N_1234);
and U5945 (N_5945,N_663,N_2046);
or U5946 (N_5946,N_1950,N_165);
or U5947 (N_5947,N_187,N_2087);
or U5948 (N_5948,N_75,N_1039);
and U5949 (N_5949,N_952,N_2042);
and U5950 (N_5950,N_2510,N_1741);
or U5951 (N_5951,N_2052,N_2474);
and U5952 (N_5952,N_1434,N_694);
nor U5953 (N_5953,N_287,N_906);
and U5954 (N_5954,N_480,N_1646);
and U5955 (N_5955,N_111,N_2809);
nor U5956 (N_5956,N_2658,N_2729);
and U5957 (N_5957,N_905,N_2462);
xor U5958 (N_5958,N_575,N_28);
nor U5959 (N_5959,N_1122,N_2465);
nor U5960 (N_5960,N_960,N_1446);
nor U5961 (N_5961,N_2004,N_1376);
nand U5962 (N_5962,N_1881,N_902);
nand U5963 (N_5963,N_1706,N_2312);
nand U5964 (N_5964,N_1284,N_198);
nor U5965 (N_5965,N_23,N_2314);
nor U5966 (N_5966,N_1678,N_14);
and U5967 (N_5967,N_938,N_1295);
nor U5968 (N_5968,N_2578,N_2710);
nand U5969 (N_5969,N_408,N_536);
and U5970 (N_5970,N_838,N_1490);
and U5971 (N_5971,N_2570,N_1375);
nor U5972 (N_5972,N_1521,N_146);
and U5973 (N_5973,N_310,N_381);
nor U5974 (N_5974,N_1843,N_1690);
and U5975 (N_5975,N_2775,N_5);
nor U5976 (N_5976,N_1768,N_1577);
nand U5977 (N_5977,N_2680,N_2813);
or U5978 (N_5978,N_4,N_1256);
nand U5979 (N_5979,N_2529,N_1932);
xnor U5980 (N_5980,N_1706,N_2645);
xnor U5981 (N_5981,N_732,N_1854);
and U5982 (N_5982,N_989,N_2864);
nand U5983 (N_5983,N_1097,N_1640);
xor U5984 (N_5984,N_775,N_798);
nor U5985 (N_5985,N_902,N_1577);
or U5986 (N_5986,N_400,N_269);
nor U5987 (N_5987,N_824,N_2098);
or U5988 (N_5988,N_62,N_1709);
nor U5989 (N_5989,N_2582,N_2719);
nand U5990 (N_5990,N_1996,N_2292);
nor U5991 (N_5991,N_2190,N_851);
or U5992 (N_5992,N_1479,N_2307);
or U5993 (N_5993,N_2042,N_795);
nor U5994 (N_5994,N_2855,N_1447);
and U5995 (N_5995,N_960,N_431);
nand U5996 (N_5996,N_2539,N_298);
and U5997 (N_5997,N_1819,N_2507);
nand U5998 (N_5998,N_1707,N_2598);
nor U5999 (N_5999,N_12,N_546);
nand U6000 (N_6000,N_4860,N_5755);
or U6001 (N_6001,N_4080,N_5134);
nor U6002 (N_6002,N_3351,N_3792);
nor U6003 (N_6003,N_4527,N_5746);
or U6004 (N_6004,N_3610,N_4116);
nand U6005 (N_6005,N_3898,N_3735);
xnor U6006 (N_6006,N_4970,N_4456);
xnor U6007 (N_6007,N_4735,N_4337);
xor U6008 (N_6008,N_3818,N_4831);
xnor U6009 (N_6009,N_3376,N_4914);
and U6010 (N_6010,N_5520,N_3903);
nand U6011 (N_6011,N_4239,N_4324);
nand U6012 (N_6012,N_3862,N_4237);
or U6013 (N_6013,N_4119,N_5562);
nor U6014 (N_6014,N_3358,N_5944);
or U6015 (N_6015,N_4511,N_4316);
or U6016 (N_6016,N_4790,N_5108);
nor U6017 (N_6017,N_3773,N_5922);
and U6018 (N_6018,N_5574,N_3262);
xnor U6019 (N_6019,N_4624,N_4664);
xnor U6020 (N_6020,N_3266,N_4933);
nor U6021 (N_6021,N_5978,N_3033);
nand U6022 (N_6022,N_5006,N_3016);
nor U6023 (N_6023,N_4408,N_5340);
xnor U6024 (N_6024,N_5770,N_3528);
xor U6025 (N_6025,N_3323,N_3057);
and U6026 (N_6026,N_3018,N_3196);
and U6027 (N_6027,N_3024,N_4270);
or U6028 (N_6028,N_3430,N_5396);
xor U6029 (N_6029,N_3680,N_3447);
and U6030 (N_6030,N_4290,N_4996);
xor U6031 (N_6031,N_5205,N_4857);
nor U6032 (N_6032,N_4631,N_4365);
nand U6033 (N_6033,N_3642,N_3150);
xnor U6034 (N_6034,N_4490,N_5661);
or U6035 (N_6035,N_4530,N_4562);
or U6036 (N_6036,N_5934,N_4172);
nand U6037 (N_6037,N_5993,N_4120);
and U6038 (N_6038,N_3381,N_5336);
and U6039 (N_6039,N_3516,N_4249);
nor U6040 (N_6040,N_3488,N_3041);
or U6041 (N_6041,N_5100,N_4174);
xnor U6042 (N_6042,N_3989,N_3404);
xor U6043 (N_6043,N_4158,N_3184);
xor U6044 (N_6044,N_5779,N_3225);
nor U6045 (N_6045,N_5435,N_4342);
or U6046 (N_6046,N_5794,N_4386);
and U6047 (N_6047,N_5639,N_4060);
nor U6048 (N_6048,N_5596,N_4839);
nor U6049 (N_6049,N_4704,N_3585);
xor U6050 (N_6050,N_3367,N_4400);
nor U6051 (N_6051,N_5584,N_5069);
and U6052 (N_6052,N_3101,N_5615);
xnor U6053 (N_6053,N_3526,N_4668);
or U6054 (N_6054,N_3475,N_3620);
and U6055 (N_6055,N_5690,N_3461);
nand U6056 (N_6056,N_3649,N_3967);
nand U6057 (N_6057,N_4495,N_4039);
or U6058 (N_6058,N_4001,N_5912);
nor U6059 (N_6059,N_4332,N_4619);
or U6060 (N_6060,N_4247,N_4462);
nor U6061 (N_6061,N_5239,N_4707);
nor U6062 (N_6062,N_4100,N_4881);
and U6063 (N_6063,N_4723,N_5478);
xor U6064 (N_6064,N_5885,N_3491);
nand U6065 (N_6065,N_5333,N_4805);
and U6066 (N_6066,N_4508,N_4955);
nor U6067 (N_6067,N_5614,N_4561);
or U6068 (N_6068,N_3242,N_3696);
and U6069 (N_6069,N_5074,N_5876);
nor U6070 (N_6070,N_3863,N_5405);
or U6071 (N_6071,N_3343,N_4637);
or U6072 (N_6072,N_3256,N_5242);
and U6073 (N_6073,N_5228,N_5706);
and U6074 (N_6074,N_3954,N_5059);
nor U6075 (N_6075,N_4801,N_4146);
nor U6076 (N_6076,N_4677,N_3207);
or U6077 (N_6077,N_5730,N_5905);
nor U6078 (N_6078,N_3556,N_4278);
nor U6079 (N_6079,N_3678,N_3065);
or U6080 (N_6080,N_3513,N_5888);
and U6081 (N_6081,N_5994,N_5629);
or U6082 (N_6082,N_5650,N_4979);
nand U6083 (N_6083,N_5973,N_5692);
and U6084 (N_6084,N_5728,N_4096);
xor U6085 (N_6085,N_3036,N_5966);
nor U6086 (N_6086,N_5810,N_4416);
nand U6087 (N_6087,N_5747,N_3174);
nor U6088 (N_6088,N_4653,N_3825);
and U6089 (N_6089,N_3807,N_3572);
nand U6090 (N_6090,N_5272,N_4851);
or U6091 (N_6091,N_5687,N_3474);
or U6092 (N_6092,N_5426,N_3754);
xnor U6093 (N_6093,N_4563,N_4098);
xnor U6094 (N_6094,N_4433,N_4409);
nand U6095 (N_6095,N_5214,N_5185);
and U6096 (N_6096,N_3464,N_5036);
xor U6097 (N_6097,N_4727,N_3647);
or U6098 (N_6098,N_4049,N_5578);
nor U6099 (N_6099,N_4225,N_4545);
and U6100 (N_6100,N_4378,N_3548);
xnor U6101 (N_6101,N_5081,N_3719);
nand U6102 (N_6102,N_3438,N_5600);
nand U6103 (N_6103,N_3428,N_4868);
and U6104 (N_6104,N_5937,N_3922);
and U6105 (N_6105,N_5724,N_3440);
nand U6106 (N_6106,N_3766,N_4110);
and U6107 (N_6107,N_4605,N_3843);
nand U6108 (N_6108,N_3154,N_5399);
nand U6109 (N_6109,N_3177,N_4756);
xnor U6110 (N_6110,N_3896,N_5416);
nor U6111 (N_6111,N_5590,N_3763);
or U6112 (N_6112,N_5060,N_4683);
and U6113 (N_6113,N_4055,N_5750);
or U6114 (N_6114,N_3940,N_4772);
nor U6115 (N_6115,N_4929,N_4256);
nand U6116 (N_6116,N_4223,N_5822);
nor U6117 (N_6117,N_4101,N_3672);
xnor U6118 (N_6118,N_3597,N_3919);
or U6119 (N_6119,N_4730,N_5097);
nand U6120 (N_6120,N_4688,N_5261);
nand U6121 (N_6121,N_5855,N_4579);
nand U6122 (N_6122,N_3992,N_3145);
or U6123 (N_6123,N_3870,N_4635);
and U6124 (N_6124,N_4632,N_4824);
nand U6125 (N_6125,N_4414,N_5860);
or U6126 (N_6126,N_4732,N_3124);
nor U6127 (N_6127,N_4016,N_5575);
nor U6128 (N_6128,N_3176,N_5155);
nor U6129 (N_6129,N_4746,N_3129);
xnor U6130 (N_6130,N_3623,N_3293);
nor U6131 (N_6131,N_5249,N_3549);
xor U6132 (N_6132,N_5436,N_3013);
nor U6133 (N_6133,N_3340,N_5339);
nand U6134 (N_6134,N_4912,N_3749);
or U6135 (N_6135,N_3088,N_4775);
and U6136 (N_6136,N_3268,N_3525);
and U6137 (N_6137,N_3917,N_4476);
nor U6138 (N_6138,N_3045,N_4213);
nor U6139 (N_6139,N_4678,N_3155);
nor U6140 (N_6140,N_4984,N_5094);
nor U6141 (N_6141,N_5296,N_4082);
xnor U6142 (N_6142,N_5653,N_5041);
and U6143 (N_6143,N_4309,N_5087);
nand U6144 (N_6144,N_4760,N_4852);
or U6145 (N_6145,N_5714,N_5581);
and U6146 (N_6146,N_4622,N_3031);
nand U6147 (N_6147,N_4250,N_4969);
xor U6148 (N_6148,N_5982,N_3717);
or U6149 (N_6149,N_4892,N_3729);
xor U6150 (N_6150,N_4361,N_4965);
nor U6151 (N_6151,N_3830,N_5243);
nand U6152 (N_6152,N_5015,N_3644);
or U6153 (N_6153,N_4583,N_4672);
and U6154 (N_6154,N_5818,N_4017);
nor U6155 (N_6155,N_4949,N_4443);
and U6156 (N_6156,N_5259,N_3891);
xnor U6157 (N_6157,N_5902,N_5450);
nand U6158 (N_6158,N_4021,N_4124);
nand U6159 (N_6159,N_4064,N_4904);
or U6160 (N_6160,N_3973,N_5553);
or U6161 (N_6161,N_3675,N_3684);
xnor U6162 (N_6162,N_4516,N_3867);
xor U6163 (N_6163,N_3589,N_4159);
nor U6164 (N_6164,N_4370,N_5326);
nor U6165 (N_6165,N_5641,N_4321);
nand U6166 (N_6166,N_4499,N_4380);
nor U6167 (N_6167,N_3044,N_3755);
and U6168 (N_6168,N_4796,N_5114);
or U6169 (N_6169,N_5224,N_4422);
nor U6170 (N_6170,N_4828,N_4734);
nand U6171 (N_6171,N_4795,N_3083);
or U6172 (N_6172,N_5162,N_4600);
xnor U6173 (N_6173,N_4097,N_3732);
nor U6174 (N_6174,N_5572,N_4216);
or U6175 (N_6175,N_3550,N_3198);
and U6176 (N_6176,N_4510,N_4419);
nand U6177 (N_6177,N_5704,N_3402);
or U6178 (N_6178,N_4057,N_3598);
xor U6179 (N_6179,N_4701,N_4383);
nor U6180 (N_6180,N_5991,N_4126);
nand U6181 (N_6181,N_3512,N_5762);
nand U6182 (N_6182,N_4924,N_4178);
nand U6183 (N_6183,N_4133,N_5351);
or U6184 (N_6184,N_5234,N_3227);
nand U6185 (N_6185,N_4236,N_3361);
and U6186 (N_6186,N_5664,N_3181);
nor U6187 (N_6187,N_4451,N_4572);
nand U6188 (N_6188,N_5979,N_4663);
xor U6189 (N_6189,N_4267,N_5218);
or U6190 (N_6190,N_3591,N_5383);
nor U6191 (N_6191,N_4432,N_4791);
nor U6192 (N_6192,N_3694,N_5168);
xor U6193 (N_6193,N_3047,N_3864);
and U6194 (N_6194,N_5569,N_3422);
xor U6195 (N_6195,N_4586,N_5352);
xor U6196 (N_6196,N_3854,N_3350);
nor U6197 (N_6197,N_3325,N_3626);
and U6198 (N_6198,N_5680,N_3128);
xnor U6199 (N_6199,N_3582,N_4502);
or U6200 (N_6200,N_5962,N_5096);
or U6201 (N_6201,N_4343,N_3220);
or U6202 (N_6202,N_3835,N_3654);
xor U6203 (N_6203,N_5588,N_3179);
and U6204 (N_6204,N_5723,N_3799);
xor U6205 (N_6205,N_4072,N_4128);
nor U6206 (N_6206,N_4122,N_5131);
nor U6207 (N_6207,N_5460,N_5532);
nor U6208 (N_6208,N_5874,N_5184);
nor U6209 (N_6209,N_5579,N_4610);
nand U6210 (N_6210,N_3728,N_3393);
or U6211 (N_6211,N_4715,N_5656);
nor U6212 (N_6212,N_5718,N_5908);
and U6213 (N_6213,N_4621,N_3650);
nor U6214 (N_6214,N_5867,N_3206);
nand U6215 (N_6215,N_5945,N_3403);
nand U6216 (N_6216,N_5439,N_4388);
and U6217 (N_6217,N_5619,N_5480);
xor U6218 (N_6218,N_5211,N_5761);
or U6219 (N_6219,N_3514,N_3751);
nand U6220 (N_6220,N_3126,N_4713);
nor U6221 (N_6221,N_5857,N_3977);
nor U6222 (N_6222,N_4389,N_5288);
or U6223 (N_6223,N_3302,N_4402);
nand U6224 (N_6224,N_3506,N_5031);
nand U6225 (N_6225,N_3166,N_4764);
nor U6226 (N_6226,N_4165,N_5274);
nand U6227 (N_6227,N_5899,N_3079);
nor U6228 (N_6228,N_5491,N_3169);
xnor U6229 (N_6229,N_4463,N_4037);
and U6230 (N_6230,N_3700,N_5140);
xor U6231 (N_6231,N_3094,N_5645);
xnor U6232 (N_6232,N_4373,N_3733);
nor U6233 (N_6233,N_5144,N_5281);
and U6234 (N_6234,N_3312,N_4850);
and U6235 (N_6235,N_4837,N_3673);
and U6236 (N_6236,N_5148,N_3353);
or U6237 (N_6237,N_5726,N_5901);
nor U6238 (N_6238,N_4015,N_4010);
and U6239 (N_6239,N_3478,N_3373);
nand U6240 (N_6240,N_4488,N_4331);
or U6241 (N_6241,N_3743,N_3406);
and U6242 (N_6242,N_4272,N_3379);
nor U6243 (N_6243,N_4861,N_4887);
nand U6244 (N_6244,N_4345,N_5318);
or U6245 (N_6245,N_3153,N_3275);
xnor U6246 (N_6246,N_5915,N_3244);
nor U6247 (N_6247,N_4685,N_4196);
xor U6248 (N_6248,N_4131,N_5890);
xnor U6249 (N_6249,N_3286,N_3076);
nand U6250 (N_6250,N_3806,N_4595);
or U6251 (N_6251,N_4125,N_4604);
nand U6252 (N_6252,N_3490,N_5988);
and U6253 (N_6253,N_3541,N_4977);
and U6254 (N_6254,N_3905,N_3892);
xnor U6255 (N_6255,N_3923,N_4415);
xnor U6256 (N_6256,N_3061,N_5943);
or U6257 (N_6257,N_5796,N_3934);
nand U6258 (N_6258,N_5987,N_4152);
nand U6259 (N_6259,N_3183,N_3303);
and U6260 (N_6260,N_5275,N_3502);
and U6261 (N_6261,N_3646,N_3075);
xor U6262 (N_6262,N_3398,N_5844);
nor U6263 (N_6263,N_3131,N_5585);
xnor U6264 (N_6264,N_4574,N_4944);
xor U6265 (N_6265,N_3715,N_5063);
or U6266 (N_6266,N_3054,N_3636);
xor U6267 (N_6267,N_3364,N_4556);
nand U6268 (N_6268,N_5422,N_4564);
and U6269 (N_6269,N_3148,N_3968);
xor U6270 (N_6270,N_4325,N_3747);
and U6271 (N_6271,N_3296,N_4493);
xor U6272 (N_6272,N_4738,N_5486);
or U6273 (N_6273,N_5538,N_5132);
nand U6274 (N_6274,N_4173,N_5229);
or U6275 (N_6275,N_4243,N_4763);
and U6276 (N_6276,N_4496,N_5284);
or U6277 (N_6277,N_4138,N_4395);
nand U6278 (N_6278,N_4136,N_5699);
xor U6279 (N_6279,N_5289,N_4749);
nor U6280 (N_6280,N_5760,N_5252);
nand U6281 (N_6281,N_5010,N_3449);
or U6282 (N_6282,N_3042,N_5180);
nand U6283 (N_6283,N_3856,N_5283);
or U6284 (N_6284,N_5149,N_5671);
xor U6285 (N_6285,N_4694,N_5411);
or U6286 (N_6286,N_5567,N_5642);
nor U6287 (N_6287,N_4156,N_3055);
and U6288 (N_6288,N_4578,N_3942);
xor U6289 (N_6289,N_4457,N_4210);
xnor U6290 (N_6290,N_5171,N_3264);
nand U6291 (N_6291,N_4265,N_5996);
or U6292 (N_6292,N_3705,N_5636);
nor U6293 (N_6293,N_3910,N_3938);
nand U6294 (N_6294,N_4088,N_5102);
or U6295 (N_6295,N_3685,N_3710);
nor U6296 (N_6296,N_3049,N_4822);
nor U6297 (N_6297,N_4848,N_4872);
xnor U6298 (N_6298,N_5152,N_5291);
nor U6299 (N_6299,N_5852,N_5095);
and U6300 (N_6300,N_3238,N_5278);
or U6301 (N_6301,N_5861,N_3877);
xnor U6302 (N_6302,N_4051,N_4222);
or U6303 (N_6303,N_4960,N_5128);
nand U6304 (N_6304,N_3232,N_5332);
nand U6305 (N_6305,N_4534,N_4903);
or U6306 (N_6306,N_5540,N_4020);
nor U6307 (N_6307,N_5547,N_5964);
and U6308 (N_6308,N_5388,N_3161);
or U6309 (N_6309,N_3342,N_4834);
nor U6310 (N_6310,N_4441,N_4742);
and U6311 (N_6311,N_3897,N_4407);
and U6312 (N_6312,N_4477,N_4973);
or U6313 (N_6313,N_5508,N_3889);
or U6314 (N_6314,N_3921,N_4033);
nor U6315 (N_6315,N_4844,N_5147);
xor U6316 (N_6316,N_3439,N_4728);
nor U6317 (N_6317,N_5217,N_3215);
and U6318 (N_6318,N_5008,N_4843);
and U6319 (N_6319,N_4575,N_3297);
nand U6320 (N_6320,N_5795,N_4665);
nand U6321 (N_6321,N_4468,N_4818);
nor U6322 (N_6322,N_4648,N_5143);
xor U6323 (N_6323,N_5929,N_4004);
or U6324 (N_6324,N_4202,N_4470);
and U6325 (N_6325,N_3035,N_3239);
nand U6326 (N_6326,N_4226,N_4838);
and U6327 (N_6327,N_4177,N_5971);
and U6328 (N_6328,N_3282,N_5630);
and U6329 (N_6329,N_3831,N_3643);
nand U6330 (N_6330,N_4864,N_5196);
or U6331 (N_6331,N_3738,N_5892);
xnor U6332 (N_6332,N_3767,N_4030);
or U6333 (N_6333,N_3368,N_4987);
nor U6334 (N_6334,N_5904,N_5782);
or U6335 (N_6335,N_3105,N_4875);
and U6336 (N_6336,N_4306,N_5362);
nand U6337 (N_6337,N_3151,N_5141);
and U6338 (N_6338,N_4642,N_5787);
nor U6339 (N_6339,N_3466,N_5887);
nand U6340 (N_6340,N_4691,N_3857);
xnor U6341 (N_6341,N_3087,N_5829);
nor U6342 (N_6342,N_4608,N_5846);
nor U6343 (N_6343,N_5990,N_5722);
or U6344 (N_6344,N_4209,N_4918);
nand U6345 (N_6345,N_5047,N_4207);
nand U6346 (N_6346,N_4334,N_4961);
and U6347 (N_6347,N_4859,N_4964);
nor U6348 (N_6348,N_4641,N_3002);
or U6349 (N_6349,N_5900,N_3140);
xor U6350 (N_6350,N_5624,N_5398);
or U6351 (N_6351,N_3639,N_4939);
and U6352 (N_6352,N_3691,N_3943);
and U6353 (N_6353,N_5024,N_3969);
and U6354 (N_6354,N_5977,N_4821);
nand U6355 (N_6355,N_4638,N_5517);
nor U6356 (N_6356,N_5448,N_4279);
nand U6357 (N_6357,N_4139,N_3682);
or U6358 (N_6358,N_5297,N_5920);
and U6359 (N_6359,N_3362,N_4926);
nand U6360 (N_6360,N_3027,N_5000);
and U6361 (N_6361,N_3432,N_4271);
xnor U6362 (N_6362,N_3566,N_4498);
and U6363 (N_6363,N_3359,N_3911);
nand U6364 (N_6364,N_4971,N_3454);
xnor U6365 (N_6365,N_3378,N_3100);
nor U6366 (N_6366,N_5186,N_4931);
or U6367 (N_6367,N_3819,N_4520);
xnor U6368 (N_6368,N_5985,N_3927);
and U6369 (N_6369,N_5367,N_4454);
xor U6370 (N_6370,N_5560,N_4189);
and U6371 (N_6371,N_3690,N_5542);
xnor U6372 (N_6372,N_5374,N_3498);
xor U6373 (N_6373,N_4467,N_5007);
or U6374 (N_6374,N_4000,N_3741);
and U6375 (N_6375,N_4639,N_5194);
xor U6376 (N_6376,N_4291,N_3666);
nand U6377 (N_6377,N_5053,N_3987);
nand U6378 (N_6378,N_3926,N_4765);
nor U6379 (N_6379,N_4863,N_5043);
and U6380 (N_6380,N_5707,N_4771);
nor U6381 (N_6381,N_4366,N_5372);
nor U6382 (N_6382,N_5471,N_5223);
nand U6383 (N_6383,N_5247,N_5678);
xnor U6384 (N_6384,N_5682,N_3584);
or U6385 (N_6385,N_3462,N_5836);
or U6386 (N_6386,N_4132,N_3060);
and U6387 (N_6387,N_5798,N_4895);
and U6388 (N_6388,N_3245,N_3269);
nand U6389 (N_6389,N_4698,N_5365);
nor U6390 (N_6390,N_3193,N_4399);
xor U6391 (N_6391,N_4761,N_5368);
or U6392 (N_6392,N_5535,N_4479);
nand U6393 (N_6393,N_4420,N_5044);
nand U6394 (N_6394,N_5566,N_3292);
xnor U6395 (N_6395,N_3431,N_4482);
nand U6396 (N_6396,N_4492,N_3985);
xor U6397 (N_6397,N_3394,N_3133);
nor U6398 (N_6398,N_4460,N_3117);
or U6399 (N_6399,N_5705,N_4450);
and U6400 (N_6400,N_5174,N_5745);
and U6401 (N_6401,N_4783,N_4606);
or U6402 (N_6402,N_3413,N_5627);
and U6403 (N_6403,N_3291,N_3116);
nand U6404 (N_6404,N_5648,N_5703);
or U6405 (N_6405,N_4846,N_3609);
and U6406 (N_6406,N_3504,N_4745);
or U6407 (N_6407,N_4046,N_4336);
and U6408 (N_6408,N_3663,N_5769);
nor U6409 (N_6409,N_5764,N_4878);
and U6410 (N_6410,N_3546,N_3383);
nand U6411 (N_6411,N_3357,N_3723);
or U6412 (N_6412,N_3909,N_4073);
nand U6413 (N_6413,N_5456,N_4221);
or U6414 (N_6414,N_5522,N_5033);
xnor U6415 (N_6415,N_3507,N_4932);
nand U6416 (N_6416,N_5913,N_4814);
nand U6417 (N_6417,N_4779,N_5858);
nor U6418 (N_6418,N_4351,N_3958);
and U6419 (N_6419,N_5129,N_3382);
xnor U6420 (N_6420,N_4589,N_3789);
xnor U6421 (N_6421,N_4503,N_5441);
xor U6422 (N_6422,N_4473,N_4014);
and U6423 (N_6423,N_4435,N_5752);
nand U6424 (N_6424,N_3883,N_3633);
nor U6425 (N_6425,N_3495,N_5206);
xnor U6426 (N_6426,N_3536,N_3544);
xor U6427 (N_6427,N_3095,N_5485);
xnor U6428 (N_6428,N_5733,N_5158);
nor U6429 (N_6429,N_4031,N_4829);
nor U6430 (N_6430,N_3852,N_5067);
or U6431 (N_6431,N_5638,N_4118);
and U6432 (N_6432,N_5894,N_4948);
xnor U6433 (N_6433,N_5428,N_5591);
and U6434 (N_6434,N_5772,N_5077);
and U6435 (N_6435,N_3539,N_3509);
or U6436 (N_6436,N_5086,N_4023);
nand U6437 (N_6437,N_3668,N_5935);
and U6438 (N_6438,N_4153,N_3731);
and U6439 (N_6439,N_4353,N_4986);
xor U6440 (N_6440,N_5354,N_5222);
or U6441 (N_6441,N_5269,N_3697);
and U6442 (N_6442,N_3604,N_4296);
nor U6443 (N_6443,N_5257,N_5369);
and U6444 (N_6444,N_4776,N_5871);
nor U6445 (N_6445,N_5446,N_4712);
and U6446 (N_6446,N_4594,N_4774);
nand U6447 (N_6447,N_4806,N_4930);
and U6448 (N_6448,N_3756,N_3552);
xor U6449 (N_6449,N_4991,N_3190);
or U6450 (N_6450,N_5974,N_4349);
nor U6451 (N_6451,N_5090,N_5421);
xnor U6452 (N_6452,N_5919,N_5592);
nand U6453 (N_6453,N_3981,N_3028);
and U6454 (N_6454,N_4780,N_4338);
nand U6455 (N_6455,N_5482,N_4203);
xor U6456 (N_6456,N_3706,N_3841);
xor U6457 (N_6457,N_4359,N_4328);
and U6458 (N_6458,N_4645,N_5493);
and U6459 (N_6459,N_4792,N_3267);
nor U6460 (N_6460,N_5835,N_3826);
or U6461 (N_6461,N_5343,N_4440);
and U6462 (N_6462,N_3662,N_4257);
xnor U6463 (N_6463,N_3932,N_5071);
xor U6464 (N_6464,N_3019,N_5187);
nor U6465 (N_6465,N_4640,N_4882);
xnor U6466 (N_6466,N_3764,N_3064);
or U6467 (N_6467,N_5092,N_5055);
or U6468 (N_6468,N_3071,N_5774);
xor U6469 (N_6469,N_5536,N_5942);
nor U6470 (N_6470,N_5049,N_5666);
nor U6471 (N_6471,N_5866,N_5341);
or U6472 (N_6472,N_3152,N_4559);
and U6473 (N_6473,N_3580,N_5777);
or U6474 (N_6474,N_4231,N_3614);
nor U6475 (N_6475,N_3974,N_4945);
nor U6476 (N_6476,N_4248,N_3470);
nor U6477 (N_6477,N_4319,N_4438);
nor U6478 (N_6478,N_5972,N_5568);
nor U6479 (N_6479,N_5376,N_5231);
nand U6480 (N_6480,N_3226,N_3070);
or U6481 (N_6481,N_4938,N_4849);
nand U6482 (N_6482,N_4167,N_3011);
xor U6483 (N_6483,N_3562,N_4008);
or U6484 (N_6484,N_3217,N_4013);
and U6485 (N_6485,N_5713,N_4856);
nand U6486 (N_6486,N_4940,N_3624);
and U6487 (N_6487,N_4092,N_5440);
nand U6488 (N_6488,N_5295,N_5506);
xnor U6489 (N_6489,N_4617,N_5999);
xnor U6490 (N_6490,N_4628,N_3659);
or U6491 (N_6491,N_4487,N_5394);
nand U6492 (N_6492,N_4323,N_5812);
xor U6493 (N_6493,N_3059,N_3429);
or U6494 (N_6494,N_5315,N_5612);
xnor U6495 (N_6495,N_3540,N_5895);
nand U6496 (N_6496,N_5729,N_5181);
or U6497 (N_6497,N_3319,N_4983);
and U6498 (N_6498,N_3698,N_3622);
nand U6499 (N_6499,N_4269,N_5375);
nor U6500 (N_6500,N_4782,N_5119);
and U6501 (N_6501,N_3842,N_4777);
xnor U6502 (N_6502,N_4618,N_4817);
and U6503 (N_6503,N_4826,N_4669);
nor U6504 (N_6504,N_3778,N_4254);
xnor U6505 (N_6505,N_3976,N_3637);
nand U6506 (N_6506,N_3115,N_5410);
and U6507 (N_6507,N_5361,N_5731);
and U6508 (N_6508,N_3410,N_5101);
nand U6509 (N_6509,N_5453,N_3468);
nor U6510 (N_6510,N_4150,N_3999);
nor U6511 (N_6511,N_4293,N_5427);
nand U6512 (N_6512,N_3336,N_3660);
and U6513 (N_6513,N_3522,N_5534);
nand U6514 (N_6514,N_5019,N_4382);
nand U6515 (N_6515,N_4117,N_4211);
and U6516 (N_6516,N_4748,N_5954);
xor U6517 (N_6517,N_5470,N_3017);
and U6518 (N_6518,N_5521,N_5558);
or U6519 (N_6519,N_5120,N_3021);
nor U6520 (N_6520,N_3072,N_3501);
nor U6521 (N_6521,N_4217,N_4307);
or U6522 (N_6522,N_4992,N_3270);
nand U6523 (N_6523,N_5415,N_4842);
nor U6524 (N_6524,N_5488,N_4106);
nor U6525 (N_6525,N_5788,N_3858);
xor U6526 (N_6526,N_5622,N_3186);
and U6527 (N_6527,N_4999,N_3228);
nand U6528 (N_6528,N_3619,N_4890);
nor U6529 (N_6529,N_4246,N_5387);
nand U6530 (N_6530,N_5827,N_3103);
or U6531 (N_6531,N_5580,N_4840);
xnor U6532 (N_6532,N_3670,N_4870);
xnor U6533 (N_6533,N_3010,N_4959);
or U6534 (N_6534,N_5492,N_4729);
nand U6535 (N_6535,N_5940,N_3524);
nand U6536 (N_6536,N_4358,N_3878);
or U6537 (N_6537,N_3020,N_3775);
or U6538 (N_6538,N_5864,N_5749);
or U6539 (N_6539,N_3607,N_3314);
or U6540 (N_6540,N_3545,N_5317);
xnor U6541 (N_6541,N_3156,N_3313);
or U6542 (N_6542,N_3606,N_3953);
or U6543 (N_6543,N_3203,N_4350);
or U6544 (N_6544,N_5595,N_4967);
and U6545 (N_6545,N_3446,N_3801);
nand U6546 (N_6546,N_4115,N_3485);
xnor U6547 (N_6547,N_5476,N_5337);
nand U6548 (N_6548,N_3593,N_4411);
nand U6549 (N_6549,N_4963,N_3727);
nor U6550 (N_6550,N_5625,N_4869);
xnor U6551 (N_6551,N_4535,N_3865);
nor U6552 (N_6552,N_3081,N_5740);
nor U6553 (N_6553,N_4154,N_4034);
and U6554 (N_6554,N_3257,N_4330);
nand U6555 (N_6555,N_3434,N_4050);
nand U6556 (N_6556,N_5301,N_4445);
nor U6557 (N_6557,N_3982,N_5497);
nand U6558 (N_6558,N_4005,N_4687);
and U6559 (N_6559,N_5273,N_5075);
nand U6560 (N_6560,N_5710,N_4725);
nand U6561 (N_6561,N_5425,N_3925);
and U6562 (N_6562,N_3386,N_3814);
or U6563 (N_6563,N_4372,N_5550);
nor U6564 (N_6564,N_3596,N_5013);
nor U6565 (N_6565,N_5197,N_4078);
nand U6566 (N_6566,N_3978,N_4925);
nand U6567 (N_6567,N_4998,N_4798);
and U6568 (N_6568,N_4867,N_5841);
xor U6569 (N_6569,N_5548,N_5490);
nor U6570 (N_6570,N_5349,N_5300);
xnor U6571 (N_6571,N_3739,N_5565);
nand U6572 (N_6572,N_3971,N_3347);
and U6573 (N_6573,N_5702,N_3995);
or U6574 (N_6574,N_4888,N_5685);
nand U6575 (N_6575,N_5821,N_4634);
or U6576 (N_6576,N_3770,N_5909);
nor U6577 (N_6577,N_4144,N_3613);
nand U6578 (N_6578,N_3782,N_5359);
nand U6579 (N_6579,N_5576,N_5549);
nand U6580 (N_6580,N_5121,N_5330);
or U6581 (N_6581,N_5392,N_5381);
and U6582 (N_6582,N_3533,N_3929);
xnor U6583 (N_6583,N_4737,N_4523);
and U6584 (N_6584,N_5552,N_4819);
and U6585 (N_6585,N_5452,N_5775);
xnor U6586 (N_6586,N_5851,N_3318);
and U6587 (N_6587,N_4612,N_4434);
nor U6588 (N_6588,N_5279,N_3794);
xor U6589 (N_6589,N_5122,N_4282);
or U6590 (N_6590,N_5430,N_3581);
xnor U6591 (N_6591,N_4418,N_5236);
or U6592 (N_6592,N_4149,N_3332);
nor U6593 (N_6593,N_3214,N_3221);
and U6594 (N_6594,N_4298,N_4753);
nor U6595 (N_6595,N_5854,N_4646);
nor U6596 (N_6596,N_5417,N_5378);
nor U6597 (N_6597,N_3165,N_5204);
nor U6598 (N_6598,N_3497,N_5382);
nor U6599 (N_6599,N_4067,N_5955);
and U6600 (N_6600,N_3702,N_4058);
nor U6601 (N_6601,N_3740,N_4083);
xnor U6602 (N_6602,N_4767,N_5696);
xor U6603 (N_6603,N_5800,N_4935);
and U6604 (N_6604,N_5235,N_5192);
xor U6605 (N_6605,N_4206,N_4810);
xnor U6606 (N_6606,N_4695,N_4980);
xor U6607 (N_6607,N_4876,N_5878);
xor U6608 (N_6608,N_4424,N_5429);
nand U6609 (N_6609,N_5838,N_5161);
and U6610 (N_6610,N_4405,N_5513);
xnor U6611 (N_6611,N_5462,N_4542);
and U6612 (N_6612,N_3679,N_5255);
or U6613 (N_6613,N_5136,N_3170);
xor U6614 (N_6614,N_5040,N_3811);
xor U6615 (N_6615,N_3241,N_3588);
nor U6616 (N_6616,N_4755,N_5757);
nand U6617 (N_6617,N_3025,N_5564);
xor U6618 (N_6618,N_4430,N_4662);
nor U6619 (N_6619,N_5632,N_3143);
xnor U6620 (N_6620,N_4344,N_4244);
and U6621 (N_6621,N_3029,N_4059);
nand U6622 (N_6622,N_4909,N_5366);
or U6623 (N_6623,N_3759,N_3960);
nor U6624 (N_6624,N_4448,N_4891);
and U6625 (N_6625,N_4543,N_4652);
nor U6626 (N_6626,N_3601,N_5676);
xor U6627 (N_6627,N_4941,N_4459);
nand U6628 (N_6628,N_4045,N_4346);
nor U6629 (N_6629,N_5062,N_4532);
or U6630 (N_6630,N_3832,N_4507);
xor U6631 (N_6631,N_3425,N_4573);
or U6632 (N_6632,N_5298,N_5842);
nor U6633 (N_6633,N_5969,N_4094);
nor U6634 (N_6634,N_5693,N_4649);
or U6635 (N_6635,N_3308,N_3994);
xnor U6636 (N_6636,N_5495,N_5172);
nand U6637 (N_6637,N_5391,N_3676);
nand U6638 (N_6638,N_4109,N_4786);
nand U6639 (N_6639,N_3372,N_5294);
nand U6640 (N_6640,N_3707,N_5865);
nor U6641 (N_6641,N_5780,N_3600);
nand U6642 (N_6642,N_5556,N_5084);
xnor U6643 (N_6643,N_3677,N_3850);
and U6644 (N_6644,N_5626,N_3201);
xnor U6645 (N_6645,N_4513,N_4916);
nand U6646 (N_6646,N_3908,N_3134);
nor U6647 (N_6647,N_5124,N_3421);
and U6648 (N_6648,N_4018,N_5052);
and U6649 (N_6649,N_4899,N_5959);
or U6650 (N_6650,N_3655,N_5673);
nor U6651 (N_6651,N_4897,N_5371);
nand U6652 (N_6652,N_3335,N_4708);
nor U6653 (N_6653,N_3876,N_5503);
xor U6654 (N_6654,N_5163,N_3630);
nand U6655 (N_6655,N_3753,N_5258);
and U6656 (N_6656,N_5334,N_5948);
nor U6657 (N_6657,N_4135,N_4766);
xnor U6658 (N_6658,N_3762,N_3483);
or U6659 (N_6659,N_3997,N_3538);
nand U6660 (N_6660,N_4908,N_5489);
or U6661 (N_6661,N_3602,N_3167);
nand U6662 (N_6662,N_3052,N_3839);
nor U6663 (N_6663,N_5789,N_5925);
nand U6664 (N_6664,N_3693,N_3627);
nor U6665 (N_6665,N_4990,N_3369);
nor U6666 (N_6666,N_4262,N_5323);
xnor U6667 (N_6667,N_5847,N_3936);
nand U6668 (N_6668,N_5066,N_5897);
or U6669 (N_6669,N_5928,N_3542);
or U6670 (N_6670,N_4880,N_3231);
nand U6671 (N_6671,N_4143,N_3748);
xor U6672 (N_6672,N_3744,N_5736);
xor U6673 (N_6673,N_4855,N_3515);
nor U6674 (N_6674,N_3399,N_5312);
and U6675 (N_6675,N_4182,N_3683);
or U6676 (N_6676,N_3531,N_5924);
nor U6677 (N_6677,N_5950,N_5353);
and U6678 (N_6678,N_4682,N_5302);
nor U6679 (N_6679,N_3034,N_3777);
and U6680 (N_6680,N_5939,N_4312);
and U6681 (N_6681,N_5791,N_5068);
and U6682 (N_6682,N_3686,N_3127);
nor U6683 (N_6683,N_4026,N_3638);
or U6684 (N_6684,N_5225,N_3416);
nand U6685 (N_6685,N_3420,N_4157);
nand U6686 (N_6686,N_4536,N_4596);
and U6687 (N_6687,N_3881,N_5561);
and U6688 (N_6688,N_5472,N_4962);
xnor U6689 (N_6689,N_5743,N_5716);
xnor U6690 (N_6690,N_5621,N_5266);
or U6691 (N_6691,N_4773,N_3586);
and U6692 (N_6692,N_5968,N_3924);
nor U6693 (N_6693,N_3003,N_3555);
or U6694 (N_6694,N_3671,N_3494);
nand U6695 (N_6695,N_5633,N_5831);
or U6696 (N_6696,N_4529,N_3000);
nand U6697 (N_6697,N_4541,N_4233);
nor U6698 (N_6698,N_5709,N_5306);
or U6699 (N_6699,N_5458,N_5355);
and U6700 (N_6700,N_4514,N_5833);
and U6701 (N_6701,N_4068,N_4229);
and U6702 (N_6702,N_5952,N_5451);
nand U6703 (N_6703,N_3913,N_5483);
xnor U6704 (N_6704,N_3860,N_5357);
or U6705 (N_6705,N_4198,N_4989);
nand U6706 (N_6706,N_3725,N_3499);
and U6707 (N_6707,N_4787,N_3511);
nor U6708 (N_6708,N_3793,N_5759);
and U6709 (N_6709,N_4928,N_5646);
nand U6710 (N_6710,N_3467,N_5358);
and U6711 (N_6711,N_5921,N_3817);
or U6712 (N_6712,N_4341,N_5014);
nand U6713 (N_6713,N_4758,N_3781);
nor U6714 (N_6714,N_3530,N_4444);
and U6715 (N_6715,N_5717,N_5042);
nor U6716 (N_6716,N_3861,N_3959);
nor U6717 (N_6717,N_5287,N_5203);
nor U6718 (N_6718,N_4284,N_3209);
nor U6719 (N_6719,N_3916,N_5324);
nor U6720 (N_6720,N_3893,N_5190);
xnor U6721 (N_6721,N_5079,N_4788);
xnor U6722 (N_6722,N_5021,N_3409);
xor U6723 (N_6723,N_3278,N_4762);
xor U6724 (N_6724,N_5896,N_5285);
and U6725 (N_6725,N_5884,N_5834);
and U6726 (N_6726,N_5758,N_4484);
xor U6727 (N_6727,N_4784,N_5173);
nand U6728 (N_6728,N_5674,N_4027);
and U6729 (N_6729,N_3774,N_3261);
nand U6730 (N_6730,N_5734,N_5363);
and U6731 (N_6731,N_4164,N_3653);
nor U6732 (N_6732,N_3254,N_4601);
nand U6733 (N_6733,N_3053,N_4988);
xnor U6734 (N_6734,N_4736,N_3112);
and U6735 (N_6735,N_3834,N_5213);
or U6736 (N_6736,N_5320,N_5658);
nand U6737 (N_6737,N_4593,N_4577);
or U6738 (N_6738,N_3272,N_5989);
nor U6739 (N_6739,N_4614,N_3713);
xnor U6740 (N_6740,N_3093,N_5668);
xnor U6741 (N_6741,N_3742,N_4486);
and U6742 (N_6742,N_5751,N_3592);
xor U6743 (N_6743,N_5193,N_3823);
or U6744 (N_6744,N_4019,N_4326);
nor U6745 (N_6745,N_3708,N_5479);
xor U6746 (N_6746,N_5819,N_5617);
nor U6747 (N_6747,N_3236,N_5931);
nor U6748 (N_6748,N_4393,N_3720);
and U6749 (N_6749,N_3941,N_4620);
or U6750 (N_6750,N_5377,N_3415);
nor U6751 (N_6751,N_4123,N_4981);
nor U6752 (N_6752,N_4160,N_5776);
nand U6753 (N_6753,N_4582,N_5742);
or U6754 (N_6754,N_4809,N_5524);
xnor U6755 (N_6755,N_3258,N_3354);
or U6756 (N_6756,N_5350,N_4397);
xor U6757 (N_6757,N_3391,N_4656);
or U6758 (N_6758,N_3077,N_4214);
nor U6759 (N_6759,N_4580,N_4232);
or U6760 (N_6760,N_5293,N_4464);
nor U6761 (N_6761,N_4515,N_3004);
nor U6762 (N_6762,N_5431,N_5364);
and U6763 (N_6763,N_4570,N_5806);
or U6764 (N_6764,N_5754,N_3437);
nor U6765 (N_6765,N_5393,N_4497);
or U6766 (N_6766,N_5442,N_5270);
and U6767 (N_6767,N_4105,N_4485);
nor U6768 (N_6768,N_3634,N_3991);
nand U6769 (N_6769,N_5175,N_5065);
and U6770 (N_6770,N_3274,N_3779);
nand U6771 (N_6771,N_3901,N_4011);
and U6772 (N_6772,N_4584,N_5432);
nand U6773 (N_6773,N_5058,N_3880);
xnor U6774 (N_6774,N_3508,N_5862);
nand U6775 (N_6775,N_3988,N_5933);
nand U6776 (N_6776,N_4613,N_4035);
and U6777 (N_6777,N_3543,N_4429);
and U6778 (N_6778,N_4069,N_4455);
nand U6779 (N_6779,N_3521,N_3699);
nand U6780 (N_6780,N_5863,N_4275);
nor U6781 (N_6781,N_3937,N_4107);
nand U6782 (N_6782,N_5157,N_3812);
xor U6783 (N_6783,N_5571,N_5299);
xnor U6784 (N_6784,N_3567,N_5557);
nand U6785 (N_6785,N_4854,N_4794);
or U6786 (N_6786,N_4320,N_3370);
xor U6787 (N_6787,N_5182,N_3455);
xor U6788 (N_6788,N_4335,N_5028);
nand U6789 (N_6789,N_3822,N_4410);
xor U6790 (N_6790,N_5941,N_5872);
and U6791 (N_6791,N_5914,N_4340);
or U6792 (N_6792,N_3078,N_3836);
or U6793 (N_6793,N_4830,N_4504);
xnor U6794 (N_6794,N_3529,N_3104);
nor U6795 (N_6795,N_5467,N_4716);
xor U6796 (N_6796,N_4228,N_5953);
xnor U6797 (N_6797,N_3249,N_4975);
nand U6798 (N_6798,N_5251,N_4720);
xnor U6799 (N_6799,N_4951,N_4483);
xnor U6800 (N_6800,N_3477,N_3972);
nor U6801 (N_6801,N_3787,N_3097);
or U6802 (N_6802,N_4188,N_5765);
and U6803 (N_6803,N_4710,N_5531);
nand U6804 (N_6804,N_3962,N_3564);
nand U6805 (N_6805,N_5212,N_4740);
and U6806 (N_6806,N_3389,N_4427);
xor U6807 (N_6807,N_3168,N_4475);
xnor U6808 (N_6808,N_4022,N_5370);
nand U6809 (N_6809,N_4070,N_3185);
or U6810 (N_6810,N_4681,N_5473);
or U6811 (N_6811,N_4696,N_5814);
and U6812 (N_6812,N_3871,N_5607);
xor U6813 (N_6813,N_3851,N_5686);
nor U6814 (N_6814,N_4201,N_3026);
nor U6815 (N_6815,N_4751,N_5691);
nor U6816 (N_6816,N_4099,N_5634);
nor U6817 (N_6817,N_3827,N_4915);
and U6818 (N_6818,N_4168,N_5280);
and U6819 (N_6819,N_4770,N_4379);
nor U6820 (N_6820,N_3192,N_4952);
and U6821 (N_6821,N_3594,N_4609);
nor U6822 (N_6822,N_4968,N_4185);
nand U6823 (N_6823,N_5684,N_4006);
or U6824 (N_6824,N_5610,N_3330);
xnor U6825 (N_6825,N_4029,N_4199);
nand U6826 (N_6826,N_4175,N_3348);
nor U6827 (N_6827,N_4423,N_5004);
nor U6828 (N_6828,N_3809,N_5898);
xor U6829 (N_6829,N_3527,N_3375);
xor U6830 (N_6830,N_5811,N_4437);
nand U6831 (N_6831,N_5177,N_3322);
and U6832 (N_6832,N_5346,N_4170);
xor U6833 (N_6833,N_5360,N_5807);
or U6834 (N_6834,N_5083,N_3281);
xor U6835 (N_6835,N_4238,N_5801);
nor U6836 (N_6836,N_5537,N_5655);
nand U6837 (N_6837,N_4056,N_3800);
and U6838 (N_6838,N_5125,N_3218);
xor U6839 (N_6839,N_4368,N_4276);
nor U6840 (N_6840,N_4258,N_3730);
or U6841 (N_6841,N_4137,N_4686);
and U6842 (N_6842,N_3304,N_4898);
nand U6843 (N_6843,N_3458,N_4804);
and U6844 (N_6844,N_4002,N_3273);
xnor U6845 (N_6845,N_3503,N_3046);
and U6846 (N_6846,N_5529,N_5545);
or U6847 (N_6847,N_4426,N_3426);
xnor U6848 (N_6848,N_4197,N_5679);
nor U6849 (N_6849,N_3510,N_4597);
nor U6850 (N_6850,N_5188,N_5930);
nand U6851 (N_6851,N_3912,N_5385);
and U6852 (N_6852,N_3039,N_4392);
nand U6853 (N_6853,N_5254,N_4743);
nand U6854 (N_6854,N_4289,N_4180);
or U6855 (N_6855,N_4329,N_4789);
and U6856 (N_6856,N_5926,N_4865);
nand U6857 (N_6857,N_4171,N_5221);
xnor U6858 (N_6858,N_4901,N_5654);
xor U6859 (N_6859,N_5153,N_4972);
and U6860 (N_6860,N_5413,N_5843);
nor U6861 (N_6861,N_5681,N_4651);
and U6862 (N_6862,N_4629,N_4670);
nand U6863 (N_6863,N_5468,N_3445);
and U6864 (N_6864,N_3703,N_4807);
nand U6865 (N_6865,N_4263,N_3641);
nor U6866 (N_6866,N_3998,N_4362);
nand U6867 (N_6867,N_3327,N_4658);
or U6868 (N_6868,N_5105,N_5026);
or U6869 (N_6869,N_3130,N_5072);
nor U6870 (N_6870,N_5303,N_3320);
and U6871 (N_6871,N_3718,N_4540);
nand U6872 (N_6872,N_5598,N_5030);
nand U6873 (N_6873,N_4633,N_4517);
or U6874 (N_6874,N_4679,N_5528);
and U6875 (N_6875,N_3248,N_5602);
nand U6876 (N_6876,N_4752,N_5826);
nor U6877 (N_6877,N_3277,N_4547);
and U6878 (N_6878,N_3453,N_3436);
or U6879 (N_6879,N_3493,N_4721);
xor U6880 (N_6880,N_3197,N_5305);
nor U6881 (N_6881,N_4853,N_5644);
nor U6882 (N_6882,N_4385,N_5570);
xnor U6883 (N_6883,N_5778,N_5620);
xnor U6884 (N_6884,N_3576,N_5271);
nand U6885 (N_6885,N_3408,N_5510);
and U6886 (N_6886,N_3324,N_3844);
or U6887 (N_6887,N_4112,N_3479);
nand U6888 (N_6888,N_5401,N_5848);
xor U6889 (N_6889,N_3279,N_3786);
nor U6890 (N_6890,N_3553,N_5253);
nor U6891 (N_6891,N_3289,N_3287);
nand U6892 (N_6892,N_3260,N_4193);
nor U6893 (N_6893,N_4390,N_3712);
nor U6894 (N_6894,N_5146,N_5518);
xnor U6895 (N_6895,N_3110,N_4166);
nand U6896 (N_6896,N_4264,N_5220);
nand U6897 (N_6897,N_5001,N_4218);
nand U6898 (N_6898,N_4347,N_5050);
nand U6899 (N_6899,N_3132,N_5766);
xnor U6900 (N_6900,N_5875,N_3271);
and U6901 (N_6901,N_4391,N_5526);
xor U6902 (N_6902,N_4956,N_5313);
xor U6903 (N_6903,N_3099,N_3492);
nor U6904 (N_6904,N_4893,N_4943);
and U6905 (N_6905,N_4585,N_5135);
xnor U6906 (N_6906,N_3565,N_3223);
nand U6907 (N_6907,N_3957,N_5577);
xnor U6908 (N_6908,N_3965,N_4539);
or U6909 (N_6909,N_3387,N_3537);
xor U6910 (N_6910,N_3849,N_4235);
nor U6911 (N_6911,N_5813,N_5241);
xor U6912 (N_6912,N_5215,N_3414);
or U6913 (N_6913,N_4978,N_3210);
or U6914 (N_6914,N_3202,N_3810);
xnor U6915 (N_6915,N_4724,N_5505);
nand U6916 (N_6916,N_3838,N_5660);
nand U6917 (N_6917,N_4714,N_4114);
or U6918 (N_6918,N_5056,N_5463);
or U6919 (N_6919,N_4615,N_5457);
and U6920 (N_6920,N_3894,N_5903);
nand U6921 (N_6921,N_3299,N_4381);
nor U6922 (N_6922,N_4625,N_3229);
or U6923 (N_6923,N_4474,N_3352);
or U6924 (N_6924,N_5825,N_4300);
xor U6925 (N_6925,N_5397,N_4626);
nand U6926 (N_6926,N_4048,N_4896);
nand U6927 (N_6927,N_3631,N_3073);
nand U6928 (N_6928,N_5406,N_3113);
nor U6929 (N_6929,N_3481,N_4028);
and U6930 (N_6930,N_5481,N_5737);
nor U6931 (N_6931,N_3012,N_4741);
nand U6932 (N_6932,N_3772,N_3902);
or U6933 (N_6933,N_5804,N_3895);
and U6934 (N_6934,N_4108,N_5390);
nand U6935 (N_6935,N_4047,N_5839);
nor U6936 (N_6936,N_4044,N_3191);
nand U6937 (N_6937,N_5034,N_4719);
and U6938 (N_6938,N_3456,N_4576);
or U6939 (N_6939,N_3294,N_4636);
nand U6940 (N_6940,N_5292,N_5260);
nor U6941 (N_6941,N_5328,N_5029);
nor U6942 (N_6942,N_5797,N_5245);
or U6943 (N_6943,N_3084,N_4671);
and U6944 (N_6944,N_5604,N_4571);
or U6945 (N_6945,N_3405,N_3688);
or U6946 (N_6946,N_4292,N_3963);
nand U6947 (N_6947,N_3092,N_3570);
xor U6948 (N_6948,N_4481,N_3648);
xor U6949 (N_6949,N_3326,N_4224);
and U6950 (N_6950,N_3875,N_4823);
nor U6951 (N_6951,N_3765,N_5799);
and U6952 (N_6952,N_4062,N_5189);
nor U6953 (N_6953,N_4934,N_4076);
xnor U6954 (N_6954,N_3309,N_5961);
nand U6955 (N_6955,N_4847,N_4537);
nand U6956 (N_6956,N_3307,N_3136);
xor U6957 (N_6957,N_5142,N_5409);
or U6958 (N_6958,N_5407,N_5541);
nor U6959 (N_6959,N_3603,N_5091);
nand U6960 (N_6960,N_5054,N_3785);
and U6961 (N_6961,N_3476,N_5356);
nand U6962 (N_6962,N_5016,N_5652);
xor U6963 (N_6963,N_4003,N_4994);
and U6964 (N_6964,N_4287,N_3808);
xor U6965 (N_6965,N_5786,N_5089);
or U6966 (N_6966,N_4526,N_5023);
xnor U6967 (N_6967,N_4699,N_4374);
xor U6968 (N_6968,N_5960,N_5768);
xnor U6969 (N_6969,N_4603,N_5698);
and U6970 (N_6970,N_3163,N_5907);
xor U6971 (N_6971,N_3283,N_4873);
nor U6972 (N_6972,N_3900,N_3390);
xnor U6973 (N_6973,N_4500,N_3276);
and U6974 (N_6974,N_5792,N_3955);
and U6975 (N_6975,N_4927,N_5502);
or U6976 (N_6976,N_4976,N_4333);
nand U6977 (N_6977,N_5025,N_5616);
nor U6978 (N_6978,N_5307,N_5176);
nand U6979 (N_6979,N_3821,N_4953);
or U6980 (N_6980,N_3484,N_4920);
xor U6981 (N_6981,N_3669,N_4089);
xor U6982 (N_6982,N_3873,N_4024);
nor U6983 (N_6983,N_4650,N_4816);
nor U6984 (N_6984,N_4666,N_3141);
or U6985 (N_6985,N_3149,N_5824);
or U6986 (N_6986,N_5093,N_5741);
or U6987 (N_6987,N_5662,N_5130);
nand U6988 (N_6988,N_5233,N_5395);
or U6989 (N_6989,N_3007,N_5263);
and U6990 (N_6990,N_4884,N_3734);
nor U6991 (N_6991,N_3224,N_3069);
nand U6992 (N_6992,N_3745,N_3144);
and U6993 (N_6993,N_3500,N_3114);
and U6994 (N_6994,N_5076,N_3107);
or U6995 (N_6995,N_3704,N_3486);
nor U6996 (N_6996,N_5793,N_4155);
nand U6997 (N_6997,N_5250,N_3172);
or U6998 (N_6998,N_4007,N_3805);
nor U6999 (N_6999,N_5669,N_3208);
nand U7000 (N_7000,N_4937,N_4919);
nor U7001 (N_7001,N_5554,N_4142);
nor U7002 (N_7002,N_4376,N_5501);
or U7003 (N_7003,N_5773,N_5856);
xor U7004 (N_7004,N_4194,N_4295);
xor U7005 (N_7005,N_4412,N_4705);
and U7006 (N_7006,N_4644,N_3444);
xnor U7007 (N_7007,N_5992,N_4268);
xnor U7008 (N_7008,N_4643,N_5400);
nand U7009 (N_7009,N_3388,N_4387);
nand U7010 (N_7010,N_4689,N_5589);
and U7011 (N_7011,N_5868,N_5719);
and U7012 (N_7012,N_3022,N_3802);
xor U7013 (N_7013,N_4436,N_3868);
and U7014 (N_7014,N_4722,N_4280);
xnor U7015 (N_7015,N_5179,N_5469);
and U7016 (N_7016,N_4885,N_4491);
and U7017 (N_7017,N_3970,N_4179);
and U7018 (N_7018,N_3797,N_5608);
nor U7019 (N_7019,N_4560,N_3265);
nand U7020 (N_7020,N_3469,N_5137);
nand U7021 (N_7021,N_4797,N_3776);
xor U7022 (N_7022,N_5498,N_4506);
nand U7023 (N_7023,N_3629,N_4084);
and U7024 (N_7024,N_5191,N_4208);
or U7025 (N_7025,N_3681,N_3615);
or U7026 (N_7026,N_5675,N_4403);
nand U7027 (N_7027,N_3761,N_3480);
or U7028 (N_7028,N_4191,N_4086);
nand U7029 (N_7029,N_4554,N_3063);
xor U7030 (N_7030,N_5002,N_3259);
and U7031 (N_7031,N_5208,N_4134);
and U7032 (N_7032,N_4425,N_4184);
nor U7033 (N_7033,N_4858,N_3374);
and U7034 (N_7034,N_5853,N_4151);
or U7035 (N_7035,N_5910,N_3517);
nor U7036 (N_7036,N_5070,N_3473);
and U7037 (N_7037,N_3948,N_3066);
nand U7038 (N_7038,N_3884,N_4567);
or U7039 (N_7039,N_5886,N_5290);
nand U7040 (N_7040,N_4401,N_4259);
nand U7041 (N_7041,N_3472,N_4036);
or U7042 (N_7042,N_4065,N_5651);
or U7043 (N_7043,N_4660,N_3890);
and U7044 (N_7044,N_5445,N_4439);
and U7045 (N_7045,N_4936,N_5009);
and U7046 (N_7046,N_4252,N_3949);
nor U7047 (N_7047,N_4318,N_4607);
nor U7048 (N_7048,N_3442,N_4655);
and U7049 (N_7049,N_3135,N_5459);
nor U7050 (N_7050,N_5116,N_5277);
nor U7051 (N_7051,N_3109,N_3918);
and U7052 (N_7052,N_5078,N_3632);
nor U7053 (N_7053,N_4442,N_3448);
or U7054 (N_7054,N_5967,N_5689);
nor U7055 (N_7055,N_3321,N_5594);
nand U7056 (N_7056,N_5109,N_3122);
and U7057 (N_7057,N_5165,N_4032);
and U7058 (N_7058,N_4505,N_3757);
xor U7059 (N_7059,N_5237,N_3108);
nor U7060 (N_7060,N_5635,N_4355);
or U7061 (N_7061,N_5098,N_4871);
nand U7062 (N_7062,N_3459,N_5200);
or U7063 (N_7063,N_4205,N_3085);
nor U7064 (N_7064,N_4811,N_4261);
and U7065 (N_7065,N_3006,N_5379);
nand U7066 (N_7066,N_5500,N_3371);
nand U7067 (N_7067,N_3119,N_3411);
and U7068 (N_7068,N_5039,N_3914);
nand U7069 (N_7069,N_3146,N_3828);
nand U7070 (N_7070,N_5859,N_3171);
nor U7071 (N_7071,N_3869,N_5936);
nand U7072 (N_7072,N_3345,N_3056);
or U7073 (N_7073,N_3578,N_5308);
xnor U7074 (N_7074,N_5419,N_4706);
xnor U7075 (N_7075,N_5082,N_4911);
nor U7076 (N_7076,N_4525,N_5020);
nor U7077 (N_7077,N_5256,N_3920);
xnor U7078 (N_7078,N_4673,N_5667);
and U7079 (N_7079,N_5159,N_5386);
or U7080 (N_7080,N_4759,N_5784);
or U7081 (N_7081,N_3048,N_4147);
or U7082 (N_7082,N_4548,N_5672);
and U7083 (N_7083,N_5998,N_4183);
or U7084 (N_7084,N_5230,N_4602);
or U7085 (N_7085,N_5587,N_5613);
and U7086 (N_7086,N_3695,N_4906);
or U7087 (N_7087,N_3845,N_4703);
nand U7088 (N_7088,N_4413,N_4827);
or U7089 (N_7089,N_4489,N_4590);
or U7090 (N_7090,N_3463,N_5677);
and U7091 (N_7091,N_4127,N_5035);
nand U7092 (N_7092,N_3123,N_3106);
xnor U7093 (N_7093,N_3568,N_3204);
and U7094 (N_7094,N_4769,N_4659);
nor U7095 (N_7095,N_3213,N_3194);
xnor U7096 (N_7096,N_3769,N_3944);
or U7097 (N_7097,N_4528,N_5963);
or U7098 (N_7098,N_3635,N_3714);
and U7099 (N_7099,N_3305,N_3721);
nand U7100 (N_7100,N_5700,N_5232);
xnor U7101 (N_7101,N_5169,N_4200);
or U7102 (N_7102,N_3879,N_5983);
xnor U7103 (N_7103,N_3737,N_4121);
and U7104 (N_7104,N_5167,N_3009);
xor U7105 (N_7105,N_5771,N_3251);
or U7106 (N_7106,N_4519,N_5073);
nor U7107 (N_7107,N_3263,N_4478);
or U7108 (N_7108,N_3240,N_3222);
xor U7109 (N_7109,N_3886,N_3853);
xor U7110 (N_7110,N_5321,N_3612);
or U7111 (N_7111,N_5156,N_3120);
nand U7112 (N_7112,N_3701,N_4754);
xnor U7113 (N_7113,N_3138,N_4195);
xor U7114 (N_7114,N_5981,N_5938);
or U7115 (N_7115,N_4219,N_4431);
and U7116 (N_7116,N_4835,N_3460);
nand U7117 (N_7117,N_4803,N_4709);
xor U7118 (N_7118,N_3250,N_5916);
and U7119 (N_7119,N_3058,N_3337);
or U7120 (N_7120,N_5408,N_4950);
and U7121 (N_7121,N_5389,N_3180);
nand U7122 (N_7122,N_3605,N_3306);
nand U7123 (N_7123,N_4113,N_4569);
or U7124 (N_7124,N_4557,N_4693);
nand U7125 (N_7125,N_5947,N_3579);
xor U7126 (N_7126,N_4947,N_3709);
or U7127 (N_7127,N_4266,N_3859);
and U7128 (N_7128,N_3560,N_4313);
or U7129 (N_7129,N_5335,N_5670);
nand U7130 (N_7130,N_3788,N_4384);
and U7131 (N_7131,N_5637,N_3068);
nor U7132 (N_7132,N_5384,N_3687);
nor U7133 (N_7133,N_4815,N_5048);
nand U7134 (N_7134,N_4369,N_4799);
xor U7135 (N_7135,N_5032,N_5454);
xor U7136 (N_7136,N_5316,N_3563);
and U7137 (N_7137,N_4339,N_3752);
and U7138 (N_7138,N_5304,N_5753);
and U7139 (N_7139,N_5701,N_4234);
nor U7140 (N_7140,N_3001,N_4042);
or U7141 (N_7141,N_4538,N_3246);
nor U7142 (N_7142,N_4702,N_3243);
and U7143 (N_7143,N_4676,N_4910);
or U7144 (N_7144,N_5418,N_4012);
and U7145 (N_7145,N_4104,N_5434);
nand U7146 (N_7146,N_3979,N_3724);
or U7147 (N_7147,N_3365,N_4982);
or U7148 (N_7148,N_4192,N_4690);
xor U7149 (N_7149,N_3158,N_3519);
nand U7150 (N_7150,N_3569,N_4061);
and U7151 (N_7151,N_3407,N_5850);
nand U7152 (N_7152,N_3983,N_3837);
xor U7153 (N_7153,N_4611,N_5582);
nor U7154 (N_7154,N_4245,N_4866);
nand U7155 (N_7155,N_3147,N_3098);
nor U7156 (N_7156,N_4836,N_5202);
or U7157 (N_7157,N_5543,N_5244);
nand U7158 (N_7158,N_5455,N_3758);
or U7159 (N_7159,N_5512,N_3692);
or U7160 (N_7160,N_4883,N_4750);
xor U7161 (N_7161,N_4974,N_3645);
nand U7162 (N_7162,N_3888,N_4544);
or U7163 (N_7163,N_5475,N_5744);
xnor U7164 (N_7164,N_3255,N_4304);
nor U7165 (N_7165,N_5519,N_4241);
nand U7166 (N_7166,N_5110,N_5809);
and U7167 (N_7167,N_4922,N_3188);
nand U7168 (N_7168,N_4555,N_3904);
xor U7169 (N_7169,N_3380,N_4071);
nand U7170 (N_7170,N_5104,N_3534);
and U7171 (N_7171,N_3082,N_3252);
or U7172 (N_7172,N_5195,N_5694);
xor U7173 (N_7173,N_3452,N_3930);
nor U7174 (N_7174,N_3219,N_4692);
nor U7175 (N_7175,N_5597,N_5727);
nand U7176 (N_7176,N_5618,N_3331);
or U7177 (N_7177,N_4317,N_5474);
nor U7178 (N_7178,N_5017,N_5711);
or U7179 (N_7179,N_4054,N_5708);
nor U7180 (N_7180,N_3866,N_3833);
xor U7181 (N_7181,N_3661,N_3349);
nand U7182 (N_7182,N_4509,N_3328);
or U7183 (N_7183,N_4942,N_3928);
nor U7184 (N_7184,N_3667,N_4802);
or U7185 (N_7185,N_3595,N_5657);
nor U7186 (N_7186,N_4832,N_3051);
or U7187 (N_7187,N_5647,N_4398);
nand U7188 (N_7188,N_5697,N_5816);
nand U7189 (N_7189,N_5238,N_5127);
and U7190 (N_7190,N_3037,N_5970);
nand U7191 (N_7191,N_5268,N_5609);
xnor U7192 (N_7192,N_3573,N_4375);
and U7193 (N_7193,N_4551,N_5511);
nand U7194 (N_7194,N_5732,N_4825);
and U7195 (N_7195,N_4565,N_4040);
xor U7196 (N_7196,N_4494,N_3301);
or U7197 (N_7197,N_3795,N_5601);
and U7198 (N_7198,N_3950,N_5038);
nor U7199 (N_7199,N_3230,N_5046);
and U7200 (N_7200,N_5683,N_4654);
nand U7201 (N_7201,N_5465,N_5160);
nand U7202 (N_7202,N_5525,N_3952);
nor U7203 (N_7203,N_4091,N_4009);
or U7204 (N_7204,N_3780,N_4187);
and U7205 (N_7205,N_4285,N_4522);
xnor U7206 (N_7206,N_3882,N_3824);
nor U7207 (N_7207,N_4081,N_5984);
and U7208 (N_7208,N_5123,N_5932);
and U7209 (N_7209,N_4053,N_5986);
or U7210 (N_7210,N_5037,N_5965);
or U7211 (N_7211,N_4598,N_4130);
nand U7212 (N_7212,N_4215,N_5976);
xor U7213 (N_7213,N_4103,N_5523);
nor U7214 (N_7214,N_3187,N_5282);
xor U7215 (N_7215,N_4394,N_4627);
and U7216 (N_7216,N_5264,N_5011);
xnor U7217 (N_7217,N_5331,N_5325);
xor U7218 (N_7218,N_3212,N_5957);
or U7219 (N_7219,N_3616,N_4921);
nor U7220 (N_7220,N_3505,N_3885);
or U7221 (N_7221,N_5790,N_4907);
or U7222 (N_7222,N_4552,N_4501);
xor U7223 (N_7223,N_4322,N_5447);
and U7224 (N_7224,N_5404,N_5199);
or U7225 (N_7225,N_5869,N_4176);
xnor U7226 (N_7226,N_5164,N_4997);
nand U7227 (N_7227,N_4360,N_5663);
and U7228 (N_7228,N_3621,N_4889);
nand U7229 (N_7229,N_3443,N_5209);
or U7230 (N_7230,N_4954,N_4902);
nor U7231 (N_7231,N_4066,N_4253);
nor U7232 (N_7232,N_3796,N_3665);
nand U7233 (N_7233,N_5544,N_3162);
xnor U7234 (N_7234,N_5080,N_4680);
nand U7235 (N_7235,N_3118,N_3658);
and U7236 (N_7236,N_3067,N_3111);
nor U7237 (N_7237,N_3199,N_5126);
nor U7238 (N_7238,N_5464,N_3433);
and U7239 (N_7239,N_3142,N_3427);
nand U7240 (N_7240,N_5088,N_5643);
nand U7241 (N_7241,N_5563,N_4161);
nand U7242 (N_7242,N_3288,N_5767);
nor U7243 (N_7243,N_4684,N_5437);
nand U7244 (N_7244,N_5433,N_4090);
or U7245 (N_7245,N_5113,N_4647);
nand U7246 (N_7246,N_5227,N_5466);
and U7247 (N_7247,N_4521,N_3674);
xor U7248 (N_7248,N_4141,N_3990);
nor U7249 (N_7249,N_3160,N_5599);
and U7250 (N_7250,N_4204,N_4558);
nor U7251 (N_7251,N_5849,N_5783);
xor U7252 (N_7252,N_5551,N_4421);
nand U7253 (N_7253,N_5688,N_3074);
and U7254 (N_7254,N_3189,N_3611);
xor U7255 (N_7255,N_5012,N_4074);
nor U7256 (N_7256,N_3829,N_4357);
nand U7257 (N_7257,N_4808,N_5045);
and U7258 (N_7258,N_3625,N_3195);
nor U7259 (N_7259,N_5918,N_5606);
and U7260 (N_7260,N_4327,N_5873);
xnor U7261 (N_7261,N_4162,N_4697);
nand U7262 (N_7262,N_4833,N_3846);
nand U7263 (N_7263,N_5198,N_5891);
nor U7264 (N_7264,N_5956,N_3102);
nor U7265 (N_7265,N_4587,N_4447);
or U7266 (N_7266,N_5889,N_4277);
nand U7267 (N_7267,N_3334,N_3008);
or U7268 (N_7268,N_3435,N_3583);
or U7269 (N_7269,N_4025,N_4917);
or U7270 (N_7270,N_4145,N_5586);
and U7271 (N_7271,N_3487,N_3315);
or U7272 (N_7272,N_4377,N_4308);
nand U7273 (N_7273,N_5823,N_5240);
xnor U7274 (N_7274,N_3746,N_3344);
and U7275 (N_7275,N_5145,N_5348);
nor U7276 (N_7276,N_4169,N_3392);
or U7277 (N_7277,N_4471,N_5309);
nor U7278 (N_7278,N_3750,N_5226);
and U7279 (N_7279,N_4995,N_3178);
xnor U7280 (N_7280,N_3961,N_5837);
and U7281 (N_7281,N_4820,N_5830);
nand U7282 (N_7282,N_4311,N_5201);
or U7283 (N_7283,N_5344,N_4085);
or U7284 (N_7284,N_5319,N_5803);
nor U7285 (N_7285,N_3121,N_5623);
xnor U7286 (N_7286,N_5107,N_5845);
xor U7287 (N_7287,N_5477,N_3441);
and U7288 (N_7288,N_5373,N_5018);
or U7289 (N_7289,N_5516,N_5631);
nor U7290 (N_7290,N_4813,N_5877);
nand U7291 (N_7291,N_3559,N_5338);
xnor U7292 (N_7292,N_3419,N_4310);
xnor U7293 (N_7293,N_5530,N_3716);
and U7294 (N_7294,N_5949,N_4075);
and U7295 (N_7295,N_4731,N_4985);
nand U7296 (N_7296,N_3040,N_3300);
or U7297 (N_7297,N_5748,N_3182);
xor U7298 (N_7298,N_4599,N_4356);
nand U7299 (N_7299,N_4354,N_4785);
and U7300 (N_7300,N_5403,N_5150);
nor U7301 (N_7301,N_5820,N_4446);
and U7302 (N_7302,N_5573,N_3547);
or U7303 (N_7303,N_3726,N_3173);
xor U7304 (N_7304,N_4111,N_3090);
or U7305 (N_7305,N_4093,N_4518);
and U7306 (N_7306,N_4186,N_4480);
xnor U7307 (N_7307,N_5946,N_3014);
xnor U7308 (N_7308,N_5499,N_5659);
nand U7309 (N_7309,N_5117,N_4862);
or U7310 (N_7310,N_5828,N_3235);
and U7311 (N_7311,N_3377,N_5507);
nor U7312 (N_7312,N_3417,N_4717);
xnor U7313 (N_7313,N_4661,N_4531);
xnor U7314 (N_7314,N_3253,N_5781);
nand U7315 (N_7315,N_3451,N_3395);
and U7316 (N_7316,N_3813,N_5881);
nor U7317 (N_7317,N_5870,N_3791);
and U7318 (N_7318,N_5695,N_4524);
or U7319 (N_7319,N_4043,N_3551);
nand U7320 (N_7320,N_3984,N_4630);
and U7321 (N_7321,N_4301,N_4592);
nor U7322 (N_7322,N_3652,N_5756);
nand U7323 (N_7323,N_4913,N_3532);
and U7324 (N_7324,N_4305,N_3355);
and U7325 (N_7325,N_5515,N_5311);
nand U7326 (N_7326,N_4077,N_4616);
and U7327 (N_7327,N_3043,N_4294);
or U7328 (N_7328,N_5509,N_4718);
nand U7329 (N_7329,N_5443,N_3518);
or U7330 (N_7330,N_5329,N_3234);
nor U7331 (N_7331,N_5879,N_4469);
xnor U7332 (N_7332,N_4315,N_3561);
and U7333 (N_7333,N_5154,N_5815);
or U7334 (N_7334,N_3557,N_3139);
and U7335 (N_7335,N_3520,N_3907);
nor U7336 (N_7336,N_4900,N_3310);
nand U7337 (N_7337,N_4227,N_4675);
xnor U7338 (N_7338,N_4297,N_4894);
or U7339 (N_7339,N_5262,N_4966);
nand U7340 (N_7340,N_4623,N_4181);
xor U7341 (N_7341,N_3205,N_3996);
and U7342 (N_7342,N_4220,N_4453);
nand U7343 (N_7343,N_3840,N_4472);
xnor U7344 (N_7344,N_4281,N_5115);
nor U7345 (N_7345,N_4879,N_4739);
and U7346 (N_7346,N_5133,N_4667);
nor U7347 (N_7347,N_5449,N_3736);
nand U7348 (N_7348,N_3760,N_4299);
and U7349 (N_7349,N_3200,N_4886);
and U7350 (N_7350,N_4700,N_5840);
nor U7351 (N_7351,N_3628,N_3125);
xor U7352 (N_7352,N_4283,N_3157);
xor U7353 (N_7353,N_4079,N_5559);
xnor U7354 (N_7354,N_3050,N_3768);
xnor U7355 (N_7355,N_5906,N_5112);
or U7356 (N_7356,N_4255,N_3689);
nand U7357 (N_7357,N_4367,N_4274);
nand U7358 (N_7358,N_5605,N_5246);
nor U7359 (N_7359,N_5151,N_3401);
and U7360 (N_7360,N_5883,N_3784);
xnor U7361 (N_7361,N_5444,N_3664);
nor U7362 (N_7362,N_4288,N_4190);
xor U7363 (N_7363,N_4302,N_3657);
xnor U7364 (N_7364,N_3032,N_4711);
and U7365 (N_7365,N_5210,N_3617);
or U7366 (N_7366,N_3247,N_5712);
nand U7367 (N_7367,N_5997,N_4923);
xor U7368 (N_7368,N_3360,N_5423);
or U7369 (N_7369,N_4404,N_3523);
nor U7370 (N_7370,N_5219,N_3482);
or U7371 (N_7371,N_3285,N_4364);
or U7372 (N_7372,N_5715,N_5583);
and U7373 (N_7373,N_5484,N_5342);
xnor U7374 (N_7374,N_5027,N_4874);
nor U7375 (N_7375,N_5286,N_4363);
nand U7376 (N_7376,N_3164,N_5649);
nor U7377 (N_7377,N_4038,N_5721);
nand U7378 (N_7378,N_4747,N_3899);
xnor U7379 (N_7379,N_4449,N_3820);
or U7380 (N_7380,N_5923,N_5980);
and U7381 (N_7381,N_5170,N_3815);
xor U7382 (N_7382,N_5911,N_4095);
xor U7383 (N_7383,N_3947,N_4102);
or U7384 (N_7384,N_5802,N_3945);
xnor U7385 (N_7385,N_3575,N_5927);
xor U7386 (N_7386,N_3086,N_4371);
and U7387 (N_7387,N_5420,N_3237);
or U7388 (N_7388,N_4129,N_4744);
or U7389 (N_7389,N_4757,N_4428);
xor U7390 (N_7390,N_3872,N_4546);
xor U7391 (N_7391,N_3855,N_4778);
and U7392 (N_7392,N_3030,N_5593);
and U7393 (N_7393,N_3137,N_3015);
nand U7394 (N_7394,N_5347,N_3975);
nor U7395 (N_7395,N_3722,N_3956);
xnor U7396 (N_7396,N_3280,N_5882);
nor U7397 (N_7397,N_5832,N_3233);
nor U7398 (N_7398,N_3096,N_3771);
nand U7399 (N_7399,N_4466,N_5461);
or U7400 (N_7400,N_4553,N_4793);
and U7401 (N_7401,N_3317,N_3651);
nor U7402 (N_7402,N_3848,N_4148);
or U7403 (N_7403,N_4260,N_3397);
nand U7404 (N_7404,N_5628,N_5546);
or U7405 (N_7405,N_3608,N_4512);
nor U7406 (N_7406,N_5527,N_3175);
nor U7407 (N_7407,N_3366,N_4087);
xnor U7408 (N_7408,N_3496,N_3424);
nand U7409 (N_7409,N_5111,N_3656);
nor U7410 (N_7410,N_5808,N_3339);
or U7411 (N_7411,N_4877,N_5805);
xor U7412 (N_7412,N_3363,N_5763);
nand U7413 (N_7413,N_5739,N_3338);
nand U7414 (N_7414,N_3333,N_3062);
and U7415 (N_7415,N_3711,N_3964);
xnor U7416 (N_7416,N_4768,N_3993);
nor U7417 (N_7417,N_4286,N_5178);
nand U7418 (N_7418,N_3571,N_5958);
or U7419 (N_7419,N_4733,N_5496);
xor U7420 (N_7420,N_4352,N_5487);
or U7421 (N_7421,N_5817,N_5106);
or U7422 (N_7422,N_5603,N_4841);
and U7423 (N_7423,N_5103,N_3396);
nor U7424 (N_7424,N_5738,N_3816);
xnor U7425 (N_7425,N_3356,N_3284);
nand U7426 (N_7426,N_3946,N_3906);
and U7427 (N_7427,N_5720,N_5735);
nand U7428 (N_7428,N_5494,N_4591);
nor U7429 (N_7429,N_5207,N_4588);
xnor U7430 (N_7430,N_4406,N_3939);
or U7431 (N_7431,N_5539,N_5725);
or U7432 (N_7432,N_3329,N_4140);
nand U7433 (N_7433,N_3798,N_3384);
nor U7434 (N_7434,N_4303,N_4461);
nor U7435 (N_7435,N_5085,N_3080);
nor U7436 (N_7436,N_5051,N_3577);
xor U7437 (N_7437,N_3535,N_5555);
nor U7438 (N_7438,N_3803,N_3295);
nand U7439 (N_7439,N_5003,N_5640);
and U7440 (N_7440,N_3554,N_4052);
xor U7441 (N_7441,N_4396,N_3640);
and U7442 (N_7442,N_3986,N_3489);
or U7443 (N_7443,N_3005,N_4417);
or U7444 (N_7444,N_5345,N_5533);
or U7445 (N_7445,N_4800,N_3558);
nor U7446 (N_7446,N_5951,N_4163);
nor U7447 (N_7447,N_4657,N_3400);
or U7448 (N_7448,N_5380,N_3089);
xor U7449 (N_7449,N_3038,N_3790);
xor U7450 (N_7450,N_3587,N_5166);
or U7451 (N_7451,N_3574,N_5022);
or U7452 (N_7452,N_3216,N_5665);
or U7453 (N_7453,N_5057,N_4946);
or U7454 (N_7454,N_5267,N_3887);
and U7455 (N_7455,N_3023,N_3450);
and U7456 (N_7456,N_3298,N_3311);
nor U7457 (N_7457,N_4465,N_4581);
and U7458 (N_7458,N_5414,N_5276);
nor U7459 (N_7459,N_3931,N_5183);
nor U7460 (N_7460,N_3316,N_5061);
xnor U7461 (N_7461,N_5880,N_3847);
or U7462 (N_7462,N_5893,N_3346);
or U7463 (N_7463,N_5327,N_5424);
xnor U7464 (N_7464,N_3385,N_3874);
nor U7465 (N_7465,N_5099,N_5064);
and U7466 (N_7466,N_4458,N_3091);
and U7467 (N_7467,N_4566,N_4533);
or U7468 (N_7468,N_4958,N_5138);
and U7469 (N_7469,N_4812,N_3159);
and U7470 (N_7470,N_5785,N_5438);
xor U7471 (N_7471,N_5139,N_4314);
nand U7472 (N_7472,N_3915,N_5216);
and U7473 (N_7473,N_5314,N_5504);
nor U7474 (N_7474,N_5611,N_3804);
and U7475 (N_7475,N_3412,N_3457);
or U7476 (N_7476,N_4063,N_4993);
and U7477 (N_7477,N_3590,N_5265);
or U7478 (N_7478,N_3211,N_3980);
nand U7479 (N_7479,N_4957,N_5514);
xor U7480 (N_7480,N_5248,N_4212);
and U7481 (N_7481,N_4273,N_5005);
xnor U7482 (N_7482,N_3783,N_3966);
xnor U7483 (N_7483,N_5402,N_5118);
nand U7484 (N_7484,N_4674,N_4240);
xor U7485 (N_7485,N_4549,N_3935);
or U7486 (N_7486,N_5917,N_4568);
nor U7487 (N_7487,N_3341,N_4845);
xor U7488 (N_7488,N_3599,N_3465);
nand U7489 (N_7489,N_4726,N_5975);
xnor U7490 (N_7490,N_3933,N_4452);
xnor U7491 (N_7491,N_4242,N_5412);
xor U7492 (N_7492,N_3618,N_5310);
or U7493 (N_7493,N_4251,N_4041);
and U7494 (N_7494,N_4905,N_3423);
nand U7495 (N_7495,N_3471,N_3418);
nand U7496 (N_7496,N_3290,N_5322);
or U7497 (N_7497,N_4781,N_3951);
or U7498 (N_7498,N_4230,N_4550);
and U7499 (N_7499,N_5995,N_4348);
nor U7500 (N_7500,N_4183,N_3368);
or U7501 (N_7501,N_3942,N_4793);
xor U7502 (N_7502,N_5052,N_3335);
xnor U7503 (N_7503,N_3384,N_5787);
or U7504 (N_7504,N_3132,N_5136);
and U7505 (N_7505,N_5561,N_3075);
or U7506 (N_7506,N_3337,N_5990);
or U7507 (N_7507,N_3671,N_3480);
nand U7508 (N_7508,N_5246,N_3312);
and U7509 (N_7509,N_4748,N_5341);
and U7510 (N_7510,N_4824,N_4271);
nand U7511 (N_7511,N_3134,N_4674);
xnor U7512 (N_7512,N_3173,N_5337);
xor U7513 (N_7513,N_3419,N_3836);
nand U7514 (N_7514,N_5314,N_3010);
and U7515 (N_7515,N_5865,N_5604);
or U7516 (N_7516,N_4481,N_5382);
or U7517 (N_7517,N_3694,N_5685);
xnor U7518 (N_7518,N_5420,N_3240);
or U7519 (N_7519,N_5878,N_3182);
and U7520 (N_7520,N_5508,N_3725);
or U7521 (N_7521,N_5170,N_4883);
nor U7522 (N_7522,N_3179,N_4323);
or U7523 (N_7523,N_4641,N_3560);
nand U7524 (N_7524,N_5550,N_4889);
and U7525 (N_7525,N_5815,N_4479);
and U7526 (N_7526,N_4155,N_5177);
or U7527 (N_7527,N_5289,N_3076);
nand U7528 (N_7528,N_3188,N_5467);
or U7529 (N_7529,N_4999,N_3604);
and U7530 (N_7530,N_3681,N_4019);
or U7531 (N_7531,N_3341,N_5585);
nand U7532 (N_7532,N_3215,N_5578);
and U7533 (N_7533,N_3351,N_5589);
and U7534 (N_7534,N_4252,N_5519);
xnor U7535 (N_7535,N_5867,N_4786);
xor U7536 (N_7536,N_3856,N_5549);
and U7537 (N_7537,N_5959,N_3074);
nor U7538 (N_7538,N_4732,N_3660);
xnor U7539 (N_7539,N_4933,N_3604);
nor U7540 (N_7540,N_4543,N_5392);
and U7541 (N_7541,N_4786,N_5627);
nor U7542 (N_7542,N_3656,N_3292);
and U7543 (N_7543,N_4812,N_4396);
nor U7544 (N_7544,N_3582,N_4605);
nor U7545 (N_7545,N_4989,N_4224);
nor U7546 (N_7546,N_3330,N_4647);
and U7547 (N_7547,N_5840,N_4471);
and U7548 (N_7548,N_4161,N_3888);
xor U7549 (N_7549,N_5017,N_4630);
nor U7550 (N_7550,N_3610,N_3005);
nor U7551 (N_7551,N_3149,N_5520);
nand U7552 (N_7552,N_3955,N_4255);
and U7553 (N_7553,N_3647,N_4659);
xnor U7554 (N_7554,N_4061,N_4162);
nor U7555 (N_7555,N_4886,N_3921);
nand U7556 (N_7556,N_5493,N_5799);
xor U7557 (N_7557,N_5054,N_3643);
xor U7558 (N_7558,N_4488,N_5695);
nand U7559 (N_7559,N_4918,N_3941);
nand U7560 (N_7560,N_5053,N_4145);
nand U7561 (N_7561,N_4776,N_4606);
and U7562 (N_7562,N_4925,N_4566);
and U7563 (N_7563,N_5704,N_3057);
and U7564 (N_7564,N_4890,N_3435);
or U7565 (N_7565,N_4484,N_4430);
or U7566 (N_7566,N_3917,N_5781);
or U7567 (N_7567,N_5826,N_4419);
nor U7568 (N_7568,N_3741,N_5229);
and U7569 (N_7569,N_5436,N_4735);
or U7570 (N_7570,N_3081,N_4003);
and U7571 (N_7571,N_4135,N_3454);
xor U7572 (N_7572,N_3367,N_4373);
nand U7573 (N_7573,N_5374,N_3666);
xnor U7574 (N_7574,N_4023,N_5205);
xor U7575 (N_7575,N_5956,N_4456);
and U7576 (N_7576,N_3739,N_3478);
nor U7577 (N_7577,N_3571,N_5945);
or U7578 (N_7578,N_5603,N_4252);
nor U7579 (N_7579,N_3846,N_3865);
nor U7580 (N_7580,N_4610,N_4157);
nand U7581 (N_7581,N_5693,N_5391);
xnor U7582 (N_7582,N_3096,N_3250);
xnor U7583 (N_7583,N_5891,N_5602);
nand U7584 (N_7584,N_5851,N_4596);
or U7585 (N_7585,N_4341,N_5367);
nor U7586 (N_7586,N_5660,N_4510);
or U7587 (N_7587,N_5822,N_3737);
and U7588 (N_7588,N_3358,N_4741);
xor U7589 (N_7589,N_4512,N_4313);
nor U7590 (N_7590,N_5202,N_5904);
nand U7591 (N_7591,N_3539,N_4632);
xnor U7592 (N_7592,N_4069,N_5452);
nand U7593 (N_7593,N_3262,N_4729);
and U7594 (N_7594,N_5006,N_5635);
and U7595 (N_7595,N_3436,N_3945);
nand U7596 (N_7596,N_4221,N_5754);
nor U7597 (N_7597,N_4249,N_5938);
nand U7598 (N_7598,N_3453,N_4261);
nand U7599 (N_7599,N_5621,N_3624);
nor U7600 (N_7600,N_4528,N_5953);
xnor U7601 (N_7601,N_3929,N_5130);
nand U7602 (N_7602,N_3463,N_5980);
xnor U7603 (N_7603,N_5240,N_5534);
nand U7604 (N_7604,N_3798,N_3103);
xnor U7605 (N_7605,N_4469,N_3225);
nor U7606 (N_7606,N_3955,N_5075);
xnor U7607 (N_7607,N_5673,N_4614);
nor U7608 (N_7608,N_3865,N_3932);
and U7609 (N_7609,N_4929,N_4985);
nand U7610 (N_7610,N_3058,N_4814);
and U7611 (N_7611,N_4534,N_3761);
and U7612 (N_7612,N_3629,N_5241);
xor U7613 (N_7613,N_4693,N_5954);
nor U7614 (N_7614,N_3361,N_3338);
and U7615 (N_7615,N_4001,N_4569);
nand U7616 (N_7616,N_5761,N_5541);
xor U7617 (N_7617,N_3122,N_5295);
and U7618 (N_7618,N_3791,N_5393);
and U7619 (N_7619,N_4990,N_4773);
or U7620 (N_7620,N_5116,N_3553);
nor U7621 (N_7621,N_5360,N_4965);
xor U7622 (N_7622,N_3927,N_3329);
xnor U7623 (N_7623,N_3232,N_4520);
nand U7624 (N_7624,N_5265,N_3247);
or U7625 (N_7625,N_4792,N_3371);
and U7626 (N_7626,N_3796,N_3393);
and U7627 (N_7627,N_3711,N_5381);
or U7628 (N_7628,N_3457,N_4464);
nand U7629 (N_7629,N_4183,N_5542);
or U7630 (N_7630,N_4115,N_4190);
xnor U7631 (N_7631,N_4448,N_4103);
or U7632 (N_7632,N_5364,N_3274);
and U7633 (N_7633,N_4495,N_4716);
nor U7634 (N_7634,N_5029,N_3069);
or U7635 (N_7635,N_3353,N_4626);
or U7636 (N_7636,N_4787,N_5003);
nor U7637 (N_7637,N_3383,N_3962);
and U7638 (N_7638,N_4342,N_3685);
nand U7639 (N_7639,N_3891,N_5618);
nand U7640 (N_7640,N_4089,N_5062);
nor U7641 (N_7641,N_3415,N_3940);
nand U7642 (N_7642,N_5116,N_3100);
nor U7643 (N_7643,N_4758,N_5144);
nand U7644 (N_7644,N_5693,N_5524);
nor U7645 (N_7645,N_4715,N_4812);
or U7646 (N_7646,N_3661,N_4849);
nand U7647 (N_7647,N_4115,N_5730);
and U7648 (N_7648,N_4806,N_3196);
or U7649 (N_7649,N_5436,N_4125);
nor U7650 (N_7650,N_3821,N_3183);
or U7651 (N_7651,N_4570,N_5380);
and U7652 (N_7652,N_3820,N_5820);
xnor U7653 (N_7653,N_5456,N_3455);
or U7654 (N_7654,N_3359,N_3635);
or U7655 (N_7655,N_4413,N_4605);
and U7656 (N_7656,N_5221,N_5241);
nand U7657 (N_7657,N_5317,N_3605);
nor U7658 (N_7658,N_3293,N_5545);
nor U7659 (N_7659,N_5696,N_5956);
nor U7660 (N_7660,N_5811,N_3306);
nand U7661 (N_7661,N_5936,N_3588);
and U7662 (N_7662,N_3848,N_5355);
nor U7663 (N_7663,N_5462,N_3516);
and U7664 (N_7664,N_4478,N_3455);
and U7665 (N_7665,N_3295,N_5899);
and U7666 (N_7666,N_5438,N_4997);
or U7667 (N_7667,N_4897,N_5305);
or U7668 (N_7668,N_5116,N_4464);
or U7669 (N_7669,N_4289,N_3561);
and U7670 (N_7670,N_5302,N_3076);
or U7671 (N_7671,N_4032,N_5690);
or U7672 (N_7672,N_5674,N_4071);
nand U7673 (N_7673,N_3017,N_5242);
nand U7674 (N_7674,N_5371,N_3899);
and U7675 (N_7675,N_3729,N_3349);
nor U7676 (N_7676,N_4753,N_4092);
nand U7677 (N_7677,N_5416,N_3985);
and U7678 (N_7678,N_4493,N_3694);
nand U7679 (N_7679,N_3354,N_5269);
nor U7680 (N_7680,N_4607,N_5689);
xor U7681 (N_7681,N_3235,N_3314);
nand U7682 (N_7682,N_5630,N_5522);
xnor U7683 (N_7683,N_5604,N_4330);
xor U7684 (N_7684,N_3897,N_3628);
nor U7685 (N_7685,N_3052,N_4122);
nor U7686 (N_7686,N_4705,N_3062);
xnor U7687 (N_7687,N_5792,N_3272);
nor U7688 (N_7688,N_3705,N_5604);
and U7689 (N_7689,N_4914,N_3101);
nor U7690 (N_7690,N_4749,N_4614);
and U7691 (N_7691,N_3782,N_5529);
and U7692 (N_7692,N_4144,N_4423);
or U7693 (N_7693,N_4186,N_5143);
nor U7694 (N_7694,N_5973,N_4323);
or U7695 (N_7695,N_3372,N_4853);
nand U7696 (N_7696,N_5363,N_4162);
and U7697 (N_7697,N_5360,N_4904);
nor U7698 (N_7698,N_4355,N_3640);
nand U7699 (N_7699,N_5298,N_5831);
xor U7700 (N_7700,N_3803,N_3432);
nand U7701 (N_7701,N_4330,N_4464);
or U7702 (N_7702,N_4482,N_3811);
or U7703 (N_7703,N_5453,N_4991);
nand U7704 (N_7704,N_3668,N_3127);
and U7705 (N_7705,N_4378,N_4417);
and U7706 (N_7706,N_4657,N_3238);
and U7707 (N_7707,N_4582,N_3078);
or U7708 (N_7708,N_3792,N_4929);
nand U7709 (N_7709,N_5415,N_5150);
or U7710 (N_7710,N_4747,N_5765);
xor U7711 (N_7711,N_3038,N_3988);
xnor U7712 (N_7712,N_4108,N_4387);
or U7713 (N_7713,N_3759,N_5429);
nand U7714 (N_7714,N_3950,N_3911);
nor U7715 (N_7715,N_3517,N_5318);
and U7716 (N_7716,N_3705,N_3016);
and U7717 (N_7717,N_3788,N_5238);
or U7718 (N_7718,N_3910,N_4351);
nand U7719 (N_7719,N_3484,N_3836);
xnor U7720 (N_7720,N_5730,N_3311);
nor U7721 (N_7721,N_5464,N_5313);
nand U7722 (N_7722,N_3570,N_4832);
or U7723 (N_7723,N_4073,N_4231);
xnor U7724 (N_7724,N_5422,N_3686);
nor U7725 (N_7725,N_3097,N_3548);
or U7726 (N_7726,N_3092,N_3228);
or U7727 (N_7727,N_3318,N_4670);
nor U7728 (N_7728,N_4609,N_5879);
nand U7729 (N_7729,N_3008,N_5995);
or U7730 (N_7730,N_4215,N_4747);
and U7731 (N_7731,N_5157,N_4431);
nand U7732 (N_7732,N_4308,N_5637);
nand U7733 (N_7733,N_3179,N_3442);
nand U7734 (N_7734,N_4433,N_4357);
and U7735 (N_7735,N_3421,N_4739);
or U7736 (N_7736,N_3341,N_4689);
xor U7737 (N_7737,N_4753,N_3679);
or U7738 (N_7738,N_4129,N_5670);
and U7739 (N_7739,N_4594,N_4804);
nor U7740 (N_7740,N_3179,N_5913);
nor U7741 (N_7741,N_5890,N_5959);
nor U7742 (N_7742,N_4290,N_3550);
nor U7743 (N_7743,N_3200,N_3331);
xnor U7744 (N_7744,N_5804,N_5296);
nor U7745 (N_7745,N_5568,N_4497);
or U7746 (N_7746,N_3135,N_4063);
nor U7747 (N_7747,N_4404,N_4034);
nor U7748 (N_7748,N_5084,N_4425);
and U7749 (N_7749,N_5812,N_5311);
or U7750 (N_7750,N_3104,N_4547);
nor U7751 (N_7751,N_3658,N_5031);
and U7752 (N_7752,N_4973,N_5703);
or U7753 (N_7753,N_4465,N_3875);
nand U7754 (N_7754,N_5251,N_3948);
and U7755 (N_7755,N_3884,N_3940);
and U7756 (N_7756,N_3567,N_5361);
and U7757 (N_7757,N_5988,N_4060);
or U7758 (N_7758,N_5610,N_3641);
nor U7759 (N_7759,N_4548,N_5632);
nor U7760 (N_7760,N_3332,N_3553);
nor U7761 (N_7761,N_4437,N_3698);
and U7762 (N_7762,N_4532,N_5792);
xor U7763 (N_7763,N_4783,N_3038);
nand U7764 (N_7764,N_5533,N_4147);
nand U7765 (N_7765,N_3610,N_3769);
nor U7766 (N_7766,N_5992,N_3495);
or U7767 (N_7767,N_3401,N_3640);
xor U7768 (N_7768,N_3432,N_4363);
nor U7769 (N_7769,N_4413,N_5636);
xnor U7770 (N_7770,N_5598,N_4169);
nand U7771 (N_7771,N_5321,N_5495);
nand U7772 (N_7772,N_3036,N_3916);
nand U7773 (N_7773,N_4710,N_3945);
nor U7774 (N_7774,N_3401,N_3583);
nand U7775 (N_7775,N_4170,N_3409);
nor U7776 (N_7776,N_3733,N_3495);
nor U7777 (N_7777,N_3903,N_3103);
and U7778 (N_7778,N_5652,N_4126);
or U7779 (N_7779,N_4635,N_4960);
or U7780 (N_7780,N_3629,N_5997);
xor U7781 (N_7781,N_5313,N_5195);
xnor U7782 (N_7782,N_3800,N_4392);
xor U7783 (N_7783,N_4241,N_5201);
or U7784 (N_7784,N_4916,N_4079);
nor U7785 (N_7785,N_5953,N_3145);
nor U7786 (N_7786,N_4267,N_4059);
or U7787 (N_7787,N_4120,N_3113);
nor U7788 (N_7788,N_3978,N_3554);
and U7789 (N_7789,N_5834,N_5688);
nor U7790 (N_7790,N_5265,N_5305);
nand U7791 (N_7791,N_5935,N_4192);
nor U7792 (N_7792,N_4798,N_3630);
or U7793 (N_7793,N_4681,N_5692);
nor U7794 (N_7794,N_5695,N_5150);
and U7795 (N_7795,N_3067,N_3468);
xnor U7796 (N_7796,N_3147,N_3485);
xnor U7797 (N_7797,N_3745,N_5953);
nand U7798 (N_7798,N_3603,N_5607);
or U7799 (N_7799,N_3120,N_4002);
nand U7800 (N_7800,N_5692,N_3750);
and U7801 (N_7801,N_3736,N_4608);
nand U7802 (N_7802,N_4169,N_3022);
xor U7803 (N_7803,N_3099,N_5849);
xnor U7804 (N_7804,N_4150,N_4646);
nor U7805 (N_7805,N_4322,N_5633);
or U7806 (N_7806,N_4748,N_5439);
and U7807 (N_7807,N_3335,N_4069);
nand U7808 (N_7808,N_3715,N_5080);
and U7809 (N_7809,N_5221,N_3196);
nand U7810 (N_7810,N_3756,N_5260);
or U7811 (N_7811,N_5598,N_4479);
nand U7812 (N_7812,N_3574,N_3917);
or U7813 (N_7813,N_5371,N_5595);
nor U7814 (N_7814,N_3986,N_5237);
or U7815 (N_7815,N_3267,N_3561);
nor U7816 (N_7816,N_3801,N_5629);
nand U7817 (N_7817,N_3597,N_5404);
nor U7818 (N_7818,N_5695,N_5740);
xor U7819 (N_7819,N_3219,N_4346);
nor U7820 (N_7820,N_3961,N_4138);
nor U7821 (N_7821,N_5388,N_4323);
and U7822 (N_7822,N_4680,N_3957);
nor U7823 (N_7823,N_5073,N_4817);
xor U7824 (N_7824,N_3404,N_4856);
xor U7825 (N_7825,N_4872,N_5641);
and U7826 (N_7826,N_4366,N_3735);
and U7827 (N_7827,N_5383,N_4172);
or U7828 (N_7828,N_5734,N_4312);
nand U7829 (N_7829,N_4708,N_4929);
nand U7830 (N_7830,N_3698,N_3201);
xor U7831 (N_7831,N_4346,N_4282);
nor U7832 (N_7832,N_5069,N_5798);
nand U7833 (N_7833,N_4758,N_5678);
nand U7834 (N_7834,N_5450,N_3587);
nor U7835 (N_7835,N_4104,N_4600);
xnor U7836 (N_7836,N_3564,N_3146);
nand U7837 (N_7837,N_5184,N_3667);
or U7838 (N_7838,N_3476,N_4696);
xnor U7839 (N_7839,N_3312,N_3381);
or U7840 (N_7840,N_4784,N_5190);
or U7841 (N_7841,N_5534,N_4289);
xnor U7842 (N_7842,N_3941,N_4341);
nor U7843 (N_7843,N_5419,N_5098);
and U7844 (N_7844,N_5904,N_3229);
nor U7845 (N_7845,N_3118,N_3092);
or U7846 (N_7846,N_4033,N_5750);
nor U7847 (N_7847,N_5656,N_4145);
nand U7848 (N_7848,N_3984,N_3548);
or U7849 (N_7849,N_4889,N_5739);
and U7850 (N_7850,N_4988,N_3054);
and U7851 (N_7851,N_3823,N_3266);
and U7852 (N_7852,N_4110,N_4756);
nand U7853 (N_7853,N_4099,N_5299);
xnor U7854 (N_7854,N_5630,N_5801);
or U7855 (N_7855,N_4925,N_3739);
nand U7856 (N_7856,N_5608,N_4596);
xor U7857 (N_7857,N_4854,N_5622);
or U7858 (N_7858,N_4404,N_5733);
nand U7859 (N_7859,N_5674,N_3267);
xor U7860 (N_7860,N_3206,N_3798);
nor U7861 (N_7861,N_3561,N_3896);
nand U7862 (N_7862,N_5353,N_3992);
nand U7863 (N_7863,N_3690,N_4434);
xor U7864 (N_7864,N_4764,N_3206);
nand U7865 (N_7865,N_3301,N_3964);
xnor U7866 (N_7866,N_5212,N_3092);
nand U7867 (N_7867,N_4838,N_4794);
and U7868 (N_7868,N_5643,N_5001);
or U7869 (N_7869,N_5202,N_3948);
xnor U7870 (N_7870,N_5715,N_5843);
and U7871 (N_7871,N_5698,N_5105);
and U7872 (N_7872,N_5477,N_4156);
and U7873 (N_7873,N_3315,N_5597);
nor U7874 (N_7874,N_3525,N_4624);
or U7875 (N_7875,N_3649,N_3079);
and U7876 (N_7876,N_5609,N_4088);
or U7877 (N_7877,N_3507,N_5356);
and U7878 (N_7878,N_5404,N_5086);
xor U7879 (N_7879,N_3778,N_4919);
or U7880 (N_7880,N_4450,N_4053);
nand U7881 (N_7881,N_5214,N_4479);
and U7882 (N_7882,N_3584,N_3735);
and U7883 (N_7883,N_4567,N_5825);
xor U7884 (N_7884,N_3722,N_5417);
or U7885 (N_7885,N_5341,N_4813);
nor U7886 (N_7886,N_5248,N_4028);
xor U7887 (N_7887,N_5630,N_4268);
and U7888 (N_7888,N_3738,N_3558);
nand U7889 (N_7889,N_4915,N_4896);
xor U7890 (N_7890,N_3180,N_5367);
or U7891 (N_7891,N_4975,N_4798);
nor U7892 (N_7892,N_5156,N_3649);
and U7893 (N_7893,N_3555,N_4709);
or U7894 (N_7894,N_4308,N_4608);
or U7895 (N_7895,N_4145,N_3636);
nand U7896 (N_7896,N_5295,N_5011);
nand U7897 (N_7897,N_4867,N_5977);
xor U7898 (N_7898,N_4313,N_3817);
and U7899 (N_7899,N_4202,N_3628);
nand U7900 (N_7900,N_4097,N_5867);
nor U7901 (N_7901,N_3438,N_5481);
nand U7902 (N_7902,N_3477,N_3704);
and U7903 (N_7903,N_4064,N_3284);
nand U7904 (N_7904,N_3625,N_3800);
and U7905 (N_7905,N_3435,N_3674);
nor U7906 (N_7906,N_4042,N_3385);
or U7907 (N_7907,N_4053,N_4072);
or U7908 (N_7908,N_3467,N_4247);
nand U7909 (N_7909,N_5562,N_3183);
nor U7910 (N_7910,N_4719,N_4516);
nor U7911 (N_7911,N_5537,N_4522);
nor U7912 (N_7912,N_4835,N_5422);
nand U7913 (N_7913,N_3049,N_5057);
or U7914 (N_7914,N_4907,N_5408);
or U7915 (N_7915,N_4185,N_5880);
nand U7916 (N_7916,N_5091,N_5254);
xor U7917 (N_7917,N_4577,N_5394);
or U7918 (N_7918,N_5705,N_4985);
and U7919 (N_7919,N_4191,N_3683);
and U7920 (N_7920,N_3766,N_4266);
or U7921 (N_7921,N_4362,N_5811);
nand U7922 (N_7922,N_3655,N_4076);
nand U7923 (N_7923,N_3431,N_5863);
or U7924 (N_7924,N_3994,N_3378);
or U7925 (N_7925,N_3653,N_5986);
nor U7926 (N_7926,N_5191,N_4820);
nand U7927 (N_7927,N_5467,N_3999);
nor U7928 (N_7928,N_5001,N_4379);
xnor U7929 (N_7929,N_5401,N_4329);
nand U7930 (N_7930,N_4828,N_4565);
nor U7931 (N_7931,N_4540,N_5822);
and U7932 (N_7932,N_5827,N_3872);
and U7933 (N_7933,N_5223,N_5999);
xnor U7934 (N_7934,N_3890,N_4495);
xor U7935 (N_7935,N_4675,N_5837);
nor U7936 (N_7936,N_3863,N_3901);
nand U7937 (N_7937,N_3319,N_3696);
nand U7938 (N_7938,N_4994,N_4159);
nand U7939 (N_7939,N_5787,N_4099);
xnor U7940 (N_7940,N_4591,N_5323);
nand U7941 (N_7941,N_4881,N_3851);
nand U7942 (N_7942,N_4883,N_3167);
nand U7943 (N_7943,N_4637,N_3065);
or U7944 (N_7944,N_4595,N_3215);
xnor U7945 (N_7945,N_3989,N_5164);
nand U7946 (N_7946,N_4892,N_5972);
nand U7947 (N_7947,N_4643,N_4232);
xor U7948 (N_7948,N_3890,N_5149);
nor U7949 (N_7949,N_3413,N_3870);
nor U7950 (N_7950,N_5672,N_4684);
xor U7951 (N_7951,N_4921,N_3691);
xnor U7952 (N_7952,N_5907,N_5704);
xnor U7953 (N_7953,N_4876,N_3132);
and U7954 (N_7954,N_3288,N_3243);
nand U7955 (N_7955,N_5995,N_4377);
and U7956 (N_7956,N_3695,N_5442);
or U7957 (N_7957,N_4927,N_4383);
nand U7958 (N_7958,N_4573,N_4630);
or U7959 (N_7959,N_4885,N_5513);
or U7960 (N_7960,N_4569,N_3235);
nor U7961 (N_7961,N_5841,N_3949);
or U7962 (N_7962,N_3067,N_5369);
xor U7963 (N_7963,N_5456,N_5936);
and U7964 (N_7964,N_4201,N_4813);
xnor U7965 (N_7965,N_5798,N_4992);
xor U7966 (N_7966,N_5554,N_3388);
or U7967 (N_7967,N_5896,N_5621);
or U7968 (N_7968,N_4837,N_5085);
nand U7969 (N_7969,N_5778,N_5726);
nor U7970 (N_7970,N_4494,N_5549);
nand U7971 (N_7971,N_3542,N_5221);
nor U7972 (N_7972,N_5128,N_5188);
nand U7973 (N_7973,N_5062,N_3270);
and U7974 (N_7974,N_4802,N_3380);
nor U7975 (N_7975,N_5170,N_4264);
and U7976 (N_7976,N_4529,N_3773);
xor U7977 (N_7977,N_4827,N_4466);
nor U7978 (N_7978,N_4467,N_3428);
nor U7979 (N_7979,N_5865,N_5440);
nand U7980 (N_7980,N_3622,N_5944);
or U7981 (N_7981,N_5284,N_3651);
or U7982 (N_7982,N_5219,N_4538);
nor U7983 (N_7983,N_3008,N_3070);
or U7984 (N_7984,N_4837,N_3165);
xnor U7985 (N_7985,N_3739,N_3918);
xor U7986 (N_7986,N_5623,N_3429);
nor U7987 (N_7987,N_5730,N_5246);
nand U7988 (N_7988,N_4897,N_3505);
nand U7989 (N_7989,N_3226,N_4602);
xor U7990 (N_7990,N_3960,N_3057);
or U7991 (N_7991,N_5542,N_3383);
nand U7992 (N_7992,N_3459,N_3363);
xor U7993 (N_7993,N_4143,N_5409);
or U7994 (N_7994,N_4101,N_3138);
nor U7995 (N_7995,N_4488,N_5259);
and U7996 (N_7996,N_3621,N_4957);
nor U7997 (N_7997,N_5370,N_4265);
or U7998 (N_7998,N_5981,N_3477);
and U7999 (N_7999,N_4114,N_5608);
xnor U8000 (N_8000,N_3784,N_4820);
and U8001 (N_8001,N_5376,N_4867);
and U8002 (N_8002,N_5326,N_3416);
or U8003 (N_8003,N_5156,N_5033);
and U8004 (N_8004,N_5018,N_4317);
nand U8005 (N_8005,N_4621,N_4042);
nor U8006 (N_8006,N_5868,N_4119);
and U8007 (N_8007,N_4212,N_5892);
xor U8008 (N_8008,N_5842,N_4174);
xor U8009 (N_8009,N_3235,N_5779);
nor U8010 (N_8010,N_3185,N_4644);
xor U8011 (N_8011,N_5192,N_3869);
nand U8012 (N_8012,N_3671,N_4091);
or U8013 (N_8013,N_5913,N_3739);
nand U8014 (N_8014,N_4985,N_4956);
nor U8015 (N_8015,N_5938,N_5269);
and U8016 (N_8016,N_5251,N_5860);
nor U8017 (N_8017,N_5443,N_5155);
xor U8018 (N_8018,N_5197,N_5465);
and U8019 (N_8019,N_4088,N_4224);
or U8020 (N_8020,N_5718,N_5451);
nor U8021 (N_8021,N_3619,N_5548);
nand U8022 (N_8022,N_5260,N_4617);
nor U8023 (N_8023,N_4847,N_3069);
nand U8024 (N_8024,N_5432,N_3941);
nor U8025 (N_8025,N_4755,N_5092);
or U8026 (N_8026,N_3660,N_4689);
nand U8027 (N_8027,N_3664,N_5292);
or U8028 (N_8028,N_5138,N_3819);
or U8029 (N_8029,N_4490,N_3133);
and U8030 (N_8030,N_4536,N_3604);
nor U8031 (N_8031,N_4685,N_4833);
nand U8032 (N_8032,N_5707,N_4668);
or U8033 (N_8033,N_5138,N_4540);
nor U8034 (N_8034,N_5172,N_3476);
xnor U8035 (N_8035,N_4474,N_3082);
xor U8036 (N_8036,N_5756,N_3572);
and U8037 (N_8037,N_3759,N_4222);
nor U8038 (N_8038,N_5527,N_4636);
or U8039 (N_8039,N_4547,N_3323);
xnor U8040 (N_8040,N_3365,N_5119);
nand U8041 (N_8041,N_4740,N_3228);
xnor U8042 (N_8042,N_3179,N_3276);
nand U8043 (N_8043,N_3340,N_3200);
and U8044 (N_8044,N_5865,N_4705);
nand U8045 (N_8045,N_5406,N_4942);
nor U8046 (N_8046,N_5877,N_3585);
nor U8047 (N_8047,N_4894,N_4228);
xor U8048 (N_8048,N_4554,N_3879);
nand U8049 (N_8049,N_4659,N_5455);
nor U8050 (N_8050,N_4688,N_3755);
and U8051 (N_8051,N_4041,N_3839);
nor U8052 (N_8052,N_4042,N_5036);
nand U8053 (N_8053,N_3127,N_4887);
nand U8054 (N_8054,N_4117,N_5542);
nand U8055 (N_8055,N_3603,N_4163);
or U8056 (N_8056,N_3284,N_4486);
nor U8057 (N_8057,N_3614,N_5412);
or U8058 (N_8058,N_4967,N_5040);
nor U8059 (N_8059,N_3564,N_3618);
xnor U8060 (N_8060,N_4842,N_4425);
xnor U8061 (N_8061,N_3716,N_4964);
and U8062 (N_8062,N_3479,N_5443);
and U8063 (N_8063,N_5621,N_3520);
and U8064 (N_8064,N_4665,N_3654);
xor U8065 (N_8065,N_4972,N_5588);
and U8066 (N_8066,N_4360,N_3056);
xnor U8067 (N_8067,N_4611,N_5604);
nor U8068 (N_8068,N_3019,N_3434);
and U8069 (N_8069,N_5655,N_5123);
nor U8070 (N_8070,N_3277,N_4994);
xor U8071 (N_8071,N_5622,N_4722);
xnor U8072 (N_8072,N_3550,N_5487);
xnor U8073 (N_8073,N_5148,N_5589);
xor U8074 (N_8074,N_4306,N_5039);
and U8075 (N_8075,N_3040,N_3976);
nor U8076 (N_8076,N_3393,N_3368);
xor U8077 (N_8077,N_5112,N_5735);
nor U8078 (N_8078,N_5809,N_4386);
nor U8079 (N_8079,N_5797,N_3209);
or U8080 (N_8080,N_3611,N_3084);
nand U8081 (N_8081,N_3444,N_5484);
nor U8082 (N_8082,N_3125,N_4673);
and U8083 (N_8083,N_4833,N_4188);
xnor U8084 (N_8084,N_4227,N_4304);
and U8085 (N_8085,N_4501,N_4473);
nand U8086 (N_8086,N_4773,N_3407);
or U8087 (N_8087,N_5219,N_3251);
and U8088 (N_8088,N_4247,N_4249);
nand U8089 (N_8089,N_4434,N_5903);
and U8090 (N_8090,N_3064,N_5342);
nand U8091 (N_8091,N_3103,N_4467);
and U8092 (N_8092,N_3206,N_3593);
nand U8093 (N_8093,N_3862,N_4706);
and U8094 (N_8094,N_4595,N_3677);
nand U8095 (N_8095,N_5695,N_4414);
or U8096 (N_8096,N_4779,N_4398);
nor U8097 (N_8097,N_4407,N_5460);
xnor U8098 (N_8098,N_5684,N_4098);
nand U8099 (N_8099,N_4213,N_4980);
or U8100 (N_8100,N_5142,N_4694);
nor U8101 (N_8101,N_4351,N_5229);
or U8102 (N_8102,N_4756,N_4735);
nand U8103 (N_8103,N_4939,N_5388);
xor U8104 (N_8104,N_5924,N_5897);
and U8105 (N_8105,N_4986,N_5493);
nand U8106 (N_8106,N_3482,N_4157);
xnor U8107 (N_8107,N_4705,N_5749);
and U8108 (N_8108,N_4373,N_5114);
xor U8109 (N_8109,N_5820,N_3352);
nand U8110 (N_8110,N_4358,N_4655);
and U8111 (N_8111,N_3823,N_5054);
or U8112 (N_8112,N_5164,N_5043);
or U8113 (N_8113,N_5538,N_4277);
nor U8114 (N_8114,N_4712,N_5397);
or U8115 (N_8115,N_3980,N_4798);
xnor U8116 (N_8116,N_4971,N_3941);
xnor U8117 (N_8117,N_5767,N_3543);
nor U8118 (N_8118,N_5320,N_3004);
nor U8119 (N_8119,N_5628,N_5220);
and U8120 (N_8120,N_5549,N_4282);
nand U8121 (N_8121,N_4450,N_4141);
and U8122 (N_8122,N_4088,N_4511);
xor U8123 (N_8123,N_4890,N_4523);
and U8124 (N_8124,N_5577,N_3867);
nand U8125 (N_8125,N_5516,N_3293);
and U8126 (N_8126,N_5551,N_5893);
nand U8127 (N_8127,N_3186,N_5421);
xnor U8128 (N_8128,N_5629,N_3520);
nor U8129 (N_8129,N_5471,N_4275);
nand U8130 (N_8130,N_5416,N_3234);
nor U8131 (N_8131,N_5473,N_5347);
or U8132 (N_8132,N_5420,N_5184);
nor U8133 (N_8133,N_4051,N_5752);
or U8134 (N_8134,N_5468,N_4738);
and U8135 (N_8135,N_3662,N_5792);
nand U8136 (N_8136,N_5394,N_3230);
and U8137 (N_8137,N_3927,N_4369);
and U8138 (N_8138,N_4786,N_5469);
and U8139 (N_8139,N_4588,N_3630);
xor U8140 (N_8140,N_4136,N_5555);
nor U8141 (N_8141,N_3350,N_4814);
and U8142 (N_8142,N_4379,N_3106);
nand U8143 (N_8143,N_4466,N_4095);
nor U8144 (N_8144,N_4585,N_4354);
and U8145 (N_8145,N_4933,N_3072);
nand U8146 (N_8146,N_3075,N_4518);
or U8147 (N_8147,N_3594,N_4487);
xnor U8148 (N_8148,N_3466,N_4684);
nor U8149 (N_8149,N_5842,N_5573);
nor U8150 (N_8150,N_5732,N_3994);
xor U8151 (N_8151,N_5039,N_5186);
nand U8152 (N_8152,N_5430,N_4519);
nor U8153 (N_8153,N_4830,N_5378);
nor U8154 (N_8154,N_3493,N_4460);
nor U8155 (N_8155,N_4026,N_3292);
nand U8156 (N_8156,N_5748,N_4522);
nand U8157 (N_8157,N_4918,N_5724);
xnor U8158 (N_8158,N_3240,N_5883);
or U8159 (N_8159,N_3687,N_4261);
nand U8160 (N_8160,N_4903,N_3017);
xnor U8161 (N_8161,N_3980,N_5647);
nand U8162 (N_8162,N_3706,N_3082);
and U8163 (N_8163,N_4078,N_4139);
and U8164 (N_8164,N_5183,N_3692);
nand U8165 (N_8165,N_4633,N_5743);
or U8166 (N_8166,N_4110,N_5483);
or U8167 (N_8167,N_3886,N_3592);
or U8168 (N_8168,N_4619,N_3627);
xor U8169 (N_8169,N_3977,N_5842);
xnor U8170 (N_8170,N_4054,N_3686);
and U8171 (N_8171,N_5886,N_5323);
nand U8172 (N_8172,N_4693,N_3661);
xnor U8173 (N_8173,N_3857,N_4430);
and U8174 (N_8174,N_3666,N_3401);
nand U8175 (N_8175,N_3540,N_5196);
nand U8176 (N_8176,N_5260,N_4705);
and U8177 (N_8177,N_5938,N_5020);
or U8178 (N_8178,N_3747,N_5999);
and U8179 (N_8179,N_4007,N_5680);
nor U8180 (N_8180,N_5309,N_3779);
xor U8181 (N_8181,N_5202,N_4450);
and U8182 (N_8182,N_3035,N_4417);
and U8183 (N_8183,N_4160,N_4013);
nand U8184 (N_8184,N_5632,N_3718);
xor U8185 (N_8185,N_3045,N_5234);
nor U8186 (N_8186,N_4606,N_3627);
nand U8187 (N_8187,N_3773,N_5490);
nand U8188 (N_8188,N_4927,N_4425);
nand U8189 (N_8189,N_5344,N_4235);
or U8190 (N_8190,N_3436,N_3639);
nand U8191 (N_8191,N_5130,N_4481);
nand U8192 (N_8192,N_3899,N_5280);
or U8193 (N_8193,N_4684,N_5214);
nor U8194 (N_8194,N_3177,N_5998);
xnor U8195 (N_8195,N_3999,N_5334);
or U8196 (N_8196,N_4621,N_4270);
nand U8197 (N_8197,N_4085,N_5316);
or U8198 (N_8198,N_3598,N_4832);
nor U8199 (N_8199,N_4675,N_5317);
or U8200 (N_8200,N_5967,N_3981);
or U8201 (N_8201,N_3267,N_5380);
or U8202 (N_8202,N_3816,N_3887);
and U8203 (N_8203,N_4051,N_3463);
xor U8204 (N_8204,N_5100,N_5600);
or U8205 (N_8205,N_4188,N_5591);
xnor U8206 (N_8206,N_5733,N_5032);
xnor U8207 (N_8207,N_3083,N_3209);
or U8208 (N_8208,N_5059,N_3771);
nor U8209 (N_8209,N_4873,N_5066);
xor U8210 (N_8210,N_3242,N_3138);
or U8211 (N_8211,N_3935,N_4048);
xor U8212 (N_8212,N_3463,N_5848);
xor U8213 (N_8213,N_4261,N_4076);
and U8214 (N_8214,N_3558,N_3598);
and U8215 (N_8215,N_3199,N_3914);
nor U8216 (N_8216,N_4250,N_5828);
nand U8217 (N_8217,N_5862,N_3491);
or U8218 (N_8218,N_4921,N_3767);
nor U8219 (N_8219,N_4105,N_4666);
nor U8220 (N_8220,N_5978,N_5131);
or U8221 (N_8221,N_5714,N_5616);
and U8222 (N_8222,N_3849,N_5946);
nand U8223 (N_8223,N_4728,N_3931);
xor U8224 (N_8224,N_3712,N_5683);
or U8225 (N_8225,N_3075,N_4616);
nand U8226 (N_8226,N_5689,N_3839);
xor U8227 (N_8227,N_4254,N_3959);
xor U8228 (N_8228,N_4682,N_5896);
or U8229 (N_8229,N_5386,N_3749);
xor U8230 (N_8230,N_3080,N_5415);
xnor U8231 (N_8231,N_3961,N_4131);
nand U8232 (N_8232,N_5281,N_3081);
nor U8233 (N_8233,N_5142,N_5086);
nand U8234 (N_8234,N_5196,N_5204);
or U8235 (N_8235,N_3033,N_3721);
nand U8236 (N_8236,N_3524,N_5087);
and U8237 (N_8237,N_3890,N_3938);
nand U8238 (N_8238,N_3158,N_5310);
and U8239 (N_8239,N_3258,N_4653);
nor U8240 (N_8240,N_3289,N_4853);
xnor U8241 (N_8241,N_4242,N_4139);
nand U8242 (N_8242,N_4475,N_3514);
or U8243 (N_8243,N_5290,N_3012);
xnor U8244 (N_8244,N_5914,N_5427);
or U8245 (N_8245,N_4889,N_3801);
and U8246 (N_8246,N_5761,N_4993);
xor U8247 (N_8247,N_4782,N_3371);
and U8248 (N_8248,N_4552,N_5650);
and U8249 (N_8249,N_4704,N_4965);
or U8250 (N_8250,N_4864,N_5193);
and U8251 (N_8251,N_5365,N_5993);
nor U8252 (N_8252,N_4947,N_3940);
and U8253 (N_8253,N_4524,N_3907);
xnor U8254 (N_8254,N_5535,N_5194);
nand U8255 (N_8255,N_4122,N_4946);
nor U8256 (N_8256,N_5330,N_3339);
xor U8257 (N_8257,N_4126,N_4736);
and U8258 (N_8258,N_4164,N_3131);
and U8259 (N_8259,N_4527,N_5102);
nor U8260 (N_8260,N_3869,N_5359);
and U8261 (N_8261,N_5194,N_5910);
nand U8262 (N_8262,N_3287,N_4381);
nor U8263 (N_8263,N_3845,N_4560);
and U8264 (N_8264,N_3770,N_4742);
or U8265 (N_8265,N_4824,N_4274);
or U8266 (N_8266,N_3313,N_4451);
nor U8267 (N_8267,N_4286,N_4672);
nand U8268 (N_8268,N_5749,N_3274);
nor U8269 (N_8269,N_5370,N_5166);
and U8270 (N_8270,N_3376,N_5408);
or U8271 (N_8271,N_5431,N_5463);
nand U8272 (N_8272,N_3301,N_5044);
or U8273 (N_8273,N_3634,N_4153);
and U8274 (N_8274,N_3655,N_3595);
nand U8275 (N_8275,N_5168,N_4222);
and U8276 (N_8276,N_3970,N_4016);
xor U8277 (N_8277,N_4906,N_5883);
and U8278 (N_8278,N_4599,N_3626);
nor U8279 (N_8279,N_4276,N_5980);
or U8280 (N_8280,N_5135,N_3400);
and U8281 (N_8281,N_4393,N_3377);
or U8282 (N_8282,N_5743,N_4398);
xor U8283 (N_8283,N_3569,N_5224);
nand U8284 (N_8284,N_4215,N_3464);
xor U8285 (N_8285,N_5157,N_4808);
xor U8286 (N_8286,N_3431,N_5771);
and U8287 (N_8287,N_4889,N_5491);
and U8288 (N_8288,N_3475,N_3415);
and U8289 (N_8289,N_3875,N_4411);
xnor U8290 (N_8290,N_5436,N_3004);
and U8291 (N_8291,N_4460,N_4517);
nand U8292 (N_8292,N_5190,N_5429);
xor U8293 (N_8293,N_4626,N_3513);
xor U8294 (N_8294,N_3569,N_4372);
nor U8295 (N_8295,N_3793,N_3819);
xor U8296 (N_8296,N_3060,N_3895);
and U8297 (N_8297,N_3291,N_4622);
or U8298 (N_8298,N_3878,N_3445);
nor U8299 (N_8299,N_3141,N_3360);
xor U8300 (N_8300,N_3876,N_5039);
xor U8301 (N_8301,N_4955,N_3121);
or U8302 (N_8302,N_3187,N_5812);
xor U8303 (N_8303,N_3297,N_4278);
nor U8304 (N_8304,N_5786,N_3049);
and U8305 (N_8305,N_5869,N_4855);
and U8306 (N_8306,N_5547,N_3391);
xor U8307 (N_8307,N_3704,N_3261);
or U8308 (N_8308,N_4686,N_4744);
nor U8309 (N_8309,N_3918,N_5080);
nand U8310 (N_8310,N_3759,N_4710);
or U8311 (N_8311,N_4772,N_3596);
xnor U8312 (N_8312,N_3960,N_4306);
or U8313 (N_8313,N_5522,N_5434);
and U8314 (N_8314,N_4981,N_3781);
nand U8315 (N_8315,N_5335,N_5328);
xor U8316 (N_8316,N_5295,N_5957);
or U8317 (N_8317,N_3556,N_5032);
nand U8318 (N_8318,N_5033,N_5929);
nand U8319 (N_8319,N_3474,N_5969);
nor U8320 (N_8320,N_4105,N_5363);
nand U8321 (N_8321,N_5944,N_5310);
xor U8322 (N_8322,N_4233,N_3574);
xnor U8323 (N_8323,N_5162,N_4796);
and U8324 (N_8324,N_4313,N_4707);
nand U8325 (N_8325,N_3114,N_4922);
nor U8326 (N_8326,N_5426,N_5701);
nand U8327 (N_8327,N_5286,N_5791);
or U8328 (N_8328,N_3801,N_3240);
nand U8329 (N_8329,N_3685,N_5727);
nor U8330 (N_8330,N_4964,N_3041);
nand U8331 (N_8331,N_5331,N_5820);
xor U8332 (N_8332,N_4239,N_3866);
xor U8333 (N_8333,N_5801,N_3427);
xnor U8334 (N_8334,N_4730,N_3530);
nand U8335 (N_8335,N_5879,N_5208);
xnor U8336 (N_8336,N_3996,N_5941);
and U8337 (N_8337,N_3273,N_4585);
and U8338 (N_8338,N_5722,N_3973);
xor U8339 (N_8339,N_5948,N_3149);
or U8340 (N_8340,N_5072,N_4012);
or U8341 (N_8341,N_5215,N_4128);
or U8342 (N_8342,N_5509,N_3240);
xor U8343 (N_8343,N_3755,N_3471);
and U8344 (N_8344,N_4992,N_4286);
nor U8345 (N_8345,N_3390,N_4681);
nand U8346 (N_8346,N_4070,N_4861);
nor U8347 (N_8347,N_3178,N_3788);
nor U8348 (N_8348,N_3941,N_4780);
nor U8349 (N_8349,N_3773,N_3005);
xor U8350 (N_8350,N_4941,N_5585);
nor U8351 (N_8351,N_3357,N_4364);
or U8352 (N_8352,N_5452,N_5052);
xnor U8353 (N_8353,N_5759,N_3772);
xnor U8354 (N_8354,N_5832,N_5930);
nand U8355 (N_8355,N_3054,N_4072);
and U8356 (N_8356,N_5772,N_3632);
or U8357 (N_8357,N_5585,N_5321);
or U8358 (N_8358,N_4675,N_4299);
or U8359 (N_8359,N_4935,N_5214);
xnor U8360 (N_8360,N_3544,N_3937);
nor U8361 (N_8361,N_3586,N_4902);
xor U8362 (N_8362,N_4559,N_3827);
or U8363 (N_8363,N_3324,N_3816);
or U8364 (N_8364,N_3679,N_3869);
and U8365 (N_8365,N_4299,N_3982);
nand U8366 (N_8366,N_4710,N_4435);
nand U8367 (N_8367,N_5594,N_3561);
xnor U8368 (N_8368,N_3974,N_5235);
or U8369 (N_8369,N_5545,N_4514);
nor U8370 (N_8370,N_5453,N_4711);
or U8371 (N_8371,N_4737,N_4228);
xnor U8372 (N_8372,N_3612,N_4211);
nand U8373 (N_8373,N_5695,N_3875);
nor U8374 (N_8374,N_4958,N_4317);
nand U8375 (N_8375,N_3701,N_3720);
and U8376 (N_8376,N_4348,N_3176);
xnor U8377 (N_8377,N_4352,N_5806);
xnor U8378 (N_8378,N_3182,N_4126);
nor U8379 (N_8379,N_4488,N_5053);
or U8380 (N_8380,N_3361,N_5595);
nor U8381 (N_8381,N_3486,N_4291);
and U8382 (N_8382,N_5297,N_3382);
nand U8383 (N_8383,N_3795,N_3038);
nor U8384 (N_8384,N_4264,N_3753);
xnor U8385 (N_8385,N_4341,N_4041);
xor U8386 (N_8386,N_3668,N_4373);
and U8387 (N_8387,N_5126,N_4794);
xnor U8388 (N_8388,N_5194,N_3788);
and U8389 (N_8389,N_3380,N_3188);
and U8390 (N_8390,N_5521,N_5718);
and U8391 (N_8391,N_4981,N_5007);
or U8392 (N_8392,N_3174,N_3420);
and U8393 (N_8393,N_3584,N_5262);
xnor U8394 (N_8394,N_5234,N_3301);
nand U8395 (N_8395,N_5031,N_5879);
or U8396 (N_8396,N_4901,N_3143);
nor U8397 (N_8397,N_4138,N_4987);
xor U8398 (N_8398,N_4404,N_5820);
xnor U8399 (N_8399,N_3900,N_4546);
or U8400 (N_8400,N_5573,N_3538);
xor U8401 (N_8401,N_4380,N_5747);
xnor U8402 (N_8402,N_5269,N_5322);
or U8403 (N_8403,N_5432,N_4301);
nor U8404 (N_8404,N_3608,N_3585);
nor U8405 (N_8405,N_4115,N_4235);
or U8406 (N_8406,N_3494,N_5695);
or U8407 (N_8407,N_5329,N_4362);
nor U8408 (N_8408,N_5837,N_4125);
nor U8409 (N_8409,N_5568,N_5893);
nand U8410 (N_8410,N_4168,N_3308);
or U8411 (N_8411,N_3410,N_4531);
nand U8412 (N_8412,N_4099,N_4394);
or U8413 (N_8413,N_4205,N_3667);
and U8414 (N_8414,N_4611,N_3334);
xnor U8415 (N_8415,N_4173,N_4433);
nand U8416 (N_8416,N_4218,N_4253);
nand U8417 (N_8417,N_5532,N_5119);
or U8418 (N_8418,N_4144,N_3159);
nor U8419 (N_8419,N_4391,N_4920);
and U8420 (N_8420,N_4855,N_4348);
nor U8421 (N_8421,N_5758,N_3478);
and U8422 (N_8422,N_5030,N_5921);
nor U8423 (N_8423,N_4695,N_5605);
nor U8424 (N_8424,N_4113,N_3058);
xnor U8425 (N_8425,N_3633,N_3530);
or U8426 (N_8426,N_3957,N_3104);
or U8427 (N_8427,N_3144,N_3344);
and U8428 (N_8428,N_4190,N_3345);
nor U8429 (N_8429,N_5926,N_3535);
nand U8430 (N_8430,N_4185,N_5334);
nand U8431 (N_8431,N_3214,N_4648);
and U8432 (N_8432,N_3325,N_4183);
xor U8433 (N_8433,N_4233,N_4531);
xnor U8434 (N_8434,N_4945,N_3233);
nor U8435 (N_8435,N_5499,N_5510);
nand U8436 (N_8436,N_4650,N_3399);
nand U8437 (N_8437,N_5010,N_3093);
nor U8438 (N_8438,N_3268,N_5402);
or U8439 (N_8439,N_3764,N_3449);
and U8440 (N_8440,N_5776,N_4907);
or U8441 (N_8441,N_5094,N_4426);
nor U8442 (N_8442,N_4876,N_3429);
or U8443 (N_8443,N_4139,N_5607);
xnor U8444 (N_8444,N_4338,N_4835);
xnor U8445 (N_8445,N_3666,N_4210);
and U8446 (N_8446,N_5360,N_3522);
xor U8447 (N_8447,N_4628,N_5838);
and U8448 (N_8448,N_5978,N_3620);
nand U8449 (N_8449,N_3415,N_3328);
nor U8450 (N_8450,N_4656,N_3619);
nor U8451 (N_8451,N_5534,N_4833);
nor U8452 (N_8452,N_5238,N_5260);
or U8453 (N_8453,N_4090,N_5398);
nand U8454 (N_8454,N_3987,N_5204);
or U8455 (N_8455,N_5770,N_4903);
or U8456 (N_8456,N_4658,N_5558);
and U8457 (N_8457,N_5028,N_4423);
xnor U8458 (N_8458,N_5868,N_4363);
and U8459 (N_8459,N_4366,N_4933);
nor U8460 (N_8460,N_3730,N_5559);
or U8461 (N_8461,N_3796,N_5000);
nor U8462 (N_8462,N_5956,N_3909);
nor U8463 (N_8463,N_4698,N_3825);
nand U8464 (N_8464,N_3386,N_5386);
nand U8465 (N_8465,N_4806,N_4414);
or U8466 (N_8466,N_3773,N_5013);
and U8467 (N_8467,N_3787,N_5294);
xnor U8468 (N_8468,N_3079,N_4942);
nand U8469 (N_8469,N_3160,N_4586);
or U8470 (N_8470,N_3163,N_4559);
or U8471 (N_8471,N_3413,N_5537);
nand U8472 (N_8472,N_5823,N_5571);
and U8473 (N_8473,N_3987,N_5328);
and U8474 (N_8474,N_3491,N_3157);
xnor U8475 (N_8475,N_5754,N_5882);
nor U8476 (N_8476,N_4337,N_4011);
xnor U8477 (N_8477,N_3468,N_4590);
or U8478 (N_8478,N_4213,N_3758);
or U8479 (N_8479,N_3295,N_5596);
or U8480 (N_8480,N_3392,N_3382);
nand U8481 (N_8481,N_3113,N_3963);
nand U8482 (N_8482,N_5292,N_4277);
xor U8483 (N_8483,N_5170,N_4204);
xnor U8484 (N_8484,N_3171,N_4290);
nor U8485 (N_8485,N_4078,N_3610);
and U8486 (N_8486,N_3357,N_5474);
xor U8487 (N_8487,N_5590,N_5625);
nor U8488 (N_8488,N_4554,N_5948);
nand U8489 (N_8489,N_5143,N_4371);
and U8490 (N_8490,N_4218,N_5539);
or U8491 (N_8491,N_4155,N_5697);
nand U8492 (N_8492,N_3513,N_5166);
nor U8493 (N_8493,N_3755,N_3215);
and U8494 (N_8494,N_3411,N_5273);
and U8495 (N_8495,N_5248,N_4388);
or U8496 (N_8496,N_4275,N_3081);
and U8497 (N_8497,N_5566,N_3740);
and U8498 (N_8498,N_5876,N_5928);
nand U8499 (N_8499,N_5047,N_4138);
and U8500 (N_8500,N_4588,N_4619);
xor U8501 (N_8501,N_4755,N_3834);
nor U8502 (N_8502,N_4200,N_4986);
nand U8503 (N_8503,N_5259,N_4592);
nand U8504 (N_8504,N_5411,N_4740);
or U8505 (N_8505,N_3723,N_5178);
or U8506 (N_8506,N_3739,N_3616);
nor U8507 (N_8507,N_4698,N_5206);
xor U8508 (N_8508,N_4668,N_4085);
and U8509 (N_8509,N_5050,N_5116);
nor U8510 (N_8510,N_3281,N_3287);
xnor U8511 (N_8511,N_5472,N_3595);
or U8512 (N_8512,N_3110,N_5863);
nor U8513 (N_8513,N_5982,N_5072);
nor U8514 (N_8514,N_3811,N_5777);
xor U8515 (N_8515,N_3555,N_3063);
nand U8516 (N_8516,N_3654,N_3388);
and U8517 (N_8517,N_4493,N_5211);
nand U8518 (N_8518,N_4789,N_5326);
xnor U8519 (N_8519,N_4321,N_4937);
nor U8520 (N_8520,N_3737,N_5991);
nor U8521 (N_8521,N_5883,N_5111);
nor U8522 (N_8522,N_4630,N_5708);
xor U8523 (N_8523,N_5308,N_4306);
or U8524 (N_8524,N_4039,N_3324);
xor U8525 (N_8525,N_3242,N_5731);
nor U8526 (N_8526,N_3682,N_3503);
nand U8527 (N_8527,N_5244,N_4633);
xnor U8528 (N_8528,N_5304,N_4067);
nand U8529 (N_8529,N_4813,N_5205);
or U8530 (N_8530,N_5331,N_3335);
and U8531 (N_8531,N_4915,N_5048);
or U8532 (N_8532,N_5618,N_3665);
xnor U8533 (N_8533,N_5512,N_3580);
and U8534 (N_8534,N_5863,N_3091);
and U8535 (N_8535,N_5965,N_5149);
nor U8536 (N_8536,N_5426,N_4552);
and U8537 (N_8537,N_4641,N_4942);
nor U8538 (N_8538,N_5793,N_4571);
nor U8539 (N_8539,N_3681,N_4435);
or U8540 (N_8540,N_4904,N_3354);
or U8541 (N_8541,N_5189,N_5555);
or U8542 (N_8542,N_4314,N_4095);
and U8543 (N_8543,N_4615,N_5685);
xnor U8544 (N_8544,N_4326,N_5536);
xor U8545 (N_8545,N_4544,N_5116);
and U8546 (N_8546,N_5236,N_4582);
or U8547 (N_8547,N_5277,N_4983);
or U8548 (N_8548,N_4750,N_4077);
or U8549 (N_8549,N_5636,N_3999);
or U8550 (N_8550,N_5951,N_3529);
or U8551 (N_8551,N_5428,N_5662);
xor U8552 (N_8552,N_3737,N_5719);
xor U8553 (N_8553,N_4423,N_3407);
nand U8554 (N_8554,N_5857,N_3270);
xor U8555 (N_8555,N_5119,N_3805);
nand U8556 (N_8556,N_5226,N_5207);
nand U8557 (N_8557,N_5105,N_5173);
and U8558 (N_8558,N_5369,N_3350);
and U8559 (N_8559,N_5650,N_5850);
and U8560 (N_8560,N_3097,N_5080);
nor U8561 (N_8561,N_4570,N_4290);
and U8562 (N_8562,N_3150,N_5680);
nand U8563 (N_8563,N_3446,N_3837);
nand U8564 (N_8564,N_4344,N_5224);
nand U8565 (N_8565,N_5961,N_3259);
and U8566 (N_8566,N_5166,N_5010);
and U8567 (N_8567,N_4895,N_3597);
and U8568 (N_8568,N_3583,N_3545);
or U8569 (N_8569,N_5963,N_5170);
and U8570 (N_8570,N_3214,N_3329);
nand U8571 (N_8571,N_3708,N_3556);
xor U8572 (N_8572,N_3214,N_4417);
or U8573 (N_8573,N_3757,N_3595);
or U8574 (N_8574,N_5022,N_3704);
xnor U8575 (N_8575,N_5506,N_4946);
and U8576 (N_8576,N_3532,N_5706);
or U8577 (N_8577,N_3193,N_5419);
or U8578 (N_8578,N_4600,N_3477);
nor U8579 (N_8579,N_5889,N_3276);
or U8580 (N_8580,N_5842,N_3086);
or U8581 (N_8581,N_4603,N_3452);
or U8582 (N_8582,N_5255,N_4549);
and U8583 (N_8583,N_5528,N_4606);
xor U8584 (N_8584,N_3515,N_4871);
nand U8585 (N_8585,N_4591,N_3039);
nor U8586 (N_8586,N_4339,N_4359);
and U8587 (N_8587,N_5031,N_4913);
and U8588 (N_8588,N_3155,N_5568);
nand U8589 (N_8589,N_5389,N_3920);
and U8590 (N_8590,N_4320,N_4872);
nor U8591 (N_8591,N_4233,N_3803);
and U8592 (N_8592,N_4157,N_5737);
xor U8593 (N_8593,N_4220,N_5576);
and U8594 (N_8594,N_4718,N_4175);
or U8595 (N_8595,N_4356,N_5772);
nor U8596 (N_8596,N_4399,N_3570);
xnor U8597 (N_8597,N_3923,N_3399);
or U8598 (N_8598,N_4441,N_4759);
nand U8599 (N_8599,N_5302,N_4675);
and U8600 (N_8600,N_4846,N_5232);
xnor U8601 (N_8601,N_4601,N_3157);
or U8602 (N_8602,N_3315,N_5783);
xnor U8603 (N_8603,N_4079,N_5045);
xor U8604 (N_8604,N_5753,N_5910);
nand U8605 (N_8605,N_4256,N_4745);
nor U8606 (N_8606,N_4595,N_4456);
or U8607 (N_8607,N_3842,N_5124);
nand U8608 (N_8608,N_5676,N_5544);
or U8609 (N_8609,N_3584,N_3029);
nand U8610 (N_8610,N_5089,N_3171);
and U8611 (N_8611,N_4894,N_5868);
nand U8612 (N_8612,N_5638,N_5705);
nor U8613 (N_8613,N_4762,N_3551);
nor U8614 (N_8614,N_5767,N_3490);
or U8615 (N_8615,N_4932,N_4097);
or U8616 (N_8616,N_5057,N_5987);
and U8617 (N_8617,N_5081,N_4919);
nor U8618 (N_8618,N_3910,N_5364);
nand U8619 (N_8619,N_3722,N_3021);
nor U8620 (N_8620,N_5406,N_4668);
nand U8621 (N_8621,N_5537,N_5770);
and U8622 (N_8622,N_3487,N_4844);
nor U8623 (N_8623,N_5621,N_4396);
xor U8624 (N_8624,N_3308,N_5118);
xor U8625 (N_8625,N_3809,N_3728);
nor U8626 (N_8626,N_4720,N_5183);
and U8627 (N_8627,N_3149,N_5839);
and U8628 (N_8628,N_5030,N_4399);
or U8629 (N_8629,N_3582,N_3092);
and U8630 (N_8630,N_3291,N_5994);
and U8631 (N_8631,N_5109,N_3267);
and U8632 (N_8632,N_5699,N_4833);
and U8633 (N_8633,N_5259,N_5386);
and U8634 (N_8634,N_3580,N_4172);
and U8635 (N_8635,N_5753,N_3744);
nor U8636 (N_8636,N_5964,N_3591);
nand U8637 (N_8637,N_4745,N_4145);
xor U8638 (N_8638,N_5578,N_4971);
nor U8639 (N_8639,N_3044,N_3888);
xnor U8640 (N_8640,N_4540,N_4172);
nand U8641 (N_8641,N_5945,N_5286);
nand U8642 (N_8642,N_4920,N_4156);
or U8643 (N_8643,N_4777,N_4937);
nand U8644 (N_8644,N_4888,N_4159);
and U8645 (N_8645,N_4236,N_5090);
or U8646 (N_8646,N_5678,N_5630);
or U8647 (N_8647,N_4778,N_3106);
xnor U8648 (N_8648,N_5816,N_5554);
or U8649 (N_8649,N_3382,N_3560);
nor U8650 (N_8650,N_4682,N_3096);
xnor U8651 (N_8651,N_5758,N_4941);
and U8652 (N_8652,N_4313,N_5677);
xor U8653 (N_8653,N_5105,N_3952);
xor U8654 (N_8654,N_4038,N_4244);
or U8655 (N_8655,N_4158,N_4456);
xor U8656 (N_8656,N_3506,N_5735);
nand U8657 (N_8657,N_3067,N_4183);
nand U8658 (N_8658,N_4813,N_4534);
xor U8659 (N_8659,N_5973,N_5208);
nor U8660 (N_8660,N_4036,N_5484);
nand U8661 (N_8661,N_5856,N_4236);
or U8662 (N_8662,N_3576,N_3150);
xor U8663 (N_8663,N_5417,N_5664);
nand U8664 (N_8664,N_5151,N_4453);
nor U8665 (N_8665,N_4704,N_3030);
or U8666 (N_8666,N_3551,N_5695);
xnor U8667 (N_8667,N_4217,N_5784);
and U8668 (N_8668,N_3904,N_3376);
and U8669 (N_8669,N_3993,N_3821);
xnor U8670 (N_8670,N_5876,N_4763);
xnor U8671 (N_8671,N_5172,N_3781);
xnor U8672 (N_8672,N_5078,N_5665);
nand U8673 (N_8673,N_3717,N_3331);
xor U8674 (N_8674,N_5213,N_3619);
or U8675 (N_8675,N_4250,N_4417);
nand U8676 (N_8676,N_5773,N_3284);
nor U8677 (N_8677,N_5289,N_5748);
nor U8678 (N_8678,N_5436,N_3894);
nand U8679 (N_8679,N_3782,N_4675);
xnor U8680 (N_8680,N_4062,N_4566);
nor U8681 (N_8681,N_3466,N_5991);
xor U8682 (N_8682,N_5704,N_5081);
nor U8683 (N_8683,N_3759,N_3107);
nor U8684 (N_8684,N_4821,N_5333);
nor U8685 (N_8685,N_3155,N_4293);
xnor U8686 (N_8686,N_5459,N_3462);
xnor U8687 (N_8687,N_3822,N_5802);
nor U8688 (N_8688,N_4355,N_5575);
nor U8689 (N_8689,N_5932,N_5687);
xnor U8690 (N_8690,N_3911,N_3961);
xnor U8691 (N_8691,N_5929,N_4251);
or U8692 (N_8692,N_5800,N_3451);
xnor U8693 (N_8693,N_3834,N_3428);
xnor U8694 (N_8694,N_3685,N_4385);
nand U8695 (N_8695,N_5169,N_5395);
nand U8696 (N_8696,N_5249,N_5548);
xor U8697 (N_8697,N_4820,N_5670);
and U8698 (N_8698,N_3769,N_4053);
xnor U8699 (N_8699,N_3549,N_5215);
nand U8700 (N_8700,N_5674,N_4680);
or U8701 (N_8701,N_3931,N_4005);
nand U8702 (N_8702,N_5480,N_5278);
xor U8703 (N_8703,N_4227,N_5921);
or U8704 (N_8704,N_4651,N_5600);
nand U8705 (N_8705,N_3440,N_4851);
nor U8706 (N_8706,N_5643,N_4047);
nor U8707 (N_8707,N_4447,N_3877);
xnor U8708 (N_8708,N_4443,N_4485);
nor U8709 (N_8709,N_5102,N_3996);
or U8710 (N_8710,N_5810,N_3539);
and U8711 (N_8711,N_3452,N_3971);
or U8712 (N_8712,N_3450,N_5783);
and U8713 (N_8713,N_4321,N_3454);
or U8714 (N_8714,N_5327,N_4739);
xnor U8715 (N_8715,N_3294,N_4114);
and U8716 (N_8716,N_3403,N_3540);
or U8717 (N_8717,N_4971,N_4194);
or U8718 (N_8718,N_4680,N_4705);
nor U8719 (N_8719,N_4635,N_4618);
or U8720 (N_8720,N_5797,N_3114);
nor U8721 (N_8721,N_4461,N_4779);
or U8722 (N_8722,N_4545,N_4883);
nor U8723 (N_8723,N_5883,N_5799);
nand U8724 (N_8724,N_5928,N_3496);
nor U8725 (N_8725,N_4968,N_3978);
nand U8726 (N_8726,N_5007,N_5107);
nor U8727 (N_8727,N_4214,N_5222);
and U8728 (N_8728,N_5219,N_3349);
and U8729 (N_8729,N_5358,N_5630);
nand U8730 (N_8730,N_5791,N_4696);
nor U8731 (N_8731,N_5139,N_5044);
nor U8732 (N_8732,N_3030,N_4754);
or U8733 (N_8733,N_4544,N_3995);
or U8734 (N_8734,N_4959,N_4727);
and U8735 (N_8735,N_3418,N_4447);
xnor U8736 (N_8736,N_3749,N_5952);
or U8737 (N_8737,N_3694,N_3358);
xnor U8738 (N_8738,N_3495,N_4351);
nor U8739 (N_8739,N_5802,N_3877);
and U8740 (N_8740,N_3480,N_4329);
nand U8741 (N_8741,N_4953,N_3656);
nor U8742 (N_8742,N_5506,N_5488);
and U8743 (N_8743,N_3225,N_5408);
nor U8744 (N_8744,N_5903,N_3334);
nand U8745 (N_8745,N_3287,N_4389);
nor U8746 (N_8746,N_4934,N_4101);
and U8747 (N_8747,N_5499,N_4759);
nand U8748 (N_8748,N_4941,N_4644);
and U8749 (N_8749,N_4199,N_4120);
nand U8750 (N_8750,N_3797,N_5611);
nor U8751 (N_8751,N_5456,N_5899);
xnor U8752 (N_8752,N_4777,N_4769);
nor U8753 (N_8753,N_4200,N_4603);
nor U8754 (N_8754,N_3915,N_3754);
or U8755 (N_8755,N_5214,N_4610);
or U8756 (N_8756,N_4792,N_4399);
or U8757 (N_8757,N_5588,N_5528);
or U8758 (N_8758,N_5296,N_5278);
nand U8759 (N_8759,N_5698,N_4080);
xor U8760 (N_8760,N_3454,N_5082);
xor U8761 (N_8761,N_4983,N_4097);
and U8762 (N_8762,N_5039,N_3453);
and U8763 (N_8763,N_3683,N_3884);
nor U8764 (N_8764,N_5744,N_5590);
and U8765 (N_8765,N_4443,N_5260);
and U8766 (N_8766,N_3945,N_4216);
xnor U8767 (N_8767,N_3986,N_4549);
nand U8768 (N_8768,N_3962,N_4099);
xnor U8769 (N_8769,N_5908,N_4739);
xor U8770 (N_8770,N_3632,N_5052);
and U8771 (N_8771,N_4874,N_4267);
nand U8772 (N_8772,N_5114,N_4815);
and U8773 (N_8773,N_4549,N_5173);
and U8774 (N_8774,N_3008,N_5306);
and U8775 (N_8775,N_5418,N_4014);
nand U8776 (N_8776,N_5837,N_5183);
nand U8777 (N_8777,N_5918,N_4391);
xnor U8778 (N_8778,N_3862,N_5406);
nor U8779 (N_8779,N_4171,N_5544);
or U8780 (N_8780,N_5698,N_5362);
nand U8781 (N_8781,N_4911,N_5775);
xor U8782 (N_8782,N_5118,N_4627);
or U8783 (N_8783,N_5232,N_3129);
nor U8784 (N_8784,N_5123,N_4128);
xor U8785 (N_8785,N_5927,N_3625);
or U8786 (N_8786,N_4736,N_3764);
nand U8787 (N_8787,N_5110,N_3088);
nand U8788 (N_8788,N_4472,N_3122);
nand U8789 (N_8789,N_5148,N_3857);
nor U8790 (N_8790,N_4886,N_5782);
nand U8791 (N_8791,N_3076,N_4512);
xnor U8792 (N_8792,N_4548,N_5192);
xnor U8793 (N_8793,N_3115,N_5764);
nor U8794 (N_8794,N_5722,N_5028);
and U8795 (N_8795,N_3425,N_3313);
nand U8796 (N_8796,N_4594,N_5276);
or U8797 (N_8797,N_5143,N_5333);
nor U8798 (N_8798,N_4432,N_5952);
or U8799 (N_8799,N_5021,N_4124);
nor U8800 (N_8800,N_5157,N_4122);
nand U8801 (N_8801,N_3022,N_3637);
and U8802 (N_8802,N_5333,N_4920);
xnor U8803 (N_8803,N_3162,N_3556);
and U8804 (N_8804,N_4296,N_3360);
and U8805 (N_8805,N_5114,N_5792);
nand U8806 (N_8806,N_3693,N_5275);
nand U8807 (N_8807,N_3726,N_3076);
nor U8808 (N_8808,N_5591,N_4573);
nand U8809 (N_8809,N_4265,N_5080);
and U8810 (N_8810,N_5602,N_4331);
and U8811 (N_8811,N_5828,N_3999);
or U8812 (N_8812,N_5866,N_3986);
and U8813 (N_8813,N_4276,N_5213);
or U8814 (N_8814,N_4478,N_4159);
nor U8815 (N_8815,N_3767,N_3899);
nor U8816 (N_8816,N_4702,N_5651);
nand U8817 (N_8817,N_4786,N_5178);
xnor U8818 (N_8818,N_3505,N_3988);
or U8819 (N_8819,N_4295,N_5717);
xnor U8820 (N_8820,N_5391,N_5357);
and U8821 (N_8821,N_3875,N_5021);
and U8822 (N_8822,N_5742,N_4815);
nor U8823 (N_8823,N_3430,N_5529);
nand U8824 (N_8824,N_4660,N_4017);
or U8825 (N_8825,N_4344,N_5717);
nand U8826 (N_8826,N_4214,N_4209);
and U8827 (N_8827,N_5855,N_5571);
nand U8828 (N_8828,N_3922,N_4943);
xnor U8829 (N_8829,N_3663,N_4224);
nor U8830 (N_8830,N_4650,N_4289);
and U8831 (N_8831,N_5859,N_3844);
nand U8832 (N_8832,N_5974,N_4294);
or U8833 (N_8833,N_5812,N_3059);
xor U8834 (N_8834,N_3300,N_3782);
nand U8835 (N_8835,N_4065,N_4414);
nand U8836 (N_8836,N_5306,N_3641);
or U8837 (N_8837,N_5734,N_3425);
nor U8838 (N_8838,N_5226,N_5622);
nand U8839 (N_8839,N_5227,N_4325);
nor U8840 (N_8840,N_3032,N_3804);
and U8841 (N_8841,N_3366,N_5814);
nor U8842 (N_8842,N_3441,N_5630);
xor U8843 (N_8843,N_4846,N_5263);
nand U8844 (N_8844,N_5574,N_4148);
xor U8845 (N_8845,N_4712,N_5265);
nand U8846 (N_8846,N_3272,N_4627);
nand U8847 (N_8847,N_3652,N_3210);
or U8848 (N_8848,N_3270,N_3327);
nor U8849 (N_8849,N_4446,N_5430);
and U8850 (N_8850,N_3339,N_3108);
nor U8851 (N_8851,N_3471,N_4420);
or U8852 (N_8852,N_3538,N_3262);
nor U8853 (N_8853,N_3167,N_5685);
nor U8854 (N_8854,N_5339,N_4717);
xnor U8855 (N_8855,N_3465,N_3866);
or U8856 (N_8856,N_5883,N_5078);
nor U8857 (N_8857,N_4321,N_3689);
nand U8858 (N_8858,N_3147,N_3357);
xor U8859 (N_8859,N_4652,N_4607);
nand U8860 (N_8860,N_4442,N_4476);
and U8861 (N_8861,N_3854,N_5203);
or U8862 (N_8862,N_4577,N_5336);
nand U8863 (N_8863,N_3692,N_5283);
or U8864 (N_8864,N_5052,N_5931);
and U8865 (N_8865,N_3909,N_3258);
nor U8866 (N_8866,N_5055,N_5240);
or U8867 (N_8867,N_5905,N_3467);
nand U8868 (N_8868,N_4884,N_3687);
or U8869 (N_8869,N_5800,N_3515);
or U8870 (N_8870,N_5932,N_3046);
nand U8871 (N_8871,N_5023,N_5646);
xnor U8872 (N_8872,N_4739,N_4247);
nand U8873 (N_8873,N_4208,N_4252);
and U8874 (N_8874,N_3850,N_3471);
nor U8875 (N_8875,N_4639,N_4189);
xnor U8876 (N_8876,N_3887,N_3341);
or U8877 (N_8877,N_4538,N_4450);
and U8878 (N_8878,N_3146,N_4055);
or U8879 (N_8879,N_4514,N_3222);
and U8880 (N_8880,N_4058,N_3332);
nand U8881 (N_8881,N_5979,N_5610);
and U8882 (N_8882,N_3494,N_5701);
xnor U8883 (N_8883,N_4400,N_4674);
or U8884 (N_8884,N_3515,N_3155);
and U8885 (N_8885,N_4223,N_5612);
or U8886 (N_8886,N_5822,N_5491);
xor U8887 (N_8887,N_4459,N_3454);
nand U8888 (N_8888,N_4743,N_5191);
or U8889 (N_8889,N_3277,N_5392);
nor U8890 (N_8890,N_5046,N_4191);
or U8891 (N_8891,N_5038,N_4248);
nor U8892 (N_8892,N_5814,N_5622);
or U8893 (N_8893,N_4025,N_4933);
or U8894 (N_8894,N_5257,N_3858);
and U8895 (N_8895,N_3230,N_3637);
nor U8896 (N_8896,N_5036,N_5955);
and U8897 (N_8897,N_4416,N_4682);
or U8898 (N_8898,N_5246,N_4506);
nor U8899 (N_8899,N_3914,N_4651);
nor U8900 (N_8900,N_4688,N_5759);
or U8901 (N_8901,N_4358,N_3834);
or U8902 (N_8902,N_3116,N_5244);
or U8903 (N_8903,N_5849,N_5611);
xnor U8904 (N_8904,N_4937,N_5265);
and U8905 (N_8905,N_4380,N_5120);
nand U8906 (N_8906,N_4756,N_5526);
or U8907 (N_8907,N_4649,N_4289);
xor U8908 (N_8908,N_3604,N_3288);
and U8909 (N_8909,N_3548,N_5604);
nor U8910 (N_8910,N_3489,N_5089);
and U8911 (N_8911,N_3314,N_3073);
or U8912 (N_8912,N_5058,N_5576);
nor U8913 (N_8913,N_3133,N_4102);
nand U8914 (N_8914,N_4520,N_3443);
and U8915 (N_8915,N_3705,N_3037);
and U8916 (N_8916,N_5952,N_3606);
or U8917 (N_8917,N_4135,N_3910);
nand U8918 (N_8918,N_5302,N_5336);
or U8919 (N_8919,N_4389,N_3289);
nor U8920 (N_8920,N_5135,N_5804);
nand U8921 (N_8921,N_4784,N_5410);
or U8922 (N_8922,N_4631,N_5417);
and U8923 (N_8923,N_4991,N_4612);
and U8924 (N_8924,N_4454,N_5292);
nor U8925 (N_8925,N_3465,N_4623);
or U8926 (N_8926,N_4252,N_5613);
nand U8927 (N_8927,N_4266,N_5967);
nor U8928 (N_8928,N_4940,N_4007);
nand U8929 (N_8929,N_4327,N_5927);
and U8930 (N_8930,N_4448,N_3103);
and U8931 (N_8931,N_3672,N_3311);
or U8932 (N_8932,N_5847,N_5114);
or U8933 (N_8933,N_3327,N_5494);
and U8934 (N_8934,N_4758,N_4102);
nor U8935 (N_8935,N_4049,N_3040);
nand U8936 (N_8936,N_5359,N_5215);
nand U8937 (N_8937,N_4504,N_3028);
and U8938 (N_8938,N_5573,N_3436);
and U8939 (N_8939,N_4083,N_3278);
nand U8940 (N_8940,N_4226,N_3859);
or U8941 (N_8941,N_3657,N_5875);
xnor U8942 (N_8942,N_5973,N_3739);
nor U8943 (N_8943,N_4059,N_5718);
nor U8944 (N_8944,N_5259,N_4168);
xor U8945 (N_8945,N_4647,N_4990);
and U8946 (N_8946,N_5703,N_5723);
nor U8947 (N_8947,N_3735,N_3672);
and U8948 (N_8948,N_4964,N_5520);
or U8949 (N_8949,N_5470,N_5566);
nand U8950 (N_8950,N_3273,N_5161);
and U8951 (N_8951,N_4749,N_3096);
nor U8952 (N_8952,N_3434,N_5986);
nor U8953 (N_8953,N_4149,N_4948);
nand U8954 (N_8954,N_3805,N_5718);
xor U8955 (N_8955,N_3575,N_5203);
nand U8956 (N_8956,N_3823,N_5316);
nor U8957 (N_8957,N_5651,N_5578);
nand U8958 (N_8958,N_5860,N_4449);
xor U8959 (N_8959,N_3938,N_3148);
and U8960 (N_8960,N_4372,N_3738);
xor U8961 (N_8961,N_4763,N_4525);
nor U8962 (N_8962,N_3006,N_4003);
nand U8963 (N_8963,N_4131,N_4563);
nand U8964 (N_8964,N_3980,N_3089);
nand U8965 (N_8965,N_4963,N_4721);
or U8966 (N_8966,N_5267,N_5920);
and U8967 (N_8967,N_5170,N_3701);
xor U8968 (N_8968,N_5271,N_5547);
xnor U8969 (N_8969,N_3396,N_3977);
or U8970 (N_8970,N_4093,N_4517);
or U8971 (N_8971,N_5311,N_4326);
nand U8972 (N_8972,N_5922,N_5490);
nor U8973 (N_8973,N_4965,N_3504);
and U8974 (N_8974,N_5040,N_4035);
xnor U8975 (N_8975,N_4326,N_3040);
or U8976 (N_8976,N_4090,N_4349);
or U8977 (N_8977,N_4076,N_4508);
nand U8978 (N_8978,N_5158,N_5616);
nand U8979 (N_8979,N_3024,N_3675);
nor U8980 (N_8980,N_4366,N_4652);
nand U8981 (N_8981,N_3483,N_5920);
xor U8982 (N_8982,N_3243,N_3934);
and U8983 (N_8983,N_4002,N_3182);
nor U8984 (N_8984,N_3002,N_3377);
nand U8985 (N_8985,N_5687,N_3954);
xnor U8986 (N_8986,N_4850,N_4133);
nor U8987 (N_8987,N_4744,N_3302);
xnor U8988 (N_8988,N_4005,N_5627);
and U8989 (N_8989,N_5801,N_5951);
and U8990 (N_8990,N_4776,N_4930);
nor U8991 (N_8991,N_5177,N_5599);
and U8992 (N_8992,N_3295,N_5700);
and U8993 (N_8993,N_5169,N_3361);
and U8994 (N_8994,N_3913,N_3796);
nand U8995 (N_8995,N_3889,N_5527);
nand U8996 (N_8996,N_5870,N_3352);
and U8997 (N_8997,N_3959,N_4753);
xnor U8998 (N_8998,N_3631,N_4756);
xor U8999 (N_8999,N_5164,N_4666);
nand U9000 (N_9000,N_7890,N_8115);
or U9001 (N_9001,N_7101,N_6240);
and U9002 (N_9002,N_7387,N_8769);
or U9003 (N_9003,N_6473,N_6187);
nor U9004 (N_9004,N_8009,N_8415);
nand U9005 (N_9005,N_7122,N_8167);
nor U9006 (N_9006,N_7845,N_6341);
nor U9007 (N_9007,N_6074,N_8621);
and U9008 (N_9008,N_7451,N_6602);
nor U9009 (N_9009,N_7084,N_6077);
and U9010 (N_9010,N_8835,N_8714);
nand U9011 (N_9011,N_6418,N_6351);
or U9012 (N_9012,N_8512,N_8157);
xnor U9013 (N_9013,N_6133,N_8248);
nor U9014 (N_9014,N_6304,N_8855);
nor U9015 (N_9015,N_8149,N_8561);
or U9016 (N_9016,N_6619,N_7734);
xnor U9017 (N_9017,N_7566,N_7558);
nor U9018 (N_9018,N_7386,N_8224);
nor U9019 (N_9019,N_8152,N_8554);
xnor U9020 (N_9020,N_8449,N_8334);
nand U9021 (N_9021,N_6655,N_7538);
xnor U9022 (N_9022,N_7365,N_6224);
nand U9023 (N_9023,N_6821,N_8631);
xnor U9024 (N_9024,N_6366,N_6663);
or U9025 (N_9025,N_8284,N_7415);
and U9026 (N_9026,N_7917,N_8087);
nor U9027 (N_9027,N_6108,N_7051);
and U9028 (N_9028,N_7202,N_6671);
nor U9029 (N_9029,N_7668,N_8367);
xnor U9030 (N_9030,N_7254,N_7870);
nand U9031 (N_9031,N_7424,N_7326);
xor U9032 (N_9032,N_7401,N_8303);
and U9033 (N_9033,N_7267,N_8520);
nand U9034 (N_9034,N_7186,N_8864);
nand U9035 (N_9035,N_7049,N_6135);
xor U9036 (N_9036,N_7394,N_7716);
and U9037 (N_9037,N_6317,N_6298);
xnor U9038 (N_9038,N_6612,N_8468);
nand U9039 (N_9039,N_7550,N_7212);
nand U9040 (N_9040,N_8885,N_7209);
nand U9041 (N_9041,N_8050,N_6168);
or U9042 (N_9042,N_6220,N_8223);
nand U9043 (N_9043,N_8814,N_7653);
nor U9044 (N_9044,N_6360,N_7712);
nand U9045 (N_9045,N_6729,N_7277);
nand U9046 (N_9046,N_7696,N_7025);
nor U9047 (N_9047,N_6182,N_8822);
xnor U9048 (N_9048,N_7602,N_8859);
and U9049 (N_9049,N_7982,N_6834);
xor U9050 (N_9050,N_8282,N_7536);
xor U9051 (N_9051,N_7891,N_6264);
or U9052 (N_9052,N_6871,N_6794);
nand U9053 (N_9053,N_7299,N_8083);
and U9054 (N_9054,N_6175,N_8884);
nor U9055 (N_9055,N_7247,N_6845);
xor U9056 (N_9056,N_8307,N_8811);
and U9057 (N_9057,N_7400,N_6557);
or U9058 (N_9058,N_7858,N_6183);
nand U9059 (N_9059,N_6722,N_7929);
nand U9060 (N_9060,N_6326,N_8498);
or U9061 (N_9061,N_8943,N_7809);
or U9062 (N_9062,N_7249,N_6858);
nor U9063 (N_9063,N_8955,N_6402);
xor U9064 (N_9064,N_8827,N_7239);
nor U9065 (N_9065,N_7573,N_7810);
nand U9066 (N_9066,N_6032,N_7062);
xnor U9067 (N_9067,N_8292,N_8857);
or U9068 (N_9068,N_7147,N_8636);
nand U9069 (N_9069,N_6842,N_8688);
and U9070 (N_9070,N_8099,N_8608);
or U9071 (N_9071,N_7083,N_7069);
nand U9072 (N_9072,N_6772,N_7989);
nand U9073 (N_9073,N_6892,N_8339);
and U9074 (N_9074,N_6007,N_6931);
nor U9075 (N_9075,N_8966,N_8557);
nor U9076 (N_9076,N_6451,N_7193);
or U9077 (N_9077,N_8024,N_6814);
nand U9078 (N_9078,N_8685,N_7624);
nand U9079 (N_9079,N_7606,N_7152);
and U9080 (N_9080,N_8027,N_8288);
nor U9081 (N_9081,N_6695,N_7555);
and U9082 (N_9082,N_6614,N_8493);
nor U9083 (N_9083,N_7360,N_6866);
and U9084 (N_9084,N_8926,N_8328);
nor U9085 (N_9085,N_8915,N_6202);
xnor U9086 (N_9086,N_8194,N_6422);
nor U9087 (N_9087,N_6361,N_6258);
or U9088 (N_9088,N_7919,N_7698);
or U9089 (N_9089,N_6376,N_6434);
nor U9090 (N_9090,N_6006,N_7674);
nor U9091 (N_9091,N_8635,N_7375);
and U9092 (N_9092,N_7578,N_7708);
nor U9093 (N_9093,N_6862,N_8191);
and U9094 (N_9094,N_7786,N_7508);
nand U9095 (N_9095,N_7746,N_6539);
nand U9096 (N_9096,N_7001,N_6825);
and U9097 (N_9097,N_6398,N_7397);
xor U9098 (N_9098,N_6761,N_6248);
nand U9099 (N_9099,N_7077,N_7681);
or U9100 (N_9100,N_8077,N_7070);
and U9101 (N_9101,N_8150,N_7645);
xnor U9102 (N_9102,N_7347,N_7704);
xnor U9103 (N_9103,N_8613,N_8438);
nor U9104 (N_9104,N_8136,N_6767);
nor U9105 (N_9105,N_7865,N_8564);
or U9106 (N_9106,N_7175,N_7851);
nand U9107 (N_9107,N_6705,N_7385);
nand U9108 (N_9108,N_7440,N_6420);
nand U9109 (N_9109,N_7279,N_6920);
or U9110 (N_9110,N_6324,N_7224);
or U9111 (N_9111,N_7906,N_7913);
nand U9112 (N_9112,N_8416,N_7967);
xor U9113 (N_9113,N_6868,N_6629);
xor U9114 (N_9114,N_8285,N_8421);
nor U9115 (N_9115,N_8126,N_8865);
nand U9116 (N_9116,N_8264,N_7446);
and U9117 (N_9117,N_7633,N_8940);
nand U9118 (N_9118,N_8779,N_7198);
or U9119 (N_9119,N_8957,N_7951);
nor U9120 (N_9120,N_6469,N_7769);
or U9121 (N_9121,N_6838,N_7887);
nor U9122 (N_9122,N_8364,N_8302);
and U9123 (N_9123,N_8450,N_8826);
or U9124 (N_9124,N_7987,N_8134);
nor U9125 (N_9125,N_7315,N_8251);
nand U9126 (N_9126,N_6070,N_8005);
xor U9127 (N_9127,N_8469,N_8403);
and U9128 (N_9128,N_6397,N_7842);
nor U9129 (N_9129,N_8732,N_6573);
or U9130 (N_9130,N_6743,N_6562);
or U9131 (N_9131,N_8791,N_6054);
nand U9132 (N_9132,N_7996,N_7369);
nand U9133 (N_9133,N_8122,N_6346);
or U9134 (N_9134,N_8394,N_6698);
nor U9135 (N_9135,N_7591,N_7110);
and U9136 (N_9136,N_8457,N_6273);
or U9137 (N_9137,N_8017,N_7355);
nor U9138 (N_9138,N_8369,N_7126);
and U9139 (N_9139,N_6714,N_7133);
xor U9140 (N_9140,N_6064,N_6977);
nand U9141 (N_9141,N_8413,N_8553);
and U9142 (N_9142,N_7530,N_6140);
xnor U9143 (N_9143,N_6738,N_8916);
xnor U9144 (N_9144,N_7148,N_8593);
xor U9145 (N_9145,N_7431,N_6918);
nand U9146 (N_9146,N_6606,N_8405);
xnor U9147 (N_9147,N_8383,N_6560);
or U9148 (N_9148,N_7030,N_8343);
and U9149 (N_9149,N_7767,N_7378);
xnor U9150 (N_9150,N_7690,N_6900);
xnor U9151 (N_9151,N_8423,N_6494);
nor U9152 (N_9152,N_6633,N_6253);
xnor U9153 (N_9153,N_8552,N_8802);
xor U9154 (N_9154,N_8500,N_6869);
and U9155 (N_9155,N_8116,N_7035);
and U9156 (N_9156,N_7151,N_7611);
xor U9157 (N_9157,N_7603,N_6975);
nand U9158 (N_9158,N_8333,N_7200);
xnor U9159 (N_9159,N_7398,N_7532);
nand U9160 (N_9160,N_8853,N_7302);
xor U9161 (N_9161,N_8962,N_7664);
or U9162 (N_9162,N_7737,N_7628);
nor U9163 (N_9163,N_8910,N_6957);
nand U9164 (N_9164,N_7004,N_8010);
and U9165 (N_9165,N_6748,N_7937);
or U9166 (N_9166,N_7998,N_7751);
or U9167 (N_9167,N_6826,N_7739);
nor U9168 (N_9168,N_8013,N_7017);
nor U9169 (N_9169,N_6238,N_7372);
nand U9170 (N_9170,N_8868,N_6086);
nor U9171 (N_9171,N_6198,N_8379);
nand U9172 (N_9172,N_6245,N_8794);
xor U9173 (N_9173,N_6340,N_7461);
nand U9174 (N_9174,N_6699,N_8776);
and U9175 (N_9175,N_7112,N_8053);
nor U9176 (N_9176,N_6137,N_7984);
nor U9177 (N_9177,N_8001,N_8588);
nand U9178 (N_9178,N_6459,N_6526);
or U9179 (N_9179,N_8983,N_7777);
nand U9180 (N_9180,N_8491,N_8754);
nor U9181 (N_9181,N_7968,N_7284);
nor U9182 (N_9182,N_7881,N_8075);
and U9183 (N_9183,N_8014,N_6058);
xnor U9184 (N_9184,N_8159,N_7564);
nand U9185 (N_9185,N_7185,N_7918);
and U9186 (N_9186,N_8929,N_7228);
and U9187 (N_9187,N_6713,N_8121);
xor U9188 (N_9188,N_6724,N_6684);
and U9189 (N_9189,N_8020,N_8816);
and U9190 (N_9190,N_6396,N_6157);
xnor U9191 (N_9191,N_8874,N_6085);
xor U9192 (N_9192,N_6964,N_8625);
nor U9193 (N_9193,N_7731,N_8569);
xnor U9194 (N_9194,N_8390,N_8591);
nand U9195 (N_9195,N_6437,N_7509);
or U9196 (N_9196,N_8870,N_8205);
or U9197 (N_9197,N_6255,N_6073);
and U9198 (N_9198,N_6783,N_6582);
nand U9199 (N_9199,N_7620,N_7502);
nor U9200 (N_9200,N_6912,N_8900);
nor U9201 (N_9201,N_8353,N_7297);
xnor U9202 (N_9202,N_7685,N_6408);
or U9203 (N_9203,N_8660,N_7325);
nand U9204 (N_9204,N_6590,N_8479);
or U9205 (N_9205,N_6711,N_6847);
and U9206 (N_9206,N_8495,N_6903);
xnor U9207 (N_9207,N_7539,N_7097);
and U9208 (N_9208,N_8630,N_6488);
nand U9209 (N_9209,N_7003,N_8725);
and U9210 (N_9210,N_6899,N_6696);
and U9211 (N_9211,N_6493,N_8861);
xnor U9212 (N_9212,N_6604,N_7684);
nand U9213 (N_9213,N_7971,N_8540);
or U9214 (N_9214,N_7854,N_6929);
xor U9215 (N_9215,N_6307,N_7163);
nand U9216 (N_9216,N_7484,N_7406);
nand U9217 (N_9217,N_8742,N_6116);
nor U9218 (N_9218,N_7172,N_8187);
and U9219 (N_9219,N_6667,N_6063);
and U9220 (N_9220,N_7912,N_8699);
nor U9221 (N_9221,N_6372,N_7165);
and U9222 (N_9222,N_7453,N_6803);
and U9223 (N_9223,N_6647,N_7039);
xnor U9224 (N_9224,N_6342,N_6822);
xnor U9225 (N_9225,N_6263,N_6512);
or U9226 (N_9226,N_8104,N_7817);
or U9227 (N_9227,N_6867,N_6286);
xnor U9228 (N_9228,N_6109,N_8833);
nor U9229 (N_9229,N_6158,N_7506);
nor U9230 (N_9230,N_8033,N_8108);
and U9231 (N_9231,N_8237,N_7104);
nor U9232 (N_9232,N_8756,N_7150);
nand U9233 (N_9233,N_8290,N_7371);
nand U9234 (N_9234,N_7142,N_8674);
xnor U9235 (N_9235,N_8072,N_6712);
or U9236 (N_9236,N_7309,N_8628);
xnor U9237 (N_9237,N_7100,N_6002);
xor U9238 (N_9238,N_8101,N_6840);
nand U9239 (N_9239,N_8120,N_7487);
nor U9240 (N_9240,N_8797,N_8444);
or U9241 (N_9241,N_8329,N_6913);
nand U9242 (N_9242,N_6855,N_6887);
nand U9243 (N_9243,N_8546,N_6678);
nand U9244 (N_9244,N_7547,N_7710);
nand U9245 (N_9245,N_6019,N_7534);
nor U9246 (N_9246,N_8891,N_6670);
xor U9247 (N_9247,N_8718,N_8375);
and U9248 (N_9248,N_7503,N_6148);
xor U9249 (N_9249,N_6078,N_7518);
or U9250 (N_9250,N_7529,N_6546);
nand U9251 (N_9251,N_7659,N_6830);
or U9252 (N_9252,N_6672,N_7208);
nand U9253 (N_9253,N_6289,N_7635);
xnor U9254 (N_9254,N_8793,N_8559);
xor U9255 (N_9255,N_6156,N_6444);
or U9256 (N_9256,N_8085,N_6125);
xnor U9257 (N_9257,N_6436,N_8509);
nor U9258 (N_9258,N_7825,N_8642);
xnor U9259 (N_9259,N_6679,N_8841);
nand U9260 (N_9260,N_8888,N_7044);
or U9261 (N_9261,N_6501,N_8417);
nor U9262 (N_9262,N_7362,N_8587);
or U9263 (N_9263,N_6336,N_7513);
xor U9264 (N_9264,N_8501,N_7679);
xnor U9265 (N_9265,N_7457,N_6476);
nand U9266 (N_9266,N_7333,N_8872);
nand U9267 (N_9267,N_8357,N_7584);
xor U9268 (N_9268,N_6204,N_6233);
nor U9269 (N_9269,N_6262,N_6736);
nor U9270 (N_9270,N_7806,N_7310);
nand U9271 (N_9271,N_8633,N_6201);
nor U9272 (N_9272,N_6642,N_7059);
xor U9273 (N_9273,N_7233,N_7115);
nand U9274 (N_9274,N_8456,N_6591);
xnor U9275 (N_9275,N_7949,N_6645);
xor U9276 (N_9276,N_7352,N_7318);
nor U9277 (N_9277,N_6164,N_6160);
xnor U9278 (N_9278,N_6940,N_8453);
nand U9279 (N_9279,N_8103,N_7724);
xnor U9280 (N_9280,N_7376,N_6214);
and U9281 (N_9281,N_7293,N_7693);
nor U9282 (N_9282,N_7849,N_6856);
nand U9283 (N_9283,N_8110,N_8098);
or U9284 (N_9284,N_8984,N_7976);
and U9285 (N_9285,N_6643,N_8039);
nor U9286 (N_9286,N_8186,N_7833);
nor U9287 (N_9287,N_7818,N_7742);
or U9288 (N_9288,N_7441,N_6104);
and U9289 (N_9289,N_6400,N_8766);
and U9290 (N_9290,N_6723,N_6260);
nor U9291 (N_9291,N_8492,N_8620);
nor U9292 (N_9292,N_8942,N_7923);
and U9293 (N_9293,N_7066,N_7229);
nand U9294 (N_9294,N_7834,N_8645);
and U9295 (N_9295,N_7839,N_7311);
nor U9296 (N_9296,N_7242,N_6951);
nand U9297 (N_9297,N_7182,N_6159);
or U9298 (N_9298,N_7661,N_8052);
or U9299 (N_9299,N_8174,N_8429);
nor U9300 (N_9300,N_7480,N_7308);
and U9301 (N_9301,N_8722,N_7540);
nor U9302 (N_9302,N_7535,N_8499);
nand U9303 (N_9303,N_6517,N_8536);
nand U9304 (N_9304,N_7885,N_8063);
or U9305 (N_9305,N_7493,N_7094);
or U9306 (N_9306,N_6066,N_8892);
xor U9307 (N_9307,N_8578,N_6211);
nand U9308 (N_9308,N_6394,N_6014);
xor U9309 (N_9309,N_8040,N_7468);
nor U9310 (N_9310,N_7301,N_6507);
nand U9311 (N_9311,N_8312,N_6807);
xnor U9312 (N_9312,N_7648,N_8238);
and U9313 (N_9313,N_7711,N_7986);
nor U9314 (N_9314,N_8580,N_8852);
nand U9315 (N_9315,N_7304,N_8084);
xnor U9316 (N_9316,N_6190,N_8476);
nor U9317 (N_9317,N_8004,N_6297);
or U9318 (N_9318,N_7978,N_8740);
nor U9319 (N_9319,N_8330,N_6901);
xor U9320 (N_9320,N_6854,N_6735);
xnor U9321 (N_9321,N_8177,N_6680);
xnor U9322 (N_9322,N_6257,N_7459);
and U9323 (N_9323,N_8597,N_6658);
xor U9324 (N_9324,N_8135,N_7064);
or U9325 (N_9325,N_8064,N_6254);
or U9326 (N_9326,N_8694,N_8189);
or U9327 (N_9327,N_8951,N_7735);
nor U9328 (N_9328,N_8477,N_7541);
xnor U9329 (N_9329,N_6999,N_8373);
nor U9330 (N_9330,N_7879,N_7181);
xnor U9331 (N_9331,N_8350,N_7383);
xnor U9332 (N_9332,N_8474,N_6831);
nand U9333 (N_9333,N_6091,N_8650);
and U9334 (N_9334,N_7482,N_8678);
nor U9335 (N_9335,N_6305,N_8480);
nor U9336 (N_9336,N_8012,N_7837);
nor U9337 (N_9337,N_6449,N_6448);
nand U9338 (N_9338,N_8676,N_7481);
nor U9339 (N_9339,N_7013,N_7907);
and U9340 (N_9340,N_6985,N_7449);
nor U9341 (N_9341,N_8978,N_8335);
nor U9342 (N_9342,N_7802,N_6122);
nor U9343 (N_9343,N_8679,N_7957);
nor U9344 (N_9344,N_8031,N_6581);
or U9345 (N_9345,N_8547,N_8619);
nand U9346 (N_9346,N_8397,N_8686);
or U9347 (N_9347,N_7350,N_8575);
nand U9348 (N_9348,N_8968,N_8148);
xnor U9349 (N_9349,N_6259,N_8213);
nand U9350 (N_9350,N_7382,N_8374);
nor U9351 (N_9351,N_7814,N_6112);
or U9352 (N_9352,N_8400,N_8834);
or U9353 (N_9353,N_8018,N_7332);
nand U9354 (N_9354,N_7156,N_6513);
nor U9355 (N_9355,N_7761,N_6504);
nand U9356 (N_9356,N_6313,N_7426);
or U9357 (N_9357,N_6768,N_6318);
nor U9358 (N_9358,N_7280,N_6242);
or U9359 (N_9359,N_7991,N_6098);
or U9360 (N_9360,N_8022,N_7447);
or U9361 (N_9361,N_7168,N_7510);
nand U9362 (N_9362,N_8930,N_7463);
nor U9363 (N_9363,N_6849,N_8412);
nand U9364 (N_9364,N_7791,N_7812);
and U9365 (N_9365,N_8704,N_8418);
xnor U9366 (N_9366,N_6719,N_8875);
and U9367 (N_9367,N_8651,N_6335);
and U9368 (N_9368,N_6333,N_6595);
or U9369 (N_9369,N_8629,N_8804);
nand U9370 (N_9370,N_6235,N_8617);
xor U9371 (N_9371,N_6483,N_7599);
nand U9372 (N_9372,N_6843,N_6456);
and U9373 (N_9373,N_6447,N_7292);
nand U9374 (N_9374,N_8850,N_7469);
nand U9375 (N_9375,N_8646,N_7335);
or U9376 (N_9376,N_6720,N_7617);
xnor U9377 (N_9377,N_8858,N_7119);
nor U9378 (N_9378,N_6439,N_8311);
and U9379 (N_9379,N_8076,N_6495);
nand U9380 (N_9380,N_8585,N_7046);
and U9381 (N_9381,N_8551,N_8911);
nor U9382 (N_9382,N_8511,N_8082);
or U9383 (N_9383,N_8549,N_7373);
and U9384 (N_9384,N_6725,N_6668);
nand U9385 (N_9385,N_8784,N_7222);
xnor U9386 (N_9386,N_8935,N_6005);
xor U9387 (N_9387,N_7807,N_7354);
and U9388 (N_9388,N_8706,N_8703);
nand U9389 (N_9389,N_8556,N_8466);
or U9390 (N_9390,N_8781,N_6580);
xnor U9391 (N_9391,N_7725,N_7927);
nand U9392 (N_9392,N_7056,N_8181);
xor U9393 (N_9393,N_8927,N_8602);
xor U9394 (N_9394,N_7052,N_7959);
xor U9395 (N_9395,N_6615,N_8934);
and U9396 (N_9396,N_7939,N_8941);
xnor U9397 (N_9397,N_6545,N_8320);
and U9398 (N_9398,N_8021,N_8259);
and U9399 (N_9399,N_7798,N_6395);
or U9400 (N_9400,N_6100,N_6778);
nand U9401 (N_9401,N_6654,N_6171);
nor U9402 (N_9402,N_6811,N_7883);
nor U9403 (N_9403,N_8147,N_8598);
and U9404 (N_9404,N_8690,N_6056);
nand U9405 (N_9405,N_8961,N_7638);
xnor U9406 (N_9406,N_6250,N_7336);
and U9407 (N_9407,N_8319,N_8089);
xnor U9408 (N_9408,N_8830,N_7847);
nand U9409 (N_9409,N_8296,N_6217);
xnor U9410 (N_9410,N_6067,N_6609);
nand U9411 (N_9411,N_6636,N_8939);
or U9412 (N_9412,N_8821,N_6824);
and U9413 (N_9413,N_6308,N_8372);
nand U9414 (N_9414,N_6045,N_8442);
nor U9415 (N_9415,N_8204,N_6191);
nor U9416 (N_9416,N_7632,N_8097);
and U9417 (N_9417,N_8572,N_7811);
xnor U9418 (N_9418,N_7423,N_8595);
nor U9419 (N_9419,N_7238,N_6648);
or U9420 (N_9420,N_8963,N_6674);
or U9421 (N_9421,N_8356,N_6919);
and U9422 (N_9422,N_7892,N_8171);
and U9423 (N_9423,N_6432,N_7138);
nor U9424 (N_9424,N_7639,N_7464);
nand U9425 (N_9425,N_7730,N_6344);
and U9426 (N_9426,N_7889,N_6121);
nor U9427 (N_9427,N_7637,N_7067);
nor U9428 (N_9428,N_7250,N_7214);
or U9429 (N_9429,N_6290,N_8483);
nor U9430 (N_9430,N_6890,N_7295);
or U9431 (N_9431,N_8661,N_6411);
and U9432 (N_9432,N_8436,N_8749);
xor U9433 (N_9433,N_7585,N_8848);
xnor U9434 (N_9434,N_8153,N_6509);
or U9435 (N_9435,N_8484,N_7546);
nor U9436 (N_9436,N_6320,N_7257);
and U9437 (N_9437,N_6563,N_8521);
xnor U9438 (N_9438,N_7577,N_6029);
nor U9439 (N_9439,N_6142,N_8663);
xnor U9440 (N_9440,N_7896,N_8516);
and U9441 (N_9441,N_7246,N_6928);
nand U9442 (N_9442,N_8565,N_7367);
or U9443 (N_9443,N_6246,N_8216);
or U9444 (N_9444,N_7264,N_7970);
or U9445 (N_9445,N_6206,N_7932);
or U9446 (N_9446,N_6564,N_7473);
xnor U9447 (N_9447,N_7691,N_6130);
or U9448 (N_9448,N_8698,N_8658);
nand U9449 (N_9449,N_7521,N_7655);
or U9450 (N_9450,N_6886,N_7060);
or U9451 (N_9451,N_7328,N_8041);
or U9452 (N_9452,N_7205,N_8971);
or U9453 (N_9453,N_7033,N_8139);
or U9454 (N_9454,N_6022,N_6229);
nor U9455 (N_9455,N_7341,N_7680);
nand U9456 (N_9456,N_7960,N_6661);
and U9457 (N_9457,N_6981,N_6758);
or U9458 (N_9458,N_8158,N_8839);
nor U9459 (N_9459,N_8964,N_8355);
xnor U9460 (N_9460,N_6195,N_8151);
nor U9461 (N_9461,N_7947,N_8592);
or U9462 (N_9462,N_7132,N_6367);
nor U9463 (N_9463,N_6927,N_8051);
xnor U9464 (N_9464,N_8812,N_8573);
nand U9465 (N_9465,N_7569,N_6487);
or U9466 (N_9466,N_7794,N_7211);
nor U9467 (N_9467,N_6948,N_8904);
xnor U9468 (N_9468,N_8346,N_8026);
nor U9469 (N_9469,N_7090,N_8730);
nor U9470 (N_9470,N_6071,N_7993);
nor U9471 (N_9471,N_8252,N_6416);
nor U9472 (N_9472,N_6793,N_7269);
xor U9473 (N_9473,N_6425,N_7894);
or U9474 (N_9474,N_6092,N_8867);
and U9475 (N_9475,N_8972,N_6544);
and U9476 (N_9476,N_7861,N_6079);
or U9477 (N_9477,N_6385,N_6052);
or U9478 (N_9478,N_8287,N_6616);
xor U9479 (N_9479,N_6549,N_6124);
xnor U9480 (N_9480,N_6287,N_6480);
nand U9481 (N_9481,N_8815,N_8127);
nand U9482 (N_9482,N_7241,N_8384);
nand U9483 (N_9483,N_6357,N_6710);
nor U9484 (N_9484,N_8154,N_8295);
and U9485 (N_9485,N_7721,N_7765);
or U9486 (N_9486,N_8970,N_6355);
or U9487 (N_9487,N_7590,N_6910);
and U9488 (N_9488,N_6089,N_6804);
and U9489 (N_9489,N_6417,N_8649);
nand U9490 (N_9490,N_7728,N_8519);
and U9491 (N_9491,N_6316,N_6129);
and U9492 (N_9492,N_6863,N_7930);
nor U9493 (N_9493,N_7501,N_8785);
and U9494 (N_9494,N_6252,N_8684);
xnor U9495 (N_9495,N_6799,N_6628);
nor U9496 (N_9496,N_7225,N_6631);
nand U9497 (N_9497,N_7985,N_7687);
or U9498 (N_9498,N_7219,N_8234);
nor U9499 (N_9499,N_6584,N_8432);
and U9500 (N_9500,N_6055,N_7210);
nor U9501 (N_9501,N_8341,N_7650);
xnor U9502 (N_9502,N_8998,N_7291);
nor U9503 (N_9503,N_7629,N_8192);
nand U9504 (N_9504,N_7149,N_6350);
and U9505 (N_9505,N_7404,N_8316);
and U9506 (N_9506,N_7324,N_8318);
xor U9507 (N_9507,N_6765,N_8772);
or U9508 (N_9508,N_6013,N_6044);
or U9509 (N_9509,N_8215,N_8399);
or U9510 (N_9510,N_8060,N_7941);
and U9511 (N_9511,N_6419,N_8472);
and U9512 (N_9512,N_7448,N_6393);
nor U9513 (N_9513,N_8568,N_7203);
nor U9514 (N_9514,N_6176,N_6115);
nor U9515 (N_9515,N_8199,N_7327);
and U9516 (N_9516,N_6503,N_6345);
and U9517 (N_9517,N_8866,N_8952);
xnor U9518 (N_9518,N_7544,N_6440);
or U9519 (N_9519,N_8377,N_6084);
nand U9520 (N_9520,N_8701,N_6199);
nand U9521 (N_9521,N_8178,N_7427);
and U9522 (N_9522,N_8210,N_7570);
nand U9523 (N_9523,N_6010,N_8596);
nand U9524 (N_9524,N_7549,N_7995);
xnor U9525 (N_9525,N_8693,N_7779);
nor U9526 (N_9526,N_8354,N_8969);
nand U9527 (N_9527,N_6944,N_7497);
or U9528 (N_9528,N_8166,N_7827);
nor U9529 (N_9529,N_8548,N_8677);
xor U9530 (N_9530,N_6755,N_8283);
or U9531 (N_9531,N_8475,N_7283);
nor U9532 (N_9532,N_7492,N_6585);
xnor U9533 (N_9533,N_6823,N_6623);
nor U9534 (N_9534,N_8304,N_8297);
xnor U9535 (N_9535,N_8571,N_8081);
nor U9536 (N_9536,N_8993,N_7750);
nor U9537 (N_9537,N_6382,N_6813);
or U9538 (N_9538,N_8239,N_8624);
or U9539 (N_9539,N_7820,N_7667);
or U9540 (N_9540,N_6935,N_7741);
nand U9541 (N_9541,N_7091,N_7012);
nor U9542 (N_9542,N_8535,N_7815);
nand U9543 (N_9543,N_8030,N_8043);
xnor U9544 (N_9544,N_6567,N_6916);
nor U9545 (N_9545,N_7405,N_8753);
or U9546 (N_9546,N_7718,N_6737);
and U9547 (N_9547,N_7934,N_6216);
or U9548 (N_9548,N_7034,N_6276);
nand U9549 (N_9549,N_6475,N_6482);
and U9550 (N_9550,N_8755,N_6530);
nand U9551 (N_9551,N_6676,N_6038);
or U9552 (N_9552,N_6659,N_6787);
or U9553 (N_9553,N_6547,N_8527);
nor U9554 (N_9554,N_7800,N_8879);
nor U9555 (N_9555,N_6174,N_6872);
xnor U9556 (N_9556,N_7675,N_6008);
or U9557 (N_9557,N_7412,N_7207);
nand U9558 (N_9558,N_7478,N_6579);
xnor U9559 (N_9559,N_7184,N_6034);
xor U9560 (N_9560,N_8305,N_8321);
or U9561 (N_9561,N_6465,N_6709);
or U9562 (N_9562,N_6586,N_7528);
nand U9563 (N_9563,N_7963,N_6638);
nand U9564 (N_9564,N_6572,N_7719);
and U9565 (N_9565,N_8623,N_8281);
nor U9566 (N_9566,N_7232,N_6461);
or U9567 (N_9567,N_8562,N_8173);
xnor U9568 (N_9568,N_7206,N_7723);
xor U9569 (N_9569,N_6354,N_6181);
xor U9570 (N_9570,N_6173,N_6953);
or U9571 (N_9571,N_6797,N_6889);
nand U9572 (N_9572,N_7144,N_7433);
nand U9573 (N_9573,N_7038,N_7079);
nand U9574 (N_9574,N_8293,N_7623);
or U9575 (N_9575,N_6053,N_8100);
nor U9576 (N_9576,N_6523,N_7490);
or U9577 (N_9577,N_6337,N_7343);
xnor U9578 (N_9578,N_6261,N_8576);
nor U9579 (N_9579,N_6165,N_7096);
or U9580 (N_9580,N_7409,N_6939);
and U9581 (N_9581,N_8140,N_8836);
nor U9582 (N_9582,N_6911,N_6649);
or U9583 (N_9583,N_8317,N_7613);
and U9584 (N_9584,N_7980,N_7054);
or U9585 (N_9585,N_8249,N_7878);
and U9586 (N_9586,N_7136,N_6618);
xor U9587 (N_9587,N_8124,N_6365);
or U9588 (N_9588,N_8818,N_8410);
and U9589 (N_9589,N_6285,N_8708);
and U9590 (N_9590,N_7874,N_6080);
nand U9591 (N_9591,N_8482,N_6763);
and U9592 (N_9592,N_8856,N_7312);
and U9593 (N_9593,N_6596,N_7141);
nand U9594 (N_9594,N_7342,N_7384);
or U9595 (N_9595,N_6334,N_7475);
nor U9596 (N_9596,N_6943,N_6859);
or U9597 (N_9597,N_8670,N_7275);
nand U9598 (N_9598,N_6293,N_8680);
nand U9599 (N_9599,N_8513,N_7895);
xor U9600 (N_9600,N_6409,N_6020);
or U9601 (N_9601,N_7288,N_6101);
or U9602 (N_9602,N_8666,N_6841);
nand U9603 (N_9603,N_6474,N_7127);
xnor U9604 (N_9604,N_8228,N_7568);
nor U9605 (N_9605,N_6373,N_8751);
xor U9606 (N_9606,N_6926,N_8743);
and U9607 (N_9607,N_8395,N_6151);
nand U9608 (N_9608,N_7793,N_7491);
nand U9609 (N_9609,N_7792,N_8225);
or U9610 (N_9610,N_8409,N_8905);
and U9611 (N_9611,N_7676,N_8214);
nand U9612 (N_9612,N_6491,N_6144);
and U9613 (N_9613,N_7533,N_8895);
xor U9614 (N_9614,N_8849,N_7022);
and U9615 (N_9615,N_7908,N_6088);
or U9616 (N_9616,N_8525,N_7155);
and U9617 (N_9617,N_6511,N_7788);
xor U9618 (N_9618,N_8542,N_8419);
nor U9619 (N_9619,N_8144,N_8783);
xnor U9620 (N_9620,N_7770,N_7485);
nor U9621 (N_9621,N_7313,N_6424);
nor U9622 (N_9622,N_8738,N_6702);
nor U9623 (N_9623,N_7099,N_8717);
nand U9624 (N_9624,N_7187,N_7443);
xor U9625 (N_9625,N_7626,N_7007);
or U9626 (N_9626,N_7768,N_8696);
nand U9627 (N_9627,N_6374,N_7672);
and U9628 (N_9628,N_7559,N_8447);
xnor U9629 (N_9629,N_6639,N_8925);
xor U9630 (N_9630,N_8455,N_8058);
nor U9631 (N_9631,N_6734,N_7036);
nor U9632 (N_9632,N_6846,N_8634);
nor U9633 (N_9633,N_7160,N_8074);
and U9634 (N_9634,N_8131,N_7065);
or U9635 (N_9635,N_6681,N_8193);
nor U9636 (N_9636,N_8002,N_8665);
nand U9637 (N_9637,N_6392,N_7088);
or U9638 (N_9638,N_6906,N_8486);
nand U9639 (N_9639,N_7425,N_8528);
nand U9640 (N_9640,N_7909,N_7709);
xnor U9641 (N_9641,N_8770,N_7024);
nand U9642 (N_9642,N_7922,N_6952);
nand U9643 (N_9643,N_6568,N_6178);
xor U9644 (N_9644,N_6971,N_8654);
nor U9645 (N_9645,N_7699,N_8803);
and U9646 (N_9646,N_6210,N_6715);
and U9647 (N_9647,N_7230,N_8838);
or U9648 (N_9648,N_8744,N_8982);
and U9649 (N_9649,N_6945,N_7169);
xnor U9650 (N_9650,N_8070,N_8757);
nor U9651 (N_9651,N_6792,N_6068);
and U9652 (N_9652,N_8376,N_6861);
or U9653 (N_9653,N_7763,N_7582);
or U9654 (N_9654,N_6274,N_6508);
nand U9655 (N_9655,N_6356,N_8898);
nand U9656 (N_9656,N_6477,N_6731);
nor U9657 (N_9657,N_8828,N_6302);
xnor U9658 (N_9658,N_8366,N_6976);
or U9659 (N_9659,N_7429,N_8775);
nand U9660 (N_9660,N_8908,N_8627);
and U9661 (N_9661,N_8632,N_7109);
or U9662 (N_9662,N_6384,N_8990);
xnor U9663 (N_9663,N_8203,N_7621);
nand U9664 (N_9664,N_8401,N_7130);
or U9665 (N_9665,N_7220,N_8129);
nor U9666 (N_9666,N_8411,N_6241);
xnor U9667 (N_9667,N_8824,N_6662);
xor U9668 (N_9668,N_7268,N_7260);
nor U9669 (N_9669,N_7616,N_8049);
or U9670 (N_9670,N_8581,N_7647);
nand U9671 (N_9671,N_7002,N_6136);
and U9672 (N_9672,N_8338,N_7732);
and U9673 (N_9673,N_7303,N_8746);
or U9674 (N_9674,N_7388,N_7527);
or U9675 (N_9675,N_7966,N_7435);
nor U9676 (N_9676,N_7251,N_8953);
or U9677 (N_9677,N_6788,N_6817);
nor U9678 (N_9678,N_6893,N_6865);
xnor U9679 (N_9679,N_7795,N_7450);
xor U9680 (N_9680,N_7472,N_8382);
and U9681 (N_9681,N_6706,N_8107);
xnor U9682 (N_9682,N_8331,N_6707);
and U9683 (N_9683,N_8426,N_6898);
nand U9684 (N_9684,N_6134,N_8380);
xor U9685 (N_9685,N_6990,N_6270);
or U9686 (N_9686,N_8638,N_7216);
xnor U9687 (N_9687,N_8119,N_8558);
nand U9688 (N_9688,N_8428,N_8887);
or U9689 (N_9689,N_7467,N_6251);
nor U9690 (N_9690,N_6894,N_7901);
xor U9691 (N_9691,N_6404,N_7579);
xnor U9692 (N_9692,N_7396,N_7413);
or U9693 (N_9693,N_7819,N_8143);
nand U9694 (N_9694,N_6770,N_6601);
or U9695 (N_9695,N_8219,N_8197);
nand U9696 (N_9696,N_8459,N_7726);
nor U9697 (N_9697,N_8876,N_7722);
nor U9698 (N_9698,N_6377,N_6727);
or U9699 (N_9699,N_6611,N_6594);
or U9700 (N_9700,N_8061,N_7531);
nand U9701 (N_9701,N_8526,N_7563);
or U9702 (N_9702,N_7643,N_8946);
nand U9703 (N_9703,N_6980,N_7381);
or U9704 (N_9704,N_7418,N_6492);
xor U9705 (N_9705,N_6496,N_8913);
and U9706 (N_9706,N_7784,N_7348);
xnor U9707 (N_9707,N_7074,N_8997);
nand U9708 (N_9708,N_8422,N_7262);
nor U9709 (N_9709,N_8726,N_6577);
and U9710 (N_9710,N_8705,N_8359);
or U9711 (N_9711,N_6265,N_8878);
nand U9712 (N_9712,N_6632,N_6172);
xnor U9713 (N_9713,N_7331,N_6490);
or U9714 (N_9714,N_7636,N_8948);
xnor U9715 (N_9715,N_7121,N_6769);
or U9716 (N_9716,N_7201,N_7964);
xor U9717 (N_9717,N_7474,N_6653);
nor U9718 (N_9718,N_8539,N_6888);
nand U9719 (N_9719,N_6207,N_6150);
nor U9720 (N_9720,N_8042,N_7021);
xnor U9721 (N_9721,N_8047,N_8464);
or U9722 (N_9722,N_7043,N_7120);
nand U9723 (N_9723,N_8989,N_6048);
nand U9724 (N_9724,N_7143,N_8188);
nand U9725 (N_9725,N_7697,N_6617);
nor U9726 (N_9726,N_7128,N_8274);
or U9727 (N_9727,N_7042,N_8172);
xnor U9728 (N_9728,N_7285,N_8733);
xor U9729 (N_9729,N_7938,N_6836);
or U9730 (N_9730,N_7933,N_8768);
nor U9731 (N_9731,N_7618,N_6030);
xor U9732 (N_9732,N_8724,N_7057);
nand U9733 (N_9733,N_6554,N_8737);
xor U9734 (N_9734,N_6962,N_7754);
or U9735 (N_9735,N_8894,N_8351);
xor U9736 (N_9736,N_8924,N_8425);
and U9737 (N_9737,N_8954,N_7720);
nor U9738 (N_9738,N_6773,N_7145);
nand U9739 (N_9739,N_6300,N_8687);
nor U9740 (N_9740,N_6850,N_8496);
and U9741 (N_9741,N_6796,N_6464);
xor U9742 (N_9742,N_8168,N_6072);
and U9743 (N_9743,N_8257,N_7026);
nor U9744 (N_9744,N_8146,N_6791);
nand U9745 (N_9745,N_6347,N_8844);
nand U9746 (N_9746,N_7204,N_8796);
nor U9747 (N_9747,N_7320,N_7856);
or U9748 (N_9748,N_8125,N_8950);
and U9749 (N_9749,N_7432,N_8272);
and U9750 (N_9750,N_7171,N_6904);
or U9751 (N_9751,N_8657,N_7391);
xnor U9752 (N_9752,N_8949,N_7588);
nand U9753 (N_9753,N_8226,N_7395);
xnor U9754 (N_9754,N_6818,N_6162);
and U9755 (N_9755,N_6505,N_7266);
and U9756 (N_9756,N_7265,N_7023);
nand U9757 (N_9757,N_8209,N_6498);
nor U9758 (N_9758,N_8640,N_6558);
and U9759 (N_9759,N_7926,N_7824);
or U9760 (N_9760,N_7771,N_8889);
xnor U9761 (N_9761,N_6021,N_6339);
xnor U9762 (N_9762,N_6777,N_6428);
nand U9763 (N_9763,N_7511,N_8062);
or U9764 (N_9764,N_8032,N_7990);
nand U9765 (N_9765,N_6051,N_7673);
nand U9766 (N_9766,N_7235,N_8923);
xnor U9767 (N_9767,N_8681,N_6046);
nor U9768 (N_9768,N_7113,N_7565);
nor U9769 (N_9769,N_7974,N_7707);
xor U9770 (N_9770,N_7316,N_8995);
nor U9771 (N_9771,N_7068,N_7276);
nor U9772 (N_9772,N_8604,N_8221);
nor U9773 (N_9773,N_6972,N_7592);
xor U9774 (N_9774,N_8141,N_6749);
xnor U9775 (N_9775,N_6610,N_7713);
nor U9776 (N_9776,N_8424,N_8386);
nor U9777 (N_9777,N_8912,N_8368);
nand U9778 (N_9778,N_8798,N_8242);
xnor U9779 (N_9779,N_6060,N_8985);
nor U9780 (N_9780,N_7775,N_6152);
nand U9781 (N_9781,N_6379,N_7961);
or U9782 (N_9782,N_6744,N_7797);
nor U9783 (N_9783,N_8071,N_6550);
xor U9784 (N_9784,N_6878,N_6519);
xor U9785 (N_9785,N_8467,N_8370);
nor U9786 (N_9786,N_7942,N_7105);
xor U9787 (N_9787,N_7619,N_6065);
and U9788 (N_9788,N_8590,N_7747);
nor U9789 (N_9789,N_7783,N_7551);
xor U9790 (N_9790,N_6386,N_6540);
nand U9791 (N_9791,N_8601,N_8406);
nand U9792 (N_9792,N_6764,N_6757);
or U9793 (N_9793,N_6090,N_8999);
nor U9794 (N_9794,N_7498,N_6809);
or U9795 (N_9795,N_8435,N_7574);
xor U9796 (N_9796,N_6237,N_7411);
and U9797 (N_9797,N_6154,N_7634);
and U9798 (N_9798,N_8358,N_7857);
or U9799 (N_9799,N_8471,N_6352);
nor U9800 (N_9800,N_6880,N_6779);
nor U9801 (N_9801,N_8402,N_6527);
and U9802 (N_9802,N_6640,N_6691);
and U9803 (N_9803,N_6096,N_8979);
xor U9804 (N_9804,N_7666,N_6942);
xor U9805 (N_9805,N_6995,N_6113);
nand U9806 (N_9806,N_7608,N_7014);
and U9807 (N_9807,N_6897,N_8460);
nand U9808 (N_9808,N_8713,N_6454);
nor U9809 (N_9809,N_6876,N_6747);
or U9810 (N_9810,N_6288,N_8928);
nor U9811 (N_9811,N_8336,N_6740);
xnor U9812 (N_9812,N_6117,N_7273);
nand U9813 (N_9813,N_7271,N_6947);
nor U9814 (N_9814,N_8408,N_8446);
xor U9815 (N_9815,N_8615,N_8488);
or U9816 (N_9816,N_7944,N_6001);
nor U9817 (N_9817,N_8431,N_6970);
xnor U9818 (N_9818,N_8016,N_8490);
nor U9819 (N_9819,N_6275,N_8505);
and U9820 (N_9820,N_8048,N_7689);
or U9821 (N_9821,N_8862,N_6348);
or U9822 (N_9822,N_8156,N_7692);
nand U9823 (N_9823,N_8728,N_6588);
or U9824 (N_9824,N_6227,N_6213);
or U9825 (N_9825,N_7701,N_6315);
nand U9826 (N_9826,N_7173,N_6209);
and U9827 (N_9827,N_6808,N_7595);
xor U9828 (N_9828,N_8396,N_7189);
nor U9829 (N_9829,N_7678,N_6282);
xor U9830 (N_9830,N_8445,N_6111);
nand U9831 (N_9831,N_6120,N_6949);
nand U9832 (N_9832,N_8847,N_7364);
nand U9833 (N_9833,N_6277,N_6555);
and U9834 (N_9834,N_7240,N_6798);
or U9835 (N_9835,N_7363,N_6081);
xor U9836 (N_9836,N_6651,N_7972);
nand U9837 (N_9837,N_8778,N_6383);
or U9838 (N_9838,N_8407,N_6969);
or U9839 (N_9839,N_6401,N_6790);
xor U9840 (N_9840,N_6185,N_7134);
and U9841 (N_9841,N_7377,N_8771);
xor U9842 (N_9842,N_7828,N_7174);
or U9843 (N_9843,N_6622,N_7597);
nor U9844 (N_9844,N_6531,N_6370);
or U9845 (N_9845,N_8745,N_6576);
and U9846 (N_9846,N_8902,N_7281);
nand U9847 (N_9847,N_7580,N_8533);
or U9848 (N_9848,N_7159,N_6922);
nor U9849 (N_9849,N_6486,N_6605);
and U9850 (N_9850,N_8245,N_6161);
nor U9851 (N_9851,N_8437,N_7753);
nand U9852 (N_9852,N_7695,N_6754);
xor U9853 (N_9853,N_7146,N_7270);
or U9854 (N_9854,N_8255,N_7899);
and U9855 (N_9855,N_6278,N_8360);
and U9856 (N_9856,N_8371,N_6812);
nor U9857 (N_9857,N_8265,N_8227);
nand U9858 (N_9858,N_8169,N_6532);
nor U9859 (N_9859,N_7129,N_6881);
nor U9860 (N_9860,N_7975,N_8387);
or U9861 (N_9861,N_6413,N_8773);
or U9862 (N_9862,N_6598,N_8327);
nor U9863 (N_9863,N_8015,N_6177);
nand U9864 (N_9864,N_6896,N_7272);
xor U9865 (N_9865,N_6279,N_6857);
and U9866 (N_9866,N_8667,N_7981);
or U9867 (N_9867,N_6406,N_8462);
xor U9868 (N_9868,N_8268,N_8105);
or U9869 (N_9869,N_7598,N_6954);
xor U9870 (N_9870,N_8389,N_6219);
nand U9871 (N_9871,N_6870,N_7848);
xnor U9872 (N_9872,N_8931,N_7361);
or U9873 (N_9873,N_7740,N_8987);
xor U9874 (N_9874,N_6291,N_6042);
or U9875 (N_9875,N_8662,N_6806);
nand U9876 (N_9876,N_6169,N_6956);
xnor U9877 (N_9877,N_7319,N_8006);
nand U9878 (N_9878,N_6524,N_8639);
nand U9879 (N_9879,N_6095,N_6327);
xor U9880 (N_9880,N_8782,N_8727);
nor U9881 (N_9881,N_8668,N_8555);
nand U9882 (N_9882,N_6369,N_7408);
xor U9883 (N_9883,N_8871,N_8807);
or U9884 (N_9884,N_8945,N_6311);
or U9885 (N_9885,N_6244,N_8731);
nor U9886 (N_9886,N_8981,N_6815);
and U9887 (N_9887,N_7743,N_8161);
nor U9888 (N_9888,N_7850,N_6011);
nor U9889 (N_9889,N_8202,N_6759);
xnor U9890 (N_9890,N_7863,N_8786);
or U9891 (N_9891,N_8315,N_6902);
and U9892 (N_9892,N_6225,N_6460);
and U9893 (N_9893,N_6566,N_7733);
nor U9894 (N_9894,N_8381,N_6212);
nor U9895 (N_9895,N_7390,N_8764);
xnor U9896 (N_9896,N_8200,N_8207);
xor U9897 (N_9897,N_8566,N_7061);
or U9898 (N_9898,N_6589,N_6131);
or U9899 (N_9899,N_6446,N_7075);
and U9900 (N_9900,N_7078,N_8277);
and U9901 (N_9901,N_7905,N_6694);
xor U9902 (N_9902,N_8922,N_7609);
nor U9903 (N_9903,N_6689,N_6998);
and U9904 (N_9904,N_7465,N_8529);
or U9905 (N_9905,N_8919,N_6785);
nor U9906 (N_9906,N_8734,N_7231);
nand U9907 (N_9907,N_8736,N_8869);
nand U9908 (N_9908,N_7560,N_6266);
nor U9909 (N_9909,N_7873,N_6082);
or U9910 (N_9910,N_6996,N_7290);
nor U9911 (N_9911,N_8054,N_8719);
and U9912 (N_9912,N_8854,N_7682);
nor U9913 (N_9913,N_6215,N_7428);
and U9914 (N_9914,N_7261,N_6321);
and U9915 (N_9915,N_6762,N_6193);
nor U9916 (N_9916,N_6294,N_6127);
or U9917 (N_9917,N_6368,N_7183);
or U9918 (N_9918,N_8683,N_7862);
and U9919 (N_9919,N_6033,N_8201);
and U9920 (N_9920,N_8777,N_6700);
and U9921 (N_9921,N_8463,N_6023);
nand U9922 (N_9922,N_7006,N_6537);
or U9923 (N_9923,N_6331,N_6025);
or U9924 (N_9924,N_7593,N_8795);
or U9925 (N_9925,N_7359,N_7339);
and U9926 (N_9926,N_8996,N_6256);
and U9927 (N_9927,N_8609,N_8697);
nor U9928 (N_9928,N_7790,N_7581);
xnor U9929 (N_9929,N_7522,N_8883);
and U9930 (N_9930,N_7766,N_8232);
and U9931 (N_9931,N_6637,N_7166);
nand U9932 (N_9932,N_6685,N_7234);
xnor U9933 (N_9933,N_8448,N_6816);
or U9934 (N_9934,N_8813,N_6593);
nor U9935 (N_9935,N_8170,N_7029);
xnor U9936 (N_9936,N_8078,N_7314);
nand U9937 (N_9937,N_6535,N_6874);
xor U9938 (N_9938,N_8799,N_6358);
nor U9939 (N_9939,N_7752,N_6548);
nor U9940 (N_9940,N_6330,N_8767);
nor U9941 (N_9941,N_7640,N_7194);
nor U9942 (N_9942,N_8441,N_7191);
xor U9943 (N_9943,N_8510,N_6378);
xnor U9944 (N_9944,N_8896,N_8616);
or U9945 (N_9945,N_8392,N_8716);
nor U9946 (N_9946,N_6155,N_6565);
xor U9947 (N_9947,N_8233,N_7526);
nor U9948 (N_9948,N_8196,N_6110);
nor U9949 (N_9949,N_8045,N_7829);
nor U9950 (N_9950,N_8388,N_6041);
nor U9951 (N_9951,N_6353,N_6445);
and U9952 (N_9952,N_6431,N_6784);
and U9953 (N_9953,N_8260,N_7683);
xor U9954 (N_9954,N_6103,N_6141);
nand U9955 (N_9955,N_7715,N_7630);
nor U9956 (N_9956,N_8138,N_8029);
or U9957 (N_9957,N_7663,N_7774);
nor U9958 (N_9958,N_8430,N_6864);
and U9959 (N_9959,N_8647,N_6426);
xor U9960 (N_9960,N_8992,N_7436);
xor U9961 (N_9961,N_6885,N_7671);
and U9962 (N_9962,N_7955,N_8545);
xor U9963 (N_9963,N_7223,N_8890);
xor U9964 (N_9964,N_8057,N_6664);
or U9965 (N_9965,N_6466,N_7157);
xor U9966 (N_9966,N_8439,N_8267);
nand U9967 (N_9967,N_7946,N_8179);
xnor U9968 (N_9968,N_6442,N_6533);
or U9969 (N_9969,N_7197,N_8659);
or U9970 (N_9970,N_6819,N_6343);
xor U9971 (N_9971,N_7190,N_7379);
nand U9972 (N_9972,N_8133,N_7841);
or U9973 (N_9973,N_6844,N_7554);
and U9974 (N_9974,N_6750,N_8741);
nand U9975 (N_9975,N_6621,N_6543);
and U9976 (N_9976,N_6934,N_8599);
and U9977 (N_9977,N_8675,N_7495);
nand U9978 (N_9978,N_6875,N_8903);
nor U9979 (N_9979,N_8788,N_6800);
nor U9980 (N_9980,N_8973,N_6410);
xnor U9981 (N_9981,N_8308,N_7567);
nand U9982 (N_9982,N_7399,N_8729);
and U9983 (N_9983,N_6203,N_8808);
and U9984 (N_9984,N_6399,N_6967);
or U9985 (N_9985,N_8262,N_6988);
or U9986 (N_9986,N_7622,N_6405);
and U9987 (N_9987,N_8825,N_7973);
and U9988 (N_9988,N_6040,N_8975);
nand U9989 (N_9989,N_8300,N_7063);
or U9990 (N_9990,N_8128,N_7782);
nand U9991 (N_9991,N_6984,N_7729);
xnor U9992 (N_9992,N_8497,N_8537);
and U9993 (N_9993,N_8007,N_7139);
xor U9994 (N_9994,N_8936,N_8899);
xor U9995 (N_9995,N_7519,N_6578);
or U9996 (N_9996,N_8988,N_6771);
xnor U9997 (N_9997,N_8502,N_6688);
nor U9998 (N_9998,N_7717,N_7322);
or U9999 (N_9999,N_8739,N_8823);
or U10000 (N_10000,N_7102,N_8937);
xnor U10001 (N_10001,N_7085,N_6281);
nor U10002 (N_10002,N_8352,N_7705);
nor U10003 (N_10003,N_7512,N_6987);
and U10004 (N_10004,N_8461,N_7840);
nand U10005 (N_10005,N_8175,N_7125);
or U10006 (N_10006,N_8059,N_6915);
or U10007 (N_10007,N_8176,N_6057);
and U10008 (N_10008,N_8735,N_8909);
or U10009 (N_10009,N_7796,N_7389);
or U10010 (N_10010,N_7915,N_6848);
or U10011 (N_10011,N_6457,N_7596);
nand U10012 (N_10012,N_6879,N_6597);
and U10013 (N_10013,N_8261,N_6600);
or U10014 (N_10014,N_6965,N_7496);
and U10015 (N_10015,N_8485,N_7871);
or U10016 (N_10016,N_8067,N_6683);
nor U10017 (N_10017,N_8579,N_6380);
nand U10018 (N_10018,N_8036,N_6721);
nor U10019 (N_10019,N_6925,N_8789);
xnor U10020 (N_10020,N_7799,N_8361);
xnor U10021 (N_10021,N_7738,N_8322);
nand U10022 (N_10022,N_7196,N_6810);
or U10023 (N_10023,N_6634,N_8612);
or U10024 (N_10024,N_7422,N_7880);
and U10025 (N_10025,N_6974,N_8761);
and U10026 (N_10026,N_7455,N_7338);
xnor U10027 (N_10027,N_6625,N_7421);
nor U10028 (N_10028,N_8280,N_8298);
or U10029 (N_10029,N_6024,N_8710);
or U10030 (N_10030,N_6828,N_7462);
or U10031 (N_10031,N_7557,N_7920);
nor U10032 (N_10032,N_8977,N_7430);
or U10033 (N_10033,N_6170,N_8810);
or U10034 (N_10034,N_8643,N_6004);
and U10035 (N_10035,N_8183,N_7773);
nor U10036 (N_10036,N_8217,N_6884);
nand U10037 (N_10037,N_8514,N_6701);
and U10038 (N_10038,N_6139,N_7289);
nand U10039 (N_10039,N_6955,N_7300);
nor U10040 (N_10040,N_8594,N_6283);
nor U10041 (N_10041,N_8538,N_8792);
nor U10042 (N_10042,N_8873,N_7846);
nand U10043 (N_10043,N_6035,N_8508);
xor U10044 (N_10044,N_8689,N_8185);
xor U10045 (N_10045,N_7703,N_7872);
nor U10046 (N_10046,N_8507,N_8515);
or U10047 (N_10047,N_8231,N_7082);
nor U10048 (N_10048,N_6462,N_8079);
nand U10049 (N_10049,N_6478,N_6966);
and U10050 (N_10050,N_7483,N_8068);
nand U10051 (N_10051,N_7921,N_8263);
or U10052 (N_10052,N_7706,N_6485);
nand U10053 (N_10053,N_8752,N_8747);
and U10054 (N_10054,N_7402,N_8605);
and U10055 (N_10055,N_8114,N_6075);
and U10056 (N_10056,N_7867,N_6166);
and U10057 (N_10057,N_6873,N_8028);
xnor U10058 (N_10058,N_7380,N_6741);
nand U10059 (N_10059,N_8470,N_6414);
or U10060 (N_10060,N_7248,N_7749);
or U10061 (N_10061,N_6692,N_8958);
xnor U10062 (N_10062,N_7924,N_8610);
xnor U10063 (N_10063,N_8465,N_8583);
xnor U10064 (N_10064,N_8829,N_7999);
nor U10065 (N_10065,N_8243,N_6801);
nor U10066 (N_10066,N_6938,N_7256);
xor U10067 (N_10067,N_8275,N_6789);
and U10068 (N_10068,N_6551,N_8008);
or U10069 (N_10069,N_7153,N_6959);
or U10070 (N_10070,N_6292,N_6499);
nand U10071 (N_10071,N_7108,N_8440);
nand U10072 (N_10072,N_7914,N_6646);
and U10073 (N_10073,N_6299,N_8088);
xor U10074 (N_10074,N_8363,N_6435);
or U10075 (N_10075,N_7657,N_6268);
nand U10076 (N_10076,N_8111,N_7041);
nand U10077 (N_10077,N_8208,N_8117);
and U10078 (N_10078,N_7307,N_7050);
nor U10079 (N_10079,N_8092,N_7460);
or U10080 (N_10080,N_7822,N_6310);
nand U10081 (N_10081,N_8278,N_8817);
xor U10082 (N_10082,N_7306,N_8819);
nor U10083 (N_10083,N_7803,N_8893);
nand U10084 (N_10084,N_8034,N_6708);
or U10085 (N_10085,N_6062,N_6827);
xor U10086 (N_10086,N_7562,N_7523);
xnor U10087 (N_10087,N_7123,N_8299);
nand U10088 (N_10088,N_8365,N_6732);
nand U10089 (N_10089,N_7500,N_7103);
xor U10090 (N_10090,N_8534,N_8560);
or U10091 (N_10091,N_6933,N_7329);
or U10092 (N_10092,N_6665,N_7016);
or U10093 (N_10093,N_8544,N_6782);
nand U10094 (N_10094,N_6666,N_8800);
xnor U10095 (N_10095,N_7414,N_6323);
or U10096 (N_10096,N_7756,N_7252);
or U10097 (N_10097,N_7875,N_8504);
or U10098 (N_10098,N_8434,N_6774);
nor U10099 (N_10099,N_8881,N_7997);
nor U10100 (N_10100,N_8503,N_7263);
or U10101 (N_10101,N_6463,N_8325);
nor U10102 (N_10102,N_6644,N_8289);
xnor U10103 (N_10103,N_7816,N_6039);
and U10104 (N_10104,N_6107,N_6742);
nand U10105 (N_10105,N_8637,N_7296);
and U10106 (N_10106,N_7950,N_8212);
nand U10107 (N_10107,N_8306,N_6118);
xor U10108 (N_10108,N_8246,N_7903);
nand U10109 (N_10109,N_7259,N_7553);
xnor U10110 (N_10110,N_8664,N_7346);
nand U10111 (N_10111,N_7994,N_7488);
nand U10112 (N_10112,N_7877,N_6069);
and U10113 (N_10113,N_7940,N_6186);
and U10114 (N_10114,N_8606,N_7407);
or U10115 (N_10115,N_8760,N_6963);
or U10116 (N_10116,N_8720,N_8206);
xnor U10117 (N_10117,N_7058,N_6050);
and U10118 (N_10118,N_7969,N_7860);
nor U10119 (N_10119,N_7282,N_6930);
and U10120 (N_10120,N_7625,N_7080);
nor U10121 (N_10121,N_6119,N_7935);
or U10122 (N_10122,N_6652,N_8748);
nand U10123 (N_10123,N_6123,N_6739);
or U10124 (N_10124,N_8655,N_7852);
and U10125 (N_10125,N_7218,N_8965);
nor U10126 (N_10126,N_6883,N_7992);
nand U10127 (N_10127,N_6997,N_7215);
nor U10128 (N_10128,N_7073,N_6028);
nand U10129 (N_10129,N_8286,N_8886);
and U10130 (N_10130,N_6363,N_6853);
or U10131 (N_10131,N_7403,N_8809);
nor U10132 (N_10132,N_7548,N_7018);
nor U10133 (N_10133,N_8019,N_7958);
xnor U10134 (N_10134,N_6592,N_6322);
nor U10135 (N_10135,N_7537,N_7454);
nand U10136 (N_10136,N_8056,N_8762);
nand U10137 (N_10137,N_8917,N_7028);
and U10138 (N_10138,N_8860,N_6452);
nor U10139 (N_10139,N_7864,N_6149);
or U10140 (N_10140,N_7954,N_6514);
and U10141 (N_10141,N_6049,N_8314);
xor U10142 (N_10142,N_6184,N_6704);
or U10143 (N_10143,N_6992,N_7600);
nor U10144 (N_10144,N_6231,N_6852);
nor U10145 (N_10145,N_8222,N_7755);
xnor U10146 (N_10146,N_8543,N_7504);
xor U10147 (N_10147,N_8427,N_6000);
xnor U10148 (N_10148,N_6973,N_8080);
and U10149 (N_10149,N_6102,N_7868);
nor U10150 (N_10150,N_8235,N_7778);
nor U10151 (N_10151,N_6891,N_8614);
nor U10152 (N_10152,N_8478,N_7344);
nand U10153 (N_10153,N_7000,N_8102);
and U10154 (N_10154,N_8607,N_7095);
or U10155 (N_10155,N_6506,N_6559);
nor U10156 (N_10156,N_8691,N_8182);
nor U10157 (N_10157,N_8863,N_8541);
xnor U10158 (N_10158,N_8137,N_7137);
nand U10159 (N_10159,N_7180,N_7337);
nor U10160 (N_10160,N_8096,N_8712);
and U10161 (N_10161,N_7610,N_7008);
nand U10162 (N_10162,N_7244,N_7665);
nand U10163 (N_10163,N_7702,N_8641);
nor U10164 (N_10164,N_7287,N_7340);
and U10165 (N_10165,N_6983,N_6415);
nor U10166 (N_10166,N_6236,N_6026);
and U10167 (N_10167,N_6895,N_6003);
nand U10168 (N_10168,N_6391,N_8707);
and U10169 (N_10169,N_7356,N_6205);
and U10170 (N_10170,N_6536,N_8787);
nand U10171 (N_10171,N_6218,N_6624);
xnor U10172 (N_10172,N_8266,N_7445);
nor U10173 (N_10173,N_6921,N_8244);
or U10174 (N_10174,N_8230,N_7416);
and U10175 (N_10175,N_8851,N_8611);
xor U10176 (N_10176,N_8095,N_8780);
and U10177 (N_10177,N_8451,N_6375);
nor U10178 (N_10178,N_8037,N_6269);
or U10179 (N_10179,N_8348,N_6180);
nand U10180 (N_10180,N_6453,N_7089);
nor U10181 (N_10181,N_6362,N_8723);
or U10182 (N_10182,N_6472,N_7965);
nand U10183 (N_10183,N_7114,N_8145);
nand U10184 (N_10184,N_8393,N_6138);
nor U10185 (N_10185,N_8914,N_8473);
or U10186 (N_10186,N_6687,N_6455);
nor U10187 (N_10187,N_7140,N_6234);
nor U10188 (N_10188,N_7677,N_8160);
nand U10189 (N_10189,N_6924,N_8309);
or U10190 (N_10190,N_6613,N_7884);
xor U10191 (N_10191,N_7368,N_6015);
xnor U10192 (N_10192,N_6570,N_7952);
and U10193 (N_10193,N_8517,N_7161);
nand U10194 (N_10194,N_6950,N_7821);
and U10195 (N_10195,N_8291,N_8066);
and U10196 (N_10196,N_7651,N_8324);
or U10197 (N_10197,N_6295,N_7977);
or U10198 (N_10198,N_6690,N_6607);
nand U10199 (N_10199,N_8332,N_6528);
or U10200 (N_10200,N_8310,N_6458);
or U10201 (N_10201,N_8184,N_7525);
and U10202 (N_10202,N_7131,N_7274);
or U10203 (N_10203,N_8846,N_8155);
nand U10204 (N_10204,N_7826,N_8906);
nand U10205 (N_10205,N_8270,N_6114);
nand U10206 (N_10206,N_8938,N_6249);
and U10207 (N_10207,N_8065,N_8715);
xor U10208 (N_10208,N_7658,N_7656);
xor U10209 (N_10209,N_7217,N_8820);
nand U10210 (N_10210,N_6923,N_7943);
nor U10211 (N_10211,N_7572,N_6443);
nand U10212 (N_10212,N_7853,N_6728);
and U10213 (N_10213,N_7321,N_7911);
or U10214 (N_10214,N_7607,N_8648);
and U10215 (N_10215,N_8301,N_8947);
or U10216 (N_10216,N_7458,N_8253);
and U10217 (N_10217,N_7199,N_7192);
or U10218 (N_10218,N_7477,N_6905);
or U10219 (N_10219,N_8220,N_6860);
or U10220 (N_10220,N_8574,N_6960);
nand U10221 (N_10221,N_6329,N_6438);
nand U10222 (N_10222,N_7886,N_7253);
xnor U10223 (N_10223,N_8326,N_7830);
nand U10224 (N_10224,N_6877,N_8256);
nor U10225 (N_10225,N_8038,N_8069);
xnor U10226 (N_10226,N_7583,N_8750);
and U10227 (N_10227,N_7785,N_7586);
nand U10228 (N_10228,N_7838,N_7237);
nand U10229 (N_10229,N_7576,N_8831);
xor U10230 (N_10230,N_7660,N_6332);
xor U10231 (N_10231,N_6941,N_7744);
xnor U10232 (N_10232,N_6917,N_6693);
or U10233 (N_10233,N_8932,N_8960);
xor U10234 (N_10234,N_7167,N_6230);
nand U10235 (N_10235,N_8843,N_7466);
nor U10236 (N_10236,N_8584,N_8240);
and U10237 (N_10237,N_7154,N_6907);
xor U10238 (N_10238,N_7646,N_7505);
nor U10239 (N_10239,N_7670,N_6914);
nand U10240 (N_10240,N_6989,N_7444);
nor U10241 (N_10241,N_8123,N_8011);
and U10242 (N_10242,N_6697,N_6450);
nand U10243 (N_10243,N_8709,N_8845);
xnor U10244 (N_10244,N_7124,N_7542);
nor U10245 (N_10245,N_8586,N_8530);
nand U10246 (N_10246,N_6746,N_6936);
and U10247 (N_10247,N_8165,N_7177);
and U10248 (N_10248,N_6319,N_8524);
nor U10249 (N_10249,N_6534,N_7047);
and U10250 (N_10250,N_6556,N_7900);
and U10251 (N_10251,N_7392,N_6017);
or U10252 (N_10252,N_8113,N_6421);
or U10253 (N_10253,N_6829,N_7438);
nand U10254 (N_10254,N_6208,N_6016);
xor U10255 (N_10255,N_8195,N_7442);
nand U10256 (N_10256,N_8805,N_7893);
or U10257 (N_10257,N_6780,N_8091);
or U10258 (N_10258,N_6968,N_8093);
nand U10259 (N_10259,N_8711,N_6221);
or U10260 (N_10260,N_6371,N_8758);
nand U10261 (N_10261,N_6153,N_6510);
and U10262 (N_10262,N_6603,N_7334);
xor U10263 (N_10263,N_6994,N_8673);
nand U10264 (N_10264,N_7759,N_6194);
and U10265 (N_10265,N_6525,N_8236);
and U10266 (N_10266,N_7866,N_6429);
and U10267 (N_10267,N_6388,N_8044);
xor U10268 (N_10268,N_6937,N_7823);
xor U10269 (N_10269,N_7366,N_7813);
nor U10270 (N_10270,N_7048,N_6128);
or U10271 (N_10271,N_7258,N_6575);
nor U10272 (N_10272,N_7092,N_7662);
xnor U10273 (N_10273,N_6635,N_8142);
or U10274 (N_10274,N_8832,N_7010);
or U10275 (N_10275,N_8130,N_7587);
nand U10276 (N_10276,N_7517,N_8700);
nor U10277 (N_10277,N_7869,N_7575);
nand U10278 (N_10278,N_7948,N_7370);
nor U10279 (N_10279,N_7093,N_8023);
or U10280 (N_10280,N_6522,N_6226);
nand U10281 (N_10281,N_6043,N_8073);
or U10282 (N_10282,N_8344,N_6179);
xnor U10283 (N_10283,N_7801,N_7642);
nand U10284 (N_10284,N_7844,N_7641);
and U10285 (N_10285,N_6571,N_8025);
or U10286 (N_10286,N_6730,N_6031);
and U10287 (N_10287,N_7945,N_7601);
nor U10288 (N_10288,N_6751,N_6753);
nor U10289 (N_10289,N_7644,N_7053);
nand U10290 (N_10290,N_8626,N_6433);
or U10291 (N_10291,N_6143,N_8443);
and U10292 (N_10292,N_6247,N_6303);
or U10293 (N_10293,N_7176,N_7748);
nor U10294 (N_10294,N_6228,N_7353);
or U10295 (N_10295,N_8532,N_6146);
or U10296 (N_10296,N_7781,N_7524);
nand U10297 (N_10297,N_6716,N_8323);
nor U10298 (N_10298,N_8790,N_8522);
nand U10299 (N_10299,N_7164,N_7979);
xor U10300 (N_10300,N_8672,N_7086);
or U10301 (N_10301,N_7654,N_6192);
or U10302 (N_10302,N_8920,N_8523);
nand U10303 (N_10303,N_6958,N_6932);
xnor U10304 (N_10304,N_6839,N_8986);
nor U10305 (N_10305,N_7571,N_8765);
nand U10306 (N_10306,N_7452,N_7294);
nand U10307 (N_10307,N_7831,N_6500);
nand U10308 (N_10308,N_8644,N_7076);
nand U10309 (N_10309,N_6908,N_6752);
nand U10310 (N_10310,N_6776,N_6835);
nand U10311 (N_10311,N_7071,N_8563);
and U10312 (N_10312,N_7479,N_7925);
or U10313 (N_10313,N_7898,N_6390);
nor U10314 (N_10314,N_6760,N_6222);
xor U10315 (N_10315,N_7694,N_8391);
nand U10316 (N_10316,N_6781,N_7417);
nand U10317 (N_10317,N_8682,N_7437);
xnor U10318 (N_10318,N_7772,N_7614);
and U10319 (N_10319,N_6502,N_6059);
nor U10320 (N_10320,N_6145,N_8842);
or U10321 (N_10321,N_8494,N_7686);
nand U10322 (N_10322,N_7808,N_8897);
and U10323 (N_10323,N_6314,N_6381);
nand U10324 (N_10324,N_8003,N_7843);
xnor U10325 (N_10325,N_6479,N_6542);
xor U10326 (N_10326,N_7764,N_7015);
or U10327 (N_10327,N_6097,N_8000);
and U10328 (N_10328,N_6325,N_8801);
or U10329 (N_10329,N_6766,N_6561);
nand U10330 (N_10330,N_8653,N_8347);
nand U10331 (N_10331,N_6087,N_8991);
nand U10332 (N_10332,N_7087,N_7507);
nand U10333 (N_10333,N_6993,N_8481);
or U10334 (N_10334,N_8269,N_6328);
nor U10335 (N_10335,N_6991,N_7928);
or U10336 (N_10336,N_6630,N_7278);
xnor U10337 (N_10337,N_8118,N_8806);
or U10338 (N_10338,N_6468,N_7170);
and U10339 (N_10339,N_6882,N_8229);
nor U10340 (N_10340,N_6037,N_6197);
xnor U10341 (N_10341,N_7855,N_7323);
and U10342 (N_10342,N_7604,N_6820);
xor U10343 (N_10343,N_7107,N_8918);
and U10344 (N_10344,N_7514,N_6583);
xor U10345 (N_10345,N_7470,N_7027);
xor U10346 (N_10346,N_7135,N_6541);
and U10347 (N_10347,N_7345,N_8378);
xor U10348 (N_10348,N_7489,N_7298);
xor U10349 (N_10349,N_8692,N_7652);
or U10350 (N_10350,N_6271,N_6786);
nand U10351 (N_10351,N_7213,N_7098);
and U10352 (N_10352,N_7627,N_7162);
nor U10353 (N_10353,N_8046,N_7888);
nor U10354 (N_10354,N_7736,N_8162);
and U10355 (N_10355,N_8404,N_6364);
or U10356 (N_10356,N_8618,N_8180);
or U10357 (N_10357,N_8840,N_7931);
nor U10358 (N_10358,N_8603,N_6946);
nor U10359 (N_10359,N_6961,N_7055);
or U10360 (N_10360,N_6626,N_8241);
xnor U10361 (N_10361,N_6309,N_6359);
and U10362 (N_10362,N_7552,N_6189);
xnor U10363 (N_10363,N_8340,N_6484);
xor U10364 (N_10364,N_7032,N_6686);
nor U10365 (N_10365,N_7556,N_7031);
or U10366 (N_10366,N_6471,N_8273);
or U10367 (N_10367,N_6239,N_8518);
nor U10368 (N_10368,N_7916,N_7910);
or U10369 (N_10369,N_7953,N_7832);
xor U10370 (N_10370,N_6009,N_6833);
or U10371 (N_10371,N_7988,N_6641);
and U10372 (N_10372,N_7700,N_8420);
or U10373 (N_10373,N_7962,N_6726);
nor U10374 (N_10374,N_7594,N_8337);
or U10375 (N_10375,N_6267,N_6795);
and U10376 (N_10376,N_6718,N_7714);
or U10377 (N_10377,N_6832,N_6200);
or U10378 (N_10378,N_8211,N_8276);
nor U10379 (N_10379,N_6673,N_6423);
nand U10380 (N_10380,N_6126,N_6627);
xor U10381 (N_10381,N_6430,N_7543);
xnor U10382 (N_10382,N_6569,N_8094);
xor U10383 (N_10383,N_6196,N_6349);
nand U10384 (N_10384,N_7471,N_7118);
and U10385 (N_10385,N_7245,N_7374);
nand U10386 (N_10386,N_8487,N_7349);
nand U10387 (N_10387,N_7787,N_6407);
nor U10388 (N_10388,N_7393,N_6389);
xnor U10389 (N_10389,N_7688,N_8652);
and U10390 (N_10390,N_8774,N_6733);
or U10391 (N_10391,N_7882,N_7561);
or U10392 (N_10392,N_6223,N_7243);
xor U10393 (N_10393,N_7936,N_8901);
and U10394 (N_10394,N_8385,N_6099);
nand U10395 (N_10395,N_8582,N_8956);
nor U10396 (N_10396,N_8294,N_6296);
and U10397 (N_10397,N_6982,N_6553);
nor U10398 (N_10398,N_8109,N_6076);
nand U10399 (N_10399,N_7317,N_6306);
nor U10400 (N_10400,N_7876,N_7757);
and U10401 (N_10401,N_7727,N_6163);
xnor U10402 (N_10402,N_8974,N_7045);
nor U10403 (N_10403,N_7836,N_6599);
nor U10404 (N_10404,N_7476,N_7019);
or U10405 (N_10405,N_8414,N_7305);
xnor U10406 (N_10406,N_7081,N_7897);
and U10407 (N_10407,N_7745,N_8759);
nor U10408 (N_10408,N_7116,N_7009);
or U10409 (N_10409,N_7956,N_7117);
or U10410 (N_10410,N_6574,N_6338);
nor U10411 (N_10411,N_6094,N_8669);
or U10412 (N_10412,N_7011,N_6521);
xor U10413 (N_10413,N_8702,N_6837);
nand U10414 (N_10414,N_7545,N_8506);
nand U10415 (N_10415,N_8342,N_7236);
and U10416 (N_10416,N_7494,N_7859);
xnor U10417 (N_10417,N_6012,N_8600);
or U10418 (N_10418,N_6412,N_7983);
nand U10419 (N_10419,N_6756,N_6284);
or U10420 (N_10420,N_7106,N_8454);
xnor U10421 (N_10421,N_7612,N_6470);
nand U10422 (N_10422,N_7649,N_7904);
nand U10423 (N_10423,N_7037,N_7351);
nand U10424 (N_10424,N_6656,N_8313);
xnor U10425 (N_10425,N_8218,N_7020);
nand U10426 (N_10426,N_7195,N_6587);
or U10427 (N_10427,N_7762,N_7226);
and U10428 (N_10428,N_6675,N_6387);
nand U10429 (N_10429,N_8921,N_6301);
nor U10430 (N_10430,N_6083,N_8907);
and U10431 (N_10431,N_8622,N_6188);
or U10432 (N_10432,N_6515,N_6986);
nor U10433 (N_10433,N_6802,N_7072);
nor U10434 (N_10434,N_8550,N_7439);
or U10435 (N_10435,N_6518,N_8589);
nand U10436 (N_10436,N_7520,N_8247);
nand U10437 (N_10437,N_8279,N_8190);
nor U10438 (N_10438,N_8763,N_7499);
and U10439 (N_10439,N_6147,N_6745);
nor U10440 (N_10440,N_8721,N_7111);
nand U10441 (N_10441,N_7330,N_7835);
nand U10442 (N_10442,N_8980,N_8959);
or U10443 (N_10443,N_6538,N_8163);
nor U10444 (N_10444,N_6497,N_6660);
or U10445 (N_10445,N_7419,N_6620);
xor U10446 (N_10446,N_6650,N_8567);
nor U10447 (N_10447,N_7040,N_6403);
xnor U10448 (N_10448,N_8837,N_6978);
nor U10449 (N_10449,N_6717,N_7005);
and U10450 (N_10450,N_6132,N_6093);
or U10451 (N_10451,N_7760,N_7486);
xor U10452 (N_10452,N_7804,N_7589);
or U10453 (N_10453,N_6909,N_6427);
and U10454 (N_10454,N_7758,N_8345);
nand U10455 (N_10455,N_8458,N_8880);
nand U10456 (N_10456,N_6312,N_8944);
or U10457 (N_10457,N_6677,N_8106);
or U10458 (N_10458,N_6481,N_7358);
nand U10459 (N_10459,N_7515,N_6036);
and U10460 (N_10460,N_8531,N_7420);
and U10461 (N_10461,N_6669,N_8349);
and U10462 (N_10462,N_8250,N_6106);
nand U10463 (N_10463,N_6703,N_8695);
nand U10464 (N_10464,N_6489,N_8882);
and U10465 (N_10465,N_7158,N_6280);
and U10466 (N_10466,N_6441,N_7516);
nand U10467 (N_10467,N_6272,N_6105);
nand U10468 (N_10468,N_7631,N_7178);
or U10469 (N_10469,N_8967,N_6657);
nand U10470 (N_10470,N_8489,N_6805);
and U10471 (N_10471,N_6027,N_8258);
nor U10472 (N_10472,N_6047,N_7456);
xnor U10473 (N_10473,N_6516,N_6167);
xnor U10474 (N_10474,N_7780,N_8398);
nor U10475 (N_10475,N_7357,N_6552);
or U10476 (N_10476,N_7434,N_8577);
nand U10477 (N_10477,N_6232,N_7615);
or U10478 (N_10478,N_8933,N_8994);
or U10479 (N_10479,N_8362,N_7221);
and U10480 (N_10480,N_7605,N_6243);
xnor U10481 (N_10481,N_6018,N_7255);
nand U10482 (N_10482,N_8671,N_7227);
and U10483 (N_10483,N_8656,N_7789);
nor U10484 (N_10484,N_8976,N_6061);
or U10485 (N_10485,N_6608,N_7286);
and U10486 (N_10486,N_8164,N_7188);
or U10487 (N_10487,N_8271,N_8254);
nor U10488 (N_10488,N_8132,N_8433);
and U10489 (N_10489,N_8198,N_8112);
and U10490 (N_10490,N_7805,N_6979);
or U10491 (N_10491,N_7902,N_8877);
nand U10492 (N_10492,N_8055,N_6467);
or U10493 (N_10493,N_7776,N_6775);
and U10494 (N_10494,N_6682,N_6851);
and U10495 (N_10495,N_7179,N_8086);
or U10496 (N_10496,N_8090,N_6529);
nand U10497 (N_10497,N_8452,N_6520);
and U10498 (N_10498,N_8035,N_7669);
nand U10499 (N_10499,N_7410,N_8570);
nand U10500 (N_10500,N_7442,N_7246);
nor U10501 (N_10501,N_8029,N_6507);
nor U10502 (N_10502,N_6495,N_7415);
xnor U10503 (N_10503,N_8266,N_6600);
and U10504 (N_10504,N_7741,N_8013);
or U10505 (N_10505,N_6693,N_8004);
or U10506 (N_10506,N_7631,N_8117);
and U10507 (N_10507,N_6829,N_8305);
and U10508 (N_10508,N_7105,N_6182);
nor U10509 (N_10509,N_6837,N_8630);
or U10510 (N_10510,N_6198,N_6891);
or U10511 (N_10511,N_7507,N_8801);
nor U10512 (N_10512,N_8310,N_6591);
xnor U10513 (N_10513,N_8898,N_8283);
xnor U10514 (N_10514,N_6859,N_8774);
or U10515 (N_10515,N_8213,N_6190);
or U10516 (N_10516,N_8170,N_6075);
or U10517 (N_10517,N_8285,N_7122);
nor U10518 (N_10518,N_8583,N_8396);
nor U10519 (N_10519,N_8862,N_6450);
nor U10520 (N_10520,N_7982,N_6645);
nand U10521 (N_10521,N_6464,N_7760);
xor U10522 (N_10522,N_7876,N_8598);
and U10523 (N_10523,N_7985,N_6439);
and U10524 (N_10524,N_8077,N_8308);
nor U10525 (N_10525,N_8143,N_8961);
or U10526 (N_10526,N_6910,N_7458);
nand U10527 (N_10527,N_7850,N_6433);
xnor U10528 (N_10528,N_8264,N_6839);
nand U10529 (N_10529,N_7356,N_6557);
or U10530 (N_10530,N_7005,N_7681);
nand U10531 (N_10531,N_8696,N_6125);
xnor U10532 (N_10532,N_6093,N_7980);
nor U10533 (N_10533,N_8639,N_7501);
and U10534 (N_10534,N_8637,N_6088);
nand U10535 (N_10535,N_7155,N_7093);
or U10536 (N_10536,N_6254,N_7054);
or U10537 (N_10537,N_7647,N_6381);
nand U10538 (N_10538,N_6009,N_6283);
nand U10539 (N_10539,N_7531,N_6927);
and U10540 (N_10540,N_8425,N_8065);
xnor U10541 (N_10541,N_7638,N_7824);
or U10542 (N_10542,N_8451,N_7941);
or U10543 (N_10543,N_6714,N_7339);
nand U10544 (N_10544,N_6895,N_8771);
nand U10545 (N_10545,N_6252,N_8617);
or U10546 (N_10546,N_8740,N_8561);
or U10547 (N_10547,N_6278,N_8446);
nor U10548 (N_10548,N_7630,N_6739);
xor U10549 (N_10549,N_8084,N_7360);
nand U10550 (N_10550,N_7300,N_6387);
and U10551 (N_10551,N_7863,N_6384);
nand U10552 (N_10552,N_7090,N_8979);
or U10553 (N_10553,N_6435,N_7961);
xor U10554 (N_10554,N_8738,N_6090);
xnor U10555 (N_10555,N_6878,N_8911);
or U10556 (N_10556,N_8575,N_6212);
nand U10557 (N_10557,N_7504,N_7300);
and U10558 (N_10558,N_8155,N_7903);
nor U10559 (N_10559,N_6924,N_6135);
and U10560 (N_10560,N_6916,N_6918);
or U10561 (N_10561,N_8868,N_8049);
nand U10562 (N_10562,N_7057,N_7574);
nand U10563 (N_10563,N_8482,N_6534);
xnor U10564 (N_10564,N_6063,N_6751);
nand U10565 (N_10565,N_6397,N_7222);
xor U10566 (N_10566,N_7923,N_8258);
or U10567 (N_10567,N_6332,N_7248);
xnor U10568 (N_10568,N_8124,N_7414);
xnor U10569 (N_10569,N_6540,N_7554);
xnor U10570 (N_10570,N_8937,N_7078);
nor U10571 (N_10571,N_6696,N_6091);
and U10572 (N_10572,N_8543,N_7303);
and U10573 (N_10573,N_8559,N_6311);
nand U10574 (N_10574,N_7132,N_6386);
and U10575 (N_10575,N_6865,N_7926);
nand U10576 (N_10576,N_8107,N_6301);
xnor U10577 (N_10577,N_7659,N_8823);
xor U10578 (N_10578,N_8083,N_6570);
and U10579 (N_10579,N_6592,N_7253);
and U10580 (N_10580,N_7549,N_8604);
or U10581 (N_10581,N_8822,N_6425);
and U10582 (N_10582,N_7511,N_6560);
or U10583 (N_10583,N_8657,N_7229);
and U10584 (N_10584,N_7443,N_8020);
or U10585 (N_10585,N_7804,N_6377);
or U10586 (N_10586,N_6646,N_6099);
nand U10587 (N_10587,N_8991,N_8921);
and U10588 (N_10588,N_6020,N_6208);
and U10589 (N_10589,N_8803,N_8594);
and U10590 (N_10590,N_7491,N_8253);
nor U10591 (N_10591,N_7836,N_7357);
nor U10592 (N_10592,N_7609,N_6660);
or U10593 (N_10593,N_6066,N_6912);
nor U10594 (N_10594,N_8050,N_6525);
and U10595 (N_10595,N_6669,N_6488);
xor U10596 (N_10596,N_6065,N_8549);
nand U10597 (N_10597,N_7213,N_8255);
and U10598 (N_10598,N_7944,N_7759);
and U10599 (N_10599,N_6059,N_7801);
and U10600 (N_10600,N_6491,N_8085);
nor U10601 (N_10601,N_8494,N_7369);
xnor U10602 (N_10602,N_7112,N_8252);
nor U10603 (N_10603,N_7554,N_8016);
or U10604 (N_10604,N_7581,N_6943);
or U10605 (N_10605,N_8800,N_7862);
and U10606 (N_10606,N_6960,N_6955);
nor U10607 (N_10607,N_6953,N_6072);
or U10608 (N_10608,N_6036,N_8452);
nand U10609 (N_10609,N_6001,N_6583);
nand U10610 (N_10610,N_6024,N_7870);
nor U10611 (N_10611,N_6870,N_6245);
and U10612 (N_10612,N_7156,N_6303);
and U10613 (N_10613,N_7106,N_8076);
or U10614 (N_10614,N_7019,N_6544);
nor U10615 (N_10615,N_8115,N_8031);
and U10616 (N_10616,N_7648,N_6975);
nand U10617 (N_10617,N_6464,N_7789);
nor U10618 (N_10618,N_8217,N_6717);
nor U10619 (N_10619,N_6475,N_7131);
nor U10620 (N_10620,N_7095,N_6920);
nor U10621 (N_10621,N_8439,N_8519);
and U10622 (N_10622,N_8659,N_7638);
and U10623 (N_10623,N_8681,N_6510);
nor U10624 (N_10624,N_8261,N_8404);
xnor U10625 (N_10625,N_7412,N_7441);
and U10626 (N_10626,N_8796,N_7674);
nor U10627 (N_10627,N_6196,N_6796);
nor U10628 (N_10628,N_7916,N_6632);
nand U10629 (N_10629,N_8630,N_8202);
nor U10630 (N_10630,N_8591,N_6266);
and U10631 (N_10631,N_7502,N_7827);
or U10632 (N_10632,N_6605,N_6806);
or U10633 (N_10633,N_6601,N_8453);
nor U10634 (N_10634,N_8854,N_6634);
nand U10635 (N_10635,N_8465,N_8407);
or U10636 (N_10636,N_7218,N_6895);
xor U10637 (N_10637,N_7932,N_8899);
nand U10638 (N_10638,N_8082,N_7743);
nor U10639 (N_10639,N_7587,N_7821);
nor U10640 (N_10640,N_7561,N_7330);
nor U10641 (N_10641,N_6276,N_7897);
nand U10642 (N_10642,N_6727,N_6215);
nor U10643 (N_10643,N_6478,N_8691);
xor U10644 (N_10644,N_8123,N_7855);
xnor U10645 (N_10645,N_7621,N_7025);
nor U10646 (N_10646,N_6074,N_7271);
nand U10647 (N_10647,N_7347,N_6010);
nand U10648 (N_10648,N_6503,N_8568);
and U10649 (N_10649,N_7136,N_6267);
xnor U10650 (N_10650,N_6907,N_7812);
nand U10651 (N_10651,N_8703,N_6005);
nand U10652 (N_10652,N_8104,N_8588);
xnor U10653 (N_10653,N_6804,N_8485);
nand U10654 (N_10654,N_8456,N_7000);
nor U10655 (N_10655,N_7711,N_6241);
nand U10656 (N_10656,N_8052,N_7797);
xor U10657 (N_10657,N_6212,N_8034);
nor U10658 (N_10658,N_7109,N_6459);
xor U10659 (N_10659,N_6283,N_7901);
nand U10660 (N_10660,N_7145,N_7140);
nor U10661 (N_10661,N_8046,N_6414);
and U10662 (N_10662,N_8598,N_7751);
nor U10663 (N_10663,N_6703,N_6456);
or U10664 (N_10664,N_6334,N_8108);
nand U10665 (N_10665,N_8685,N_6014);
and U10666 (N_10666,N_8619,N_6068);
xnor U10667 (N_10667,N_6483,N_6445);
and U10668 (N_10668,N_6542,N_6506);
or U10669 (N_10669,N_7342,N_7319);
or U10670 (N_10670,N_7775,N_6524);
and U10671 (N_10671,N_7059,N_7946);
and U10672 (N_10672,N_8907,N_7697);
xnor U10673 (N_10673,N_6922,N_6950);
nor U10674 (N_10674,N_7903,N_6247);
nand U10675 (N_10675,N_7970,N_7883);
and U10676 (N_10676,N_7025,N_8173);
xor U10677 (N_10677,N_6892,N_6423);
or U10678 (N_10678,N_8276,N_6211);
nor U10679 (N_10679,N_8234,N_7775);
nor U10680 (N_10680,N_8251,N_6578);
xnor U10681 (N_10681,N_7513,N_7191);
and U10682 (N_10682,N_8639,N_7412);
nand U10683 (N_10683,N_7668,N_6665);
nor U10684 (N_10684,N_7983,N_8265);
nand U10685 (N_10685,N_7244,N_6750);
or U10686 (N_10686,N_7534,N_8728);
and U10687 (N_10687,N_7171,N_6844);
or U10688 (N_10688,N_7114,N_7355);
and U10689 (N_10689,N_8781,N_7929);
or U10690 (N_10690,N_6247,N_8080);
nor U10691 (N_10691,N_8823,N_8483);
and U10692 (N_10692,N_6048,N_6307);
or U10693 (N_10693,N_6635,N_6606);
and U10694 (N_10694,N_8134,N_8973);
xnor U10695 (N_10695,N_6002,N_6975);
or U10696 (N_10696,N_6516,N_6538);
and U10697 (N_10697,N_7885,N_8805);
xor U10698 (N_10698,N_8976,N_8187);
and U10699 (N_10699,N_6615,N_6733);
and U10700 (N_10700,N_8757,N_6412);
xor U10701 (N_10701,N_8162,N_6865);
or U10702 (N_10702,N_8022,N_8849);
nand U10703 (N_10703,N_7159,N_6442);
nor U10704 (N_10704,N_6999,N_8649);
or U10705 (N_10705,N_8204,N_6710);
xnor U10706 (N_10706,N_6505,N_7052);
nor U10707 (N_10707,N_8889,N_6346);
or U10708 (N_10708,N_7588,N_6774);
or U10709 (N_10709,N_8341,N_6864);
nor U10710 (N_10710,N_8785,N_8852);
nand U10711 (N_10711,N_7551,N_6906);
or U10712 (N_10712,N_8250,N_8071);
and U10713 (N_10713,N_8108,N_8406);
or U10714 (N_10714,N_7151,N_6654);
xnor U10715 (N_10715,N_7045,N_7517);
and U10716 (N_10716,N_8840,N_6843);
nor U10717 (N_10717,N_7040,N_6569);
nor U10718 (N_10718,N_7653,N_8987);
nor U10719 (N_10719,N_7759,N_6771);
nand U10720 (N_10720,N_8767,N_6500);
or U10721 (N_10721,N_8644,N_6490);
or U10722 (N_10722,N_6552,N_6966);
and U10723 (N_10723,N_6745,N_6624);
or U10724 (N_10724,N_6443,N_6535);
nand U10725 (N_10725,N_8031,N_7094);
and U10726 (N_10726,N_6746,N_8000);
nand U10727 (N_10727,N_7323,N_7937);
or U10728 (N_10728,N_7723,N_8874);
nor U10729 (N_10729,N_6814,N_7961);
nand U10730 (N_10730,N_6642,N_7565);
nand U10731 (N_10731,N_6288,N_8140);
or U10732 (N_10732,N_6728,N_8524);
nor U10733 (N_10733,N_7368,N_7890);
or U10734 (N_10734,N_6017,N_7691);
xor U10735 (N_10735,N_6947,N_8623);
nand U10736 (N_10736,N_7613,N_6512);
xnor U10737 (N_10737,N_7458,N_6753);
and U10738 (N_10738,N_8669,N_7751);
nand U10739 (N_10739,N_8178,N_7181);
nand U10740 (N_10740,N_7976,N_7022);
xor U10741 (N_10741,N_8266,N_7891);
xnor U10742 (N_10742,N_7881,N_7929);
nand U10743 (N_10743,N_7780,N_8574);
and U10744 (N_10744,N_8829,N_7484);
xor U10745 (N_10745,N_8745,N_7698);
or U10746 (N_10746,N_6397,N_7216);
and U10747 (N_10747,N_7022,N_6486);
xnor U10748 (N_10748,N_7526,N_7535);
and U10749 (N_10749,N_7246,N_8611);
nand U10750 (N_10750,N_7061,N_7491);
or U10751 (N_10751,N_6513,N_8769);
xor U10752 (N_10752,N_6959,N_7869);
or U10753 (N_10753,N_7749,N_7230);
nand U10754 (N_10754,N_6667,N_8786);
xnor U10755 (N_10755,N_6544,N_6280);
nand U10756 (N_10756,N_8845,N_7763);
and U10757 (N_10757,N_7792,N_8181);
or U10758 (N_10758,N_6966,N_7089);
and U10759 (N_10759,N_7253,N_6600);
and U10760 (N_10760,N_7185,N_8858);
nor U10761 (N_10761,N_8658,N_6810);
or U10762 (N_10762,N_8577,N_7601);
or U10763 (N_10763,N_6601,N_7636);
or U10764 (N_10764,N_8519,N_6853);
nor U10765 (N_10765,N_6380,N_8469);
or U10766 (N_10766,N_7463,N_7715);
nor U10767 (N_10767,N_8654,N_6522);
nor U10768 (N_10768,N_7135,N_8935);
nand U10769 (N_10769,N_8632,N_6444);
nor U10770 (N_10770,N_6509,N_7090);
xor U10771 (N_10771,N_8250,N_8231);
and U10772 (N_10772,N_8812,N_8912);
and U10773 (N_10773,N_8994,N_8540);
and U10774 (N_10774,N_7099,N_7607);
nor U10775 (N_10775,N_6271,N_6420);
and U10776 (N_10776,N_7300,N_7490);
or U10777 (N_10777,N_6280,N_8415);
or U10778 (N_10778,N_6755,N_6501);
and U10779 (N_10779,N_6782,N_8785);
and U10780 (N_10780,N_7744,N_7286);
xor U10781 (N_10781,N_7314,N_7161);
xor U10782 (N_10782,N_6524,N_8768);
and U10783 (N_10783,N_6525,N_7308);
and U10784 (N_10784,N_7336,N_7839);
nor U10785 (N_10785,N_7834,N_8915);
and U10786 (N_10786,N_8157,N_8271);
nor U10787 (N_10787,N_7911,N_7105);
nor U10788 (N_10788,N_6495,N_6236);
and U10789 (N_10789,N_6217,N_6009);
nand U10790 (N_10790,N_8976,N_6931);
nor U10791 (N_10791,N_7286,N_7358);
nand U10792 (N_10792,N_8738,N_8541);
or U10793 (N_10793,N_8090,N_7801);
nand U10794 (N_10794,N_6941,N_7394);
or U10795 (N_10795,N_6384,N_6060);
and U10796 (N_10796,N_6481,N_6485);
nor U10797 (N_10797,N_6198,N_6112);
or U10798 (N_10798,N_8686,N_7841);
or U10799 (N_10799,N_6419,N_8234);
xnor U10800 (N_10800,N_6856,N_8161);
nor U10801 (N_10801,N_6386,N_7340);
or U10802 (N_10802,N_7812,N_8147);
nand U10803 (N_10803,N_7086,N_6558);
and U10804 (N_10804,N_6594,N_7606);
nor U10805 (N_10805,N_6237,N_6597);
nand U10806 (N_10806,N_7839,N_7038);
nor U10807 (N_10807,N_7862,N_7082);
and U10808 (N_10808,N_7623,N_7442);
nand U10809 (N_10809,N_8700,N_8156);
and U10810 (N_10810,N_6762,N_7930);
xnor U10811 (N_10811,N_8189,N_6494);
nor U10812 (N_10812,N_8897,N_8838);
xnor U10813 (N_10813,N_8551,N_7473);
and U10814 (N_10814,N_6226,N_6277);
nand U10815 (N_10815,N_7993,N_8767);
and U10816 (N_10816,N_7759,N_8736);
xor U10817 (N_10817,N_8274,N_7438);
nor U10818 (N_10818,N_8486,N_8423);
nand U10819 (N_10819,N_8612,N_8169);
and U10820 (N_10820,N_6220,N_7305);
nand U10821 (N_10821,N_6127,N_8622);
nand U10822 (N_10822,N_6965,N_8934);
xnor U10823 (N_10823,N_8822,N_6220);
nor U10824 (N_10824,N_7366,N_8744);
or U10825 (N_10825,N_7575,N_7487);
and U10826 (N_10826,N_8417,N_6630);
nor U10827 (N_10827,N_6232,N_7682);
xnor U10828 (N_10828,N_7348,N_6767);
and U10829 (N_10829,N_7645,N_6037);
xnor U10830 (N_10830,N_6304,N_7586);
xor U10831 (N_10831,N_8941,N_8569);
nand U10832 (N_10832,N_6980,N_7031);
and U10833 (N_10833,N_6734,N_8266);
xnor U10834 (N_10834,N_6073,N_7080);
nor U10835 (N_10835,N_7924,N_8223);
nor U10836 (N_10836,N_8506,N_6537);
or U10837 (N_10837,N_7274,N_7361);
nor U10838 (N_10838,N_7762,N_6877);
or U10839 (N_10839,N_6462,N_7471);
and U10840 (N_10840,N_6880,N_6443);
xnor U10841 (N_10841,N_8600,N_7273);
nor U10842 (N_10842,N_8562,N_6760);
xor U10843 (N_10843,N_6636,N_7440);
nand U10844 (N_10844,N_8059,N_6523);
and U10845 (N_10845,N_6857,N_8674);
xnor U10846 (N_10846,N_8072,N_7550);
nor U10847 (N_10847,N_6736,N_6833);
nor U10848 (N_10848,N_7530,N_8781);
or U10849 (N_10849,N_6298,N_8008);
nor U10850 (N_10850,N_6059,N_6642);
xnor U10851 (N_10851,N_7337,N_6212);
nor U10852 (N_10852,N_6539,N_7350);
and U10853 (N_10853,N_6643,N_6623);
nor U10854 (N_10854,N_8374,N_6925);
and U10855 (N_10855,N_7039,N_6648);
xor U10856 (N_10856,N_8063,N_7146);
nand U10857 (N_10857,N_6543,N_7077);
nand U10858 (N_10858,N_6587,N_7329);
xnor U10859 (N_10859,N_8248,N_8586);
xor U10860 (N_10860,N_7786,N_8555);
xor U10861 (N_10861,N_7635,N_7645);
xor U10862 (N_10862,N_8469,N_6230);
xnor U10863 (N_10863,N_8318,N_8496);
or U10864 (N_10864,N_7928,N_7319);
nand U10865 (N_10865,N_8107,N_8316);
and U10866 (N_10866,N_7227,N_6198);
xnor U10867 (N_10867,N_7147,N_8046);
nand U10868 (N_10868,N_7208,N_8487);
nor U10869 (N_10869,N_7741,N_8928);
nor U10870 (N_10870,N_6383,N_7154);
or U10871 (N_10871,N_6842,N_6220);
nor U10872 (N_10872,N_8010,N_7664);
xor U10873 (N_10873,N_8735,N_7504);
nand U10874 (N_10874,N_6085,N_7409);
or U10875 (N_10875,N_7742,N_6324);
xor U10876 (N_10876,N_8219,N_6924);
or U10877 (N_10877,N_7526,N_8241);
nand U10878 (N_10878,N_6406,N_6011);
or U10879 (N_10879,N_8363,N_7908);
or U10880 (N_10880,N_6322,N_7675);
nor U10881 (N_10881,N_8269,N_8008);
or U10882 (N_10882,N_6746,N_8544);
nand U10883 (N_10883,N_6580,N_6025);
nand U10884 (N_10884,N_8398,N_6507);
xnor U10885 (N_10885,N_6086,N_7517);
nor U10886 (N_10886,N_8308,N_7235);
xor U10887 (N_10887,N_6822,N_6107);
nand U10888 (N_10888,N_6482,N_6076);
nand U10889 (N_10889,N_7269,N_8327);
nor U10890 (N_10890,N_8447,N_8850);
nor U10891 (N_10891,N_6737,N_6375);
nor U10892 (N_10892,N_6847,N_6624);
or U10893 (N_10893,N_8758,N_8053);
or U10894 (N_10894,N_7639,N_7486);
nor U10895 (N_10895,N_6246,N_6612);
and U10896 (N_10896,N_7136,N_6865);
nor U10897 (N_10897,N_7476,N_7190);
nand U10898 (N_10898,N_8406,N_8013);
nor U10899 (N_10899,N_8608,N_7421);
nand U10900 (N_10900,N_8373,N_8844);
nand U10901 (N_10901,N_6762,N_6523);
xnor U10902 (N_10902,N_8998,N_8930);
nand U10903 (N_10903,N_8956,N_8567);
xnor U10904 (N_10904,N_8772,N_7850);
nand U10905 (N_10905,N_7924,N_6011);
and U10906 (N_10906,N_8474,N_8436);
xor U10907 (N_10907,N_7580,N_7566);
nor U10908 (N_10908,N_7231,N_6860);
nand U10909 (N_10909,N_8083,N_6163);
or U10910 (N_10910,N_8746,N_6704);
nor U10911 (N_10911,N_7028,N_7325);
nand U10912 (N_10912,N_6859,N_7682);
nor U10913 (N_10913,N_8684,N_7090);
nand U10914 (N_10914,N_6739,N_8808);
xnor U10915 (N_10915,N_8506,N_7575);
xor U10916 (N_10916,N_6785,N_8272);
nand U10917 (N_10917,N_8537,N_8681);
nor U10918 (N_10918,N_7950,N_7884);
nor U10919 (N_10919,N_7212,N_6355);
nand U10920 (N_10920,N_8772,N_7867);
and U10921 (N_10921,N_7543,N_8601);
nand U10922 (N_10922,N_6581,N_8378);
nor U10923 (N_10923,N_6429,N_8873);
and U10924 (N_10924,N_8690,N_6629);
nor U10925 (N_10925,N_8059,N_6990);
and U10926 (N_10926,N_7485,N_8972);
and U10927 (N_10927,N_7858,N_7412);
nand U10928 (N_10928,N_8116,N_8013);
nor U10929 (N_10929,N_6647,N_8550);
xnor U10930 (N_10930,N_6265,N_6074);
nand U10931 (N_10931,N_6152,N_6374);
nand U10932 (N_10932,N_8042,N_8198);
or U10933 (N_10933,N_8616,N_7105);
nor U10934 (N_10934,N_7724,N_7282);
nand U10935 (N_10935,N_7723,N_8608);
nand U10936 (N_10936,N_7987,N_8433);
nand U10937 (N_10937,N_8096,N_7768);
xnor U10938 (N_10938,N_8766,N_7178);
xnor U10939 (N_10939,N_8929,N_8980);
or U10940 (N_10940,N_8782,N_6929);
nand U10941 (N_10941,N_7529,N_7961);
and U10942 (N_10942,N_8819,N_6056);
nand U10943 (N_10943,N_6492,N_7148);
and U10944 (N_10944,N_7579,N_7782);
xor U10945 (N_10945,N_6647,N_6530);
nor U10946 (N_10946,N_7057,N_6257);
or U10947 (N_10947,N_6742,N_7580);
xor U10948 (N_10948,N_8085,N_6080);
xnor U10949 (N_10949,N_6671,N_6866);
nor U10950 (N_10950,N_7698,N_8426);
nor U10951 (N_10951,N_8338,N_8895);
or U10952 (N_10952,N_8635,N_6158);
nor U10953 (N_10953,N_8889,N_7732);
xor U10954 (N_10954,N_7825,N_6799);
nand U10955 (N_10955,N_8293,N_7261);
xor U10956 (N_10956,N_7404,N_8006);
and U10957 (N_10957,N_7178,N_8944);
or U10958 (N_10958,N_8092,N_8382);
nor U10959 (N_10959,N_8969,N_7818);
and U10960 (N_10960,N_6993,N_6222);
or U10961 (N_10961,N_8997,N_8241);
nand U10962 (N_10962,N_8942,N_6766);
nand U10963 (N_10963,N_7728,N_7931);
nor U10964 (N_10964,N_6702,N_8517);
nor U10965 (N_10965,N_8399,N_6833);
and U10966 (N_10966,N_6871,N_8563);
nor U10967 (N_10967,N_7083,N_7410);
nor U10968 (N_10968,N_7669,N_6351);
xnor U10969 (N_10969,N_7416,N_7453);
and U10970 (N_10970,N_8557,N_7811);
nor U10971 (N_10971,N_6648,N_8238);
nand U10972 (N_10972,N_7795,N_8349);
nor U10973 (N_10973,N_7764,N_6418);
xor U10974 (N_10974,N_8251,N_7934);
and U10975 (N_10975,N_6785,N_8200);
or U10976 (N_10976,N_7875,N_6863);
xor U10977 (N_10977,N_7883,N_8006);
or U10978 (N_10978,N_7894,N_6084);
xnor U10979 (N_10979,N_6661,N_8675);
xor U10980 (N_10980,N_8406,N_6397);
xor U10981 (N_10981,N_6897,N_8875);
or U10982 (N_10982,N_7569,N_6137);
and U10983 (N_10983,N_8512,N_6664);
nor U10984 (N_10984,N_6358,N_8044);
nand U10985 (N_10985,N_7243,N_8976);
nor U10986 (N_10986,N_6519,N_6653);
and U10987 (N_10987,N_8770,N_8203);
nand U10988 (N_10988,N_6385,N_6437);
or U10989 (N_10989,N_7756,N_8242);
xnor U10990 (N_10990,N_6740,N_7311);
xnor U10991 (N_10991,N_7611,N_6280);
or U10992 (N_10992,N_7174,N_7551);
nand U10993 (N_10993,N_8506,N_8318);
or U10994 (N_10994,N_7090,N_7792);
nand U10995 (N_10995,N_7838,N_6343);
nor U10996 (N_10996,N_8626,N_8763);
or U10997 (N_10997,N_7058,N_7673);
xnor U10998 (N_10998,N_7428,N_7643);
xnor U10999 (N_10999,N_6183,N_8752);
and U11000 (N_11000,N_8845,N_6865);
or U11001 (N_11001,N_7596,N_8433);
and U11002 (N_11002,N_7162,N_6914);
nor U11003 (N_11003,N_6391,N_6346);
nand U11004 (N_11004,N_7261,N_7099);
xnor U11005 (N_11005,N_6520,N_6781);
or U11006 (N_11006,N_8454,N_8852);
nor U11007 (N_11007,N_8962,N_6957);
nand U11008 (N_11008,N_6713,N_6666);
nor U11009 (N_11009,N_6429,N_8883);
or U11010 (N_11010,N_6752,N_6705);
and U11011 (N_11011,N_8493,N_7469);
nand U11012 (N_11012,N_6752,N_7610);
nor U11013 (N_11013,N_6569,N_7535);
nor U11014 (N_11014,N_6661,N_7158);
or U11015 (N_11015,N_6053,N_6879);
nor U11016 (N_11016,N_6003,N_8112);
xnor U11017 (N_11017,N_6703,N_8230);
and U11018 (N_11018,N_7895,N_6697);
xnor U11019 (N_11019,N_7859,N_6940);
and U11020 (N_11020,N_7035,N_6554);
or U11021 (N_11021,N_7701,N_7775);
or U11022 (N_11022,N_7237,N_7361);
and U11023 (N_11023,N_7993,N_8230);
nor U11024 (N_11024,N_6666,N_7189);
and U11025 (N_11025,N_6360,N_7134);
nand U11026 (N_11026,N_7335,N_8490);
or U11027 (N_11027,N_6372,N_7127);
or U11028 (N_11028,N_8817,N_8313);
or U11029 (N_11029,N_7882,N_8859);
nor U11030 (N_11030,N_7058,N_7844);
xnor U11031 (N_11031,N_6689,N_7403);
xor U11032 (N_11032,N_8299,N_6008);
nand U11033 (N_11033,N_6572,N_8141);
nor U11034 (N_11034,N_8727,N_7386);
or U11035 (N_11035,N_6071,N_8265);
and U11036 (N_11036,N_6172,N_8862);
xor U11037 (N_11037,N_8108,N_6886);
nand U11038 (N_11038,N_6031,N_6677);
and U11039 (N_11039,N_8163,N_6119);
and U11040 (N_11040,N_6374,N_7154);
and U11041 (N_11041,N_7044,N_7998);
nand U11042 (N_11042,N_6571,N_8876);
or U11043 (N_11043,N_6596,N_6299);
or U11044 (N_11044,N_7258,N_7960);
nor U11045 (N_11045,N_6444,N_8985);
or U11046 (N_11046,N_8343,N_7271);
nand U11047 (N_11047,N_6700,N_7593);
nand U11048 (N_11048,N_8110,N_8612);
and U11049 (N_11049,N_8801,N_6819);
xnor U11050 (N_11050,N_8148,N_6391);
and U11051 (N_11051,N_8300,N_6239);
nor U11052 (N_11052,N_8355,N_8411);
and U11053 (N_11053,N_7856,N_8420);
and U11054 (N_11054,N_6644,N_6214);
or U11055 (N_11055,N_7146,N_8164);
nand U11056 (N_11056,N_6685,N_7051);
nand U11057 (N_11057,N_6740,N_6895);
and U11058 (N_11058,N_7092,N_6424);
and U11059 (N_11059,N_6783,N_8146);
xnor U11060 (N_11060,N_7388,N_6531);
or U11061 (N_11061,N_7529,N_7899);
nand U11062 (N_11062,N_7360,N_7898);
xor U11063 (N_11063,N_8998,N_7067);
nand U11064 (N_11064,N_8702,N_7704);
xnor U11065 (N_11065,N_8574,N_8656);
or U11066 (N_11066,N_6478,N_6443);
and U11067 (N_11067,N_8589,N_8446);
or U11068 (N_11068,N_7602,N_7973);
nand U11069 (N_11069,N_7278,N_6612);
nand U11070 (N_11070,N_7528,N_6069);
xor U11071 (N_11071,N_8327,N_6805);
or U11072 (N_11072,N_8339,N_6832);
nor U11073 (N_11073,N_6305,N_8046);
or U11074 (N_11074,N_8239,N_7043);
or U11075 (N_11075,N_8079,N_7521);
nor U11076 (N_11076,N_8482,N_6742);
and U11077 (N_11077,N_7752,N_6576);
xor U11078 (N_11078,N_8189,N_6180);
nor U11079 (N_11079,N_8081,N_6858);
nor U11080 (N_11080,N_8945,N_8728);
nor U11081 (N_11081,N_8891,N_8441);
nand U11082 (N_11082,N_6111,N_7941);
nand U11083 (N_11083,N_8756,N_7136);
nor U11084 (N_11084,N_6184,N_7951);
or U11085 (N_11085,N_7952,N_8771);
xor U11086 (N_11086,N_7234,N_8449);
or U11087 (N_11087,N_6232,N_8244);
and U11088 (N_11088,N_8275,N_6240);
and U11089 (N_11089,N_6744,N_6422);
nor U11090 (N_11090,N_6935,N_7099);
nand U11091 (N_11091,N_6128,N_7305);
and U11092 (N_11092,N_6322,N_7515);
xor U11093 (N_11093,N_6761,N_8444);
nor U11094 (N_11094,N_8851,N_7425);
nand U11095 (N_11095,N_8572,N_8356);
xor U11096 (N_11096,N_6656,N_6948);
nor U11097 (N_11097,N_6892,N_7599);
nand U11098 (N_11098,N_7177,N_6754);
nor U11099 (N_11099,N_8101,N_8471);
nand U11100 (N_11100,N_6289,N_8275);
nor U11101 (N_11101,N_8513,N_6041);
nor U11102 (N_11102,N_6014,N_7719);
and U11103 (N_11103,N_6643,N_7249);
or U11104 (N_11104,N_8604,N_8361);
nand U11105 (N_11105,N_7441,N_6819);
nand U11106 (N_11106,N_6889,N_6447);
xnor U11107 (N_11107,N_6445,N_6457);
nor U11108 (N_11108,N_7674,N_8206);
or U11109 (N_11109,N_7896,N_6373);
nand U11110 (N_11110,N_8420,N_6999);
or U11111 (N_11111,N_6921,N_7701);
xor U11112 (N_11112,N_7896,N_7826);
and U11113 (N_11113,N_8007,N_7470);
or U11114 (N_11114,N_6032,N_6205);
and U11115 (N_11115,N_8414,N_6333);
xor U11116 (N_11116,N_7571,N_6569);
and U11117 (N_11117,N_6583,N_6896);
or U11118 (N_11118,N_6890,N_6650);
nand U11119 (N_11119,N_7125,N_8712);
and U11120 (N_11120,N_6726,N_6632);
xor U11121 (N_11121,N_8189,N_7041);
and U11122 (N_11122,N_8945,N_6370);
and U11123 (N_11123,N_8223,N_6522);
or U11124 (N_11124,N_7481,N_6968);
xor U11125 (N_11125,N_6371,N_6032);
or U11126 (N_11126,N_6226,N_6467);
nor U11127 (N_11127,N_8768,N_6125);
or U11128 (N_11128,N_8435,N_7178);
xor U11129 (N_11129,N_8124,N_8553);
nor U11130 (N_11130,N_6972,N_7483);
nand U11131 (N_11131,N_8529,N_6026);
nor U11132 (N_11132,N_7918,N_7039);
and U11133 (N_11133,N_7234,N_8292);
or U11134 (N_11134,N_7136,N_7187);
xnor U11135 (N_11135,N_6030,N_8367);
or U11136 (N_11136,N_7636,N_8768);
xor U11137 (N_11137,N_7269,N_7696);
and U11138 (N_11138,N_6942,N_7737);
or U11139 (N_11139,N_8376,N_7162);
nand U11140 (N_11140,N_7458,N_8820);
xnor U11141 (N_11141,N_6927,N_6646);
nor U11142 (N_11142,N_8980,N_8033);
or U11143 (N_11143,N_6621,N_8364);
or U11144 (N_11144,N_7955,N_8815);
or U11145 (N_11145,N_6364,N_7129);
or U11146 (N_11146,N_7007,N_8756);
and U11147 (N_11147,N_7924,N_7850);
and U11148 (N_11148,N_8562,N_8922);
nor U11149 (N_11149,N_6903,N_8362);
nor U11150 (N_11150,N_6153,N_6305);
xnor U11151 (N_11151,N_7307,N_6336);
nand U11152 (N_11152,N_6188,N_8010);
or U11153 (N_11153,N_7841,N_8413);
nor U11154 (N_11154,N_8904,N_8576);
nor U11155 (N_11155,N_7787,N_7295);
nand U11156 (N_11156,N_6334,N_6593);
or U11157 (N_11157,N_6906,N_7758);
and U11158 (N_11158,N_8080,N_6952);
or U11159 (N_11159,N_8002,N_8890);
and U11160 (N_11160,N_6503,N_8896);
nor U11161 (N_11161,N_8675,N_8630);
and U11162 (N_11162,N_8276,N_7352);
xnor U11163 (N_11163,N_8750,N_8286);
nor U11164 (N_11164,N_6289,N_7904);
nor U11165 (N_11165,N_8244,N_6230);
and U11166 (N_11166,N_7380,N_8092);
and U11167 (N_11167,N_8630,N_8856);
nand U11168 (N_11168,N_8659,N_8828);
or U11169 (N_11169,N_8927,N_6998);
or U11170 (N_11170,N_8654,N_8298);
nand U11171 (N_11171,N_7250,N_6347);
nand U11172 (N_11172,N_8259,N_6325);
nand U11173 (N_11173,N_8476,N_8902);
nand U11174 (N_11174,N_7611,N_7169);
nand U11175 (N_11175,N_6874,N_6935);
nand U11176 (N_11176,N_8051,N_7749);
or U11177 (N_11177,N_8878,N_6007);
and U11178 (N_11178,N_7803,N_6791);
or U11179 (N_11179,N_8867,N_6659);
nor U11180 (N_11180,N_6504,N_8089);
nand U11181 (N_11181,N_7241,N_8452);
or U11182 (N_11182,N_6229,N_7788);
nor U11183 (N_11183,N_7637,N_7411);
xnor U11184 (N_11184,N_7077,N_8193);
nor U11185 (N_11185,N_6987,N_6204);
and U11186 (N_11186,N_8110,N_8388);
or U11187 (N_11187,N_8603,N_7946);
and U11188 (N_11188,N_6942,N_8387);
and U11189 (N_11189,N_7428,N_8792);
nand U11190 (N_11190,N_8831,N_8910);
nand U11191 (N_11191,N_8293,N_7685);
and U11192 (N_11192,N_8967,N_8093);
xnor U11193 (N_11193,N_8271,N_7021);
xnor U11194 (N_11194,N_6744,N_8385);
or U11195 (N_11195,N_6158,N_7664);
nor U11196 (N_11196,N_7116,N_7407);
or U11197 (N_11197,N_7339,N_8007);
and U11198 (N_11198,N_6987,N_6675);
and U11199 (N_11199,N_8435,N_6653);
and U11200 (N_11200,N_8985,N_7967);
xor U11201 (N_11201,N_7660,N_8496);
or U11202 (N_11202,N_6927,N_8105);
and U11203 (N_11203,N_6143,N_8600);
and U11204 (N_11204,N_7406,N_7833);
and U11205 (N_11205,N_6206,N_8741);
and U11206 (N_11206,N_8282,N_8572);
and U11207 (N_11207,N_8456,N_6506);
or U11208 (N_11208,N_8797,N_7053);
nand U11209 (N_11209,N_6068,N_6184);
and U11210 (N_11210,N_8491,N_7130);
or U11211 (N_11211,N_6690,N_6538);
nand U11212 (N_11212,N_8156,N_8688);
and U11213 (N_11213,N_6858,N_6066);
xnor U11214 (N_11214,N_6741,N_8269);
xor U11215 (N_11215,N_8395,N_7592);
nand U11216 (N_11216,N_7824,N_6101);
nand U11217 (N_11217,N_7111,N_6251);
xor U11218 (N_11218,N_8542,N_6513);
and U11219 (N_11219,N_7846,N_6086);
xor U11220 (N_11220,N_7401,N_8881);
and U11221 (N_11221,N_6738,N_8345);
and U11222 (N_11222,N_7144,N_6270);
xor U11223 (N_11223,N_6535,N_6490);
or U11224 (N_11224,N_7282,N_6276);
xnor U11225 (N_11225,N_6409,N_8045);
nor U11226 (N_11226,N_8205,N_8735);
nand U11227 (N_11227,N_6142,N_8362);
nor U11228 (N_11228,N_7499,N_7970);
nor U11229 (N_11229,N_8080,N_8206);
and U11230 (N_11230,N_7784,N_7746);
xnor U11231 (N_11231,N_8959,N_6517);
nand U11232 (N_11232,N_7960,N_7565);
and U11233 (N_11233,N_8429,N_7349);
or U11234 (N_11234,N_6060,N_8895);
or U11235 (N_11235,N_6401,N_6247);
nand U11236 (N_11236,N_6703,N_7386);
xor U11237 (N_11237,N_6633,N_7259);
nor U11238 (N_11238,N_7990,N_6133);
and U11239 (N_11239,N_7179,N_6432);
xor U11240 (N_11240,N_7626,N_7021);
and U11241 (N_11241,N_6045,N_8457);
nor U11242 (N_11242,N_7083,N_7753);
nor U11243 (N_11243,N_7696,N_8492);
xnor U11244 (N_11244,N_8307,N_6456);
xor U11245 (N_11245,N_7533,N_8844);
or U11246 (N_11246,N_8696,N_8711);
and U11247 (N_11247,N_7283,N_7001);
and U11248 (N_11248,N_7040,N_8304);
nand U11249 (N_11249,N_6500,N_7123);
nor U11250 (N_11250,N_7087,N_7021);
or U11251 (N_11251,N_6934,N_7223);
nand U11252 (N_11252,N_6552,N_7708);
nor U11253 (N_11253,N_7543,N_7600);
xor U11254 (N_11254,N_8303,N_8532);
or U11255 (N_11255,N_7078,N_8898);
nand U11256 (N_11256,N_7908,N_8774);
nand U11257 (N_11257,N_7459,N_8067);
xnor U11258 (N_11258,N_7605,N_6113);
xnor U11259 (N_11259,N_8478,N_8097);
nand U11260 (N_11260,N_8226,N_7090);
or U11261 (N_11261,N_7797,N_7182);
xor U11262 (N_11262,N_7607,N_7925);
nor U11263 (N_11263,N_7081,N_8784);
or U11264 (N_11264,N_6374,N_6817);
xor U11265 (N_11265,N_7930,N_8178);
nand U11266 (N_11266,N_7484,N_8795);
and U11267 (N_11267,N_6770,N_7186);
nand U11268 (N_11268,N_7836,N_7607);
and U11269 (N_11269,N_8062,N_7958);
or U11270 (N_11270,N_7954,N_8212);
xnor U11271 (N_11271,N_6325,N_8347);
xor U11272 (N_11272,N_7762,N_8240);
or U11273 (N_11273,N_8386,N_6205);
nor U11274 (N_11274,N_7622,N_6021);
xor U11275 (N_11275,N_7318,N_7956);
xor U11276 (N_11276,N_8476,N_6749);
nor U11277 (N_11277,N_7986,N_8607);
xnor U11278 (N_11278,N_6951,N_8119);
and U11279 (N_11279,N_7828,N_7978);
xnor U11280 (N_11280,N_6275,N_7654);
nor U11281 (N_11281,N_6732,N_8008);
xor U11282 (N_11282,N_8202,N_7736);
and U11283 (N_11283,N_7604,N_7433);
nand U11284 (N_11284,N_6418,N_8838);
nor U11285 (N_11285,N_7562,N_8832);
xnor U11286 (N_11286,N_7652,N_8019);
nor U11287 (N_11287,N_8728,N_8619);
and U11288 (N_11288,N_8348,N_8989);
nor U11289 (N_11289,N_8638,N_7113);
nor U11290 (N_11290,N_7262,N_8912);
xnor U11291 (N_11291,N_8973,N_8126);
or U11292 (N_11292,N_7201,N_7345);
or U11293 (N_11293,N_7911,N_8881);
and U11294 (N_11294,N_6564,N_7563);
nor U11295 (N_11295,N_6533,N_6744);
and U11296 (N_11296,N_7745,N_8295);
and U11297 (N_11297,N_6955,N_6682);
xnor U11298 (N_11298,N_8549,N_8195);
or U11299 (N_11299,N_6955,N_8054);
xor U11300 (N_11300,N_6627,N_6708);
nor U11301 (N_11301,N_7627,N_6595);
or U11302 (N_11302,N_7386,N_6119);
nand U11303 (N_11303,N_6534,N_7335);
or U11304 (N_11304,N_7901,N_7722);
nand U11305 (N_11305,N_6960,N_6006);
xor U11306 (N_11306,N_8006,N_8241);
or U11307 (N_11307,N_7717,N_8880);
xor U11308 (N_11308,N_8896,N_7482);
xor U11309 (N_11309,N_8330,N_8677);
or U11310 (N_11310,N_8632,N_7294);
or U11311 (N_11311,N_8137,N_7705);
and U11312 (N_11312,N_7959,N_7282);
and U11313 (N_11313,N_8451,N_7875);
nand U11314 (N_11314,N_6965,N_6931);
xor U11315 (N_11315,N_8588,N_8623);
nand U11316 (N_11316,N_7400,N_6637);
nand U11317 (N_11317,N_6860,N_7730);
nor U11318 (N_11318,N_6579,N_7671);
nand U11319 (N_11319,N_8158,N_8872);
or U11320 (N_11320,N_8143,N_8771);
nand U11321 (N_11321,N_6208,N_7447);
or U11322 (N_11322,N_7687,N_7366);
nand U11323 (N_11323,N_7086,N_8994);
and U11324 (N_11324,N_6040,N_7968);
nand U11325 (N_11325,N_7570,N_6562);
xnor U11326 (N_11326,N_6206,N_6777);
nand U11327 (N_11327,N_6788,N_8733);
xnor U11328 (N_11328,N_8272,N_7204);
nor U11329 (N_11329,N_7947,N_7055);
xor U11330 (N_11330,N_8993,N_8153);
xor U11331 (N_11331,N_7065,N_8873);
or U11332 (N_11332,N_6628,N_7762);
or U11333 (N_11333,N_7096,N_7681);
xnor U11334 (N_11334,N_6716,N_7042);
nor U11335 (N_11335,N_8531,N_7932);
nand U11336 (N_11336,N_8751,N_6401);
and U11337 (N_11337,N_8419,N_6928);
or U11338 (N_11338,N_8058,N_7410);
or U11339 (N_11339,N_8447,N_8955);
xnor U11340 (N_11340,N_7367,N_7071);
xnor U11341 (N_11341,N_6182,N_7982);
xor U11342 (N_11342,N_7044,N_7076);
or U11343 (N_11343,N_6264,N_8063);
xor U11344 (N_11344,N_6330,N_6475);
nor U11345 (N_11345,N_7714,N_6511);
xor U11346 (N_11346,N_7410,N_7830);
xnor U11347 (N_11347,N_7163,N_6434);
xnor U11348 (N_11348,N_8836,N_6305);
and U11349 (N_11349,N_8501,N_7058);
xnor U11350 (N_11350,N_6968,N_7264);
xnor U11351 (N_11351,N_6820,N_7594);
or U11352 (N_11352,N_7145,N_6996);
xor U11353 (N_11353,N_7155,N_8098);
or U11354 (N_11354,N_6382,N_8336);
nand U11355 (N_11355,N_6663,N_7500);
nor U11356 (N_11356,N_6423,N_6034);
nor U11357 (N_11357,N_8019,N_7111);
nand U11358 (N_11358,N_7439,N_8734);
nor U11359 (N_11359,N_6440,N_6849);
and U11360 (N_11360,N_6810,N_7976);
nand U11361 (N_11361,N_7652,N_7111);
and U11362 (N_11362,N_6908,N_8811);
xnor U11363 (N_11363,N_7874,N_8452);
and U11364 (N_11364,N_8407,N_6210);
xor U11365 (N_11365,N_7072,N_6157);
or U11366 (N_11366,N_6317,N_8734);
nor U11367 (N_11367,N_6334,N_7211);
nor U11368 (N_11368,N_7228,N_7708);
and U11369 (N_11369,N_6151,N_6448);
and U11370 (N_11370,N_6642,N_6793);
nor U11371 (N_11371,N_6649,N_6296);
or U11372 (N_11372,N_8686,N_8934);
xor U11373 (N_11373,N_6111,N_6041);
xor U11374 (N_11374,N_8655,N_6115);
xnor U11375 (N_11375,N_8642,N_6720);
xor U11376 (N_11376,N_8688,N_8066);
nor U11377 (N_11377,N_6076,N_7115);
nor U11378 (N_11378,N_6986,N_8640);
and U11379 (N_11379,N_7562,N_8252);
and U11380 (N_11380,N_8835,N_7375);
nor U11381 (N_11381,N_8762,N_7959);
nand U11382 (N_11382,N_8513,N_8167);
or U11383 (N_11383,N_6985,N_8226);
xnor U11384 (N_11384,N_7306,N_6229);
and U11385 (N_11385,N_8958,N_7285);
and U11386 (N_11386,N_8365,N_6133);
xnor U11387 (N_11387,N_6859,N_8154);
nand U11388 (N_11388,N_8951,N_7577);
nor U11389 (N_11389,N_6916,N_6804);
or U11390 (N_11390,N_7933,N_6033);
xor U11391 (N_11391,N_6005,N_7860);
nand U11392 (N_11392,N_6455,N_8124);
nor U11393 (N_11393,N_8212,N_6055);
or U11394 (N_11394,N_8259,N_7550);
nor U11395 (N_11395,N_6195,N_7634);
nand U11396 (N_11396,N_8116,N_7978);
xor U11397 (N_11397,N_8419,N_6169);
xor U11398 (N_11398,N_7518,N_7471);
nand U11399 (N_11399,N_7367,N_8474);
and U11400 (N_11400,N_6515,N_8969);
or U11401 (N_11401,N_6126,N_6501);
xor U11402 (N_11402,N_7815,N_8132);
xnor U11403 (N_11403,N_8480,N_6029);
and U11404 (N_11404,N_6710,N_6791);
and U11405 (N_11405,N_8117,N_6350);
xnor U11406 (N_11406,N_6871,N_8179);
xnor U11407 (N_11407,N_7759,N_6283);
xor U11408 (N_11408,N_8634,N_7338);
nor U11409 (N_11409,N_7546,N_6231);
nand U11410 (N_11410,N_8879,N_8447);
xnor U11411 (N_11411,N_7520,N_6566);
nor U11412 (N_11412,N_7548,N_6436);
or U11413 (N_11413,N_8860,N_8836);
or U11414 (N_11414,N_6316,N_6311);
nor U11415 (N_11415,N_6680,N_6937);
and U11416 (N_11416,N_6234,N_6075);
or U11417 (N_11417,N_6758,N_7729);
nor U11418 (N_11418,N_8426,N_8890);
nor U11419 (N_11419,N_7232,N_6263);
and U11420 (N_11420,N_8214,N_6492);
nor U11421 (N_11421,N_8994,N_7525);
xnor U11422 (N_11422,N_6198,N_8156);
and U11423 (N_11423,N_8683,N_8169);
xnor U11424 (N_11424,N_7391,N_8249);
nand U11425 (N_11425,N_7192,N_6896);
nor U11426 (N_11426,N_7674,N_8011);
or U11427 (N_11427,N_6940,N_8853);
or U11428 (N_11428,N_8421,N_6417);
and U11429 (N_11429,N_8525,N_6486);
nor U11430 (N_11430,N_6226,N_7891);
xnor U11431 (N_11431,N_8944,N_7896);
nand U11432 (N_11432,N_7020,N_7883);
nand U11433 (N_11433,N_7067,N_6502);
nor U11434 (N_11434,N_6061,N_6128);
or U11435 (N_11435,N_6491,N_6659);
or U11436 (N_11436,N_6351,N_8662);
nor U11437 (N_11437,N_6180,N_8078);
or U11438 (N_11438,N_6072,N_6306);
and U11439 (N_11439,N_8106,N_6822);
or U11440 (N_11440,N_8199,N_6112);
and U11441 (N_11441,N_8946,N_6580);
nand U11442 (N_11442,N_7203,N_6565);
nor U11443 (N_11443,N_6216,N_8270);
and U11444 (N_11444,N_6372,N_6838);
nor U11445 (N_11445,N_7817,N_6827);
nand U11446 (N_11446,N_7979,N_8741);
and U11447 (N_11447,N_8145,N_6354);
and U11448 (N_11448,N_6289,N_6300);
and U11449 (N_11449,N_7311,N_6666);
nand U11450 (N_11450,N_7953,N_7330);
nor U11451 (N_11451,N_7440,N_6631);
and U11452 (N_11452,N_8794,N_8821);
or U11453 (N_11453,N_8403,N_7408);
xnor U11454 (N_11454,N_6940,N_6759);
or U11455 (N_11455,N_7244,N_6811);
and U11456 (N_11456,N_8802,N_8081);
xor U11457 (N_11457,N_7246,N_8843);
xnor U11458 (N_11458,N_8308,N_7404);
nor U11459 (N_11459,N_8388,N_8207);
xnor U11460 (N_11460,N_8266,N_6402);
xor U11461 (N_11461,N_8761,N_8840);
and U11462 (N_11462,N_6298,N_7115);
nor U11463 (N_11463,N_6354,N_8030);
nor U11464 (N_11464,N_6767,N_7993);
nand U11465 (N_11465,N_8803,N_7205);
and U11466 (N_11466,N_7079,N_8723);
xor U11467 (N_11467,N_7227,N_6794);
xor U11468 (N_11468,N_7918,N_8852);
and U11469 (N_11469,N_6777,N_8590);
xnor U11470 (N_11470,N_6005,N_7242);
xor U11471 (N_11471,N_6218,N_8098);
nand U11472 (N_11472,N_7587,N_8249);
xnor U11473 (N_11473,N_6967,N_7175);
nor U11474 (N_11474,N_7662,N_6202);
nand U11475 (N_11475,N_8256,N_8816);
nor U11476 (N_11476,N_6176,N_7652);
and U11477 (N_11477,N_6016,N_6219);
and U11478 (N_11478,N_8253,N_6125);
nand U11479 (N_11479,N_7459,N_7492);
xor U11480 (N_11480,N_7730,N_7029);
or U11481 (N_11481,N_6842,N_6161);
nor U11482 (N_11482,N_6879,N_8003);
xor U11483 (N_11483,N_7047,N_8988);
nor U11484 (N_11484,N_8335,N_6616);
and U11485 (N_11485,N_6676,N_7851);
nand U11486 (N_11486,N_6760,N_7499);
nand U11487 (N_11487,N_8644,N_6420);
and U11488 (N_11488,N_8632,N_7931);
nor U11489 (N_11489,N_6235,N_7897);
and U11490 (N_11490,N_7496,N_8960);
or U11491 (N_11491,N_7821,N_8056);
or U11492 (N_11492,N_7579,N_8945);
and U11493 (N_11493,N_7657,N_7477);
and U11494 (N_11494,N_8944,N_6887);
nand U11495 (N_11495,N_8774,N_7539);
and U11496 (N_11496,N_6409,N_8165);
xnor U11497 (N_11497,N_8046,N_6606);
nor U11498 (N_11498,N_7091,N_6215);
nor U11499 (N_11499,N_7547,N_6237);
nor U11500 (N_11500,N_8493,N_6573);
xor U11501 (N_11501,N_6414,N_7612);
and U11502 (N_11502,N_6490,N_7309);
and U11503 (N_11503,N_8223,N_8508);
nand U11504 (N_11504,N_7481,N_6675);
and U11505 (N_11505,N_6171,N_8188);
nor U11506 (N_11506,N_6786,N_7372);
nor U11507 (N_11507,N_7797,N_7717);
nand U11508 (N_11508,N_7153,N_8540);
xnor U11509 (N_11509,N_6552,N_6050);
nor U11510 (N_11510,N_6828,N_6342);
or U11511 (N_11511,N_7131,N_6730);
xor U11512 (N_11512,N_8709,N_6544);
and U11513 (N_11513,N_6310,N_8428);
or U11514 (N_11514,N_7730,N_7602);
and U11515 (N_11515,N_7188,N_8144);
xnor U11516 (N_11516,N_7887,N_6363);
or U11517 (N_11517,N_8853,N_7974);
xnor U11518 (N_11518,N_8034,N_7220);
and U11519 (N_11519,N_6469,N_7325);
and U11520 (N_11520,N_7802,N_7791);
and U11521 (N_11521,N_7500,N_8174);
and U11522 (N_11522,N_6037,N_8279);
and U11523 (N_11523,N_8836,N_8541);
nor U11524 (N_11524,N_8740,N_8712);
nor U11525 (N_11525,N_7578,N_8701);
xnor U11526 (N_11526,N_6434,N_7664);
nor U11527 (N_11527,N_6341,N_6540);
nand U11528 (N_11528,N_8125,N_7906);
xor U11529 (N_11529,N_8665,N_8861);
or U11530 (N_11530,N_8153,N_8141);
xnor U11531 (N_11531,N_6317,N_6135);
nor U11532 (N_11532,N_7598,N_6027);
or U11533 (N_11533,N_8362,N_7939);
xnor U11534 (N_11534,N_8892,N_6819);
xor U11535 (N_11535,N_7598,N_8207);
xnor U11536 (N_11536,N_8453,N_6875);
xor U11537 (N_11537,N_7852,N_8346);
nand U11538 (N_11538,N_8941,N_6627);
nand U11539 (N_11539,N_8815,N_8063);
xor U11540 (N_11540,N_7810,N_6778);
and U11541 (N_11541,N_6836,N_8289);
nand U11542 (N_11542,N_6718,N_7115);
nand U11543 (N_11543,N_6622,N_7393);
and U11544 (N_11544,N_6460,N_6361);
xnor U11545 (N_11545,N_7008,N_8272);
and U11546 (N_11546,N_8389,N_7447);
or U11547 (N_11547,N_6243,N_8038);
nor U11548 (N_11548,N_8742,N_8758);
nor U11549 (N_11549,N_7462,N_7018);
and U11550 (N_11550,N_7814,N_8260);
and U11551 (N_11551,N_6284,N_8880);
or U11552 (N_11552,N_8803,N_7499);
or U11553 (N_11553,N_6004,N_8996);
nor U11554 (N_11554,N_6590,N_6498);
xor U11555 (N_11555,N_7705,N_8739);
nor U11556 (N_11556,N_6536,N_8068);
nand U11557 (N_11557,N_6211,N_6357);
or U11558 (N_11558,N_6331,N_8808);
xnor U11559 (N_11559,N_6583,N_8636);
nor U11560 (N_11560,N_6694,N_7962);
nor U11561 (N_11561,N_6846,N_6573);
nor U11562 (N_11562,N_6349,N_8101);
nand U11563 (N_11563,N_7566,N_6885);
nor U11564 (N_11564,N_6173,N_8752);
nor U11565 (N_11565,N_6192,N_7903);
and U11566 (N_11566,N_7524,N_6866);
nand U11567 (N_11567,N_6972,N_8116);
nand U11568 (N_11568,N_8779,N_8915);
nand U11569 (N_11569,N_8682,N_8280);
nand U11570 (N_11570,N_8195,N_6869);
nand U11571 (N_11571,N_7110,N_8062);
nor U11572 (N_11572,N_7314,N_8746);
or U11573 (N_11573,N_7708,N_8355);
nand U11574 (N_11574,N_6724,N_7681);
xor U11575 (N_11575,N_8391,N_7402);
and U11576 (N_11576,N_6834,N_8852);
nor U11577 (N_11577,N_6468,N_8769);
or U11578 (N_11578,N_6880,N_8582);
or U11579 (N_11579,N_6123,N_7579);
xnor U11580 (N_11580,N_8340,N_7517);
and U11581 (N_11581,N_7728,N_7773);
nand U11582 (N_11582,N_8412,N_8491);
nor U11583 (N_11583,N_8396,N_6353);
or U11584 (N_11584,N_8237,N_6078);
nand U11585 (N_11585,N_6278,N_7111);
nand U11586 (N_11586,N_7844,N_8137);
nand U11587 (N_11587,N_6985,N_8427);
nor U11588 (N_11588,N_6805,N_8423);
xor U11589 (N_11589,N_6535,N_8102);
xor U11590 (N_11590,N_6511,N_6533);
and U11591 (N_11591,N_7268,N_8980);
xor U11592 (N_11592,N_7709,N_8103);
xnor U11593 (N_11593,N_7159,N_8245);
nand U11594 (N_11594,N_6743,N_8731);
and U11595 (N_11595,N_8600,N_6061);
nor U11596 (N_11596,N_7960,N_6975);
or U11597 (N_11597,N_6678,N_8178);
and U11598 (N_11598,N_7164,N_6423);
or U11599 (N_11599,N_8907,N_8879);
or U11600 (N_11600,N_8214,N_8094);
nor U11601 (N_11601,N_6826,N_8438);
xor U11602 (N_11602,N_6855,N_8619);
nor U11603 (N_11603,N_6380,N_7894);
nor U11604 (N_11604,N_7087,N_7124);
nor U11605 (N_11605,N_8431,N_8329);
nand U11606 (N_11606,N_7083,N_8376);
and U11607 (N_11607,N_7958,N_6943);
or U11608 (N_11608,N_6730,N_7089);
nor U11609 (N_11609,N_7389,N_6136);
or U11610 (N_11610,N_8416,N_8110);
and U11611 (N_11611,N_7822,N_7537);
nand U11612 (N_11612,N_6094,N_7897);
nand U11613 (N_11613,N_6599,N_8116);
nor U11614 (N_11614,N_7099,N_6640);
or U11615 (N_11615,N_8701,N_6066);
and U11616 (N_11616,N_6019,N_7195);
and U11617 (N_11617,N_6102,N_7284);
or U11618 (N_11618,N_7422,N_7054);
and U11619 (N_11619,N_7497,N_7609);
and U11620 (N_11620,N_8941,N_8902);
and U11621 (N_11621,N_6034,N_8277);
nor U11622 (N_11622,N_6260,N_6146);
nor U11623 (N_11623,N_6339,N_6907);
xor U11624 (N_11624,N_6259,N_8559);
or U11625 (N_11625,N_8450,N_8724);
or U11626 (N_11626,N_7820,N_7120);
nor U11627 (N_11627,N_7344,N_7137);
nor U11628 (N_11628,N_6218,N_7576);
xnor U11629 (N_11629,N_6940,N_8136);
xnor U11630 (N_11630,N_6187,N_6629);
and U11631 (N_11631,N_8337,N_8969);
nand U11632 (N_11632,N_6830,N_8080);
nor U11633 (N_11633,N_6617,N_8366);
and U11634 (N_11634,N_7493,N_7339);
nor U11635 (N_11635,N_8563,N_8815);
nor U11636 (N_11636,N_6181,N_6735);
or U11637 (N_11637,N_8184,N_7426);
xnor U11638 (N_11638,N_6287,N_7375);
and U11639 (N_11639,N_6282,N_7634);
or U11640 (N_11640,N_7213,N_7095);
or U11641 (N_11641,N_8401,N_8418);
nand U11642 (N_11642,N_8035,N_6519);
nor U11643 (N_11643,N_6233,N_6983);
xor U11644 (N_11644,N_6184,N_8096);
and U11645 (N_11645,N_6305,N_6075);
or U11646 (N_11646,N_7577,N_8532);
and U11647 (N_11647,N_7003,N_7768);
xnor U11648 (N_11648,N_8469,N_7132);
nor U11649 (N_11649,N_8465,N_7625);
and U11650 (N_11650,N_8042,N_6467);
and U11651 (N_11651,N_8751,N_8773);
nor U11652 (N_11652,N_7777,N_8200);
and U11653 (N_11653,N_8933,N_7044);
nor U11654 (N_11654,N_7170,N_6885);
nand U11655 (N_11655,N_8137,N_6181);
xor U11656 (N_11656,N_7528,N_6203);
or U11657 (N_11657,N_7028,N_6155);
or U11658 (N_11658,N_8747,N_8318);
nor U11659 (N_11659,N_6807,N_8514);
and U11660 (N_11660,N_7341,N_6843);
xnor U11661 (N_11661,N_8292,N_7947);
xor U11662 (N_11662,N_7758,N_8134);
or U11663 (N_11663,N_8112,N_6191);
or U11664 (N_11664,N_6810,N_8689);
or U11665 (N_11665,N_6274,N_7384);
and U11666 (N_11666,N_7916,N_6513);
nor U11667 (N_11667,N_8968,N_8633);
xnor U11668 (N_11668,N_6716,N_6093);
xor U11669 (N_11669,N_8625,N_8916);
nor U11670 (N_11670,N_8557,N_8379);
nand U11671 (N_11671,N_7379,N_8087);
nand U11672 (N_11672,N_7257,N_7953);
xor U11673 (N_11673,N_8650,N_6443);
or U11674 (N_11674,N_8045,N_7203);
xor U11675 (N_11675,N_7043,N_7615);
and U11676 (N_11676,N_7998,N_8102);
nor U11677 (N_11677,N_7928,N_8618);
nor U11678 (N_11678,N_7407,N_6101);
or U11679 (N_11679,N_6340,N_8786);
nand U11680 (N_11680,N_8810,N_8703);
xor U11681 (N_11681,N_8362,N_7576);
or U11682 (N_11682,N_7883,N_6654);
and U11683 (N_11683,N_7689,N_6184);
xnor U11684 (N_11684,N_8170,N_7675);
nand U11685 (N_11685,N_8542,N_6455);
and U11686 (N_11686,N_8665,N_8048);
or U11687 (N_11687,N_7441,N_8130);
xor U11688 (N_11688,N_6083,N_7901);
or U11689 (N_11689,N_7260,N_6559);
xnor U11690 (N_11690,N_6831,N_6430);
xor U11691 (N_11691,N_7518,N_6567);
or U11692 (N_11692,N_8552,N_6097);
xnor U11693 (N_11693,N_8389,N_7688);
and U11694 (N_11694,N_7191,N_7976);
or U11695 (N_11695,N_8315,N_6349);
nor U11696 (N_11696,N_7832,N_8970);
nor U11697 (N_11697,N_8128,N_7160);
nand U11698 (N_11698,N_7924,N_6696);
and U11699 (N_11699,N_6906,N_6832);
nand U11700 (N_11700,N_6480,N_7505);
and U11701 (N_11701,N_7431,N_8668);
and U11702 (N_11702,N_8045,N_7858);
or U11703 (N_11703,N_8341,N_8780);
xnor U11704 (N_11704,N_8292,N_6075);
and U11705 (N_11705,N_6127,N_8805);
or U11706 (N_11706,N_7817,N_8575);
nor U11707 (N_11707,N_7763,N_8701);
xor U11708 (N_11708,N_6606,N_7703);
nor U11709 (N_11709,N_8844,N_6659);
and U11710 (N_11710,N_7412,N_6799);
or U11711 (N_11711,N_6537,N_8080);
nand U11712 (N_11712,N_8096,N_7257);
or U11713 (N_11713,N_8025,N_7196);
nand U11714 (N_11714,N_8380,N_7990);
or U11715 (N_11715,N_8373,N_7053);
xor U11716 (N_11716,N_7283,N_8232);
nor U11717 (N_11717,N_8714,N_6704);
and U11718 (N_11718,N_6270,N_6559);
nand U11719 (N_11719,N_7721,N_6356);
and U11720 (N_11720,N_8438,N_8875);
nor U11721 (N_11721,N_6887,N_7051);
or U11722 (N_11722,N_8666,N_6666);
xnor U11723 (N_11723,N_7871,N_6704);
xnor U11724 (N_11724,N_6373,N_7833);
and U11725 (N_11725,N_7385,N_8868);
nor U11726 (N_11726,N_7198,N_8349);
xnor U11727 (N_11727,N_7814,N_8945);
or U11728 (N_11728,N_6788,N_7147);
xnor U11729 (N_11729,N_7191,N_7433);
xnor U11730 (N_11730,N_8773,N_8196);
nor U11731 (N_11731,N_8602,N_8447);
xnor U11732 (N_11732,N_8924,N_8416);
nand U11733 (N_11733,N_7534,N_8929);
and U11734 (N_11734,N_7369,N_6538);
nor U11735 (N_11735,N_6941,N_8697);
nor U11736 (N_11736,N_7199,N_8412);
or U11737 (N_11737,N_7976,N_6257);
xnor U11738 (N_11738,N_7932,N_6100);
nor U11739 (N_11739,N_6881,N_7889);
nand U11740 (N_11740,N_8884,N_8532);
and U11741 (N_11741,N_8250,N_8721);
nor U11742 (N_11742,N_6374,N_7492);
and U11743 (N_11743,N_8295,N_6948);
nand U11744 (N_11744,N_6227,N_6648);
nand U11745 (N_11745,N_8403,N_6866);
nand U11746 (N_11746,N_6916,N_7774);
and U11747 (N_11747,N_6377,N_6840);
xor U11748 (N_11748,N_7761,N_7960);
nor U11749 (N_11749,N_8126,N_8711);
or U11750 (N_11750,N_6751,N_8658);
nand U11751 (N_11751,N_8951,N_8215);
and U11752 (N_11752,N_8588,N_7825);
and U11753 (N_11753,N_8055,N_8513);
or U11754 (N_11754,N_7120,N_8302);
and U11755 (N_11755,N_7921,N_6437);
xor U11756 (N_11756,N_6131,N_7835);
xor U11757 (N_11757,N_7514,N_8369);
and U11758 (N_11758,N_7848,N_7272);
or U11759 (N_11759,N_7639,N_8937);
or U11760 (N_11760,N_7389,N_7175);
or U11761 (N_11761,N_6632,N_7851);
xor U11762 (N_11762,N_7969,N_7104);
and U11763 (N_11763,N_8195,N_8418);
nand U11764 (N_11764,N_8667,N_8673);
xnor U11765 (N_11765,N_6284,N_7803);
nand U11766 (N_11766,N_8805,N_6472);
nand U11767 (N_11767,N_7418,N_8704);
and U11768 (N_11768,N_8812,N_8607);
or U11769 (N_11769,N_8973,N_8250);
nand U11770 (N_11770,N_7248,N_7896);
nand U11771 (N_11771,N_7445,N_7452);
nor U11772 (N_11772,N_7315,N_6379);
and U11773 (N_11773,N_7968,N_7713);
nor U11774 (N_11774,N_8656,N_8645);
xor U11775 (N_11775,N_6649,N_8416);
nor U11776 (N_11776,N_6300,N_6508);
nor U11777 (N_11777,N_8111,N_7413);
nand U11778 (N_11778,N_8644,N_6314);
nand U11779 (N_11779,N_6952,N_7019);
xnor U11780 (N_11780,N_6236,N_8140);
or U11781 (N_11781,N_6969,N_7216);
and U11782 (N_11782,N_8089,N_8478);
xnor U11783 (N_11783,N_8014,N_6757);
nor U11784 (N_11784,N_6131,N_6731);
or U11785 (N_11785,N_7494,N_8684);
or U11786 (N_11786,N_7886,N_8888);
and U11787 (N_11787,N_8978,N_6084);
nand U11788 (N_11788,N_8615,N_7095);
nor U11789 (N_11789,N_6673,N_8281);
xnor U11790 (N_11790,N_6356,N_8934);
nor U11791 (N_11791,N_6135,N_7703);
and U11792 (N_11792,N_6913,N_7377);
nor U11793 (N_11793,N_6666,N_7651);
or U11794 (N_11794,N_6590,N_6684);
nand U11795 (N_11795,N_6319,N_6059);
or U11796 (N_11796,N_7093,N_6596);
and U11797 (N_11797,N_6010,N_7504);
nand U11798 (N_11798,N_6589,N_8336);
nand U11799 (N_11799,N_8613,N_6430);
nand U11800 (N_11800,N_8174,N_8102);
xor U11801 (N_11801,N_7911,N_7142);
nand U11802 (N_11802,N_6487,N_8075);
or U11803 (N_11803,N_7443,N_8648);
nand U11804 (N_11804,N_7195,N_7270);
or U11805 (N_11805,N_6252,N_8916);
or U11806 (N_11806,N_7392,N_7893);
or U11807 (N_11807,N_6239,N_7995);
xnor U11808 (N_11808,N_8856,N_7001);
xnor U11809 (N_11809,N_6101,N_7668);
or U11810 (N_11810,N_7960,N_8590);
xnor U11811 (N_11811,N_8256,N_6302);
nor U11812 (N_11812,N_7117,N_8376);
nor U11813 (N_11813,N_7498,N_6526);
and U11814 (N_11814,N_7403,N_7673);
and U11815 (N_11815,N_7992,N_6679);
nor U11816 (N_11816,N_7243,N_6651);
xnor U11817 (N_11817,N_8206,N_8928);
nand U11818 (N_11818,N_8976,N_8048);
nor U11819 (N_11819,N_6816,N_6349);
nand U11820 (N_11820,N_8320,N_8068);
or U11821 (N_11821,N_6004,N_7293);
and U11822 (N_11822,N_7881,N_8547);
and U11823 (N_11823,N_6501,N_6651);
nor U11824 (N_11824,N_8889,N_7187);
nand U11825 (N_11825,N_7050,N_6547);
nand U11826 (N_11826,N_8735,N_8667);
nor U11827 (N_11827,N_6641,N_6413);
nor U11828 (N_11828,N_6199,N_7061);
nor U11829 (N_11829,N_7653,N_7763);
xor U11830 (N_11830,N_8340,N_7444);
nand U11831 (N_11831,N_8908,N_6664);
xor U11832 (N_11832,N_6825,N_7247);
nand U11833 (N_11833,N_7079,N_6316);
or U11834 (N_11834,N_7754,N_7999);
xnor U11835 (N_11835,N_6635,N_6490);
and U11836 (N_11836,N_6708,N_7640);
xor U11837 (N_11837,N_6713,N_8963);
nor U11838 (N_11838,N_7959,N_7766);
nor U11839 (N_11839,N_7321,N_6466);
and U11840 (N_11840,N_7710,N_8994);
nand U11841 (N_11841,N_6930,N_7286);
nand U11842 (N_11842,N_6580,N_8692);
xor U11843 (N_11843,N_7460,N_8347);
nand U11844 (N_11844,N_8307,N_6512);
xor U11845 (N_11845,N_7742,N_8790);
nor U11846 (N_11846,N_7471,N_8754);
nor U11847 (N_11847,N_8013,N_8727);
nor U11848 (N_11848,N_6925,N_8620);
and U11849 (N_11849,N_8226,N_8371);
and U11850 (N_11850,N_8227,N_6537);
nor U11851 (N_11851,N_6417,N_6657);
nor U11852 (N_11852,N_8128,N_7489);
xnor U11853 (N_11853,N_6112,N_7682);
nand U11854 (N_11854,N_7643,N_6597);
xor U11855 (N_11855,N_7598,N_6363);
or U11856 (N_11856,N_6815,N_8977);
or U11857 (N_11857,N_7297,N_8505);
nand U11858 (N_11858,N_7904,N_8307);
nand U11859 (N_11859,N_6920,N_8829);
xnor U11860 (N_11860,N_6367,N_7547);
and U11861 (N_11861,N_8983,N_7111);
nand U11862 (N_11862,N_6516,N_6245);
xnor U11863 (N_11863,N_6706,N_7679);
nand U11864 (N_11864,N_7815,N_6242);
xnor U11865 (N_11865,N_8759,N_7207);
and U11866 (N_11866,N_6058,N_6321);
or U11867 (N_11867,N_8394,N_7174);
xor U11868 (N_11868,N_8242,N_6413);
nor U11869 (N_11869,N_8703,N_7208);
and U11870 (N_11870,N_6742,N_7431);
and U11871 (N_11871,N_6868,N_8908);
or U11872 (N_11872,N_6642,N_6566);
and U11873 (N_11873,N_8770,N_6130);
xnor U11874 (N_11874,N_6998,N_6258);
nand U11875 (N_11875,N_6381,N_6831);
nor U11876 (N_11876,N_6205,N_6963);
xor U11877 (N_11877,N_6964,N_8399);
or U11878 (N_11878,N_6206,N_8075);
nor U11879 (N_11879,N_7981,N_8272);
nand U11880 (N_11880,N_7826,N_7756);
and U11881 (N_11881,N_7206,N_7905);
nand U11882 (N_11882,N_7486,N_6178);
nor U11883 (N_11883,N_8232,N_7296);
xnor U11884 (N_11884,N_6252,N_6237);
xor U11885 (N_11885,N_7012,N_8869);
nor U11886 (N_11886,N_7039,N_8667);
and U11887 (N_11887,N_7495,N_6727);
xor U11888 (N_11888,N_7912,N_7328);
xor U11889 (N_11889,N_8379,N_8682);
nand U11890 (N_11890,N_8977,N_6182);
nand U11891 (N_11891,N_8850,N_8911);
nor U11892 (N_11892,N_8593,N_6548);
nand U11893 (N_11893,N_8549,N_7781);
and U11894 (N_11894,N_6597,N_6378);
nor U11895 (N_11895,N_8893,N_6108);
or U11896 (N_11896,N_8243,N_7584);
or U11897 (N_11897,N_6489,N_8941);
or U11898 (N_11898,N_8743,N_7097);
nor U11899 (N_11899,N_8856,N_7937);
and U11900 (N_11900,N_8110,N_7274);
xnor U11901 (N_11901,N_7180,N_7840);
xnor U11902 (N_11902,N_6616,N_8073);
nor U11903 (N_11903,N_7176,N_6063);
and U11904 (N_11904,N_6583,N_6679);
and U11905 (N_11905,N_8194,N_7391);
nand U11906 (N_11906,N_8299,N_8741);
nor U11907 (N_11907,N_8488,N_6770);
or U11908 (N_11908,N_8505,N_7278);
nor U11909 (N_11909,N_7210,N_7081);
nand U11910 (N_11910,N_8671,N_7110);
xor U11911 (N_11911,N_8324,N_6219);
nand U11912 (N_11912,N_7392,N_6844);
xor U11913 (N_11913,N_7468,N_7970);
xnor U11914 (N_11914,N_8287,N_6070);
nand U11915 (N_11915,N_6967,N_8424);
xnor U11916 (N_11916,N_8632,N_7526);
and U11917 (N_11917,N_7694,N_8166);
xnor U11918 (N_11918,N_6276,N_6698);
nand U11919 (N_11919,N_8111,N_8453);
and U11920 (N_11920,N_8198,N_7620);
xnor U11921 (N_11921,N_6778,N_6106);
nand U11922 (N_11922,N_6579,N_7918);
or U11923 (N_11923,N_7023,N_8377);
xor U11924 (N_11924,N_8937,N_6663);
or U11925 (N_11925,N_7149,N_6624);
nor U11926 (N_11926,N_8161,N_6456);
and U11927 (N_11927,N_7418,N_6640);
nand U11928 (N_11928,N_8370,N_6234);
xor U11929 (N_11929,N_8088,N_7559);
nor U11930 (N_11930,N_8507,N_8138);
and U11931 (N_11931,N_6422,N_7145);
and U11932 (N_11932,N_7076,N_8086);
or U11933 (N_11933,N_7645,N_6047);
xnor U11934 (N_11934,N_7284,N_8539);
or U11935 (N_11935,N_7601,N_7064);
nand U11936 (N_11936,N_8448,N_7386);
nand U11937 (N_11937,N_6956,N_6474);
xor U11938 (N_11938,N_6563,N_7366);
and U11939 (N_11939,N_8107,N_6329);
and U11940 (N_11940,N_8825,N_8832);
nand U11941 (N_11941,N_8844,N_7672);
and U11942 (N_11942,N_6186,N_7123);
nand U11943 (N_11943,N_6425,N_7078);
xor U11944 (N_11944,N_7101,N_8581);
nor U11945 (N_11945,N_8326,N_7475);
and U11946 (N_11946,N_6238,N_8157);
nor U11947 (N_11947,N_8697,N_8687);
and U11948 (N_11948,N_6477,N_7340);
xnor U11949 (N_11949,N_7868,N_8404);
nor U11950 (N_11950,N_6136,N_7646);
xnor U11951 (N_11951,N_8636,N_7151);
or U11952 (N_11952,N_7914,N_7833);
and U11953 (N_11953,N_7063,N_7281);
nor U11954 (N_11954,N_6788,N_8969);
xnor U11955 (N_11955,N_8472,N_6993);
xor U11956 (N_11956,N_6720,N_6019);
nor U11957 (N_11957,N_6729,N_8458);
nor U11958 (N_11958,N_6291,N_6632);
and U11959 (N_11959,N_7531,N_7054);
and U11960 (N_11960,N_8453,N_6407);
nor U11961 (N_11961,N_6943,N_7699);
or U11962 (N_11962,N_8132,N_8416);
xor U11963 (N_11963,N_8055,N_6497);
and U11964 (N_11964,N_6725,N_6520);
or U11965 (N_11965,N_6801,N_7865);
xnor U11966 (N_11966,N_8720,N_6466);
xnor U11967 (N_11967,N_6925,N_8161);
and U11968 (N_11968,N_8321,N_8224);
and U11969 (N_11969,N_6593,N_6173);
and U11970 (N_11970,N_8204,N_7041);
nand U11971 (N_11971,N_6092,N_8414);
nand U11972 (N_11972,N_6773,N_8803);
or U11973 (N_11973,N_6367,N_7011);
and U11974 (N_11974,N_6713,N_8551);
nand U11975 (N_11975,N_7237,N_8856);
xor U11976 (N_11976,N_7325,N_8600);
xnor U11977 (N_11977,N_8273,N_6987);
nand U11978 (N_11978,N_7435,N_8433);
nand U11979 (N_11979,N_7341,N_8035);
nor U11980 (N_11980,N_8406,N_6768);
xor U11981 (N_11981,N_7480,N_7415);
nand U11982 (N_11982,N_6010,N_7400);
and U11983 (N_11983,N_7363,N_8704);
xnor U11984 (N_11984,N_8074,N_8400);
xnor U11985 (N_11985,N_6975,N_7875);
and U11986 (N_11986,N_8082,N_8972);
nand U11987 (N_11987,N_8171,N_7993);
or U11988 (N_11988,N_8047,N_8901);
xnor U11989 (N_11989,N_7372,N_6232);
nor U11990 (N_11990,N_6657,N_8190);
xor U11991 (N_11991,N_6922,N_7102);
nor U11992 (N_11992,N_7274,N_7073);
and U11993 (N_11993,N_6932,N_6197);
and U11994 (N_11994,N_7921,N_7407);
or U11995 (N_11995,N_6558,N_7080);
or U11996 (N_11996,N_8204,N_7841);
or U11997 (N_11997,N_6352,N_6077);
nand U11998 (N_11998,N_7755,N_7941);
xnor U11999 (N_11999,N_8815,N_7378);
or U12000 (N_12000,N_9440,N_10340);
nor U12001 (N_12001,N_11649,N_11100);
nand U12002 (N_12002,N_10166,N_11782);
xnor U12003 (N_12003,N_9639,N_10032);
nor U12004 (N_12004,N_10000,N_10426);
nand U12005 (N_12005,N_9545,N_11970);
nor U12006 (N_12006,N_10809,N_11459);
and U12007 (N_12007,N_10288,N_11546);
xor U12008 (N_12008,N_9073,N_9830);
or U12009 (N_12009,N_10037,N_11984);
or U12010 (N_12010,N_10967,N_9121);
or U12011 (N_12011,N_10041,N_11929);
or U12012 (N_12012,N_11201,N_9862);
and U12013 (N_12013,N_9857,N_9616);
nand U12014 (N_12014,N_10575,N_11237);
nand U12015 (N_12015,N_11294,N_11739);
nand U12016 (N_12016,N_10866,N_11851);
nor U12017 (N_12017,N_9134,N_11961);
xor U12018 (N_12018,N_11416,N_11230);
xor U12019 (N_12019,N_11058,N_11719);
nand U12020 (N_12020,N_9676,N_9068);
nand U12021 (N_12021,N_10714,N_11919);
or U12022 (N_12022,N_9125,N_10752);
nor U12023 (N_12023,N_9624,N_10653);
or U12024 (N_12024,N_10318,N_9167);
or U12025 (N_12025,N_9299,N_11872);
nor U12026 (N_12026,N_11926,N_10349);
and U12027 (N_12027,N_10883,N_9426);
xnor U12028 (N_12028,N_9209,N_10030);
xnor U12029 (N_12029,N_9527,N_10603);
nand U12030 (N_12030,N_9228,N_10027);
nand U12031 (N_12031,N_10812,N_11659);
nor U12032 (N_12032,N_9765,N_10211);
and U12033 (N_12033,N_10573,N_11461);
xor U12034 (N_12034,N_11270,N_10673);
nor U12035 (N_12035,N_10863,N_11381);
nand U12036 (N_12036,N_10501,N_9164);
or U12037 (N_12037,N_10721,N_11646);
nor U12038 (N_12038,N_9985,N_9280);
nor U12039 (N_12039,N_9013,N_9691);
nand U12040 (N_12040,N_9330,N_9204);
xor U12041 (N_12041,N_11091,N_9022);
or U12042 (N_12042,N_10710,N_11636);
and U12043 (N_12043,N_9752,N_9455);
or U12044 (N_12044,N_9343,N_10947);
nor U12045 (N_12045,N_10156,N_9700);
xnor U12046 (N_12046,N_9395,N_9664);
xor U12047 (N_12047,N_10221,N_11401);
and U12048 (N_12048,N_9914,N_10567);
nor U12049 (N_12049,N_9482,N_10640);
and U12050 (N_12050,N_10429,N_11253);
or U12051 (N_12051,N_11802,N_11738);
nor U12052 (N_12052,N_10989,N_11674);
or U12053 (N_12053,N_11409,N_10043);
nand U12054 (N_12054,N_10411,N_9520);
nor U12055 (N_12055,N_10216,N_9655);
and U12056 (N_12056,N_11785,N_11711);
xor U12057 (N_12057,N_10851,N_9900);
and U12058 (N_12058,N_11562,N_10317);
xor U12059 (N_12059,N_9665,N_10869);
nor U12060 (N_12060,N_10615,N_10168);
and U12061 (N_12061,N_11937,N_10888);
or U12062 (N_12062,N_10786,N_11763);
or U12063 (N_12063,N_10552,N_10528);
nand U12064 (N_12064,N_10960,N_11330);
nand U12065 (N_12065,N_11614,N_9881);
nand U12066 (N_12066,N_11819,N_10337);
nor U12067 (N_12067,N_9709,N_9263);
or U12068 (N_12068,N_10824,N_9838);
xnor U12069 (N_12069,N_11348,N_9064);
nand U12070 (N_12070,N_10572,N_10867);
nor U12071 (N_12071,N_9824,N_9433);
xor U12072 (N_12072,N_9511,N_9849);
or U12073 (N_12073,N_11542,N_10008);
nand U12074 (N_12074,N_10144,N_10180);
or U12075 (N_12075,N_9138,N_11626);
and U12076 (N_12076,N_10915,N_11104);
and U12077 (N_12077,N_10601,N_11177);
or U12078 (N_12078,N_10988,N_11506);
xor U12079 (N_12079,N_11988,N_11033);
nor U12080 (N_12080,N_11728,N_9126);
xnor U12081 (N_12081,N_9226,N_11315);
xor U12082 (N_12082,N_10397,N_11087);
nor U12083 (N_12083,N_9929,N_11193);
nand U12084 (N_12084,N_11223,N_11466);
and U12085 (N_12085,N_10483,N_11267);
or U12086 (N_12086,N_10647,N_10906);
nor U12087 (N_12087,N_11020,N_9858);
or U12088 (N_12088,N_11602,N_10806);
nand U12089 (N_12089,N_10649,N_10686);
nand U12090 (N_12090,N_9763,N_11651);
xor U12091 (N_12091,N_11697,N_11999);
nand U12092 (N_12092,N_11972,N_11685);
and U12093 (N_12093,N_10197,N_11451);
xnor U12094 (N_12094,N_11879,N_9633);
nand U12095 (N_12095,N_11203,N_11307);
and U12096 (N_12096,N_11120,N_9649);
and U12097 (N_12097,N_11118,N_11301);
and U12098 (N_12098,N_10245,N_9724);
xor U12099 (N_12099,N_10362,N_11303);
or U12100 (N_12100,N_11245,N_11045);
xor U12101 (N_12101,N_11325,N_11268);
and U12102 (N_12102,N_10038,N_11340);
or U12103 (N_12103,N_9868,N_10305);
xor U12104 (N_12104,N_9074,N_10323);
and U12105 (N_12105,N_10777,N_9778);
xor U12106 (N_12106,N_10466,N_10918);
nor U12107 (N_12107,N_9019,N_9034);
nor U12108 (N_12108,N_11948,N_11582);
nand U12109 (N_12109,N_10847,N_10013);
nand U12110 (N_12110,N_9173,N_11904);
and U12111 (N_12111,N_11577,N_10258);
or U12112 (N_12112,N_10623,N_11527);
or U12113 (N_12113,N_11210,N_11310);
nand U12114 (N_12114,N_11709,N_11876);
nor U12115 (N_12115,N_10844,N_9131);
or U12116 (N_12116,N_10113,N_11629);
nor U12117 (N_12117,N_11313,N_9158);
or U12118 (N_12118,N_11573,N_10100);
or U12119 (N_12119,N_9947,N_9523);
or U12120 (N_12120,N_10331,N_11766);
or U12121 (N_12121,N_10188,N_9365);
nor U12122 (N_12122,N_11930,N_11918);
nor U12123 (N_12123,N_9350,N_9797);
nand U12124 (N_12124,N_9287,N_11593);
nand U12125 (N_12125,N_10772,N_9327);
nand U12126 (N_12126,N_9853,N_11551);
nor U12127 (N_12127,N_11894,N_9470);
xnor U12128 (N_12128,N_11634,N_10415);
nand U12129 (N_12129,N_10205,N_11842);
and U12130 (N_12130,N_9311,N_10252);
xor U12131 (N_12131,N_11680,N_11367);
nand U12132 (N_12132,N_9057,N_10941);
nand U12133 (N_12133,N_10278,N_9518);
xor U12134 (N_12134,N_9419,N_11262);
xor U12135 (N_12135,N_9532,N_10808);
nor U12136 (N_12136,N_9092,N_9932);
or U12137 (N_12137,N_10176,N_10478);
and U12138 (N_12138,N_11947,N_9420);
and U12139 (N_12139,N_10994,N_11714);
nor U12140 (N_12140,N_10834,N_11713);
nand U12141 (N_12141,N_11533,N_10875);
nand U12142 (N_12142,N_11922,N_11150);
nor U12143 (N_12143,N_9669,N_10021);
and U12144 (N_12144,N_9203,N_9850);
and U12145 (N_12145,N_11304,N_9104);
and U12146 (N_12146,N_11579,N_11457);
nor U12147 (N_12147,N_11857,N_10063);
xor U12148 (N_12148,N_9942,N_10081);
or U12149 (N_12149,N_10525,N_10914);
xor U12150 (N_12150,N_11271,N_9854);
or U12151 (N_12151,N_10079,N_9609);
and U12152 (N_12152,N_11965,N_9811);
and U12153 (N_12153,N_9539,N_9396);
nor U12154 (N_12154,N_9562,N_11339);
and U12155 (N_12155,N_10890,N_10213);
nor U12156 (N_12156,N_10486,N_9613);
xor U12157 (N_12157,N_11165,N_9690);
and U12158 (N_12158,N_11326,N_10532);
or U12159 (N_12159,N_9447,N_11356);
nor U12160 (N_12160,N_11027,N_9494);
nand U12161 (N_12161,N_11050,N_11153);
nand U12162 (N_12162,N_10018,N_10031);
nor U12163 (N_12163,N_10745,N_11891);
and U12164 (N_12164,N_11638,N_11928);
nand U12165 (N_12165,N_11895,N_10419);
nand U12166 (N_12166,N_10167,N_9042);
nor U12167 (N_12167,N_11694,N_9187);
or U12168 (N_12168,N_9959,N_10660);
nor U12169 (N_12169,N_11426,N_10028);
nor U12170 (N_12170,N_11693,N_11154);
xor U12171 (N_12171,N_10073,N_11324);
or U12172 (N_12172,N_10292,N_11557);
and U12173 (N_12173,N_11232,N_9493);
nor U12174 (N_12174,N_10789,N_9973);
nand U12175 (N_12175,N_9356,N_11881);
or U12176 (N_12176,N_11216,N_11159);
nor U12177 (N_12177,N_10823,N_11822);
nor U12178 (N_12178,N_11102,N_11034);
nand U12179 (N_12179,N_9958,N_9738);
or U12180 (N_12180,N_11239,N_11944);
and U12181 (N_12181,N_9542,N_11804);
or U12182 (N_12182,N_9040,N_11215);
nand U12183 (N_12183,N_10974,N_9546);
and U12184 (N_12184,N_9867,N_10129);
xnor U12185 (N_12185,N_9557,N_11060);
nor U12186 (N_12186,N_9784,N_9317);
nand U12187 (N_12187,N_11521,N_10282);
or U12188 (N_12188,N_9645,N_10407);
xnor U12189 (N_12189,N_11513,N_11700);
or U12190 (N_12190,N_9840,N_9109);
or U12191 (N_12191,N_9928,N_9364);
xor U12192 (N_12192,N_10227,N_10469);
nand U12193 (N_12193,N_10428,N_10629);
nand U12194 (N_12194,N_10372,N_10384);
nand U12195 (N_12195,N_10519,N_9988);
nand U12196 (N_12196,N_9878,N_10247);
and U12197 (N_12197,N_9592,N_9439);
nand U12198 (N_12198,N_11587,N_10161);
nor U12199 (N_12199,N_11666,N_10695);
and U12200 (N_12200,N_10099,N_9253);
nor U12201 (N_12201,N_11250,N_10708);
and U12202 (N_12202,N_11632,N_11379);
nand U12203 (N_12203,N_9171,N_10389);
nand U12204 (N_12204,N_10973,N_10942);
or U12205 (N_12205,N_10932,N_11292);
or U12206 (N_12206,N_10706,N_11204);
nand U12207 (N_12207,N_11344,N_11959);
nor U12208 (N_12208,N_10594,N_11962);
or U12209 (N_12209,N_9047,N_9653);
xnor U12210 (N_12210,N_11143,N_11350);
or U12211 (N_12211,N_9197,N_11181);
nand U12212 (N_12212,N_11195,N_9175);
xor U12213 (N_12213,N_9247,N_11996);
and U12214 (N_12214,N_9681,N_9835);
and U12215 (N_12215,N_10271,N_11067);
xor U12216 (N_12216,N_9291,N_9541);
nand U12217 (N_12217,N_10223,N_10754);
and U12218 (N_12218,N_11142,N_11683);
or U12219 (N_12219,N_10052,N_11093);
or U12220 (N_12220,N_9575,N_9926);
nor U12221 (N_12221,N_9847,N_9190);
or U12222 (N_12222,N_11661,N_11125);
or U12223 (N_12223,N_10365,N_11731);
and U12224 (N_12224,N_10001,N_11920);
nor U12225 (N_12225,N_9295,N_10566);
or U12226 (N_12226,N_10103,N_11859);
nor U12227 (N_12227,N_9274,N_11349);
nor U12228 (N_12228,N_10122,N_10529);
and U12229 (N_12229,N_10451,N_10533);
or U12230 (N_12230,N_9646,N_9922);
nand U12231 (N_12231,N_9904,N_11371);
or U12232 (N_12232,N_9048,N_11830);
nand U12233 (N_12233,N_9003,N_10599);
xnor U12234 (N_12234,N_9901,N_9252);
or U12235 (N_12235,N_10865,N_11425);
or U12236 (N_12236,N_11180,N_11064);
xnor U12237 (N_12237,N_9516,N_9314);
nand U12238 (N_12238,N_11952,N_9597);
nor U12239 (N_12239,N_9035,N_11380);
nand U12240 (N_12240,N_11537,N_10404);
and U12241 (N_12241,N_11158,N_11853);
xnor U12242 (N_12242,N_9787,N_9895);
and U12243 (N_12243,N_9186,N_11721);
nand U12244 (N_12244,N_11848,N_10402);
xor U12245 (N_12245,N_9483,N_11075);
nor U12246 (N_12246,N_11943,N_11498);
or U12247 (N_12247,N_9451,N_9711);
nand U12248 (N_12248,N_9355,N_11799);
xnor U12249 (N_12249,N_10782,N_10321);
xnor U12250 (N_12250,N_10509,N_11431);
xor U12251 (N_12251,N_11096,N_9033);
xnor U12252 (N_12252,N_9225,N_9010);
nor U12253 (N_12253,N_10713,N_10148);
and U12254 (N_12254,N_11905,N_10217);
nand U12255 (N_12255,N_11317,N_10226);
and U12256 (N_12256,N_11890,N_9999);
nand U12257 (N_12257,N_9931,N_9231);
or U12258 (N_12258,N_9256,N_11565);
or U12259 (N_12259,N_10393,N_9887);
and U12260 (N_12260,N_9678,N_9662);
nor U12261 (N_12261,N_11227,N_9406);
xnor U12262 (N_12262,N_9168,N_9250);
or U12263 (N_12263,N_10412,N_11524);
nor U12264 (N_12264,N_10667,N_9829);
nor U12265 (N_12265,N_9178,N_9208);
and U12266 (N_12266,N_10473,N_10837);
nand U12267 (N_12267,N_11559,N_11529);
nand U12268 (N_12268,N_11287,N_11433);
or U12269 (N_12269,N_11811,N_11809);
nand U12270 (N_12270,N_11375,N_9336);
or U12271 (N_12271,N_11743,N_10881);
nand U12272 (N_12272,N_9332,N_11188);
or U12273 (N_12273,N_9983,N_9737);
and U12274 (N_12274,N_11191,N_9870);
nand U12275 (N_12275,N_11411,N_9257);
nand U12276 (N_12276,N_11089,N_10380);
xor U12277 (N_12277,N_10361,N_11974);
or U12278 (N_12278,N_9462,N_10904);
nor U12279 (N_12279,N_11949,N_10984);
nand U12280 (N_12280,N_10265,N_9487);
xor U12281 (N_12281,N_9801,N_9227);
nor U12282 (N_12282,N_11917,N_11778);
nor U12283 (N_12283,N_10938,N_9303);
and U12284 (N_12284,N_9563,N_10878);
xor U12285 (N_12285,N_11211,N_9151);
and U12286 (N_12286,N_11532,N_11915);
and U12287 (N_12287,N_9558,N_9725);
xor U12288 (N_12288,N_10071,N_9316);
nor U12289 (N_12289,N_11885,N_9195);
or U12290 (N_12290,N_11718,N_9113);
nand U12291 (N_12291,N_11708,N_10900);
and U12292 (N_12292,N_11690,N_9605);
nor U12293 (N_12293,N_11733,N_10759);
nand U12294 (N_12294,N_11376,N_9372);
nor U12295 (N_12295,N_11660,N_10933);
nand U12296 (N_12296,N_9800,N_11276);
and U12297 (N_12297,N_11953,N_11222);
nand U12298 (N_12298,N_9803,N_10804);
or U12299 (N_12299,N_10236,N_11906);
xnor U12300 (N_12300,N_9969,N_9436);
or U12301 (N_12301,N_10325,N_9990);
and U12302 (N_12302,N_10876,N_9307);
and U12303 (N_12303,N_11595,N_10554);
or U12304 (N_12304,N_9907,N_11497);
and U12305 (N_12305,N_10283,N_11128);
and U12306 (N_12306,N_10756,N_11190);
nand U12307 (N_12307,N_10978,N_11363);
or U12308 (N_12308,N_11553,N_10198);
nand U12309 (N_12309,N_11535,N_9943);
nor U12310 (N_12310,N_11530,N_9792);
nand U12311 (N_12311,N_10657,N_9590);
or U12312 (N_12312,N_9020,N_11921);
xnor U12313 (N_12313,N_11662,N_10681);
and U12314 (N_12314,N_10608,N_10704);
nand U12315 (N_12315,N_9385,N_10518);
nor U12316 (N_12316,N_11074,N_10555);
nand U12317 (N_12317,N_10231,N_11572);
nor U12318 (N_12318,N_10889,N_11892);
or U12319 (N_12319,N_11954,N_10650);
xnor U12320 (N_12320,N_9561,N_10576);
or U12321 (N_12321,N_11980,N_10956);
and U12322 (N_12322,N_9415,N_11775);
nand U12323 (N_12323,N_9775,N_9052);
and U12324 (N_12324,N_11162,N_9018);
or U12325 (N_12325,N_9755,N_10208);
nor U12326 (N_12326,N_11789,N_11194);
xor U12327 (N_12327,N_10320,N_10836);
nand U12328 (N_12328,N_10955,N_11772);
or U12329 (N_12329,N_9255,N_11950);
xnor U12330 (N_12330,N_10753,N_11092);
and U12331 (N_12331,N_10443,N_9438);
nand U12332 (N_12332,N_11297,N_11351);
xnor U12333 (N_12333,N_11520,N_9923);
xor U12334 (N_12334,N_11456,N_11070);
xor U12335 (N_12335,N_10302,N_11273);
or U12336 (N_12336,N_11185,N_10537);
nor U12337 (N_12337,N_11453,N_11810);
nand U12338 (N_12338,N_9242,N_11359);
and U12339 (N_12339,N_9086,N_10577);
nor U12340 (N_12340,N_9703,N_10774);
xnor U12341 (N_12341,N_11938,N_11698);
xor U12342 (N_12342,N_10170,N_9341);
xnor U12343 (N_12343,N_9993,N_9089);
nand U12344 (N_12344,N_11011,N_9407);
xnor U12345 (N_12345,N_11609,N_9729);
nor U12346 (N_12346,N_9697,N_11392);
nand U12347 (N_12347,N_11327,N_11839);
and U12348 (N_12348,N_11318,N_9181);
xor U12349 (N_12349,N_10948,N_11654);
xnor U12350 (N_12350,N_10687,N_10061);
nor U12351 (N_12351,N_11244,N_10017);
or U12352 (N_12352,N_9404,N_10585);
nand U12353 (N_12353,N_9855,N_10489);
nor U12354 (N_12354,N_10606,N_10445);
or U12355 (N_12355,N_11114,N_11445);
and U12356 (N_12356,N_11862,N_10831);
and U12357 (N_12357,N_10237,N_10734);
or U12358 (N_12358,N_9754,N_11823);
or U12359 (N_12359,N_11975,N_9095);
nor U12360 (N_12360,N_9917,N_11323);
nand U12361 (N_12361,N_9704,N_10453);
nand U12362 (N_12362,N_9476,N_10479);
xnor U12363 (N_12363,N_9304,N_10634);
xnor U12364 (N_12364,N_11419,N_10935);
nor U12365 (N_12365,N_9996,N_11333);
nor U12366 (N_12366,N_11995,N_10140);
xor U12367 (N_12367,N_11669,N_10444);
or U12368 (N_12368,N_9179,N_9381);
nand U12369 (N_12369,N_9566,N_9046);
nor U12370 (N_12370,N_10097,N_10977);
and U12371 (N_12371,N_10467,N_10279);
or U12372 (N_12372,N_9460,N_10244);
or U12373 (N_12373,N_11979,N_9261);
nand U12374 (N_12374,N_11540,N_10474);
or U12375 (N_12375,N_10626,N_11771);
nor U12376 (N_12376,N_10674,N_11347);
nand U12377 (N_12377,N_10589,N_9601);
or U12378 (N_12378,N_10506,N_10239);
xnor U12379 (N_12379,N_10654,N_10996);
or U12380 (N_12380,N_11820,N_9962);
or U12381 (N_12381,N_9919,N_10382);
or U12382 (N_12382,N_10461,N_9182);
nand U12383 (N_12383,N_10979,N_10424);
or U12384 (N_12384,N_11645,N_10084);
nor U12385 (N_12385,N_10108,N_9667);
nor U12386 (N_12386,N_9631,N_11973);
and U12387 (N_12387,N_10701,N_9686);
and U12388 (N_12388,N_9534,N_9863);
xor U12389 (N_12389,N_11960,N_9389);
xor U12390 (N_12390,N_10338,N_11834);
xor U12391 (N_12391,N_11840,N_10294);
and U12392 (N_12392,N_11914,N_9454);
nand U12393 (N_12393,N_11212,N_9500);
and U12394 (N_12394,N_11808,N_10187);
xnor U12395 (N_12395,N_9169,N_10946);
or U12396 (N_12396,N_9856,N_9379);
xor U12397 (N_12397,N_10276,N_10791);
and U12398 (N_12398,N_11776,N_9145);
xnor U12399 (N_12399,N_9489,N_11171);
xnor U12400 (N_12400,N_9107,N_9465);
nand U12401 (N_12401,N_9568,N_10926);
nor U12402 (N_12402,N_11243,N_10742);
xnor U12403 (N_12403,N_11168,N_10307);
nand U12404 (N_12404,N_10718,N_10363);
nand U12405 (N_12405,N_10559,N_9206);
and U12406 (N_12406,N_9553,N_11336);
or U12407 (N_12407,N_11389,N_11902);
nand U12408 (N_12408,N_9258,N_9490);
xor U12409 (N_12409,N_9744,N_9728);
nor U12410 (N_12410,N_10551,N_9425);
nor U12411 (N_12411,N_10449,N_9194);
or U12412 (N_12412,N_11173,N_11044);
nor U12413 (N_12413,N_11696,N_11130);
nand U12414 (N_12414,N_9521,N_10193);
nor U12415 (N_12415,N_10007,N_11751);
xnor U12416 (N_12416,N_9449,N_11338);
xor U12417 (N_12417,N_9920,N_9589);
and U12418 (N_12418,N_11394,N_9444);
nor U12419 (N_12419,N_11023,N_10229);
nor U12420 (N_12420,N_9758,N_11755);
nor U12421 (N_12421,N_10376,N_11653);
xnor U12422 (N_12422,N_11838,N_10431);
nand U12423 (N_12423,N_10123,N_11555);
xor U12424 (N_12424,N_9069,N_11507);
nor U12425 (N_12425,N_10503,N_10499);
xnor U12426 (N_12426,N_10699,N_10709);
or U12427 (N_12427,N_10126,N_9743);
xor U12428 (N_12428,N_11071,N_9484);
and U12429 (N_12429,N_11600,N_11489);
nand U12430 (N_12430,N_9882,N_10785);
xnor U12431 (N_12431,N_9891,N_10711);
and U12432 (N_12432,N_9051,N_9071);
or U12433 (N_12433,N_9132,N_10983);
and U12434 (N_12434,N_10970,N_11812);
nor U12435 (N_12435,N_10417,N_11737);
xor U12436 (N_12436,N_10535,N_9525);
or U12437 (N_12437,N_10818,N_11467);
or U12438 (N_12438,N_10997,N_10563);
nand U12439 (N_12439,N_9995,N_9495);
nand U12440 (N_12440,N_10300,N_9344);
or U12441 (N_12441,N_9359,N_10348);
or U12442 (N_12442,N_10086,N_10420);
nor U12443 (N_12443,N_11406,N_10998);
nand U12444 (N_12444,N_9997,N_9417);
nand U12445 (N_12445,N_11783,N_9320);
nand U12446 (N_12446,N_9129,N_11824);
nand U12447 (N_12447,N_9224,N_9550);
and U12448 (N_12448,N_10848,N_11736);
or U12449 (N_12449,N_9611,N_11945);
xnor U12450 (N_12450,N_11676,N_10620);
nand U12451 (N_12451,N_9049,N_10976);
xor U12452 (N_12452,N_10940,N_11382);
and U12453 (N_12453,N_11396,N_9302);
and U12454 (N_12454,N_11288,N_9706);
and U12455 (N_12455,N_9230,N_9952);
nor U12456 (N_12456,N_11004,N_9458);
nand U12457 (N_12457,N_9726,N_10342);
or U12458 (N_12458,N_9687,N_10735);
nor U12459 (N_12459,N_9079,N_11368);
or U12460 (N_12460,N_11679,N_10690);
and U12461 (N_12461,N_11441,N_9422);
nor U12462 (N_12462,N_9098,N_9466);
and U12463 (N_12463,N_10512,N_9761);
nand U12464 (N_12464,N_11192,N_10134);
or U12465 (N_12465,N_10995,N_11205);
nand U12466 (N_12466,N_9955,N_9670);
nor U12467 (N_12467,N_10327,N_10481);
or U12468 (N_12468,N_10820,N_9289);
and U12469 (N_12469,N_10476,N_10700);
xnor U12470 (N_12470,N_11377,N_10862);
nor U12471 (N_12471,N_11576,N_11094);
and U12472 (N_12472,N_9939,N_10455);
nand U12473 (N_12473,N_11689,N_11552);
nand U12474 (N_12474,N_10157,N_10329);
nand U12475 (N_12475,N_9799,N_10261);
and U12476 (N_12476,N_9698,N_9428);
xor U12477 (N_12477,N_11051,N_11078);
or U12478 (N_12478,N_11152,N_11670);
and U12479 (N_12479,N_9298,N_9628);
nand U12480 (N_12480,N_9638,N_9409);
or U12481 (N_12481,N_11101,N_11309);
and U12482 (N_12482,N_10614,N_9220);
or U12483 (N_12483,N_10006,N_9342);
xnor U12484 (N_12484,N_10556,N_11258);
or U12485 (N_12485,N_11671,N_9960);
nor U12486 (N_12486,N_9281,N_9282);
nor U12487 (N_12487,N_11833,N_9083);
nor U12488 (N_12488,N_11502,N_10816);
or U12489 (N_12489,N_9037,N_11306);
and U12490 (N_12490,N_10858,N_11813);
xnor U12491 (N_12491,N_10720,N_11873);
nand U12492 (N_12492,N_9360,N_9573);
and U12493 (N_12493,N_9654,N_10843);
xnor U12494 (N_12494,N_11657,N_10500);
or U12495 (N_12495,N_10313,N_10901);
xor U12496 (N_12496,N_10328,N_10788);
or U12497 (N_12497,N_9938,N_11934);
xor U12498 (N_12498,N_10138,N_10927);
or U12499 (N_12499,N_9598,N_9762);
or U12500 (N_12500,N_10177,N_11725);
nor U12501 (N_12501,N_9100,N_11642);
xnor U12502 (N_12502,N_9093,N_10290);
nor U12503 (N_12503,N_10255,N_9883);
and U12504 (N_12504,N_10341,N_10475);
nand U12505 (N_12505,N_9632,N_10104);
nor U12506 (N_12506,N_11059,N_10128);
nand U12507 (N_12507,N_10204,N_11247);
xor U12508 (N_12508,N_9576,N_9629);
and U12509 (N_12509,N_9140,N_11568);
and U12510 (N_12510,N_9453,N_11706);
xnor U12511 (N_12511,N_10838,N_11856);
xor U12512 (N_12512,N_10740,N_10980);
nand U12513 (N_12513,N_11978,N_10117);
xor U12514 (N_12514,N_10083,N_9822);
nor U12515 (N_12515,N_11598,N_10693);
nand U12516 (N_12516,N_11992,N_9467);
xnor U12517 (N_12517,N_10975,N_9702);
nor U12518 (N_12518,N_9199,N_11012);
or U12519 (N_12519,N_11283,N_10536);
xnor U12520 (N_12520,N_11429,N_10910);
nand U12521 (N_12521,N_11637,N_11298);
nor U12522 (N_12522,N_11983,N_11644);
nor U12523 (N_12523,N_9659,N_9397);
and U12524 (N_12524,N_9305,N_10845);
or U12525 (N_12525,N_11378,N_10639);
nand U12526 (N_12526,N_9688,N_9717);
nor U12527 (N_12527,N_11882,N_10521);
xor U12528 (N_12528,N_9567,N_11115);
xnor U12529 (N_12529,N_11724,N_11854);
nor U12530 (N_12530,N_9786,N_11608);
xnor U12531 (N_12531,N_10621,N_9866);
nand U12532 (N_12532,N_10702,N_11242);
nor U12533 (N_12533,N_10195,N_10403);
nor U12534 (N_12534,N_10142,N_11624);
nor U12535 (N_12535,N_11291,N_11462);
nor U12536 (N_12536,N_9423,N_11176);
xor U12537 (N_12537,N_11618,N_10301);
and U12538 (N_12538,N_10115,N_10335);
xor U12539 (N_12539,N_11987,N_10002);
nor U12540 (N_12540,N_9041,N_10581);
nand U12541 (N_12541,N_11985,N_10511);
nand U12542 (N_12542,N_10548,N_10215);
nor U12543 (N_12543,N_9477,N_10874);
and U12544 (N_12544,N_10541,N_10602);
or U12545 (N_12545,N_9223,N_9469);
xor U12546 (N_12546,N_9705,N_11554);
and U12547 (N_12547,N_9894,N_9971);
nand U12548 (N_12548,N_9643,N_10438);
xor U12549 (N_12549,N_11874,N_11069);
nand U12550 (N_12550,N_10540,N_9352);
or U12551 (N_12551,N_9833,N_11747);
nor U12552 (N_12552,N_11105,N_10539);
nor U12553 (N_12553,N_10648,N_10937);
nand U12554 (N_12554,N_11113,N_10643);
and U12555 (N_12555,N_11673,N_11365);
nand U12556 (N_12556,N_10102,N_11888);
or U12557 (N_12557,N_9021,N_10569);
or U12558 (N_12558,N_10171,N_9392);
and U12559 (N_12559,N_11030,N_9964);
and U12560 (N_12560,N_11005,N_11612);
nand U12561 (N_12561,N_10109,N_11219);
or U12562 (N_12562,N_9783,N_9127);
nor U12563 (N_12563,N_9414,N_11366);
nor U12564 (N_12564,N_9615,N_9239);
nor U12565 (N_12565,N_10055,N_11729);
or U12566 (N_12566,N_9940,N_10163);
or U12567 (N_12567,N_9346,N_10359);
or U12568 (N_12568,N_11131,N_11770);
xnor U12569 (N_12569,N_10087,N_10815);
xnor U12570 (N_12570,N_10886,N_11913);
xor U12571 (N_12571,N_11073,N_11218);
nand U12572 (N_12572,N_11599,N_9976);
or U12573 (N_12573,N_11014,N_9347);
or U12574 (N_12574,N_10136,N_11487);
nor U12575 (N_12575,N_9292,N_9549);
nand U12576 (N_12576,N_10413,N_9579);
nand U12577 (N_12577,N_9268,N_9512);
nor U12578 (N_12578,N_10224,N_10636);
or U12579 (N_12579,N_10641,N_11877);
xor U12580 (N_12580,N_11652,N_11329);
nand U12581 (N_12581,N_11296,N_10682);
or U12582 (N_12582,N_9585,N_9249);
nand U12583 (N_12583,N_10561,N_10972);
and U12584 (N_12584,N_10879,N_10607);
and U12585 (N_12585,N_9215,N_10155);
nand U12586 (N_12586,N_11925,N_9399);
nand U12587 (N_12587,N_11370,N_9871);
and U12588 (N_12588,N_9183,N_10295);
nor U12589 (N_12589,N_9080,N_11134);
nor U12590 (N_12590,N_9236,N_9810);
nand U12591 (N_12591,N_9004,N_9581);
or U12592 (N_12592,N_9766,N_9066);
nand U12593 (N_12593,N_10057,N_10923);
or U12594 (N_12594,N_9028,N_10352);
nand U12595 (N_12595,N_11641,N_11124);
or U12596 (N_12596,N_9806,N_11421);
xnor U12597 (N_12597,N_9637,N_11648);
nor U12598 (N_12598,N_11427,N_10736);
or U12599 (N_12599,N_10592,N_10374);
or U12600 (N_12600,N_10958,N_10291);
or U12601 (N_12601,N_11858,N_10746);
or U12602 (N_12602,N_11558,N_11111);
nor U12603 (N_12603,N_10762,N_10131);
and U12604 (N_12604,N_11076,N_9910);
xnor U12605 (N_12605,N_11787,N_9533);
nor U12606 (N_12606,N_10462,N_11119);
or U12607 (N_12607,N_9948,N_11534);
nor U12608 (N_12608,N_11797,N_9730);
nor U12609 (N_12609,N_10547,N_10056);
and U12610 (N_12610,N_10965,N_10578);
and U12611 (N_12611,N_9689,N_11903);
and U12612 (N_12612,N_10184,N_10894);
xnor U12613 (N_12613,N_9680,N_10270);
or U12614 (N_12614,N_9421,N_9953);
nand U12615 (N_12615,N_11932,N_11065);
nand U12616 (N_12616,N_10202,N_11607);
xnor U12617 (N_12617,N_10480,N_11161);
nor U12618 (N_12618,N_9832,N_10943);
and U12619 (N_12619,N_11850,N_9951);
and U12620 (N_12620,N_9890,N_11052);
and U12621 (N_12621,N_10873,N_11702);
or U12622 (N_12622,N_10827,N_10825);
and U12623 (N_12623,N_9393,N_10014);
nand U12624 (N_12624,N_9720,N_10574);
xor U12625 (N_12625,N_11164,N_10199);
and U12626 (N_12626,N_9027,N_9827);
or U12627 (N_12627,N_11767,N_11561);
xnor U12628 (N_12628,N_11290,N_9656);
nor U12629 (N_12629,N_10460,N_9536);
and U12630 (N_12630,N_9782,N_10936);
nand U12631 (N_12631,N_10768,N_9749);
xor U12632 (N_12632,N_9233,N_11682);
or U12633 (N_12633,N_9497,N_9275);
nor U12634 (N_12634,N_10093,N_11635);
nand U12635 (N_12635,N_11865,N_11256);
nor U12636 (N_12636,N_11897,N_9842);
and U12637 (N_12637,N_10659,N_10234);
and U12638 (N_12638,N_11765,N_11997);
nand U12639 (N_12639,N_9193,N_9005);
and U12640 (N_12640,N_9588,N_11864);
nand U12641 (N_12641,N_9159,N_11443);
and U12642 (N_12642,N_9087,N_10651);
or U12643 (N_12643,N_9620,N_9987);
or U12644 (N_12644,N_11571,N_9845);
nor U12645 (N_12645,N_11374,N_11884);
and U12646 (N_12646,N_11844,N_10810);
or U12647 (N_12647,N_10596,N_11490);
nor U12648 (N_12648,N_9157,N_9577);
xnor U12649 (N_12649,N_11605,N_10959);
nand U12650 (N_12650,N_9122,N_10304);
and U12651 (N_12651,N_11141,N_11174);
nand U12652 (N_12652,N_10584,N_9701);
nand U12653 (N_12653,N_10684,N_10619);
xor U12654 (N_12654,N_9816,N_9886);
or U12655 (N_12655,N_9506,N_10173);
nand U12656 (N_12656,N_11019,N_10726);
and U12657 (N_12657,N_10605,N_9499);
xor U12658 (N_12658,N_10683,N_9641);
xor U12659 (N_12659,N_9055,N_9229);
nor U12660 (N_12660,N_9361,N_10089);
or U12661 (N_12661,N_10609,N_9099);
xor U12662 (N_12662,N_10251,N_10091);
nor U12663 (N_12663,N_11432,N_10857);
and U12664 (N_12664,N_10829,N_11505);
nor U12665 (N_12665,N_10846,N_10246);
and U12666 (N_12666,N_11182,N_10395);
or U12667 (N_12667,N_11107,N_10441);
and U12668 (N_12668,N_9463,N_11900);
xnor U12669 (N_12669,N_10916,N_9039);
xor U12670 (N_12670,N_9285,N_10309);
and U12671 (N_12671,N_11342,N_11525);
and U12672 (N_12672,N_10414,N_11302);
nor U12673 (N_12673,N_10256,N_10871);
nor U12674 (N_12674,N_10580,N_11257);
nor U12675 (N_12675,N_9714,N_9510);
and U12676 (N_12676,N_11255,N_10744);
and U12677 (N_12677,N_10819,N_11870);
and U12678 (N_12678,N_11630,N_11048);
nand U12679 (N_12679,N_9374,N_11847);
xnor U12680 (N_12680,N_10066,N_10423);
nor U12681 (N_12681,N_10698,N_10840);
and U12682 (N_12682,N_11871,N_9739);
or U12683 (N_12683,N_10939,N_11939);
nor U12684 (N_12684,N_11035,N_9143);
nor U12685 (N_12685,N_10671,N_10542);
and U12686 (N_12686,N_11517,N_9216);
nor U12687 (N_12687,N_10730,N_10611);
or U12688 (N_12688,N_9219,N_9461);
xor U12689 (N_12689,N_9767,N_9719);
nor U12690 (N_12690,N_9693,N_10637);
or U12691 (N_12691,N_11077,N_10391);
xnor U12692 (N_12692,N_10464,N_11523);
or U12693 (N_12693,N_10053,N_10880);
xor U12694 (N_12694,N_10968,N_11135);
or U12695 (N_12695,N_9984,N_10147);
nand U12696 (N_12696,N_10892,N_10269);
nand U12697 (N_12697,N_9387,N_10920);
or U12698 (N_12698,N_10666,N_11664);
nor U12699 (N_12699,N_10333,N_9082);
and U12700 (N_12700,N_10044,N_9334);
nor U12701 (N_12701,N_11606,N_11748);
and U12702 (N_12702,N_11699,N_10371);
nand U12703 (N_12703,N_9750,N_11088);
nor U12704 (N_12704,N_11604,N_9986);
and U12705 (N_12705,N_10143,N_9614);
and U12706 (N_12706,N_10860,N_10897);
nor U12707 (N_12707,N_10549,N_11454);
xnor U12708 (N_12708,N_10792,N_9024);
nor U12709 (N_12709,N_10760,N_9012);
or U12710 (N_12710,N_10877,N_9437);
or U12711 (N_12711,N_9240,N_9682);
nor U12712 (N_12712,N_9481,N_9781);
nand U12713 (N_12713,N_10902,N_11354);
or U12714 (N_12714,N_11656,N_9551);
xor U12715 (N_12715,N_10612,N_10800);
and U12716 (N_12716,N_9528,N_11655);
nand U12717 (N_12717,N_10439,N_11663);
xnor U12718 (N_12718,N_9053,N_11956);
nand U12719 (N_12719,N_9630,N_11149);
nand U12720 (N_12720,N_11849,N_11701);
nor U12721 (N_12721,N_10078,N_10094);
and U12722 (N_12722,N_9635,N_9595);
nand U12723 (N_12723,N_9529,N_10421);
nand U12724 (N_12724,N_9991,N_11321);
xor U12725 (N_12725,N_9627,N_10757);
nand U12726 (N_12726,N_10763,N_10228);
nor U12727 (N_12727,N_9603,N_10530);
xor U12728 (N_12728,N_11183,N_11063);
and U12729 (N_12729,N_9309,N_10598);
and U12730 (N_12730,N_9294,N_9116);
and U12731 (N_12731,N_9232,N_11707);
xor U12732 (N_12732,N_11029,N_9464);
or U12733 (N_12733,N_11726,N_10952);
nand U12734 (N_12734,N_11252,N_10855);
or U12735 (N_12735,N_9443,N_10538);
nor U12736 (N_12736,N_11269,N_11951);
xnor U12737 (N_12737,N_9912,N_11860);
and U12738 (N_12738,N_9284,N_9565);
nor U12739 (N_12739,N_9110,N_10758);
nand U12740 (N_12740,N_9201,N_11675);
nor U12741 (N_12741,N_10822,N_10287);
and U12742 (N_12742,N_11758,N_9814);
nand U12743 (N_12743,N_10096,N_9058);
or U12744 (N_12744,N_11720,N_11199);
nor U12745 (N_12745,N_11829,N_11424);
nor U12746 (N_12746,N_10797,N_9478);
nand U12747 (N_12747,N_9288,N_9727);
and U12748 (N_12748,N_11079,N_10285);
xnor U12749 (N_12749,N_9760,N_11681);
nor U12750 (N_12750,N_11756,N_11584);
xnor U12751 (N_12751,N_11387,N_9410);
nor U12752 (N_12752,N_10151,N_9967);
and U12753 (N_12753,N_10343,N_11619);
xor U12754 (N_12754,N_9009,N_10493);
xor U12755 (N_12755,N_9780,N_11418);
and U12756 (N_12756,N_9424,N_10326);
nor U12757 (N_12757,N_11692,N_11967);
and U12758 (N_12758,N_11734,N_10924);
nor U12759 (N_12759,N_10303,N_11013);
or U12760 (N_12760,N_11621,N_11026);
or U12761 (N_12761,N_9380,N_9076);
or U12762 (N_12762,N_10872,N_10595);
or U12763 (N_12763,N_11556,N_11277);
nor U12764 (N_12764,N_11746,N_10390);
nor U12765 (N_12765,N_11438,N_9804);
nand U12766 (N_12766,N_10405,N_9474);
and U12767 (N_12767,N_10670,N_11509);
xor U12768 (N_12768,N_10765,N_9128);
or U12769 (N_12769,N_10111,N_11486);
nand U12770 (N_12770,N_10570,N_10842);
or U12771 (N_12771,N_9198,N_11826);
nand U12772 (N_12772,N_11494,N_11806);
nand U12773 (N_12773,N_11448,N_11062);
xor U12774 (N_12774,N_9696,N_10191);
xor U12775 (N_12775,N_11235,N_11761);
nand U12776 (N_12776,N_9898,N_9488);
and U12777 (N_12777,N_9559,N_11186);
and U12778 (N_12778,N_9507,N_11869);
nand U12779 (N_12779,N_9769,N_11145);
xnor U12780 (N_12780,N_9277,N_9248);
xor U12781 (N_12781,N_9308,N_10440);
nand U12782 (N_12782,N_11982,N_11249);
or U12783 (N_12783,N_11855,N_11570);
nand U12784 (N_12784,N_11966,N_11328);
nor U12785 (N_12785,N_9323,N_10495);
nand U12786 (N_12786,N_11022,N_11893);
or U12787 (N_12787,N_9555,N_9622);
or U12788 (N_12788,N_10150,N_9902);
nor U12789 (N_12789,N_11541,N_10350);
nor U12790 (N_12790,N_10381,N_11831);
or U12791 (N_12791,N_11796,N_9286);
nand U12792 (N_12792,N_9934,N_10488);
or U12793 (N_12793,N_11722,N_11184);
nand U12794 (N_12794,N_10766,N_9335);
nor U12795 (N_12795,N_10770,N_10379);
and U12796 (N_12796,N_9384,N_11442);
nand U12797 (N_12797,N_10121,N_9505);
and U12798 (N_12798,N_10023,N_9063);
nand U12799 (N_12799,N_9578,N_9596);
and U12800 (N_12800,N_9513,N_10811);
or U12801 (N_12801,N_9067,N_9954);
and U12802 (N_12802,N_11491,N_10345);
nand U12803 (N_12803,N_9981,N_9452);
xor U12804 (N_12804,N_11971,N_10020);
xor U12805 (N_12805,N_10491,N_9945);
xnor U12806 (N_12806,N_11678,N_10448);
xor U12807 (N_12807,N_11410,N_11788);
nand U12808 (N_12808,N_11007,N_10903);
nand U12809 (N_12809,N_10158,N_9032);
or U12810 (N_12810,N_11311,N_9106);
and U12811 (N_12811,N_9944,N_9710);
or U12812 (N_12812,N_11545,N_11485);
xor U12813 (N_12813,N_11479,N_11886);
and U12814 (N_12814,N_11055,N_10727);
and U12815 (N_12815,N_11408,N_10133);
or U12816 (N_12816,N_10394,N_10625);
nor U12817 (N_12817,N_11189,N_9339);
or U12818 (N_12818,N_11407,N_10799);
nand U12819 (N_12819,N_9222,N_11594);
or U12820 (N_12820,N_10468,N_10127);
xor U12821 (N_12821,N_9519,N_10330);
xnor U12822 (N_12822,N_11592,N_9166);
or U12823 (N_12823,N_10033,N_9570);
nor U12824 (N_12824,N_11197,N_10907);
xnor U12825 (N_12825,N_11358,N_9105);
or U12826 (N_12826,N_10494,N_10747);
nor U12827 (N_12827,N_11405,N_9675);
or U12828 (N_12828,N_10406,N_9679);
nor U12829 (N_12829,N_9587,N_11260);
or U12830 (N_12830,N_10985,N_9722);
xor U12831 (N_12831,N_10990,N_10787);
and U12832 (N_12832,N_11516,N_10112);
nor U12833 (N_12833,N_9259,N_10969);
and U12834 (N_12834,N_9176,N_10776);
nand U12835 (N_12835,N_11428,N_11832);
nor U12836 (N_12836,N_10262,N_10242);
xnor U12837 (N_12837,N_9353,N_9293);
and U12838 (N_12838,N_11550,N_10238);
and U12839 (N_12839,N_9877,N_9927);
or U12840 (N_12840,N_9218,N_11633);
nand U12841 (N_12841,N_9269,N_10314);
nor U12842 (N_12842,N_11898,N_11403);
xnor U12843 (N_12843,N_9879,N_10266);
and U12844 (N_12844,N_10891,N_9315);
nor U12845 (N_12845,N_11837,N_11388);
or U12846 (N_12846,N_10433,N_10010);
nor U12847 (N_12847,N_11295,N_9805);
nor U12848 (N_12848,N_11352,N_10324);
nand U12849 (N_12849,N_9191,N_10591);
or U12850 (N_12850,N_11417,N_9357);
and U12851 (N_12851,N_10691,N_11061);
nand U12852 (N_12852,N_11160,N_11108);
nor U12853 (N_12853,N_9322,N_9977);
nand U12854 (N_12854,N_9823,N_11493);
nand U12855 (N_12855,N_10731,N_10725);
nand U12856 (N_12856,N_11117,N_11278);
nand U12857 (N_12857,N_10531,N_9150);
or U12858 (N_12858,N_11780,N_9260);
nand U12859 (N_12859,N_9090,N_9924);
or U12860 (N_12860,N_10436,N_11266);
or U12861 (N_12861,N_10677,N_11519);
nand U12862 (N_12862,N_10470,N_11547);
xnor U12863 (N_12863,N_10807,N_10497);
or U12864 (N_12864,N_11384,N_10617);
xor U12865 (N_12865,N_11977,N_9272);
nor U12866 (N_12866,N_10045,N_11395);
or U12867 (N_12867,N_11081,N_10373);
or U12868 (N_12868,N_11046,N_9599);
nand U12869 (N_12869,N_9772,N_9607);
or U12870 (N_12870,N_11567,N_10964);
or U12871 (N_12871,N_11735,N_10597);
nor U12872 (N_12872,N_11248,N_10610);
nand U12873 (N_12873,N_10919,N_9774);
and U12874 (N_12874,N_10369,N_11792);
nor U12875 (N_12875,N_10738,N_11536);
nand U12876 (N_12876,N_9217,N_10425);
and U12877 (N_12877,N_11727,N_9707);
xnor U12878 (N_12878,N_10676,N_10813);
nor U12879 (N_12879,N_11597,N_11639);
xnor U12880 (N_12880,N_9980,N_11843);
or U12881 (N_12881,N_10986,N_11021);
nand U12882 (N_12882,N_9685,N_10418);
nor U12883 (N_12883,N_9663,N_10463);
xnor U12884 (N_12884,N_11156,N_10662);
and U12885 (N_12885,N_10296,N_9721);
nand U12886 (N_12886,N_10332,N_11238);
xor U12887 (N_12887,N_11715,N_10898);
or U12888 (N_12888,N_10259,N_10152);
nor U12889 (N_12889,N_11314,N_9376);
nand U12890 (N_12890,N_9837,N_10884);
and U12891 (N_12891,N_10859,N_9821);
and U12892 (N_12892,N_11450,N_10398);
nor U12893 (N_12893,N_10050,N_9779);
nor U12894 (N_12894,N_9974,N_9363);
xor U12895 (N_12895,N_10344,N_9695);
nand U12896 (N_12896,N_10230,N_11345);
or U12897 (N_12897,N_9537,N_10360);
and U12898 (N_12898,N_9283,N_11560);
and U12899 (N_12899,N_11279,N_11024);
xor U12900 (N_12900,N_10737,N_9556);
or U12901 (N_12901,N_10534,N_11151);
or U12902 (N_12902,N_11643,N_10856);
nor U12903 (N_12903,N_10067,N_9008);
xor U12904 (N_12904,N_10077,N_11814);
xnor U12905 (N_12905,N_9961,N_9747);
xor U12906 (N_12906,N_9941,N_10101);
xor U12907 (N_12907,N_11293,N_11460);
or U12908 (N_12908,N_9192,N_11226);
or U12909 (N_12909,N_10565,N_11110);
and U12910 (N_12910,N_9936,N_9016);
nand U12911 (N_12911,N_9809,N_9030);
nand U12912 (N_12912,N_11001,N_10917);
xor U12913 (N_12913,N_9300,N_10750);
xor U12914 (N_12914,N_10210,N_10739);
nor U12915 (N_12915,N_10656,N_11566);
nand U12916 (N_12916,N_9813,N_10257);
and U12917 (N_12917,N_9059,N_11139);
nand U12918 (N_12918,N_9535,N_9234);
nor U12919 (N_12919,N_9137,N_9368);
nand U12920 (N_12920,N_9648,N_9788);
nand U12921 (N_12921,N_11704,N_9552);
nand U12922 (N_12922,N_10299,N_9957);
nand U12923 (N_12923,N_11794,N_9014);
xnor U12924 (N_12924,N_9876,N_10364);
nand U12925 (N_12925,N_9860,N_10011);
and U12926 (N_12926,N_9235,N_11846);
xnor U12927 (N_12927,N_9580,N_11470);
nor U12928 (N_12928,N_10135,N_10465);
xor U12929 (N_12929,N_10868,N_10120);
nor U12930 (N_12930,N_9594,N_9448);
or U12931 (N_12931,N_9370,N_9077);
nor U12932 (N_12932,N_10850,N_9899);
nor U12933 (N_12933,N_11129,N_10145);
or U12934 (N_12934,N_11768,N_9369);
nand U12935 (N_12935,N_11803,N_9318);
nand U12936 (N_12936,N_9221,N_10905);
nand U12937 (N_12937,N_9918,N_11753);
nand U12938 (N_12938,N_10409,N_9238);
xor U12939 (N_12939,N_10367,N_9970);
and U12940 (N_12940,N_9174,N_11166);
nor U12941 (N_12941,N_10024,N_9817);
nor U12942 (N_12942,N_11126,N_10353);
xnor U12943 (N_12943,N_10114,N_9301);
xnor U12944 (N_12944,N_10668,N_11712);
xor U12945 (N_12945,N_11994,N_9262);
nor U12946 (N_12946,N_11686,N_11818);
or U12947 (N_12947,N_11444,N_10839);
xnor U12948 (N_12948,N_9103,N_10821);
nand U12949 (N_12949,N_9736,N_9264);
nor U12950 (N_12950,N_10545,N_10207);
and U12951 (N_12951,N_11901,N_9818);
and U12952 (N_12952,N_10779,N_9279);
or U12953 (N_12953,N_11665,N_9794);
nor U12954 (N_12954,N_11968,N_10795);
nor U12955 (N_12955,N_10505,N_9446);
xnor U12956 (N_12956,N_9418,N_9061);
nand U12957 (N_12957,N_11435,N_11032);
and U12958 (N_12958,N_9716,N_9313);
or U12959 (N_12959,N_10688,N_11603);
nor U12960 (N_12960,N_10631,N_9826);
nand U12961 (N_12961,N_9189,N_11246);
and U12962 (N_12962,N_11178,N_11620);
nor U12963 (N_12963,N_11742,N_11764);
or U12964 (N_12964,N_11136,N_9514);
nor U12965 (N_12965,N_11991,N_9276);
and U12966 (N_12966,N_9574,N_11095);
and U12967 (N_12967,N_9432,N_10064);
or U12968 (N_12968,N_9154,N_10446);
nand U12969 (N_12969,N_9133,N_11543);
or U12970 (N_12970,N_11878,N_11691);
or U12971 (N_12971,N_11157,N_10125);
xnor U12972 (N_12972,N_9658,N_10805);
and U12973 (N_12973,N_10035,N_11828);
nand U12974 (N_12974,N_9405,N_9602);
xnor U12975 (N_12975,N_10678,N_9972);
nand U12976 (N_12976,N_11167,N_9084);
nor U12977 (N_12977,N_9184,N_11285);
nand U12978 (N_12978,N_10764,N_10334);
nand U12979 (N_12979,N_10712,N_10523);
xnor U12980 (N_12980,N_9756,N_11795);
and U12981 (N_12981,N_10286,N_11025);
or U12982 (N_12982,N_11228,N_10558);
nand U12983 (N_12983,N_10560,N_9411);
xor U12984 (N_12984,N_11821,N_9088);
xnor U12985 (N_12985,N_10354,N_9111);
nor U12986 (N_12986,N_9892,N_10672);
or U12987 (N_12987,N_11221,N_10209);
nor U12988 (N_12988,N_11003,N_9427);
xor U12989 (N_12989,N_10264,N_10849);
xnor U12990 (N_12990,N_10780,N_9608);
xnor U12991 (N_12991,N_10019,N_9735);
xor U12992 (N_12992,N_9509,N_11286);
nor U12993 (N_12993,N_11225,N_9650);
or U12994 (N_12994,N_9600,N_9905);
or U12995 (N_12995,N_10092,N_10080);
nand U12996 (N_12996,N_9692,N_11591);
nor U12997 (N_12997,N_10182,N_9142);
xnor U12998 (N_12998,N_11964,N_10319);
nor U12999 (N_12999,N_9802,N_11617);
nand U13000 (N_13000,N_10514,N_10587);
xnor U13001 (N_13001,N_11744,N_10496);
xor U13002 (N_13002,N_9978,N_11163);
nand U13003 (N_13003,N_11449,N_11146);
and U13004 (N_13004,N_11518,N_10098);
and U13005 (N_13005,N_10386,N_11816);
nor U13006 (N_13006,N_9241,N_9170);
and U13007 (N_13007,N_9486,N_10966);
nor U13008 (N_13008,N_10058,N_10298);
nand U13009 (N_13009,N_11815,N_11798);
xnor U13010 (N_13010,N_10854,N_9965);
nor U13011 (N_13011,N_11037,N_9625);
nor U13012 (N_13012,N_11774,N_10437);
nor U13013 (N_13013,N_11473,N_9773);
nor U13014 (N_13014,N_10722,N_11017);
or U13015 (N_13015,N_10277,N_11147);
nand U13016 (N_13016,N_9865,N_10435);
nand U13017 (N_13017,N_11343,N_11923);
xor U13018 (N_13018,N_9640,N_9177);
nor U13019 (N_13019,N_10793,N_10961);
or U13020 (N_13020,N_9498,N_11175);
xor U13021 (N_13021,N_10749,N_10358);
and U13022 (N_13022,N_11455,N_11200);
and U13023 (N_13023,N_11549,N_10962);
or U13024 (N_13024,N_10105,N_11539);
and U13025 (N_13025,N_10543,N_11585);
or U13026 (N_13026,N_11622,N_10773);
or U13027 (N_13027,N_10925,N_11372);
nor U13028 (N_13028,N_11478,N_10297);
and U13029 (N_13029,N_9036,N_10922);
nor U13030 (N_13030,N_10571,N_9982);
xnor U13031 (N_13031,N_9091,N_9290);
xor U13032 (N_13032,N_11208,N_11817);
xnor U13033 (N_13033,N_11492,N_11331);
xnor U13034 (N_13034,N_11084,N_10685);
or U13035 (N_13035,N_9270,N_11749);
or U13036 (N_13036,N_11667,N_11476);
xor U13037 (N_13037,N_10751,N_11845);
and U13038 (N_13038,N_9626,N_11040);
nand U13039 (N_13039,N_11750,N_10040);
nand U13040 (N_13040,N_9610,N_11206);
xor U13041 (N_13041,N_11169,N_9254);
xnor U13042 (N_13042,N_9072,N_10899);
nand U13043 (N_13043,N_10452,N_9768);
or U13044 (N_13044,N_10306,N_10378);
or U13045 (N_13045,N_10357,N_10508);
xor U13046 (N_13046,N_10110,N_11907);
nor U13047 (N_13047,N_11981,N_9897);
nor U13048 (N_13048,N_10392,N_9949);
nand U13049 (N_13049,N_9375,N_10502);
xnor U13050 (N_13050,N_11123,N_10771);
and U13051 (N_13051,N_9916,N_9096);
and U13052 (N_13052,N_11369,N_10513);
nor U13053 (N_13053,N_10396,N_11423);
and U13054 (N_13054,N_9153,N_11575);
and U13055 (N_13055,N_9906,N_11495);
xor U13056 (N_13056,N_11710,N_10522);
nand U13057 (N_13057,N_10911,N_10049);
nor U13058 (N_13058,N_10068,N_11446);
and U13059 (N_13059,N_9382,N_9992);
nand U13060 (N_13060,N_10046,N_10692);
nand U13061 (N_13061,N_9884,N_9412);
nand U13062 (N_13062,N_10346,N_9297);
and U13063 (N_13063,N_9348,N_11140);
nor U13064 (N_13064,N_10663,N_9502);
and U13065 (N_13065,N_9874,N_11916);
or U13066 (N_13066,N_9130,N_11241);
or U13067 (N_13067,N_11510,N_10293);
nor U13068 (N_13068,N_10992,N_11623);
and U13069 (N_13069,N_9351,N_11414);
xor U13070 (N_13070,N_10472,N_9354);
nor U13071 (N_13071,N_9139,N_9043);
nor U13072 (N_13072,N_11072,N_9745);
nor U13073 (N_13073,N_10582,N_11016);
and U13074 (N_13074,N_11969,N_10174);
and U13075 (N_13075,N_10249,N_11998);
nand U13076 (N_13076,N_9473,N_10835);
nor U13077 (N_13077,N_9101,N_9070);
xor U13078 (N_13078,N_11233,N_11628);
xor U13079 (N_13079,N_9400,N_9333);
xor U13080 (N_13080,N_9503,N_10963);
nor U13081 (N_13081,N_11263,N_10029);
nand U13082 (N_13082,N_9776,N_10356);
xnor U13083 (N_13083,N_9060,N_9251);
and U13084 (N_13084,N_11137,N_11909);
or U13085 (N_13085,N_11413,N_11705);
nand U13086 (N_13086,N_10172,N_11716);
or U13087 (N_13087,N_11868,N_9056);
xnor U13088 (N_13088,N_9712,N_9403);
xor U13089 (N_13089,N_11386,N_10991);
or U13090 (N_13090,N_11308,N_9196);
nor U13091 (N_13091,N_11740,N_11041);
nand U13092 (N_13092,N_10085,N_10642);
xnor U13093 (N_13093,N_9746,N_11958);
xor U13094 (N_13094,N_10814,N_9038);
nor U13095 (N_13095,N_10116,N_10828);
nand U13096 (N_13096,N_9475,N_10861);
or U13097 (N_13097,N_10164,N_11986);
nand U13098 (N_13098,N_10724,N_10160);
nand U13099 (N_13099,N_10527,N_9211);
or U13100 (N_13100,N_11912,N_9831);
and U13101 (N_13101,N_10315,N_9310);
xnor U13102 (N_13102,N_9398,N_11412);
or U13103 (N_13103,N_9435,N_10909);
or U13104 (N_13104,N_11099,N_9586);
nand U13105 (N_13105,N_10921,N_10062);
and U13106 (N_13106,N_11647,N_9097);
nand U13107 (N_13107,N_11800,N_9328);
nor U13108 (N_13108,N_11390,N_10817);
nor U13109 (N_13109,N_9296,N_11103);
and U13110 (N_13110,N_9155,N_11548);
nand U13111 (N_13111,N_10130,N_10456);
nand U13112 (N_13112,N_11942,N_10928);
nand U13113 (N_13113,N_9998,N_11924);
and U13114 (N_13114,N_11483,N_9515);
and U13115 (N_13115,N_11580,N_11106);
nand U13116 (N_13116,N_9963,N_9718);
or U13117 (N_13117,N_10248,N_9115);
nor U13118 (N_13118,N_9402,N_9522);
and U13119 (N_13119,N_11760,N_11762);
nand U13120 (N_13120,N_9144,N_10275);
or U13121 (N_13121,N_10281,N_9582);
or U13122 (N_13122,N_9025,N_9117);
nor U13123 (N_13123,N_9759,N_11957);
nor U13124 (N_13124,N_9349,N_9583);
nand U13125 (N_13125,N_11875,N_10149);
nor U13126 (N_13126,N_9340,N_11468);
nor U13127 (N_13127,N_9366,N_10944);
xor U13128 (N_13128,N_10783,N_9933);
nor U13129 (N_13129,N_11018,N_11791);
and U13130 (N_13130,N_9429,N_10482);
xnor U13131 (N_13131,N_11863,N_11259);
or U13132 (N_13132,N_9968,N_11578);
nand U13133 (N_13133,N_10022,N_10604);
or U13134 (N_13134,N_10316,N_9383);
xnor U13135 (N_13135,N_9937,N_11397);
and U13136 (N_13136,N_9734,N_10222);
nand U13137 (N_13137,N_10400,N_9114);
nand U13138 (N_13138,N_11899,N_9045);
xnor U13139 (N_13139,N_10945,N_10088);
or U13140 (N_13140,N_9770,N_9909);
or U13141 (N_13141,N_9325,N_10185);
nand U13142 (N_13142,N_11801,N_10661);
nand U13143 (N_13143,N_9119,N_10218);
and U13144 (N_13144,N_10912,N_11688);
or U13145 (N_13145,N_10190,N_10696);
and U13146 (N_13146,N_9846,N_9921);
xor U13147 (N_13147,N_10957,N_10253);
xor U13148 (N_13148,N_10971,N_11187);
xor U13149 (N_13149,N_10370,N_11793);
or U13150 (N_13150,N_9245,N_9445);
or U13151 (N_13151,N_11305,N_10981);
or U13152 (N_13152,N_11399,N_9118);
or U13153 (N_13153,N_10219,N_9757);
and U13154 (N_13154,N_9841,N_10769);
nor U13155 (N_13155,N_9416,N_11574);
xnor U13156 (N_13156,N_9593,N_10633);
xor U13157 (N_13157,N_9394,N_11695);
xnor U13158 (N_13158,N_9172,N_10179);
xnor U13159 (N_13159,N_10427,N_11362);
nor U13160 (N_13160,N_11229,N_10999);
nand U13161 (N_13161,N_11745,N_9979);
or U13162 (N_13162,N_11911,N_11896);
nor U13163 (N_13163,N_11133,N_9740);
nand U13164 (N_13164,N_10870,N_10159);
and U13165 (N_13165,N_10588,N_10484);
nand U13166 (N_13166,N_9885,N_11337);
and U13167 (N_13167,N_10655,N_11990);
nor U13168 (N_13168,N_9023,N_11522);
or U13169 (N_13169,N_10784,N_11057);
or U13170 (N_13170,N_9377,N_10526);
xnor U13171 (N_13171,N_9848,N_9146);
and U13172 (N_13172,N_9844,N_10459);
xnor U13173 (N_13173,N_11475,N_9378);
or U13174 (N_13174,N_11264,N_9050);
or U13175 (N_13175,N_10645,N_9480);
and U13176 (N_13176,N_9836,N_10054);
and U13177 (N_13177,N_9358,N_10273);
and U13178 (N_13178,N_9265,N_9666);
and U13179 (N_13179,N_9815,N_10485);
or U13180 (N_13180,N_9789,N_9180);
nand U13181 (N_13181,N_10347,N_11889);
and U13182 (N_13182,N_9873,N_9683);
nand U13183 (N_13183,N_10586,N_9946);
and U13184 (N_13184,N_11080,N_10169);
and U13185 (N_13185,N_11008,N_10593);
nand U13186 (N_13186,N_10680,N_9094);
and U13187 (N_13187,N_11404,N_11047);
and U13188 (N_13188,N_9000,N_9371);
nor U13189 (N_13189,N_11503,N_10694);
nand U13190 (N_13190,N_11908,N_10841);
nor U13191 (N_13191,N_9185,N_10124);
nor U13192 (N_13192,N_9869,N_9913);
nor U13193 (N_13193,N_9825,N_9492);
and U13194 (N_13194,N_9530,N_11511);
nand U13195 (N_13195,N_11933,N_11322);
xor U13196 (N_13196,N_11284,N_11732);
or U13197 (N_13197,N_10515,N_10430);
xnor U13198 (N_13198,N_11082,N_11261);
xnor U13199 (N_13199,N_10833,N_11640);
nand U13200 (N_13200,N_10477,N_9753);
xor U13201 (N_13201,N_11741,N_9647);
nor U13202 (N_13202,N_11482,N_10042);
nand U13203 (N_13203,N_11480,N_11723);
nand U13204 (N_13204,N_9141,N_9319);
or U13205 (N_13205,N_11779,N_10454);
nand U13206 (N_13206,N_9011,N_11880);
xnor U13207 (N_13207,N_11447,N_11422);
nor U13208 (N_13208,N_10183,N_10408);
or U13209 (N_13209,N_9321,N_11391);
or U13210 (N_13210,N_10895,N_11098);
nand U13211 (N_13211,N_9915,N_9408);
and U13212 (N_13212,N_10658,N_9819);
xnor U13213 (N_13213,N_10490,N_11955);
nor U13214 (N_13214,N_9966,N_11272);
nor U13215 (N_13215,N_9472,N_10638);
nand U13216 (N_13216,N_11009,N_10308);
or U13217 (N_13217,N_9764,N_11312);
or U13218 (N_13218,N_9329,N_11217);
nor U13219 (N_13219,N_9434,N_11364);
or U13220 (N_13220,N_10225,N_10274);
nand U13221 (N_13221,N_11097,N_9459);
xor U13222 (N_13222,N_9617,N_9450);
nand U13223 (N_13223,N_11214,N_9684);
nor U13224 (N_13224,N_10212,N_10272);
or U13225 (N_13225,N_11807,N_11043);
or U13226 (N_13226,N_10492,N_10853);
and U13227 (N_13227,N_9621,N_10432);
or U13228 (N_13228,N_10951,N_9612);
xnor U13229 (N_13229,N_10368,N_11941);
xor U13230 (N_13230,N_9501,N_9636);
nand U13231 (N_13231,N_11254,N_9001);
nor U13232 (N_13232,N_11138,N_11109);
nand U13233 (N_13233,N_9925,N_9386);
or U13234 (N_13234,N_10882,N_9163);
and U13235 (N_13235,N_9930,N_11684);
and U13236 (N_13236,N_11841,N_10852);
and U13237 (N_13237,N_10194,N_10240);
nand U13238 (N_13238,N_11398,N_10399);
nor U13239 (N_13239,N_10715,N_11730);
or U13240 (N_13240,N_9152,N_11508);
or U13241 (N_13241,N_9273,N_9148);
nand U13242 (N_13242,N_9210,N_10993);
and U13243 (N_13243,N_10377,N_9634);
xor U13244 (N_13244,N_11332,N_10665);
nor U13245 (N_13245,N_9456,N_10471);
or U13246 (N_13246,N_9560,N_10072);
nor U13247 (N_13247,N_10387,N_10798);
nand U13248 (N_13248,N_11677,N_11006);
xor U13249 (N_13249,N_9267,N_11852);
nand U13250 (N_13250,N_10235,N_10723);
nor U13251 (N_13251,N_11910,N_11144);
nor U13252 (N_13252,N_10401,N_11148);
and U13253 (N_13253,N_9908,N_9903);
xor U13254 (N_13254,N_9102,N_10375);
or U13255 (N_13255,N_11066,N_10250);
or U13256 (N_13256,N_11360,N_9006);
xnor U13257 (N_13257,N_9834,N_11474);
nor U13258 (N_13258,N_10507,N_9156);
or U13259 (N_13259,N_11931,N_9391);
or U13260 (N_13260,N_9007,N_10263);
or U13261 (N_13261,N_10689,N_11083);
and U13262 (N_13262,N_9120,N_11757);
xnor U13263 (N_13263,N_10107,N_9526);
xnor U13264 (N_13264,N_9808,N_10646);
or U13265 (N_13265,N_10913,N_9202);
xor U13266 (N_13266,N_10366,N_9732);
and U13267 (N_13267,N_9243,N_11341);
nand U13268 (N_13268,N_9554,N_10669);
xnor U13269 (N_13269,N_11400,N_9657);
xnor U13270 (N_13270,N_10047,N_10280);
and U13271 (N_13271,N_9839,N_10339);
nand U13272 (N_13272,N_9345,N_11989);
or U13273 (N_13273,N_9828,N_9200);
nand U13274 (N_13274,N_10039,N_11465);
and U13275 (N_13275,N_9571,N_9538);
nor U13276 (N_13276,N_9324,N_9564);
xor U13277 (N_13277,N_9950,N_10388);
nand U13278 (N_13278,N_9751,N_10717);
nand U13279 (N_13279,N_9205,N_10803);
xnor U13280 (N_13280,N_11616,N_9441);
nor U13281 (N_13281,N_9244,N_9362);
or U13282 (N_13282,N_11861,N_10012);
nand U13283 (N_13283,N_9207,N_11488);
xor U13284 (N_13284,N_11002,N_11687);
and U13285 (N_13285,N_10982,N_9584);
or U13286 (N_13286,N_11439,N_10422);
xnor U13287 (N_13287,N_11752,N_9108);
nand U13288 (N_13288,N_9591,N_10716);
and U13289 (N_13289,N_10767,N_11538);
nand U13290 (N_13290,N_9893,N_10630);
nand U13291 (N_13291,N_9017,N_11116);
or U13292 (N_13292,N_10553,N_10733);
xnor U13293 (N_13293,N_11346,N_9081);
nand U13294 (N_13294,N_10550,N_10622);
and U13295 (N_13295,N_9054,N_11068);
nand U13296 (N_13296,N_10026,N_10790);
and U13297 (N_13297,N_11085,N_11373);
xnor U13298 (N_13298,N_9852,N_11759);
and U13299 (N_13299,N_9785,N_10206);
nor U13300 (N_13300,N_11544,N_11289);
and U13301 (N_13301,N_11198,N_9812);
nand U13302 (N_13302,N_10748,N_10864);
nand U13303 (N_13303,N_9112,N_10755);
xnor U13304 (N_13304,N_9213,N_11053);
or U13305 (N_13305,N_10383,N_10048);
xnor U13306 (N_13306,N_9331,N_10761);
xor U13307 (N_13307,N_10457,N_11202);
xnor U13308 (N_13308,N_10106,N_10616);
or U13309 (N_13309,N_10090,N_10796);
nand U13310 (N_13310,N_11036,N_11420);
xnor U13311 (N_13311,N_11236,N_10442);
nor U13312 (N_13312,N_9859,N_10564);
xor U13313 (N_13313,N_9135,N_9326);
or U13314 (N_13314,N_9713,N_11631);
nor U13315 (N_13315,N_10201,N_10517);
and U13316 (N_13316,N_10896,N_9791);
xnor U13317 (N_13317,N_10516,N_11282);
and U13318 (N_13318,N_9989,N_10504);
nand U13319 (N_13319,N_11393,N_11213);
or U13320 (N_13320,N_11090,N_10243);
xor U13321 (N_13321,N_10025,N_11581);
or U13322 (N_13322,N_9795,N_10268);
or U13323 (N_13323,N_10613,N_10154);
nand U13324 (N_13324,N_10743,N_9015);
xnor U13325 (N_13325,N_10705,N_9367);
nor U13326 (N_13326,N_11601,N_9677);
nor U13327 (N_13327,N_11299,N_11112);
nor U13328 (N_13328,N_9442,N_11383);
or U13329 (N_13329,N_9694,N_10741);
nor U13330 (N_13330,N_11717,N_11155);
nor U13331 (N_13331,N_9508,N_11224);
xor U13332 (N_13332,N_10385,N_11827);
nand U13333 (N_13333,N_9026,N_11436);
nor U13334 (N_13334,N_10181,N_10009);
and U13335 (N_13335,N_9708,N_10241);
and U13336 (N_13336,N_9413,N_11615);
and U13337 (N_13337,N_10076,N_9338);
and U13338 (N_13338,N_10778,N_9547);
and U13339 (N_13339,N_11275,N_10095);
xnor U13340 (N_13340,N_11769,N_11499);
nand U13341 (N_13341,N_11357,N_10065);
xnor U13342 (N_13342,N_11790,N_9661);
nor U13343 (N_13343,N_11355,N_11481);
and U13344 (N_13344,N_9798,N_9431);
nand U13345 (N_13345,N_9569,N_11122);
nor U13346 (N_13346,N_9306,N_11477);
nor U13347 (N_13347,N_10664,N_10450);
nand U13348 (N_13348,N_10950,N_9843);
xor U13349 (N_13349,N_11319,N_9872);
or U13350 (N_13350,N_9491,N_11625);
xor U13351 (N_13351,N_9430,N_9124);
xor U13352 (N_13352,N_9741,N_10016);
xnor U13353 (N_13353,N_11251,N_11504);
or U13354 (N_13354,N_9388,N_11179);
and U13355 (N_13355,N_11563,N_10355);
nand U13356 (N_13356,N_10679,N_11015);
nand U13357 (N_13357,N_10075,N_9517);
xnor U13358 (N_13358,N_9642,N_10322);
nor U13359 (N_13359,N_11927,N_11805);
nand U13360 (N_13360,N_9880,N_9644);
nand U13361 (N_13361,N_10175,N_9975);
nand U13362 (N_13362,N_9742,N_11588);
and U13363 (N_13363,N_9668,N_10051);
nand U13364 (N_13364,N_9312,N_9246);
nor U13365 (N_13365,N_11835,N_9889);
nand U13366 (N_13366,N_10447,N_9572);
and U13367 (N_13367,N_9457,N_10284);
xnor U13368 (N_13368,N_11385,N_10003);
and U13369 (N_13369,N_10893,N_10416);
xnor U13370 (N_13370,N_11049,N_11781);
and U13371 (N_13371,N_11000,N_10675);
and U13372 (N_13372,N_11668,N_11596);
xor U13373 (N_13373,N_11627,N_11786);
nor U13374 (N_13374,N_9672,N_9790);
nand U13375 (N_13375,N_10546,N_10953);
and U13376 (N_13376,N_11589,N_11056);
and U13377 (N_13377,N_10781,N_10458);
and U13378 (N_13378,N_9524,N_11703);
nand U13379 (N_13379,N_10568,N_11472);
nand U13380 (N_13380,N_10070,N_11658);
or U13381 (N_13381,N_9875,N_10826);
nor U13382 (N_13382,N_9161,N_11437);
xnor U13383 (N_13383,N_10930,N_11883);
or U13384 (N_13384,N_11434,N_10832);
nor U13385 (N_13385,N_9733,N_10498);
nand U13386 (N_13386,N_11825,N_10524);
nand U13387 (N_13387,N_11172,N_10074);
xnor U13388 (N_13388,N_9723,N_11936);
xnor U13389 (N_13389,N_10310,N_11127);
and U13390 (N_13390,N_10200,N_11569);
nor U13391 (N_13391,N_11512,N_9029);
or U13392 (N_13392,N_11496,N_11207);
and U13393 (N_13393,N_9660,N_10015);
or U13394 (N_13394,N_11300,N_10801);
nand U13395 (N_13395,N_11121,N_11031);
nand U13396 (N_13396,N_11196,N_9085);
nor U13397 (N_13397,N_11231,N_10487);
and U13398 (N_13398,N_10220,N_11415);
xnor U13399 (N_13399,N_10336,N_10034);
nor U13400 (N_13400,N_10410,N_11528);
nand U13401 (N_13401,N_10137,N_9390);
xnor U13402 (N_13402,N_11440,N_11265);
and U13403 (N_13403,N_10954,N_10132);
nand U13404 (N_13404,N_9956,N_10141);
xor U13405 (N_13405,N_11501,N_9935);
or U13406 (N_13406,N_11777,N_10059);
nand U13407 (N_13407,N_10312,N_11784);
nand U13408 (N_13408,N_10703,N_10802);
nand U13409 (N_13409,N_10119,N_10562);
and U13410 (N_13410,N_10203,N_10775);
or U13411 (N_13411,N_9619,N_11458);
nand U13412 (N_13412,N_9237,N_9793);
nand U13413 (N_13413,N_10830,N_9896);
or U13414 (N_13414,N_9888,N_11086);
nand U13415 (N_13415,N_9266,N_11650);
xnor U13416 (N_13416,N_9123,N_11281);
nor U13417 (N_13417,N_11402,N_11240);
nand U13418 (N_13418,N_11471,N_9044);
and U13419 (N_13419,N_9471,N_9544);
nor U13420 (N_13420,N_10178,N_11672);
nand U13421 (N_13421,N_11361,N_9777);
or U13422 (N_13422,N_10036,N_10728);
nand U13423 (N_13423,N_11613,N_11754);
or U13424 (N_13424,N_10887,N_11334);
or U13425 (N_13425,N_10254,N_11993);
nand U13426 (N_13426,N_9401,N_10118);
nand U13427 (N_13427,N_10644,N_11039);
nor U13428 (N_13428,N_10908,N_9136);
nand U13429 (N_13429,N_11887,N_9911);
nor U13430 (N_13430,N_10196,N_9861);
and U13431 (N_13431,N_10139,N_10635);
nand U13432 (N_13432,N_10351,N_10627);
or U13433 (N_13433,N_10289,N_9673);
nor U13434 (N_13434,N_11500,N_10583);
or U13435 (N_13435,N_9652,N_9165);
xnor U13436 (N_13436,N_11430,N_9468);
nor U13437 (N_13437,N_10624,N_11132);
nand U13438 (N_13438,N_10311,N_9149);
xor U13439 (N_13439,N_11976,N_9031);
nand U13440 (N_13440,N_9373,N_9062);
xor U13441 (N_13441,N_11316,N_10186);
and U13442 (N_13442,N_10214,N_11335);
and U13443 (N_13443,N_10146,N_10060);
or U13444 (N_13444,N_9214,N_10082);
nand U13445 (N_13445,N_10260,N_9674);
and U13446 (N_13446,N_10590,N_9496);
and U13447 (N_13447,N_9807,N_9160);
nand U13448 (N_13448,N_10707,N_10434);
nand U13449 (N_13449,N_9162,N_9731);
xor U13450 (N_13450,N_9147,N_9479);
xnor U13451 (N_13451,N_11234,N_11452);
nand U13452 (N_13452,N_11611,N_11564);
xnor U13453 (N_13453,N_10885,N_10004);
and U13454 (N_13454,N_11935,N_10934);
xor U13455 (N_13455,N_10931,N_11963);
or U13456 (N_13456,N_9796,N_11320);
and U13457 (N_13457,N_9699,N_9851);
nor U13458 (N_13458,N_11514,N_11940);
and U13459 (N_13459,N_11274,N_9337);
or U13460 (N_13460,N_9623,N_10600);
xor U13461 (N_13461,N_10632,N_9531);
xnor U13462 (N_13462,N_11515,N_10557);
or U13463 (N_13463,N_10233,N_10069);
or U13464 (N_13464,N_9606,N_9485);
nand U13465 (N_13465,N_9820,N_11526);
or U13466 (N_13466,N_9748,N_9651);
nand U13467 (N_13467,N_10949,N_9212);
or U13468 (N_13468,N_11946,N_9002);
or U13469 (N_13469,N_9504,N_9543);
and U13470 (N_13470,N_11010,N_9771);
and U13471 (N_13471,N_11610,N_11170);
and U13472 (N_13472,N_11586,N_10652);
nor U13473 (N_13473,N_10732,N_10719);
nor U13474 (N_13474,N_11042,N_9994);
xor U13475 (N_13475,N_10544,N_11038);
nand U13476 (N_13476,N_10267,N_11583);
xor U13477 (N_13477,N_10162,N_11484);
and U13478 (N_13478,N_9540,N_11280);
and U13479 (N_13479,N_10729,N_9715);
nand U13480 (N_13480,N_10189,N_11463);
or U13481 (N_13481,N_10697,N_11836);
xor U13482 (N_13482,N_9188,N_10165);
and U13483 (N_13483,N_10618,N_9271);
xor U13484 (N_13484,N_9278,N_10929);
nand U13485 (N_13485,N_10579,N_9075);
or U13486 (N_13486,N_9065,N_11773);
or U13487 (N_13487,N_11209,N_10987);
nor U13488 (N_13488,N_10005,N_11054);
nand U13489 (N_13489,N_9078,N_9618);
nand U13490 (N_13490,N_11469,N_11464);
nand U13491 (N_13491,N_11028,N_10232);
or U13492 (N_13492,N_11866,N_11353);
or U13493 (N_13493,N_9864,N_10520);
nor U13494 (N_13494,N_9548,N_10794);
nor U13495 (N_13495,N_11867,N_9671);
or U13496 (N_13496,N_10153,N_11531);
xnor U13497 (N_13497,N_10192,N_10510);
and U13498 (N_13498,N_11220,N_11590);
nand U13499 (N_13499,N_9604,N_10628);
xnor U13500 (N_13500,N_11936,N_9562);
xor U13501 (N_13501,N_10706,N_10310);
and U13502 (N_13502,N_9943,N_11162);
and U13503 (N_13503,N_11405,N_11579);
nand U13504 (N_13504,N_10057,N_11974);
or U13505 (N_13505,N_9770,N_9472);
nand U13506 (N_13506,N_9636,N_9022);
nand U13507 (N_13507,N_11538,N_9425);
or U13508 (N_13508,N_11850,N_9737);
and U13509 (N_13509,N_11667,N_9151);
or U13510 (N_13510,N_9409,N_9310);
nand U13511 (N_13511,N_9194,N_11355);
xnor U13512 (N_13512,N_10235,N_11682);
nor U13513 (N_13513,N_11088,N_11859);
and U13514 (N_13514,N_9885,N_10073);
and U13515 (N_13515,N_10492,N_11347);
xor U13516 (N_13516,N_9705,N_9301);
xor U13517 (N_13517,N_11206,N_10279);
nand U13518 (N_13518,N_9615,N_9254);
and U13519 (N_13519,N_11715,N_11341);
and U13520 (N_13520,N_9426,N_9128);
xnor U13521 (N_13521,N_9921,N_10738);
nor U13522 (N_13522,N_11642,N_11688);
or U13523 (N_13523,N_10499,N_11192);
xnor U13524 (N_13524,N_11918,N_9264);
xor U13525 (N_13525,N_10087,N_10195);
nand U13526 (N_13526,N_11037,N_10754);
and U13527 (N_13527,N_11314,N_9489);
or U13528 (N_13528,N_11942,N_11255);
xor U13529 (N_13529,N_11434,N_10529);
nor U13530 (N_13530,N_11970,N_11170);
or U13531 (N_13531,N_10653,N_11165);
nand U13532 (N_13532,N_10109,N_10242);
and U13533 (N_13533,N_11679,N_10427);
nand U13534 (N_13534,N_11288,N_10428);
xor U13535 (N_13535,N_11376,N_11878);
xnor U13536 (N_13536,N_10440,N_9981);
nor U13537 (N_13537,N_11204,N_9029);
or U13538 (N_13538,N_9762,N_9489);
and U13539 (N_13539,N_10729,N_9888);
and U13540 (N_13540,N_11279,N_11382);
and U13541 (N_13541,N_10688,N_9534);
and U13542 (N_13542,N_10504,N_10406);
xnor U13543 (N_13543,N_9234,N_9749);
nor U13544 (N_13544,N_10378,N_9766);
and U13545 (N_13545,N_11210,N_9429);
nor U13546 (N_13546,N_10160,N_9340);
or U13547 (N_13547,N_9547,N_11131);
nand U13548 (N_13548,N_9978,N_11157);
nand U13549 (N_13549,N_11715,N_11841);
and U13550 (N_13550,N_10717,N_9776);
nand U13551 (N_13551,N_9650,N_11072);
or U13552 (N_13552,N_11576,N_11273);
nand U13553 (N_13553,N_9885,N_11672);
xor U13554 (N_13554,N_9862,N_9322);
or U13555 (N_13555,N_11232,N_11358);
nor U13556 (N_13556,N_11387,N_10715);
or U13557 (N_13557,N_9115,N_9650);
or U13558 (N_13558,N_9321,N_9730);
nor U13559 (N_13559,N_11610,N_11151);
nor U13560 (N_13560,N_11254,N_10085);
nand U13561 (N_13561,N_9191,N_11104);
and U13562 (N_13562,N_10050,N_9550);
nor U13563 (N_13563,N_9878,N_11326);
nor U13564 (N_13564,N_9033,N_11583);
nand U13565 (N_13565,N_10671,N_11971);
or U13566 (N_13566,N_9027,N_11389);
nor U13567 (N_13567,N_11754,N_11755);
nor U13568 (N_13568,N_9451,N_10415);
nor U13569 (N_13569,N_10884,N_11036);
nand U13570 (N_13570,N_11852,N_10788);
nor U13571 (N_13571,N_11136,N_11583);
or U13572 (N_13572,N_9615,N_9896);
nand U13573 (N_13573,N_9483,N_11791);
nor U13574 (N_13574,N_9078,N_9123);
and U13575 (N_13575,N_10564,N_9623);
and U13576 (N_13576,N_10201,N_11422);
or U13577 (N_13577,N_9370,N_10030);
nor U13578 (N_13578,N_11093,N_11170);
nand U13579 (N_13579,N_10567,N_11776);
xnor U13580 (N_13580,N_11468,N_9991);
nor U13581 (N_13581,N_9929,N_11303);
xor U13582 (N_13582,N_9329,N_9752);
and U13583 (N_13583,N_10664,N_9419);
and U13584 (N_13584,N_9903,N_11322);
nor U13585 (N_13585,N_9444,N_9730);
nand U13586 (N_13586,N_10415,N_9940);
or U13587 (N_13587,N_10358,N_11423);
or U13588 (N_13588,N_10047,N_10237);
xor U13589 (N_13589,N_9105,N_10777);
and U13590 (N_13590,N_10554,N_9649);
and U13591 (N_13591,N_11069,N_11750);
xor U13592 (N_13592,N_10264,N_9515);
and U13593 (N_13593,N_9504,N_11347);
or U13594 (N_13594,N_10683,N_10489);
xor U13595 (N_13595,N_10674,N_10969);
and U13596 (N_13596,N_9154,N_11839);
nand U13597 (N_13597,N_11141,N_11367);
nand U13598 (N_13598,N_11561,N_11150);
xor U13599 (N_13599,N_11533,N_11308);
xnor U13600 (N_13600,N_11869,N_10908);
nand U13601 (N_13601,N_11196,N_9473);
nor U13602 (N_13602,N_10886,N_11523);
or U13603 (N_13603,N_10419,N_11462);
and U13604 (N_13604,N_9348,N_11917);
and U13605 (N_13605,N_11013,N_9442);
and U13606 (N_13606,N_11477,N_10847);
or U13607 (N_13607,N_11311,N_9303);
nand U13608 (N_13608,N_11098,N_10085);
nand U13609 (N_13609,N_11122,N_10733);
and U13610 (N_13610,N_10427,N_10638);
nor U13611 (N_13611,N_10402,N_10216);
nor U13612 (N_13612,N_9739,N_9457);
or U13613 (N_13613,N_10451,N_9480);
or U13614 (N_13614,N_9439,N_11755);
nand U13615 (N_13615,N_9717,N_10302);
or U13616 (N_13616,N_11212,N_10961);
xor U13617 (N_13617,N_10522,N_9302);
xnor U13618 (N_13618,N_10905,N_9110);
or U13619 (N_13619,N_10399,N_9094);
and U13620 (N_13620,N_11001,N_11135);
xnor U13621 (N_13621,N_10434,N_9262);
xnor U13622 (N_13622,N_11525,N_11390);
nor U13623 (N_13623,N_11748,N_11485);
nand U13624 (N_13624,N_9507,N_11989);
and U13625 (N_13625,N_11967,N_9026);
xnor U13626 (N_13626,N_9915,N_10180);
or U13627 (N_13627,N_10087,N_10166);
and U13628 (N_13628,N_10343,N_10459);
or U13629 (N_13629,N_9023,N_10893);
and U13630 (N_13630,N_10679,N_9177);
nand U13631 (N_13631,N_11919,N_11314);
nand U13632 (N_13632,N_10500,N_11496);
nor U13633 (N_13633,N_9908,N_9623);
xnor U13634 (N_13634,N_9554,N_10542);
xor U13635 (N_13635,N_9067,N_10112);
nand U13636 (N_13636,N_9610,N_11011);
nand U13637 (N_13637,N_9074,N_9283);
or U13638 (N_13638,N_10363,N_10823);
and U13639 (N_13639,N_9811,N_9262);
nand U13640 (N_13640,N_10392,N_9644);
and U13641 (N_13641,N_11362,N_11898);
xor U13642 (N_13642,N_10147,N_11889);
nand U13643 (N_13643,N_10940,N_10515);
nor U13644 (N_13644,N_10562,N_11574);
nor U13645 (N_13645,N_9273,N_11409);
xor U13646 (N_13646,N_10572,N_10671);
or U13647 (N_13647,N_9899,N_11739);
nand U13648 (N_13648,N_11240,N_11617);
or U13649 (N_13649,N_10616,N_9433);
xnor U13650 (N_13650,N_9563,N_9907);
nand U13651 (N_13651,N_9238,N_11872);
nor U13652 (N_13652,N_10391,N_10715);
and U13653 (N_13653,N_11150,N_11433);
and U13654 (N_13654,N_10827,N_9446);
and U13655 (N_13655,N_9660,N_10284);
and U13656 (N_13656,N_9127,N_10565);
and U13657 (N_13657,N_11820,N_10153);
or U13658 (N_13658,N_10099,N_9002);
and U13659 (N_13659,N_9642,N_11228);
xnor U13660 (N_13660,N_9291,N_11871);
xor U13661 (N_13661,N_9130,N_9014);
or U13662 (N_13662,N_9121,N_10738);
nor U13663 (N_13663,N_10838,N_10002);
xor U13664 (N_13664,N_9671,N_9473);
or U13665 (N_13665,N_11445,N_9172);
and U13666 (N_13666,N_9636,N_10029);
xor U13667 (N_13667,N_9213,N_9831);
and U13668 (N_13668,N_11050,N_11544);
xor U13669 (N_13669,N_10968,N_10280);
and U13670 (N_13670,N_10720,N_11975);
and U13671 (N_13671,N_11637,N_10462);
nand U13672 (N_13672,N_10092,N_9302);
xor U13673 (N_13673,N_9715,N_10802);
and U13674 (N_13674,N_11686,N_11768);
nor U13675 (N_13675,N_10581,N_11567);
xnor U13676 (N_13676,N_10734,N_9607);
nor U13677 (N_13677,N_10429,N_9972);
nor U13678 (N_13678,N_11884,N_9626);
xnor U13679 (N_13679,N_11383,N_10077);
xor U13680 (N_13680,N_11315,N_10557);
or U13681 (N_13681,N_10257,N_9054);
nor U13682 (N_13682,N_11858,N_10884);
nor U13683 (N_13683,N_11237,N_10793);
nor U13684 (N_13684,N_11440,N_9354);
nand U13685 (N_13685,N_11735,N_10425);
nand U13686 (N_13686,N_11308,N_9068);
nor U13687 (N_13687,N_10625,N_9478);
and U13688 (N_13688,N_9033,N_10662);
and U13689 (N_13689,N_10397,N_9463);
xor U13690 (N_13690,N_10072,N_9097);
nand U13691 (N_13691,N_10552,N_9209);
nand U13692 (N_13692,N_11499,N_9169);
nand U13693 (N_13693,N_10585,N_11096);
xor U13694 (N_13694,N_10317,N_10779);
xor U13695 (N_13695,N_11299,N_10436);
nand U13696 (N_13696,N_10545,N_11819);
nor U13697 (N_13697,N_11179,N_9310);
nor U13698 (N_13698,N_11711,N_11604);
nor U13699 (N_13699,N_11784,N_9599);
nor U13700 (N_13700,N_9754,N_10502);
or U13701 (N_13701,N_11396,N_10604);
and U13702 (N_13702,N_10945,N_11094);
nand U13703 (N_13703,N_10227,N_10719);
xor U13704 (N_13704,N_9589,N_9806);
and U13705 (N_13705,N_10096,N_11759);
or U13706 (N_13706,N_9848,N_11244);
and U13707 (N_13707,N_10387,N_11072);
xor U13708 (N_13708,N_11468,N_11781);
or U13709 (N_13709,N_9682,N_9050);
nand U13710 (N_13710,N_10649,N_10084);
or U13711 (N_13711,N_10773,N_11662);
xor U13712 (N_13712,N_11048,N_11384);
or U13713 (N_13713,N_9240,N_11516);
or U13714 (N_13714,N_10554,N_11358);
xnor U13715 (N_13715,N_10078,N_11221);
and U13716 (N_13716,N_9190,N_11684);
nand U13717 (N_13717,N_11782,N_9998);
or U13718 (N_13718,N_11980,N_9637);
or U13719 (N_13719,N_10766,N_11246);
xor U13720 (N_13720,N_10371,N_10970);
nor U13721 (N_13721,N_10239,N_10074);
and U13722 (N_13722,N_10476,N_9527);
nor U13723 (N_13723,N_9536,N_10477);
nor U13724 (N_13724,N_9491,N_10015);
nand U13725 (N_13725,N_10917,N_9446);
xor U13726 (N_13726,N_11763,N_9393);
nand U13727 (N_13727,N_11113,N_10143);
and U13728 (N_13728,N_9668,N_9225);
nand U13729 (N_13729,N_9897,N_11554);
and U13730 (N_13730,N_10818,N_9632);
nand U13731 (N_13731,N_10456,N_9230);
nor U13732 (N_13732,N_11175,N_9374);
nor U13733 (N_13733,N_10410,N_9036);
xnor U13734 (N_13734,N_11419,N_10380);
and U13735 (N_13735,N_10130,N_10303);
nand U13736 (N_13736,N_10236,N_10337);
nor U13737 (N_13737,N_9952,N_10705);
or U13738 (N_13738,N_11135,N_10180);
or U13739 (N_13739,N_10301,N_10471);
xnor U13740 (N_13740,N_9588,N_9869);
and U13741 (N_13741,N_10639,N_9337);
and U13742 (N_13742,N_9111,N_11537);
or U13743 (N_13743,N_9489,N_10696);
nor U13744 (N_13744,N_11841,N_11861);
nor U13745 (N_13745,N_11473,N_9881);
nor U13746 (N_13746,N_9919,N_10509);
or U13747 (N_13747,N_10156,N_9724);
and U13748 (N_13748,N_9491,N_9308);
and U13749 (N_13749,N_10073,N_9878);
and U13750 (N_13750,N_11379,N_11242);
xnor U13751 (N_13751,N_10980,N_9367);
and U13752 (N_13752,N_9270,N_9175);
or U13753 (N_13753,N_11342,N_11116);
nor U13754 (N_13754,N_10593,N_9177);
and U13755 (N_13755,N_10444,N_9539);
and U13756 (N_13756,N_10807,N_9789);
xnor U13757 (N_13757,N_9358,N_9491);
nand U13758 (N_13758,N_9499,N_10599);
or U13759 (N_13759,N_11766,N_9016);
xor U13760 (N_13760,N_9318,N_9218);
and U13761 (N_13761,N_11933,N_11294);
and U13762 (N_13762,N_10953,N_9645);
nor U13763 (N_13763,N_9238,N_11689);
and U13764 (N_13764,N_10049,N_9559);
nand U13765 (N_13765,N_10136,N_10538);
or U13766 (N_13766,N_9710,N_9918);
xor U13767 (N_13767,N_10585,N_9529);
nand U13768 (N_13768,N_10371,N_11373);
nor U13769 (N_13769,N_9867,N_11954);
or U13770 (N_13770,N_9842,N_10786);
or U13771 (N_13771,N_9978,N_9873);
and U13772 (N_13772,N_11661,N_9857);
nor U13773 (N_13773,N_11472,N_11947);
or U13774 (N_13774,N_11423,N_10111);
nor U13775 (N_13775,N_11338,N_9797);
and U13776 (N_13776,N_11475,N_9179);
nor U13777 (N_13777,N_10671,N_10195);
nor U13778 (N_13778,N_11554,N_10772);
and U13779 (N_13779,N_11877,N_10036);
and U13780 (N_13780,N_11422,N_10858);
xor U13781 (N_13781,N_10000,N_11838);
or U13782 (N_13782,N_10363,N_9928);
or U13783 (N_13783,N_11190,N_11454);
nand U13784 (N_13784,N_10430,N_11879);
nand U13785 (N_13785,N_11901,N_11350);
and U13786 (N_13786,N_10554,N_11256);
and U13787 (N_13787,N_11205,N_9035);
xor U13788 (N_13788,N_9503,N_11449);
and U13789 (N_13789,N_9560,N_11759);
nand U13790 (N_13790,N_10646,N_11133);
xnor U13791 (N_13791,N_11080,N_11769);
nand U13792 (N_13792,N_9700,N_10562);
xnor U13793 (N_13793,N_11614,N_10444);
nand U13794 (N_13794,N_9154,N_9229);
or U13795 (N_13795,N_9464,N_11240);
nand U13796 (N_13796,N_10106,N_9422);
nand U13797 (N_13797,N_11034,N_11230);
and U13798 (N_13798,N_11272,N_11620);
nor U13799 (N_13799,N_11097,N_11654);
nand U13800 (N_13800,N_11768,N_9344);
nor U13801 (N_13801,N_10678,N_11839);
xor U13802 (N_13802,N_11612,N_11348);
and U13803 (N_13803,N_9034,N_9087);
nand U13804 (N_13804,N_11508,N_10428);
xnor U13805 (N_13805,N_10969,N_9143);
and U13806 (N_13806,N_10836,N_9998);
or U13807 (N_13807,N_10556,N_11860);
nand U13808 (N_13808,N_11852,N_10124);
nand U13809 (N_13809,N_10367,N_9252);
and U13810 (N_13810,N_9721,N_10617);
and U13811 (N_13811,N_9124,N_9151);
or U13812 (N_13812,N_10591,N_10977);
and U13813 (N_13813,N_10177,N_10033);
nor U13814 (N_13814,N_9843,N_11224);
nor U13815 (N_13815,N_11262,N_11686);
xnor U13816 (N_13816,N_11548,N_11368);
nand U13817 (N_13817,N_9829,N_11944);
nor U13818 (N_13818,N_10915,N_10480);
nand U13819 (N_13819,N_9383,N_9119);
nor U13820 (N_13820,N_10664,N_10123);
xnor U13821 (N_13821,N_9291,N_9544);
nand U13822 (N_13822,N_9795,N_9178);
or U13823 (N_13823,N_10876,N_9003);
or U13824 (N_13824,N_9770,N_11780);
and U13825 (N_13825,N_10872,N_9360);
nand U13826 (N_13826,N_9111,N_10087);
nand U13827 (N_13827,N_11525,N_9090);
xnor U13828 (N_13828,N_10873,N_10263);
or U13829 (N_13829,N_11145,N_9622);
xor U13830 (N_13830,N_10625,N_10655);
or U13831 (N_13831,N_9311,N_11994);
and U13832 (N_13832,N_10233,N_10144);
nand U13833 (N_13833,N_10196,N_10809);
or U13834 (N_13834,N_9491,N_10355);
nor U13835 (N_13835,N_11890,N_10231);
nand U13836 (N_13836,N_10402,N_10238);
or U13837 (N_13837,N_9852,N_11542);
nor U13838 (N_13838,N_11233,N_9077);
xnor U13839 (N_13839,N_10099,N_10444);
nand U13840 (N_13840,N_10367,N_11044);
nor U13841 (N_13841,N_11049,N_10665);
nor U13842 (N_13842,N_9913,N_10374);
xor U13843 (N_13843,N_10326,N_9521);
or U13844 (N_13844,N_9032,N_9567);
nor U13845 (N_13845,N_9191,N_10972);
and U13846 (N_13846,N_11280,N_10081);
xnor U13847 (N_13847,N_11857,N_10337);
xor U13848 (N_13848,N_10217,N_10611);
nor U13849 (N_13849,N_10928,N_9284);
xnor U13850 (N_13850,N_11603,N_9186);
xor U13851 (N_13851,N_9423,N_9501);
xor U13852 (N_13852,N_10203,N_11295);
nand U13853 (N_13853,N_9000,N_9928);
xnor U13854 (N_13854,N_10130,N_10851);
nand U13855 (N_13855,N_9424,N_9796);
or U13856 (N_13856,N_10442,N_11770);
nor U13857 (N_13857,N_11491,N_9835);
nor U13858 (N_13858,N_9014,N_11937);
nand U13859 (N_13859,N_11293,N_11123);
nor U13860 (N_13860,N_11975,N_11705);
xor U13861 (N_13861,N_10367,N_9797);
xor U13862 (N_13862,N_11600,N_10440);
xnor U13863 (N_13863,N_11622,N_9861);
nor U13864 (N_13864,N_10907,N_10444);
and U13865 (N_13865,N_11923,N_11251);
or U13866 (N_13866,N_11202,N_11117);
nor U13867 (N_13867,N_10858,N_10371);
and U13868 (N_13868,N_9714,N_10865);
or U13869 (N_13869,N_11823,N_11004);
xnor U13870 (N_13870,N_9177,N_9102);
xnor U13871 (N_13871,N_9808,N_10454);
nand U13872 (N_13872,N_10089,N_9294);
nor U13873 (N_13873,N_11007,N_9341);
nor U13874 (N_13874,N_10979,N_10166);
nor U13875 (N_13875,N_10280,N_11524);
or U13876 (N_13876,N_10122,N_10709);
or U13877 (N_13877,N_11982,N_11824);
nand U13878 (N_13878,N_9915,N_10803);
xor U13879 (N_13879,N_9961,N_11605);
or U13880 (N_13880,N_9597,N_11164);
and U13881 (N_13881,N_11028,N_10590);
and U13882 (N_13882,N_10649,N_9260);
or U13883 (N_13883,N_10271,N_11750);
and U13884 (N_13884,N_11704,N_9190);
or U13885 (N_13885,N_10216,N_10522);
nor U13886 (N_13886,N_9496,N_11631);
xor U13887 (N_13887,N_10524,N_11042);
and U13888 (N_13888,N_10806,N_11764);
or U13889 (N_13889,N_11676,N_11422);
and U13890 (N_13890,N_11556,N_10214);
nor U13891 (N_13891,N_10410,N_10293);
or U13892 (N_13892,N_9527,N_11947);
xor U13893 (N_13893,N_11968,N_11677);
xor U13894 (N_13894,N_11061,N_10265);
nor U13895 (N_13895,N_11742,N_9859);
nand U13896 (N_13896,N_10017,N_11384);
nand U13897 (N_13897,N_11039,N_10799);
and U13898 (N_13898,N_10670,N_9483);
and U13899 (N_13899,N_10759,N_9471);
nor U13900 (N_13900,N_9475,N_11118);
or U13901 (N_13901,N_9756,N_10086);
or U13902 (N_13902,N_11698,N_10382);
nor U13903 (N_13903,N_11067,N_9730);
nand U13904 (N_13904,N_10871,N_11167);
nand U13905 (N_13905,N_10757,N_10427);
and U13906 (N_13906,N_11829,N_11780);
nor U13907 (N_13907,N_9624,N_10313);
nand U13908 (N_13908,N_10434,N_9668);
or U13909 (N_13909,N_10249,N_9939);
or U13910 (N_13910,N_10638,N_10558);
nand U13911 (N_13911,N_11774,N_9698);
xnor U13912 (N_13912,N_9743,N_9807);
xor U13913 (N_13913,N_9515,N_10049);
nand U13914 (N_13914,N_11391,N_11235);
nor U13915 (N_13915,N_10458,N_10628);
xor U13916 (N_13916,N_9993,N_9413);
xor U13917 (N_13917,N_10048,N_10302);
and U13918 (N_13918,N_10074,N_9128);
xor U13919 (N_13919,N_10201,N_9884);
nand U13920 (N_13920,N_11149,N_11419);
xnor U13921 (N_13921,N_10555,N_9551);
nor U13922 (N_13922,N_9954,N_10100);
nand U13923 (N_13923,N_11004,N_11226);
nor U13924 (N_13924,N_9351,N_11409);
nor U13925 (N_13925,N_11522,N_10751);
nand U13926 (N_13926,N_11844,N_9131);
and U13927 (N_13927,N_9630,N_11867);
and U13928 (N_13928,N_10111,N_11540);
nor U13929 (N_13929,N_9569,N_10502);
and U13930 (N_13930,N_11957,N_11798);
or U13931 (N_13931,N_10763,N_10878);
nor U13932 (N_13932,N_10933,N_11697);
and U13933 (N_13933,N_10786,N_9187);
and U13934 (N_13934,N_9892,N_10429);
xor U13935 (N_13935,N_11839,N_10012);
xor U13936 (N_13936,N_10932,N_9397);
nor U13937 (N_13937,N_11774,N_9373);
or U13938 (N_13938,N_9724,N_11065);
nand U13939 (N_13939,N_11155,N_9409);
or U13940 (N_13940,N_11137,N_10665);
xor U13941 (N_13941,N_9603,N_10103);
and U13942 (N_13942,N_10206,N_10327);
or U13943 (N_13943,N_9976,N_10122);
xor U13944 (N_13944,N_10960,N_11332);
or U13945 (N_13945,N_11754,N_11426);
nor U13946 (N_13946,N_9337,N_11985);
nand U13947 (N_13947,N_10328,N_11727);
and U13948 (N_13948,N_9909,N_11284);
nor U13949 (N_13949,N_11551,N_11322);
nand U13950 (N_13950,N_10050,N_11286);
and U13951 (N_13951,N_10353,N_11619);
and U13952 (N_13952,N_9945,N_11249);
or U13953 (N_13953,N_10482,N_10060);
and U13954 (N_13954,N_10920,N_9911);
or U13955 (N_13955,N_11818,N_11185);
xor U13956 (N_13956,N_11085,N_9495);
and U13957 (N_13957,N_9435,N_9516);
or U13958 (N_13958,N_11602,N_11111);
and U13959 (N_13959,N_11109,N_10536);
nand U13960 (N_13960,N_10771,N_9313);
and U13961 (N_13961,N_10154,N_11058);
nand U13962 (N_13962,N_9772,N_11563);
nand U13963 (N_13963,N_9049,N_9848);
or U13964 (N_13964,N_9563,N_10576);
or U13965 (N_13965,N_9231,N_9565);
xor U13966 (N_13966,N_10297,N_9018);
nand U13967 (N_13967,N_11669,N_9016);
nand U13968 (N_13968,N_9693,N_11604);
or U13969 (N_13969,N_10778,N_11207);
xor U13970 (N_13970,N_11117,N_10491);
nand U13971 (N_13971,N_10158,N_9149);
or U13972 (N_13972,N_10906,N_10419);
nor U13973 (N_13973,N_11829,N_9381);
and U13974 (N_13974,N_11975,N_10308);
or U13975 (N_13975,N_10232,N_9532);
nand U13976 (N_13976,N_9941,N_9450);
and U13977 (N_13977,N_9744,N_11318);
and U13978 (N_13978,N_9324,N_10047);
nand U13979 (N_13979,N_11191,N_10951);
nand U13980 (N_13980,N_9960,N_11700);
and U13981 (N_13981,N_9652,N_11193);
nand U13982 (N_13982,N_9793,N_11016);
nor U13983 (N_13983,N_10869,N_11110);
nor U13984 (N_13984,N_9193,N_10870);
nand U13985 (N_13985,N_10261,N_11685);
xor U13986 (N_13986,N_9616,N_11673);
or U13987 (N_13987,N_10305,N_10528);
or U13988 (N_13988,N_10702,N_9009);
and U13989 (N_13989,N_9120,N_10822);
or U13990 (N_13990,N_9922,N_9769);
or U13991 (N_13991,N_10858,N_11356);
xor U13992 (N_13992,N_11097,N_10996);
nor U13993 (N_13993,N_10855,N_10602);
or U13994 (N_13994,N_9405,N_10480);
xor U13995 (N_13995,N_10477,N_9440);
nor U13996 (N_13996,N_9457,N_10504);
nand U13997 (N_13997,N_11653,N_10513);
or U13998 (N_13998,N_11071,N_11953);
nor U13999 (N_13999,N_10765,N_10054);
xor U14000 (N_14000,N_9106,N_9694);
xor U14001 (N_14001,N_11444,N_9871);
and U14002 (N_14002,N_11629,N_9832);
nor U14003 (N_14003,N_11534,N_11208);
and U14004 (N_14004,N_9026,N_9126);
and U14005 (N_14005,N_9045,N_10949);
nor U14006 (N_14006,N_11572,N_10030);
nand U14007 (N_14007,N_11337,N_11382);
nand U14008 (N_14008,N_9607,N_9125);
nand U14009 (N_14009,N_11185,N_11077);
nor U14010 (N_14010,N_10579,N_10732);
xnor U14011 (N_14011,N_9223,N_9813);
or U14012 (N_14012,N_11559,N_10510);
nand U14013 (N_14013,N_9211,N_11600);
or U14014 (N_14014,N_11851,N_11453);
xor U14015 (N_14015,N_9039,N_9489);
xnor U14016 (N_14016,N_11648,N_11063);
nand U14017 (N_14017,N_9893,N_11617);
nand U14018 (N_14018,N_10286,N_10960);
or U14019 (N_14019,N_11213,N_9447);
xnor U14020 (N_14020,N_9003,N_11060);
xnor U14021 (N_14021,N_11976,N_9584);
nand U14022 (N_14022,N_11374,N_9513);
xnor U14023 (N_14023,N_11130,N_11867);
xnor U14024 (N_14024,N_9468,N_11085);
nor U14025 (N_14025,N_11930,N_9943);
nand U14026 (N_14026,N_11830,N_10402);
and U14027 (N_14027,N_10868,N_9281);
or U14028 (N_14028,N_10082,N_10146);
or U14029 (N_14029,N_11220,N_10937);
nand U14030 (N_14030,N_10069,N_11362);
xor U14031 (N_14031,N_10499,N_11325);
nor U14032 (N_14032,N_10790,N_9076);
nand U14033 (N_14033,N_9757,N_9345);
nand U14034 (N_14034,N_11646,N_9520);
nand U14035 (N_14035,N_11079,N_11956);
or U14036 (N_14036,N_10429,N_11653);
nand U14037 (N_14037,N_10070,N_11627);
or U14038 (N_14038,N_9923,N_10494);
and U14039 (N_14039,N_9776,N_11597);
xnor U14040 (N_14040,N_9551,N_11009);
xnor U14041 (N_14041,N_11139,N_10288);
nand U14042 (N_14042,N_11753,N_10309);
or U14043 (N_14043,N_10684,N_9874);
nand U14044 (N_14044,N_9567,N_10895);
xnor U14045 (N_14045,N_9949,N_9570);
nor U14046 (N_14046,N_10582,N_9994);
nor U14047 (N_14047,N_10928,N_11868);
nor U14048 (N_14048,N_10682,N_11603);
xnor U14049 (N_14049,N_10234,N_9274);
nand U14050 (N_14050,N_10053,N_10702);
nand U14051 (N_14051,N_11686,N_11241);
or U14052 (N_14052,N_10554,N_9448);
nor U14053 (N_14053,N_10249,N_9769);
nand U14054 (N_14054,N_9715,N_11432);
nand U14055 (N_14055,N_9443,N_11300);
xnor U14056 (N_14056,N_9856,N_10779);
and U14057 (N_14057,N_9819,N_9692);
nor U14058 (N_14058,N_11021,N_10440);
xnor U14059 (N_14059,N_9944,N_10079);
xnor U14060 (N_14060,N_9132,N_10197);
xor U14061 (N_14061,N_11818,N_9969);
and U14062 (N_14062,N_9122,N_11882);
and U14063 (N_14063,N_9208,N_10368);
nand U14064 (N_14064,N_11838,N_11670);
nor U14065 (N_14065,N_11123,N_9173);
and U14066 (N_14066,N_10974,N_9219);
nor U14067 (N_14067,N_9794,N_11903);
or U14068 (N_14068,N_9994,N_11518);
or U14069 (N_14069,N_11348,N_11132);
nand U14070 (N_14070,N_11927,N_10877);
nand U14071 (N_14071,N_9379,N_10451);
xor U14072 (N_14072,N_9587,N_11812);
or U14073 (N_14073,N_11331,N_10791);
xnor U14074 (N_14074,N_9343,N_9101);
and U14075 (N_14075,N_11887,N_11566);
xor U14076 (N_14076,N_11363,N_9831);
nor U14077 (N_14077,N_11799,N_10680);
and U14078 (N_14078,N_11914,N_11368);
xnor U14079 (N_14079,N_10889,N_10508);
nor U14080 (N_14080,N_11906,N_11323);
xor U14081 (N_14081,N_9628,N_11892);
xnor U14082 (N_14082,N_10063,N_10054);
xor U14083 (N_14083,N_11811,N_9733);
and U14084 (N_14084,N_11488,N_11881);
and U14085 (N_14085,N_11205,N_10410);
or U14086 (N_14086,N_11027,N_10129);
xor U14087 (N_14087,N_9630,N_11709);
or U14088 (N_14088,N_11552,N_11606);
nand U14089 (N_14089,N_9779,N_11060);
nand U14090 (N_14090,N_11013,N_11098);
and U14091 (N_14091,N_11107,N_9470);
nor U14092 (N_14092,N_10229,N_11679);
or U14093 (N_14093,N_11381,N_11049);
nand U14094 (N_14094,N_11242,N_10026);
nor U14095 (N_14095,N_9241,N_9459);
nand U14096 (N_14096,N_11232,N_11122);
nor U14097 (N_14097,N_11257,N_10480);
and U14098 (N_14098,N_11644,N_11335);
nor U14099 (N_14099,N_9444,N_9595);
and U14100 (N_14100,N_9948,N_11835);
or U14101 (N_14101,N_10334,N_9252);
nor U14102 (N_14102,N_11811,N_11086);
and U14103 (N_14103,N_10103,N_9390);
or U14104 (N_14104,N_9620,N_9208);
and U14105 (N_14105,N_11357,N_10558);
nand U14106 (N_14106,N_11551,N_10452);
and U14107 (N_14107,N_11931,N_10434);
xnor U14108 (N_14108,N_10952,N_11431);
and U14109 (N_14109,N_9565,N_11387);
and U14110 (N_14110,N_11148,N_11374);
nor U14111 (N_14111,N_10560,N_11976);
nor U14112 (N_14112,N_9461,N_11610);
or U14113 (N_14113,N_9071,N_11123);
xnor U14114 (N_14114,N_11025,N_9815);
and U14115 (N_14115,N_10643,N_11740);
xnor U14116 (N_14116,N_10530,N_9782);
and U14117 (N_14117,N_10688,N_11648);
xnor U14118 (N_14118,N_9822,N_11039);
nand U14119 (N_14119,N_10456,N_9047);
xor U14120 (N_14120,N_10117,N_10479);
nand U14121 (N_14121,N_10287,N_9769);
nand U14122 (N_14122,N_9128,N_9500);
or U14123 (N_14123,N_9035,N_11869);
nand U14124 (N_14124,N_9730,N_10464);
nand U14125 (N_14125,N_11829,N_9252);
nand U14126 (N_14126,N_10295,N_9179);
xor U14127 (N_14127,N_10247,N_9972);
or U14128 (N_14128,N_10879,N_9625);
nor U14129 (N_14129,N_9778,N_9947);
xor U14130 (N_14130,N_11563,N_11671);
nand U14131 (N_14131,N_9932,N_10925);
or U14132 (N_14132,N_11758,N_11062);
and U14133 (N_14133,N_10578,N_9810);
and U14134 (N_14134,N_11122,N_9291);
or U14135 (N_14135,N_11168,N_9756);
and U14136 (N_14136,N_9707,N_10781);
xor U14137 (N_14137,N_10715,N_9725);
nor U14138 (N_14138,N_11211,N_10766);
or U14139 (N_14139,N_10951,N_9772);
and U14140 (N_14140,N_11568,N_11291);
xor U14141 (N_14141,N_10025,N_9878);
nand U14142 (N_14142,N_11997,N_10950);
nand U14143 (N_14143,N_11548,N_10451);
or U14144 (N_14144,N_10020,N_11616);
nor U14145 (N_14145,N_10101,N_9275);
and U14146 (N_14146,N_10234,N_11304);
xor U14147 (N_14147,N_9508,N_11601);
xor U14148 (N_14148,N_9357,N_11843);
or U14149 (N_14149,N_10916,N_9752);
nor U14150 (N_14150,N_10136,N_10592);
or U14151 (N_14151,N_11304,N_10095);
nand U14152 (N_14152,N_10255,N_10467);
nor U14153 (N_14153,N_10628,N_9807);
nor U14154 (N_14154,N_11104,N_10930);
and U14155 (N_14155,N_10718,N_10328);
nor U14156 (N_14156,N_9044,N_9979);
or U14157 (N_14157,N_11149,N_9575);
or U14158 (N_14158,N_9116,N_10302);
nand U14159 (N_14159,N_11755,N_10046);
or U14160 (N_14160,N_11202,N_10336);
nor U14161 (N_14161,N_11532,N_11593);
nand U14162 (N_14162,N_9757,N_9363);
and U14163 (N_14163,N_10207,N_9649);
xnor U14164 (N_14164,N_11089,N_11450);
or U14165 (N_14165,N_11751,N_9863);
or U14166 (N_14166,N_9825,N_11990);
nand U14167 (N_14167,N_9217,N_11136);
nand U14168 (N_14168,N_9174,N_10649);
nand U14169 (N_14169,N_9861,N_11299);
nand U14170 (N_14170,N_9680,N_9362);
nor U14171 (N_14171,N_11673,N_9236);
or U14172 (N_14172,N_9586,N_9075);
xnor U14173 (N_14173,N_11854,N_11782);
xnor U14174 (N_14174,N_11389,N_11407);
xnor U14175 (N_14175,N_11952,N_9696);
xor U14176 (N_14176,N_10393,N_11380);
nand U14177 (N_14177,N_10929,N_11633);
xnor U14178 (N_14178,N_9231,N_9306);
or U14179 (N_14179,N_9613,N_9271);
nor U14180 (N_14180,N_9862,N_11877);
xor U14181 (N_14181,N_10902,N_10376);
or U14182 (N_14182,N_9648,N_11203);
xor U14183 (N_14183,N_10055,N_11713);
or U14184 (N_14184,N_11016,N_9465);
nor U14185 (N_14185,N_10705,N_10555);
nand U14186 (N_14186,N_11236,N_10681);
nor U14187 (N_14187,N_11467,N_11145);
nand U14188 (N_14188,N_11863,N_9605);
or U14189 (N_14189,N_9173,N_11688);
nor U14190 (N_14190,N_10361,N_11358);
nor U14191 (N_14191,N_10563,N_10614);
and U14192 (N_14192,N_10016,N_9870);
nand U14193 (N_14193,N_11587,N_10395);
nand U14194 (N_14194,N_9721,N_11624);
or U14195 (N_14195,N_11823,N_10444);
nor U14196 (N_14196,N_11940,N_9928);
xor U14197 (N_14197,N_9999,N_9501);
nand U14198 (N_14198,N_10144,N_11822);
or U14199 (N_14199,N_9526,N_9330);
and U14200 (N_14200,N_10859,N_9149);
nor U14201 (N_14201,N_11064,N_10467);
xnor U14202 (N_14202,N_11307,N_10050);
nand U14203 (N_14203,N_9931,N_11399);
nand U14204 (N_14204,N_10369,N_11160);
nor U14205 (N_14205,N_9277,N_11878);
nor U14206 (N_14206,N_10865,N_10677);
or U14207 (N_14207,N_11064,N_11488);
or U14208 (N_14208,N_9827,N_11273);
xnor U14209 (N_14209,N_10434,N_9037);
nor U14210 (N_14210,N_9389,N_11431);
nand U14211 (N_14211,N_11911,N_10462);
nand U14212 (N_14212,N_11136,N_10372);
nand U14213 (N_14213,N_9760,N_9435);
xor U14214 (N_14214,N_10836,N_9505);
and U14215 (N_14215,N_9950,N_10190);
or U14216 (N_14216,N_10423,N_10342);
xor U14217 (N_14217,N_9137,N_11770);
or U14218 (N_14218,N_9924,N_9789);
and U14219 (N_14219,N_11768,N_10857);
or U14220 (N_14220,N_10275,N_9080);
nor U14221 (N_14221,N_11709,N_9593);
and U14222 (N_14222,N_11754,N_9924);
and U14223 (N_14223,N_9822,N_10728);
or U14224 (N_14224,N_10487,N_10740);
or U14225 (N_14225,N_10429,N_10281);
nand U14226 (N_14226,N_11467,N_11118);
or U14227 (N_14227,N_10931,N_9647);
or U14228 (N_14228,N_10048,N_10556);
nor U14229 (N_14229,N_9700,N_9143);
xnor U14230 (N_14230,N_11088,N_11878);
nor U14231 (N_14231,N_9550,N_11384);
xor U14232 (N_14232,N_10658,N_11894);
nor U14233 (N_14233,N_10507,N_10775);
or U14234 (N_14234,N_9054,N_11022);
and U14235 (N_14235,N_9824,N_10477);
xor U14236 (N_14236,N_11000,N_9343);
or U14237 (N_14237,N_10500,N_10069);
or U14238 (N_14238,N_11875,N_9612);
xnor U14239 (N_14239,N_11295,N_10308);
or U14240 (N_14240,N_10098,N_11327);
xnor U14241 (N_14241,N_10779,N_10248);
and U14242 (N_14242,N_10692,N_9508);
and U14243 (N_14243,N_10958,N_11275);
or U14244 (N_14244,N_10780,N_9509);
nand U14245 (N_14245,N_11538,N_10672);
and U14246 (N_14246,N_9052,N_10326);
or U14247 (N_14247,N_9834,N_9071);
nor U14248 (N_14248,N_9504,N_10569);
or U14249 (N_14249,N_11537,N_9334);
nor U14250 (N_14250,N_10117,N_9499);
and U14251 (N_14251,N_10699,N_11205);
nor U14252 (N_14252,N_11038,N_10341);
and U14253 (N_14253,N_9409,N_10839);
xnor U14254 (N_14254,N_9596,N_11858);
nor U14255 (N_14255,N_11096,N_11140);
xor U14256 (N_14256,N_9668,N_9238);
nor U14257 (N_14257,N_9171,N_10227);
nand U14258 (N_14258,N_10134,N_10097);
nor U14259 (N_14259,N_10652,N_10136);
xnor U14260 (N_14260,N_10101,N_11770);
and U14261 (N_14261,N_11961,N_9086);
or U14262 (N_14262,N_10228,N_11520);
nand U14263 (N_14263,N_9888,N_10844);
and U14264 (N_14264,N_11110,N_10943);
xor U14265 (N_14265,N_9454,N_9550);
nand U14266 (N_14266,N_9022,N_9883);
nand U14267 (N_14267,N_11805,N_11664);
nor U14268 (N_14268,N_10415,N_9660);
and U14269 (N_14269,N_11414,N_9100);
nand U14270 (N_14270,N_9015,N_10331);
or U14271 (N_14271,N_9163,N_10779);
and U14272 (N_14272,N_9718,N_10246);
and U14273 (N_14273,N_9887,N_9678);
nor U14274 (N_14274,N_9008,N_10126);
or U14275 (N_14275,N_10683,N_9079);
nand U14276 (N_14276,N_9733,N_11749);
xor U14277 (N_14277,N_11698,N_11870);
and U14278 (N_14278,N_11574,N_9901);
xor U14279 (N_14279,N_9136,N_9472);
nor U14280 (N_14280,N_9379,N_10562);
nand U14281 (N_14281,N_11160,N_11196);
nor U14282 (N_14282,N_11342,N_10371);
nor U14283 (N_14283,N_11676,N_11751);
and U14284 (N_14284,N_10599,N_11563);
xor U14285 (N_14285,N_10932,N_11551);
nor U14286 (N_14286,N_11109,N_9526);
nor U14287 (N_14287,N_10068,N_9967);
xnor U14288 (N_14288,N_9173,N_10299);
or U14289 (N_14289,N_9570,N_9165);
nor U14290 (N_14290,N_9671,N_10613);
nand U14291 (N_14291,N_11197,N_9233);
xnor U14292 (N_14292,N_11636,N_10439);
nor U14293 (N_14293,N_9152,N_11308);
and U14294 (N_14294,N_9836,N_11642);
xnor U14295 (N_14295,N_10504,N_11849);
nor U14296 (N_14296,N_9043,N_11154);
or U14297 (N_14297,N_10242,N_10897);
and U14298 (N_14298,N_10742,N_9332);
xor U14299 (N_14299,N_11116,N_9879);
or U14300 (N_14300,N_9770,N_9510);
nor U14301 (N_14301,N_11376,N_10750);
nand U14302 (N_14302,N_11035,N_9731);
xnor U14303 (N_14303,N_11511,N_10762);
and U14304 (N_14304,N_9179,N_10514);
nor U14305 (N_14305,N_9823,N_11688);
nor U14306 (N_14306,N_11981,N_11589);
nand U14307 (N_14307,N_9159,N_10221);
xnor U14308 (N_14308,N_11773,N_9305);
xor U14309 (N_14309,N_10218,N_10883);
and U14310 (N_14310,N_9136,N_10957);
nor U14311 (N_14311,N_11423,N_11926);
or U14312 (N_14312,N_9540,N_9630);
and U14313 (N_14313,N_11017,N_9296);
xnor U14314 (N_14314,N_9920,N_11297);
xnor U14315 (N_14315,N_11355,N_11090);
or U14316 (N_14316,N_11262,N_10045);
xnor U14317 (N_14317,N_11905,N_11097);
nand U14318 (N_14318,N_11782,N_10740);
xnor U14319 (N_14319,N_11760,N_9834);
nand U14320 (N_14320,N_10821,N_11563);
or U14321 (N_14321,N_11011,N_10149);
or U14322 (N_14322,N_10820,N_9546);
xor U14323 (N_14323,N_11760,N_11060);
or U14324 (N_14324,N_10520,N_10781);
nand U14325 (N_14325,N_9142,N_10426);
or U14326 (N_14326,N_9577,N_9824);
xor U14327 (N_14327,N_9604,N_9827);
nand U14328 (N_14328,N_11210,N_11168);
nand U14329 (N_14329,N_9532,N_11265);
nand U14330 (N_14330,N_9722,N_10889);
xnor U14331 (N_14331,N_11693,N_10782);
nor U14332 (N_14332,N_10317,N_11902);
or U14333 (N_14333,N_10609,N_9252);
xnor U14334 (N_14334,N_9796,N_11748);
xor U14335 (N_14335,N_10320,N_10295);
or U14336 (N_14336,N_11133,N_10603);
and U14337 (N_14337,N_10805,N_11691);
xnor U14338 (N_14338,N_9654,N_11517);
xor U14339 (N_14339,N_9188,N_11879);
xor U14340 (N_14340,N_9895,N_10905);
nand U14341 (N_14341,N_9532,N_10133);
nand U14342 (N_14342,N_9652,N_10175);
nor U14343 (N_14343,N_9601,N_11409);
xor U14344 (N_14344,N_10755,N_9558);
or U14345 (N_14345,N_9251,N_10453);
nand U14346 (N_14346,N_10209,N_10753);
nand U14347 (N_14347,N_9677,N_9428);
or U14348 (N_14348,N_9706,N_11196);
nor U14349 (N_14349,N_10059,N_11691);
xnor U14350 (N_14350,N_10698,N_9668);
and U14351 (N_14351,N_11636,N_9888);
and U14352 (N_14352,N_11949,N_9973);
nand U14353 (N_14353,N_9121,N_11653);
nor U14354 (N_14354,N_10026,N_10982);
nor U14355 (N_14355,N_11664,N_9772);
xor U14356 (N_14356,N_9453,N_11655);
and U14357 (N_14357,N_10011,N_10748);
and U14358 (N_14358,N_10209,N_10671);
xor U14359 (N_14359,N_11097,N_9876);
nand U14360 (N_14360,N_9485,N_11828);
or U14361 (N_14361,N_11393,N_9800);
nor U14362 (N_14362,N_9592,N_11615);
xnor U14363 (N_14363,N_9415,N_10160);
xnor U14364 (N_14364,N_9775,N_10806);
nand U14365 (N_14365,N_11040,N_10503);
xor U14366 (N_14366,N_11751,N_10219);
nor U14367 (N_14367,N_9968,N_10428);
xor U14368 (N_14368,N_10892,N_11258);
or U14369 (N_14369,N_11646,N_10610);
or U14370 (N_14370,N_11987,N_9415);
nand U14371 (N_14371,N_10994,N_10408);
or U14372 (N_14372,N_11326,N_10962);
nor U14373 (N_14373,N_9421,N_11241);
nor U14374 (N_14374,N_10647,N_11687);
or U14375 (N_14375,N_11327,N_10831);
nand U14376 (N_14376,N_11862,N_11361);
and U14377 (N_14377,N_10089,N_10414);
nor U14378 (N_14378,N_11148,N_9326);
and U14379 (N_14379,N_11263,N_9698);
nand U14380 (N_14380,N_9806,N_10185);
xnor U14381 (N_14381,N_10930,N_10712);
or U14382 (N_14382,N_10686,N_9965);
or U14383 (N_14383,N_11017,N_10892);
nand U14384 (N_14384,N_9406,N_11368);
and U14385 (N_14385,N_11360,N_11358);
nor U14386 (N_14386,N_11316,N_10544);
nor U14387 (N_14387,N_11815,N_10687);
and U14388 (N_14388,N_9326,N_10740);
and U14389 (N_14389,N_10625,N_10016);
nor U14390 (N_14390,N_11815,N_11004);
or U14391 (N_14391,N_11505,N_10840);
nor U14392 (N_14392,N_11170,N_10532);
xor U14393 (N_14393,N_10500,N_9614);
xor U14394 (N_14394,N_10872,N_11734);
and U14395 (N_14395,N_9483,N_10955);
and U14396 (N_14396,N_10333,N_9435);
xnor U14397 (N_14397,N_11822,N_11097);
or U14398 (N_14398,N_10391,N_10793);
and U14399 (N_14399,N_9242,N_10865);
nor U14400 (N_14400,N_9116,N_11533);
nor U14401 (N_14401,N_9820,N_11602);
nor U14402 (N_14402,N_10522,N_11217);
nand U14403 (N_14403,N_9832,N_11137);
nor U14404 (N_14404,N_11880,N_9824);
nand U14405 (N_14405,N_9900,N_9171);
nor U14406 (N_14406,N_10950,N_10002);
nor U14407 (N_14407,N_11897,N_10651);
or U14408 (N_14408,N_9506,N_11776);
and U14409 (N_14409,N_9056,N_10180);
and U14410 (N_14410,N_11134,N_9587);
nand U14411 (N_14411,N_10721,N_11787);
nor U14412 (N_14412,N_10520,N_9814);
nor U14413 (N_14413,N_9027,N_9620);
xnor U14414 (N_14414,N_11344,N_11312);
and U14415 (N_14415,N_9100,N_9444);
or U14416 (N_14416,N_11436,N_11422);
and U14417 (N_14417,N_11892,N_11521);
and U14418 (N_14418,N_10677,N_9491);
nor U14419 (N_14419,N_10607,N_9591);
nor U14420 (N_14420,N_11953,N_9197);
nor U14421 (N_14421,N_9667,N_11881);
or U14422 (N_14422,N_10766,N_11515);
or U14423 (N_14423,N_11983,N_11103);
nor U14424 (N_14424,N_11903,N_9956);
and U14425 (N_14425,N_11364,N_9122);
nand U14426 (N_14426,N_11482,N_9957);
xor U14427 (N_14427,N_9946,N_9300);
or U14428 (N_14428,N_9163,N_10139);
or U14429 (N_14429,N_11917,N_10994);
and U14430 (N_14430,N_9044,N_9562);
or U14431 (N_14431,N_11606,N_10720);
nand U14432 (N_14432,N_9396,N_11714);
and U14433 (N_14433,N_10822,N_11616);
nand U14434 (N_14434,N_9888,N_10994);
or U14435 (N_14435,N_11096,N_10296);
nand U14436 (N_14436,N_9837,N_10942);
or U14437 (N_14437,N_10869,N_9017);
nor U14438 (N_14438,N_9320,N_9250);
or U14439 (N_14439,N_10799,N_9902);
or U14440 (N_14440,N_11971,N_11043);
xnor U14441 (N_14441,N_9530,N_11072);
and U14442 (N_14442,N_9992,N_9792);
xor U14443 (N_14443,N_10459,N_9203);
or U14444 (N_14444,N_9886,N_11068);
xnor U14445 (N_14445,N_9973,N_10554);
and U14446 (N_14446,N_10495,N_11445);
xor U14447 (N_14447,N_9913,N_10823);
and U14448 (N_14448,N_11475,N_9230);
and U14449 (N_14449,N_10477,N_11016);
or U14450 (N_14450,N_10827,N_10581);
nand U14451 (N_14451,N_11571,N_11102);
or U14452 (N_14452,N_10810,N_11909);
nor U14453 (N_14453,N_10999,N_10696);
and U14454 (N_14454,N_9220,N_10448);
nand U14455 (N_14455,N_11617,N_10646);
and U14456 (N_14456,N_11489,N_10811);
xor U14457 (N_14457,N_11097,N_11786);
nand U14458 (N_14458,N_9328,N_9823);
nand U14459 (N_14459,N_10005,N_9859);
nand U14460 (N_14460,N_9474,N_9720);
or U14461 (N_14461,N_9624,N_9061);
nand U14462 (N_14462,N_10642,N_10089);
nor U14463 (N_14463,N_9783,N_9884);
nand U14464 (N_14464,N_10974,N_9243);
and U14465 (N_14465,N_11578,N_11553);
or U14466 (N_14466,N_9810,N_10125);
nand U14467 (N_14467,N_11895,N_9864);
nand U14468 (N_14468,N_11889,N_9514);
or U14469 (N_14469,N_11903,N_11734);
or U14470 (N_14470,N_9822,N_9351);
xnor U14471 (N_14471,N_10757,N_10005);
xnor U14472 (N_14472,N_10019,N_10760);
nand U14473 (N_14473,N_10051,N_9566);
xor U14474 (N_14474,N_11187,N_10917);
xnor U14475 (N_14475,N_9323,N_10233);
or U14476 (N_14476,N_11283,N_10701);
nor U14477 (N_14477,N_11025,N_9893);
nand U14478 (N_14478,N_10334,N_10615);
nor U14479 (N_14479,N_11147,N_10424);
or U14480 (N_14480,N_10289,N_11700);
or U14481 (N_14481,N_11247,N_10603);
and U14482 (N_14482,N_11602,N_9172);
nand U14483 (N_14483,N_10492,N_11556);
nor U14484 (N_14484,N_9184,N_9664);
xor U14485 (N_14485,N_11900,N_10361);
xor U14486 (N_14486,N_9915,N_10792);
xnor U14487 (N_14487,N_10090,N_10886);
xnor U14488 (N_14488,N_11144,N_11975);
xnor U14489 (N_14489,N_10116,N_10104);
and U14490 (N_14490,N_11910,N_11060);
or U14491 (N_14491,N_10672,N_10706);
or U14492 (N_14492,N_10878,N_9331);
and U14493 (N_14493,N_9684,N_11304);
or U14494 (N_14494,N_10985,N_10299);
nand U14495 (N_14495,N_11104,N_10348);
nor U14496 (N_14496,N_9500,N_11304);
and U14497 (N_14497,N_11906,N_11547);
nand U14498 (N_14498,N_9254,N_9949);
nor U14499 (N_14499,N_11524,N_11411);
nand U14500 (N_14500,N_11489,N_10007);
nand U14501 (N_14501,N_9754,N_10319);
xnor U14502 (N_14502,N_11684,N_9295);
and U14503 (N_14503,N_9443,N_10012);
xor U14504 (N_14504,N_11743,N_10322);
xor U14505 (N_14505,N_9659,N_9870);
or U14506 (N_14506,N_9252,N_9469);
xnor U14507 (N_14507,N_9755,N_9021);
nor U14508 (N_14508,N_10228,N_11301);
nor U14509 (N_14509,N_9440,N_9003);
and U14510 (N_14510,N_10633,N_11870);
and U14511 (N_14511,N_10285,N_10375);
and U14512 (N_14512,N_10821,N_9455);
or U14513 (N_14513,N_10082,N_9495);
xnor U14514 (N_14514,N_11659,N_10087);
nand U14515 (N_14515,N_9953,N_9350);
and U14516 (N_14516,N_10364,N_9626);
xnor U14517 (N_14517,N_11650,N_10403);
xor U14518 (N_14518,N_11870,N_11982);
or U14519 (N_14519,N_11279,N_9266);
nand U14520 (N_14520,N_11584,N_11667);
or U14521 (N_14521,N_10711,N_9643);
or U14522 (N_14522,N_10628,N_10760);
nor U14523 (N_14523,N_9463,N_9935);
or U14524 (N_14524,N_9376,N_11814);
nor U14525 (N_14525,N_9260,N_10029);
xnor U14526 (N_14526,N_9354,N_11729);
and U14527 (N_14527,N_11592,N_9165);
xnor U14528 (N_14528,N_11320,N_10875);
and U14529 (N_14529,N_11192,N_9792);
or U14530 (N_14530,N_9538,N_9835);
nand U14531 (N_14531,N_11332,N_10405);
and U14532 (N_14532,N_11605,N_9266);
nor U14533 (N_14533,N_9993,N_9281);
and U14534 (N_14534,N_11652,N_11684);
and U14535 (N_14535,N_10223,N_9364);
or U14536 (N_14536,N_11165,N_11378);
xor U14537 (N_14537,N_10972,N_9171);
xor U14538 (N_14538,N_9965,N_10244);
xor U14539 (N_14539,N_9958,N_9945);
xor U14540 (N_14540,N_9831,N_11669);
and U14541 (N_14541,N_11246,N_10213);
or U14542 (N_14542,N_10003,N_11995);
nor U14543 (N_14543,N_11362,N_9696);
or U14544 (N_14544,N_11309,N_11590);
xor U14545 (N_14545,N_10077,N_10641);
nor U14546 (N_14546,N_11928,N_11111);
xor U14547 (N_14547,N_10216,N_10169);
or U14548 (N_14548,N_9407,N_9492);
and U14549 (N_14549,N_10093,N_11705);
and U14550 (N_14550,N_10703,N_10354);
nand U14551 (N_14551,N_9292,N_11638);
nand U14552 (N_14552,N_11318,N_9467);
nand U14553 (N_14553,N_11478,N_9391);
and U14554 (N_14554,N_10919,N_11692);
nand U14555 (N_14555,N_9806,N_11948);
or U14556 (N_14556,N_10293,N_9615);
or U14557 (N_14557,N_9078,N_11197);
and U14558 (N_14558,N_10859,N_11367);
nand U14559 (N_14559,N_10119,N_10874);
and U14560 (N_14560,N_10319,N_9426);
nand U14561 (N_14561,N_9175,N_9991);
nor U14562 (N_14562,N_10023,N_9765);
nor U14563 (N_14563,N_10859,N_9692);
and U14564 (N_14564,N_11001,N_11819);
and U14565 (N_14565,N_9615,N_10836);
xnor U14566 (N_14566,N_11969,N_9381);
or U14567 (N_14567,N_11198,N_10474);
nor U14568 (N_14568,N_10744,N_10106);
nand U14569 (N_14569,N_9247,N_9682);
or U14570 (N_14570,N_11161,N_10804);
and U14571 (N_14571,N_11321,N_9584);
nand U14572 (N_14572,N_10610,N_11952);
nand U14573 (N_14573,N_9644,N_11963);
and U14574 (N_14574,N_11105,N_11663);
nor U14575 (N_14575,N_9857,N_11839);
or U14576 (N_14576,N_9242,N_11079);
nand U14577 (N_14577,N_11034,N_10413);
or U14578 (N_14578,N_10686,N_11435);
or U14579 (N_14579,N_9690,N_9652);
or U14580 (N_14580,N_10131,N_9917);
nand U14581 (N_14581,N_10709,N_11097);
nor U14582 (N_14582,N_9100,N_9470);
nor U14583 (N_14583,N_11277,N_10971);
nor U14584 (N_14584,N_10526,N_9564);
nor U14585 (N_14585,N_9108,N_9212);
nand U14586 (N_14586,N_11547,N_10400);
nand U14587 (N_14587,N_10910,N_10396);
nor U14588 (N_14588,N_11754,N_10216);
xnor U14589 (N_14589,N_11598,N_9522);
and U14590 (N_14590,N_9353,N_10881);
xnor U14591 (N_14591,N_11118,N_11743);
nand U14592 (N_14592,N_9897,N_9002);
xor U14593 (N_14593,N_11340,N_9825);
nor U14594 (N_14594,N_10368,N_9770);
xnor U14595 (N_14595,N_9240,N_11452);
or U14596 (N_14596,N_11892,N_11471);
nand U14597 (N_14597,N_9008,N_11383);
xor U14598 (N_14598,N_11256,N_11492);
or U14599 (N_14599,N_10075,N_10481);
nand U14600 (N_14600,N_9033,N_9984);
or U14601 (N_14601,N_10613,N_10277);
xor U14602 (N_14602,N_10090,N_9024);
xor U14603 (N_14603,N_11608,N_11924);
nor U14604 (N_14604,N_10559,N_9495);
nor U14605 (N_14605,N_9423,N_10809);
nand U14606 (N_14606,N_10973,N_10741);
and U14607 (N_14607,N_9785,N_9339);
and U14608 (N_14608,N_10367,N_11643);
xnor U14609 (N_14609,N_11405,N_11863);
nor U14610 (N_14610,N_10611,N_9546);
or U14611 (N_14611,N_9271,N_11442);
and U14612 (N_14612,N_11195,N_11808);
nor U14613 (N_14613,N_10179,N_9687);
or U14614 (N_14614,N_10098,N_10331);
xnor U14615 (N_14615,N_10080,N_10689);
nand U14616 (N_14616,N_11601,N_11830);
nand U14617 (N_14617,N_10983,N_10853);
nand U14618 (N_14618,N_9559,N_9143);
nand U14619 (N_14619,N_11432,N_10810);
nand U14620 (N_14620,N_10972,N_11398);
nand U14621 (N_14621,N_9378,N_10610);
xor U14622 (N_14622,N_9227,N_9470);
or U14623 (N_14623,N_10964,N_9600);
and U14624 (N_14624,N_10574,N_9118);
or U14625 (N_14625,N_9415,N_10474);
nand U14626 (N_14626,N_9362,N_9386);
nor U14627 (N_14627,N_10830,N_11722);
xnor U14628 (N_14628,N_10589,N_11797);
nand U14629 (N_14629,N_9412,N_11054);
or U14630 (N_14630,N_11358,N_9789);
and U14631 (N_14631,N_11583,N_9854);
or U14632 (N_14632,N_9086,N_11478);
nor U14633 (N_14633,N_9878,N_9445);
and U14634 (N_14634,N_9271,N_11010);
and U14635 (N_14635,N_11457,N_9783);
or U14636 (N_14636,N_9885,N_11873);
or U14637 (N_14637,N_10482,N_11463);
nand U14638 (N_14638,N_9487,N_11837);
or U14639 (N_14639,N_9245,N_11597);
nor U14640 (N_14640,N_10668,N_10449);
nand U14641 (N_14641,N_11849,N_11862);
nor U14642 (N_14642,N_11723,N_9249);
nand U14643 (N_14643,N_9198,N_11122);
and U14644 (N_14644,N_9254,N_10424);
nor U14645 (N_14645,N_9419,N_11760);
nor U14646 (N_14646,N_9354,N_10769);
or U14647 (N_14647,N_10935,N_10731);
or U14648 (N_14648,N_11786,N_9374);
nor U14649 (N_14649,N_9964,N_10658);
nand U14650 (N_14650,N_11645,N_10795);
and U14651 (N_14651,N_11183,N_11819);
or U14652 (N_14652,N_10158,N_11033);
and U14653 (N_14653,N_10871,N_11711);
or U14654 (N_14654,N_9233,N_11223);
nand U14655 (N_14655,N_10262,N_10922);
xor U14656 (N_14656,N_9860,N_10075);
nand U14657 (N_14657,N_10527,N_9324);
nand U14658 (N_14658,N_9259,N_10983);
and U14659 (N_14659,N_11325,N_9135);
nand U14660 (N_14660,N_9005,N_11625);
and U14661 (N_14661,N_11026,N_9702);
and U14662 (N_14662,N_9734,N_11257);
xnor U14663 (N_14663,N_10411,N_11283);
nor U14664 (N_14664,N_11154,N_10997);
and U14665 (N_14665,N_10481,N_9082);
or U14666 (N_14666,N_10079,N_9674);
nor U14667 (N_14667,N_9248,N_10985);
nand U14668 (N_14668,N_9333,N_9831);
and U14669 (N_14669,N_11127,N_11841);
and U14670 (N_14670,N_9943,N_9574);
xnor U14671 (N_14671,N_10574,N_11728);
and U14672 (N_14672,N_10005,N_11413);
or U14673 (N_14673,N_11247,N_11867);
xor U14674 (N_14674,N_9433,N_11401);
nand U14675 (N_14675,N_11416,N_9953);
nand U14676 (N_14676,N_10546,N_10873);
nor U14677 (N_14677,N_9336,N_11033);
nor U14678 (N_14678,N_10817,N_10308);
nor U14679 (N_14679,N_9031,N_10571);
and U14680 (N_14680,N_11029,N_11608);
nand U14681 (N_14681,N_11793,N_11189);
xnor U14682 (N_14682,N_9544,N_9970);
nor U14683 (N_14683,N_10250,N_10702);
xnor U14684 (N_14684,N_10355,N_9334);
nor U14685 (N_14685,N_9477,N_11158);
nor U14686 (N_14686,N_9147,N_11790);
and U14687 (N_14687,N_11090,N_9878);
nor U14688 (N_14688,N_11584,N_11355);
and U14689 (N_14689,N_9912,N_11252);
nand U14690 (N_14690,N_9261,N_10161);
and U14691 (N_14691,N_9763,N_10957);
xor U14692 (N_14692,N_10149,N_9536);
nand U14693 (N_14693,N_9361,N_10184);
xor U14694 (N_14694,N_9586,N_11679);
nand U14695 (N_14695,N_10087,N_11600);
xor U14696 (N_14696,N_11908,N_9713);
xnor U14697 (N_14697,N_9497,N_11333);
or U14698 (N_14698,N_9256,N_9854);
nand U14699 (N_14699,N_10048,N_9415);
nand U14700 (N_14700,N_10919,N_11196);
and U14701 (N_14701,N_10656,N_11729);
nand U14702 (N_14702,N_10325,N_11169);
nand U14703 (N_14703,N_9017,N_9431);
xnor U14704 (N_14704,N_11619,N_11896);
nor U14705 (N_14705,N_9676,N_9969);
and U14706 (N_14706,N_11500,N_10281);
xnor U14707 (N_14707,N_11715,N_9147);
nand U14708 (N_14708,N_11483,N_11084);
nor U14709 (N_14709,N_11016,N_9018);
and U14710 (N_14710,N_10886,N_10277);
or U14711 (N_14711,N_10224,N_10579);
nand U14712 (N_14712,N_11406,N_11240);
nor U14713 (N_14713,N_11885,N_11181);
xnor U14714 (N_14714,N_10090,N_10692);
xnor U14715 (N_14715,N_11725,N_9993);
nor U14716 (N_14716,N_9811,N_10469);
nor U14717 (N_14717,N_9490,N_10930);
nor U14718 (N_14718,N_9445,N_11383);
xnor U14719 (N_14719,N_9980,N_10076);
nor U14720 (N_14720,N_10495,N_11840);
nand U14721 (N_14721,N_11752,N_10360);
nor U14722 (N_14722,N_11033,N_9956);
nand U14723 (N_14723,N_10232,N_11532);
and U14724 (N_14724,N_11850,N_9485);
nor U14725 (N_14725,N_9586,N_11574);
and U14726 (N_14726,N_10407,N_11749);
or U14727 (N_14727,N_11383,N_9836);
and U14728 (N_14728,N_11287,N_11194);
nor U14729 (N_14729,N_10802,N_10556);
nor U14730 (N_14730,N_10055,N_10256);
and U14731 (N_14731,N_10086,N_11057);
and U14732 (N_14732,N_10430,N_9443);
and U14733 (N_14733,N_10590,N_11630);
xor U14734 (N_14734,N_10538,N_11897);
and U14735 (N_14735,N_10060,N_11287);
nor U14736 (N_14736,N_11281,N_10734);
or U14737 (N_14737,N_10333,N_10895);
xnor U14738 (N_14738,N_11962,N_10642);
nor U14739 (N_14739,N_9461,N_9862);
or U14740 (N_14740,N_11419,N_9394);
xor U14741 (N_14741,N_10560,N_9079);
nor U14742 (N_14742,N_9652,N_11793);
nand U14743 (N_14743,N_11455,N_10108);
nand U14744 (N_14744,N_9874,N_9601);
and U14745 (N_14745,N_10573,N_11383);
nor U14746 (N_14746,N_9810,N_11710);
nand U14747 (N_14747,N_9711,N_11546);
xor U14748 (N_14748,N_11624,N_9402);
or U14749 (N_14749,N_10596,N_11543);
or U14750 (N_14750,N_10365,N_9233);
xnor U14751 (N_14751,N_11851,N_9080);
nand U14752 (N_14752,N_10082,N_9096);
xnor U14753 (N_14753,N_9850,N_10861);
nor U14754 (N_14754,N_11293,N_11876);
or U14755 (N_14755,N_11778,N_10134);
xor U14756 (N_14756,N_11973,N_10579);
xnor U14757 (N_14757,N_9481,N_11226);
nand U14758 (N_14758,N_11633,N_10061);
and U14759 (N_14759,N_9713,N_11175);
nor U14760 (N_14760,N_10853,N_10476);
xnor U14761 (N_14761,N_9681,N_9363);
nor U14762 (N_14762,N_10605,N_9028);
nand U14763 (N_14763,N_10734,N_10863);
and U14764 (N_14764,N_11375,N_10204);
nand U14765 (N_14765,N_10031,N_10909);
or U14766 (N_14766,N_11512,N_11609);
nor U14767 (N_14767,N_9553,N_9725);
and U14768 (N_14768,N_11651,N_10827);
nand U14769 (N_14769,N_9211,N_9336);
nand U14770 (N_14770,N_10799,N_11201);
nand U14771 (N_14771,N_9847,N_10856);
and U14772 (N_14772,N_9970,N_10068);
and U14773 (N_14773,N_9739,N_10488);
nor U14774 (N_14774,N_10353,N_9497);
nor U14775 (N_14775,N_10276,N_11748);
or U14776 (N_14776,N_11771,N_9488);
and U14777 (N_14777,N_10609,N_11462);
nor U14778 (N_14778,N_10656,N_10012);
or U14779 (N_14779,N_9490,N_11926);
nand U14780 (N_14780,N_11573,N_10373);
nand U14781 (N_14781,N_9357,N_9040);
nand U14782 (N_14782,N_11809,N_10331);
or U14783 (N_14783,N_9763,N_10275);
nand U14784 (N_14784,N_11623,N_9675);
nand U14785 (N_14785,N_11639,N_10289);
or U14786 (N_14786,N_10539,N_9123);
or U14787 (N_14787,N_11616,N_11201);
or U14788 (N_14788,N_11140,N_9431);
nor U14789 (N_14789,N_9119,N_10234);
and U14790 (N_14790,N_11102,N_9384);
and U14791 (N_14791,N_11012,N_9008);
nand U14792 (N_14792,N_9228,N_11314);
or U14793 (N_14793,N_11467,N_11131);
and U14794 (N_14794,N_11356,N_10157);
nor U14795 (N_14795,N_9707,N_11197);
or U14796 (N_14796,N_9317,N_11861);
xor U14797 (N_14797,N_9886,N_10138);
or U14798 (N_14798,N_9667,N_9600);
nor U14799 (N_14799,N_9085,N_11198);
nand U14800 (N_14800,N_11759,N_10761);
and U14801 (N_14801,N_10706,N_10714);
or U14802 (N_14802,N_9191,N_11429);
and U14803 (N_14803,N_11824,N_9270);
nand U14804 (N_14804,N_9460,N_9475);
nand U14805 (N_14805,N_10180,N_11167);
or U14806 (N_14806,N_9666,N_9684);
and U14807 (N_14807,N_11120,N_10924);
xnor U14808 (N_14808,N_11532,N_9094);
nand U14809 (N_14809,N_11267,N_11835);
nor U14810 (N_14810,N_11392,N_10406);
xnor U14811 (N_14811,N_11627,N_9569);
nand U14812 (N_14812,N_10883,N_9320);
and U14813 (N_14813,N_9843,N_9628);
nand U14814 (N_14814,N_10836,N_9043);
and U14815 (N_14815,N_10465,N_9882);
and U14816 (N_14816,N_10152,N_9636);
or U14817 (N_14817,N_10732,N_10890);
and U14818 (N_14818,N_10590,N_9048);
or U14819 (N_14819,N_10580,N_11860);
or U14820 (N_14820,N_9370,N_9421);
and U14821 (N_14821,N_10510,N_10095);
nand U14822 (N_14822,N_9955,N_11663);
nor U14823 (N_14823,N_9879,N_10326);
xnor U14824 (N_14824,N_11830,N_10108);
nor U14825 (N_14825,N_10865,N_9192);
nor U14826 (N_14826,N_9394,N_11969);
nor U14827 (N_14827,N_11173,N_9469);
and U14828 (N_14828,N_10380,N_9206);
nor U14829 (N_14829,N_11123,N_11851);
and U14830 (N_14830,N_10868,N_10327);
and U14831 (N_14831,N_11674,N_11361);
or U14832 (N_14832,N_9231,N_11518);
nand U14833 (N_14833,N_10116,N_10547);
or U14834 (N_14834,N_10475,N_9051);
or U14835 (N_14835,N_10711,N_9429);
nor U14836 (N_14836,N_11148,N_10023);
nor U14837 (N_14837,N_11367,N_10600);
or U14838 (N_14838,N_10720,N_11116);
nand U14839 (N_14839,N_10647,N_11825);
or U14840 (N_14840,N_9384,N_11422);
nor U14841 (N_14841,N_10897,N_9356);
nor U14842 (N_14842,N_10266,N_9420);
nor U14843 (N_14843,N_9068,N_9016);
nand U14844 (N_14844,N_9830,N_10652);
and U14845 (N_14845,N_10049,N_10170);
and U14846 (N_14846,N_9363,N_11484);
or U14847 (N_14847,N_11525,N_10497);
nor U14848 (N_14848,N_10305,N_9490);
nor U14849 (N_14849,N_9312,N_9369);
nor U14850 (N_14850,N_9175,N_9763);
and U14851 (N_14851,N_11407,N_9675);
and U14852 (N_14852,N_10969,N_10439);
xor U14853 (N_14853,N_9510,N_9118);
and U14854 (N_14854,N_10117,N_9258);
nor U14855 (N_14855,N_10488,N_11660);
or U14856 (N_14856,N_11890,N_10487);
nand U14857 (N_14857,N_9637,N_11615);
nor U14858 (N_14858,N_10395,N_9123);
xnor U14859 (N_14859,N_11495,N_11263);
and U14860 (N_14860,N_10104,N_11831);
xor U14861 (N_14861,N_10474,N_10449);
nand U14862 (N_14862,N_10163,N_10203);
nor U14863 (N_14863,N_9585,N_11541);
or U14864 (N_14864,N_9625,N_9315);
nand U14865 (N_14865,N_9891,N_9991);
nand U14866 (N_14866,N_11862,N_11145);
nor U14867 (N_14867,N_9718,N_10334);
nor U14868 (N_14868,N_9392,N_10289);
and U14869 (N_14869,N_9865,N_9665);
and U14870 (N_14870,N_11176,N_9057);
nor U14871 (N_14871,N_11461,N_9604);
or U14872 (N_14872,N_10489,N_11536);
nor U14873 (N_14873,N_10744,N_9383);
nand U14874 (N_14874,N_11588,N_9067);
or U14875 (N_14875,N_11317,N_9369);
xnor U14876 (N_14876,N_9409,N_9383);
xnor U14877 (N_14877,N_9141,N_9427);
or U14878 (N_14878,N_9124,N_10490);
or U14879 (N_14879,N_10334,N_10817);
or U14880 (N_14880,N_11465,N_9695);
nor U14881 (N_14881,N_9193,N_9661);
nor U14882 (N_14882,N_9688,N_9292);
or U14883 (N_14883,N_11549,N_10650);
nand U14884 (N_14884,N_10017,N_9725);
and U14885 (N_14885,N_10483,N_11709);
nand U14886 (N_14886,N_11709,N_10768);
and U14887 (N_14887,N_10836,N_11629);
or U14888 (N_14888,N_10470,N_9896);
or U14889 (N_14889,N_9723,N_9636);
nand U14890 (N_14890,N_9641,N_9075);
nand U14891 (N_14891,N_10076,N_10191);
or U14892 (N_14892,N_10502,N_10823);
nor U14893 (N_14893,N_10744,N_9108);
or U14894 (N_14894,N_11272,N_10385);
and U14895 (N_14895,N_9405,N_11348);
and U14896 (N_14896,N_9208,N_11380);
nand U14897 (N_14897,N_9673,N_11305);
or U14898 (N_14898,N_9696,N_11079);
or U14899 (N_14899,N_10880,N_11256);
nor U14900 (N_14900,N_10952,N_11582);
nor U14901 (N_14901,N_10103,N_9839);
nor U14902 (N_14902,N_11533,N_11233);
nor U14903 (N_14903,N_10305,N_9285);
nor U14904 (N_14904,N_11928,N_11184);
nand U14905 (N_14905,N_11175,N_10060);
xnor U14906 (N_14906,N_10399,N_9953);
nor U14907 (N_14907,N_10570,N_10320);
nor U14908 (N_14908,N_11922,N_11296);
xor U14909 (N_14909,N_11607,N_9559);
xnor U14910 (N_14910,N_11933,N_11525);
nand U14911 (N_14911,N_11730,N_9395);
nand U14912 (N_14912,N_11485,N_11124);
nand U14913 (N_14913,N_10196,N_10126);
nor U14914 (N_14914,N_11659,N_10580);
xnor U14915 (N_14915,N_10403,N_9883);
nor U14916 (N_14916,N_9178,N_11230);
nor U14917 (N_14917,N_9995,N_10276);
xnor U14918 (N_14918,N_10718,N_9945);
nand U14919 (N_14919,N_9743,N_10460);
nor U14920 (N_14920,N_9222,N_10854);
or U14921 (N_14921,N_10352,N_10225);
nor U14922 (N_14922,N_11234,N_9430);
nor U14923 (N_14923,N_11765,N_9615);
nand U14924 (N_14924,N_9275,N_11662);
xor U14925 (N_14925,N_11485,N_11695);
and U14926 (N_14926,N_9094,N_10145);
nor U14927 (N_14927,N_11613,N_9410);
nand U14928 (N_14928,N_9387,N_11436);
nand U14929 (N_14929,N_10652,N_10310);
or U14930 (N_14930,N_10490,N_9304);
or U14931 (N_14931,N_10491,N_10084);
xnor U14932 (N_14932,N_11644,N_11990);
nand U14933 (N_14933,N_11203,N_11830);
nor U14934 (N_14934,N_9202,N_9473);
nand U14935 (N_14935,N_10681,N_9840);
nand U14936 (N_14936,N_9416,N_11565);
and U14937 (N_14937,N_11789,N_11244);
xor U14938 (N_14938,N_10755,N_9565);
or U14939 (N_14939,N_9959,N_9654);
and U14940 (N_14940,N_11699,N_11367);
and U14941 (N_14941,N_9420,N_11587);
xor U14942 (N_14942,N_9298,N_11648);
nor U14943 (N_14943,N_10573,N_10536);
xor U14944 (N_14944,N_9974,N_9817);
and U14945 (N_14945,N_11830,N_10506);
nor U14946 (N_14946,N_10790,N_9868);
nor U14947 (N_14947,N_10919,N_11353);
xor U14948 (N_14948,N_9209,N_9680);
nor U14949 (N_14949,N_9637,N_11057);
and U14950 (N_14950,N_9348,N_9937);
nand U14951 (N_14951,N_11827,N_10619);
xnor U14952 (N_14952,N_11402,N_10795);
or U14953 (N_14953,N_10034,N_9090);
nor U14954 (N_14954,N_11136,N_11824);
nand U14955 (N_14955,N_11328,N_11085);
and U14956 (N_14956,N_10562,N_9157);
xnor U14957 (N_14957,N_9568,N_11137);
or U14958 (N_14958,N_11603,N_9144);
or U14959 (N_14959,N_11495,N_10563);
xor U14960 (N_14960,N_9110,N_11145);
xor U14961 (N_14961,N_11804,N_10998);
nand U14962 (N_14962,N_11632,N_9590);
and U14963 (N_14963,N_10796,N_10119);
nand U14964 (N_14964,N_10662,N_11671);
or U14965 (N_14965,N_10830,N_11319);
or U14966 (N_14966,N_9447,N_10833);
or U14967 (N_14967,N_11383,N_10906);
xor U14968 (N_14968,N_10111,N_10823);
nor U14969 (N_14969,N_11509,N_10114);
nor U14970 (N_14970,N_10899,N_9246);
nor U14971 (N_14971,N_10334,N_9184);
or U14972 (N_14972,N_10735,N_11149);
nand U14973 (N_14973,N_10229,N_11905);
or U14974 (N_14974,N_10726,N_10128);
nor U14975 (N_14975,N_9395,N_10258);
or U14976 (N_14976,N_9856,N_11368);
and U14977 (N_14977,N_11131,N_9013);
and U14978 (N_14978,N_10400,N_9990);
nand U14979 (N_14979,N_9628,N_11210);
nor U14980 (N_14980,N_11714,N_10758);
xnor U14981 (N_14981,N_11659,N_9526);
nor U14982 (N_14982,N_11926,N_11902);
xnor U14983 (N_14983,N_11471,N_9219);
nor U14984 (N_14984,N_11740,N_10232);
and U14985 (N_14985,N_9680,N_9559);
and U14986 (N_14986,N_9188,N_9702);
and U14987 (N_14987,N_11132,N_10259);
xor U14988 (N_14988,N_9797,N_11007);
nor U14989 (N_14989,N_9063,N_9510);
nor U14990 (N_14990,N_10934,N_9782);
xor U14991 (N_14991,N_11073,N_9785);
or U14992 (N_14992,N_9661,N_9977);
or U14993 (N_14993,N_10875,N_9982);
xnor U14994 (N_14994,N_11138,N_9194);
and U14995 (N_14995,N_11796,N_10396);
nand U14996 (N_14996,N_11520,N_9735);
xnor U14997 (N_14997,N_9417,N_11420);
and U14998 (N_14998,N_9187,N_10452);
nand U14999 (N_14999,N_11184,N_10610);
nor UO_0 (O_0,N_14393,N_12145);
nand UO_1 (O_1,N_14538,N_14130);
nor UO_2 (O_2,N_13630,N_14469);
nand UO_3 (O_3,N_13045,N_12804);
xnor UO_4 (O_4,N_12686,N_12822);
and UO_5 (O_5,N_12632,N_13599);
nand UO_6 (O_6,N_12799,N_12338);
nor UO_7 (O_7,N_14265,N_14631);
xor UO_8 (O_8,N_13104,N_13488);
xor UO_9 (O_9,N_14923,N_13881);
nand UO_10 (O_10,N_14616,N_12645);
nand UO_11 (O_11,N_14438,N_12668);
nand UO_12 (O_12,N_13604,N_14384);
nor UO_13 (O_13,N_12718,N_14780);
or UO_14 (O_14,N_14811,N_14871);
nand UO_15 (O_15,N_14793,N_12960);
or UO_16 (O_16,N_14127,N_13213);
or UO_17 (O_17,N_13959,N_13974);
or UO_18 (O_18,N_12448,N_12133);
nand UO_19 (O_19,N_14693,N_13467);
nand UO_20 (O_20,N_13675,N_13149);
nor UO_21 (O_21,N_12655,N_13920);
xnor UO_22 (O_22,N_12923,N_13862);
nor UO_23 (O_23,N_13007,N_13124);
nand UO_24 (O_24,N_12347,N_14574);
nor UO_25 (O_25,N_13473,N_13432);
xor UO_26 (O_26,N_13896,N_12814);
nand UO_27 (O_27,N_14168,N_14266);
nor UO_28 (O_28,N_12545,N_12083);
or UO_29 (O_29,N_14726,N_12281);
and UO_30 (O_30,N_13309,N_12297);
nand UO_31 (O_31,N_14660,N_14097);
or UO_32 (O_32,N_14535,N_13852);
and UO_33 (O_33,N_13736,N_13402);
nor UO_34 (O_34,N_14657,N_12089);
or UO_35 (O_35,N_12303,N_14433);
nand UO_36 (O_36,N_13468,N_14710);
and UO_37 (O_37,N_14861,N_13631);
and UO_38 (O_38,N_12029,N_14490);
xor UO_39 (O_39,N_14475,N_12916);
or UO_40 (O_40,N_12166,N_13368);
nor UO_41 (O_41,N_13747,N_12802);
and UO_42 (O_42,N_12220,N_14706);
or UO_43 (O_43,N_12955,N_13365);
nor UO_44 (O_44,N_14379,N_12383);
xor UO_45 (O_45,N_12865,N_14652);
and UO_46 (O_46,N_14675,N_14319);
and UO_47 (O_47,N_13263,N_14741);
nand UO_48 (O_48,N_14863,N_12940);
nor UO_49 (O_49,N_14397,N_12310);
nor UO_50 (O_50,N_14434,N_13031);
and UO_51 (O_51,N_14594,N_13932);
nand UO_52 (O_52,N_13012,N_13995);
nand UO_53 (O_53,N_13633,N_14640);
nand UO_54 (O_54,N_14872,N_13443);
or UO_55 (O_55,N_14177,N_14653);
or UO_56 (O_56,N_13378,N_13154);
nor UO_57 (O_57,N_12922,N_12333);
xnor UO_58 (O_58,N_13634,N_12816);
nor UO_59 (O_59,N_14483,N_13192);
nor UO_60 (O_60,N_12437,N_14100);
nand UO_61 (O_61,N_14381,N_14910);
nand UO_62 (O_62,N_14610,N_14868);
xor UO_63 (O_63,N_12237,N_13440);
and UO_64 (O_64,N_12409,N_12501);
nor UO_65 (O_65,N_14427,N_13186);
or UO_66 (O_66,N_12439,N_13581);
nand UO_67 (O_67,N_14200,N_14015);
xor UO_68 (O_68,N_13010,N_12336);
nor UO_69 (O_69,N_13724,N_14011);
and UO_70 (O_70,N_12641,N_14961);
xor UO_71 (O_71,N_13891,N_13883);
or UO_72 (O_72,N_12432,N_14738);
nand UO_73 (O_73,N_12877,N_13543);
or UO_74 (O_74,N_14019,N_12987);
nor UO_75 (O_75,N_13827,N_14751);
nand UO_76 (O_76,N_12457,N_12101);
xnor UO_77 (O_77,N_13865,N_14830);
and UO_78 (O_78,N_14807,N_13002);
nor UO_79 (O_79,N_13254,N_14358);
xnor UO_80 (O_80,N_12376,N_13755);
and UO_81 (O_81,N_12359,N_12839);
nand UO_82 (O_82,N_13704,N_14152);
nand UO_83 (O_83,N_13737,N_12837);
and UO_84 (O_84,N_13541,N_13588);
xnor UO_85 (O_85,N_12714,N_13300);
nand UO_86 (O_86,N_12722,N_12984);
or UO_87 (O_87,N_14786,N_13344);
xnor UO_88 (O_88,N_12163,N_14238);
xor UO_89 (O_89,N_12570,N_12765);
nand UO_90 (O_90,N_13572,N_14676);
and UO_91 (O_91,N_13810,N_12709);
and UO_92 (O_92,N_13579,N_12646);
xnor UO_93 (O_93,N_13870,N_14017);
or UO_94 (O_94,N_12526,N_13693);
or UO_95 (O_95,N_14398,N_13076);
nand UO_96 (O_96,N_13683,N_14083);
nand UO_97 (O_97,N_14271,N_12048);
nand UO_98 (O_98,N_13938,N_12241);
nand UO_99 (O_99,N_14138,N_14282);
and UO_100 (O_100,N_14367,N_14905);
nor UO_101 (O_101,N_12497,N_14079);
or UO_102 (O_102,N_14988,N_12047);
nor UO_103 (O_103,N_14092,N_12793);
and UO_104 (O_104,N_13009,N_13127);
nor UO_105 (O_105,N_12650,N_13939);
and UO_106 (O_106,N_14170,N_14355);
nor UO_107 (O_107,N_14175,N_14805);
xnor UO_108 (O_108,N_13113,N_12609);
or UO_109 (O_109,N_13266,N_12482);
or UO_110 (O_110,N_14413,N_13478);
xor UO_111 (O_111,N_13702,N_13105);
nor UO_112 (O_112,N_14553,N_13426);
nor UO_113 (O_113,N_13397,N_12104);
or UO_114 (O_114,N_14783,N_13719);
nand UO_115 (O_115,N_13767,N_13503);
nor UO_116 (O_116,N_12342,N_14982);
nor UO_117 (O_117,N_13350,N_14990);
nand UO_118 (O_118,N_14522,N_12164);
or UO_119 (O_119,N_13484,N_14534);
nor UO_120 (O_120,N_12546,N_13976);
xor UO_121 (O_121,N_13385,N_13661);
nor UO_122 (O_122,N_12531,N_13603);
or UO_123 (O_123,N_14328,N_12943);
and UO_124 (O_124,N_13398,N_14400);
xnor UO_125 (O_125,N_13394,N_12597);
or UO_126 (O_126,N_14135,N_12337);
nand UO_127 (O_127,N_14629,N_14246);
or UO_128 (O_128,N_13132,N_13744);
nand UO_129 (O_129,N_12175,N_12659);
xnor UO_130 (O_130,N_14778,N_12543);
or UO_131 (O_131,N_13612,N_13008);
nor UO_132 (O_132,N_12446,N_13898);
and UO_133 (O_133,N_12717,N_14554);
or UO_134 (O_134,N_14188,N_13003);
or UO_135 (O_135,N_13166,N_12433);
nand UO_136 (O_136,N_14006,N_12422);
nand UO_137 (O_137,N_12548,N_13274);
nand UO_138 (O_138,N_12130,N_14699);
nor UO_139 (O_139,N_12615,N_13799);
or UO_140 (O_140,N_14440,N_12592);
nor UO_141 (O_141,N_14387,N_13487);
and UO_142 (O_142,N_13297,N_13109);
nand UO_143 (O_143,N_14263,N_12013);
nand UO_144 (O_144,N_12859,N_13751);
or UO_145 (O_145,N_14285,N_13598);
xor UO_146 (O_146,N_12040,N_12680);
or UO_147 (O_147,N_14161,N_13268);
nand UO_148 (O_148,N_13221,N_13700);
xnor UO_149 (O_149,N_13392,N_13319);
nand UO_150 (O_150,N_12348,N_12560);
or UO_151 (O_151,N_14678,N_12181);
and UO_152 (O_152,N_14069,N_12456);
or UO_153 (O_153,N_14145,N_13670);
or UO_154 (O_154,N_13427,N_14312);
nand UO_155 (O_155,N_13998,N_13231);
nand UO_156 (O_156,N_14442,N_13051);
nand UO_157 (O_157,N_14211,N_13270);
or UO_158 (O_158,N_12774,N_14583);
nand UO_159 (O_159,N_13387,N_14102);
and UO_160 (O_160,N_14300,N_12931);
nand UO_161 (O_161,N_14541,N_14792);
xnor UO_162 (O_162,N_14421,N_12840);
and UO_163 (O_163,N_13228,N_14112);
or UO_164 (O_164,N_13449,N_13840);
and UO_165 (O_165,N_14273,N_13514);
nor UO_166 (O_166,N_12605,N_13046);
xor UO_167 (O_167,N_14390,N_13899);
nand UO_168 (O_168,N_12519,N_12986);
nand UO_169 (O_169,N_12229,N_14620);
xnor UO_170 (O_170,N_12569,N_12852);
xor UO_171 (O_171,N_12999,N_14096);
nand UO_172 (O_172,N_14194,N_13438);
nor UO_173 (O_173,N_12428,N_12478);
nor UO_174 (O_174,N_14321,N_12801);
xnor UO_175 (O_175,N_12584,N_14885);
and UO_176 (O_176,N_13321,N_13346);
xnor UO_177 (O_177,N_13477,N_13894);
nand UO_178 (O_178,N_12851,N_12387);
nand UO_179 (O_179,N_12442,N_12735);
nand UO_180 (O_180,N_13022,N_14545);
nand UO_181 (O_181,N_12624,N_14494);
nor UO_182 (O_182,N_14394,N_14153);
and UO_183 (O_183,N_13617,N_14325);
and UO_184 (O_184,N_14997,N_12990);
nand UO_185 (O_185,N_13320,N_14409);
nor UO_186 (O_186,N_12065,N_13660);
and UO_187 (O_187,N_14721,N_12012);
nor UO_188 (O_188,N_13262,N_13897);
or UO_189 (O_189,N_14295,N_13963);
or UO_190 (O_190,N_12156,N_13622);
nand UO_191 (O_191,N_12716,N_12466);
nand UO_192 (O_192,N_14163,N_12092);
or UO_193 (O_193,N_13406,N_13817);
xor UO_194 (O_194,N_13833,N_13712);
xor UO_195 (O_195,N_13367,N_12567);
and UO_196 (O_196,N_14318,N_14294);
nor UO_197 (O_197,N_14301,N_13929);
or UO_198 (O_198,N_12389,N_14256);
nor UO_199 (O_199,N_13966,N_12614);
nand UO_200 (O_200,N_14895,N_12918);
nand UO_201 (O_201,N_12970,N_12664);
xnor UO_202 (O_202,N_14497,N_14424);
nor UO_203 (O_203,N_13925,N_12232);
or UO_204 (O_204,N_12557,N_12746);
and UO_205 (O_205,N_13716,N_12964);
or UO_206 (O_206,N_14189,N_14980);
and UO_207 (O_207,N_14985,N_13510);
xor UO_208 (O_208,N_14316,N_12926);
xor UO_209 (O_209,N_13548,N_14991);
xor UO_210 (O_210,N_12407,N_14502);
xor UO_211 (O_211,N_13429,N_12930);
xnor UO_212 (O_212,N_13190,N_12425);
or UO_213 (O_213,N_13874,N_13323);
nor UO_214 (O_214,N_12062,N_14231);
nor UO_215 (O_215,N_14904,N_14503);
nand UO_216 (O_216,N_13928,N_14129);
nor UO_217 (O_217,N_14280,N_12262);
or UO_218 (O_218,N_12351,N_12553);
nand UO_219 (O_219,N_14436,N_12893);
nor UO_220 (O_220,N_12087,N_14714);
nand UO_221 (O_221,N_14853,N_14873);
nor UO_222 (O_222,N_14713,N_12134);
and UO_223 (O_223,N_14758,N_14234);
xor UO_224 (O_224,N_14925,N_13695);
xnor UO_225 (O_225,N_12973,N_13999);
and UO_226 (O_226,N_14578,N_12042);
nor UO_227 (O_227,N_14731,N_12275);
or UO_228 (O_228,N_14334,N_12451);
nand UO_229 (O_229,N_14186,N_13841);
or UO_230 (O_230,N_12972,N_14378);
nand UO_231 (O_231,N_13033,N_14979);
xor UO_232 (O_232,N_13260,N_14917);
nor UO_233 (O_233,N_14255,N_14643);
nor UO_234 (O_234,N_12537,N_14812);
and UO_235 (O_235,N_14298,N_13259);
nand UO_236 (O_236,N_13778,N_14766);
and UO_237 (O_237,N_14317,N_12218);
xnor UO_238 (O_238,N_12654,N_13194);
nand UO_239 (O_239,N_13222,N_12139);
or UO_240 (O_240,N_12097,N_13439);
xor UO_241 (O_241,N_13979,N_14169);
nand UO_242 (O_242,N_12658,N_13621);
or UO_243 (O_243,N_12663,N_13084);
nand UO_244 (O_244,N_14728,N_14945);
nand UO_245 (O_245,N_14279,N_13129);
and UO_246 (O_246,N_14665,N_12544);
xor UO_247 (O_247,N_13591,N_12606);
or UO_248 (O_248,N_12226,N_13685);
nand UO_249 (O_249,N_12132,N_14411);
xnor UO_250 (O_250,N_12630,N_13561);
nand UO_251 (O_251,N_12678,N_12721);
nand UO_252 (O_252,N_14612,N_12200);
nor UO_253 (O_253,N_12054,N_12881);
xor UO_254 (O_254,N_12011,N_12094);
nand UO_255 (O_255,N_13264,N_12240);
and UO_256 (O_256,N_14897,N_14426);
xnor UO_257 (O_257,N_13812,N_14582);
xor UO_258 (O_258,N_12810,N_14500);
xnor UO_259 (O_259,N_13821,N_14829);
xor UO_260 (O_260,N_13411,N_12071);
or UO_261 (O_261,N_13533,N_12364);
xnor UO_262 (O_262,N_12749,N_14386);
and UO_263 (O_263,N_12265,N_12915);
nand UO_264 (O_264,N_14195,N_14484);
nor UO_265 (O_265,N_12397,N_14599);
nand UO_266 (O_266,N_14581,N_12707);
nor UO_267 (O_267,N_12627,N_13142);
or UO_268 (O_268,N_12800,N_12935);
nand UO_269 (O_269,N_13613,N_13880);
and UO_270 (O_270,N_14226,N_13752);
nand UO_271 (O_271,N_13066,N_13527);
xnor UO_272 (O_272,N_12136,N_14931);
xor UO_273 (O_273,N_13493,N_14906);
xor UO_274 (O_274,N_14790,N_13182);
nor UO_275 (O_275,N_14313,N_13994);
xnor UO_276 (O_276,N_13990,N_12157);
nor UO_277 (O_277,N_14042,N_13667);
xnor UO_278 (O_278,N_12014,N_14405);
nand UO_279 (O_279,N_12015,N_12622);
or UO_280 (O_280,N_12669,N_13694);
xnor UO_281 (O_281,N_12248,N_14528);
nand UO_282 (O_282,N_13566,N_13520);
xnor UO_283 (O_283,N_13483,N_13526);
nand UO_284 (O_284,N_13909,N_12667);
or UO_285 (O_285,N_14128,N_12920);
nand UO_286 (O_286,N_14047,N_13506);
and UO_287 (O_287,N_13576,N_14477);
nor UO_288 (O_288,N_14619,N_14890);
nor UO_289 (O_289,N_12599,N_14929);
and UO_290 (O_290,N_14350,N_13472);
and UO_291 (O_291,N_13969,N_13011);
or UO_292 (O_292,N_12562,N_12171);
nand UO_293 (O_293,N_14674,N_13734);
and UO_294 (O_294,N_14399,N_14349);
and UO_295 (O_295,N_14344,N_12867);
and UO_296 (O_296,N_12533,N_13644);
nor UO_297 (O_297,N_13057,N_13814);
xor UO_298 (O_298,N_12891,N_13546);
nor UO_299 (O_299,N_13216,N_14134);
xor UO_300 (O_300,N_12400,N_14037);
nand UO_301 (O_301,N_14351,N_12203);
nor UO_302 (O_302,N_14272,N_14966);
nor UO_303 (O_303,N_13442,N_13165);
nor UO_304 (O_304,N_12027,N_14289);
or UO_305 (O_305,N_13403,N_12514);
nor UO_306 (O_306,N_14839,N_13768);
nor UO_307 (O_307,N_13082,N_12408);
nand UO_308 (O_308,N_13304,N_14458);
nand UO_309 (O_309,N_14600,N_13653);
and UO_310 (O_310,N_14197,N_14977);
and UO_311 (O_311,N_13509,N_13791);
nand UO_312 (O_312,N_13404,N_14156);
or UO_313 (O_313,N_14382,N_12561);
nand UO_314 (O_314,N_13048,N_13776);
and UO_315 (O_315,N_14471,N_12410);
nor UO_316 (O_316,N_12957,N_14029);
nor UO_317 (O_317,N_14401,N_14291);
nand UO_318 (O_318,N_14315,N_14566);
nand UO_319 (O_319,N_14043,N_14605);
nand UO_320 (O_320,N_13199,N_13416);
xnor UO_321 (O_321,N_13957,N_14539);
nand UO_322 (O_322,N_13239,N_12170);
nor UO_323 (O_323,N_12813,N_13948);
and UO_324 (O_324,N_13041,N_12204);
xor UO_325 (O_325,N_12868,N_14335);
and UO_326 (O_326,N_13339,N_14457);
and UO_327 (O_327,N_12302,N_12512);
and UO_328 (O_328,N_13972,N_14377);
and UO_329 (O_329,N_13749,N_13762);
or UO_330 (O_330,N_12496,N_13686);
xor UO_331 (O_331,N_14274,N_14067);
or UO_332 (O_332,N_13656,N_12788);
and UO_333 (O_333,N_12998,N_14396);
nor UO_334 (O_334,N_12515,N_12063);
nor UO_335 (O_335,N_12435,N_13708);
and UO_336 (O_336,N_14008,N_13600);
or UO_337 (O_337,N_13793,N_12480);
nor UO_338 (O_338,N_14235,N_12450);
or UO_339 (O_339,N_13530,N_12023);
or UO_340 (O_340,N_13121,N_12230);
or UO_341 (O_341,N_14488,N_12454);
and UO_342 (O_342,N_12264,N_13682);
xor UO_343 (O_343,N_12616,N_12542);
nor UO_344 (O_344,N_14821,N_14144);
xor UO_345 (O_345,N_13914,N_14647);
nor UO_346 (O_346,N_14088,N_13459);
and UO_347 (O_347,N_12197,N_12684);
xor UO_348 (O_348,N_12950,N_13742);
and UO_349 (O_349,N_12811,N_12843);
and UO_350 (O_350,N_12574,N_13445);
and UO_351 (O_351,N_13373,N_12601);
xnor UO_352 (O_352,N_14262,N_14455);
or UO_353 (O_353,N_14199,N_14824);
xor UO_354 (O_354,N_13607,N_13931);
or UO_355 (O_355,N_12997,N_13872);
nor UO_356 (O_356,N_12559,N_14408);
and UO_357 (O_357,N_12385,N_13668);
nand UO_358 (O_358,N_12008,N_14115);
nor UO_359 (O_359,N_13207,N_12963);
or UO_360 (O_360,N_12739,N_12805);
nand UO_361 (O_361,N_13563,N_13180);
nor UO_362 (O_362,N_13804,N_13352);
nor UO_363 (O_363,N_14989,N_14942);
nand UO_364 (O_364,N_13725,N_13940);
and UO_365 (O_365,N_13244,N_13987);
nor UO_366 (O_366,N_13962,N_12331);
and UO_367 (O_367,N_14076,N_14908);
xnor UO_368 (O_368,N_14712,N_14843);
xnor UO_369 (O_369,N_13981,N_14504);
nor UO_370 (O_370,N_14984,N_12625);
nor UO_371 (O_371,N_12866,N_14449);
nand UO_372 (O_372,N_12864,N_13291);
or UO_373 (O_373,N_14846,N_13044);
nand UO_374 (O_374,N_13669,N_14532);
nor UO_375 (O_375,N_14834,N_12789);
nand UO_376 (O_376,N_13167,N_12039);
nand UO_377 (O_377,N_14700,N_14040);
nand UO_378 (O_378,N_14743,N_12534);
and UO_379 (O_379,N_14463,N_13281);
and UO_380 (O_380,N_13726,N_12234);
and UO_381 (O_381,N_14412,N_12118);
nand UO_382 (O_382,N_12880,N_12556);
and UO_383 (O_383,N_12377,N_12731);
nor UO_384 (O_384,N_12135,N_14452);
nand UO_385 (O_385,N_12072,N_12100);
nor UO_386 (O_386,N_12776,N_13771);
nand UO_387 (O_387,N_14555,N_12242);
xnor UO_388 (O_388,N_12193,N_14810);
and UO_389 (O_389,N_13508,N_13265);
and UO_390 (O_390,N_12892,N_14462);
nand UO_391 (O_391,N_14509,N_14607);
or UO_392 (O_392,N_12525,N_13955);
or UO_393 (O_393,N_13413,N_13623);
nand UO_394 (O_394,N_12443,N_12890);
or UO_395 (O_395,N_12563,N_14866);
xnor UO_396 (O_396,N_13795,N_12849);
nand UO_397 (O_397,N_12607,N_14320);
xnor UO_398 (O_398,N_13900,N_12883);
nor UO_399 (O_399,N_13678,N_14962);
or UO_400 (O_400,N_12452,N_12492);
and UO_401 (O_401,N_13727,N_13333);
xnor UO_402 (O_402,N_13032,N_14116);
xnor UO_403 (O_403,N_14587,N_14951);
nand UO_404 (O_404,N_14891,N_12856);
nand UO_405 (O_405,N_14656,N_14995);
or UO_406 (O_406,N_12142,N_12225);
and UO_407 (O_407,N_13240,N_12058);
and UO_408 (O_408,N_14617,N_13887);
and UO_409 (O_409,N_13504,N_13460);
xnor UO_410 (O_410,N_12182,N_14027);
nor UO_411 (O_411,N_13172,N_14330);
or UO_412 (O_412,N_12540,N_12921);
xnor UO_413 (O_413,N_12976,N_13071);
and UO_414 (O_414,N_12770,N_12585);
nand UO_415 (O_415,N_12114,N_12979);
or UO_416 (O_416,N_13131,N_12413);
nand UO_417 (O_417,N_13220,N_14841);
nor UO_418 (O_418,N_12794,N_13362);
nor UO_419 (O_419,N_14292,N_13829);
and UO_420 (O_420,N_12099,N_14403);
nand UO_421 (O_421,N_12939,N_13024);
xnor UO_422 (O_422,N_13096,N_13619);
and UO_423 (O_423,N_12313,N_13334);
nand UO_424 (O_424,N_14930,N_12860);
nor UO_425 (O_425,N_14303,N_12300);
nor UO_426 (O_426,N_13692,N_12024);
xnor UO_427 (O_427,N_12745,N_13209);
or UO_428 (O_428,N_14789,N_13068);
xnor UO_429 (O_429,N_14150,N_12291);
or UO_430 (O_430,N_13494,N_14340);
nand UO_431 (O_431,N_12284,N_13673);
and UO_432 (O_432,N_14049,N_12199);
and UO_433 (O_433,N_13597,N_13278);
xnor UO_434 (O_434,N_12855,N_13884);
nor UO_435 (O_435,N_12706,N_13707);
and UO_436 (O_436,N_13711,N_12373);
or UO_437 (O_437,N_13714,N_13913);
nor UO_438 (O_438,N_14091,N_14418);
xor UO_439 (O_439,N_12110,N_12418);
nand UO_440 (O_440,N_13237,N_12894);
and UO_441 (O_441,N_13189,N_12677);
or UO_442 (O_442,N_14098,N_13163);
xnor UO_443 (O_443,N_14219,N_12080);
or UO_444 (O_444,N_14921,N_13087);
nand UO_445 (O_445,N_12761,N_12445);
or UO_446 (O_446,N_12289,N_12060);
xnor UO_447 (O_447,N_14852,N_12572);
nor UO_448 (O_448,N_12500,N_13836);
and UO_449 (O_449,N_13075,N_12978);
and UO_450 (O_450,N_14536,N_13395);
and UO_451 (O_451,N_14972,N_14190);
xor UO_452 (O_452,N_14080,N_14870);
xnor UO_453 (O_453,N_13890,N_13978);
nand UO_454 (O_454,N_12869,N_13060);
nand UO_455 (O_455,N_14252,N_13792);
or UO_456 (O_456,N_12103,N_12633);
xor UO_457 (O_457,N_13956,N_14898);
nand UO_458 (O_458,N_14845,N_12688);
and UO_459 (O_459,N_14109,N_14139);
nor UO_460 (O_460,N_14529,N_13232);
or UO_461 (O_461,N_13141,N_13851);
nand UO_462 (O_462,N_13037,N_14548);
and UO_463 (O_463,N_13536,N_13754);
and UO_464 (O_464,N_12028,N_12223);
xnor UO_465 (O_465,N_13696,N_13335);
nand UO_466 (O_466,N_14470,N_13122);
nand UO_467 (O_467,N_12854,N_12649);
xor UO_468 (O_468,N_12812,N_14896);
and UO_469 (O_469,N_14105,N_12549);
and UO_470 (O_470,N_13951,N_12712);
nand UO_471 (O_471,N_12273,N_14004);
and UO_472 (O_472,N_13625,N_14205);
xnor UO_473 (O_473,N_14874,N_13521);
or UO_474 (O_474,N_14228,N_14697);
and UO_475 (O_475,N_12090,N_14402);
xnor UO_476 (O_476,N_12243,N_14798);
xor UO_477 (O_477,N_13203,N_12610);
and UO_478 (O_478,N_13174,N_13377);
nor UO_479 (O_479,N_12910,N_12460);
nand UO_480 (O_480,N_12876,N_14276);
xor UO_481 (O_481,N_13433,N_14530);
or UO_482 (O_482,N_12644,N_12259);
xnor UO_483 (O_483,N_12186,N_14165);
or UO_484 (O_484,N_13583,N_12681);
xor UO_485 (O_485,N_13168,N_12470);
nor UO_486 (O_486,N_12954,N_12696);
or UO_487 (O_487,N_12844,N_12536);
nand UO_488 (O_488,N_12675,N_14533);
and UO_489 (O_489,N_12326,N_13544);
or UO_490 (O_490,N_14887,N_14865);
nand UO_491 (O_491,N_14293,N_14767);
and UO_492 (O_492,N_13162,N_14201);
nor UO_493 (O_493,N_13691,N_13567);
and UO_494 (O_494,N_14425,N_14137);
nand UO_495 (O_495,N_14309,N_13225);
or UO_496 (O_496,N_12272,N_12151);
or UO_497 (O_497,N_14095,N_12059);
and UO_498 (O_498,N_14692,N_12577);
xor UO_499 (O_499,N_14249,N_12825);
nor UO_500 (O_500,N_14359,N_14847);
nor UO_501 (O_501,N_14270,N_12917);
nor UO_502 (O_502,N_14007,N_13481);
nor UO_503 (O_503,N_12693,N_13743);
or UO_504 (O_504,N_13906,N_13205);
nor UO_505 (O_505,N_12538,N_14577);
and UO_506 (O_506,N_14341,N_14597);
and UO_507 (O_507,N_12141,N_14924);
or UO_508 (O_508,N_14453,N_12356);
xor UO_509 (O_509,N_14021,N_14524);
nand UO_510 (O_510,N_13425,N_13126);
xor UO_511 (O_511,N_14407,N_14311);
nor UO_512 (O_512,N_14760,N_13482);
nand UO_513 (O_513,N_14590,N_13034);
and UO_514 (O_514,N_13242,N_14523);
or UO_515 (O_515,N_14779,N_14644);
nand UO_516 (O_516,N_14446,N_14071);
nor UO_517 (O_517,N_14927,N_12415);
nor UO_518 (O_518,N_12755,N_12623);
nor UO_519 (O_519,N_12091,N_14033);
and UO_520 (O_520,N_13992,N_14207);
or UO_521 (O_521,N_13086,N_13293);
or UO_522 (O_522,N_14247,N_13844);
nand UO_523 (O_523,N_14243,N_12473);
xor UO_524 (O_524,N_13164,N_12494);
nand UO_525 (O_525,N_12513,N_12929);
and UO_526 (O_526,N_13434,N_12098);
nor UO_527 (O_527,N_14915,N_13973);
nand UO_528 (O_528,N_13364,N_14869);
or UO_529 (O_529,N_14264,N_14218);
xnor UO_530 (O_530,N_13454,N_13666);
nand UO_531 (O_531,N_12991,N_14456);
nand UO_532 (O_532,N_14467,N_12944);
nand UO_533 (O_533,N_13813,N_14167);
or UO_534 (O_534,N_14118,N_13092);
nand UO_535 (O_535,N_13230,N_13638);
nand UO_536 (O_536,N_13098,N_14748);
nor UO_537 (O_537,N_13206,N_12255);
xor UO_538 (O_538,N_12870,N_12049);
nor UO_539 (O_539,N_12613,N_13272);
xor UO_540 (O_540,N_12682,N_13571);
nor UO_541 (O_541,N_13933,N_13765);
nand UO_542 (O_542,N_14461,N_14451);
or UO_543 (O_543,N_14975,N_12033);
xnor UO_544 (O_544,N_13447,N_13238);
nor UO_545 (O_545,N_14525,N_12018);
nand UO_546 (O_546,N_13441,N_12873);
and UO_547 (O_547,N_14907,N_14448);
and UO_548 (O_548,N_12612,N_13001);
xor UO_549 (O_549,N_14229,N_13722);
xnor UO_550 (O_550,N_13780,N_14416);
or UO_551 (O_551,N_13295,N_14063);
xnor UO_552 (O_552,N_14310,N_13436);
or UO_553 (O_553,N_13681,N_14698);
nor UO_554 (O_554,N_14663,N_13689);
xor UO_555 (O_555,N_14928,N_14441);
or UO_556 (O_556,N_13279,N_13059);
nor UO_557 (O_557,N_13296,N_13179);
nor UO_558 (O_558,N_12334,N_12581);
or UO_559 (O_559,N_13642,N_13147);
nand UO_560 (O_560,N_12838,N_13892);
nor UO_561 (O_561,N_12155,N_12863);
nor UO_562 (O_562,N_12330,N_12848);
and UO_563 (O_563,N_14969,N_12784);
xor UO_564 (O_564,N_12143,N_13620);
nor UO_565 (O_565,N_13713,N_12455);
and UO_566 (O_566,N_13038,N_12490);
or UO_567 (O_567,N_13358,N_12252);
and UO_568 (O_568,N_14217,N_12552);
xor UO_569 (O_569,N_14957,N_13655);
nor UO_570 (O_570,N_13953,N_14181);
and UO_571 (O_571,N_13986,N_14081);
nor UO_572 (O_572,N_12932,N_12207);
xor UO_573 (O_573,N_13537,N_13340);
or UO_574 (O_574,N_12343,N_14099);
nor UO_575 (O_575,N_14034,N_12245);
xor UO_576 (O_576,N_13677,N_14077);
nor UO_577 (O_577,N_13945,N_13039);
nor UO_578 (O_578,N_14797,N_12394);
nand UO_579 (O_579,N_12046,N_14662);
nor UO_580 (O_580,N_12176,N_13097);
or UO_581 (O_581,N_12057,N_12412);
and UO_582 (O_582,N_14518,N_14782);
xnor UO_583 (O_583,N_13155,N_14689);
nor UO_584 (O_584,N_14571,N_14588);
and UO_585 (O_585,N_12416,N_12591);
xnor UO_586 (O_586,N_12959,N_13006);
nand UO_587 (O_587,N_14479,N_13025);
or UO_588 (O_588,N_14711,N_14827);
or UO_589 (O_589,N_14749,N_14764);
nand UO_590 (O_590,N_12423,N_14762);
and UO_591 (O_591,N_12589,N_14375);
nor UO_592 (O_592,N_14914,N_13569);
nor UO_593 (O_593,N_13464,N_13964);
xnor UO_594 (O_594,N_12982,N_12773);
or UO_595 (O_595,N_13028,N_13376);
xor UO_596 (O_596,N_14608,N_12202);
or UO_597 (O_597,N_14388,N_12088);
and UO_598 (O_598,N_12192,N_13705);
xor UO_599 (O_599,N_12766,N_13366);
xnor UO_600 (O_600,N_14550,N_14030);
and UO_601 (O_601,N_13252,N_14709);
and UO_602 (O_602,N_14806,N_12493);
or UO_603 (O_603,N_12723,N_14720);
and UO_604 (O_604,N_12580,N_14283);
nor UO_605 (O_605,N_13553,N_13201);
nand UO_606 (O_606,N_14232,N_12983);
and UO_607 (O_607,N_14489,N_14090);
nand UO_608 (O_608,N_13699,N_12578);
or UO_609 (O_609,N_13636,N_12661);
nand UO_610 (O_610,N_13868,N_13405);
xor UO_611 (O_611,N_13056,N_14992);
nand UO_612 (O_612,N_14552,N_14860);
nand UO_613 (O_613,N_13256,N_13187);
and UO_614 (O_614,N_13674,N_14058);
and UO_615 (O_615,N_12551,N_12149);
and UO_616 (O_616,N_14024,N_13349);
nand UO_617 (O_617,N_13214,N_13233);
nor UO_618 (O_618,N_12674,N_13107);
xnor UO_619 (O_619,N_13106,N_12951);
xor UO_620 (O_620,N_12969,N_14196);
or UO_621 (O_621,N_14346,N_14822);
nand UO_622 (O_622,N_12498,N_12320);
nand UO_623 (O_623,N_13807,N_14593);
nor UO_624 (O_624,N_14075,N_13390);
and UO_625 (O_625,N_13605,N_13657);
xnor UO_626 (O_626,N_13875,N_12108);
or UO_627 (O_627,N_12701,N_12477);
or UO_628 (O_628,N_12586,N_14848);
xor UO_629 (O_629,N_13248,N_12508);
xnor UO_630 (O_630,N_12558,N_13885);
or UO_631 (O_631,N_14254,N_14682);
and UO_632 (O_632,N_14185,N_12958);
nand UO_633 (O_633,N_12127,N_12732);
xor UO_634 (O_634,N_14624,N_12109);
nand UO_635 (O_635,N_14825,N_14093);
nand UO_636 (O_636,N_13080,N_13159);
and UO_637 (O_637,N_12692,N_13253);
nor UO_638 (O_638,N_12231,N_13257);
or UO_639 (O_639,N_12535,N_14973);
nor UO_640 (O_640,N_13361,N_13181);
and UO_641 (O_641,N_12520,N_13798);
xnor UO_642 (O_642,N_13800,N_13301);
nand UO_643 (O_643,N_13997,N_14983);
or UO_644 (O_644,N_14670,N_14038);
or UO_645 (O_645,N_14473,N_13921);
xnor UO_646 (O_646,N_13735,N_12640);
xor UO_647 (O_647,N_14703,N_12263);
xnor UO_648 (O_648,N_13314,N_13169);
nor UO_649 (O_649,N_13730,N_13299);
xnor UO_650 (O_650,N_12938,N_14078);
or UO_651 (O_651,N_12541,N_14801);
nor UO_652 (O_652,N_14986,N_14770);
nor UO_653 (O_653,N_12213,N_12122);
or UO_654 (O_654,N_12790,N_13505);
nand UO_655 (O_655,N_12847,N_14596);
nand UO_656 (O_656,N_14968,N_13781);
and UO_657 (O_657,N_12711,N_14369);
or UO_658 (O_658,N_13061,N_14506);
nor UO_659 (O_659,N_14936,N_14362);
and UO_660 (O_660,N_13152,N_13489);
nand UO_661 (O_661,N_14661,N_13849);
and UO_662 (O_662,N_13801,N_13977);
xnor UO_663 (O_663,N_12296,N_13383);
or UO_664 (O_664,N_13063,N_12222);
nor UO_665 (O_665,N_13280,N_13784);
or UO_666 (O_666,N_13360,N_14820);
or UO_667 (O_667,N_12462,N_14543);
xor UO_668 (O_668,N_12523,N_13593);
or UO_669 (O_669,N_14208,N_13641);
xor UO_670 (O_670,N_12566,N_12250);
nor UO_671 (O_671,N_13474,N_14883);
nor UO_672 (O_672,N_12573,N_14242);
xor UO_673 (O_673,N_13235,N_12074);
nand UO_674 (O_674,N_12846,N_12952);
and UO_675 (O_675,N_13284,N_13115);
nor UO_676 (O_676,N_13927,N_12635);
nand UO_677 (O_677,N_12173,N_12271);
or UO_678 (O_678,N_12832,N_13176);
or UO_679 (O_679,N_13942,N_12936);
xor UO_680 (O_680,N_13717,N_12705);
or UO_681 (O_681,N_14752,N_14389);
xnor UO_682 (O_682,N_14556,N_14939);
nand UO_683 (O_683,N_14251,N_12321);
or UO_684 (O_684,N_13258,N_14512);
nand UO_685 (O_685,N_13329,N_12595);
or UO_686 (O_686,N_13355,N_13845);
nand UO_687 (O_687,N_13069,N_14673);
xor UO_688 (O_688,N_14336,N_12366);
or UO_689 (O_689,N_14066,N_12323);
nand UO_690 (O_690,N_14203,N_14955);
nand UO_691 (O_691,N_13351,N_12238);
nand UO_692 (O_692,N_12777,N_13282);
xnor UO_693 (O_693,N_13095,N_12153);
nor UO_694 (O_694,N_14472,N_13595);
nor UO_695 (O_695,N_14338,N_13889);
and UO_696 (O_696,N_12227,N_14106);
or UO_697 (O_697,N_12665,N_13050);
xor UO_698 (O_698,N_14974,N_14601);
xor UO_699 (O_699,N_14250,N_13837);
nor UO_700 (O_700,N_12025,N_14443);
nand UO_701 (O_701,N_14591,N_13229);
and UO_702 (O_702,N_14326,N_14499);
nor UO_703 (O_703,N_12115,N_14892);
or UO_704 (O_704,N_12760,N_14410);
xor UO_705 (O_705,N_13480,N_12956);
xnor UO_706 (O_706,N_14956,N_13965);
nand UO_707 (O_707,N_12003,N_12386);
or UO_708 (O_708,N_12928,N_13277);
and UO_709 (O_709,N_14788,N_14278);
xnor UO_710 (O_710,N_13227,N_13135);
nand UO_711 (O_711,N_13306,N_12905);
xnor UO_712 (O_712,N_12140,N_14753);
or UO_713 (O_713,N_13843,N_13511);
or UO_714 (O_714,N_12345,N_12683);
or UO_715 (O_715,N_12704,N_13573);
or UO_716 (O_716,N_12634,N_12685);
or UO_717 (O_717,N_13200,N_14772);
xor UO_718 (O_718,N_12842,N_14178);
nor UO_719 (O_719,N_12128,N_14646);
or UO_720 (O_720,N_14561,N_14391);
nand UO_721 (O_721,N_14052,N_12638);
nand UO_722 (O_722,N_13557,N_13241);
nor UO_723 (O_723,N_13594,N_12603);
xnor UO_724 (O_724,N_14184,N_13303);
nor UO_725 (O_725,N_14193,N_12362);
or UO_726 (O_726,N_13609,N_12555);
and UO_727 (O_727,N_12524,N_14304);
nor UO_728 (O_728,N_13523,N_12628);
nand UO_729 (O_729,N_14513,N_12438);
xor UO_730 (O_730,N_14916,N_12381);
nand UO_731 (O_731,N_13728,N_12069);
nor UO_732 (O_732,N_12319,N_14836);
nand UO_733 (O_733,N_13822,N_12393);
nand UO_734 (O_734,N_14212,N_13937);
and UO_735 (O_735,N_12215,N_12474);
nor UO_736 (O_736,N_14630,N_14542);
nor UO_737 (O_737,N_12352,N_13029);
or UO_738 (O_738,N_14108,N_12210);
or UO_739 (O_739,N_12301,N_13458);
and UO_740 (O_740,N_14649,N_14147);
xnor UO_741 (O_741,N_13869,N_14745);
xnor UO_742 (O_742,N_12835,N_12224);
and UO_743 (O_743,N_12311,N_14435);
and UO_744 (O_744,N_14527,N_13400);
or UO_745 (O_745,N_13067,N_12401);
xor UO_746 (O_746,N_14671,N_13302);
and UO_747 (O_747,N_13662,N_12949);
xor UO_748 (O_748,N_13902,N_14819);
xnor UO_749 (O_749,N_13457,N_12499);
xor UO_750 (O_750,N_12823,N_13312);
xnor UO_751 (O_751,N_14919,N_14684);
nand UO_752 (O_752,N_12587,N_12274);
and UO_753 (O_753,N_14946,N_14694);
and UO_754 (O_754,N_13156,N_13420);
nor UO_755 (O_755,N_12710,N_12829);
and UO_756 (O_756,N_12744,N_12036);
nand UO_757 (O_757,N_13359,N_12269);
nor UO_758 (O_758,N_13943,N_14707);
nor UO_759 (O_759,N_12648,N_14893);
nand UO_760 (O_760,N_12741,N_13535);
and UO_761 (O_761,N_14976,N_12747);
nand UO_762 (O_762,N_12022,N_14215);
nand UO_763 (O_763,N_12953,N_12335);
xnor UO_764 (O_764,N_13391,N_12738);
or UO_765 (O_765,N_12602,N_13519);
nand UO_766 (O_766,N_13993,N_13040);
xor UO_767 (O_767,N_14636,N_12249);
nand UO_768 (O_768,N_14383,N_12085);
and UO_769 (O_769,N_13215,N_14965);
or UO_770 (O_770,N_13065,N_14795);
and UO_771 (O_771,N_14632,N_12417);
or UO_772 (O_772,N_13381,N_13552);
xor UO_773 (O_773,N_12371,N_14900);
or UO_774 (O_774,N_13471,N_13842);
nor UO_775 (O_775,N_14679,N_14028);
or UO_776 (O_776,N_13004,N_14241);
and UO_777 (O_777,N_14487,N_12244);
or UO_778 (O_778,N_14450,N_14216);
and UO_779 (O_779,N_13226,N_13175);
and UO_780 (O_780,N_13679,N_13325);
and UO_781 (O_781,N_12734,N_14223);
nand UO_782 (O_782,N_14365,N_13119);
xor UO_783 (O_783,N_13085,N_13125);
and UO_784 (O_784,N_13659,N_12279);
or UO_785 (O_785,N_13018,N_13853);
xor UO_786 (O_786,N_12598,N_12751);
or UO_787 (O_787,N_12152,N_12374);
or UO_788 (O_788,N_12106,N_14911);
or UO_789 (O_789,N_14213,N_13290);
xnor UO_790 (O_790,N_13123,N_13748);
and UO_791 (O_791,N_13815,N_14507);
and UO_792 (O_792,N_14814,N_14062);
nand UO_793 (O_793,N_14800,N_14437);
nor UO_794 (O_794,N_12608,N_12827);
or UO_795 (O_795,N_14909,N_14171);
and UO_796 (O_796,N_14485,N_14005);
and UO_797 (O_797,N_12516,N_12005);
xnor UO_798 (O_798,N_12180,N_13802);
and UO_799 (O_799,N_13102,N_14198);
nor UO_800 (O_800,N_14889,N_13137);
xnor UO_801 (O_801,N_12752,N_14172);
and UO_802 (O_802,N_13564,N_13904);
xnor UO_803 (O_803,N_13545,N_12792);
and UO_804 (O_804,N_13386,N_14025);
nand UO_805 (O_805,N_13372,N_12441);
xnor UO_806 (O_806,N_13565,N_14835);
nor UO_807 (O_807,N_14329,N_13450);
and UO_808 (O_808,N_13327,N_14064);
or UO_809 (O_809,N_13093,N_12817);
xnor UO_810 (O_810,N_13054,N_14950);
and UO_811 (O_811,N_14009,N_13318);
and UO_812 (O_812,N_12031,N_13139);
nor UO_813 (O_813,N_12528,N_14864);
xor UO_814 (O_814,N_12312,N_13435);
nor UO_815 (O_815,N_12160,N_12165);
nor UO_816 (O_816,N_13741,N_14000);
or UO_817 (O_817,N_14056,N_13052);
nand UO_818 (O_818,N_14589,N_12340);
nor UO_819 (O_819,N_12565,N_13342);
nand UO_820 (O_820,N_12901,N_12430);
or UO_821 (O_821,N_12191,N_12576);
and UO_822 (O_822,N_13907,N_14584);
xor UO_823 (O_823,N_12521,N_14306);
nor UO_824 (O_824,N_12299,N_13663);
xor UO_825 (O_825,N_12068,N_13246);
nand UO_826 (O_826,N_12575,N_14142);
xor UO_827 (O_827,N_14771,N_12285);
or UO_828 (O_828,N_12495,N_14938);
nand UO_829 (O_829,N_12082,N_14068);
nor UO_830 (O_830,N_12503,N_12161);
or UO_831 (O_831,N_12298,N_14683);
xnor UO_832 (O_832,N_13100,N_14686);
xor UO_833 (O_833,N_13984,N_13624);
nand UO_834 (O_834,N_14773,N_14559);
or UO_835 (O_835,N_13797,N_14696);
and UO_836 (O_836,N_13103,N_13456);
and UO_837 (O_837,N_12096,N_13157);
or UO_838 (O_838,N_13671,N_13648);
or UO_839 (O_839,N_12502,N_13664);
and UO_840 (O_840,N_12458,N_13158);
and UO_841 (O_841,N_12725,N_14650);
or UO_842 (O_842,N_14659,N_13446);
or UO_843 (O_843,N_14685,N_12174);
nand UO_844 (O_844,N_12070,N_12977);
nand UO_845 (O_845,N_13217,N_12828);
xnor UO_846 (O_846,N_14087,N_13839);
or UO_847 (O_847,N_13049,N_12485);
and UO_848 (O_848,N_14476,N_12332);
xnor UO_849 (O_849,N_14718,N_13160);
nor UO_850 (O_850,N_12305,N_14074);
nor UO_851 (O_851,N_13950,N_12857);
or UO_852 (O_852,N_13861,N_14374);
xor UO_853 (O_853,N_14505,N_14903);
or UO_854 (O_854,N_12898,N_14734);
or UO_855 (O_855,N_14808,N_14514);
xnor UO_856 (O_856,N_13924,N_13408);
xor UO_857 (O_857,N_13701,N_12102);
or UO_858 (O_858,N_14342,N_14417);
or UO_859 (O_859,N_14122,N_12483);
nand UO_860 (O_860,N_13850,N_13211);
xor UO_861 (O_861,N_13418,N_13183);
and UO_862 (O_862,N_12044,N_13047);
and UO_863 (O_863,N_14901,N_14609);
xnor UO_864 (O_864,N_12144,N_12511);
and UO_865 (O_865,N_12737,N_13860);
or UO_866 (O_866,N_14765,N_14716);
and UO_867 (O_867,N_14119,N_14623);
xnor UO_868 (O_868,N_14493,N_13697);
xor UO_869 (O_869,N_12360,N_13785);
nor UO_870 (O_870,N_13687,N_13326);
or UO_871 (O_871,N_13988,N_14680);
or UO_872 (O_872,N_13036,N_12154);
or UO_873 (O_873,N_12506,N_13560);
or UO_874 (O_874,N_12043,N_14776);
xor UO_875 (O_875,N_12185,N_13763);
or UO_876 (O_876,N_13832,N_12257);
or UO_877 (O_877,N_14376,N_14308);
nand UO_878 (O_878,N_12125,N_14740);
nor UO_879 (O_879,N_13072,N_12993);
and UO_880 (O_880,N_13492,N_13534);
and UO_881 (O_881,N_14104,N_12927);
or UO_882 (O_882,N_14002,N_13916);
and UO_883 (O_883,N_14763,N_12995);
xor UO_884 (O_884,N_14227,N_12206);
nand UO_885 (O_885,N_12651,N_12414);
nand UO_886 (O_886,N_13879,N_14658);
or UO_887 (O_887,N_12055,N_13968);
or UO_888 (O_888,N_13575,N_13414);
and UO_889 (O_889,N_12420,N_14875);
and UO_890 (O_890,N_12639,N_12689);
and UO_891 (O_891,N_14691,N_13877);
or UO_892 (O_892,N_14333,N_14645);
or UO_893 (O_893,N_14288,N_14373);
xor UO_894 (O_894,N_13985,N_13542);
and UO_895 (O_895,N_13568,N_13733);
nor UO_896 (O_896,N_13782,N_13089);
or UO_897 (O_897,N_13665,N_12429);
nor UO_898 (O_898,N_13499,N_13601);
nand UO_899 (O_899,N_12626,N_12962);
nand UO_900 (O_900,N_12020,N_13876);
nor UO_901 (O_901,N_14121,N_12779);
or UO_902 (O_902,N_12742,N_13073);
nor UO_903 (O_903,N_14060,N_14041);
xnor UO_904 (O_904,N_13019,N_12214);
or UO_905 (O_905,N_14828,N_13500);
and UO_906 (O_906,N_13580,N_13422);
and UO_907 (O_907,N_14744,N_12937);
nor UO_908 (O_908,N_14486,N_13111);
xor UO_909 (O_909,N_13739,N_14569);
nand UO_910 (O_910,N_13989,N_14781);
and UO_911 (O_911,N_14978,N_14192);
or UO_912 (O_912,N_14182,N_14065);
xnor UO_913 (O_913,N_13777,N_14073);
nand UO_914 (O_914,N_14057,N_13606);
nand UO_915 (O_915,N_13602,N_13292);
or UO_916 (O_916,N_14259,N_13971);
or UO_917 (O_917,N_13703,N_14867);
nor UO_918 (O_918,N_12845,N_14054);
nand UO_919 (O_919,N_12339,N_12084);
nor UO_920 (O_920,N_12369,N_14032);
nor UO_921 (O_921,N_13219,N_12504);
xor UO_922 (O_922,N_14547,N_14563);
or UO_923 (O_923,N_13658,N_12945);
nand UO_924 (O_924,N_13091,N_14173);
nand UO_925 (O_925,N_14361,N_14048);
nand UO_926 (O_926,N_12775,N_14324);
nand UO_927 (O_927,N_14053,N_12889);
nand UO_928 (O_928,N_13549,N_13723);
nand UO_929 (O_929,N_13415,N_14576);
or UO_930 (O_930,N_13064,N_14445);
and UO_931 (O_931,N_14715,N_14204);
nor UO_932 (O_932,N_12254,N_14615);
or UO_933 (O_933,N_12126,N_14785);
or UO_934 (O_934,N_13516,N_13140);
and UO_935 (O_935,N_12489,N_13130);
or UO_936 (O_936,N_13740,N_12329);
or UO_937 (O_937,N_13709,N_13864);
xnor UO_938 (O_938,N_12620,N_14305);
nand UO_939 (O_939,N_13393,N_13960);
nor UO_940 (O_940,N_12906,N_13070);
xnor UO_941 (O_941,N_13324,N_12179);
or UO_942 (O_942,N_14981,N_14347);
xnor UO_943 (O_943,N_14439,N_13173);
nor UO_944 (O_944,N_14708,N_13110);
nand UO_945 (O_945,N_14746,N_13196);
or UO_946 (O_946,N_12720,N_14343);
and UO_947 (O_947,N_12196,N_14086);
and UO_948 (O_948,N_13788,N_14492);
and UO_949 (O_949,N_13461,N_13556);
and UO_950 (O_950,N_13396,N_13469);
xnor UO_951 (O_951,N_13779,N_14478);
and UO_952 (O_952,N_13643,N_14495);
xor UO_953 (O_953,N_13958,N_13847);
and UO_954 (O_954,N_13863,N_14572);
xor UO_955 (O_955,N_12066,N_14613);
and UO_956 (O_956,N_13466,N_14160);
and UO_957 (O_957,N_13455,N_13732);
xor UO_958 (O_958,N_14039,N_13590);
nand UO_959 (O_959,N_13578,N_12826);
xor UO_960 (O_960,N_14117,N_14755);
nand UO_961 (O_961,N_12221,N_14774);
or UO_962 (O_962,N_12507,N_13382);
nor UO_963 (O_963,N_12965,N_14736);
or UO_964 (O_964,N_12286,N_13410);
nand UO_965 (O_965,N_13858,N_14844);
and UO_966 (O_966,N_12396,N_13202);
xnor UO_967 (O_967,N_12947,N_12037);
xor UO_968 (O_968,N_12032,N_12395);
xor UO_969 (O_969,N_13375,N_14816);
xnor UO_970 (O_970,N_12205,N_14158);
and UO_971 (O_971,N_13551,N_12107);
nor UO_972 (O_972,N_13337,N_14690);
xnor UO_973 (O_973,N_12621,N_12925);
or UO_974 (O_974,N_13307,N_14747);
xor UO_975 (O_975,N_12278,N_12975);
and UO_976 (O_976,N_12158,N_12554);
or UO_977 (O_977,N_12809,N_14103);
nand UO_978 (O_978,N_13369,N_12316);
xnor UO_979 (O_979,N_13574,N_12195);
nand UO_980 (O_980,N_14430,N_12600);
or UO_981 (O_981,N_14637,N_14459);
nand UO_982 (O_982,N_13608,N_12933);
or UO_983 (O_983,N_13746,N_13786);
xor UO_984 (O_984,N_14110,N_12687);
xnor UO_985 (O_985,N_14799,N_12836);
nand UO_986 (O_986,N_12948,N_12219);
nand UO_987 (O_987,N_12778,N_12590);
nand UO_988 (O_988,N_14854,N_14918);
nor UO_989 (O_989,N_13629,N_12187);
xnor UO_990 (O_990,N_14468,N_12378);
xnor UO_991 (O_991,N_14858,N_14926);
nor UO_992 (O_992,N_14082,N_12019);
xnor UO_993 (O_993,N_14368,N_14756);
or UO_994 (O_994,N_13363,N_14920);
nor UO_995 (O_995,N_14603,N_12636);
or UO_996 (O_996,N_14415,N_13143);
and UO_997 (O_997,N_13261,N_14406);
nor UO_998 (O_998,N_13627,N_13013);
or UO_999 (O_999,N_12753,N_14001);
nor UO_1000 (O_1000,N_13772,N_12349);
xor UO_1001 (O_1001,N_13090,N_13146);
xnor UO_1002 (O_1002,N_12662,N_14881);
xor UO_1003 (O_1003,N_12188,N_13774);
nor UO_1004 (O_1004,N_12653,N_13271);
and UO_1005 (O_1005,N_13341,N_13559);
nand UO_1006 (O_1006,N_13191,N_13848);
nor UO_1007 (O_1007,N_12787,N_14248);
nor UO_1008 (O_1008,N_12850,N_14592);
and UO_1009 (O_1009,N_13401,N_14940);
nor UO_1010 (O_1010,N_13148,N_14944);
xnor UO_1011 (O_1011,N_12026,N_14954);
nor UO_1012 (O_1012,N_12355,N_14949);
nor UO_1013 (O_1013,N_13347,N_14677);
xor UO_1014 (O_1014,N_12270,N_14287);
nor UO_1015 (O_1015,N_13094,N_14179);
and UO_1016 (O_1016,N_12934,N_14269);
or UO_1017 (O_1017,N_14277,N_14803);
xnor UO_1018 (O_1018,N_14013,N_12253);
or UO_1019 (O_1019,N_14611,N_14432);
nor UO_1020 (O_1020,N_13635,N_14428);
or UO_1021 (O_1021,N_13582,N_14544);
nand UO_1022 (O_1022,N_13626,N_13805);
nor UO_1023 (O_1023,N_13824,N_14284);
and UO_1024 (O_1024,N_14857,N_12292);
or UO_1025 (O_1025,N_12402,N_14567);
nand UO_1026 (O_1026,N_12798,N_12797);
or UO_1027 (O_1027,N_12475,N_12113);
nor UO_1028 (O_1028,N_14557,N_14183);
nor UO_1029 (O_1029,N_12819,N_12772);
xor UO_1030 (O_1030,N_12280,N_12463);
nor UO_1031 (O_1031,N_12002,N_13540);
and UO_1032 (O_1032,N_14761,N_13161);
nor UO_1033 (O_1033,N_14880,N_12261);
or UO_1034 (O_1034,N_14187,N_12831);
or UO_1035 (O_1035,N_13491,N_12246);
nor UO_1036 (O_1036,N_13275,N_14704);
xor UO_1037 (O_1037,N_14520,N_13243);
nor UO_1038 (O_1038,N_14878,N_14526);
nor UO_1039 (O_1039,N_13475,N_12967);
xnor UO_1040 (O_1040,N_14565,N_14510);
and UO_1041 (O_1041,N_12277,N_12518);
nor UO_1042 (O_1042,N_14960,N_14655);
xor UO_1043 (O_1043,N_13554,N_12713);
nor UO_1044 (O_1044,N_12703,N_14061);
and UO_1045 (O_1045,N_14055,N_12833);
nor UO_1046 (O_1046,N_13423,N_13255);
and UO_1047 (O_1047,N_13117,N_13151);
or UO_1048 (O_1048,N_14757,N_13251);
nor UO_1049 (O_1049,N_14072,N_12079);
xor UO_1050 (O_1050,N_13819,N_12403);
or UO_1051 (O_1051,N_13370,N_12444);
xnor UO_1052 (O_1052,N_13133,N_13961);
nand UO_1053 (O_1053,N_14143,N_12440);
nand UO_1054 (O_1054,N_13513,N_14958);
nand UO_1055 (O_1055,N_14546,N_14737);
or UO_1056 (O_1056,N_14964,N_13294);
nand UO_1057 (O_1057,N_13308,N_14260);
and UO_1058 (O_1058,N_12780,N_14996);
or UO_1059 (O_1059,N_13923,N_14862);
nor UO_1060 (O_1060,N_14531,N_12974);
xor UO_1061 (O_1061,N_12064,N_14348);
xor UO_1062 (O_1062,N_14750,N_12167);
nor UO_1063 (O_1063,N_13476,N_14855);
xor UO_1064 (O_1064,N_12902,N_14125);
nand UO_1065 (O_1065,N_13193,N_14667);
and UO_1066 (O_1066,N_14240,N_13371);
nor UO_1067 (O_1067,N_13954,N_14666);
xnor UO_1068 (O_1068,N_14084,N_12009);
and UO_1069 (O_1069,N_12258,N_12771);
nand UO_1070 (O_1070,N_12985,N_13195);
and UO_1071 (O_1071,N_13721,N_14558);
xor UO_1072 (O_1072,N_13592,N_14999);
nor UO_1073 (O_1073,N_12449,N_12617);
or UO_1074 (O_1074,N_14286,N_13354);
or UO_1075 (O_1075,N_12147,N_14654);
xor UO_1076 (O_1076,N_12322,N_12017);
or UO_1077 (O_1077,N_14036,N_14474);
nand UO_1078 (O_1078,N_14133,N_14840);
xor UO_1079 (O_1079,N_13764,N_12426);
nor UO_1080 (O_1080,N_14339,N_14245);
nor UO_1081 (O_1081,N_12233,N_13286);
and UO_1082 (O_1082,N_13081,N_14352);
or UO_1083 (O_1083,N_14354,N_13996);
nor UO_1084 (O_1084,N_12830,N_13794);
nor UO_1085 (O_1085,N_12642,N_12129);
and UO_1086 (O_1086,N_14856,N_14851);
or UO_1087 (O_1087,N_13645,N_14003);
and UO_1088 (O_1088,N_12652,N_14959);
nand UO_1089 (O_1089,N_13688,N_12034);
and UO_1090 (O_1090,N_12700,N_12370);
nand UO_1091 (O_1091,N_12672,N_12368);
and UO_1092 (O_1092,N_13407,N_12530);
nand UO_1093 (O_1093,N_13866,N_12086);
xor UO_1094 (O_1094,N_12808,N_13419);
nand UO_1095 (O_1095,N_13834,N_14429);
xnor UO_1096 (O_1096,N_12510,N_13210);
nor UO_1097 (O_1097,N_13766,N_12900);
xnor UO_1098 (O_1098,N_13854,N_12476);
or UO_1099 (O_1099,N_12872,N_14668);
or UO_1100 (O_1100,N_14562,N_13983);
or UO_1101 (O_1101,N_13903,N_13030);
and UO_1102 (O_1102,N_12637,N_12406);
xnor UO_1103 (O_1103,N_12268,N_12878);
xnor UO_1104 (O_1104,N_12821,N_13496);
nor UO_1105 (O_1105,N_12861,N_12119);
nor UO_1106 (O_1106,N_14059,N_12719);
xor UO_1107 (O_1107,N_13136,N_13305);
or UO_1108 (O_1108,N_13185,N_14464);
and UO_1109 (O_1109,N_12216,N_12404);
and UO_1110 (O_1110,N_12375,N_12006);
nor UO_1111 (O_1111,N_12123,N_14733);
nor UO_1112 (O_1112,N_14886,N_14837);
nand UO_1113 (O_1113,N_12769,N_12411);
nor UO_1114 (O_1114,N_14970,N_13888);
xor UO_1115 (O_1115,N_12758,N_13417);
or UO_1116 (O_1116,N_13720,N_13917);
xor UO_1117 (O_1117,N_12382,N_12532);
xnor UO_1118 (O_1118,N_14261,N_12994);
nor UO_1119 (O_1119,N_13871,N_14360);
or UO_1120 (O_1120,N_13758,N_14498);
and UO_1121 (O_1121,N_12131,N_14879);
xor UO_1122 (O_1122,N_14356,N_14422);
or UO_1123 (O_1123,N_14573,N_12727);
and UO_1124 (O_1124,N_14899,N_14281);
nand UO_1125 (O_1125,N_12919,N_12884);
and UO_1126 (O_1126,N_12657,N_13273);
nor UO_1127 (O_1127,N_14963,N_12434);
nand UO_1128 (O_1128,N_14560,N_13528);
nor UO_1129 (O_1129,N_13611,N_12571);
or UO_1130 (O_1130,N_14551,N_13343);
and UO_1131 (O_1131,N_14322,N_14236);
or UO_1132 (O_1132,N_14162,N_12841);
or UO_1133 (O_1133,N_14395,N_13878);
or UO_1134 (O_1134,N_12093,N_14935);
xnor UO_1135 (O_1135,N_12853,N_14638);
and UO_1136 (O_1136,N_13718,N_12075);
nor UO_1137 (O_1137,N_13234,N_13745);
or UO_1138 (O_1138,N_13596,N_12317);
xnor UO_1139 (O_1139,N_13374,N_14815);
nor UO_1140 (O_1140,N_12911,N_14268);
and UO_1141 (O_1141,N_12459,N_13796);
and UO_1142 (O_1142,N_14113,N_13831);
nor UO_1143 (O_1143,N_13515,N_12697);
xor UO_1144 (O_1144,N_14606,N_13867);
xnor UO_1145 (O_1145,N_14826,N_12698);
nand UO_1146 (O_1146,N_13118,N_14902);
and UO_1147 (O_1147,N_12372,N_12469);
nand UO_1148 (O_1148,N_14016,N_14501);
xor UO_1149 (O_1149,N_13315,N_14508);
xor UO_1150 (O_1150,N_13332,N_13384);
xnor UO_1151 (O_1151,N_12596,N_13615);
nor UO_1152 (O_1152,N_14491,N_12052);
xor UO_1153 (O_1153,N_13886,N_12361);
nor UO_1154 (O_1154,N_14419,N_13823);
nand UO_1155 (O_1155,N_12228,N_13112);
nand UO_1156 (O_1156,N_12324,N_12818);
or UO_1157 (O_1157,N_13005,N_13589);
nor UO_1158 (O_1158,N_14626,N_13283);
and UO_1159 (O_1159,N_12796,N_12251);
nor UO_1160 (O_1160,N_12629,N_13731);
xnor UO_1161 (O_1161,N_14913,N_13336);
nand UO_1162 (O_1162,N_12795,N_14838);
or UO_1163 (O_1163,N_12465,N_12882);
or UO_1164 (O_1164,N_13317,N_12367);
or UO_1165 (O_1165,N_13826,N_13463);
nor UO_1166 (O_1166,N_14516,N_14705);
nand UO_1167 (O_1167,N_12315,N_12579);
and UO_1168 (O_1168,N_12124,N_13570);
nor UO_1169 (O_1169,N_12887,N_14220);
xnor UO_1170 (O_1170,N_13647,N_12505);
and UO_1171 (O_1171,N_12618,N_14813);
nand UO_1172 (O_1172,N_13915,N_14166);
nor UO_1173 (O_1173,N_14431,N_12379);
nor UO_1174 (O_1174,N_12421,N_13223);
nor UO_1175 (O_1175,N_14831,N_14314);
and UO_1176 (O_1176,N_13448,N_14018);
and UO_1177 (O_1177,N_14296,N_12471);
nor UO_1178 (O_1178,N_14237,N_14877);
nand UO_1179 (O_1179,N_12116,N_14210);
nand UO_1180 (O_1180,N_14717,N_14725);
or UO_1181 (O_1181,N_12708,N_12067);
or UO_1182 (O_1182,N_13970,N_12051);
and UO_1183 (O_1183,N_13083,N_13328);
nand UO_1184 (O_1184,N_13895,N_13558);
xor UO_1185 (O_1185,N_12194,N_12318);
nor UO_1186 (O_1186,N_14149,N_13470);
xnor UO_1187 (O_1187,N_12568,N_13610);
and UO_1188 (O_1188,N_12314,N_13912);
nand UO_1189 (O_1189,N_13715,N_13835);
nor UO_1190 (O_1190,N_12527,N_12988);
or UO_1191 (O_1191,N_13276,N_14126);
or UO_1192 (O_1192,N_12946,N_14775);
or UO_1193 (O_1193,N_14012,N_12276);
xnor UO_1194 (O_1194,N_14739,N_12858);
or UO_1195 (O_1195,N_12754,N_13330);
nand UO_1196 (O_1196,N_13547,N_14154);
xnor UO_1197 (O_1197,N_13811,N_12148);
nand UO_1198 (O_1198,N_13424,N_12690);
xnor UO_1199 (O_1199,N_12740,N_14120);
nor UO_1200 (O_1200,N_12095,N_12875);
and UO_1201 (O_1201,N_12041,N_13208);
xor UO_1202 (O_1202,N_14253,N_14466);
xor UO_1203 (O_1203,N_13444,N_12896);
or UO_1204 (O_1204,N_12307,N_13949);
xor UO_1205 (O_1205,N_12346,N_13532);
and UO_1206 (O_1206,N_13062,N_14370);
nor UO_1207 (O_1207,N_14371,N_13585);
and UO_1208 (O_1208,N_13023,N_13651);
nor UO_1209 (O_1209,N_13486,N_12729);
xor UO_1210 (O_1210,N_13322,N_14614);
xor UO_1211 (O_1211,N_13399,N_13882);
or UO_1212 (O_1212,N_13116,N_12803);
nor UO_1213 (O_1213,N_13982,N_13838);
xnor UO_1214 (O_1214,N_14729,N_12611);
nor UO_1215 (O_1215,N_13331,N_13017);
or UO_1216 (O_1216,N_12992,N_12509);
nor UO_1217 (O_1217,N_14225,N_14796);
nand UO_1218 (O_1218,N_12980,N_14191);
or UO_1219 (O_1219,N_13501,N_14380);
nor UO_1220 (O_1220,N_13941,N_12564);
nor UO_1221 (O_1221,N_12288,N_14549);
or UO_1222 (O_1222,N_14146,N_13465);
xnor UO_1223 (O_1223,N_14618,N_14759);
xnor UO_1224 (O_1224,N_14651,N_13918);
and UO_1225 (O_1225,N_12756,N_12785);
or UO_1226 (O_1226,N_14784,N_13150);
xnor UO_1227 (O_1227,N_12782,N_12168);
nor UO_1228 (O_1228,N_13910,N_12895);
and UO_1229 (O_1229,N_14804,N_12384);
xnor UO_1230 (O_1230,N_12996,N_13710);
nor UO_1231 (O_1231,N_12903,N_12016);
nand UO_1232 (O_1232,N_12190,N_12398);
nor UO_1233 (O_1233,N_12169,N_13498);
nor UO_1234 (O_1234,N_14621,N_14258);
nor UO_1235 (O_1235,N_12786,N_14672);
xnor UO_1236 (O_1236,N_14404,N_13911);
xnor UO_1237 (O_1237,N_12053,N_13316);
nor UO_1238 (O_1238,N_14818,N_13698);
and UO_1239 (O_1239,N_12235,N_13584);
and UO_1240 (O_1240,N_14642,N_13773);
or UO_1241 (O_1241,N_14634,N_12178);
xnor UO_1242 (O_1242,N_13789,N_13452);
nor UO_1243 (O_1243,N_13077,N_14046);
nor UO_1244 (O_1244,N_12453,N_13078);
and UO_1245 (O_1245,N_13616,N_13197);
xnor UO_1246 (O_1246,N_14026,N_14817);
or UO_1247 (O_1247,N_12550,N_13632);
xor UO_1248 (O_1248,N_12807,N_12112);
nand UO_1249 (O_1249,N_14681,N_14136);
or UO_1250 (O_1250,N_14850,N_12325);
or UO_1251 (O_1251,N_14447,N_14465);
xnor UO_1252 (O_1252,N_13357,N_12647);
or UO_1253 (O_1253,N_12424,N_13014);
and UO_1254 (O_1254,N_14123,N_12172);
or UO_1255 (O_1255,N_12942,N_13015);
nor UO_1256 (O_1256,N_13269,N_13421);
and UO_1257 (O_1257,N_12673,N_13212);
xor UO_1258 (O_1258,N_12736,N_12724);
nand UO_1259 (O_1259,N_12050,N_12899);
xor UO_1260 (O_1260,N_12357,N_14934);
and UO_1261 (O_1261,N_12699,N_14297);
and UO_1262 (O_1262,N_13639,N_14423);
xnor UO_1263 (O_1263,N_13430,N_13684);
nand UO_1264 (O_1264,N_13101,N_13249);
or UO_1265 (O_1265,N_13128,N_13144);
xor UO_1266 (O_1266,N_13055,N_14480);
xor UO_1267 (O_1267,N_14628,N_12247);
nor UO_1268 (O_1268,N_14967,N_12702);
or UO_1269 (O_1269,N_12643,N_14922);
or UO_1270 (O_1270,N_12162,N_13828);
xor UO_1271 (O_1271,N_13750,N_13512);
and UO_1272 (O_1272,N_13495,N_13026);
nor UO_1273 (O_1273,N_12267,N_12447);
xnor UO_1274 (O_1274,N_13000,N_13353);
and UO_1275 (O_1275,N_14894,N_14586);
or UO_1276 (O_1276,N_14777,N_13676);
nor UO_1277 (O_1277,N_14669,N_12073);
and UO_1278 (O_1278,N_12344,N_12021);
or UO_1279 (O_1279,N_14050,N_14392);
or UO_1280 (O_1280,N_13153,N_12733);
nand UO_1281 (O_1281,N_13522,N_13818);
nor UO_1282 (O_1282,N_13453,N_14570);
or UO_1283 (O_1283,N_13919,N_14598);
xnor UO_1284 (O_1284,N_12358,N_12472);
xnor UO_1285 (O_1285,N_13637,N_14496);
nand UO_1286 (O_1286,N_14994,N_12791);
nor UO_1287 (O_1287,N_12117,N_12365);
and UO_1288 (O_1288,N_14364,N_14357);
nand UO_1289 (O_1289,N_12308,N_13905);
nand UO_1290 (O_1290,N_14998,N_12529);
and UO_1291 (O_1291,N_12293,N_13952);
and UO_1292 (O_1292,N_12871,N_12879);
and UO_1293 (O_1293,N_12488,N_12399);
and UO_1294 (O_1294,N_13184,N_12256);
nor UO_1295 (O_1295,N_13267,N_12522);
and UO_1296 (O_1296,N_12904,N_12120);
nor UO_1297 (O_1297,N_12691,N_13550);
xnor UO_1298 (O_1298,N_12076,N_13170);
xnor UO_1299 (O_1299,N_13908,N_14604);
nand UO_1300 (O_1300,N_14327,N_14363);
and UO_1301 (O_1301,N_12913,N_14742);
or UO_1302 (O_1302,N_12405,N_13497);
nand UO_1303 (O_1303,N_14481,N_12328);
nand UO_1304 (O_1304,N_13079,N_14888);
nand UO_1305 (O_1305,N_12966,N_12594);
or UO_1306 (O_1306,N_12888,N_13313);
xor UO_1307 (O_1307,N_13218,N_14202);
nand UO_1308 (O_1308,N_13485,N_14933);
and UO_1309 (O_1309,N_12111,N_12209);
nor UO_1310 (O_1310,N_12759,N_12078);
xor UO_1311 (O_1311,N_13787,N_12350);
nor UO_1312 (O_1312,N_14164,N_14876);
nand UO_1313 (O_1313,N_13138,N_12000);
xnor UO_1314 (O_1314,N_14111,N_14222);
and UO_1315 (O_1315,N_13856,N_14209);
xnor UO_1316 (O_1316,N_14727,N_12757);
and UO_1317 (O_1317,N_14833,N_14299);
nand UO_1318 (O_1318,N_14214,N_13338);
xor UO_1319 (O_1319,N_13035,N_13134);
nand UO_1320 (O_1320,N_12035,N_14385);
and UO_1321 (O_1321,N_14947,N_14420);
xnor UO_1322 (O_1322,N_13020,N_12464);
xor UO_1323 (O_1323,N_12436,N_14045);
nand UO_1324 (O_1324,N_14157,N_12363);
nor UO_1325 (O_1325,N_14787,N_14575);
or UO_1326 (O_1326,N_12419,N_12217);
nand UO_1327 (O_1327,N_13759,N_14912);
and UO_1328 (O_1328,N_13356,N_12481);
nand UO_1329 (O_1329,N_14832,N_13857);
and UO_1330 (O_1330,N_14701,N_13761);
and UO_1331 (O_1331,N_12619,N_13672);
and UO_1332 (O_1332,N_12547,N_12715);
nand UO_1333 (O_1333,N_14267,N_14802);
or UO_1334 (O_1334,N_14482,N_14859);
nor UO_1335 (O_1335,N_14020,N_13783);
and UO_1336 (O_1336,N_12961,N_14337);
nand UO_1337 (O_1337,N_12479,N_12061);
xnor UO_1338 (O_1338,N_12750,N_13756);
and UO_1339 (O_1339,N_12467,N_14585);
xor UO_1340 (O_1340,N_14971,N_12885);
xnor UO_1341 (O_1341,N_12309,N_14221);
and UO_1342 (O_1342,N_14579,N_12726);
nand UO_1343 (O_1343,N_13529,N_13760);
nor UO_1344 (O_1344,N_12968,N_12427);
nand UO_1345 (O_1345,N_14937,N_12604);
nand UO_1346 (O_1346,N_14635,N_13462);
xor UO_1347 (O_1347,N_13311,N_12001);
xor UO_1348 (O_1348,N_13967,N_14151);
nor UO_1349 (O_1349,N_13820,N_13409);
xnor UO_1350 (O_1350,N_13236,N_12909);
and UO_1351 (O_1351,N_13120,N_12484);
and UO_1352 (O_1352,N_13803,N_12304);
or UO_1353 (O_1353,N_14014,N_13171);
or UO_1354 (O_1354,N_13980,N_14722);
nand UO_1355 (O_1355,N_12941,N_14943);
xor UO_1356 (O_1356,N_14180,N_13289);
and UO_1357 (O_1357,N_12914,N_14754);
nand UO_1358 (O_1358,N_12874,N_12212);
or UO_1359 (O_1359,N_13198,N_12354);
nand UO_1360 (O_1360,N_12762,N_13479);
or UO_1361 (O_1361,N_13310,N_13428);
xor UO_1362 (O_1362,N_14206,N_12728);
nor UO_1363 (O_1363,N_14323,N_13088);
nand UO_1364 (O_1364,N_14332,N_14622);
xor UO_1365 (O_1365,N_12121,N_12491);
and UO_1366 (O_1366,N_12007,N_12198);
or UO_1367 (O_1367,N_12694,N_13114);
or UO_1368 (O_1368,N_14023,N_14176);
nand UO_1369 (O_1369,N_12030,N_12056);
xnor UO_1370 (O_1370,N_12380,N_13936);
nor UO_1371 (O_1371,N_12390,N_14331);
nor UO_1372 (O_1372,N_13790,N_13016);
and UO_1373 (O_1373,N_14044,N_13562);
and UO_1374 (O_1374,N_14794,N_12748);
nand UO_1375 (O_1375,N_14114,N_14723);
xor UO_1376 (O_1376,N_14031,N_13431);
nand UO_1377 (O_1377,N_13389,N_14345);
xnor UO_1378 (O_1378,N_13348,N_12184);
and UO_1379 (O_1379,N_13188,N_12010);
xnor UO_1380 (O_1380,N_13490,N_14022);
nor UO_1381 (O_1381,N_13680,N_12912);
and UO_1382 (O_1382,N_13729,N_12886);
nor UO_1383 (O_1383,N_12767,N_14519);
nor UO_1384 (O_1384,N_14732,N_13204);
nand UO_1385 (O_1385,N_13946,N_12306);
or UO_1386 (O_1386,N_13646,N_14568);
xor UO_1387 (O_1387,N_13654,N_14372);
nor UO_1388 (O_1388,N_12660,N_12517);
nand UO_1389 (O_1389,N_14882,N_14521);
or UO_1390 (O_1390,N_13021,N_12283);
or UO_1391 (O_1391,N_14131,N_14769);
and UO_1392 (O_1392,N_13628,N_14627);
nor UO_1393 (O_1393,N_13652,N_13507);
nand UO_1394 (O_1394,N_14224,N_12679);
or UO_1395 (O_1395,N_14602,N_12353);
xor UO_1396 (O_1396,N_12593,N_13706);
and UO_1397 (O_1397,N_14174,N_13738);
nor UO_1398 (O_1398,N_12908,N_12695);
xor UO_1399 (O_1399,N_12468,N_12290);
nor UO_1400 (O_1400,N_12038,N_13108);
and UO_1401 (O_1401,N_12150,N_14987);
and UO_1402 (O_1402,N_14932,N_14625);
and UO_1403 (O_1403,N_13538,N_12327);
and UO_1404 (O_1404,N_14140,N_14159);
and UO_1405 (O_1405,N_12177,N_13846);
nor UO_1406 (O_1406,N_12239,N_12670);
and UO_1407 (O_1407,N_12631,N_13873);
nor UO_1408 (O_1408,N_12208,N_12201);
or UO_1409 (O_1409,N_12146,N_13855);
and UO_1410 (O_1410,N_12820,N_14639);
xor UO_1411 (O_1411,N_12081,N_12294);
and UO_1412 (O_1412,N_13926,N_12138);
nand UO_1413 (O_1413,N_13893,N_12671);
xor UO_1414 (O_1414,N_14580,N_13587);
or UO_1415 (O_1415,N_13245,N_14688);
nand UO_1416 (O_1416,N_14993,N_14641);
xor UO_1417 (O_1417,N_13775,N_14035);
or UO_1418 (O_1418,N_12183,N_14948);
or UO_1419 (O_1419,N_12971,N_13525);
nor UO_1420 (O_1420,N_14094,N_14132);
nor UO_1421 (O_1421,N_13816,N_13058);
and UO_1422 (O_1422,N_14070,N_14540);
or UO_1423 (O_1423,N_13806,N_14849);
nor UO_1424 (O_1424,N_13935,N_12897);
nor UO_1425 (O_1425,N_12341,N_13690);
xnor UO_1426 (O_1426,N_12077,N_14537);
xnor UO_1427 (O_1427,N_13451,N_14648);
and UO_1428 (O_1428,N_13379,N_14148);
xor UO_1429 (O_1429,N_12989,N_13502);
nor UO_1430 (O_1430,N_14239,N_14444);
nor UO_1431 (O_1431,N_13145,N_13809);
nand UO_1432 (O_1432,N_13901,N_14730);
and UO_1433 (O_1433,N_13074,N_14768);
xnor UO_1434 (O_1434,N_12781,N_12392);
nand UO_1435 (O_1435,N_13388,N_12582);
and UO_1436 (O_1436,N_13531,N_12730);
nand UO_1437 (O_1437,N_13437,N_14257);
nand UO_1438 (O_1438,N_13769,N_14141);
nand UO_1439 (O_1439,N_13287,N_13517);
nand UO_1440 (O_1440,N_12295,N_12806);
nand UO_1441 (O_1441,N_14941,N_14089);
nand UO_1442 (O_1442,N_12260,N_12004);
or UO_1443 (O_1443,N_12768,N_12783);
nand UO_1444 (O_1444,N_12981,N_13618);
and UO_1445 (O_1445,N_13288,N_13298);
and UO_1446 (O_1446,N_14275,N_13991);
and UO_1447 (O_1447,N_12189,N_14230);
and UO_1448 (O_1448,N_13944,N_14595);
xor UO_1449 (O_1449,N_13178,N_12764);
xor UO_1450 (O_1450,N_13650,N_12486);
nor UO_1451 (O_1451,N_12907,N_14051);
xor UO_1452 (O_1452,N_13753,N_12287);
xor UO_1453 (O_1453,N_14695,N_13922);
nor UO_1454 (O_1454,N_12539,N_13555);
xnor UO_1455 (O_1455,N_12743,N_13043);
nor UO_1456 (O_1456,N_13285,N_14290);
nor UO_1457 (O_1457,N_12862,N_14302);
and UO_1458 (O_1458,N_12388,N_13649);
nand UO_1459 (O_1459,N_13345,N_13539);
and UO_1460 (O_1460,N_13177,N_14244);
nand UO_1461 (O_1461,N_12282,N_12391);
or UO_1462 (O_1462,N_14460,N_12588);
or UO_1463 (O_1463,N_13859,N_13250);
xnor UO_1464 (O_1464,N_14010,N_12236);
nand UO_1465 (O_1465,N_14366,N_13099);
nand UO_1466 (O_1466,N_12487,N_14842);
and UO_1467 (O_1467,N_14101,N_14953);
and UO_1468 (O_1468,N_14791,N_12105);
nor UO_1469 (O_1469,N_13757,N_14884);
nand UO_1470 (O_1470,N_14517,N_13975);
xor UO_1471 (O_1471,N_13027,N_14124);
or UO_1472 (O_1472,N_12676,N_13586);
or UO_1473 (O_1473,N_13247,N_12159);
or UO_1474 (O_1474,N_14353,N_14233);
xor UO_1475 (O_1475,N_12045,N_13053);
nor UO_1476 (O_1476,N_12924,N_14687);
or UO_1477 (O_1477,N_14809,N_12211);
xor UO_1478 (O_1478,N_12461,N_14564);
or UO_1479 (O_1479,N_13825,N_14735);
nand UO_1480 (O_1480,N_13577,N_14155);
or UO_1481 (O_1481,N_12763,N_13947);
and UO_1482 (O_1482,N_14085,N_14454);
xor UO_1483 (O_1483,N_12266,N_12666);
xor UO_1484 (O_1484,N_13930,N_14307);
or UO_1485 (O_1485,N_12431,N_13830);
or UO_1486 (O_1486,N_14719,N_13224);
nor UO_1487 (O_1487,N_14823,N_13524);
and UO_1488 (O_1488,N_13614,N_13808);
xnor UO_1489 (O_1489,N_13770,N_14511);
xnor UO_1490 (O_1490,N_14952,N_14414);
and UO_1491 (O_1491,N_14724,N_12815);
and UO_1492 (O_1492,N_13042,N_14702);
or UO_1493 (O_1493,N_12583,N_13934);
nor UO_1494 (O_1494,N_13518,N_13640);
or UO_1495 (O_1495,N_13412,N_12137);
nand UO_1496 (O_1496,N_14515,N_13380);
and UO_1497 (O_1497,N_14107,N_12834);
nand UO_1498 (O_1498,N_12824,N_12656);
xor UO_1499 (O_1499,N_14664,N_14633);
xnor UO_1500 (O_1500,N_14660,N_12609);
nor UO_1501 (O_1501,N_12027,N_14685);
nand UO_1502 (O_1502,N_14988,N_12990);
nor UO_1503 (O_1503,N_12422,N_14919);
nand UO_1504 (O_1504,N_12500,N_13196);
or UO_1505 (O_1505,N_14494,N_14702);
nand UO_1506 (O_1506,N_13475,N_12882);
xnor UO_1507 (O_1507,N_12614,N_12954);
and UO_1508 (O_1508,N_13043,N_14219);
or UO_1509 (O_1509,N_13908,N_13545);
nand UO_1510 (O_1510,N_14199,N_13385);
nand UO_1511 (O_1511,N_13981,N_13125);
nand UO_1512 (O_1512,N_12658,N_12405);
nor UO_1513 (O_1513,N_12173,N_13696);
and UO_1514 (O_1514,N_12072,N_13892);
or UO_1515 (O_1515,N_14061,N_14527);
xor UO_1516 (O_1516,N_14556,N_14086);
or UO_1517 (O_1517,N_14700,N_12315);
xnor UO_1518 (O_1518,N_12405,N_12993);
nor UO_1519 (O_1519,N_13673,N_13105);
and UO_1520 (O_1520,N_12674,N_12394);
and UO_1521 (O_1521,N_14760,N_14721);
nand UO_1522 (O_1522,N_14844,N_14723);
nor UO_1523 (O_1523,N_14663,N_12523);
xnor UO_1524 (O_1524,N_12966,N_12821);
and UO_1525 (O_1525,N_14638,N_13415);
nand UO_1526 (O_1526,N_13624,N_13492);
and UO_1527 (O_1527,N_13773,N_13823);
and UO_1528 (O_1528,N_14845,N_13354);
nand UO_1529 (O_1529,N_14228,N_12265);
nor UO_1530 (O_1530,N_12207,N_13429);
and UO_1531 (O_1531,N_13259,N_12239);
nand UO_1532 (O_1532,N_14602,N_13618);
and UO_1533 (O_1533,N_12785,N_13315);
xor UO_1534 (O_1534,N_12982,N_14400);
xnor UO_1535 (O_1535,N_14850,N_13278);
nor UO_1536 (O_1536,N_12269,N_12449);
nor UO_1537 (O_1537,N_13431,N_14885);
xor UO_1538 (O_1538,N_14941,N_14444);
or UO_1539 (O_1539,N_14324,N_14905);
nand UO_1540 (O_1540,N_13999,N_14673);
nor UO_1541 (O_1541,N_14774,N_14829);
nand UO_1542 (O_1542,N_13280,N_12235);
and UO_1543 (O_1543,N_12124,N_14627);
or UO_1544 (O_1544,N_13908,N_14413);
or UO_1545 (O_1545,N_14651,N_14262);
nand UO_1546 (O_1546,N_14968,N_13472);
nand UO_1547 (O_1547,N_12362,N_12947);
xnor UO_1548 (O_1548,N_13197,N_12358);
nor UO_1549 (O_1549,N_12078,N_12607);
nor UO_1550 (O_1550,N_12494,N_12866);
or UO_1551 (O_1551,N_14666,N_13812);
nand UO_1552 (O_1552,N_13678,N_12214);
and UO_1553 (O_1553,N_13282,N_13988);
or UO_1554 (O_1554,N_12730,N_12898);
or UO_1555 (O_1555,N_13998,N_13407);
or UO_1556 (O_1556,N_14339,N_12382);
or UO_1557 (O_1557,N_13712,N_13989);
and UO_1558 (O_1558,N_14548,N_12630);
or UO_1559 (O_1559,N_12612,N_14381);
nor UO_1560 (O_1560,N_14760,N_14229);
xnor UO_1561 (O_1561,N_12066,N_13685);
and UO_1562 (O_1562,N_14573,N_14272);
nor UO_1563 (O_1563,N_13784,N_12143);
nor UO_1564 (O_1564,N_12964,N_14929);
nor UO_1565 (O_1565,N_12627,N_14098);
nor UO_1566 (O_1566,N_12213,N_12620);
and UO_1567 (O_1567,N_14413,N_12973);
xor UO_1568 (O_1568,N_14498,N_14153);
nand UO_1569 (O_1569,N_12313,N_13052);
xnor UO_1570 (O_1570,N_13146,N_13363);
and UO_1571 (O_1571,N_14305,N_14307);
and UO_1572 (O_1572,N_14802,N_13386);
nand UO_1573 (O_1573,N_12816,N_14392);
nor UO_1574 (O_1574,N_13723,N_14230);
xnor UO_1575 (O_1575,N_12705,N_13583);
and UO_1576 (O_1576,N_14917,N_14586);
or UO_1577 (O_1577,N_12103,N_12316);
nand UO_1578 (O_1578,N_13911,N_13499);
and UO_1579 (O_1579,N_13093,N_12726);
xor UO_1580 (O_1580,N_12058,N_14828);
and UO_1581 (O_1581,N_13660,N_13449);
or UO_1582 (O_1582,N_13540,N_13875);
xor UO_1583 (O_1583,N_12512,N_13484);
and UO_1584 (O_1584,N_14153,N_12600);
or UO_1585 (O_1585,N_12492,N_12073);
xnor UO_1586 (O_1586,N_12938,N_14867);
nand UO_1587 (O_1587,N_12747,N_14881);
or UO_1588 (O_1588,N_13072,N_13006);
xnor UO_1589 (O_1589,N_14494,N_13307);
or UO_1590 (O_1590,N_13013,N_12976);
nand UO_1591 (O_1591,N_12838,N_13398);
or UO_1592 (O_1592,N_14671,N_14654);
or UO_1593 (O_1593,N_14266,N_12147);
or UO_1594 (O_1594,N_14542,N_13934);
xnor UO_1595 (O_1595,N_13761,N_12598);
nor UO_1596 (O_1596,N_13654,N_12127);
nor UO_1597 (O_1597,N_13555,N_13201);
or UO_1598 (O_1598,N_12919,N_14460);
nand UO_1599 (O_1599,N_12385,N_12113);
nor UO_1600 (O_1600,N_13790,N_12348);
xnor UO_1601 (O_1601,N_12277,N_14417);
nand UO_1602 (O_1602,N_13718,N_13323);
nand UO_1603 (O_1603,N_12456,N_14620);
or UO_1604 (O_1604,N_12015,N_12064);
and UO_1605 (O_1605,N_13929,N_12114);
nand UO_1606 (O_1606,N_14197,N_13937);
nand UO_1607 (O_1607,N_13073,N_13672);
and UO_1608 (O_1608,N_13250,N_12863);
nor UO_1609 (O_1609,N_13737,N_13268);
or UO_1610 (O_1610,N_13963,N_14209);
and UO_1611 (O_1611,N_14478,N_12466);
or UO_1612 (O_1612,N_13166,N_13807);
and UO_1613 (O_1613,N_14701,N_13399);
or UO_1614 (O_1614,N_14588,N_14212);
and UO_1615 (O_1615,N_13623,N_14435);
or UO_1616 (O_1616,N_14528,N_12138);
xnor UO_1617 (O_1617,N_13233,N_14812);
xor UO_1618 (O_1618,N_13710,N_12706);
xnor UO_1619 (O_1619,N_14782,N_13266);
nor UO_1620 (O_1620,N_12969,N_13713);
nor UO_1621 (O_1621,N_12669,N_13730);
nand UO_1622 (O_1622,N_14158,N_12174);
and UO_1623 (O_1623,N_12982,N_12355);
or UO_1624 (O_1624,N_12249,N_14778);
or UO_1625 (O_1625,N_13849,N_12320);
or UO_1626 (O_1626,N_14387,N_12935);
xor UO_1627 (O_1627,N_12314,N_14522);
and UO_1628 (O_1628,N_13934,N_13222);
nand UO_1629 (O_1629,N_12628,N_14183);
xnor UO_1630 (O_1630,N_13111,N_14030);
or UO_1631 (O_1631,N_14092,N_12373);
nand UO_1632 (O_1632,N_14931,N_14764);
nor UO_1633 (O_1633,N_12976,N_13973);
and UO_1634 (O_1634,N_12062,N_13308);
xnor UO_1635 (O_1635,N_14820,N_13290);
xor UO_1636 (O_1636,N_14456,N_14336);
or UO_1637 (O_1637,N_14451,N_14674);
nor UO_1638 (O_1638,N_13481,N_14825);
nor UO_1639 (O_1639,N_12491,N_13716);
nand UO_1640 (O_1640,N_13759,N_13813);
or UO_1641 (O_1641,N_14249,N_14584);
or UO_1642 (O_1642,N_14248,N_14310);
xnor UO_1643 (O_1643,N_12225,N_14237);
and UO_1644 (O_1644,N_13989,N_14959);
and UO_1645 (O_1645,N_14489,N_12985);
xnor UO_1646 (O_1646,N_13430,N_13244);
or UO_1647 (O_1647,N_14447,N_13199);
and UO_1648 (O_1648,N_13703,N_13476);
nand UO_1649 (O_1649,N_12001,N_13312);
xor UO_1650 (O_1650,N_13761,N_13146);
nor UO_1651 (O_1651,N_14952,N_12684);
nand UO_1652 (O_1652,N_13752,N_13693);
nand UO_1653 (O_1653,N_13979,N_13016);
xnor UO_1654 (O_1654,N_12033,N_12778);
xor UO_1655 (O_1655,N_12385,N_12256);
and UO_1656 (O_1656,N_14814,N_14223);
or UO_1657 (O_1657,N_14616,N_13911);
xnor UO_1658 (O_1658,N_12718,N_12102);
and UO_1659 (O_1659,N_13943,N_12743);
xnor UO_1660 (O_1660,N_12203,N_14677);
xor UO_1661 (O_1661,N_12139,N_13644);
nor UO_1662 (O_1662,N_14503,N_12555);
and UO_1663 (O_1663,N_12163,N_14205);
or UO_1664 (O_1664,N_13796,N_13276);
xor UO_1665 (O_1665,N_13369,N_13405);
and UO_1666 (O_1666,N_13273,N_13199);
xor UO_1667 (O_1667,N_12518,N_12498);
and UO_1668 (O_1668,N_12819,N_13084);
nor UO_1669 (O_1669,N_13000,N_12394);
nor UO_1670 (O_1670,N_12610,N_13699);
xor UO_1671 (O_1671,N_14574,N_14727);
and UO_1672 (O_1672,N_12795,N_13220);
nand UO_1673 (O_1673,N_14612,N_12254);
or UO_1674 (O_1674,N_14824,N_14709);
or UO_1675 (O_1675,N_14588,N_13900);
xnor UO_1676 (O_1676,N_12364,N_14678);
nor UO_1677 (O_1677,N_12988,N_12564);
or UO_1678 (O_1678,N_13465,N_12101);
and UO_1679 (O_1679,N_14229,N_13928);
nor UO_1680 (O_1680,N_12088,N_12146);
nand UO_1681 (O_1681,N_13015,N_12588);
nor UO_1682 (O_1682,N_14174,N_13230);
xor UO_1683 (O_1683,N_13328,N_12610);
and UO_1684 (O_1684,N_13089,N_13555);
nor UO_1685 (O_1685,N_12087,N_12812);
xor UO_1686 (O_1686,N_13745,N_13135);
and UO_1687 (O_1687,N_14397,N_14303);
and UO_1688 (O_1688,N_13902,N_13536);
or UO_1689 (O_1689,N_12116,N_13015);
nand UO_1690 (O_1690,N_14308,N_14752);
or UO_1691 (O_1691,N_12165,N_12354);
nor UO_1692 (O_1692,N_13537,N_14618);
nor UO_1693 (O_1693,N_12921,N_13021);
xor UO_1694 (O_1694,N_14751,N_12419);
nand UO_1695 (O_1695,N_13725,N_13381);
and UO_1696 (O_1696,N_14513,N_12564);
nand UO_1697 (O_1697,N_14453,N_13452);
xor UO_1698 (O_1698,N_14357,N_13398);
nor UO_1699 (O_1699,N_13723,N_13753);
xor UO_1700 (O_1700,N_14719,N_14174);
xor UO_1701 (O_1701,N_14272,N_12348);
nand UO_1702 (O_1702,N_14219,N_13982);
nand UO_1703 (O_1703,N_14161,N_13466);
or UO_1704 (O_1704,N_14562,N_14950);
and UO_1705 (O_1705,N_12264,N_13897);
nand UO_1706 (O_1706,N_14736,N_12607);
xor UO_1707 (O_1707,N_12693,N_12681);
and UO_1708 (O_1708,N_14124,N_14659);
nor UO_1709 (O_1709,N_14831,N_13265);
nand UO_1710 (O_1710,N_13340,N_12575);
xor UO_1711 (O_1711,N_14564,N_14769);
or UO_1712 (O_1712,N_14804,N_12772);
nand UO_1713 (O_1713,N_14275,N_12062);
xor UO_1714 (O_1714,N_12514,N_12652);
or UO_1715 (O_1715,N_12832,N_13633);
xnor UO_1716 (O_1716,N_12618,N_13703);
and UO_1717 (O_1717,N_13375,N_12801);
nand UO_1718 (O_1718,N_13688,N_14379);
nand UO_1719 (O_1719,N_12765,N_13547);
xnor UO_1720 (O_1720,N_13576,N_12556);
or UO_1721 (O_1721,N_12363,N_14703);
nand UO_1722 (O_1722,N_13481,N_13610);
or UO_1723 (O_1723,N_13337,N_14606);
nand UO_1724 (O_1724,N_13412,N_14913);
xnor UO_1725 (O_1725,N_14357,N_13152);
nor UO_1726 (O_1726,N_12329,N_13322);
xor UO_1727 (O_1727,N_13666,N_13646);
nor UO_1728 (O_1728,N_13843,N_13057);
xor UO_1729 (O_1729,N_14656,N_13854);
nand UO_1730 (O_1730,N_13115,N_14711);
nand UO_1731 (O_1731,N_13720,N_12414);
or UO_1732 (O_1732,N_12540,N_14200);
nor UO_1733 (O_1733,N_13927,N_13624);
xnor UO_1734 (O_1734,N_14498,N_12885);
nor UO_1735 (O_1735,N_14561,N_13043);
nor UO_1736 (O_1736,N_12177,N_14748);
nand UO_1737 (O_1737,N_13388,N_12517);
or UO_1738 (O_1738,N_13648,N_12069);
and UO_1739 (O_1739,N_14741,N_13545);
and UO_1740 (O_1740,N_12634,N_14630);
or UO_1741 (O_1741,N_14696,N_13893);
nor UO_1742 (O_1742,N_13393,N_13658);
xnor UO_1743 (O_1743,N_14007,N_12000);
or UO_1744 (O_1744,N_12195,N_13590);
xnor UO_1745 (O_1745,N_14622,N_14458);
nand UO_1746 (O_1746,N_12462,N_14638);
or UO_1747 (O_1747,N_12254,N_14797);
xnor UO_1748 (O_1748,N_12216,N_14596);
nand UO_1749 (O_1749,N_12747,N_13306);
or UO_1750 (O_1750,N_14880,N_12495);
xor UO_1751 (O_1751,N_12753,N_14525);
nand UO_1752 (O_1752,N_13302,N_13190);
nand UO_1753 (O_1753,N_14076,N_12844);
nand UO_1754 (O_1754,N_14834,N_13303);
nor UO_1755 (O_1755,N_14149,N_13091);
or UO_1756 (O_1756,N_13760,N_12598);
nor UO_1757 (O_1757,N_13589,N_13246);
and UO_1758 (O_1758,N_14573,N_12059);
or UO_1759 (O_1759,N_14647,N_12572);
and UO_1760 (O_1760,N_13999,N_12886);
and UO_1761 (O_1761,N_13598,N_14819);
nand UO_1762 (O_1762,N_12493,N_12144);
nand UO_1763 (O_1763,N_13393,N_12541);
or UO_1764 (O_1764,N_13179,N_14619);
or UO_1765 (O_1765,N_13396,N_13625);
and UO_1766 (O_1766,N_14092,N_14468);
nand UO_1767 (O_1767,N_14003,N_13579);
or UO_1768 (O_1768,N_13857,N_13224);
or UO_1769 (O_1769,N_12082,N_14759);
and UO_1770 (O_1770,N_12138,N_12246);
nor UO_1771 (O_1771,N_14363,N_14199);
nor UO_1772 (O_1772,N_13728,N_12888);
nand UO_1773 (O_1773,N_12626,N_12409);
nor UO_1774 (O_1774,N_12611,N_14133);
xnor UO_1775 (O_1775,N_13465,N_12183);
and UO_1776 (O_1776,N_12966,N_13690);
or UO_1777 (O_1777,N_13104,N_12780);
and UO_1778 (O_1778,N_14280,N_12497);
nor UO_1779 (O_1779,N_12216,N_14365);
or UO_1780 (O_1780,N_14139,N_12615);
xor UO_1781 (O_1781,N_14614,N_12458);
and UO_1782 (O_1782,N_14932,N_12278);
xor UO_1783 (O_1783,N_13586,N_12546);
xnor UO_1784 (O_1784,N_12410,N_13070);
nor UO_1785 (O_1785,N_14932,N_13500);
nor UO_1786 (O_1786,N_13107,N_12431);
or UO_1787 (O_1787,N_13717,N_14061);
or UO_1788 (O_1788,N_13223,N_12617);
xnor UO_1789 (O_1789,N_13146,N_14557);
nand UO_1790 (O_1790,N_12099,N_13509);
or UO_1791 (O_1791,N_14374,N_14795);
nor UO_1792 (O_1792,N_13451,N_13148);
nor UO_1793 (O_1793,N_14725,N_13530);
nand UO_1794 (O_1794,N_14695,N_14173);
and UO_1795 (O_1795,N_12005,N_13708);
nand UO_1796 (O_1796,N_12046,N_14922);
xnor UO_1797 (O_1797,N_13230,N_13168);
nand UO_1798 (O_1798,N_12642,N_12017);
nor UO_1799 (O_1799,N_13554,N_14185);
nor UO_1800 (O_1800,N_13285,N_14178);
or UO_1801 (O_1801,N_13623,N_14527);
xnor UO_1802 (O_1802,N_12604,N_12435);
or UO_1803 (O_1803,N_13351,N_12159);
or UO_1804 (O_1804,N_13989,N_13796);
nor UO_1805 (O_1805,N_12163,N_14224);
or UO_1806 (O_1806,N_13003,N_12723);
and UO_1807 (O_1807,N_14675,N_12181);
nand UO_1808 (O_1808,N_13763,N_13020);
nor UO_1809 (O_1809,N_13832,N_12883);
nand UO_1810 (O_1810,N_13664,N_14534);
nor UO_1811 (O_1811,N_12316,N_14786);
or UO_1812 (O_1812,N_14227,N_14664);
nor UO_1813 (O_1813,N_14147,N_14207);
nand UO_1814 (O_1814,N_13011,N_12465);
or UO_1815 (O_1815,N_12529,N_14636);
xor UO_1816 (O_1816,N_12410,N_14807);
nor UO_1817 (O_1817,N_13991,N_12176);
or UO_1818 (O_1818,N_14391,N_14454);
and UO_1819 (O_1819,N_13121,N_13973);
xor UO_1820 (O_1820,N_12932,N_12363);
nand UO_1821 (O_1821,N_12693,N_13844);
xor UO_1822 (O_1822,N_14376,N_12253);
nor UO_1823 (O_1823,N_13122,N_14429);
xnor UO_1824 (O_1824,N_14884,N_13747);
nor UO_1825 (O_1825,N_12596,N_12923);
or UO_1826 (O_1826,N_13772,N_13297);
nor UO_1827 (O_1827,N_13568,N_14767);
xnor UO_1828 (O_1828,N_13755,N_14944);
nor UO_1829 (O_1829,N_12201,N_13694);
nand UO_1830 (O_1830,N_12726,N_12214);
and UO_1831 (O_1831,N_12165,N_13049);
or UO_1832 (O_1832,N_12140,N_14724);
nor UO_1833 (O_1833,N_12345,N_13760);
or UO_1834 (O_1834,N_12402,N_14365);
nor UO_1835 (O_1835,N_12122,N_13584);
xnor UO_1836 (O_1836,N_12771,N_14056);
xor UO_1837 (O_1837,N_12932,N_14002);
nand UO_1838 (O_1838,N_13747,N_13850);
and UO_1839 (O_1839,N_13080,N_14268);
or UO_1840 (O_1840,N_14054,N_14901);
nor UO_1841 (O_1841,N_13395,N_12303);
or UO_1842 (O_1842,N_13889,N_14262);
or UO_1843 (O_1843,N_13640,N_12045);
nand UO_1844 (O_1844,N_14965,N_12422);
nand UO_1845 (O_1845,N_13905,N_13957);
and UO_1846 (O_1846,N_13938,N_14321);
nand UO_1847 (O_1847,N_13263,N_13320);
nor UO_1848 (O_1848,N_12162,N_12121);
or UO_1849 (O_1849,N_14137,N_14101);
nor UO_1850 (O_1850,N_14651,N_14846);
xnor UO_1851 (O_1851,N_13414,N_14584);
nor UO_1852 (O_1852,N_13183,N_12923);
or UO_1853 (O_1853,N_13095,N_13157);
xnor UO_1854 (O_1854,N_13320,N_14086);
and UO_1855 (O_1855,N_12539,N_14462);
nor UO_1856 (O_1856,N_13162,N_12764);
xnor UO_1857 (O_1857,N_14294,N_12613);
nor UO_1858 (O_1858,N_12912,N_14592);
and UO_1859 (O_1859,N_14750,N_12998);
nor UO_1860 (O_1860,N_12238,N_13475);
or UO_1861 (O_1861,N_14448,N_14109);
xnor UO_1862 (O_1862,N_14227,N_13290);
and UO_1863 (O_1863,N_12763,N_14843);
or UO_1864 (O_1864,N_13743,N_12746);
or UO_1865 (O_1865,N_12092,N_12578);
xor UO_1866 (O_1866,N_12986,N_12427);
nand UO_1867 (O_1867,N_13502,N_12763);
nor UO_1868 (O_1868,N_13946,N_12327);
xor UO_1869 (O_1869,N_12998,N_13654);
and UO_1870 (O_1870,N_13976,N_14415);
or UO_1871 (O_1871,N_12231,N_14205);
nor UO_1872 (O_1872,N_12872,N_14679);
nor UO_1873 (O_1873,N_13328,N_14220);
and UO_1874 (O_1874,N_12360,N_13227);
nor UO_1875 (O_1875,N_13292,N_14410);
nand UO_1876 (O_1876,N_13548,N_13833);
or UO_1877 (O_1877,N_14726,N_13954);
nand UO_1878 (O_1878,N_13141,N_12793);
nor UO_1879 (O_1879,N_13221,N_12458);
nand UO_1880 (O_1880,N_14721,N_12715);
or UO_1881 (O_1881,N_12913,N_13788);
and UO_1882 (O_1882,N_14002,N_13305);
nand UO_1883 (O_1883,N_12957,N_14368);
and UO_1884 (O_1884,N_14131,N_12386);
and UO_1885 (O_1885,N_12412,N_12446);
or UO_1886 (O_1886,N_13295,N_12888);
xnor UO_1887 (O_1887,N_13034,N_13774);
nand UO_1888 (O_1888,N_12849,N_14216);
and UO_1889 (O_1889,N_12289,N_12857);
and UO_1890 (O_1890,N_12205,N_12155);
xor UO_1891 (O_1891,N_12898,N_14895);
xnor UO_1892 (O_1892,N_12553,N_13359);
xor UO_1893 (O_1893,N_12161,N_12420);
or UO_1894 (O_1894,N_13898,N_12610);
nor UO_1895 (O_1895,N_13179,N_12039);
xnor UO_1896 (O_1896,N_14382,N_14642);
xor UO_1897 (O_1897,N_12869,N_14149);
nor UO_1898 (O_1898,N_13803,N_13274);
and UO_1899 (O_1899,N_12499,N_13968);
xor UO_1900 (O_1900,N_12511,N_13422);
xor UO_1901 (O_1901,N_12432,N_12772);
nor UO_1902 (O_1902,N_13887,N_13383);
or UO_1903 (O_1903,N_12387,N_12987);
or UO_1904 (O_1904,N_14426,N_12861);
nor UO_1905 (O_1905,N_12065,N_13572);
nor UO_1906 (O_1906,N_14724,N_13138);
xnor UO_1907 (O_1907,N_14130,N_13396);
nor UO_1908 (O_1908,N_13865,N_13365);
or UO_1909 (O_1909,N_14082,N_12272);
or UO_1910 (O_1910,N_13045,N_14806);
xnor UO_1911 (O_1911,N_13311,N_12792);
xor UO_1912 (O_1912,N_12290,N_12397);
or UO_1913 (O_1913,N_12488,N_13670);
or UO_1914 (O_1914,N_13755,N_14631);
nor UO_1915 (O_1915,N_13793,N_13604);
nor UO_1916 (O_1916,N_14738,N_12674);
or UO_1917 (O_1917,N_12578,N_13334);
and UO_1918 (O_1918,N_14550,N_14822);
nor UO_1919 (O_1919,N_13175,N_12272);
or UO_1920 (O_1920,N_13233,N_12951);
and UO_1921 (O_1921,N_13945,N_12115);
or UO_1922 (O_1922,N_14759,N_12619);
or UO_1923 (O_1923,N_14098,N_13015);
xnor UO_1924 (O_1924,N_14133,N_14267);
xnor UO_1925 (O_1925,N_13802,N_13797);
and UO_1926 (O_1926,N_13647,N_14246);
or UO_1927 (O_1927,N_12392,N_12572);
nand UO_1928 (O_1928,N_14255,N_14634);
or UO_1929 (O_1929,N_12499,N_13191);
xor UO_1930 (O_1930,N_14414,N_12463);
xnor UO_1931 (O_1931,N_14684,N_12757);
or UO_1932 (O_1932,N_13908,N_13459);
nor UO_1933 (O_1933,N_12783,N_12679);
nand UO_1934 (O_1934,N_14485,N_13829);
xnor UO_1935 (O_1935,N_13673,N_14116);
nand UO_1936 (O_1936,N_13320,N_14285);
nor UO_1937 (O_1937,N_12167,N_14581);
and UO_1938 (O_1938,N_12404,N_14989);
nor UO_1939 (O_1939,N_12423,N_12860);
nand UO_1940 (O_1940,N_12019,N_13643);
and UO_1941 (O_1941,N_12979,N_14249);
nand UO_1942 (O_1942,N_14250,N_12953);
xnor UO_1943 (O_1943,N_12995,N_13602);
xor UO_1944 (O_1944,N_12139,N_14466);
xnor UO_1945 (O_1945,N_12730,N_13132);
nor UO_1946 (O_1946,N_12150,N_14742);
nand UO_1947 (O_1947,N_13843,N_13863);
and UO_1948 (O_1948,N_12971,N_13216);
xnor UO_1949 (O_1949,N_12439,N_12049);
xor UO_1950 (O_1950,N_13083,N_12362);
xnor UO_1951 (O_1951,N_14642,N_12746);
and UO_1952 (O_1952,N_13312,N_13602);
xnor UO_1953 (O_1953,N_13218,N_13939);
nor UO_1954 (O_1954,N_14961,N_12389);
nand UO_1955 (O_1955,N_13954,N_14779);
and UO_1956 (O_1956,N_14288,N_14038);
nor UO_1957 (O_1957,N_12176,N_12499);
and UO_1958 (O_1958,N_14883,N_12411);
nor UO_1959 (O_1959,N_14209,N_12552);
or UO_1960 (O_1960,N_12651,N_12585);
nor UO_1961 (O_1961,N_12284,N_14319);
nor UO_1962 (O_1962,N_14199,N_12155);
nand UO_1963 (O_1963,N_12991,N_13462);
xnor UO_1964 (O_1964,N_12717,N_14438);
nand UO_1965 (O_1965,N_14689,N_13707);
and UO_1966 (O_1966,N_12665,N_14208);
nor UO_1967 (O_1967,N_13948,N_13671);
nor UO_1968 (O_1968,N_12132,N_13309);
or UO_1969 (O_1969,N_12352,N_14986);
xnor UO_1970 (O_1970,N_12129,N_13347);
nand UO_1971 (O_1971,N_12783,N_12753);
or UO_1972 (O_1972,N_13095,N_12919);
and UO_1973 (O_1973,N_13300,N_12886);
and UO_1974 (O_1974,N_13229,N_14211);
and UO_1975 (O_1975,N_13985,N_14610);
or UO_1976 (O_1976,N_14708,N_14693);
and UO_1977 (O_1977,N_13290,N_12056);
or UO_1978 (O_1978,N_14709,N_12448);
and UO_1979 (O_1979,N_14080,N_12862);
xnor UO_1980 (O_1980,N_13491,N_12744);
nand UO_1981 (O_1981,N_13370,N_13172);
or UO_1982 (O_1982,N_14247,N_12599);
nor UO_1983 (O_1983,N_12368,N_12294);
nor UO_1984 (O_1984,N_14678,N_14549);
xnor UO_1985 (O_1985,N_12717,N_14324);
and UO_1986 (O_1986,N_14687,N_12857);
or UO_1987 (O_1987,N_12460,N_14414);
xor UO_1988 (O_1988,N_12962,N_14229);
nand UO_1989 (O_1989,N_12928,N_14112);
nand UO_1990 (O_1990,N_13346,N_13558);
nor UO_1991 (O_1991,N_13210,N_14357);
xor UO_1992 (O_1992,N_12171,N_14023);
nor UO_1993 (O_1993,N_14096,N_14011);
and UO_1994 (O_1994,N_14982,N_14933);
xor UO_1995 (O_1995,N_13853,N_12257);
nor UO_1996 (O_1996,N_13050,N_12046);
and UO_1997 (O_1997,N_12283,N_13511);
xor UO_1998 (O_1998,N_14692,N_12250);
xor UO_1999 (O_1999,N_14445,N_14225);
endmodule