module basic_750_5000_1000_25_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_345,In_27);
and U1 (N_1,In_463,In_662);
nand U2 (N_2,In_230,In_568);
xor U3 (N_3,In_421,In_563);
xnor U4 (N_4,In_613,In_212);
or U5 (N_5,In_469,In_665);
xnor U6 (N_6,In_497,In_521);
nand U7 (N_7,In_78,In_383);
nor U8 (N_8,In_475,In_362);
nand U9 (N_9,In_347,In_399);
nor U10 (N_10,In_446,In_524);
xnor U11 (N_11,In_645,In_299);
or U12 (N_12,In_151,In_242);
and U13 (N_13,In_710,In_107);
and U14 (N_14,In_20,In_92);
nand U15 (N_15,In_677,In_629);
and U16 (N_16,In_682,In_284);
nand U17 (N_17,In_19,In_402);
and U18 (N_18,In_360,In_201);
and U19 (N_19,In_684,In_44);
and U20 (N_20,In_105,In_511);
or U21 (N_21,In_174,In_584);
nor U22 (N_22,In_149,In_651);
nand U23 (N_23,In_1,In_24);
or U24 (N_24,In_111,In_11);
nand U25 (N_25,In_693,In_557);
nand U26 (N_26,In_398,In_198);
nor U27 (N_27,In_579,In_232);
nor U28 (N_28,In_413,In_499);
and U29 (N_29,In_466,In_354);
nor U30 (N_30,In_573,In_664);
or U31 (N_31,In_32,In_607);
xor U32 (N_32,In_372,In_575);
xor U33 (N_33,In_422,In_292);
or U34 (N_34,In_650,In_417);
and U35 (N_35,In_391,In_473);
nor U36 (N_36,In_685,In_88);
and U37 (N_37,In_535,In_635);
nor U38 (N_38,In_744,In_58);
nor U39 (N_39,In_28,In_152);
or U40 (N_40,In_386,In_236);
nand U41 (N_41,In_173,In_141);
xor U42 (N_42,In_237,In_87);
nand U43 (N_43,In_373,In_128);
nand U44 (N_44,In_130,In_14);
and U45 (N_45,In_458,In_508);
nor U46 (N_46,In_441,In_85);
or U47 (N_47,In_279,In_541);
nand U48 (N_48,In_51,In_135);
nor U49 (N_49,In_484,In_101);
or U50 (N_50,In_154,In_623);
nand U51 (N_51,In_226,In_95);
nor U52 (N_52,In_432,In_172);
nor U53 (N_53,In_660,In_104);
and U54 (N_54,In_216,In_166);
nand U55 (N_55,In_487,In_206);
nand U56 (N_56,In_289,In_86);
nand U57 (N_57,In_246,In_516);
nor U58 (N_58,In_145,In_188);
nor U59 (N_59,In_280,In_559);
or U60 (N_60,In_334,In_674);
nand U61 (N_61,In_640,In_83);
nor U62 (N_62,In_72,In_668);
or U63 (N_63,In_631,In_435);
and U64 (N_64,In_381,In_504);
nor U65 (N_65,In_118,In_702);
nand U66 (N_66,In_439,In_102);
nand U67 (N_67,In_15,In_453);
xnor U68 (N_68,In_485,In_672);
and U69 (N_69,In_218,In_633);
or U70 (N_70,In_554,In_278);
nand U71 (N_71,In_461,In_61);
xor U72 (N_72,In_468,In_319);
nor U73 (N_73,In_715,In_133);
nor U74 (N_74,In_594,In_273);
xnor U75 (N_75,In_711,In_643);
or U76 (N_76,In_690,In_156);
xnor U77 (N_77,In_610,In_178);
nor U78 (N_78,In_163,In_308);
nand U79 (N_79,In_406,In_423);
nor U80 (N_80,In_555,In_55);
xnor U81 (N_81,In_531,In_371);
and U82 (N_82,In_519,In_222);
xnor U83 (N_83,In_729,In_731);
nand U84 (N_84,In_300,In_169);
xor U85 (N_85,In_175,In_727);
nand U86 (N_86,In_472,In_349);
or U87 (N_87,In_726,In_3);
nand U88 (N_88,In_530,In_109);
nor U89 (N_89,In_460,In_164);
or U90 (N_90,In_741,In_589);
xnor U91 (N_91,In_408,In_36);
and U92 (N_92,In_29,In_140);
or U93 (N_93,In_696,In_125);
xnor U94 (N_94,In_316,In_547);
or U95 (N_95,In_712,In_286);
and U96 (N_96,In_50,In_378);
xnor U97 (N_97,In_576,In_407);
and U98 (N_98,In_126,In_621);
xnor U99 (N_99,In_127,In_517);
or U100 (N_100,In_444,In_411);
or U101 (N_101,In_553,In_352);
and U102 (N_102,In_46,In_358);
nand U103 (N_103,In_550,In_196);
or U104 (N_104,In_64,In_596);
or U105 (N_105,In_646,In_18);
nand U106 (N_106,In_170,In_745);
or U107 (N_107,In_90,In_619);
xnor U108 (N_108,In_561,In_418);
and U109 (N_109,In_681,In_388);
nor U110 (N_110,In_467,In_687);
nand U111 (N_111,In_451,In_338);
nor U112 (N_112,In_197,In_121);
and U113 (N_113,In_428,In_134);
and U114 (N_114,In_106,In_235);
nor U115 (N_115,In_743,In_722);
and U116 (N_116,In_179,In_243);
xnor U117 (N_117,In_602,In_65);
nand U118 (N_118,In_510,In_48);
and U119 (N_119,In_671,In_502);
xor U120 (N_120,In_465,In_481);
and U121 (N_121,In_720,In_120);
xnor U122 (N_122,In_666,In_483);
and U123 (N_123,In_667,In_476);
or U124 (N_124,In_454,In_207);
nor U125 (N_125,In_13,In_43);
nor U126 (N_126,In_376,In_260);
xor U127 (N_127,In_479,In_507);
nand U128 (N_128,In_57,In_414);
or U129 (N_129,In_425,In_724);
xnor U130 (N_130,In_182,In_480);
and U131 (N_131,In_678,In_582);
nand U132 (N_132,In_336,In_612);
or U133 (N_133,In_269,In_447);
or U134 (N_134,In_513,In_644);
and U135 (N_135,In_737,In_259);
or U136 (N_136,In_551,In_112);
xnor U137 (N_137,In_309,In_449);
or U138 (N_138,In_37,In_210);
nor U139 (N_139,In_276,In_529);
nand U140 (N_140,In_180,In_272);
and U141 (N_141,In_137,In_296);
or U142 (N_142,In_658,In_302);
nor U143 (N_143,In_615,In_231);
and U144 (N_144,In_735,In_108);
and U145 (N_145,In_680,In_177);
and U146 (N_146,In_41,In_464);
or U147 (N_147,In_605,In_515);
or U148 (N_148,In_361,In_325);
xnor U149 (N_149,In_698,In_244);
xor U150 (N_150,In_369,In_520);
xor U151 (N_151,In_707,In_62);
nand U152 (N_152,In_628,In_368);
xor U153 (N_153,In_670,In_478);
xnor U154 (N_154,In_5,In_740);
and U155 (N_155,In_595,In_155);
or U156 (N_156,In_601,In_241);
and U157 (N_157,In_733,In_139);
nor U158 (N_158,In_367,In_614);
and U159 (N_159,In_689,In_144);
xor U160 (N_160,In_291,In_574);
and U161 (N_161,In_717,In_459);
nor U162 (N_162,In_654,In_70);
nor U163 (N_163,In_305,In_626);
or U164 (N_164,In_355,In_387);
or U165 (N_165,In_577,In_617);
or U166 (N_166,In_208,In_527);
or U167 (N_167,In_142,In_719);
nor U168 (N_168,In_686,In_195);
or U169 (N_169,In_431,In_375);
nor U170 (N_170,In_624,In_749);
nand U171 (N_171,In_138,In_136);
xnor U172 (N_172,In_405,In_514);
xor U173 (N_173,In_307,In_190);
nor U174 (N_174,In_694,In_618);
and U175 (N_175,In_63,In_641);
or U176 (N_176,In_22,In_160);
xor U177 (N_177,In_56,In_261);
nor U178 (N_178,In_709,In_565);
xor U179 (N_179,In_616,In_462);
and U180 (N_180,In_233,In_181);
or U181 (N_181,In_66,In_448);
nor U182 (N_182,In_60,In_593);
nand U183 (N_183,In_532,In_587);
or U184 (N_184,In_346,In_7);
nand U185 (N_185,In_171,In_608);
and U186 (N_186,In_627,In_159);
and U187 (N_187,In_489,In_42);
or U188 (N_188,In_390,In_192);
xnor U189 (N_189,In_385,In_253);
or U190 (N_190,In_298,In_572);
xnor U191 (N_191,In_430,In_730);
and U192 (N_192,In_500,In_6);
xor U193 (N_193,In_114,In_239);
nor U194 (N_194,In_31,In_89);
and U195 (N_195,In_247,In_321);
nand U196 (N_196,In_539,In_200);
or U197 (N_197,In_392,In_356);
or U198 (N_198,In_229,In_320);
and U199 (N_199,In_679,In_315);
xor U200 (N_200,In_675,N_20);
nand U201 (N_201,In_204,N_180);
or U202 (N_202,N_114,In_344);
nand U203 (N_203,In_442,In_688);
and U204 (N_204,N_63,N_132);
and U205 (N_205,N_17,N_15);
nor U206 (N_206,In_611,In_676);
nand U207 (N_207,N_83,In_395);
xor U208 (N_208,In_124,N_98);
and U209 (N_209,N_172,In_317);
xnor U210 (N_210,In_556,In_116);
or U211 (N_211,In_223,In_394);
or U212 (N_212,In_161,N_175);
and U213 (N_213,N_141,N_120);
nor U214 (N_214,In_419,N_152);
and U215 (N_215,N_148,N_106);
and U216 (N_216,In_68,N_84);
xor U217 (N_217,In_438,In_267);
or U218 (N_218,In_420,In_49);
nor U219 (N_219,In_343,N_57);
nand U220 (N_220,N_27,In_477);
or U221 (N_221,In_429,N_131);
nor U222 (N_222,In_377,In_331);
and U223 (N_223,N_121,In_93);
xor U224 (N_224,In_250,In_512);
nor U225 (N_225,In_290,In_552);
or U226 (N_226,In_739,In_283);
nor U227 (N_227,N_3,In_488);
or U228 (N_228,In_115,In_498);
and U229 (N_229,In_40,In_699);
or U230 (N_230,N_110,In_379);
or U231 (N_231,In_363,In_692);
nand U232 (N_232,N_64,N_16);
and U233 (N_233,In_545,N_72);
xnor U234 (N_234,In_725,In_184);
nand U235 (N_235,In_673,In_25);
or U236 (N_236,In_220,N_30);
xor U237 (N_237,In_509,In_585);
nor U238 (N_238,In_205,N_52);
and U239 (N_239,N_176,N_48);
or U240 (N_240,In_649,N_150);
nor U241 (N_241,In_523,In_491);
nor U242 (N_242,In_191,N_71);
nor U243 (N_243,In_323,In_380);
nand U244 (N_244,In_281,In_546);
or U245 (N_245,In_224,In_490);
and U246 (N_246,In_333,N_80);
nor U247 (N_247,N_94,N_164);
nor U248 (N_248,In_94,N_143);
nor U249 (N_249,In_562,In_303);
and U250 (N_250,N_12,N_142);
nor U251 (N_251,In_301,In_187);
and U252 (N_252,In_350,In_400);
nand U253 (N_253,In_452,N_195);
nor U254 (N_254,In_282,In_410);
and U255 (N_255,N_101,In_322);
xor U256 (N_256,N_185,In_211);
xnor U257 (N_257,N_69,In_738);
and U258 (N_258,In_364,In_30);
or U259 (N_259,N_128,N_134);
nand U260 (N_260,N_22,In_549);
nand U261 (N_261,In_332,N_7);
or U262 (N_262,In_294,N_13);
xor U263 (N_263,In_73,N_187);
and U264 (N_264,In_655,N_79);
or U265 (N_265,In_630,In_560);
nand U266 (N_266,In_648,In_382);
nand U267 (N_267,In_374,In_335);
and U268 (N_268,N_129,In_625);
nand U269 (N_269,N_29,N_158);
nand U270 (N_270,N_124,N_100);
nor U271 (N_271,In_647,In_157);
xor U272 (N_272,In_74,In_277);
nor U273 (N_273,In_393,In_96);
nor U274 (N_274,N_126,In_34);
and U275 (N_275,In_455,In_493);
nand U276 (N_276,In_311,In_580);
or U277 (N_277,In_203,In_401);
xor U278 (N_278,N_51,In_569);
nand U279 (N_279,In_251,N_138);
nand U280 (N_280,In_2,In_21);
or U281 (N_281,In_501,N_167);
and U282 (N_282,In_265,In_295);
xor U283 (N_283,In_548,N_97);
nand U284 (N_284,In_657,N_44);
nand U285 (N_285,N_58,In_606);
nor U286 (N_286,In_132,In_542);
or U287 (N_287,In_217,In_110);
xor U288 (N_288,N_39,N_105);
nand U289 (N_289,N_122,N_75);
nor U290 (N_290,In_586,In_570);
nor U291 (N_291,In_71,In_306);
xnor U292 (N_292,N_25,N_65);
xor U293 (N_293,In_100,In_409);
xnor U294 (N_294,N_23,In_59);
nor U295 (N_295,N_137,N_36);
xor U296 (N_296,In_456,In_701);
xnor U297 (N_297,N_171,N_118);
xnor U298 (N_298,N_41,N_181);
nand U299 (N_299,N_192,In_540);
nor U300 (N_300,N_144,In_470);
xor U301 (N_301,In_434,N_182);
nor U302 (N_302,N_91,N_43);
and U303 (N_303,N_61,In_91);
nand U304 (N_304,N_32,In_329);
and U305 (N_305,N_189,N_55);
or U306 (N_306,N_37,In_318);
nor U307 (N_307,In_0,N_145);
and U308 (N_308,In_708,In_264);
nor U309 (N_309,In_440,N_6);
or U310 (N_310,In_474,In_543);
or U311 (N_311,In_638,In_496);
and U312 (N_312,In_167,In_297);
or U313 (N_313,In_162,In_252);
nor U314 (N_314,N_165,In_656);
and U315 (N_315,N_0,In_69);
or U316 (N_316,In_486,In_661);
nand U317 (N_317,N_11,In_370);
or U318 (N_318,N_92,In_691);
and U319 (N_319,N_113,N_59);
xnor U320 (N_320,In_82,In_443);
xnor U321 (N_321,N_197,N_170);
or U322 (N_322,In_716,In_12);
nand U323 (N_323,N_35,In_683);
xor U324 (N_324,In_634,In_129);
or U325 (N_325,In_35,In_457);
or U326 (N_326,N_188,In_518);
nand U327 (N_327,In_695,N_166);
and U328 (N_328,N_4,In_590);
and U329 (N_329,N_31,In_52);
xnor U330 (N_330,N_66,N_90);
xnor U331 (N_331,In_592,In_33);
and U332 (N_332,In_122,In_193);
and U333 (N_333,In_718,In_471);
and U334 (N_334,In_526,N_42);
xnor U335 (N_335,N_46,In_598);
xnor U336 (N_336,In_39,In_494);
nand U337 (N_337,In_536,In_505);
nand U338 (N_338,In_669,N_136);
xnor U339 (N_339,N_111,In_351);
or U340 (N_340,In_81,In_285);
nand U341 (N_341,In_10,N_178);
xor U342 (N_342,In_412,In_274);
or U343 (N_343,In_38,In_597);
or U344 (N_344,N_9,In_143);
nor U345 (N_345,N_47,In_583);
xor U346 (N_346,N_45,N_140);
xnor U347 (N_347,In_533,In_26);
and U348 (N_348,In_482,In_703);
and U349 (N_349,In_357,N_168);
and U350 (N_350,In_150,In_734);
nor U351 (N_351,In_433,N_119);
or U352 (N_352,In_353,In_245);
or U353 (N_353,In_45,In_339);
xnor U354 (N_354,N_40,In_263);
or U355 (N_355,N_85,In_266);
nand U356 (N_356,In_248,In_544);
and U357 (N_357,In_148,In_249);
nor U358 (N_358,In_700,N_50);
nand U359 (N_359,N_174,N_186);
nand U360 (N_360,In_168,N_70);
xor U361 (N_361,N_68,In_348);
xnor U362 (N_362,N_87,In_340);
nor U363 (N_363,N_82,In_704);
and U364 (N_364,In_564,N_160);
nand U365 (N_365,N_198,In_436);
or U366 (N_366,In_427,In_258);
nor U367 (N_367,N_67,In_47);
and U368 (N_368,N_157,N_56);
nand U369 (N_369,In_153,N_117);
nand U370 (N_370,N_155,In_659);
or U371 (N_371,In_310,In_209);
or U372 (N_372,N_112,In_271);
nand U373 (N_373,N_33,In_714);
xor U374 (N_374,N_8,N_123);
or U375 (N_375,In_77,In_99);
or U376 (N_376,In_23,In_341);
or U377 (N_377,N_151,In_642);
xnor U378 (N_378,In_663,In_558);
and U379 (N_379,In_604,In_599);
nor U380 (N_380,In_396,In_706);
and U381 (N_381,In_185,In_503);
nor U382 (N_382,N_177,In_76);
nand U383 (N_383,N_88,N_77);
nor U384 (N_384,In_653,In_293);
nor U385 (N_385,N_173,In_288);
nor U386 (N_386,N_21,In_238);
or U387 (N_387,N_73,N_1);
and U388 (N_388,In_98,In_256);
nor U389 (N_389,In_255,N_28);
and U390 (N_390,In_158,N_184);
nand U391 (N_391,In_537,In_365);
and U392 (N_392,N_18,In_213);
or U393 (N_393,N_149,In_326);
or U394 (N_394,N_179,N_146);
xnor U395 (N_395,N_89,In_747);
or U396 (N_396,In_637,N_26);
nor U397 (N_397,In_17,In_117);
nor U398 (N_398,In_591,N_163);
nand U399 (N_399,In_721,In_123);
or U400 (N_400,N_191,N_316);
nand U401 (N_401,N_78,N_34);
nand U402 (N_402,N_394,In_103);
xnor U403 (N_403,N_382,N_333);
nand U404 (N_404,N_398,N_127);
or U405 (N_405,In_609,In_84);
nand U406 (N_406,N_366,N_237);
and U407 (N_407,N_295,N_301);
nor U408 (N_408,In_732,N_246);
nor U409 (N_409,N_235,N_161);
xor U410 (N_410,N_232,N_102);
nand U411 (N_411,N_208,In_312);
and U412 (N_412,N_365,N_375);
nand U413 (N_413,In_522,N_24);
and U414 (N_414,In_257,N_213);
nand U415 (N_415,N_264,N_397);
or U416 (N_416,N_317,In_600);
and U417 (N_417,N_2,N_248);
nand U418 (N_418,N_388,In_403);
or U419 (N_419,In_525,N_153);
xnor U420 (N_420,N_247,N_254);
and U421 (N_421,N_368,N_202);
and U422 (N_422,N_193,N_271);
nand U423 (N_423,N_214,N_218);
nand U424 (N_424,N_362,N_351);
or U425 (N_425,N_199,N_139);
and U426 (N_426,N_399,N_269);
and U427 (N_427,In_622,N_305);
nand U428 (N_428,In_147,In_746);
and U429 (N_429,N_156,N_290);
and U430 (N_430,In_639,In_384);
xor U431 (N_431,N_86,N_81);
and U432 (N_432,N_201,N_336);
nand U433 (N_433,In_327,N_99);
and U434 (N_434,N_206,In_304);
nand U435 (N_435,N_209,N_328);
or U436 (N_436,N_133,In_54);
or U437 (N_437,N_329,In_404);
and U438 (N_438,N_183,N_357);
nand U439 (N_439,N_278,N_225);
xor U440 (N_440,N_342,In_221);
xor U441 (N_441,N_245,N_255);
nand U442 (N_442,N_284,N_346);
xnor U443 (N_443,In_748,N_341);
and U444 (N_444,N_239,N_349);
nand U445 (N_445,N_200,N_300);
xnor U446 (N_446,N_310,N_282);
nor U447 (N_447,In_270,In_254);
nor U448 (N_448,In_214,N_283);
nor U449 (N_449,N_240,In_697);
or U450 (N_450,In_506,N_261);
nand U451 (N_451,In_366,N_93);
nand U452 (N_452,In_342,N_306);
xnor U453 (N_453,N_391,N_147);
nor U454 (N_454,N_381,N_190);
xor U455 (N_455,N_315,In_16);
and U456 (N_456,In_571,N_376);
nand U457 (N_457,In_313,N_104);
and U458 (N_458,In_146,N_109);
nand U459 (N_459,N_49,N_277);
xnor U460 (N_460,N_262,N_258);
and U461 (N_461,N_211,In_119);
or U462 (N_462,N_249,In_189);
and U463 (N_463,N_224,N_294);
xnor U464 (N_464,In_652,In_225);
or U465 (N_465,N_361,N_108);
nand U466 (N_466,N_275,In_723);
xor U467 (N_467,In_415,In_534);
nand U468 (N_468,In_538,N_215);
or U469 (N_469,N_251,N_347);
nand U470 (N_470,In_9,N_386);
or U471 (N_471,N_267,N_221);
or U472 (N_472,In_330,In_736);
and U473 (N_473,N_266,N_228);
xor U474 (N_474,N_297,N_226);
xnor U475 (N_475,In_713,N_353);
or U476 (N_476,In_215,N_241);
or U477 (N_477,In_728,In_234);
xnor U478 (N_478,N_383,In_80);
nand U479 (N_479,N_169,N_393);
or U480 (N_480,N_270,N_319);
xnor U481 (N_481,N_358,In_227);
xor U482 (N_482,N_392,N_14);
nor U483 (N_483,N_325,N_345);
nand U484 (N_484,N_367,N_194);
xnor U485 (N_485,N_162,N_339);
or U486 (N_486,N_299,N_343);
or U487 (N_487,N_236,N_273);
and U488 (N_488,N_355,In_424);
nor U489 (N_489,N_115,N_396);
or U490 (N_490,N_116,N_304);
or U491 (N_491,In_131,N_260);
or U492 (N_492,N_356,N_332);
and U493 (N_493,N_203,In_578);
xnor U494 (N_494,N_287,N_242);
nand U495 (N_495,In_176,N_292);
and U496 (N_496,N_154,N_307);
nor U497 (N_497,N_288,In_359);
nand U498 (N_498,N_204,In_262);
xor U499 (N_499,In_199,N_289);
nor U500 (N_500,N_372,In_324);
and U501 (N_501,N_280,N_363);
nand U502 (N_502,N_370,N_373);
xnor U503 (N_503,In_566,In_275);
and U504 (N_504,N_60,N_318);
xor U505 (N_505,N_379,N_378);
nor U506 (N_506,N_377,N_107);
xor U507 (N_507,N_238,N_309);
or U508 (N_508,N_74,In_53);
xor U509 (N_509,N_229,N_308);
and U510 (N_510,N_395,N_389);
and U511 (N_511,N_354,N_265);
or U512 (N_512,N_387,N_380);
xor U513 (N_513,N_390,N_231);
and U514 (N_514,N_130,N_217);
xnor U515 (N_515,N_340,N_159);
nand U516 (N_516,N_281,In_219);
and U517 (N_517,In_8,In_437);
nand U518 (N_518,In_620,N_53);
and U519 (N_519,In_445,N_369);
and U520 (N_520,N_338,N_293);
nor U521 (N_521,N_125,N_272);
nor U522 (N_522,N_253,In_450);
or U523 (N_523,In_202,N_210);
xnor U524 (N_524,N_296,In_603);
nand U525 (N_525,In_194,N_298);
nand U526 (N_526,N_223,In_183);
nand U527 (N_527,In_287,N_359);
and U528 (N_528,In_567,N_303);
xnor U529 (N_529,N_220,In_186);
xor U530 (N_530,In_588,In_328);
nand U531 (N_531,In_426,N_360);
xor U532 (N_532,N_10,In_113);
or U533 (N_533,N_285,N_227);
nand U534 (N_534,N_313,In_97);
nor U535 (N_535,N_135,In_4);
nand U536 (N_536,N_103,In_705);
nor U537 (N_537,N_222,N_268);
nor U538 (N_538,N_38,N_196);
and U539 (N_539,N_62,In_495);
and U540 (N_540,N_302,N_311);
nor U541 (N_541,In_165,N_230);
nand U542 (N_542,N_233,N_385);
xnor U543 (N_543,N_374,N_352);
and U544 (N_544,N_279,In_75);
or U545 (N_545,N_337,In_581);
nand U546 (N_546,N_256,N_286);
nor U547 (N_547,N_364,In_240);
and U548 (N_548,In_742,N_276);
nand U549 (N_549,In_79,N_212);
nor U550 (N_550,N_320,N_257);
xor U551 (N_551,N_216,N_274);
and U552 (N_552,In_389,N_312);
and U553 (N_553,In_528,N_371);
nor U554 (N_554,N_95,In_416);
nor U555 (N_555,N_348,In_492);
or U556 (N_556,N_5,In_268);
nor U557 (N_557,N_327,N_243);
or U558 (N_558,N_326,N_76);
and U559 (N_559,In_67,N_323);
and U560 (N_560,In_636,N_259);
nand U561 (N_561,N_321,N_324);
nand U562 (N_562,N_334,N_322);
or U563 (N_563,In_228,N_207);
xor U564 (N_564,N_263,N_291);
xor U565 (N_565,N_219,In_314);
and U566 (N_566,N_234,N_205);
xnor U567 (N_567,N_96,N_54);
nor U568 (N_568,In_337,In_397);
nor U569 (N_569,N_19,N_250);
xor U570 (N_570,N_330,N_384);
nand U571 (N_571,In_632,N_350);
and U572 (N_572,N_344,N_314);
and U573 (N_573,N_252,N_244);
and U574 (N_574,N_331,N_335);
or U575 (N_575,In_327,N_311);
nor U576 (N_576,N_147,N_74);
or U577 (N_577,N_338,In_450);
nand U578 (N_578,N_204,In_415);
and U579 (N_579,In_538,In_254);
and U580 (N_580,N_222,N_249);
nand U581 (N_581,N_329,N_385);
and U582 (N_582,N_277,N_337);
nor U583 (N_583,N_220,In_194);
xnor U584 (N_584,In_342,N_243);
nand U585 (N_585,N_306,N_262);
or U586 (N_586,N_255,N_212);
and U587 (N_587,N_257,In_287);
or U588 (N_588,N_397,N_201);
xor U589 (N_589,N_337,N_393);
or U590 (N_590,N_103,N_162);
xnor U591 (N_591,N_196,N_147);
or U592 (N_592,N_359,N_313);
or U593 (N_593,N_10,N_282);
nor U594 (N_594,N_391,N_325);
and U595 (N_595,N_60,In_337);
xnor U596 (N_596,N_243,N_139);
nor U597 (N_597,N_301,N_183);
nand U598 (N_598,N_359,N_265);
and U599 (N_599,N_273,N_281);
nor U600 (N_600,N_442,N_462);
and U601 (N_601,N_595,N_479);
and U602 (N_602,N_416,N_521);
nor U603 (N_603,N_443,N_512);
nand U604 (N_604,N_426,N_507);
and U605 (N_605,N_533,N_485);
and U606 (N_606,N_432,N_567);
nor U607 (N_607,N_536,N_434);
nand U608 (N_608,N_552,N_496);
nand U609 (N_609,N_464,N_486);
xnor U610 (N_610,N_548,N_408);
xor U611 (N_611,N_428,N_430);
nor U612 (N_612,N_580,N_534);
xor U613 (N_613,N_483,N_520);
xor U614 (N_614,N_578,N_519);
xor U615 (N_615,N_538,N_511);
and U616 (N_616,N_402,N_460);
xor U617 (N_617,N_414,N_475);
nor U618 (N_618,N_532,N_421);
and U619 (N_619,N_598,N_540);
nor U620 (N_620,N_524,N_557);
nand U621 (N_621,N_528,N_467);
nor U622 (N_622,N_570,N_410);
xnor U623 (N_623,N_597,N_400);
nand U624 (N_624,N_587,N_591);
xor U625 (N_625,N_456,N_499);
xnor U626 (N_626,N_541,N_546);
xor U627 (N_627,N_577,N_437);
or U628 (N_628,N_469,N_599);
nor U629 (N_629,N_427,N_504);
xor U630 (N_630,N_429,N_545);
xor U631 (N_631,N_470,N_482);
nand U632 (N_632,N_554,N_415);
nor U633 (N_633,N_560,N_586);
nor U634 (N_634,N_596,N_403);
or U635 (N_635,N_561,N_489);
or U636 (N_636,N_503,N_539);
and U637 (N_637,N_404,N_589);
and U638 (N_638,N_530,N_413);
or U639 (N_639,N_544,N_590);
and U640 (N_640,N_463,N_592);
xor U641 (N_641,N_488,N_465);
and U642 (N_642,N_478,N_529);
or U643 (N_643,N_472,N_518);
and U644 (N_644,N_436,N_461);
xor U645 (N_645,N_513,N_526);
nand U646 (N_646,N_502,N_508);
or U647 (N_647,N_446,N_471);
or U648 (N_648,N_517,N_498);
xnor U649 (N_649,N_571,N_459);
nand U650 (N_650,N_480,N_493);
or U651 (N_651,N_476,N_457);
and U652 (N_652,N_576,N_584);
and U653 (N_653,N_468,N_523);
xor U654 (N_654,N_553,N_494);
and U655 (N_655,N_455,N_531);
nor U656 (N_656,N_433,N_439);
nor U657 (N_657,N_477,N_565);
nor U658 (N_658,N_522,N_525);
or U659 (N_659,N_527,N_572);
xnor U660 (N_660,N_448,N_481);
nor U661 (N_661,N_491,N_558);
and U662 (N_662,N_420,N_581);
xnor U663 (N_663,N_407,N_445);
and U664 (N_664,N_506,N_458);
or U665 (N_665,N_438,N_564);
xor U666 (N_666,N_454,N_419);
or U667 (N_667,N_452,N_406);
xor U668 (N_668,N_422,N_490);
xor U669 (N_669,N_574,N_516);
nand U670 (N_670,N_515,N_543);
or U671 (N_671,N_431,N_492);
xnor U672 (N_672,N_555,N_514);
or U673 (N_673,N_568,N_409);
or U674 (N_674,N_487,N_435);
xnor U675 (N_675,N_417,N_542);
xnor U676 (N_676,N_451,N_405);
and U677 (N_677,N_550,N_474);
nand U678 (N_678,N_593,N_547);
nor U679 (N_679,N_453,N_575);
nor U680 (N_680,N_579,N_569);
xor U681 (N_681,N_444,N_423);
and U682 (N_682,N_424,N_509);
and U683 (N_683,N_441,N_412);
nand U684 (N_684,N_501,N_497);
or U685 (N_685,N_450,N_537);
or U686 (N_686,N_401,N_440);
xor U687 (N_687,N_449,N_563);
or U688 (N_688,N_556,N_585);
or U689 (N_689,N_573,N_582);
nand U690 (N_690,N_500,N_559);
or U691 (N_691,N_594,N_505);
or U692 (N_692,N_535,N_562);
and U693 (N_693,N_411,N_484);
and U694 (N_694,N_588,N_495);
nand U695 (N_695,N_510,N_551);
or U696 (N_696,N_583,N_447);
or U697 (N_697,N_549,N_425);
and U698 (N_698,N_466,N_566);
nand U699 (N_699,N_418,N_473);
nand U700 (N_700,N_548,N_574);
and U701 (N_701,N_470,N_407);
nand U702 (N_702,N_568,N_435);
nand U703 (N_703,N_534,N_450);
xnor U704 (N_704,N_437,N_486);
and U705 (N_705,N_470,N_579);
nor U706 (N_706,N_449,N_425);
nand U707 (N_707,N_546,N_588);
and U708 (N_708,N_437,N_510);
and U709 (N_709,N_425,N_530);
or U710 (N_710,N_432,N_541);
and U711 (N_711,N_425,N_528);
nor U712 (N_712,N_445,N_547);
or U713 (N_713,N_480,N_437);
or U714 (N_714,N_494,N_578);
xnor U715 (N_715,N_540,N_511);
or U716 (N_716,N_431,N_468);
and U717 (N_717,N_468,N_564);
or U718 (N_718,N_585,N_599);
or U719 (N_719,N_525,N_422);
and U720 (N_720,N_502,N_461);
nand U721 (N_721,N_497,N_426);
nand U722 (N_722,N_402,N_494);
or U723 (N_723,N_400,N_474);
nor U724 (N_724,N_432,N_502);
or U725 (N_725,N_445,N_403);
nand U726 (N_726,N_410,N_459);
nand U727 (N_727,N_589,N_450);
nand U728 (N_728,N_491,N_460);
xnor U729 (N_729,N_405,N_500);
nand U730 (N_730,N_591,N_584);
nand U731 (N_731,N_519,N_508);
xor U732 (N_732,N_552,N_542);
nand U733 (N_733,N_555,N_408);
nand U734 (N_734,N_599,N_488);
or U735 (N_735,N_498,N_526);
and U736 (N_736,N_598,N_562);
nor U737 (N_737,N_537,N_557);
or U738 (N_738,N_413,N_557);
and U739 (N_739,N_460,N_538);
xor U740 (N_740,N_494,N_409);
xor U741 (N_741,N_530,N_591);
nor U742 (N_742,N_516,N_482);
or U743 (N_743,N_466,N_435);
nor U744 (N_744,N_429,N_521);
nand U745 (N_745,N_470,N_522);
nor U746 (N_746,N_487,N_449);
xnor U747 (N_747,N_442,N_516);
nor U748 (N_748,N_453,N_484);
xor U749 (N_749,N_570,N_411);
nor U750 (N_750,N_546,N_419);
or U751 (N_751,N_433,N_571);
or U752 (N_752,N_570,N_481);
xnor U753 (N_753,N_510,N_462);
or U754 (N_754,N_580,N_402);
or U755 (N_755,N_402,N_503);
xnor U756 (N_756,N_507,N_519);
nor U757 (N_757,N_401,N_526);
nand U758 (N_758,N_436,N_559);
or U759 (N_759,N_468,N_410);
or U760 (N_760,N_432,N_479);
or U761 (N_761,N_402,N_576);
or U762 (N_762,N_518,N_400);
or U763 (N_763,N_406,N_440);
or U764 (N_764,N_421,N_552);
nor U765 (N_765,N_578,N_434);
nand U766 (N_766,N_448,N_526);
nor U767 (N_767,N_554,N_470);
nor U768 (N_768,N_537,N_439);
nand U769 (N_769,N_569,N_436);
or U770 (N_770,N_505,N_419);
or U771 (N_771,N_536,N_410);
xnor U772 (N_772,N_548,N_427);
nand U773 (N_773,N_570,N_463);
nor U774 (N_774,N_454,N_455);
nor U775 (N_775,N_482,N_502);
and U776 (N_776,N_500,N_574);
nand U777 (N_777,N_516,N_441);
xor U778 (N_778,N_400,N_504);
nand U779 (N_779,N_501,N_407);
nand U780 (N_780,N_577,N_461);
and U781 (N_781,N_480,N_403);
nor U782 (N_782,N_595,N_411);
and U783 (N_783,N_426,N_533);
xnor U784 (N_784,N_555,N_530);
nand U785 (N_785,N_541,N_539);
nor U786 (N_786,N_522,N_465);
nor U787 (N_787,N_467,N_486);
or U788 (N_788,N_535,N_481);
and U789 (N_789,N_430,N_460);
xnor U790 (N_790,N_409,N_515);
and U791 (N_791,N_440,N_425);
nand U792 (N_792,N_571,N_483);
xnor U793 (N_793,N_472,N_584);
or U794 (N_794,N_533,N_470);
and U795 (N_795,N_572,N_487);
nor U796 (N_796,N_408,N_534);
and U797 (N_797,N_448,N_594);
nand U798 (N_798,N_582,N_596);
nand U799 (N_799,N_583,N_541);
xnor U800 (N_800,N_636,N_650);
and U801 (N_801,N_793,N_656);
nor U802 (N_802,N_757,N_640);
and U803 (N_803,N_672,N_699);
or U804 (N_804,N_771,N_719);
or U805 (N_805,N_775,N_697);
nor U806 (N_806,N_609,N_622);
nand U807 (N_807,N_729,N_683);
nand U808 (N_808,N_692,N_624);
nand U809 (N_809,N_687,N_666);
or U810 (N_810,N_694,N_711);
nand U811 (N_811,N_614,N_628);
or U812 (N_812,N_788,N_710);
xor U813 (N_813,N_668,N_727);
xnor U814 (N_814,N_642,N_705);
xnor U815 (N_815,N_600,N_635);
and U816 (N_816,N_619,N_760);
and U817 (N_817,N_654,N_723);
nor U818 (N_818,N_772,N_756);
and U819 (N_819,N_799,N_753);
nand U820 (N_820,N_709,N_610);
nor U821 (N_821,N_626,N_603);
nor U822 (N_822,N_637,N_716);
nand U823 (N_823,N_707,N_789);
nand U824 (N_824,N_746,N_728);
and U825 (N_825,N_665,N_675);
xor U826 (N_826,N_648,N_620);
nand U827 (N_827,N_734,N_673);
nor U828 (N_828,N_611,N_726);
or U829 (N_829,N_782,N_632);
xor U830 (N_830,N_752,N_744);
xor U831 (N_831,N_661,N_747);
or U832 (N_832,N_688,N_651);
xnor U833 (N_833,N_693,N_731);
xor U834 (N_834,N_777,N_704);
nor U835 (N_835,N_745,N_759);
xor U836 (N_836,N_794,N_714);
xnor U837 (N_837,N_658,N_778);
and U838 (N_838,N_741,N_766);
nand U839 (N_839,N_669,N_680);
nand U840 (N_840,N_722,N_779);
nor U841 (N_841,N_781,N_743);
or U842 (N_842,N_674,N_717);
and U843 (N_843,N_769,N_682);
and U844 (N_844,N_662,N_618);
nand U845 (N_845,N_736,N_602);
nor U846 (N_846,N_670,N_718);
or U847 (N_847,N_715,N_671);
xor U848 (N_848,N_785,N_627);
xnor U849 (N_849,N_787,N_708);
nor U850 (N_850,N_767,N_617);
xor U851 (N_851,N_703,N_677);
nor U852 (N_852,N_604,N_733);
or U853 (N_853,N_724,N_612);
and U854 (N_854,N_681,N_738);
or U855 (N_855,N_795,N_712);
nand U856 (N_856,N_647,N_786);
nor U857 (N_857,N_623,N_780);
nor U858 (N_858,N_601,N_755);
and U859 (N_859,N_659,N_700);
and U860 (N_860,N_737,N_685);
xor U861 (N_861,N_639,N_770);
xnor U862 (N_862,N_606,N_657);
or U863 (N_863,N_792,N_638);
nand U864 (N_864,N_776,N_684);
and U865 (N_865,N_740,N_652);
and U866 (N_866,N_720,N_774);
or U867 (N_867,N_689,N_748);
or U868 (N_868,N_631,N_633);
nand U869 (N_869,N_691,N_725);
and U870 (N_870,N_754,N_653);
nor U871 (N_871,N_762,N_742);
and U872 (N_872,N_784,N_645);
nor U873 (N_873,N_765,N_798);
nand U874 (N_874,N_695,N_615);
xnor U875 (N_875,N_750,N_732);
or U876 (N_876,N_679,N_616);
nand U877 (N_877,N_749,N_678);
xor U878 (N_878,N_644,N_758);
xor U879 (N_879,N_721,N_646);
xnor U880 (N_880,N_796,N_706);
xor U881 (N_881,N_751,N_613);
xor U882 (N_882,N_797,N_768);
xnor U883 (N_883,N_655,N_764);
xor U884 (N_884,N_791,N_713);
nor U885 (N_885,N_625,N_739);
xnor U886 (N_886,N_663,N_763);
nor U887 (N_887,N_630,N_761);
nor U888 (N_888,N_735,N_667);
or U889 (N_889,N_701,N_608);
and U890 (N_890,N_773,N_641);
nand U891 (N_891,N_702,N_698);
nand U892 (N_892,N_676,N_730);
and U893 (N_893,N_605,N_607);
and U894 (N_894,N_790,N_783);
nand U895 (N_895,N_621,N_686);
xnor U896 (N_896,N_634,N_643);
and U897 (N_897,N_629,N_660);
xnor U898 (N_898,N_649,N_696);
nor U899 (N_899,N_664,N_690);
and U900 (N_900,N_779,N_798);
or U901 (N_901,N_695,N_682);
nand U902 (N_902,N_682,N_699);
nand U903 (N_903,N_766,N_680);
or U904 (N_904,N_638,N_761);
and U905 (N_905,N_659,N_628);
xnor U906 (N_906,N_734,N_661);
and U907 (N_907,N_778,N_667);
or U908 (N_908,N_693,N_795);
nor U909 (N_909,N_722,N_669);
xnor U910 (N_910,N_683,N_709);
or U911 (N_911,N_799,N_632);
or U912 (N_912,N_689,N_606);
and U913 (N_913,N_620,N_614);
nand U914 (N_914,N_636,N_632);
nor U915 (N_915,N_646,N_774);
nor U916 (N_916,N_697,N_619);
or U917 (N_917,N_685,N_726);
and U918 (N_918,N_670,N_784);
nand U919 (N_919,N_750,N_745);
nor U920 (N_920,N_623,N_668);
nor U921 (N_921,N_730,N_615);
nor U922 (N_922,N_612,N_735);
nor U923 (N_923,N_645,N_679);
nand U924 (N_924,N_725,N_610);
or U925 (N_925,N_671,N_606);
and U926 (N_926,N_607,N_627);
and U927 (N_927,N_771,N_797);
and U928 (N_928,N_667,N_740);
and U929 (N_929,N_659,N_600);
or U930 (N_930,N_661,N_785);
nor U931 (N_931,N_783,N_620);
or U932 (N_932,N_704,N_661);
xor U933 (N_933,N_698,N_613);
and U934 (N_934,N_687,N_752);
or U935 (N_935,N_735,N_600);
xnor U936 (N_936,N_787,N_737);
xor U937 (N_937,N_605,N_697);
nand U938 (N_938,N_756,N_604);
nor U939 (N_939,N_652,N_680);
and U940 (N_940,N_722,N_751);
nand U941 (N_941,N_645,N_707);
and U942 (N_942,N_699,N_732);
xor U943 (N_943,N_619,N_787);
nand U944 (N_944,N_788,N_740);
and U945 (N_945,N_775,N_623);
xnor U946 (N_946,N_773,N_662);
nor U947 (N_947,N_740,N_683);
nor U948 (N_948,N_662,N_628);
nand U949 (N_949,N_629,N_783);
xnor U950 (N_950,N_653,N_713);
nor U951 (N_951,N_659,N_611);
or U952 (N_952,N_790,N_625);
and U953 (N_953,N_775,N_631);
and U954 (N_954,N_669,N_789);
xor U955 (N_955,N_607,N_781);
and U956 (N_956,N_656,N_657);
xnor U957 (N_957,N_794,N_604);
or U958 (N_958,N_654,N_743);
nor U959 (N_959,N_696,N_791);
or U960 (N_960,N_726,N_792);
nand U961 (N_961,N_704,N_647);
or U962 (N_962,N_767,N_613);
nand U963 (N_963,N_710,N_650);
nand U964 (N_964,N_656,N_786);
nor U965 (N_965,N_795,N_684);
nand U966 (N_966,N_763,N_764);
and U967 (N_967,N_705,N_619);
or U968 (N_968,N_617,N_678);
and U969 (N_969,N_621,N_798);
or U970 (N_970,N_634,N_749);
or U971 (N_971,N_769,N_661);
nor U972 (N_972,N_741,N_795);
nor U973 (N_973,N_730,N_758);
nor U974 (N_974,N_646,N_793);
nand U975 (N_975,N_699,N_779);
nor U976 (N_976,N_662,N_626);
or U977 (N_977,N_663,N_721);
or U978 (N_978,N_745,N_761);
and U979 (N_979,N_690,N_622);
xnor U980 (N_980,N_698,N_720);
and U981 (N_981,N_643,N_796);
nand U982 (N_982,N_771,N_699);
nand U983 (N_983,N_724,N_722);
xor U984 (N_984,N_670,N_797);
nand U985 (N_985,N_793,N_745);
nor U986 (N_986,N_758,N_763);
xor U987 (N_987,N_670,N_633);
and U988 (N_988,N_693,N_606);
nor U989 (N_989,N_666,N_749);
nor U990 (N_990,N_601,N_736);
nor U991 (N_991,N_736,N_628);
nand U992 (N_992,N_716,N_730);
or U993 (N_993,N_740,N_607);
and U994 (N_994,N_644,N_754);
or U995 (N_995,N_686,N_778);
nand U996 (N_996,N_655,N_711);
or U997 (N_997,N_604,N_627);
nand U998 (N_998,N_609,N_753);
or U999 (N_999,N_708,N_740);
or U1000 (N_1000,N_885,N_848);
nor U1001 (N_1001,N_949,N_906);
and U1002 (N_1002,N_995,N_800);
and U1003 (N_1003,N_965,N_975);
nor U1004 (N_1004,N_991,N_887);
and U1005 (N_1005,N_875,N_942);
xnor U1006 (N_1006,N_916,N_921);
xnor U1007 (N_1007,N_805,N_928);
nand U1008 (N_1008,N_852,N_815);
nand U1009 (N_1009,N_972,N_857);
and U1010 (N_1010,N_934,N_951);
nor U1011 (N_1011,N_827,N_854);
nand U1012 (N_1012,N_826,N_806);
nand U1013 (N_1013,N_859,N_932);
xnor U1014 (N_1014,N_862,N_985);
or U1015 (N_1015,N_869,N_894);
and U1016 (N_1016,N_924,N_835);
or U1017 (N_1017,N_858,N_816);
nand U1018 (N_1018,N_809,N_962);
or U1019 (N_1019,N_823,N_819);
and U1020 (N_1020,N_856,N_967);
or U1021 (N_1021,N_879,N_970);
nand U1022 (N_1022,N_910,N_804);
or U1023 (N_1023,N_944,N_919);
and U1024 (N_1024,N_867,N_889);
xor U1025 (N_1025,N_918,N_878);
or U1026 (N_1026,N_981,N_898);
or U1027 (N_1027,N_801,N_820);
nor U1028 (N_1028,N_930,N_987);
nor U1029 (N_1029,N_983,N_956);
xor U1030 (N_1030,N_937,N_817);
nor U1031 (N_1031,N_813,N_912);
or U1032 (N_1032,N_873,N_834);
nor U1033 (N_1033,N_824,N_973);
nor U1034 (N_1034,N_904,N_863);
nand U1035 (N_1035,N_832,N_961);
xor U1036 (N_1036,N_953,N_896);
and U1037 (N_1037,N_913,N_982);
nand U1038 (N_1038,N_957,N_901);
and U1039 (N_1039,N_855,N_812);
xnor U1040 (N_1040,N_980,N_891);
nand U1041 (N_1041,N_908,N_868);
nor U1042 (N_1042,N_971,N_948);
nand U1043 (N_1043,N_864,N_936);
xnor U1044 (N_1044,N_880,N_845);
nand U1045 (N_1045,N_977,N_939);
xnor U1046 (N_1046,N_844,N_822);
nand U1047 (N_1047,N_947,N_882);
nand U1048 (N_1048,N_935,N_940);
nor U1049 (N_1049,N_830,N_926);
xnor U1050 (N_1050,N_925,N_943);
or U1051 (N_1051,N_911,N_914);
and U1052 (N_1052,N_860,N_821);
xor U1053 (N_1053,N_841,N_802);
and U1054 (N_1054,N_984,N_900);
or U1055 (N_1055,N_960,N_853);
xnor U1056 (N_1056,N_994,N_877);
or U1057 (N_1057,N_883,N_837);
xnor U1058 (N_1058,N_838,N_950);
or U1059 (N_1059,N_974,N_907);
nor U1060 (N_1060,N_847,N_872);
xor U1061 (N_1061,N_811,N_929);
nor U1062 (N_1062,N_955,N_958);
or U1063 (N_1063,N_865,N_881);
or U1064 (N_1064,N_843,N_933);
xor U1065 (N_1065,N_979,N_976);
xor U1066 (N_1066,N_808,N_968);
nor U1067 (N_1067,N_861,N_902);
or U1068 (N_1068,N_818,N_836);
and U1069 (N_1069,N_825,N_897);
and U1070 (N_1070,N_874,N_903);
nor U1071 (N_1071,N_920,N_866);
or U1072 (N_1072,N_998,N_846);
and U1073 (N_1073,N_996,N_840);
xnor U1074 (N_1074,N_839,N_833);
xnor U1075 (N_1075,N_888,N_895);
nand U1076 (N_1076,N_807,N_923);
nand U1077 (N_1077,N_915,N_886);
nand U1078 (N_1078,N_990,N_952);
nand U1079 (N_1079,N_870,N_917);
xor U1080 (N_1080,N_892,N_810);
nor U1081 (N_1081,N_997,N_966);
or U1082 (N_1082,N_992,N_849);
or U1083 (N_1083,N_946,N_959);
nor U1084 (N_1084,N_941,N_803);
nor U1085 (N_1085,N_829,N_842);
nand U1086 (N_1086,N_988,N_890);
xor U1087 (N_1087,N_884,N_954);
or U1088 (N_1088,N_927,N_831);
or U1089 (N_1089,N_850,N_871);
or U1090 (N_1090,N_978,N_964);
xor U1091 (N_1091,N_876,N_938);
or U1092 (N_1092,N_905,N_909);
nor U1093 (N_1093,N_828,N_993);
or U1094 (N_1094,N_851,N_893);
nor U1095 (N_1095,N_999,N_931);
nor U1096 (N_1096,N_814,N_963);
and U1097 (N_1097,N_969,N_945);
or U1098 (N_1098,N_922,N_899);
nor U1099 (N_1099,N_986,N_989);
or U1100 (N_1100,N_810,N_991);
nor U1101 (N_1101,N_831,N_958);
and U1102 (N_1102,N_852,N_847);
xor U1103 (N_1103,N_830,N_953);
nand U1104 (N_1104,N_884,N_858);
and U1105 (N_1105,N_987,N_827);
nand U1106 (N_1106,N_829,N_865);
and U1107 (N_1107,N_930,N_840);
xor U1108 (N_1108,N_907,N_979);
nor U1109 (N_1109,N_961,N_837);
xor U1110 (N_1110,N_863,N_867);
nand U1111 (N_1111,N_857,N_841);
xnor U1112 (N_1112,N_913,N_840);
or U1113 (N_1113,N_967,N_882);
and U1114 (N_1114,N_917,N_894);
nor U1115 (N_1115,N_811,N_915);
and U1116 (N_1116,N_800,N_945);
xor U1117 (N_1117,N_991,N_949);
or U1118 (N_1118,N_931,N_802);
xnor U1119 (N_1119,N_965,N_939);
xor U1120 (N_1120,N_902,N_829);
or U1121 (N_1121,N_820,N_894);
or U1122 (N_1122,N_925,N_893);
nand U1123 (N_1123,N_852,N_876);
or U1124 (N_1124,N_979,N_832);
nand U1125 (N_1125,N_978,N_827);
nor U1126 (N_1126,N_872,N_919);
nor U1127 (N_1127,N_902,N_881);
nand U1128 (N_1128,N_992,N_981);
and U1129 (N_1129,N_912,N_961);
nand U1130 (N_1130,N_912,N_836);
nor U1131 (N_1131,N_892,N_812);
nor U1132 (N_1132,N_835,N_958);
xnor U1133 (N_1133,N_802,N_886);
nor U1134 (N_1134,N_807,N_955);
and U1135 (N_1135,N_849,N_900);
nand U1136 (N_1136,N_971,N_957);
or U1137 (N_1137,N_959,N_920);
nor U1138 (N_1138,N_920,N_976);
nand U1139 (N_1139,N_933,N_847);
and U1140 (N_1140,N_951,N_847);
nor U1141 (N_1141,N_909,N_818);
or U1142 (N_1142,N_987,N_840);
and U1143 (N_1143,N_807,N_874);
and U1144 (N_1144,N_854,N_905);
xor U1145 (N_1145,N_865,N_887);
nand U1146 (N_1146,N_929,N_898);
and U1147 (N_1147,N_841,N_883);
nand U1148 (N_1148,N_920,N_990);
and U1149 (N_1149,N_871,N_948);
and U1150 (N_1150,N_805,N_849);
nor U1151 (N_1151,N_838,N_815);
and U1152 (N_1152,N_971,N_918);
nand U1153 (N_1153,N_889,N_963);
xnor U1154 (N_1154,N_814,N_990);
nor U1155 (N_1155,N_864,N_970);
xor U1156 (N_1156,N_896,N_865);
nand U1157 (N_1157,N_869,N_800);
or U1158 (N_1158,N_841,N_990);
and U1159 (N_1159,N_965,N_802);
nand U1160 (N_1160,N_880,N_843);
nor U1161 (N_1161,N_878,N_884);
xnor U1162 (N_1162,N_905,N_982);
xor U1163 (N_1163,N_888,N_837);
xor U1164 (N_1164,N_993,N_907);
or U1165 (N_1165,N_912,N_826);
xor U1166 (N_1166,N_943,N_951);
xnor U1167 (N_1167,N_840,N_917);
and U1168 (N_1168,N_855,N_965);
and U1169 (N_1169,N_959,N_883);
nor U1170 (N_1170,N_885,N_922);
xnor U1171 (N_1171,N_939,N_962);
or U1172 (N_1172,N_933,N_930);
nor U1173 (N_1173,N_918,N_854);
nand U1174 (N_1174,N_983,N_889);
nand U1175 (N_1175,N_884,N_914);
and U1176 (N_1176,N_823,N_868);
or U1177 (N_1177,N_929,N_889);
and U1178 (N_1178,N_829,N_931);
xor U1179 (N_1179,N_823,N_933);
nor U1180 (N_1180,N_953,N_998);
nand U1181 (N_1181,N_801,N_987);
and U1182 (N_1182,N_952,N_826);
xnor U1183 (N_1183,N_889,N_820);
xor U1184 (N_1184,N_940,N_863);
xor U1185 (N_1185,N_916,N_932);
nor U1186 (N_1186,N_955,N_838);
nand U1187 (N_1187,N_929,N_999);
nand U1188 (N_1188,N_882,N_837);
or U1189 (N_1189,N_846,N_908);
or U1190 (N_1190,N_894,N_870);
or U1191 (N_1191,N_925,N_973);
nor U1192 (N_1192,N_829,N_828);
or U1193 (N_1193,N_951,N_823);
nand U1194 (N_1194,N_821,N_994);
nor U1195 (N_1195,N_895,N_877);
nor U1196 (N_1196,N_823,N_884);
nand U1197 (N_1197,N_959,N_924);
or U1198 (N_1198,N_839,N_845);
and U1199 (N_1199,N_959,N_905);
nor U1200 (N_1200,N_1180,N_1117);
or U1201 (N_1201,N_1134,N_1061);
nand U1202 (N_1202,N_1078,N_1049);
nor U1203 (N_1203,N_1146,N_1142);
nand U1204 (N_1204,N_1056,N_1009);
or U1205 (N_1205,N_1114,N_1041);
xnor U1206 (N_1206,N_1034,N_1091);
or U1207 (N_1207,N_1193,N_1046);
nand U1208 (N_1208,N_1057,N_1015);
and U1209 (N_1209,N_1025,N_1069);
or U1210 (N_1210,N_1144,N_1075);
xnor U1211 (N_1211,N_1182,N_1135);
and U1212 (N_1212,N_1185,N_1095);
xor U1213 (N_1213,N_1068,N_1081);
or U1214 (N_1214,N_1123,N_1016);
and U1215 (N_1215,N_1048,N_1105);
nand U1216 (N_1216,N_1094,N_1108);
nand U1217 (N_1217,N_1151,N_1129);
and U1218 (N_1218,N_1179,N_1101);
or U1219 (N_1219,N_1098,N_1030);
or U1220 (N_1220,N_1058,N_1038);
nand U1221 (N_1221,N_1176,N_1191);
nor U1222 (N_1222,N_1197,N_1080);
nand U1223 (N_1223,N_1178,N_1171);
nor U1224 (N_1224,N_1089,N_1035);
nand U1225 (N_1225,N_1156,N_1195);
xor U1226 (N_1226,N_1163,N_1088);
nor U1227 (N_1227,N_1115,N_1065);
nor U1228 (N_1228,N_1116,N_1145);
xnor U1229 (N_1229,N_1196,N_1022);
nand U1230 (N_1230,N_1164,N_1152);
nand U1231 (N_1231,N_1063,N_1174);
nor U1232 (N_1232,N_1060,N_1050);
and U1233 (N_1233,N_1120,N_1059);
and U1234 (N_1234,N_1051,N_1138);
nor U1235 (N_1235,N_1067,N_1160);
xor U1236 (N_1236,N_1131,N_1132);
xor U1237 (N_1237,N_1012,N_1023);
xor U1238 (N_1238,N_1110,N_1155);
nand U1239 (N_1239,N_1024,N_1139);
xor U1240 (N_1240,N_1045,N_1079);
nand U1241 (N_1241,N_1148,N_1008);
nand U1242 (N_1242,N_1154,N_1177);
nor U1243 (N_1243,N_1136,N_1133);
nand U1244 (N_1244,N_1099,N_1021);
nand U1245 (N_1245,N_1149,N_1173);
xnor U1246 (N_1246,N_1143,N_1002);
nor U1247 (N_1247,N_1090,N_1162);
nor U1248 (N_1248,N_1052,N_1043);
nor U1249 (N_1249,N_1150,N_1175);
nor U1250 (N_1250,N_1082,N_1183);
nor U1251 (N_1251,N_1184,N_1104);
nand U1252 (N_1252,N_1181,N_1093);
xnor U1253 (N_1253,N_1198,N_1033);
or U1254 (N_1254,N_1077,N_1172);
nor U1255 (N_1255,N_1076,N_1085);
nor U1256 (N_1256,N_1070,N_1097);
nor U1257 (N_1257,N_1087,N_1014);
or U1258 (N_1258,N_1168,N_1188);
and U1259 (N_1259,N_1187,N_1125);
nor U1260 (N_1260,N_1096,N_1066);
nor U1261 (N_1261,N_1007,N_1031);
and U1262 (N_1262,N_1086,N_1055);
or U1263 (N_1263,N_1074,N_1161);
nor U1264 (N_1264,N_1199,N_1166);
or U1265 (N_1265,N_1062,N_1017);
nor U1266 (N_1266,N_1092,N_1040);
or U1267 (N_1267,N_1128,N_1137);
xor U1268 (N_1268,N_1140,N_1170);
and U1269 (N_1269,N_1032,N_1047);
xnor U1270 (N_1270,N_1126,N_1109);
or U1271 (N_1271,N_1053,N_1121);
xor U1272 (N_1272,N_1122,N_1000);
and U1273 (N_1273,N_1186,N_1039);
xor U1274 (N_1274,N_1141,N_1102);
xor U1275 (N_1275,N_1036,N_1165);
and U1276 (N_1276,N_1113,N_1127);
xor U1277 (N_1277,N_1073,N_1190);
xnor U1278 (N_1278,N_1071,N_1112);
and U1279 (N_1279,N_1083,N_1153);
or U1280 (N_1280,N_1027,N_1001);
and U1281 (N_1281,N_1169,N_1064);
and U1282 (N_1282,N_1189,N_1026);
nand U1283 (N_1283,N_1100,N_1072);
and U1284 (N_1284,N_1004,N_1192);
nor U1285 (N_1285,N_1167,N_1019);
nand U1286 (N_1286,N_1107,N_1159);
nand U1287 (N_1287,N_1119,N_1084);
and U1288 (N_1288,N_1010,N_1011);
or U1289 (N_1289,N_1020,N_1005);
and U1290 (N_1290,N_1103,N_1028);
nor U1291 (N_1291,N_1018,N_1006);
xor U1292 (N_1292,N_1124,N_1111);
nand U1293 (N_1293,N_1118,N_1106);
xnor U1294 (N_1294,N_1037,N_1013);
nand U1295 (N_1295,N_1147,N_1044);
nor U1296 (N_1296,N_1194,N_1157);
nor U1297 (N_1297,N_1029,N_1130);
xor U1298 (N_1298,N_1003,N_1158);
and U1299 (N_1299,N_1042,N_1054);
xnor U1300 (N_1300,N_1025,N_1186);
or U1301 (N_1301,N_1165,N_1060);
or U1302 (N_1302,N_1027,N_1137);
or U1303 (N_1303,N_1189,N_1038);
xor U1304 (N_1304,N_1157,N_1100);
or U1305 (N_1305,N_1056,N_1143);
nand U1306 (N_1306,N_1011,N_1135);
or U1307 (N_1307,N_1113,N_1050);
or U1308 (N_1308,N_1184,N_1025);
nand U1309 (N_1309,N_1012,N_1190);
xnor U1310 (N_1310,N_1169,N_1132);
nand U1311 (N_1311,N_1006,N_1091);
xor U1312 (N_1312,N_1143,N_1040);
xnor U1313 (N_1313,N_1026,N_1034);
nand U1314 (N_1314,N_1087,N_1089);
nor U1315 (N_1315,N_1005,N_1122);
nor U1316 (N_1316,N_1100,N_1014);
nor U1317 (N_1317,N_1016,N_1177);
or U1318 (N_1318,N_1017,N_1088);
nand U1319 (N_1319,N_1075,N_1009);
or U1320 (N_1320,N_1131,N_1010);
nand U1321 (N_1321,N_1023,N_1153);
xnor U1322 (N_1322,N_1062,N_1153);
nand U1323 (N_1323,N_1005,N_1051);
xor U1324 (N_1324,N_1131,N_1178);
or U1325 (N_1325,N_1173,N_1090);
nand U1326 (N_1326,N_1176,N_1125);
xnor U1327 (N_1327,N_1053,N_1168);
and U1328 (N_1328,N_1007,N_1195);
nand U1329 (N_1329,N_1147,N_1010);
nand U1330 (N_1330,N_1152,N_1089);
or U1331 (N_1331,N_1101,N_1036);
nor U1332 (N_1332,N_1049,N_1054);
and U1333 (N_1333,N_1164,N_1079);
xor U1334 (N_1334,N_1071,N_1029);
or U1335 (N_1335,N_1115,N_1136);
nor U1336 (N_1336,N_1134,N_1090);
nor U1337 (N_1337,N_1132,N_1157);
and U1338 (N_1338,N_1131,N_1161);
xor U1339 (N_1339,N_1121,N_1150);
and U1340 (N_1340,N_1025,N_1015);
and U1341 (N_1341,N_1133,N_1164);
and U1342 (N_1342,N_1173,N_1118);
xor U1343 (N_1343,N_1042,N_1198);
nand U1344 (N_1344,N_1174,N_1079);
or U1345 (N_1345,N_1047,N_1184);
xor U1346 (N_1346,N_1044,N_1017);
xnor U1347 (N_1347,N_1066,N_1149);
or U1348 (N_1348,N_1079,N_1099);
or U1349 (N_1349,N_1128,N_1022);
and U1350 (N_1350,N_1025,N_1188);
or U1351 (N_1351,N_1056,N_1109);
or U1352 (N_1352,N_1091,N_1194);
xnor U1353 (N_1353,N_1197,N_1188);
and U1354 (N_1354,N_1178,N_1157);
nand U1355 (N_1355,N_1175,N_1064);
or U1356 (N_1356,N_1151,N_1054);
nor U1357 (N_1357,N_1052,N_1037);
nor U1358 (N_1358,N_1040,N_1019);
xor U1359 (N_1359,N_1075,N_1084);
or U1360 (N_1360,N_1111,N_1073);
xor U1361 (N_1361,N_1025,N_1077);
nor U1362 (N_1362,N_1084,N_1064);
nor U1363 (N_1363,N_1067,N_1182);
nand U1364 (N_1364,N_1019,N_1191);
and U1365 (N_1365,N_1118,N_1042);
xor U1366 (N_1366,N_1072,N_1090);
nand U1367 (N_1367,N_1059,N_1135);
nor U1368 (N_1368,N_1106,N_1157);
nand U1369 (N_1369,N_1184,N_1068);
nand U1370 (N_1370,N_1107,N_1096);
xor U1371 (N_1371,N_1098,N_1059);
and U1372 (N_1372,N_1188,N_1030);
and U1373 (N_1373,N_1010,N_1024);
xor U1374 (N_1374,N_1152,N_1173);
nand U1375 (N_1375,N_1065,N_1088);
or U1376 (N_1376,N_1015,N_1062);
and U1377 (N_1377,N_1093,N_1107);
xor U1378 (N_1378,N_1184,N_1077);
or U1379 (N_1379,N_1168,N_1009);
nor U1380 (N_1380,N_1031,N_1191);
nand U1381 (N_1381,N_1059,N_1175);
or U1382 (N_1382,N_1000,N_1078);
or U1383 (N_1383,N_1146,N_1063);
and U1384 (N_1384,N_1018,N_1110);
and U1385 (N_1385,N_1072,N_1061);
or U1386 (N_1386,N_1073,N_1171);
nand U1387 (N_1387,N_1188,N_1128);
or U1388 (N_1388,N_1183,N_1137);
nor U1389 (N_1389,N_1126,N_1054);
nand U1390 (N_1390,N_1094,N_1129);
or U1391 (N_1391,N_1197,N_1124);
and U1392 (N_1392,N_1011,N_1149);
nor U1393 (N_1393,N_1005,N_1149);
or U1394 (N_1394,N_1020,N_1067);
nand U1395 (N_1395,N_1174,N_1047);
nand U1396 (N_1396,N_1174,N_1004);
nor U1397 (N_1397,N_1013,N_1098);
or U1398 (N_1398,N_1000,N_1120);
or U1399 (N_1399,N_1137,N_1153);
nand U1400 (N_1400,N_1384,N_1282);
nand U1401 (N_1401,N_1307,N_1334);
and U1402 (N_1402,N_1323,N_1321);
or U1403 (N_1403,N_1353,N_1260);
xnor U1404 (N_1404,N_1238,N_1341);
nor U1405 (N_1405,N_1311,N_1272);
nand U1406 (N_1406,N_1225,N_1219);
nor U1407 (N_1407,N_1300,N_1333);
nor U1408 (N_1408,N_1223,N_1317);
or U1409 (N_1409,N_1395,N_1327);
or U1410 (N_1410,N_1275,N_1394);
and U1411 (N_1411,N_1257,N_1202);
nand U1412 (N_1412,N_1217,N_1383);
and U1413 (N_1413,N_1367,N_1240);
xnor U1414 (N_1414,N_1355,N_1371);
xnor U1415 (N_1415,N_1251,N_1243);
xor U1416 (N_1416,N_1269,N_1363);
xor U1417 (N_1417,N_1216,N_1369);
and U1418 (N_1418,N_1339,N_1397);
nor U1419 (N_1419,N_1350,N_1229);
nand U1420 (N_1420,N_1263,N_1280);
or U1421 (N_1421,N_1325,N_1372);
nor U1422 (N_1422,N_1283,N_1329);
and U1423 (N_1423,N_1324,N_1304);
and U1424 (N_1424,N_1297,N_1212);
or U1425 (N_1425,N_1389,N_1393);
nor U1426 (N_1426,N_1206,N_1250);
and U1427 (N_1427,N_1235,N_1390);
or U1428 (N_1428,N_1207,N_1375);
xnor U1429 (N_1429,N_1360,N_1222);
xor U1430 (N_1430,N_1302,N_1298);
nor U1431 (N_1431,N_1366,N_1278);
and U1432 (N_1432,N_1342,N_1289);
nand U1433 (N_1433,N_1335,N_1313);
or U1434 (N_1434,N_1247,N_1309);
and U1435 (N_1435,N_1274,N_1331);
and U1436 (N_1436,N_1354,N_1332);
xnor U1437 (N_1437,N_1261,N_1299);
nand U1438 (N_1438,N_1343,N_1242);
nand U1439 (N_1439,N_1239,N_1258);
and U1440 (N_1440,N_1319,N_1204);
or U1441 (N_1441,N_1200,N_1368);
or U1442 (N_1442,N_1221,N_1386);
nor U1443 (N_1443,N_1215,N_1220);
nor U1444 (N_1444,N_1320,N_1357);
xnor U1445 (N_1445,N_1381,N_1241);
and U1446 (N_1446,N_1265,N_1254);
xor U1447 (N_1447,N_1301,N_1330);
nor U1448 (N_1448,N_1249,N_1377);
nor U1449 (N_1449,N_1211,N_1271);
nor U1450 (N_1450,N_1352,N_1213);
and U1451 (N_1451,N_1234,N_1266);
and U1452 (N_1452,N_1227,N_1380);
xnor U1453 (N_1453,N_1267,N_1374);
nor U1454 (N_1454,N_1391,N_1252);
and U1455 (N_1455,N_1348,N_1293);
xnor U1456 (N_1456,N_1399,N_1295);
or U1457 (N_1457,N_1305,N_1376);
nor U1458 (N_1458,N_1387,N_1359);
or U1459 (N_1459,N_1314,N_1286);
and U1460 (N_1460,N_1396,N_1210);
xor U1461 (N_1461,N_1237,N_1315);
nand U1462 (N_1462,N_1326,N_1344);
nor U1463 (N_1463,N_1345,N_1318);
or U1464 (N_1464,N_1306,N_1218);
or U1465 (N_1465,N_1308,N_1310);
or U1466 (N_1466,N_1273,N_1287);
or U1467 (N_1467,N_1361,N_1248);
and U1468 (N_1468,N_1292,N_1370);
nor U1469 (N_1469,N_1373,N_1244);
nor U1470 (N_1470,N_1284,N_1296);
or U1471 (N_1471,N_1268,N_1285);
and U1472 (N_1472,N_1232,N_1208);
nor U1473 (N_1473,N_1236,N_1312);
xnor U1474 (N_1474,N_1346,N_1392);
nand U1475 (N_1475,N_1340,N_1362);
and U1476 (N_1476,N_1337,N_1228);
or U1477 (N_1477,N_1270,N_1253);
and U1478 (N_1478,N_1322,N_1303);
or U1479 (N_1479,N_1291,N_1262);
nor U1480 (N_1480,N_1209,N_1294);
and U1481 (N_1481,N_1214,N_1256);
xor U1482 (N_1482,N_1388,N_1288);
nor U1483 (N_1483,N_1277,N_1385);
and U1484 (N_1484,N_1351,N_1264);
or U1485 (N_1485,N_1364,N_1338);
and U1486 (N_1486,N_1233,N_1246);
and U1487 (N_1487,N_1347,N_1230);
or U1488 (N_1488,N_1382,N_1255);
xnor U1489 (N_1489,N_1281,N_1290);
or U1490 (N_1490,N_1365,N_1379);
and U1491 (N_1491,N_1378,N_1259);
xnor U1492 (N_1492,N_1226,N_1203);
or U1493 (N_1493,N_1336,N_1349);
xnor U1494 (N_1494,N_1276,N_1398);
and U1495 (N_1495,N_1231,N_1358);
xnor U1496 (N_1496,N_1245,N_1201);
or U1497 (N_1497,N_1279,N_1224);
nor U1498 (N_1498,N_1316,N_1328);
and U1499 (N_1499,N_1356,N_1205);
nand U1500 (N_1500,N_1272,N_1364);
nand U1501 (N_1501,N_1223,N_1282);
and U1502 (N_1502,N_1253,N_1223);
and U1503 (N_1503,N_1394,N_1262);
nand U1504 (N_1504,N_1357,N_1248);
nand U1505 (N_1505,N_1205,N_1258);
nand U1506 (N_1506,N_1210,N_1288);
nand U1507 (N_1507,N_1235,N_1377);
xnor U1508 (N_1508,N_1204,N_1285);
or U1509 (N_1509,N_1243,N_1344);
nor U1510 (N_1510,N_1326,N_1346);
nor U1511 (N_1511,N_1228,N_1244);
xor U1512 (N_1512,N_1352,N_1266);
or U1513 (N_1513,N_1223,N_1308);
and U1514 (N_1514,N_1242,N_1304);
xor U1515 (N_1515,N_1258,N_1342);
xor U1516 (N_1516,N_1283,N_1312);
xor U1517 (N_1517,N_1262,N_1391);
nor U1518 (N_1518,N_1288,N_1245);
and U1519 (N_1519,N_1359,N_1372);
and U1520 (N_1520,N_1385,N_1280);
nand U1521 (N_1521,N_1279,N_1275);
xnor U1522 (N_1522,N_1381,N_1340);
and U1523 (N_1523,N_1343,N_1237);
and U1524 (N_1524,N_1363,N_1367);
and U1525 (N_1525,N_1383,N_1298);
xnor U1526 (N_1526,N_1383,N_1368);
nand U1527 (N_1527,N_1279,N_1329);
xor U1528 (N_1528,N_1304,N_1338);
nor U1529 (N_1529,N_1373,N_1255);
or U1530 (N_1530,N_1222,N_1285);
nor U1531 (N_1531,N_1282,N_1247);
and U1532 (N_1532,N_1280,N_1255);
or U1533 (N_1533,N_1398,N_1221);
nor U1534 (N_1534,N_1256,N_1218);
nor U1535 (N_1535,N_1214,N_1217);
and U1536 (N_1536,N_1380,N_1217);
and U1537 (N_1537,N_1271,N_1269);
xor U1538 (N_1538,N_1328,N_1200);
nor U1539 (N_1539,N_1342,N_1389);
nor U1540 (N_1540,N_1366,N_1378);
xnor U1541 (N_1541,N_1270,N_1233);
nor U1542 (N_1542,N_1351,N_1377);
nor U1543 (N_1543,N_1280,N_1384);
and U1544 (N_1544,N_1397,N_1265);
xnor U1545 (N_1545,N_1286,N_1397);
nand U1546 (N_1546,N_1379,N_1280);
xor U1547 (N_1547,N_1278,N_1399);
xnor U1548 (N_1548,N_1378,N_1399);
nor U1549 (N_1549,N_1339,N_1343);
xnor U1550 (N_1550,N_1267,N_1395);
nand U1551 (N_1551,N_1321,N_1235);
or U1552 (N_1552,N_1250,N_1384);
and U1553 (N_1553,N_1242,N_1262);
xnor U1554 (N_1554,N_1270,N_1282);
and U1555 (N_1555,N_1377,N_1279);
and U1556 (N_1556,N_1289,N_1322);
xnor U1557 (N_1557,N_1244,N_1379);
or U1558 (N_1558,N_1275,N_1340);
nand U1559 (N_1559,N_1226,N_1363);
nand U1560 (N_1560,N_1337,N_1331);
nand U1561 (N_1561,N_1250,N_1303);
and U1562 (N_1562,N_1234,N_1220);
nand U1563 (N_1563,N_1378,N_1298);
xor U1564 (N_1564,N_1329,N_1394);
xor U1565 (N_1565,N_1292,N_1324);
xor U1566 (N_1566,N_1269,N_1281);
nor U1567 (N_1567,N_1338,N_1346);
and U1568 (N_1568,N_1260,N_1332);
xnor U1569 (N_1569,N_1306,N_1243);
nor U1570 (N_1570,N_1285,N_1332);
and U1571 (N_1571,N_1395,N_1386);
nand U1572 (N_1572,N_1372,N_1222);
and U1573 (N_1573,N_1234,N_1321);
or U1574 (N_1574,N_1234,N_1325);
nand U1575 (N_1575,N_1200,N_1309);
nor U1576 (N_1576,N_1278,N_1223);
nor U1577 (N_1577,N_1294,N_1216);
xnor U1578 (N_1578,N_1206,N_1321);
and U1579 (N_1579,N_1276,N_1271);
nand U1580 (N_1580,N_1200,N_1224);
or U1581 (N_1581,N_1256,N_1296);
nor U1582 (N_1582,N_1251,N_1204);
nand U1583 (N_1583,N_1365,N_1225);
nor U1584 (N_1584,N_1356,N_1312);
nand U1585 (N_1585,N_1376,N_1257);
nand U1586 (N_1586,N_1385,N_1292);
nand U1587 (N_1587,N_1343,N_1370);
xor U1588 (N_1588,N_1286,N_1384);
nor U1589 (N_1589,N_1365,N_1201);
nand U1590 (N_1590,N_1230,N_1226);
and U1591 (N_1591,N_1305,N_1343);
nand U1592 (N_1592,N_1351,N_1237);
xnor U1593 (N_1593,N_1294,N_1239);
xor U1594 (N_1594,N_1296,N_1377);
nand U1595 (N_1595,N_1264,N_1300);
xor U1596 (N_1596,N_1271,N_1278);
xor U1597 (N_1597,N_1258,N_1265);
nor U1598 (N_1598,N_1236,N_1235);
nand U1599 (N_1599,N_1335,N_1338);
or U1600 (N_1600,N_1506,N_1477);
nor U1601 (N_1601,N_1475,N_1539);
or U1602 (N_1602,N_1521,N_1546);
xnor U1603 (N_1603,N_1599,N_1571);
and U1604 (N_1604,N_1588,N_1509);
and U1605 (N_1605,N_1552,N_1493);
and U1606 (N_1606,N_1446,N_1514);
nand U1607 (N_1607,N_1432,N_1435);
xnor U1608 (N_1608,N_1484,N_1444);
and U1609 (N_1609,N_1587,N_1492);
or U1610 (N_1610,N_1421,N_1408);
or U1611 (N_1611,N_1445,N_1401);
nor U1612 (N_1612,N_1553,N_1410);
xnor U1613 (N_1613,N_1453,N_1544);
and U1614 (N_1614,N_1465,N_1447);
nand U1615 (N_1615,N_1481,N_1425);
nor U1616 (N_1616,N_1450,N_1551);
nor U1617 (N_1617,N_1449,N_1576);
xor U1618 (N_1618,N_1478,N_1543);
and U1619 (N_1619,N_1508,N_1547);
or U1620 (N_1620,N_1441,N_1594);
nand U1621 (N_1621,N_1554,N_1569);
nand U1622 (N_1622,N_1457,N_1461);
nor U1623 (N_1623,N_1503,N_1486);
nor U1624 (N_1624,N_1448,N_1412);
and U1625 (N_1625,N_1479,N_1504);
or U1626 (N_1626,N_1534,N_1472);
or U1627 (N_1627,N_1519,N_1419);
or U1628 (N_1628,N_1585,N_1545);
and U1629 (N_1629,N_1532,N_1557);
nand U1630 (N_1630,N_1436,N_1443);
nand U1631 (N_1631,N_1595,N_1578);
nor U1632 (N_1632,N_1499,N_1424);
xnor U1633 (N_1633,N_1411,N_1483);
nor U1634 (N_1634,N_1582,N_1538);
nand U1635 (N_1635,N_1525,N_1455);
nand U1636 (N_1636,N_1462,N_1517);
nor U1637 (N_1637,N_1418,N_1511);
nand U1638 (N_1638,N_1597,N_1530);
nor U1639 (N_1639,N_1400,N_1556);
xor U1640 (N_1640,N_1581,N_1434);
xnor U1641 (N_1641,N_1515,N_1526);
nand U1642 (N_1642,N_1560,N_1502);
or U1643 (N_1643,N_1463,N_1540);
or U1644 (N_1644,N_1409,N_1561);
and U1645 (N_1645,N_1482,N_1429);
xnor U1646 (N_1646,N_1531,N_1476);
xor U1647 (N_1647,N_1574,N_1579);
and U1648 (N_1648,N_1431,N_1420);
nor U1649 (N_1649,N_1416,N_1501);
nor U1650 (N_1650,N_1572,N_1510);
nand U1651 (N_1651,N_1584,N_1489);
or U1652 (N_1652,N_1403,N_1598);
xor U1653 (N_1653,N_1537,N_1495);
or U1654 (N_1654,N_1589,N_1550);
nor U1655 (N_1655,N_1490,N_1518);
nand U1656 (N_1656,N_1573,N_1415);
nand U1657 (N_1657,N_1440,N_1406);
xnor U1658 (N_1658,N_1563,N_1485);
or U1659 (N_1659,N_1414,N_1488);
nor U1660 (N_1660,N_1467,N_1580);
nand U1661 (N_1661,N_1459,N_1535);
or U1662 (N_1662,N_1596,N_1512);
xor U1663 (N_1663,N_1466,N_1524);
nand U1664 (N_1664,N_1570,N_1555);
nor U1665 (N_1665,N_1520,N_1558);
and U1666 (N_1666,N_1470,N_1536);
or U1667 (N_1667,N_1464,N_1591);
nor U1668 (N_1668,N_1564,N_1496);
xor U1669 (N_1669,N_1577,N_1437);
xor U1670 (N_1670,N_1423,N_1541);
or U1671 (N_1671,N_1422,N_1427);
nor U1672 (N_1672,N_1473,N_1505);
and U1673 (N_1673,N_1507,N_1417);
and U1674 (N_1674,N_1491,N_1549);
xnor U1675 (N_1675,N_1566,N_1494);
xor U1676 (N_1676,N_1480,N_1442);
xnor U1677 (N_1677,N_1528,N_1405);
nor U1678 (N_1678,N_1527,N_1533);
and U1679 (N_1679,N_1500,N_1438);
nand U1680 (N_1680,N_1548,N_1542);
nand U1681 (N_1681,N_1562,N_1586);
nor U1682 (N_1682,N_1458,N_1513);
and U1683 (N_1683,N_1565,N_1487);
nor U1684 (N_1684,N_1568,N_1590);
or U1685 (N_1685,N_1454,N_1407);
nand U1686 (N_1686,N_1469,N_1404);
nor U1687 (N_1687,N_1592,N_1460);
nand U1688 (N_1688,N_1474,N_1402);
nand U1689 (N_1689,N_1516,N_1413);
nand U1690 (N_1690,N_1529,N_1497);
nor U1691 (N_1691,N_1583,N_1428);
nor U1692 (N_1692,N_1468,N_1456);
and U1693 (N_1693,N_1567,N_1523);
or U1694 (N_1694,N_1426,N_1593);
xnor U1695 (N_1695,N_1522,N_1451);
and U1696 (N_1696,N_1430,N_1498);
or U1697 (N_1697,N_1433,N_1452);
nor U1698 (N_1698,N_1559,N_1471);
nor U1699 (N_1699,N_1439,N_1575);
and U1700 (N_1700,N_1589,N_1553);
xnor U1701 (N_1701,N_1555,N_1598);
nor U1702 (N_1702,N_1558,N_1415);
nand U1703 (N_1703,N_1448,N_1497);
or U1704 (N_1704,N_1420,N_1553);
and U1705 (N_1705,N_1422,N_1465);
nor U1706 (N_1706,N_1465,N_1585);
and U1707 (N_1707,N_1431,N_1537);
or U1708 (N_1708,N_1543,N_1436);
xnor U1709 (N_1709,N_1502,N_1451);
nand U1710 (N_1710,N_1476,N_1438);
or U1711 (N_1711,N_1552,N_1571);
nand U1712 (N_1712,N_1488,N_1536);
or U1713 (N_1713,N_1558,N_1575);
nand U1714 (N_1714,N_1525,N_1554);
xnor U1715 (N_1715,N_1508,N_1515);
nand U1716 (N_1716,N_1588,N_1482);
or U1717 (N_1717,N_1542,N_1581);
and U1718 (N_1718,N_1412,N_1517);
nand U1719 (N_1719,N_1472,N_1565);
nand U1720 (N_1720,N_1478,N_1561);
or U1721 (N_1721,N_1542,N_1575);
and U1722 (N_1722,N_1551,N_1420);
and U1723 (N_1723,N_1483,N_1434);
and U1724 (N_1724,N_1512,N_1543);
nand U1725 (N_1725,N_1560,N_1407);
xnor U1726 (N_1726,N_1556,N_1520);
xnor U1727 (N_1727,N_1473,N_1532);
nand U1728 (N_1728,N_1567,N_1483);
and U1729 (N_1729,N_1430,N_1444);
xnor U1730 (N_1730,N_1501,N_1584);
nor U1731 (N_1731,N_1551,N_1525);
nand U1732 (N_1732,N_1430,N_1586);
nand U1733 (N_1733,N_1474,N_1450);
xnor U1734 (N_1734,N_1510,N_1436);
xnor U1735 (N_1735,N_1461,N_1467);
and U1736 (N_1736,N_1416,N_1443);
nand U1737 (N_1737,N_1468,N_1449);
nor U1738 (N_1738,N_1469,N_1527);
nand U1739 (N_1739,N_1597,N_1523);
and U1740 (N_1740,N_1598,N_1484);
and U1741 (N_1741,N_1510,N_1494);
nor U1742 (N_1742,N_1453,N_1475);
nand U1743 (N_1743,N_1415,N_1492);
or U1744 (N_1744,N_1515,N_1524);
and U1745 (N_1745,N_1439,N_1505);
xor U1746 (N_1746,N_1595,N_1495);
xor U1747 (N_1747,N_1531,N_1402);
or U1748 (N_1748,N_1484,N_1517);
xor U1749 (N_1749,N_1562,N_1577);
xor U1750 (N_1750,N_1466,N_1534);
nand U1751 (N_1751,N_1505,N_1477);
and U1752 (N_1752,N_1517,N_1549);
xnor U1753 (N_1753,N_1471,N_1442);
nand U1754 (N_1754,N_1441,N_1583);
nand U1755 (N_1755,N_1442,N_1581);
nor U1756 (N_1756,N_1469,N_1598);
and U1757 (N_1757,N_1573,N_1421);
xor U1758 (N_1758,N_1407,N_1527);
xnor U1759 (N_1759,N_1469,N_1446);
nor U1760 (N_1760,N_1467,N_1562);
nor U1761 (N_1761,N_1432,N_1568);
xnor U1762 (N_1762,N_1461,N_1584);
nor U1763 (N_1763,N_1445,N_1553);
nor U1764 (N_1764,N_1587,N_1482);
xor U1765 (N_1765,N_1478,N_1520);
and U1766 (N_1766,N_1433,N_1415);
and U1767 (N_1767,N_1469,N_1433);
xor U1768 (N_1768,N_1457,N_1563);
and U1769 (N_1769,N_1508,N_1564);
xor U1770 (N_1770,N_1529,N_1522);
nor U1771 (N_1771,N_1469,N_1588);
xor U1772 (N_1772,N_1455,N_1415);
or U1773 (N_1773,N_1425,N_1552);
nor U1774 (N_1774,N_1414,N_1535);
nand U1775 (N_1775,N_1424,N_1481);
and U1776 (N_1776,N_1542,N_1459);
nor U1777 (N_1777,N_1440,N_1421);
nor U1778 (N_1778,N_1543,N_1519);
nor U1779 (N_1779,N_1447,N_1466);
nor U1780 (N_1780,N_1551,N_1463);
or U1781 (N_1781,N_1498,N_1536);
or U1782 (N_1782,N_1528,N_1487);
and U1783 (N_1783,N_1414,N_1410);
nor U1784 (N_1784,N_1538,N_1489);
nand U1785 (N_1785,N_1500,N_1497);
nor U1786 (N_1786,N_1527,N_1453);
or U1787 (N_1787,N_1450,N_1552);
nor U1788 (N_1788,N_1468,N_1508);
nand U1789 (N_1789,N_1461,N_1568);
or U1790 (N_1790,N_1417,N_1578);
xor U1791 (N_1791,N_1594,N_1537);
and U1792 (N_1792,N_1406,N_1400);
nand U1793 (N_1793,N_1512,N_1514);
or U1794 (N_1794,N_1539,N_1409);
nor U1795 (N_1795,N_1557,N_1446);
nand U1796 (N_1796,N_1476,N_1534);
or U1797 (N_1797,N_1412,N_1519);
nor U1798 (N_1798,N_1401,N_1422);
and U1799 (N_1799,N_1543,N_1528);
and U1800 (N_1800,N_1757,N_1755);
xor U1801 (N_1801,N_1669,N_1740);
and U1802 (N_1802,N_1727,N_1691);
nand U1803 (N_1803,N_1614,N_1647);
nand U1804 (N_1804,N_1653,N_1774);
xnor U1805 (N_1805,N_1686,N_1670);
or U1806 (N_1806,N_1722,N_1778);
xor U1807 (N_1807,N_1660,N_1769);
and U1808 (N_1808,N_1667,N_1662);
and U1809 (N_1809,N_1765,N_1745);
or U1810 (N_1810,N_1616,N_1751);
nor U1811 (N_1811,N_1652,N_1752);
nor U1812 (N_1812,N_1623,N_1654);
xor U1813 (N_1813,N_1761,N_1775);
xor U1814 (N_1814,N_1735,N_1634);
and U1815 (N_1815,N_1682,N_1607);
nor U1816 (N_1816,N_1631,N_1787);
nand U1817 (N_1817,N_1690,N_1693);
nand U1818 (N_1818,N_1718,N_1620);
xnor U1819 (N_1819,N_1611,N_1696);
and U1820 (N_1820,N_1663,N_1697);
nor U1821 (N_1821,N_1723,N_1759);
nand U1822 (N_1822,N_1649,N_1706);
nor U1823 (N_1823,N_1675,N_1680);
and U1824 (N_1824,N_1726,N_1685);
nor U1825 (N_1825,N_1703,N_1767);
nand U1826 (N_1826,N_1734,N_1701);
and U1827 (N_1827,N_1629,N_1694);
and U1828 (N_1828,N_1641,N_1770);
and U1829 (N_1829,N_1721,N_1799);
xor U1830 (N_1830,N_1618,N_1738);
xnor U1831 (N_1831,N_1783,N_1688);
nor U1832 (N_1832,N_1664,N_1737);
nand U1833 (N_1833,N_1602,N_1600);
and U1834 (N_1834,N_1677,N_1733);
or U1835 (N_1835,N_1635,N_1729);
nand U1836 (N_1836,N_1781,N_1754);
or U1837 (N_1837,N_1674,N_1771);
and U1838 (N_1838,N_1773,N_1743);
or U1839 (N_1839,N_1665,N_1731);
or U1840 (N_1840,N_1613,N_1687);
and U1841 (N_1841,N_1646,N_1604);
or U1842 (N_1842,N_1699,N_1668);
nand U1843 (N_1843,N_1749,N_1717);
or U1844 (N_1844,N_1782,N_1744);
nor U1845 (N_1845,N_1777,N_1753);
nand U1846 (N_1846,N_1764,N_1644);
nand U1847 (N_1847,N_1621,N_1789);
xnor U1848 (N_1848,N_1746,N_1725);
xor U1849 (N_1849,N_1756,N_1747);
or U1850 (N_1850,N_1609,N_1750);
nor U1851 (N_1851,N_1619,N_1730);
nand U1852 (N_1852,N_1772,N_1617);
xnor U1853 (N_1853,N_1788,N_1640);
nand U1854 (N_1854,N_1684,N_1624);
nand U1855 (N_1855,N_1741,N_1622);
nand U1856 (N_1856,N_1625,N_1656);
nand U1857 (N_1857,N_1608,N_1601);
and U1858 (N_1858,N_1758,N_1628);
and U1859 (N_1859,N_1681,N_1612);
xor U1860 (N_1860,N_1714,N_1712);
and U1861 (N_1861,N_1719,N_1638);
and U1862 (N_1862,N_1672,N_1704);
nand U1863 (N_1863,N_1710,N_1679);
nor U1864 (N_1864,N_1762,N_1659);
or U1865 (N_1865,N_1661,N_1713);
nand U1866 (N_1866,N_1708,N_1707);
or U1867 (N_1867,N_1716,N_1797);
xor U1868 (N_1868,N_1658,N_1705);
nand U1869 (N_1869,N_1790,N_1698);
nand U1870 (N_1870,N_1676,N_1742);
or U1871 (N_1871,N_1732,N_1780);
or U1872 (N_1872,N_1655,N_1695);
xnor U1873 (N_1873,N_1794,N_1666);
nor U1874 (N_1874,N_1648,N_1724);
nand U1875 (N_1875,N_1673,N_1798);
nand U1876 (N_1876,N_1728,N_1615);
and U1877 (N_1877,N_1636,N_1791);
nor U1878 (N_1878,N_1796,N_1650);
xor U1879 (N_1879,N_1639,N_1671);
xor U1880 (N_1880,N_1683,N_1610);
nor U1881 (N_1881,N_1763,N_1702);
or U1882 (N_1882,N_1627,N_1603);
and U1883 (N_1883,N_1720,N_1709);
nor U1884 (N_1884,N_1768,N_1633);
nand U1885 (N_1885,N_1748,N_1776);
or U1886 (N_1886,N_1766,N_1626);
xor U1887 (N_1887,N_1651,N_1711);
and U1888 (N_1888,N_1784,N_1605);
nor U1889 (N_1889,N_1795,N_1657);
or U1890 (N_1890,N_1779,N_1645);
and U1891 (N_1891,N_1606,N_1642);
nand U1892 (N_1892,N_1700,N_1692);
and U1893 (N_1893,N_1793,N_1792);
and U1894 (N_1894,N_1630,N_1715);
or U1895 (N_1895,N_1785,N_1643);
nor U1896 (N_1896,N_1678,N_1786);
nand U1897 (N_1897,N_1760,N_1632);
and U1898 (N_1898,N_1637,N_1736);
or U1899 (N_1899,N_1689,N_1739);
nor U1900 (N_1900,N_1749,N_1795);
xnor U1901 (N_1901,N_1695,N_1704);
xnor U1902 (N_1902,N_1652,N_1645);
nor U1903 (N_1903,N_1654,N_1670);
and U1904 (N_1904,N_1624,N_1651);
nand U1905 (N_1905,N_1796,N_1608);
or U1906 (N_1906,N_1793,N_1720);
xnor U1907 (N_1907,N_1690,N_1680);
and U1908 (N_1908,N_1743,N_1658);
or U1909 (N_1909,N_1737,N_1709);
nand U1910 (N_1910,N_1751,N_1772);
or U1911 (N_1911,N_1754,N_1699);
nor U1912 (N_1912,N_1646,N_1747);
nor U1913 (N_1913,N_1750,N_1783);
and U1914 (N_1914,N_1677,N_1747);
or U1915 (N_1915,N_1647,N_1612);
and U1916 (N_1916,N_1697,N_1624);
nor U1917 (N_1917,N_1779,N_1634);
and U1918 (N_1918,N_1776,N_1727);
nor U1919 (N_1919,N_1626,N_1791);
nor U1920 (N_1920,N_1660,N_1742);
nor U1921 (N_1921,N_1639,N_1637);
nor U1922 (N_1922,N_1698,N_1711);
and U1923 (N_1923,N_1750,N_1709);
or U1924 (N_1924,N_1635,N_1791);
xor U1925 (N_1925,N_1685,N_1763);
nand U1926 (N_1926,N_1667,N_1619);
and U1927 (N_1927,N_1604,N_1783);
or U1928 (N_1928,N_1672,N_1624);
nor U1929 (N_1929,N_1713,N_1784);
and U1930 (N_1930,N_1784,N_1743);
nor U1931 (N_1931,N_1603,N_1716);
nor U1932 (N_1932,N_1600,N_1773);
and U1933 (N_1933,N_1616,N_1727);
and U1934 (N_1934,N_1615,N_1651);
xnor U1935 (N_1935,N_1664,N_1780);
xor U1936 (N_1936,N_1635,N_1723);
and U1937 (N_1937,N_1776,N_1616);
nand U1938 (N_1938,N_1685,N_1784);
and U1939 (N_1939,N_1751,N_1618);
nand U1940 (N_1940,N_1693,N_1639);
and U1941 (N_1941,N_1732,N_1618);
nor U1942 (N_1942,N_1775,N_1691);
or U1943 (N_1943,N_1633,N_1662);
and U1944 (N_1944,N_1676,N_1776);
xor U1945 (N_1945,N_1704,N_1715);
nor U1946 (N_1946,N_1762,N_1627);
nor U1947 (N_1947,N_1672,N_1649);
nor U1948 (N_1948,N_1773,N_1689);
and U1949 (N_1949,N_1796,N_1730);
or U1950 (N_1950,N_1770,N_1731);
nand U1951 (N_1951,N_1668,N_1753);
xnor U1952 (N_1952,N_1661,N_1620);
xor U1953 (N_1953,N_1633,N_1601);
or U1954 (N_1954,N_1728,N_1679);
xor U1955 (N_1955,N_1772,N_1603);
and U1956 (N_1956,N_1601,N_1673);
nand U1957 (N_1957,N_1701,N_1728);
nor U1958 (N_1958,N_1726,N_1774);
nor U1959 (N_1959,N_1798,N_1601);
and U1960 (N_1960,N_1780,N_1735);
and U1961 (N_1961,N_1759,N_1725);
xor U1962 (N_1962,N_1627,N_1722);
xnor U1963 (N_1963,N_1713,N_1625);
nand U1964 (N_1964,N_1776,N_1695);
or U1965 (N_1965,N_1620,N_1649);
xnor U1966 (N_1966,N_1758,N_1705);
and U1967 (N_1967,N_1750,N_1672);
or U1968 (N_1968,N_1627,N_1780);
xnor U1969 (N_1969,N_1783,N_1744);
or U1970 (N_1970,N_1789,N_1795);
xnor U1971 (N_1971,N_1652,N_1697);
xnor U1972 (N_1972,N_1615,N_1660);
xor U1973 (N_1973,N_1780,N_1713);
nor U1974 (N_1974,N_1614,N_1657);
xnor U1975 (N_1975,N_1637,N_1692);
xnor U1976 (N_1976,N_1611,N_1752);
nor U1977 (N_1977,N_1607,N_1787);
nor U1978 (N_1978,N_1650,N_1671);
or U1979 (N_1979,N_1780,N_1604);
and U1980 (N_1980,N_1635,N_1680);
or U1981 (N_1981,N_1711,N_1683);
xnor U1982 (N_1982,N_1787,N_1740);
and U1983 (N_1983,N_1755,N_1647);
and U1984 (N_1984,N_1751,N_1661);
nor U1985 (N_1985,N_1716,N_1671);
nand U1986 (N_1986,N_1747,N_1796);
and U1987 (N_1987,N_1604,N_1637);
nor U1988 (N_1988,N_1749,N_1734);
nor U1989 (N_1989,N_1788,N_1751);
xor U1990 (N_1990,N_1773,N_1749);
nand U1991 (N_1991,N_1766,N_1614);
xor U1992 (N_1992,N_1616,N_1724);
nor U1993 (N_1993,N_1647,N_1611);
nor U1994 (N_1994,N_1734,N_1716);
and U1995 (N_1995,N_1708,N_1763);
xor U1996 (N_1996,N_1653,N_1728);
xnor U1997 (N_1997,N_1738,N_1602);
or U1998 (N_1998,N_1706,N_1670);
and U1999 (N_1999,N_1616,N_1643);
nor U2000 (N_2000,N_1978,N_1995);
and U2001 (N_2001,N_1858,N_1933);
xor U2002 (N_2002,N_1885,N_1901);
xor U2003 (N_2003,N_1824,N_1984);
and U2004 (N_2004,N_1891,N_1906);
nor U2005 (N_2005,N_1972,N_1918);
nor U2006 (N_2006,N_1864,N_1845);
nor U2007 (N_2007,N_1992,N_1828);
nand U2008 (N_2008,N_1979,N_1955);
xnor U2009 (N_2009,N_1849,N_1996);
nor U2010 (N_2010,N_1903,N_1813);
xor U2011 (N_2011,N_1865,N_1920);
nand U2012 (N_2012,N_1949,N_1836);
xnor U2013 (N_2013,N_1910,N_1905);
xnor U2014 (N_2014,N_1951,N_1954);
nor U2015 (N_2015,N_1914,N_1957);
and U2016 (N_2016,N_1988,N_1942);
xor U2017 (N_2017,N_1803,N_1938);
nor U2018 (N_2018,N_1946,N_1961);
xor U2019 (N_2019,N_1923,N_1851);
xnor U2020 (N_2020,N_1846,N_1971);
nand U2021 (N_2021,N_1983,N_1882);
xor U2022 (N_2022,N_1814,N_1963);
and U2023 (N_2023,N_1965,N_1843);
nand U2024 (N_2024,N_1835,N_1893);
and U2025 (N_2025,N_1908,N_1883);
and U2026 (N_2026,N_1856,N_1876);
or U2027 (N_2027,N_1810,N_1944);
xor U2028 (N_2028,N_1964,N_1833);
or U2029 (N_2029,N_1907,N_1982);
nor U2030 (N_2030,N_1820,N_1927);
and U2031 (N_2031,N_1838,N_1928);
xnor U2032 (N_2032,N_1808,N_1807);
xor U2033 (N_2033,N_1952,N_1853);
nor U2034 (N_2034,N_1913,N_1941);
nor U2035 (N_2035,N_1977,N_1800);
nor U2036 (N_2036,N_1950,N_1841);
nand U2037 (N_2037,N_1980,N_1956);
and U2038 (N_2038,N_1986,N_1967);
xor U2039 (N_2039,N_1870,N_1902);
xnor U2040 (N_2040,N_1840,N_1939);
nor U2041 (N_2041,N_1868,N_1811);
nand U2042 (N_2042,N_1998,N_1869);
nor U2043 (N_2043,N_1993,N_1875);
and U2044 (N_2044,N_1873,N_1847);
nand U2045 (N_2045,N_1815,N_1917);
and U2046 (N_2046,N_1943,N_1900);
nand U2047 (N_2047,N_1929,N_1960);
nand U2048 (N_2048,N_1812,N_1806);
nand U2049 (N_2049,N_1975,N_1855);
nand U2050 (N_2050,N_1987,N_1999);
and U2051 (N_2051,N_1931,N_1860);
xnor U2052 (N_2052,N_1966,N_1817);
and U2053 (N_2053,N_1916,N_1818);
or U2054 (N_2054,N_1832,N_1854);
nand U2055 (N_2055,N_1889,N_1867);
nor U2056 (N_2056,N_1879,N_1962);
or U2057 (N_2057,N_1924,N_1970);
nor U2058 (N_2058,N_1884,N_1877);
nor U2059 (N_2059,N_1852,N_1802);
or U2060 (N_2060,N_1909,N_1888);
nor U2061 (N_2061,N_1816,N_1895);
xor U2062 (N_2062,N_1899,N_1878);
xnor U2063 (N_2063,N_1890,N_1904);
nor U2064 (N_2064,N_1990,N_1837);
nor U2065 (N_2065,N_1842,N_1898);
nor U2066 (N_2066,N_1892,N_1911);
and U2067 (N_2067,N_1821,N_1915);
nand U2068 (N_2068,N_1947,N_1830);
or U2069 (N_2069,N_1872,N_1871);
and U2070 (N_2070,N_1973,N_1861);
nor U2071 (N_2071,N_1894,N_1948);
nor U2072 (N_2072,N_1922,N_1974);
nor U2073 (N_2073,N_1886,N_1862);
nand U2074 (N_2074,N_1989,N_1953);
nor U2075 (N_2075,N_1859,N_1823);
and U2076 (N_2076,N_1926,N_1805);
xnor U2077 (N_2077,N_1991,N_1925);
nand U2078 (N_2078,N_1994,N_1809);
and U2079 (N_2079,N_1827,N_1976);
xnor U2080 (N_2080,N_1968,N_1940);
and U2081 (N_2081,N_1959,N_1935);
nand U2082 (N_2082,N_1826,N_1822);
xnor U2083 (N_2083,N_1848,N_1985);
xnor U2084 (N_2084,N_1874,N_1881);
nand U2085 (N_2085,N_1936,N_1887);
nand U2086 (N_2086,N_1932,N_1921);
and U2087 (N_2087,N_1912,N_1804);
xnor U2088 (N_2088,N_1819,N_1934);
nand U2089 (N_2089,N_1829,N_1801);
and U2090 (N_2090,N_1834,N_1880);
nor U2091 (N_2091,N_1844,N_1850);
nor U2092 (N_2092,N_1937,N_1857);
and U2093 (N_2093,N_1825,N_1866);
nor U2094 (N_2094,N_1831,N_1945);
nand U2095 (N_2095,N_1839,N_1930);
nor U2096 (N_2096,N_1981,N_1919);
nand U2097 (N_2097,N_1863,N_1896);
or U2098 (N_2098,N_1897,N_1997);
or U2099 (N_2099,N_1969,N_1958);
nand U2100 (N_2100,N_1934,N_1851);
xnor U2101 (N_2101,N_1824,N_1957);
nand U2102 (N_2102,N_1849,N_1932);
or U2103 (N_2103,N_1839,N_1973);
nand U2104 (N_2104,N_1948,N_1915);
nand U2105 (N_2105,N_1920,N_1932);
and U2106 (N_2106,N_1922,N_1837);
or U2107 (N_2107,N_1904,N_1884);
nand U2108 (N_2108,N_1889,N_1857);
and U2109 (N_2109,N_1804,N_1969);
and U2110 (N_2110,N_1961,N_1803);
and U2111 (N_2111,N_1908,N_1888);
nor U2112 (N_2112,N_1876,N_1901);
or U2113 (N_2113,N_1893,N_1842);
nor U2114 (N_2114,N_1883,N_1881);
nand U2115 (N_2115,N_1925,N_1880);
and U2116 (N_2116,N_1967,N_1811);
nand U2117 (N_2117,N_1874,N_1861);
or U2118 (N_2118,N_1882,N_1843);
nand U2119 (N_2119,N_1954,N_1817);
or U2120 (N_2120,N_1814,N_1846);
nor U2121 (N_2121,N_1909,N_1998);
nand U2122 (N_2122,N_1992,N_1905);
nand U2123 (N_2123,N_1852,N_1985);
nand U2124 (N_2124,N_1825,N_1912);
nor U2125 (N_2125,N_1874,N_1862);
or U2126 (N_2126,N_1854,N_1872);
nand U2127 (N_2127,N_1954,N_1975);
or U2128 (N_2128,N_1866,N_1803);
xor U2129 (N_2129,N_1803,N_1872);
or U2130 (N_2130,N_1969,N_1839);
or U2131 (N_2131,N_1806,N_1915);
and U2132 (N_2132,N_1983,N_1843);
nand U2133 (N_2133,N_1960,N_1839);
or U2134 (N_2134,N_1948,N_1855);
nand U2135 (N_2135,N_1947,N_1823);
xnor U2136 (N_2136,N_1818,N_1842);
or U2137 (N_2137,N_1915,N_1989);
and U2138 (N_2138,N_1804,N_1920);
xor U2139 (N_2139,N_1921,N_1918);
xnor U2140 (N_2140,N_1860,N_1856);
and U2141 (N_2141,N_1999,N_1836);
nand U2142 (N_2142,N_1867,N_1973);
xnor U2143 (N_2143,N_1952,N_1984);
or U2144 (N_2144,N_1833,N_1916);
and U2145 (N_2145,N_1831,N_1916);
nor U2146 (N_2146,N_1808,N_1885);
or U2147 (N_2147,N_1824,N_1910);
nor U2148 (N_2148,N_1883,N_1904);
xnor U2149 (N_2149,N_1810,N_1904);
and U2150 (N_2150,N_1816,N_1949);
nor U2151 (N_2151,N_1873,N_1935);
nor U2152 (N_2152,N_1860,N_1936);
nor U2153 (N_2153,N_1837,N_1834);
nor U2154 (N_2154,N_1810,N_1900);
nor U2155 (N_2155,N_1834,N_1997);
nor U2156 (N_2156,N_1904,N_1827);
or U2157 (N_2157,N_1907,N_1831);
nor U2158 (N_2158,N_1835,N_1868);
nand U2159 (N_2159,N_1806,N_1978);
xnor U2160 (N_2160,N_1938,N_1888);
or U2161 (N_2161,N_1981,N_1803);
or U2162 (N_2162,N_1899,N_1806);
nor U2163 (N_2163,N_1814,N_1817);
nand U2164 (N_2164,N_1942,N_1952);
xor U2165 (N_2165,N_1839,N_1812);
nor U2166 (N_2166,N_1869,N_1909);
xor U2167 (N_2167,N_1916,N_1954);
nor U2168 (N_2168,N_1894,N_1927);
xnor U2169 (N_2169,N_1861,N_1883);
and U2170 (N_2170,N_1977,N_1816);
nor U2171 (N_2171,N_1987,N_1977);
nor U2172 (N_2172,N_1833,N_1842);
xnor U2173 (N_2173,N_1952,N_1966);
nand U2174 (N_2174,N_1875,N_1868);
nand U2175 (N_2175,N_1820,N_1955);
nand U2176 (N_2176,N_1880,N_1809);
or U2177 (N_2177,N_1848,N_1948);
or U2178 (N_2178,N_1832,N_1863);
and U2179 (N_2179,N_1840,N_1915);
and U2180 (N_2180,N_1966,N_1807);
and U2181 (N_2181,N_1954,N_1907);
xor U2182 (N_2182,N_1868,N_1834);
nor U2183 (N_2183,N_1932,N_1927);
nor U2184 (N_2184,N_1964,N_1992);
nand U2185 (N_2185,N_1904,N_1941);
nand U2186 (N_2186,N_1969,N_1899);
nor U2187 (N_2187,N_1885,N_1991);
and U2188 (N_2188,N_1982,N_1828);
and U2189 (N_2189,N_1917,N_1938);
nor U2190 (N_2190,N_1810,N_1913);
or U2191 (N_2191,N_1824,N_1817);
nor U2192 (N_2192,N_1984,N_1835);
and U2193 (N_2193,N_1985,N_1989);
xnor U2194 (N_2194,N_1827,N_1862);
nand U2195 (N_2195,N_1927,N_1851);
and U2196 (N_2196,N_1836,N_1804);
xnor U2197 (N_2197,N_1961,N_1823);
and U2198 (N_2198,N_1853,N_1811);
and U2199 (N_2199,N_1822,N_1896);
xnor U2200 (N_2200,N_2042,N_2043);
xnor U2201 (N_2201,N_2030,N_2147);
or U2202 (N_2202,N_2164,N_2077);
nand U2203 (N_2203,N_2000,N_2114);
nor U2204 (N_2204,N_2125,N_2158);
or U2205 (N_2205,N_2102,N_2083);
and U2206 (N_2206,N_2155,N_2135);
xor U2207 (N_2207,N_2103,N_2034);
and U2208 (N_2208,N_2037,N_2196);
xnor U2209 (N_2209,N_2015,N_2018);
or U2210 (N_2210,N_2048,N_2004);
and U2211 (N_2211,N_2076,N_2002);
and U2212 (N_2212,N_2169,N_2095);
nand U2213 (N_2213,N_2016,N_2163);
nor U2214 (N_2214,N_2003,N_2139);
nand U2215 (N_2215,N_2086,N_2069);
and U2216 (N_2216,N_2184,N_2143);
nand U2217 (N_2217,N_2148,N_2113);
and U2218 (N_2218,N_2185,N_2180);
nand U2219 (N_2219,N_2096,N_2072);
or U2220 (N_2220,N_2058,N_2154);
or U2221 (N_2221,N_2123,N_2105);
nand U2222 (N_2222,N_2188,N_2067);
and U2223 (N_2223,N_2142,N_2136);
or U2224 (N_2224,N_2171,N_2038);
xor U2225 (N_2225,N_2124,N_2126);
nand U2226 (N_2226,N_2179,N_2144);
nor U2227 (N_2227,N_2199,N_2146);
nand U2228 (N_2228,N_2049,N_2120);
or U2229 (N_2229,N_2014,N_2175);
nand U2230 (N_2230,N_2193,N_2010);
or U2231 (N_2231,N_2189,N_2039);
or U2232 (N_2232,N_2021,N_2156);
or U2233 (N_2233,N_2177,N_2090);
nand U2234 (N_2234,N_2036,N_2172);
xor U2235 (N_2235,N_2165,N_2050);
nand U2236 (N_2236,N_2075,N_2192);
and U2237 (N_2237,N_2109,N_2032);
nor U2238 (N_2238,N_2121,N_2088);
or U2239 (N_2239,N_2191,N_2079);
and U2240 (N_2240,N_2063,N_2106);
xnor U2241 (N_2241,N_2092,N_2137);
nor U2242 (N_2242,N_2040,N_2028);
nor U2243 (N_2243,N_2134,N_2187);
nor U2244 (N_2244,N_2005,N_2167);
or U2245 (N_2245,N_2119,N_2150);
or U2246 (N_2246,N_2197,N_2066);
xor U2247 (N_2247,N_2033,N_2046);
or U2248 (N_2248,N_2013,N_2152);
nor U2249 (N_2249,N_2007,N_2198);
nand U2250 (N_2250,N_2009,N_2031);
and U2251 (N_2251,N_2084,N_2099);
xor U2252 (N_2252,N_2195,N_2174);
nand U2253 (N_2253,N_2110,N_2026);
and U2254 (N_2254,N_2065,N_2115);
and U2255 (N_2255,N_2035,N_2054);
nand U2256 (N_2256,N_2183,N_2022);
nor U2257 (N_2257,N_2045,N_2176);
nor U2258 (N_2258,N_2168,N_2024);
xor U2259 (N_2259,N_2186,N_2089);
nor U2260 (N_2260,N_2161,N_2116);
xnor U2261 (N_2261,N_2091,N_2044);
nor U2262 (N_2262,N_2104,N_2008);
and U2263 (N_2263,N_2100,N_2057);
nor U2264 (N_2264,N_2082,N_2166);
xor U2265 (N_2265,N_2087,N_2141);
nor U2266 (N_2266,N_2162,N_2157);
nor U2267 (N_2267,N_2093,N_2078);
nor U2268 (N_2268,N_2029,N_2149);
or U2269 (N_2269,N_2061,N_2023);
and U2270 (N_2270,N_2056,N_2080);
and U2271 (N_2271,N_2059,N_2133);
nor U2272 (N_2272,N_2068,N_2012);
xor U2273 (N_2273,N_2098,N_2053);
or U2274 (N_2274,N_2041,N_2151);
or U2275 (N_2275,N_2107,N_2182);
and U2276 (N_2276,N_2085,N_2094);
xnor U2277 (N_2277,N_2160,N_2128);
or U2278 (N_2278,N_2064,N_2118);
or U2279 (N_2279,N_2178,N_2025);
xnor U2280 (N_2280,N_2073,N_2140);
and U2281 (N_2281,N_2129,N_2011);
or U2282 (N_2282,N_2159,N_2170);
and U2283 (N_2283,N_2051,N_2006);
xnor U2284 (N_2284,N_2111,N_2130);
nor U2285 (N_2285,N_2127,N_2173);
and U2286 (N_2286,N_2047,N_2017);
xnor U2287 (N_2287,N_2001,N_2131);
nor U2288 (N_2288,N_2062,N_2081);
and U2289 (N_2289,N_2052,N_2108);
nand U2290 (N_2290,N_2122,N_2145);
or U2291 (N_2291,N_2153,N_2097);
or U2292 (N_2292,N_2074,N_2181);
nor U2293 (N_2293,N_2071,N_2070);
and U2294 (N_2294,N_2019,N_2101);
or U2295 (N_2295,N_2055,N_2020);
or U2296 (N_2296,N_2112,N_2027);
xnor U2297 (N_2297,N_2194,N_2060);
or U2298 (N_2298,N_2138,N_2190);
or U2299 (N_2299,N_2132,N_2117);
nor U2300 (N_2300,N_2041,N_2014);
nor U2301 (N_2301,N_2091,N_2036);
or U2302 (N_2302,N_2007,N_2195);
or U2303 (N_2303,N_2081,N_2174);
or U2304 (N_2304,N_2003,N_2083);
or U2305 (N_2305,N_2080,N_2092);
or U2306 (N_2306,N_2138,N_2147);
or U2307 (N_2307,N_2163,N_2042);
nor U2308 (N_2308,N_2046,N_2029);
xnor U2309 (N_2309,N_2062,N_2143);
xnor U2310 (N_2310,N_2094,N_2110);
and U2311 (N_2311,N_2050,N_2035);
nand U2312 (N_2312,N_2150,N_2117);
nand U2313 (N_2313,N_2060,N_2014);
nand U2314 (N_2314,N_2089,N_2158);
or U2315 (N_2315,N_2003,N_2154);
or U2316 (N_2316,N_2120,N_2192);
nand U2317 (N_2317,N_2197,N_2073);
and U2318 (N_2318,N_2042,N_2089);
and U2319 (N_2319,N_2020,N_2159);
nand U2320 (N_2320,N_2193,N_2159);
nand U2321 (N_2321,N_2024,N_2161);
nor U2322 (N_2322,N_2128,N_2076);
xor U2323 (N_2323,N_2112,N_2186);
nor U2324 (N_2324,N_2198,N_2096);
xnor U2325 (N_2325,N_2183,N_2087);
xor U2326 (N_2326,N_2134,N_2196);
xor U2327 (N_2327,N_2003,N_2161);
or U2328 (N_2328,N_2084,N_2102);
or U2329 (N_2329,N_2084,N_2177);
or U2330 (N_2330,N_2135,N_2169);
nand U2331 (N_2331,N_2001,N_2050);
nor U2332 (N_2332,N_2155,N_2148);
and U2333 (N_2333,N_2132,N_2023);
nand U2334 (N_2334,N_2108,N_2137);
nor U2335 (N_2335,N_2003,N_2126);
nor U2336 (N_2336,N_2056,N_2032);
nand U2337 (N_2337,N_2154,N_2011);
and U2338 (N_2338,N_2022,N_2090);
nand U2339 (N_2339,N_2166,N_2063);
and U2340 (N_2340,N_2150,N_2136);
nor U2341 (N_2341,N_2037,N_2126);
nand U2342 (N_2342,N_2084,N_2157);
and U2343 (N_2343,N_2198,N_2175);
xnor U2344 (N_2344,N_2189,N_2083);
nor U2345 (N_2345,N_2137,N_2008);
nand U2346 (N_2346,N_2153,N_2118);
and U2347 (N_2347,N_2091,N_2195);
and U2348 (N_2348,N_2143,N_2112);
nor U2349 (N_2349,N_2057,N_2122);
nand U2350 (N_2350,N_2068,N_2124);
or U2351 (N_2351,N_2018,N_2019);
nand U2352 (N_2352,N_2093,N_2109);
nand U2353 (N_2353,N_2182,N_2071);
nor U2354 (N_2354,N_2155,N_2143);
or U2355 (N_2355,N_2165,N_2116);
and U2356 (N_2356,N_2046,N_2153);
nor U2357 (N_2357,N_2115,N_2127);
or U2358 (N_2358,N_2151,N_2188);
nor U2359 (N_2359,N_2171,N_2088);
xor U2360 (N_2360,N_2127,N_2162);
and U2361 (N_2361,N_2169,N_2137);
nor U2362 (N_2362,N_2129,N_2196);
and U2363 (N_2363,N_2081,N_2017);
xnor U2364 (N_2364,N_2052,N_2148);
or U2365 (N_2365,N_2068,N_2171);
or U2366 (N_2366,N_2110,N_2181);
and U2367 (N_2367,N_2013,N_2092);
and U2368 (N_2368,N_2106,N_2001);
nor U2369 (N_2369,N_2077,N_2011);
nor U2370 (N_2370,N_2153,N_2168);
nor U2371 (N_2371,N_2175,N_2117);
and U2372 (N_2372,N_2067,N_2053);
or U2373 (N_2373,N_2073,N_2059);
and U2374 (N_2374,N_2148,N_2191);
nor U2375 (N_2375,N_2102,N_2092);
or U2376 (N_2376,N_2193,N_2064);
nor U2377 (N_2377,N_2072,N_2169);
xnor U2378 (N_2378,N_2046,N_2134);
and U2379 (N_2379,N_2079,N_2165);
or U2380 (N_2380,N_2099,N_2112);
xor U2381 (N_2381,N_2001,N_2101);
nand U2382 (N_2382,N_2042,N_2142);
and U2383 (N_2383,N_2048,N_2145);
or U2384 (N_2384,N_2032,N_2073);
or U2385 (N_2385,N_2056,N_2047);
nand U2386 (N_2386,N_2051,N_2198);
and U2387 (N_2387,N_2153,N_2005);
nor U2388 (N_2388,N_2007,N_2060);
nor U2389 (N_2389,N_2062,N_2057);
nor U2390 (N_2390,N_2119,N_2009);
nor U2391 (N_2391,N_2052,N_2104);
or U2392 (N_2392,N_2059,N_2084);
or U2393 (N_2393,N_2168,N_2013);
xor U2394 (N_2394,N_2178,N_2146);
nand U2395 (N_2395,N_2054,N_2123);
or U2396 (N_2396,N_2025,N_2122);
or U2397 (N_2397,N_2120,N_2123);
nor U2398 (N_2398,N_2032,N_2030);
nand U2399 (N_2399,N_2174,N_2170);
xor U2400 (N_2400,N_2230,N_2269);
nor U2401 (N_2401,N_2323,N_2360);
nand U2402 (N_2402,N_2305,N_2262);
nor U2403 (N_2403,N_2319,N_2341);
xor U2404 (N_2404,N_2316,N_2216);
or U2405 (N_2405,N_2244,N_2368);
nor U2406 (N_2406,N_2376,N_2204);
nand U2407 (N_2407,N_2300,N_2338);
nand U2408 (N_2408,N_2245,N_2304);
and U2409 (N_2409,N_2223,N_2330);
and U2410 (N_2410,N_2308,N_2201);
or U2411 (N_2411,N_2353,N_2200);
or U2412 (N_2412,N_2354,N_2255);
or U2413 (N_2413,N_2345,N_2253);
nand U2414 (N_2414,N_2218,N_2361);
or U2415 (N_2415,N_2373,N_2347);
nor U2416 (N_2416,N_2282,N_2388);
nor U2417 (N_2417,N_2352,N_2369);
and U2418 (N_2418,N_2326,N_2383);
nor U2419 (N_2419,N_2217,N_2348);
nor U2420 (N_2420,N_2257,N_2298);
nor U2421 (N_2421,N_2233,N_2237);
or U2422 (N_2422,N_2329,N_2213);
nand U2423 (N_2423,N_2264,N_2333);
or U2424 (N_2424,N_2306,N_2232);
or U2425 (N_2425,N_2251,N_2292);
xor U2426 (N_2426,N_2349,N_2331);
xor U2427 (N_2427,N_2343,N_2210);
and U2428 (N_2428,N_2309,N_2320);
xor U2429 (N_2429,N_2211,N_2364);
and U2430 (N_2430,N_2248,N_2208);
xor U2431 (N_2431,N_2278,N_2273);
nor U2432 (N_2432,N_2385,N_2327);
or U2433 (N_2433,N_2214,N_2365);
or U2434 (N_2434,N_2382,N_2293);
nor U2435 (N_2435,N_2272,N_2342);
or U2436 (N_2436,N_2259,N_2283);
and U2437 (N_2437,N_2243,N_2377);
nor U2438 (N_2438,N_2371,N_2275);
nor U2439 (N_2439,N_2266,N_2398);
nand U2440 (N_2440,N_2378,N_2222);
xor U2441 (N_2441,N_2337,N_2241);
xor U2442 (N_2442,N_2209,N_2286);
xor U2443 (N_2443,N_2386,N_2372);
nand U2444 (N_2444,N_2261,N_2399);
nand U2445 (N_2445,N_2226,N_2370);
nor U2446 (N_2446,N_2393,N_2307);
nand U2447 (N_2447,N_2271,N_2231);
xnor U2448 (N_2448,N_2351,N_2202);
and U2449 (N_2449,N_2362,N_2205);
xor U2450 (N_2450,N_2215,N_2284);
or U2451 (N_2451,N_2287,N_2391);
nor U2452 (N_2452,N_2274,N_2260);
nor U2453 (N_2453,N_2355,N_2268);
and U2454 (N_2454,N_2270,N_2297);
nand U2455 (N_2455,N_2240,N_2313);
nand U2456 (N_2456,N_2367,N_2350);
or U2457 (N_2457,N_2267,N_2375);
nor U2458 (N_2458,N_2390,N_2289);
and U2459 (N_2459,N_2249,N_2285);
and U2460 (N_2460,N_2225,N_2247);
and U2461 (N_2461,N_2280,N_2258);
and U2462 (N_2462,N_2265,N_2238);
and U2463 (N_2463,N_2229,N_2392);
nand U2464 (N_2464,N_2325,N_2318);
nor U2465 (N_2465,N_2314,N_2334);
nand U2466 (N_2466,N_2221,N_2328);
nand U2467 (N_2467,N_2379,N_2219);
or U2468 (N_2468,N_2339,N_2374);
nand U2469 (N_2469,N_2358,N_2279);
nand U2470 (N_2470,N_2332,N_2394);
or U2471 (N_2471,N_2281,N_2228);
and U2472 (N_2472,N_2389,N_2324);
nor U2473 (N_2473,N_2227,N_2336);
nand U2474 (N_2474,N_2224,N_2397);
and U2475 (N_2475,N_2234,N_2288);
and U2476 (N_2476,N_2335,N_2359);
and U2477 (N_2477,N_2203,N_2296);
nor U2478 (N_2478,N_2239,N_2246);
nor U2479 (N_2479,N_2346,N_2312);
xor U2480 (N_2480,N_2256,N_2387);
nor U2481 (N_2481,N_2366,N_2276);
nor U2482 (N_2482,N_2380,N_2220);
nor U2483 (N_2483,N_2254,N_2363);
xnor U2484 (N_2484,N_2277,N_2322);
and U2485 (N_2485,N_2301,N_2340);
and U2486 (N_2486,N_2252,N_2395);
xnor U2487 (N_2487,N_2212,N_2381);
xnor U2488 (N_2488,N_2242,N_2303);
or U2489 (N_2489,N_2299,N_2294);
nor U2490 (N_2490,N_2315,N_2302);
nand U2491 (N_2491,N_2384,N_2235);
nand U2492 (N_2492,N_2295,N_2357);
nand U2493 (N_2493,N_2396,N_2207);
and U2494 (N_2494,N_2321,N_2290);
nor U2495 (N_2495,N_2311,N_2263);
nor U2496 (N_2496,N_2236,N_2310);
nand U2497 (N_2497,N_2291,N_2250);
nand U2498 (N_2498,N_2356,N_2206);
or U2499 (N_2499,N_2344,N_2317);
xnor U2500 (N_2500,N_2357,N_2371);
and U2501 (N_2501,N_2396,N_2264);
nand U2502 (N_2502,N_2237,N_2343);
nand U2503 (N_2503,N_2253,N_2228);
and U2504 (N_2504,N_2337,N_2310);
nor U2505 (N_2505,N_2282,N_2296);
and U2506 (N_2506,N_2376,N_2238);
or U2507 (N_2507,N_2340,N_2303);
or U2508 (N_2508,N_2238,N_2322);
nor U2509 (N_2509,N_2292,N_2276);
nor U2510 (N_2510,N_2325,N_2352);
nor U2511 (N_2511,N_2253,N_2214);
or U2512 (N_2512,N_2352,N_2310);
and U2513 (N_2513,N_2337,N_2346);
nor U2514 (N_2514,N_2336,N_2391);
xor U2515 (N_2515,N_2241,N_2266);
nand U2516 (N_2516,N_2343,N_2360);
xnor U2517 (N_2517,N_2228,N_2238);
xnor U2518 (N_2518,N_2369,N_2223);
nand U2519 (N_2519,N_2242,N_2233);
xor U2520 (N_2520,N_2399,N_2353);
xor U2521 (N_2521,N_2328,N_2274);
and U2522 (N_2522,N_2302,N_2204);
or U2523 (N_2523,N_2219,N_2322);
nor U2524 (N_2524,N_2370,N_2358);
xnor U2525 (N_2525,N_2205,N_2206);
xor U2526 (N_2526,N_2377,N_2226);
nor U2527 (N_2527,N_2268,N_2305);
nand U2528 (N_2528,N_2331,N_2254);
or U2529 (N_2529,N_2343,N_2321);
xnor U2530 (N_2530,N_2251,N_2206);
nand U2531 (N_2531,N_2264,N_2339);
nand U2532 (N_2532,N_2201,N_2279);
xnor U2533 (N_2533,N_2325,N_2285);
nor U2534 (N_2534,N_2247,N_2397);
and U2535 (N_2535,N_2344,N_2298);
xor U2536 (N_2536,N_2282,N_2319);
nand U2537 (N_2537,N_2307,N_2223);
xor U2538 (N_2538,N_2390,N_2353);
or U2539 (N_2539,N_2349,N_2225);
xor U2540 (N_2540,N_2306,N_2337);
and U2541 (N_2541,N_2337,N_2351);
xnor U2542 (N_2542,N_2345,N_2364);
nor U2543 (N_2543,N_2216,N_2342);
and U2544 (N_2544,N_2331,N_2394);
and U2545 (N_2545,N_2372,N_2295);
nor U2546 (N_2546,N_2242,N_2326);
nor U2547 (N_2547,N_2257,N_2247);
nand U2548 (N_2548,N_2315,N_2337);
and U2549 (N_2549,N_2215,N_2286);
nor U2550 (N_2550,N_2210,N_2202);
nand U2551 (N_2551,N_2266,N_2230);
nand U2552 (N_2552,N_2371,N_2382);
nand U2553 (N_2553,N_2364,N_2279);
or U2554 (N_2554,N_2298,N_2280);
nor U2555 (N_2555,N_2210,N_2298);
or U2556 (N_2556,N_2353,N_2328);
xor U2557 (N_2557,N_2394,N_2303);
nand U2558 (N_2558,N_2383,N_2202);
or U2559 (N_2559,N_2238,N_2384);
or U2560 (N_2560,N_2339,N_2242);
xnor U2561 (N_2561,N_2223,N_2285);
and U2562 (N_2562,N_2378,N_2390);
or U2563 (N_2563,N_2345,N_2348);
and U2564 (N_2564,N_2397,N_2311);
and U2565 (N_2565,N_2220,N_2350);
nor U2566 (N_2566,N_2246,N_2334);
or U2567 (N_2567,N_2376,N_2288);
xor U2568 (N_2568,N_2264,N_2244);
xor U2569 (N_2569,N_2252,N_2241);
nor U2570 (N_2570,N_2298,N_2365);
and U2571 (N_2571,N_2391,N_2257);
or U2572 (N_2572,N_2365,N_2284);
or U2573 (N_2573,N_2247,N_2390);
xnor U2574 (N_2574,N_2380,N_2231);
or U2575 (N_2575,N_2352,N_2394);
or U2576 (N_2576,N_2386,N_2203);
xor U2577 (N_2577,N_2384,N_2299);
nor U2578 (N_2578,N_2323,N_2320);
nor U2579 (N_2579,N_2273,N_2220);
or U2580 (N_2580,N_2396,N_2297);
nor U2581 (N_2581,N_2239,N_2232);
xnor U2582 (N_2582,N_2312,N_2270);
and U2583 (N_2583,N_2200,N_2373);
xnor U2584 (N_2584,N_2227,N_2396);
nand U2585 (N_2585,N_2393,N_2395);
nor U2586 (N_2586,N_2314,N_2246);
nand U2587 (N_2587,N_2266,N_2319);
nand U2588 (N_2588,N_2312,N_2389);
nand U2589 (N_2589,N_2200,N_2273);
xnor U2590 (N_2590,N_2248,N_2225);
and U2591 (N_2591,N_2391,N_2270);
nor U2592 (N_2592,N_2285,N_2309);
nor U2593 (N_2593,N_2369,N_2306);
and U2594 (N_2594,N_2220,N_2281);
nand U2595 (N_2595,N_2300,N_2263);
nand U2596 (N_2596,N_2205,N_2357);
xnor U2597 (N_2597,N_2348,N_2229);
or U2598 (N_2598,N_2371,N_2389);
nand U2599 (N_2599,N_2353,N_2387);
nand U2600 (N_2600,N_2418,N_2509);
nand U2601 (N_2601,N_2408,N_2569);
nand U2602 (N_2602,N_2483,N_2445);
and U2603 (N_2603,N_2546,N_2528);
xor U2604 (N_2604,N_2436,N_2543);
nand U2605 (N_2605,N_2488,N_2556);
nor U2606 (N_2606,N_2478,N_2596);
xnor U2607 (N_2607,N_2499,N_2512);
or U2608 (N_2608,N_2544,N_2498);
and U2609 (N_2609,N_2449,N_2443);
and U2610 (N_2610,N_2561,N_2555);
nand U2611 (N_2611,N_2554,N_2574);
or U2612 (N_2612,N_2417,N_2513);
nand U2613 (N_2613,N_2584,N_2414);
xnor U2614 (N_2614,N_2425,N_2593);
nand U2615 (N_2615,N_2598,N_2567);
and U2616 (N_2616,N_2494,N_2500);
nand U2617 (N_2617,N_2505,N_2429);
and U2618 (N_2618,N_2434,N_2407);
nor U2619 (N_2619,N_2573,N_2591);
nor U2620 (N_2620,N_2542,N_2475);
xnor U2621 (N_2621,N_2502,N_2508);
or U2622 (N_2622,N_2422,N_2531);
xnor U2623 (N_2623,N_2454,N_2549);
nor U2624 (N_2624,N_2452,N_2537);
xnor U2625 (N_2625,N_2575,N_2565);
nand U2626 (N_2626,N_2440,N_2446);
and U2627 (N_2627,N_2472,N_2473);
nor U2628 (N_2628,N_2587,N_2552);
and U2629 (N_2629,N_2480,N_2506);
nand U2630 (N_2630,N_2571,N_2486);
or U2631 (N_2631,N_2496,N_2525);
xnor U2632 (N_2632,N_2438,N_2507);
xor U2633 (N_2633,N_2423,N_2403);
nand U2634 (N_2634,N_2557,N_2435);
nand U2635 (N_2635,N_2419,N_2595);
nor U2636 (N_2636,N_2479,N_2402);
nor U2637 (N_2637,N_2433,N_2464);
or U2638 (N_2638,N_2437,N_2474);
nor U2639 (N_2639,N_2448,N_2583);
or U2640 (N_2640,N_2487,N_2444);
xor U2641 (N_2641,N_2468,N_2580);
or U2642 (N_2642,N_2431,N_2550);
or U2643 (N_2643,N_2497,N_2477);
nor U2644 (N_2644,N_2578,N_2430);
nor U2645 (N_2645,N_2576,N_2482);
and U2646 (N_2646,N_2427,N_2484);
or U2647 (N_2647,N_2491,N_2533);
xnor U2648 (N_2648,N_2517,N_2453);
nand U2649 (N_2649,N_2539,N_2585);
or U2650 (N_2650,N_2404,N_2426);
nor U2651 (N_2651,N_2441,N_2566);
or U2652 (N_2652,N_2467,N_2503);
nor U2653 (N_2653,N_2412,N_2493);
nor U2654 (N_2654,N_2461,N_2504);
or U2655 (N_2655,N_2447,N_2523);
nor U2656 (N_2656,N_2495,N_2589);
nor U2657 (N_2657,N_2492,N_2471);
nand U2658 (N_2658,N_2529,N_2462);
xnor U2659 (N_2659,N_2501,N_2424);
and U2660 (N_2660,N_2451,N_2560);
or U2661 (N_2661,N_2455,N_2421);
nand U2662 (N_2662,N_2463,N_2410);
or U2663 (N_2663,N_2526,N_2545);
and U2664 (N_2664,N_2551,N_2553);
nand U2665 (N_2665,N_2439,N_2538);
nand U2666 (N_2666,N_2562,N_2416);
nor U2667 (N_2667,N_2586,N_2515);
and U2668 (N_2668,N_2428,N_2522);
and U2669 (N_2669,N_2465,N_2442);
xnor U2670 (N_2670,N_2476,N_2524);
and U2671 (N_2671,N_2572,N_2582);
nor U2672 (N_2672,N_2588,N_2469);
nor U2673 (N_2673,N_2568,N_2579);
nor U2674 (N_2674,N_2409,N_2548);
xnor U2675 (N_2675,N_2456,N_2563);
and U2676 (N_2676,N_2481,N_2534);
nor U2677 (N_2677,N_2547,N_2536);
nor U2678 (N_2678,N_2581,N_2519);
nor U2679 (N_2679,N_2532,N_2516);
nor U2680 (N_2680,N_2489,N_2420);
or U2681 (N_2681,N_2450,N_2599);
nand U2682 (N_2682,N_2485,N_2527);
or U2683 (N_2683,N_2540,N_2535);
nand U2684 (N_2684,N_2406,N_2401);
xor U2685 (N_2685,N_2460,N_2530);
nand U2686 (N_2686,N_2514,N_2510);
nor U2687 (N_2687,N_2592,N_2559);
nand U2688 (N_2688,N_2490,N_2564);
nand U2689 (N_2689,N_2411,N_2558);
and U2690 (N_2690,N_2597,N_2405);
xnor U2691 (N_2691,N_2466,N_2413);
nor U2692 (N_2692,N_2594,N_2400);
nor U2693 (N_2693,N_2415,N_2432);
and U2694 (N_2694,N_2570,N_2457);
or U2695 (N_2695,N_2511,N_2470);
nor U2696 (N_2696,N_2590,N_2520);
nor U2697 (N_2697,N_2541,N_2577);
nand U2698 (N_2698,N_2459,N_2458);
xnor U2699 (N_2699,N_2521,N_2518);
xnor U2700 (N_2700,N_2560,N_2547);
or U2701 (N_2701,N_2422,N_2569);
xor U2702 (N_2702,N_2484,N_2469);
and U2703 (N_2703,N_2450,N_2524);
nand U2704 (N_2704,N_2471,N_2533);
nor U2705 (N_2705,N_2527,N_2585);
or U2706 (N_2706,N_2512,N_2422);
nor U2707 (N_2707,N_2409,N_2505);
nand U2708 (N_2708,N_2440,N_2535);
or U2709 (N_2709,N_2551,N_2572);
and U2710 (N_2710,N_2597,N_2510);
or U2711 (N_2711,N_2512,N_2559);
or U2712 (N_2712,N_2576,N_2542);
nand U2713 (N_2713,N_2540,N_2573);
xnor U2714 (N_2714,N_2509,N_2444);
and U2715 (N_2715,N_2476,N_2464);
xor U2716 (N_2716,N_2561,N_2511);
and U2717 (N_2717,N_2552,N_2516);
nor U2718 (N_2718,N_2533,N_2420);
nor U2719 (N_2719,N_2461,N_2559);
or U2720 (N_2720,N_2425,N_2539);
nand U2721 (N_2721,N_2464,N_2461);
nor U2722 (N_2722,N_2574,N_2481);
and U2723 (N_2723,N_2415,N_2572);
nor U2724 (N_2724,N_2445,N_2489);
or U2725 (N_2725,N_2457,N_2575);
xnor U2726 (N_2726,N_2467,N_2588);
or U2727 (N_2727,N_2573,N_2471);
nand U2728 (N_2728,N_2473,N_2599);
nor U2729 (N_2729,N_2504,N_2437);
nor U2730 (N_2730,N_2559,N_2464);
nor U2731 (N_2731,N_2436,N_2560);
xnor U2732 (N_2732,N_2441,N_2585);
xnor U2733 (N_2733,N_2442,N_2408);
nor U2734 (N_2734,N_2499,N_2583);
nand U2735 (N_2735,N_2519,N_2428);
xor U2736 (N_2736,N_2498,N_2405);
and U2737 (N_2737,N_2405,N_2427);
and U2738 (N_2738,N_2586,N_2555);
and U2739 (N_2739,N_2444,N_2571);
and U2740 (N_2740,N_2595,N_2500);
and U2741 (N_2741,N_2476,N_2549);
or U2742 (N_2742,N_2480,N_2564);
nor U2743 (N_2743,N_2548,N_2560);
xnor U2744 (N_2744,N_2502,N_2550);
or U2745 (N_2745,N_2595,N_2406);
or U2746 (N_2746,N_2477,N_2553);
or U2747 (N_2747,N_2537,N_2565);
xor U2748 (N_2748,N_2412,N_2517);
and U2749 (N_2749,N_2465,N_2506);
xnor U2750 (N_2750,N_2502,N_2488);
nor U2751 (N_2751,N_2568,N_2534);
xnor U2752 (N_2752,N_2567,N_2538);
or U2753 (N_2753,N_2507,N_2493);
nand U2754 (N_2754,N_2513,N_2588);
xor U2755 (N_2755,N_2598,N_2482);
nand U2756 (N_2756,N_2587,N_2551);
nand U2757 (N_2757,N_2552,N_2483);
and U2758 (N_2758,N_2509,N_2482);
and U2759 (N_2759,N_2508,N_2446);
or U2760 (N_2760,N_2410,N_2586);
nor U2761 (N_2761,N_2547,N_2569);
xor U2762 (N_2762,N_2596,N_2572);
xor U2763 (N_2763,N_2435,N_2529);
and U2764 (N_2764,N_2432,N_2542);
xnor U2765 (N_2765,N_2419,N_2456);
xor U2766 (N_2766,N_2458,N_2549);
nor U2767 (N_2767,N_2537,N_2450);
xor U2768 (N_2768,N_2427,N_2567);
nand U2769 (N_2769,N_2581,N_2464);
xor U2770 (N_2770,N_2497,N_2505);
nand U2771 (N_2771,N_2525,N_2535);
xor U2772 (N_2772,N_2599,N_2568);
nor U2773 (N_2773,N_2401,N_2521);
nand U2774 (N_2774,N_2495,N_2466);
and U2775 (N_2775,N_2481,N_2551);
or U2776 (N_2776,N_2414,N_2401);
or U2777 (N_2777,N_2524,N_2417);
and U2778 (N_2778,N_2598,N_2443);
and U2779 (N_2779,N_2428,N_2575);
nor U2780 (N_2780,N_2554,N_2542);
xnor U2781 (N_2781,N_2531,N_2549);
or U2782 (N_2782,N_2569,N_2564);
nand U2783 (N_2783,N_2593,N_2567);
xnor U2784 (N_2784,N_2494,N_2568);
and U2785 (N_2785,N_2484,N_2443);
nor U2786 (N_2786,N_2596,N_2459);
or U2787 (N_2787,N_2497,N_2561);
nor U2788 (N_2788,N_2568,N_2524);
xnor U2789 (N_2789,N_2531,N_2519);
xor U2790 (N_2790,N_2401,N_2498);
or U2791 (N_2791,N_2542,N_2424);
xor U2792 (N_2792,N_2466,N_2436);
and U2793 (N_2793,N_2413,N_2423);
nor U2794 (N_2794,N_2415,N_2402);
xnor U2795 (N_2795,N_2424,N_2508);
or U2796 (N_2796,N_2501,N_2444);
and U2797 (N_2797,N_2579,N_2553);
and U2798 (N_2798,N_2463,N_2445);
nor U2799 (N_2799,N_2552,N_2519);
xnor U2800 (N_2800,N_2660,N_2776);
xnor U2801 (N_2801,N_2671,N_2606);
nand U2802 (N_2802,N_2792,N_2691);
nor U2803 (N_2803,N_2779,N_2760);
and U2804 (N_2804,N_2688,N_2778);
or U2805 (N_2805,N_2617,N_2716);
and U2806 (N_2806,N_2708,N_2649);
nand U2807 (N_2807,N_2668,N_2678);
nor U2808 (N_2808,N_2620,N_2780);
and U2809 (N_2809,N_2629,N_2740);
nand U2810 (N_2810,N_2648,N_2765);
xnor U2811 (N_2811,N_2682,N_2784);
nand U2812 (N_2812,N_2674,N_2794);
nor U2813 (N_2813,N_2712,N_2622);
or U2814 (N_2814,N_2696,N_2675);
and U2815 (N_2815,N_2761,N_2613);
xnor U2816 (N_2816,N_2702,N_2656);
xnor U2817 (N_2817,N_2640,N_2769);
nand U2818 (N_2818,N_2681,N_2686);
xor U2819 (N_2819,N_2639,N_2717);
and U2820 (N_2820,N_2723,N_2735);
or U2821 (N_2821,N_2684,N_2755);
nand U2822 (N_2822,N_2771,N_2614);
or U2823 (N_2823,N_2752,N_2786);
or U2824 (N_2824,N_2793,N_2698);
nand U2825 (N_2825,N_2791,N_2783);
nand U2826 (N_2826,N_2730,N_2643);
nand U2827 (N_2827,N_2722,N_2676);
nand U2828 (N_2828,N_2706,N_2633);
nor U2829 (N_2829,N_2677,N_2738);
and U2830 (N_2830,N_2625,N_2713);
xnor U2831 (N_2831,N_2608,N_2766);
nand U2832 (N_2832,N_2618,N_2630);
nor U2833 (N_2833,N_2744,N_2724);
and U2834 (N_2834,N_2709,N_2754);
or U2835 (N_2835,N_2733,N_2699);
nor U2836 (N_2836,N_2601,N_2749);
nor U2837 (N_2837,N_2609,N_2720);
xor U2838 (N_2838,N_2690,N_2612);
xnor U2839 (N_2839,N_2741,N_2697);
or U2840 (N_2840,N_2634,N_2718);
nor U2841 (N_2841,N_2687,N_2750);
nand U2842 (N_2842,N_2669,N_2731);
nand U2843 (N_2843,N_2747,N_2619);
nand U2844 (N_2844,N_2727,N_2745);
nand U2845 (N_2845,N_2781,N_2683);
nor U2846 (N_2846,N_2743,N_2635);
or U2847 (N_2847,N_2616,N_2611);
nor U2848 (N_2848,N_2788,N_2605);
or U2849 (N_2849,N_2725,N_2728);
nand U2850 (N_2850,N_2645,N_2650);
nor U2851 (N_2851,N_2666,N_2600);
nor U2852 (N_2852,N_2607,N_2695);
or U2853 (N_2853,N_2644,N_2785);
nor U2854 (N_2854,N_2654,N_2604);
and U2855 (N_2855,N_2782,N_2646);
and U2856 (N_2856,N_2651,N_2753);
or U2857 (N_2857,N_2653,N_2662);
nor U2858 (N_2858,N_2758,N_2719);
nand U2859 (N_2859,N_2770,N_2773);
nand U2860 (N_2860,N_2729,N_2715);
nand U2861 (N_2861,N_2700,N_2726);
nand U2862 (N_2862,N_2667,N_2799);
nor U2863 (N_2863,N_2734,N_2721);
or U2864 (N_2864,N_2703,N_2624);
xnor U2865 (N_2865,N_2701,N_2777);
xor U2866 (N_2866,N_2672,N_2775);
or U2867 (N_2867,N_2637,N_2796);
and U2868 (N_2868,N_2751,N_2772);
nand U2869 (N_2869,N_2685,N_2659);
or U2870 (N_2870,N_2710,N_2638);
nand U2871 (N_2871,N_2665,N_2615);
nor U2872 (N_2872,N_2789,N_2642);
and U2873 (N_2873,N_2631,N_2705);
nor U2874 (N_2874,N_2657,N_2714);
or U2875 (N_2875,N_2647,N_2746);
or U2876 (N_2876,N_2787,N_2711);
or U2877 (N_2877,N_2680,N_2679);
nor U2878 (N_2878,N_2798,N_2602);
and U2879 (N_2879,N_2628,N_2693);
xnor U2880 (N_2880,N_2623,N_2768);
xor U2881 (N_2881,N_2655,N_2737);
or U2882 (N_2882,N_2663,N_2742);
nor U2883 (N_2883,N_2759,N_2652);
nand U2884 (N_2884,N_2664,N_2670);
or U2885 (N_2885,N_2795,N_2658);
and U2886 (N_2886,N_2797,N_2763);
or U2887 (N_2887,N_2732,N_2689);
nand U2888 (N_2888,N_2756,N_2692);
nand U2889 (N_2889,N_2757,N_2790);
or U2890 (N_2890,N_2627,N_2603);
nor U2891 (N_2891,N_2610,N_2739);
nor U2892 (N_2892,N_2636,N_2694);
or U2893 (N_2893,N_2626,N_2707);
nor U2894 (N_2894,N_2748,N_2641);
nand U2895 (N_2895,N_2621,N_2764);
or U2896 (N_2896,N_2767,N_2704);
and U2897 (N_2897,N_2774,N_2632);
nand U2898 (N_2898,N_2762,N_2661);
or U2899 (N_2899,N_2736,N_2673);
nor U2900 (N_2900,N_2724,N_2723);
and U2901 (N_2901,N_2743,N_2747);
xor U2902 (N_2902,N_2737,N_2636);
or U2903 (N_2903,N_2671,N_2791);
and U2904 (N_2904,N_2670,N_2739);
nor U2905 (N_2905,N_2751,N_2638);
or U2906 (N_2906,N_2664,N_2698);
nand U2907 (N_2907,N_2786,N_2638);
nor U2908 (N_2908,N_2680,N_2645);
and U2909 (N_2909,N_2731,N_2641);
xor U2910 (N_2910,N_2708,N_2790);
nor U2911 (N_2911,N_2637,N_2777);
or U2912 (N_2912,N_2798,N_2797);
xnor U2913 (N_2913,N_2624,N_2688);
nand U2914 (N_2914,N_2779,N_2654);
nor U2915 (N_2915,N_2752,N_2621);
and U2916 (N_2916,N_2780,N_2616);
nand U2917 (N_2917,N_2630,N_2745);
nand U2918 (N_2918,N_2709,N_2612);
xnor U2919 (N_2919,N_2605,N_2659);
nand U2920 (N_2920,N_2716,N_2631);
or U2921 (N_2921,N_2799,N_2671);
xnor U2922 (N_2922,N_2761,N_2777);
or U2923 (N_2923,N_2635,N_2631);
and U2924 (N_2924,N_2702,N_2614);
or U2925 (N_2925,N_2615,N_2626);
nor U2926 (N_2926,N_2764,N_2791);
xnor U2927 (N_2927,N_2646,N_2733);
or U2928 (N_2928,N_2624,N_2694);
nor U2929 (N_2929,N_2728,N_2701);
xnor U2930 (N_2930,N_2670,N_2790);
or U2931 (N_2931,N_2754,N_2738);
and U2932 (N_2932,N_2799,N_2752);
nand U2933 (N_2933,N_2700,N_2797);
or U2934 (N_2934,N_2745,N_2667);
xnor U2935 (N_2935,N_2756,N_2781);
nand U2936 (N_2936,N_2635,N_2608);
xnor U2937 (N_2937,N_2708,N_2776);
xor U2938 (N_2938,N_2782,N_2774);
and U2939 (N_2939,N_2653,N_2713);
or U2940 (N_2940,N_2688,N_2654);
xor U2941 (N_2941,N_2726,N_2629);
and U2942 (N_2942,N_2669,N_2658);
nand U2943 (N_2943,N_2677,N_2638);
nor U2944 (N_2944,N_2631,N_2698);
and U2945 (N_2945,N_2709,N_2750);
or U2946 (N_2946,N_2642,N_2628);
xor U2947 (N_2947,N_2603,N_2721);
nand U2948 (N_2948,N_2708,N_2696);
and U2949 (N_2949,N_2764,N_2731);
or U2950 (N_2950,N_2632,N_2764);
and U2951 (N_2951,N_2705,N_2760);
nor U2952 (N_2952,N_2688,N_2762);
and U2953 (N_2953,N_2720,N_2602);
and U2954 (N_2954,N_2626,N_2771);
nand U2955 (N_2955,N_2624,N_2797);
or U2956 (N_2956,N_2771,N_2684);
nor U2957 (N_2957,N_2651,N_2702);
nand U2958 (N_2958,N_2784,N_2724);
or U2959 (N_2959,N_2786,N_2619);
or U2960 (N_2960,N_2759,N_2742);
nand U2961 (N_2961,N_2782,N_2718);
xor U2962 (N_2962,N_2695,N_2625);
nor U2963 (N_2963,N_2747,N_2674);
xor U2964 (N_2964,N_2651,N_2628);
nand U2965 (N_2965,N_2613,N_2799);
or U2966 (N_2966,N_2797,N_2668);
xnor U2967 (N_2967,N_2754,N_2622);
nor U2968 (N_2968,N_2729,N_2609);
nor U2969 (N_2969,N_2793,N_2678);
and U2970 (N_2970,N_2631,N_2615);
nand U2971 (N_2971,N_2696,N_2710);
xor U2972 (N_2972,N_2615,N_2622);
nand U2973 (N_2973,N_2772,N_2656);
xnor U2974 (N_2974,N_2726,N_2756);
nand U2975 (N_2975,N_2790,N_2794);
and U2976 (N_2976,N_2617,N_2794);
xnor U2977 (N_2977,N_2707,N_2652);
nand U2978 (N_2978,N_2640,N_2638);
and U2979 (N_2979,N_2694,N_2679);
nor U2980 (N_2980,N_2759,N_2645);
xnor U2981 (N_2981,N_2690,N_2766);
or U2982 (N_2982,N_2751,N_2779);
and U2983 (N_2983,N_2660,N_2749);
or U2984 (N_2984,N_2799,N_2632);
nor U2985 (N_2985,N_2743,N_2628);
nor U2986 (N_2986,N_2764,N_2679);
nand U2987 (N_2987,N_2784,N_2701);
nand U2988 (N_2988,N_2780,N_2704);
xnor U2989 (N_2989,N_2736,N_2678);
xnor U2990 (N_2990,N_2755,N_2642);
or U2991 (N_2991,N_2702,N_2771);
nand U2992 (N_2992,N_2635,N_2629);
nand U2993 (N_2993,N_2697,N_2762);
and U2994 (N_2994,N_2782,N_2644);
nor U2995 (N_2995,N_2630,N_2738);
or U2996 (N_2996,N_2631,N_2763);
and U2997 (N_2997,N_2759,N_2704);
nor U2998 (N_2998,N_2752,N_2628);
xor U2999 (N_2999,N_2659,N_2654);
and U3000 (N_3000,N_2871,N_2852);
and U3001 (N_3001,N_2856,N_2888);
or U3002 (N_3002,N_2917,N_2859);
or U3003 (N_3003,N_2883,N_2849);
nand U3004 (N_3004,N_2900,N_2945);
nand U3005 (N_3005,N_2864,N_2861);
and U3006 (N_3006,N_2989,N_2869);
xor U3007 (N_3007,N_2826,N_2854);
and U3008 (N_3008,N_2802,N_2828);
nor U3009 (N_3009,N_2950,N_2960);
nor U3010 (N_3010,N_2927,N_2816);
nor U3011 (N_3011,N_2805,N_2990);
nand U3012 (N_3012,N_2902,N_2814);
xnor U3013 (N_3013,N_2812,N_2938);
xor U3014 (N_3014,N_2972,N_2839);
xor U3015 (N_3015,N_2890,N_2873);
nor U3016 (N_3016,N_2934,N_2949);
or U3017 (N_3017,N_2952,N_2892);
xnor U3018 (N_3018,N_2916,N_2863);
xnor U3019 (N_3019,N_2813,N_2983);
nand U3020 (N_3020,N_2842,N_2903);
xnor U3021 (N_3021,N_2884,N_2878);
and U3022 (N_3022,N_2844,N_2971);
nor U3023 (N_3023,N_2881,N_2875);
or U3024 (N_3024,N_2898,N_2882);
or U3025 (N_3025,N_2865,N_2885);
or U3026 (N_3026,N_2969,N_2820);
and U3027 (N_3027,N_2886,N_2845);
or U3028 (N_3028,N_2943,N_2906);
and U3029 (N_3029,N_2923,N_2921);
and U3030 (N_3030,N_2980,N_2880);
nor U3031 (N_3031,N_2981,N_2947);
and U3032 (N_3032,N_2841,N_2809);
and U3033 (N_3033,N_2996,N_2825);
nor U3034 (N_3034,N_2919,N_2939);
xor U3035 (N_3035,N_2922,N_2959);
nor U3036 (N_3036,N_2807,N_2867);
xor U3037 (N_3037,N_2932,N_2967);
and U3038 (N_3038,N_2979,N_2874);
or U3039 (N_3039,N_2870,N_2974);
nand U3040 (N_3040,N_2835,N_2905);
nand U3041 (N_3041,N_2817,N_2912);
nand U3042 (N_3042,N_2925,N_2926);
or U3043 (N_3043,N_2956,N_2909);
xnor U3044 (N_3044,N_2876,N_2963);
nor U3045 (N_3045,N_2953,N_2918);
nand U3046 (N_3046,N_2895,N_2958);
and U3047 (N_3047,N_2993,N_2935);
xor U3048 (N_3048,N_2868,N_2824);
and U3049 (N_3049,N_2964,N_2830);
or U3050 (N_3050,N_2995,N_2929);
nand U3051 (N_3051,N_2998,N_2977);
nand U3052 (N_3052,N_2911,N_2988);
and U3053 (N_3053,N_2847,N_2853);
nand U3054 (N_3054,N_2930,N_2818);
xor U3055 (N_3055,N_2833,N_2994);
nor U3056 (N_3056,N_2986,N_2848);
nand U3057 (N_3057,N_2931,N_2855);
or U3058 (N_3058,N_2941,N_2966);
or U3059 (N_3059,N_2999,N_2810);
or U3060 (N_3060,N_2862,N_2913);
nor U3061 (N_3061,N_2846,N_2924);
or U3062 (N_3062,N_2991,N_2928);
nor U3063 (N_3063,N_2891,N_2933);
and U3064 (N_3064,N_2879,N_2987);
nor U3065 (N_3065,N_2948,N_2978);
and U3066 (N_3066,N_2961,N_2965);
or U3067 (N_3067,N_2901,N_2985);
nor U3068 (N_3068,N_2975,N_2872);
nand U3069 (N_3069,N_2843,N_2866);
and U3070 (N_3070,N_2957,N_2942);
nand U3071 (N_3071,N_2815,N_2954);
nand U3072 (N_3072,N_2800,N_2822);
and U3073 (N_3073,N_2829,N_2887);
xnor U3074 (N_3074,N_2970,N_2857);
xnor U3075 (N_3075,N_2962,N_2946);
xnor U3076 (N_3076,N_2894,N_2889);
and U3077 (N_3077,N_2877,N_2915);
nand U3078 (N_3078,N_2803,N_2851);
nand U3079 (N_3079,N_2811,N_2937);
or U3080 (N_3080,N_2834,N_2808);
xnor U3081 (N_3081,N_2819,N_2801);
xnor U3082 (N_3082,N_2896,N_2836);
nor U3083 (N_3083,N_2860,N_2984);
or U3084 (N_3084,N_2832,N_2823);
or U3085 (N_3085,N_2955,N_2806);
xor U3086 (N_3086,N_2904,N_2858);
xor U3087 (N_3087,N_2893,N_2840);
or U3088 (N_3088,N_2976,N_2968);
or U3089 (N_3089,N_2982,N_2940);
and U3090 (N_3090,N_2951,N_2827);
xnor U3091 (N_3091,N_2997,N_2973);
xor U3092 (N_3092,N_2821,N_2897);
xnor U3093 (N_3093,N_2908,N_2992);
xor U3094 (N_3094,N_2944,N_2850);
or U3095 (N_3095,N_2920,N_2907);
and U3096 (N_3096,N_2837,N_2838);
and U3097 (N_3097,N_2804,N_2914);
nand U3098 (N_3098,N_2936,N_2831);
xor U3099 (N_3099,N_2899,N_2910);
xor U3100 (N_3100,N_2905,N_2971);
xor U3101 (N_3101,N_2875,N_2918);
nor U3102 (N_3102,N_2901,N_2804);
xor U3103 (N_3103,N_2990,N_2946);
nand U3104 (N_3104,N_2928,N_2897);
xnor U3105 (N_3105,N_2956,N_2908);
and U3106 (N_3106,N_2936,N_2914);
xor U3107 (N_3107,N_2931,N_2980);
or U3108 (N_3108,N_2903,N_2855);
and U3109 (N_3109,N_2941,N_2808);
xnor U3110 (N_3110,N_2944,N_2998);
xnor U3111 (N_3111,N_2862,N_2949);
nand U3112 (N_3112,N_2948,N_2827);
and U3113 (N_3113,N_2873,N_2834);
nand U3114 (N_3114,N_2831,N_2944);
or U3115 (N_3115,N_2865,N_2970);
xnor U3116 (N_3116,N_2997,N_2840);
and U3117 (N_3117,N_2966,N_2841);
and U3118 (N_3118,N_2817,N_2812);
nor U3119 (N_3119,N_2828,N_2980);
and U3120 (N_3120,N_2922,N_2839);
nor U3121 (N_3121,N_2802,N_2962);
and U3122 (N_3122,N_2836,N_2915);
nand U3123 (N_3123,N_2866,N_2845);
or U3124 (N_3124,N_2937,N_2938);
nor U3125 (N_3125,N_2923,N_2963);
or U3126 (N_3126,N_2959,N_2997);
xor U3127 (N_3127,N_2812,N_2839);
nand U3128 (N_3128,N_2881,N_2913);
and U3129 (N_3129,N_2802,N_2894);
or U3130 (N_3130,N_2814,N_2906);
nor U3131 (N_3131,N_2877,N_2815);
nor U3132 (N_3132,N_2846,N_2894);
and U3133 (N_3133,N_2995,N_2966);
or U3134 (N_3134,N_2960,N_2940);
and U3135 (N_3135,N_2868,N_2920);
nand U3136 (N_3136,N_2817,N_2937);
xnor U3137 (N_3137,N_2807,N_2861);
xor U3138 (N_3138,N_2960,N_2994);
xor U3139 (N_3139,N_2913,N_2839);
and U3140 (N_3140,N_2832,N_2898);
xnor U3141 (N_3141,N_2857,N_2845);
nor U3142 (N_3142,N_2876,N_2894);
nor U3143 (N_3143,N_2854,N_2880);
nor U3144 (N_3144,N_2896,N_2871);
nor U3145 (N_3145,N_2892,N_2932);
or U3146 (N_3146,N_2915,N_2980);
nand U3147 (N_3147,N_2876,N_2801);
nor U3148 (N_3148,N_2875,N_2998);
nor U3149 (N_3149,N_2953,N_2996);
or U3150 (N_3150,N_2870,N_2984);
and U3151 (N_3151,N_2909,N_2871);
or U3152 (N_3152,N_2921,N_2936);
nor U3153 (N_3153,N_2842,N_2978);
or U3154 (N_3154,N_2888,N_2855);
xnor U3155 (N_3155,N_2935,N_2945);
and U3156 (N_3156,N_2902,N_2919);
and U3157 (N_3157,N_2943,N_2965);
xor U3158 (N_3158,N_2859,N_2936);
and U3159 (N_3159,N_2836,N_2809);
or U3160 (N_3160,N_2820,N_2939);
nand U3161 (N_3161,N_2963,N_2955);
or U3162 (N_3162,N_2958,N_2839);
nor U3163 (N_3163,N_2977,N_2920);
and U3164 (N_3164,N_2965,N_2895);
and U3165 (N_3165,N_2847,N_2896);
or U3166 (N_3166,N_2824,N_2869);
or U3167 (N_3167,N_2874,N_2901);
or U3168 (N_3168,N_2811,N_2911);
xnor U3169 (N_3169,N_2914,N_2988);
nand U3170 (N_3170,N_2940,N_2801);
nor U3171 (N_3171,N_2805,N_2820);
and U3172 (N_3172,N_2871,N_2938);
and U3173 (N_3173,N_2828,N_2831);
or U3174 (N_3174,N_2919,N_2914);
or U3175 (N_3175,N_2821,N_2996);
and U3176 (N_3176,N_2967,N_2908);
nor U3177 (N_3177,N_2911,N_2907);
nand U3178 (N_3178,N_2911,N_2850);
nand U3179 (N_3179,N_2897,N_2905);
or U3180 (N_3180,N_2922,N_2979);
xor U3181 (N_3181,N_2882,N_2970);
xnor U3182 (N_3182,N_2807,N_2999);
xor U3183 (N_3183,N_2948,N_2911);
or U3184 (N_3184,N_2845,N_2981);
nand U3185 (N_3185,N_2876,N_2925);
and U3186 (N_3186,N_2830,N_2924);
nor U3187 (N_3187,N_2963,N_2956);
and U3188 (N_3188,N_2877,N_2958);
nand U3189 (N_3189,N_2827,N_2904);
nor U3190 (N_3190,N_2986,N_2917);
nand U3191 (N_3191,N_2947,N_2906);
or U3192 (N_3192,N_2835,N_2948);
and U3193 (N_3193,N_2896,N_2917);
xor U3194 (N_3194,N_2842,N_2894);
xnor U3195 (N_3195,N_2980,N_2994);
and U3196 (N_3196,N_2826,N_2852);
xor U3197 (N_3197,N_2961,N_2929);
or U3198 (N_3198,N_2822,N_2992);
nand U3199 (N_3199,N_2886,N_2958);
or U3200 (N_3200,N_3058,N_3143);
nand U3201 (N_3201,N_3067,N_3023);
nand U3202 (N_3202,N_3104,N_3073);
and U3203 (N_3203,N_3189,N_3030);
or U3204 (N_3204,N_3123,N_3169);
xnor U3205 (N_3205,N_3091,N_3177);
xnor U3206 (N_3206,N_3132,N_3157);
or U3207 (N_3207,N_3049,N_3185);
nor U3208 (N_3208,N_3061,N_3022);
nor U3209 (N_3209,N_3001,N_3198);
nand U3210 (N_3210,N_3187,N_3087);
xor U3211 (N_3211,N_3019,N_3190);
xor U3212 (N_3212,N_3074,N_3057);
and U3213 (N_3213,N_3116,N_3018);
nand U3214 (N_3214,N_3103,N_3111);
and U3215 (N_3215,N_3081,N_3011);
nor U3216 (N_3216,N_3064,N_3170);
nor U3217 (N_3217,N_3141,N_3038);
nand U3218 (N_3218,N_3046,N_3129);
or U3219 (N_3219,N_3055,N_3072);
nand U3220 (N_3220,N_3094,N_3010);
nand U3221 (N_3221,N_3056,N_3135);
nand U3222 (N_3222,N_3133,N_3100);
nand U3223 (N_3223,N_3106,N_3075);
xnor U3224 (N_3224,N_3039,N_3164);
nor U3225 (N_3225,N_3083,N_3179);
nor U3226 (N_3226,N_3137,N_3052);
nor U3227 (N_3227,N_3070,N_3199);
xor U3228 (N_3228,N_3117,N_3098);
nand U3229 (N_3229,N_3006,N_3054);
nand U3230 (N_3230,N_3167,N_3145);
nor U3231 (N_3231,N_3027,N_3159);
and U3232 (N_3232,N_3093,N_3128);
xnor U3233 (N_3233,N_3127,N_3063);
or U3234 (N_3234,N_3175,N_3048);
or U3235 (N_3235,N_3042,N_3012);
and U3236 (N_3236,N_3172,N_3174);
and U3237 (N_3237,N_3035,N_3118);
xnor U3238 (N_3238,N_3050,N_3020);
nor U3239 (N_3239,N_3125,N_3180);
nor U3240 (N_3240,N_3078,N_3031);
nor U3241 (N_3241,N_3136,N_3108);
nor U3242 (N_3242,N_3080,N_3036);
xor U3243 (N_3243,N_3090,N_3126);
or U3244 (N_3244,N_3153,N_3120);
nand U3245 (N_3245,N_3021,N_3186);
and U3246 (N_3246,N_3069,N_3053);
xnor U3247 (N_3247,N_3017,N_3124);
and U3248 (N_3248,N_3008,N_3130);
nand U3249 (N_3249,N_3051,N_3076);
or U3250 (N_3250,N_3009,N_3033);
xor U3251 (N_3251,N_3171,N_3178);
or U3252 (N_3252,N_3121,N_3071);
or U3253 (N_3253,N_3029,N_3002);
xor U3254 (N_3254,N_3184,N_3032);
or U3255 (N_3255,N_3014,N_3088);
or U3256 (N_3256,N_3044,N_3195);
nand U3257 (N_3257,N_3059,N_3139);
and U3258 (N_3258,N_3034,N_3015);
or U3259 (N_3259,N_3077,N_3144);
and U3260 (N_3260,N_3194,N_3182);
nor U3261 (N_3261,N_3131,N_3168);
nand U3262 (N_3262,N_3007,N_3003);
xor U3263 (N_3263,N_3152,N_3066);
and U3264 (N_3264,N_3173,N_3183);
or U3265 (N_3265,N_3068,N_3028);
nor U3266 (N_3266,N_3016,N_3105);
xor U3267 (N_3267,N_3160,N_3150);
xor U3268 (N_3268,N_3096,N_3084);
or U3269 (N_3269,N_3045,N_3142);
or U3270 (N_3270,N_3065,N_3146);
or U3271 (N_3271,N_3013,N_3043);
nand U3272 (N_3272,N_3176,N_3148);
or U3273 (N_3273,N_3060,N_3119);
or U3274 (N_3274,N_3040,N_3151);
and U3275 (N_3275,N_3004,N_3102);
nand U3276 (N_3276,N_3082,N_3138);
nand U3277 (N_3277,N_3041,N_3101);
nor U3278 (N_3278,N_3113,N_3154);
or U3279 (N_3279,N_3099,N_3122);
or U3280 (N_3280,N_3110,N_3158);
or U3281 (N_3281,N_3155,N_3114);
or U3282 (N_3282,N_3097,N_3047);
nor U3283 (N_3283,N_3193,N_3085);
or U3284 (N_3284,N_3163,N_3161);
and U3285 (N_3285,N_3089,N_3107);
and U3286 (N_3286,N_3147,N_3115);
xnor U3287 (N_3287,N_3025,N_3079);
nor U3288 (N_3288,N_3134,N_3156);
or U3289 (N_3289,N_3005,N_3197);
or U3290 (N_3290,N_3026,N_3140);
and U3291 (N_3291,N_3192,N_3109);
xor U3292 (N_3292,N_3112,N_3086);
or U3293 (N_3293,N_3062,N_3196);
or U3294 (N_3294,N_3166,N_3037);
or U3295 (N_3295,N_3000,N_3188);
xnor U3296 (N_3296,N_3191,N_3165);
xor U3297 (N_3297,N_3149,N_3095);
xnor U3298 (N_3298,N_3181,N_3024);
nor U3299 (N_3299,N_3162,N_3092);
or U3300 (N_3300,N_3067,N_3111);
and U3301 (N_3301,N_3179,N_3100);
nor U3302 (N_3302,N_3163,N_3065);
nor U3303 (N_3303,N_3162,N_3007);
nor U3304 (N_3304,N_3195,N_3141);
nand U3305 (N_3305,N_3062,N_3013);
nor U3306 (N_3306,N_3142,N_3018);
and U3307 (N_3307,N_3037,N_3163);
nor U3308 (N_3308,N_3025,N_3004);
nand U3309 (N_3309,N_3160,N_3020);
nand U3310 (N_3310,N_3094,N_3001);
xor U3311 (N_3311,N_3126,N_3097);
xor U3312 (N_3312,N_3049,N_3168);
nand U3313 (N_3313,N_3023,N_3065);
or U3314 (N_3314,N_3176,N_3172);
or U3315 (N_3315,N_3025,N_3061);
xnor U3316 (N_3316,N_3168,N_3053);
and U3317 (N_3317,N_3054,N_3043);
nor U3318 (N_3318,N_3169,N_3146);
or U3319 (N_3319,N_3192,N_3024);
nand U3320 (N_3320,N_3119,N_3061);
nor U3321 (N_3321,N_3159,N_3061);
xor U3322 (N_3322,N_3144,N_3081);
nor U3323 (N_3323,N_3181,N_3154);
or U3324 (N_3324,N_3034,N_3178);
xnor U3325 (N_3325,N_3158,N_3185);
xnor U3326 (N_3326,N_3114,N_3173);
and U3327 (N_3327,N_3155,N_3006);
nor U3328 (N_3328,N_3193,N_3121);
nand U3329 (N_3329,N_3151,N_3199);
or U3330 (N_3330,N_3110,N_3124);
or U3331 (N_3331,N_3182,N_3165);
xnor U3332 (N_3332,N_3086,N_3011);
and U3333 (N_3333,N_3048,N_3017);
nand U3334 (N_3334,N_3056,N_3052);
nand U3335 (N_3335,N_3081,N_3016);
nand U3336 (N_3336,N_3184,N_3049);
nand U3337 (N_3337,N_3152,N_3061);
or U3338 (N_3338,N_3074,N_3149);
nand U3339 (N_3339,N_3080,N_3086);
or U3340 (N_3340,N_3115,N_3065);
nor U3341 (N_3341,N_3193,N_3151);
and U3342 (N_3342,N_3111,N_3119);
nor U3343 (N_3343,N_3133,N_3093);
and U3344 (N_3344,N_3173,N_3108);
nor U3345 (N_3345,N_3070,N_3121);
and U3346 (N_3346,N_3046,N_3191);
nand U3347 (N_3347,N_3075,N_3101);
xor U3348 (N_3348,N_3029,N_3009);
and U3349 (N_3349,N_3175,N_3140);
nor U3350 (N_3350,N_3097,N_3125);
nand U3351 (N_3351,N_3101,N_3028);
xor U3352 (N_3352,N_3113,N_3055);
nand U3353 (N_3353,N_3158,N_3171);
nor U3354 (N_3354,N_3123,N_3097);
xor U3355 (N_3355,N_3087,N_3018);
and U3356 (N_3356,N_3093,N_3087);
nand U3357 (N_3357,N_3072,N_3117);
and U3358 (N_3358,N_3140,N_3168);
or U3359 (N_3359,N_3120,N_3049);
and U3360 (N_3360,N_3011,N_3043);
xnor U3361 (N_3361,N_3130,N_3015);
xnor U3362 (N_3362,N_3140,N_3042);
xnor U3363 (N_3363,N_3014,N_3150);
nor U3364 (N_3364,N_3162,N_3141);
xor U3365 (N_3365,N_3002,N_3077);
xnor U3366 (N_3366,N_3094,N_3130);
nor U3367 (N_3367,N_3117,N_3108);
xor U3368 (N_3368,N_3101,N_3163);
or U3369 (N_3369,N_3190,N_3032);
and U3370 (N_3370,N_3159,N_3111);
and U3371 (N_3371,N_3067,N_3158);
and U3372 (N_3372,N_3059,N_3199);
and U3373 (N_3373,N_3123,N_3027);
nor U3374 (N_3374,N_3094,N_3181);
xor U3375 (N_3375,N_3041,N_3075);
nand U3376 (N_3376,N_3178,N_3001);
nor U3377 (N_3377,N_3117,N_3080);
nor U3378 (N_3378,N_3146,N_3194);
xor U3379 (N_3379,N_3110,N_3041);
and U3380 (N_3380,N_3186,N_3092);
nand U3381 (N_3381,N_3082,N_3164);
nor U3382 (N_3382,N_3001,N_3040);
and U3383 (N_3383,N_3114,N_3139);
nor U3384 (N_3384,N_3048,N_3057);
xnor U3385 (N_3385,N_3013,N_3128);
and U3386 (N_3386,N_3086,N_3107);
or U3387 (N_3387,N_3065,N_3136);
xnor U3388 (N_3388,N_3141,N_3116);
or U3389 (N_3389,N_3116,N_3147);
or U3390 (N_3390,N_3127,N_3029);
nand U3391 (N_3391,N_3011,N_3082);
or U3392 (N_3392,N_3085,N_3045);
nand U3393 (N_3393,N_3089,N_3152);
and U3394 (N_3394,N_3105,N_3029);
xnor U3395 (N_3395,N_3176,N_3190);
and U3396 (N_3396,N_3013,N_3135);
or U3397 (N_3397,N_3062,N_3092);
nor U3398 (N_3398,N_3195,N_3086);
or U3399 (N_3399,N_3015,N_3082);
and U3400 (N_3400,N_3236,N_3309);
nand U3401 (N_3401,N_3316,N_3379);
xnor U3402 (N_3402,N_3267,N_3311);
xnor U3403 (N_3403,N_3288,N_3330);
nor U3404 (N_3404,N_3230,N_3315);
xnor U3405 (N_3405,N_3225,N_3229);
and U3406 (N_3406,N_3354,N_3301);
nor U3407 (N_3407,N_3342,N_3264);
xor U3408 (N_3408,N_3265,N_3345);
or U3409 (N_3409,N_3278,N_3241);
nor U3410 (N_3410,N_3346,N_3216);
xnor U3411 (N_3411,N_3224,N_3333);
xor U3412 (N_3412,N_3392,N_3339);
xnor U3413 (N_3413,N_3329,N_3266);
nor U3414 (N_3414,N_3271,N_3323);
and U3415 (N_3415,N_3300,N_3310);
and U3416 (N_3416,N_3356,N_3303);
xor U3417 (N_3417,N_3220,N_3270);
nor U3418 (N_3418,N_3343,N_3357);
nor U3419 (N_3419,N_3371,N_3255);
xnor U3420 (N_3420,N_3332,N_3273);
nor U3421 (N_3421,N_3295,N_3243);
and U3422 (N_3422,N_3231,N_3215);
nor U3423 (N_3423,N_3212,N_3284);
and U3424 (N_3424,N_3203,N_3279);
nor U3425 (N_3425,N_3360,N_3353);
and U3426 (N_3426,N_3268,N_3237);
nor U3427 (N_3427,N_3285,N_3364);
nor U3428 (N_3428,N_3217,N_3373);
and U3429 (N_3429,N_3256,N_3221);
xnor U3430 (N_3430,N_3366,N_3319);
nor U3431 (N_3431,N_3369,N_3349);
nor U3432 (N_3432,N_3355,N_3361);
or U3433 (N_3433,N_3351,N_3209);
xor U3434 (N_3434,N_3308,N_3235);
and U3435 (N_3435,N_3290,N_3283);
nand U3436 (N_3436,N_3200,N_3375);
nand U3437 (N_3437,N_3210,N_3334);
or U3438 (N_3438,N_3254,N_3289);
nand U3439 (N_3439,N_3382,N_3249);
nor U3440 (N_3440,N_3391,N_3370);
nor U3441 (N_3441,N_3281,N_3340);
or U3442 (N_3442,N_3247,N_3377);
nand U3443 (N_3443,N_3307,N_3350);
xor U3444 (N_3444,N_3372,N_3286);
or U3445 (N_3445,N_3344,N_3321);
nor U3446 (N_3446,N_3205,N_3302);
and U3447 (N_3447,N_3223,N_3282);
xor U3448 (N_3448,N_3232,N_3326);
xor U3449 (N_3449,N_3261,N_3386);
or U3450 (N_3450,N_3275,N_3367);
xnor U3451 (N_3451,N_3226,N_3245);
nor U3452 (N_3452,N_3234,N_3222);
and U3453 (N_3453,N_3393,N_3228);
or U3454 (N_3454,N_3335,N_3395);
or U3455 (N_3455,N_3240,N_3242);
nand U3456 (N_3456,N_3338,N_3219);
or U3457 (N_3457,N_3257,N_3263);
and U3458 (N_3458,N_3274,N_3297);
xnor U3459 (N_3459,N_3298,N_3204);
xnor U3460 (N_3460,N_3314,N_3347);
xnor U3461 (N_3461,N_3280,N_3322);
nand U3462 (N_3462,N_3380,N_3260);
xnor U3463 (N_3463,N_3238,N_3306);
nor U3464 (N_3464,N_3250,N_3244);
or U3465 (N_3465,N_3218,N_3269);
or U3466 (N_3466,N_3248,N_3388);
xor U3467 (N_3467,N_3362,N_3385);
nand U3468 (N_3468,N_3318,N_3276);
and U3469 (N_3469,N_3398,N_3201);
and U3470 (N_3470,N_3251,N_3352);
or U3471 (N_3471,N_3317,N_3384);
nor U3472 (N_3472,N_3294,N_3258);
xnor U3473 (N_3473,N_3259,N_3397);
nand U3474 (N_3474,N_3213,N_3239);
nor U3475 (N_3475,N_3394,N_3252);
nand U3476 (N_3476,N_3313,N_3292);
and U3477 (N_3477,N_3320,N_3396);
or U3478 (N_3478,N_3387,N_3272);
or U3479 (N_3479,N_3233,N_3305);
and U3480 (N_3480,N_3336,N_3358);
xnor U3481 (N_3481,N_3325,N_3246);
and U3482 (N_3482,N_3214,N_3363);
nor U3483 (N_3483,N_3381,N_3324);
xor U3484 (N_3484,N_3207,N_3348);
xor U3485 (N_3485,N_3389,N_3299);
nand U3486 (N_3486,N_3390,N_3331);
xnor U3487 (N_3487,N_3227,N_3378);
or U3488 (N_3488,N_3359,N_3312);
and U3489 (N_3489,N_3277,N_3337);
nand U3490 (N_3490,N_3211,N_3368);
or U3491 (N_3491,N_3262,N_3327);
nor U3492 (N_3492,N_3365,N_3328);
and U3493 (N_3493,N_3399,N_3341);
xnor U3494 (N_3494,N_3202,N_3296);
and U3495 (N_3495,N_3293,N_3206);
xor U3496 (N_3496,N_3291,N_3304);
or U3497 (N_3497,N_3383,N_3374);
nand U3498 (N_3498,N_3253,N_3376);
xnor U3499 (N_3499,N_3287,N_3208);
or U3500 (N_3500,N_3333,N_3295);
or U3501 (N_3501,N_3248,N_3335);
xnor U3502 (N_3502,N_3272,N_3315);
and U3503 (N_3503,N_3220,N_3225);
or U3504 (N_3504,N_3310,N_3397);
or U3505 (N_3505,N_3327,N_3345);
nand U3506 (N_3506,N_3304,N_3396);
or U3507 (N_3507,N_3210,N_3320);
or U3508 (N_3508,N_3304,N_3313);
xor U3509 (N_3509,N_3282,N_3306);
and U3510 (N_3510,N_3258,N_3228);
nand U3511 (N_3511,N_3396,N_3256);
and U3512 (N_3512,N_3286,N_3274);
xnor U3513 (N_3513,N_3298,N_3319);
or U3514 (N_3514,N_3283,N_3243);
and U3515 (N_3515,N_3219,N_3343);
xnor U3516 (N_3516,N_3281,N_3295);
nor U3517 (N_3517,N_3256,N_3212);
nand U3518 (N_3518,N_3340,N_3223);
xnor U3519 (N_3519,N_3388,N_3377);
nor U3520 (N_3520,N_3213,N_3222);
and U3521 (N_3521,N_3350,N_3269);
and U3522 (N_3522,N_3300,N_3392);
nand U3523 (N_3523,N_3328,N_3299);
nand U3524 (N_3524,N_3343,N_3252);
xnor U3525 (N_3525,N_3381,N_3357);
nand U3526 (N_3526,N_3367,N_3327);
or U3527 (N_3527,N_3329,N_3214);
xor U3528 (N_3528,N_3366,N_3380);
xor U3529 (N_3529,N_3202,N_3252);
or U3530 (N_3530,N_3307,N_3215);
nand U3531 (N_3531,N_3218,N_3315);
nand U3532 (N_3532,N_3379,N_3280);
nand U3533 (N_3533,N_3376,N_3356);
nand U3534 (N_3534,N_3313,N_3381);
xor U3535 (N_3535,N_3202,N_3312);
xor U3536 (N_3536,N_3371,N_3385);
xnor U3537 (N_3537,N_3392,N_3275);
nor U3538 (N_3538,N_3296,N_3264);
and U3539 (N_3539,N_3213,N_3372);
nand U3540 (N_3540,N_3237,N_3363);
or U3541 (N_3541,N_3259,N_3294);
and U3542 (N_3542,N_3208,N_3351);
and U3543 (N_3543,N_3363,N_3239);
or U3544 (N_3544,N_3205,N_3358);
and U3545 (N_3545,N_3316,N_3339);
nand U3546 (N_3546,N_3255,N_3383);
nand U3547 (N_3547,N_3338,N_3308);
or U3548 (N_3548,N_3264,N_3206);
and U3549 (N_3549,N_3227,N_3226);
and U3550 (N_3550,N_3319,N_3281);
nand U3551 (N_3551,N_3214,N_3341);
and U3552 (N_3552,N_3283,N_3205);
xnor U3553 (N_3553,N_3229,N_3266);
nor U3554 (N_3554,N_3213,N_3282);
xnor U3555 (N_3555,N_3231,N_3201);
xor U3556 (N_3556,N_3211,N_3255);
nand U3557 (N_3557,N_3347,N_3350);
nand U3558 (N_3558,N_3345,N_3374);
or U3559 (N_3559,N_3218,N_3329);
xor U3560 (N_3560,N_3318,N_3236);
xor U3561 (N_3561,N_3204,N_3335);
and U3562 (N_3562,N_3353,N_3300);
nor U3563 (N_3563,N_3364,N_3263);
and U3564 (N_3564,N_3237,N_3311);
and U3565 (N_3565,N_3343,N_3213);
xnor U3566 (N_3566,N_3397,N_3264);
nand U3567 (N_3567,N_3362,N_3228);
nor U3568 (N_3568,N_3212,N_3375);
nor U3569 (N_3569,N_3291,N_3337);
nand U3570 (N_3570,N_3205,N_3316);
and U3571 (N_3571,N_3353,N_3376);
nand U3572 (N_3572,N_3235,N_3283);
nand U3573 (N_3573,N_3363,N_3299);
or U3574 (N_3574,N_3259,N_3293);
and U3575 (N_3575,N_3327,N_3271);
and U3576 (N_3576,N_3356,N_3375);
xor U3577 (N_3577,N_3329,N_3318);
and U3578 (N_3578,N_3252,N_3372);
nand U3579 (N_3579,N_3280,N_3302);
xor U3580 (N_3580,N_3269,N_3292);
xnor U3581 (N_3581,N_3238,N_3285);
and U3582 (N_3582,N_3379,N_3374);
and U3583 (N_3583,N_3263,N_3324);
nand U3584 (N_3584,N_3212,N_3391);
or U3585 (N_3585,N_3210,N_3200);
xor U3586 (N_3586,N_3290,N_3256);
xnor U3587 (N_3587,N_3310,N_3305);
or U3588 (N_3588,N_3308,N_3342);
and U3589 (N_3589,N_3352,N_3214);
and U3590 (N_3590,N_3308,N_3254);
or U3591 (N_3591,N_3275,N_3271);
nor U3592 (N_3592,N_3219,N_3350);
nor U3593 (N_3593,N_3290,N_3226);
nor U3594 (N_3594,N_3310,N_3226);
and U3595 (N_3595,N_3350,N_3238);
xnor U3596 (N_3596,N_3331,N_3397);
nand U3597 (N_3597,N_3398,N_3386);
xor U3598 (N_3598,N_3310,N_3337);
and U3599 (N_3599,N_3235,N_3342);
and U3600 (N_3600,N_3570,N_3537);
or U3601 (N_3601,N_3527,N_3517);
or U3602 (N_3602,N_3405,N_3562);
nand U3603 (N_3603,N_3451,N_3524);
nor U3604 (N_3604,N_3404,N_3409);
and U3605 (N_3605,N_3473,N_3490);
nand U3606 (N_3606,N_3528,N_3478);
xnor U3607 (N_3607,N_3436,N_3550);
xnor U3608 (N_3608,N_3419,N_3509);
or U3609 (N_3609,N_3505,N_3544);
xnor U3610 (N_3610,N_3593,N_3487);
nand U3611 (N_3611,N_3424,N_3568);
nand U3612 (N_3612,N_3449,N_3591);
xor U3613 (N_3613,N_3406,N_3472);
and U3614 (N_3614,N_3563,N_3471);
nor U3615 (N_3615,N_3440,N_3486);
nor U3616 (N_3616,N_3523,N_3476);
xor U3617 (N_3617,N_3501,N_3585);
xor U3618 (N_3618,N_3598,N_3447);
nand U3619 (N_3619,N_3462,N_3431);
or U3620 (N_3620,N_3565,N_3477);
nor U3621 (N_3621,N_3519,N_3470);
xnor U3622 (N_3622,N_3457,N_3442);
and U3623 (N_3623,N_3512,N_3594);
nand U3624 (N_3624,N_3589,N_3535);
nor U3625 (N_3625,N_3588,N_3574);
xor U3626 (N_3626,N_3410,N_3450);
or U3627 (N_3627,N_3547,N_3480);
or U3628 (N_3628,N_3458,N_3564);
and U3629 (N_3629,N_3561,N_3586);
and U3630 (N_3630,N_3467,N_3448);
nand U3631 (N_3631,N_3520,N_3599);
or U3632 (N_3632,N_3533,N_3445);
xor U3633 (N_3633,N_3584,N_3554);
and U3634 (N_3634,N_3592,N_3546);
or U3635 (N_3635,N_3545,N_3485);
or U3636 (N_3636,N_3510,N_3474);
xor U3637 (N_3637,N_3414,N_3529);
nor U3638 (N_3638,N_3402,N_3465);
and U3639 (N_3639,N_3499,N_3461);
nor U3640 (N_3640,N_3515,N_3525);
and U3641 (N_3641,N_3541,N_3559);
xnor U3642 (N_3642,N_3400,N_3425);
and U3643 (N_3643,N_3569,N_3494);
and U3644 (N_3644,N_3464,N_3557);
nor U3645 (N_3645,N_3463,N_3423);
or U3646 (N_3646,N_3430,N_3567);
or U3647 (N_3647,N_3514,N_3583);
and U3648 (N_3648,N_3426,N_3548);
or U3649 (N_3649,N_3553,N_3435);
nor U3650 (N_3650,N_3444,N_3551);
xor U3651 (N_3651,N_3433,N_3502);
and U3652 (N_3652,N_3500,N_3453);
xor U3653 (N_3653,N_3498,N_3403);
or U3654 (N_3654,N_3456,N_3516);
nor U3655 (N_3655,N_3595,N_3455);
nor U3656 (N_3656,N_3488,N_3578);
nor U3657 (N_3657,N_3556,N_3532);
nor U3658 (N_3658,N_3504,N_3566);
nand U3659 (N_3659,N_3540,N_3495);
or U3660 (N_3660,N_3534,N_3596);
and U3661 (N_3661,N_3587,N_3417);
or U3662 (N_3662,N_3543,N_3446);
and U3663 (N_3663,N_3411,N_3513);
and U3664 (N_3664,N_3503,N_3580);
nor U3665 (N_3665,N_3497,N_3413);
nor U3666 (N_3666,N_3590,N_3427);
and U3667 (N_3667,N_3576,N_3522);
nand U3668 (N_3668,N_3416,N_3597);
and U3669 (N_3669,N_3518,N_3536);
nand U3670 (N_3670,N_3482,N_3454);
and U3671 (N_3671,N_3407,N_3489);
nand U3672 (N_3672,N_3466,N_3481);
or U3673 (N_3673,N_3507,N_3475);
or U3674 (N_3674,N_3452,N_3558);
or U3675 (N_3675,N_3577,N_3530);
and U3676 (N_3676,N_3496,N_3582);
and U3677 (N_3677,N_3542,N_3421);
nor U3678 (N_3678,N_3437,N_3438);
nand U3679 (N_3679,N_3538,N_3491);
xnor U3680 (N_3680,N_3555,N_3415);
xor U3681 (N_3681,N_3460,N_3401);
nand U3682 (N_3682,N_3539,N_3573);
and U3683 (N_3683,N_3429,N_3459);
or U3684 (N_3684,N_3408,N_3484);
nand U3685 (N_3685,N_3572,N_3434);
xnor U3686 (N_3686,N_3508,N_3420);
nor U3687 (N_3687,N_3441,N_3412);
and U3688 (N_3688,N_3531,N_3571);
xor U3689 (N_3689,N_3483,N_3521);
xnor U3690 (N_3690,N_3581,N_3439);
nand U3691 (N_3691,N_3493,N_3443);
xor U3692 (N_3692,N_3526,N_3418);
and U3693 (N_3693,N_3468,N_3506);
nor U3694 (N_3694,N_3479,N_3575);
and U3695 (N_3695,N_3560,N_3432);
nor U3696 (N_3696,N_3428,N_3549);
nor U3697 (N_3697,N_3492,N_3552);
nand U3698 (N_3698,N_3469,N_3422);
nand U3699 (N_3699,N_3579,N_3511);
and U3700 (N_3700,N_3487,N_3521);
or U3701 (N_3701,N_3426,N_3465);
xor U3702 (N_3702,N_3420,N_3586);
or U3703 (N_3703,N_3461,N_3584);
or U3704 (N_3704,N_3405,N_3507);
nor U3705 (N_3705,N_3479,N_3459);
xnor U3706 (N_3706,N_3491,N_3422);
and U3707 (N_3707,N_3477,N_3529);
nand U3708 (N_3708,N_3560,N_3418);
and U3709 (N_3709,N_3424,N_3593);
nor U3710 (N_3710,N_3400,N_3488);
nand U3711 (N_3711,N_3586,N_3558);
or U3712 (N_3712,N_3418,N_3516);
nand U3713 (N_3713,N_3552,N_3420);
or U3714 (N_3714,N_3522,N_3570);
or U3715 (N_3715,N_3577,N_3413);
and U3716 (N_3716,N_3512,N_3535);
or U3717 (N_3717,N_3569,N_3547);
and U3718 (N_3718,N_3550,N_3568);
nand U3719 (N_3719,N_3475,N_3540);
nor U3720 (N_3720,N_3541,N_3588);
and U3721 (N_3721,N_3486,N_3540);
xnor U3722 (N_3722,N_3406,N_3422);
xor U3723 (N_3723,N_3413,N_3430);
xor U3724 (N_3724,N_3505,N_3403);
nand U3725 (N_3725,N_3541,N_3411);
nor U3726 (N_3726,N_3563,N_3546);
nand U3727 (N_3727,N_3598,N_3539);
xnor U3728 (N_3728,N_3555,N_3462);
or U3729 (N_3729,N_3549,N_3425);
and U3730 (N_3730,N_3407,N_3580);
nor U3731 (N_3731,N_3558,N_3546);
nor U3732 (N_3732,N_3438,N_3448);
xnor U3733 (N_3733,N_3514,N_3588);
and U3734 (N_3734,N_3595,N_3536);
xor U3735 (N_3735,N_3556,N_3495);
and U3736 (N_3736,N_3521,N_3488);
or U3737 (N_3737,N_3419,N_3411);
nand U3738 (N_3738,N_3514,N_3425);
xnor U3739 (N_3739,N_3448,N_3552);
and U3740 (N_3740,N_3468,N_3492);
or U3741 (N_3741,N_3479,N_3559);
nand U3742 (N_3742,N_3400,N_3577);
xor U3743 (N_3743,N_3524,N_3543);
and U3744 (N_3744,N_3500,N_3465);
or U3745 (N_3745,N_3406,N_3514);
and U3746 (N_3746,N_3588,N_3486);
nor U3747 (N_3747,N_3539,N_3564);
and U3748 (N_3748,N_3401,N_3532);
or U3749 (N_3749,N_3498,N_3470);
nor U3750 (N_3750,N_3527,N_3407);
or U3751 (N_3751,N_3466,N_3474);
nand U3752 (N_3752,N_3426,N_3417);
nor U3753 (N_3753,N_3407,N_3425);
nor U3754 (N_3754,N_3478,N_3561);
xnor U3755 (N_3755,N_3489,N_3554);
or U3756 (N_3756,N_3429,N_3458);
or U3757 (N_3757,N_3429,N_3540);
or U3758 (N_3758,N_3562,N_3481);
nand U3759 (N_3759,N_3573,N_3470);
nor U3760 (N_3760,N_3534,N_3526);
xor U3761 (N_3761,N_3552,N_3501);
xor U3762 (N_3762,N_3424,N_3483);
nor U3763 (N_3763,N_3478,N_3557);
nand U3764 (N_3764,N_3572,N_3403);
nand U3765 (N_3765,N_3515,N_3522);
nand U3766 (N_3766,N_3420,N_3542);
nor U3767 (N_3767,N_3437,N_3522);
nand U3768 (N_3768,N_3518,N_3482);
nand U3769 (N_3769,N_3546,N_3506);
and U3770 (N_3770,N_3432,N_3536);
nor U3771 (N_3771,N_3496,N_3498);
and U3772 (N_3772,N_3576,N_3425);
nand U3773 (N_3773,N_3444,N_3574);
and U3774 (N_3774,N_3409,N_3539);
nand U3775 (N_3775,N_3441,N_3531);
nand U3776 (N_3776,N_3556,N_3509);
or U3777 (N_3777,N_3594,N_3489);
or U3778 (N_3778,N_3456,N_3410);
nor U3779 (N_3779,N_3485,N_3552);
nor U3780 (N_3780,N_3592,N_3430);
nor U3781 (N_3781,N_3586,N_3481);
or U3782 (N_3782,N_3465,N_3534);
nor U3783 (N_3783,N_3578,N_3483);
nor U3784 (N_3784,N_3421,N_3570);
nand U3785 (N_3785,N_3518,N_3545);
and U3786 (N_3786,N_3565,N_3407);
or U3787 (N_3787,N_3587,N_3542);
or U3788 (N_3788,N_3590,N_3448);
or U3789 (N_3789,N_3525,N_3558);
or U3790 (N_3790,N_3484,N_3533);
xor U3791 (N_3791,N_3566,N_3449);
and U3792 (N_3792,N_3403,N_3507);
nand U3793 (N_3793,N_3525,N_3431);
or U3794 (N_3794,N_3509,N_3482);
xor U3795 (N_3795,N_3427,N_3567);
or U3796 (N_3796,N_3552,N_3577);
nand U3797 (N_3797,N_3480,N_3478);
nand U3798 (N_3798,N_3496,N_3492);
and U3799 (N_3799,N_3575,N_3503);
xnor U3800 (N_3800,N_3799,N_3743);
or U3801 (N_3801,N_3602,N_3653);
nor U3802 (N_3802,N_3721,N_3619);
or U3803 (N_3803,N_3744,N_3682);
nand U3804 (N_3804,N_3707,N_3715);
or U3805 (N_3805,N_3639,N_3648);
xnor U3806 (N_3806,N_3696,N_3733);
nand U3807 (N_3807,N_3764,N_3643);
nand U3808 (N_3808,N_3650,N_3681);
nand U3809 (N_3809,N_3669,N_3732);
nor U3810 (N_3810,N_3644,N_3797);
nand U3811 (N_3811,N_3726,N_3772);
xor U3812 (N_3812,N_3690,N_3734);
nand U3813 (N_3813,N_3674,N_3796);
nand U3814 (N_3814,N_3634,N_3714);
and U3815 (N_3815,N_3774,N_3622);
and U3816 (N_3816,N_3710,N_3782);
and U3817 (N_3817,N_3637,N_3706);
xnor U3818 (N_3818,N_3680,N_3638);
or U3819 (N_3819,N_3646,N_3778);
xnor U3820 (N_3820,N_3686,N_3630);
nor U3821 (N_3821,N_3668,N_3738);
xnor U3822 (N_3822,N_3740,N_3728);
nand U3823 (N_3823,N_3632,N_3725);
nand U3824 (N_3824,N_3664,N_3768);
and U3825 (N_3825,N_3699,N_3709);
and U3826 (N_3826,N_3792,N_3758);
nor U3827 (N_3827,N_3687,N_3611);
nand U3828 (N_3828,N_3751,N_3749);
nand U3829 (N_3829,N_3684,N_3755);
xnor U3830 (N_3830,N_3702,N_3784);
nand U3831 (N_3831,N_3767,N_3691);
and U3832 (N_3832,N_3703,N_3727);
xor U3833 (N_3833,N_3761,N_3787);
nand U3834 (N_3834,N_3775,N_3623);
nor U3835 (N_3835,N_3616,N_3736);
or U3836 (N_3836,N_3610,N_3737);
xor U3837 (N_3837,N_3645,N_3741);
nor U3838 (N_3838,N_3695,N_3683);
and U3839 (N_3839,N_3789,N_3621);
xnor U3840 (N_3840,N_3604,N_3601);
nand U3841 (N_3841,N_3723,N_3625);
or U3842 (N_3842,N_3730,N_3688);
and U3843 (N_3843,N_3700,N_3626);
or U3844 (N_3844,N_3711,N_3641);
and U3845 (N_3845,N_3786,N_3780);
xnor U3846 (N_3846,N_3662,N_3746);
nor U3847 (N_3847,N_3658,N_3649);
xnor U3848 (N_3848,N_3615,N_3661);
nor U3849 (N_3849,N_3689,N_3605);
nor U3850 (N_3850,N_3798,N_3794);
or U3851 (N_3851,N_3779,N_3757);
and U3852 (N_3852,N_3633,N_3765);
nor U3853 (N_3853,N_3667,N_3678);
nand U3854 (N_3854,N_3716,N_3790);
nand U3855 (N_3855,N_3793,N_3675);
nand U3856 (N_3856,N_3612,N_3624);
or U3857 (N_3857,N_3693,N_3742);
xnor U3858 (N_3858,N_3747,N_3762);
nor U3859 (N_3859,N_3719,N_3676);
or U3860 (N_3860,N_3748,N_3657);
and U3861 (N_3861,N_3705,N_3607);
nand U3862 (N_3862,N_3670,N_3663);
or U3863 (N_3863,N_3692,N_3651);
nand U3864 (N_3864,N_3629,N_3773);
nand U3865 (N_3865,N_3759,N_3771);
or U3866 (N_3866,N_3631,N_3752);
or U3867 (N_3867,N_3753,N_3769);
and U3868 (N_3868,N_3788,N_3614);
or U3869 (N_3869,N_3750,N_3756);
xor U3870 (N_3870,N_3739,N_3636);
and U3871 (N_3871,N_3642,N_3729);
xor U3872 (N_3872,N_3718,N_3720);
nand U3873 (N_3873,N_3701,N_3685);
xnor U3874 (N_3874,N_3666,N_3694);
nand U3875 (N_3875,N_3618,N_3704);
xor U3876 (N_3876,N_3712,N_3665);
nor U3877 (N_3877,N_3655,N_3708);
or U3878 (N_3878,N_3766,N_3677);
and U3879 (N_3879,N_3785,N_3673);
nor U3880 (N_3880,N_3628,N_3717);
or U3881 (N_3881,N_3652,N_3640);
or U3882 (N_3882,N_3697,N_3617);
nand U3883 (N_3883,N_3776,N_3647);
xor U3884 (N_3884,N_3795,N_3613);
xnor U3885 (N_3885,N_3777,N_3783);
nand U3886 (N_3886,N_3724,N_3656);
and U3887 (N_3887,N_3671,N_3754);
nand U3888 (N_3888,N_3698,N_3620);
xnor U3889 (N_3889,N_3603,N_3672);
nand U3890 (N_3890,N_3659,N_3609);
nand U3891 (N_3891,N_3731,N_3713);
or U3892 (N_3892,N_3770,N_3760);
nand U3893 (N_3893,N_3608,N_3635);
nand U3894 (N_3894,N_3627,N_3654);
or U3895 (N_3895,N_3679,N_3722);
nor U3896 (N_3896,N_3600,N_3781);
nand U3897 (N_3897,N_3763,N_3791);
xnor U3898 (N_3898,N_3660,N_3745);
xnor U3899 (N_3899,N_3606,N_3735);
nor U3900 (N_3900,N_3604,N_3663);
xor U3901 (N_3901,N_3767,N_3686);
xor U3902 (N_3902,N_3771,N_3754);
and U3903 (N_3903,N_3784,N_3671);
xor U3904 (N_3904,N_3766,N_3784);
nand U3905 (N_3905,N_3797,N_3681);
and U3906 (N_3906,N_3675,N_3626);
nor U3907 (N_3907,N_3638,N_3742);
nor U3908 (N_3908,N_3785,N_3795);
xnor U3909 (N_3909,N_3683,N_3765);
xnor U3910 (N_3910,N_3703,N_3772);
and U3911 (N_3911,N_3726,N_3769);
xnor U3912 (N_3912,N_3750,N_3650);
or U3913 (N_3913,N_3642,N_3625);
or U3914 (N_3914,N_3602,N_3677);
xor U3915 (N_3915,N_3677,N_3701);
or U3916 (N_3916,N_3673,N_3747);
nand U3917 (N_3917,N_3672,N_3749);
nor U3918 (N_3918,N_3646,N_3787);
or U3919 (N_3919,N_3626,N_3756);
and U3920 (N_3920,N_3792,N_3786);
or U3921 (N_3921,N_3709,N_3765);
nand U3922 (N_3922,N_3687,N_3683);
and U3923 (N_3923,N_3668,N_3672);
nor U3924 (N_3924,N_3718,N_3791);
xnor U3925 (N_3925,N_3670,N_3736);
and U3926 (N_3926,N_3724,N_3683);
and U3927 (N_3927,N_3604,N_3798);
or U3928 (N_3928,N_3622,N_3706);
and U3929 (N_3929,N_3773,N_3688);
or U3930 (N_3930,N_3797,N_3732);
and U3931 (N_3931,N_3709,N_3681);
nor U3932 (N_3932,N_3605,N_3698);
and U3933 (N_3933,N_3699,N_3719);
nand U3934 (N_3934,N_3642,N_3780);
nor U3935 (N_3935,N_3712,N_3659);
xnor U3936 (N_3936,N_3713,N_3615);
or U3937 (N_3937,N_3631,N_3606);
nand U3938 (N_3938,N_3659,N_3787);
nand U3939 (N_3939,N_3695,N_3658);
or U3940 (N_3940,N_3719,N_3753);
and U3941 (N_3941,N_3689,N_3727);
or U3942 (N_3942,N_3761,N_3650);
and U3943 (N_3943,N_3723,N_3654);
and U3944 (N_3944,N_3648,N_3765);
nor U3945 (N_3945,N_3771,N_3715);
nand U3946 (N_3946,N_3792,N_3771);
and U3947 (N_3947,N_3665,N_3649);
xnor U3948 (N_3948,N_3757,N_3700);
and U3949 (N_3949,N_3681,N_3745);
nand U3950 (N_3950,N_3664,N_3790);
or U3951 (N_3951,N_3784,N_3634);
or U3952 (N_3952,N_3632,N_3652);
nand U3953 (N_3953,N_3685,N_3737);
xor U3954 (N_3954,N_3691,N_3686);
nor U3955 (N_3955,N_3713,N_3673);
nand U3956 (N_3956,N_3651,N_3610);
or U3957 (N_3957,N_3604,N_3783);
and U3958 (N_3958,N_3752,N_3647);
or U3959 (N_3959,N_3729,N_3686);
xor U3960 (N_3960,N_3761,N_3794);
and U3961 (N_3961,N_3606,N_3747);
nand U3962 (N_3962,N_3635,N_3605);
nor U3963 (N_3963,N_3692,N_3602);
or U3964 (N_3964,N_3633,N_3720);
and U3965 (N_3965,N_3792,N_3670);
or U3966 (N_3966,N_3655,N_3782);
or U3967 (N_3967,N_3620,N_3611);
and U3968 (N_3968,N_3606,N_3662);
nor U3969 (N_3969,N_3609,N_3605);
or U3970 (N_3970,N_3779,N_3778);
xnor U3971 (N_3971,N_3710,N_3625);
nand U3972 (N_3972,N_3786,N_3622);
nor U3973 (N_3973,N_3624,N_3721);
or U3974 (N_3974,N_3784,N_3619);
xor U3975 (N_3975,N_3627,N_3613);
nor U3976 (N_3976,N_3689,N_3602);
and U3977 (N_3977,N_3645,N_3694);
nor U3978 (N_3978,N_3795,N_3760);
nand U3979 (N_3979,N_3752,N_3636);
xnor U3980 (N_3980,N_3677,N_3649);
and U3981 (N_3981,N_3765,N_3647);
or U3982 (N_3982,N_3738,N_3690);
xnor U3983 (N_3983,N_3747,N_3718);
nor U3984 (N_3984,N_3664,N_3687);
xor U3985 (N_3985,N_3720,N_3644);
or U3986 (N_3986,N_3704,N_3722);
xnor U3987 (N_3987,N_3605,N_3740);
or U3988 (N_3988,N_3759,N_3668);
xor U3989 (N_3989,N_3685,N_3712);
or U3990 (N_3990,N_3663,N_3690);
nand U3991 (N_3991,N_3644,N_3740);
and U3992 (N_3992,N_3717,N_3764);
nor U3993 (N_3993,N_3715,N_3712);
and U3994 (N_3994,N_3699,N_3763);
xnor U3995 (N_3995,N_3779,N_3732);
xor U3996 (N_3996,N_3726,N_3781);
nand U3997 (N_3997,N_3664,N_3624);
nor U3998 (N_3998,N_3716,N_3611);
or U3999 (N_3999,N_3680,N_3652);
nand U4000 (N_4000,N_3961,N_3954);
or U4001 (N_4001,N_3975,N_3992);
nand U4002 (N_4002,N_3850,N_3913);
nand U4003 (N_4003,N_3957,N_3832);
xor U4004 (N_4004,N_3860,N_3906);
xor U4005 (N_4005,N_3977,N_3923);
nand U4006 (N_4006,N_3925,N_3845);
or U4007 (N_4007,N_3822,N_3971);
xnor U4008 (N_4008,N_3824,N_3878);
nand U4009 (N_4009,N_3853,N_3934);
and U4010 (N_4010,N_3836,N_3983);
xor U4011 (N_4011,N_3852,N_3919);
or U4012 (N_4012,N_3828,N_3952);
or U4013 (N_4013,N_3933,N_3938);
xor U4014 (N_4014,N_3817,N_3931);
and U4015 (N_4015,N_3901,N_3967);
nand U4016 (N_4016,N_3823,N_3902);
xnor U4017 (N_4017,N_3911,N_3985);
xnor U4018 (N_4018,N_3871,N_3995);
nor U4019 (N_4019,N_3947,N_3968);
nor U4020 (N_4020,N_3825,N_3858);
nand U4021 (N_4021,N_3873,N_3924);
or U4022 (N_4022,N_3943,N_3863);
nand U4023 (N_4023,N_3810,N_3921);
xor U4024 (N_4024,N_3955,N_3864);
nor U4025 (N_4025,N_3956,N_3887);
xor U4026 (N_4026,N_3909,N_3900);
nand U4027 (N_4027,N_3989,N_3908);
nand U4028 (N_4028,N_3907,N_3868);
nand U4029 (N_4029,N_3937,N_3833);
or U4030 (N_4030,N_3866,N_3892);
or U4031 (N_4031,N_3800,N_3942);
or U4032 (N_4032,N_3959,N_3972);
nor U4033 (N_4033,N_3939,N_3904);
or U4034 (N_4034,N_3883,N_3963);
and U4035 (N_4035,N_3946,N_3862);
nand U4036 (N_4036,N_3888,N_3842);
and U4037 (N_4037,N_3803,N_3922);
and U4038 (N_4038,N_3949,N_3918);
or U4039 (N_4039,N_3889,N_3993);
or U4040 (N_4040,N_3896,N_3827);
nand U4041 (N_4041,N_3986,N_3880);
nand U4042 (N_4042,N_3984,N_3818);
xor U4043 (N_4043,N_3802,N_3999);
nand U4044 (N_4044,N_3912,N_3806);
nor U4045 (N_4045,N_3851,N_3847);
nor U4046 (N_4046,N_3855,N_3809);
and U4047 (N_4047,N_3976,N_3990);
nor U4048 (N_4048,N_3821,N_3874);
nor U4049 (N_4049,N_3819,N_3805);
and U4050 (N_4050,N_3981,N_3848);
and U4051 (N_4051,N_3897,N_3905);
nor U4052 (N_4052,N_3885,N_3849);
and U4053 (N_4053,N_3872,N_3926);
nor U4054 (N_4054,N_3978,N_3930);
or U4055 (N_4055,N_3932,N_3870);
and U4056 (N_4056,N_3867,N_3980);
nand U4057 (N_4057,N_3996,N_3898);
or U4058 (N_4058,N_3988,N_3831);
nand U4059 (N_4059,N_3987,N_3820);
or U4060 (N_4060,N_3877,N_3935);
or U4061 (N_4061,N_3826,N_3804);
nor U4062 (N_4062,N_3953,N_3910);
or U4063 (N_4063,N_3830,N_3895);
or U4064 (N_4064,N_3839,N_3929);
and U4065 (N_4065,N_3903,N_3886);
nand U4066 (N_4066,N_3997,N_3960);
xnor U4067 (N_4067,N_3927,N_3944);
or U4068 (N_4068,N_3893,N_3974);
xor U4069 (N_4069,N_3834,N_3835);
and U4070 (N_4070,N_3884,N_3808);
nor U4071 (N_4071,N_3917,N_3916);
and U4072 (N_4072,N_3973,N_3965);
and U4073 (N_4073,N_3865,N_3915);
and U4074 (N_4074,N_3869,N_3838);
and U4075 (N_4075,N_3970,N_3844);
and U4076 (N_4076,N_3941,N_3846);
nor U4077 (N_4077,N_3890,N_3814);
nand U4078 (N_4078,N_3920,N_3801);
or U4079 (N_4079,N_3891,N_3815);
or U4080 (N_4080,N_3969,N_3881);
nand U4081 (N_4081,N_3859,N_3879);
xor U4082 (N_4082,N_3928,N_3807);
nor U4083 (N_4083,N_3982,N_3854);
or U4084 (N_4084,N_3991,N_3899);
nand U4085 (N_4085,N_3936,N_3813);
or U4086 (N_4086,N_3940,N_3966);
nor U4087 (N_4087,N_3914,N_3948);
and U4088 (N_4088,N_3876,N_3829);
xor U4089 (N_4089,N_3861,N_3857);
nand U4090 (N_4090,N_3837,N_3950);
and U4091 (N_4091,N_3840,N_3882);
xnor U4092 (N_4092,N_3894,N_3811);
nor U4093 (N_4093,N_3875,N_3962);
or U4094 (N_4094,N_3816,N_3994);
nand U4095 (N_4095,N_3812,N_3843);
nor U4096 (N_4096,N_3998,N_3964);
or U4097 (N_4097,N_3841,N_3856);
nor U4098 (N_4098,N_3945,N_3958);
xnor U4099 (N_4099,N_3979,N_3951);
xnor U4100 (N_4100,N_3918,N_3977);
nor U4101 (N_4101,N_3852,N_3922);
xnor U4102 (N_4102,N_3921,N_3851);
or U4103 (N_4103,N_3924,N_3986);
xor U4104 (N_4104,N_3928,N_3878);
nor U4105 (N_4105,N_3865,N_3935);
xnor U4106 (N_4106,N_3881,N_3937);
xor U4107 (N_4107,N_3979,N_3915);
xor U4108 (N_4108,N_3892,N_3897);
nor U4109 (N_4109,N_3962,N_3828);
nand U4110 (N_4110,N_3866,N_3970);
nand U4111 (N_4111,N_3962,N_3915);
nand U4112 (N_4112,N_3852,N_3823);
nor U4113 (N_4113,N_3935,N_3911);
and U4114 (N_4114,N_3852,N_3833);
nor U4115 (N_4115,N_3936,N_3939);
or U4116 (N_4116,N_3972,N_3946);
or U4117 (N_4117,N_3932,N_3829);
or U4118 (N_4118,N_3960,N_3845);
xnor U4119 (N_4119,N_3977,N_3919);
nand U4120 (N_4120,N_3939,N_3892);
xnor U4121 (N_4121,N_3934,N_3978);
or U4122 (N_4122,N_3928,N_3951);
nand U4123 (N_4123,N_3887,N_3908);
and U4124 (N_4124,N_3870,N_3977);
and U4125 (N_4125,N_3987,N_3841);
xnor U4126 (N_4126,N_3971,N_3873);
xnor U4127 (N_4127,N_3946,N_3836);
or U4128 (N_4128,N_3946,N_3881);
or U4129 (N_4129,N_3917,N_3872);
xor U4130 (N_4130,N_3803,N_3992);
nor U4131 (N_4131,N_3879,N_3875);
nor U4132 (N_4132,N_3990,N_3912);
or U4133 (N_4133,N_3813,N_3824);
and U4134 (N_4134,N_3853,N_3938);
and U4135 (N_4135,N_3890,N_3938);
or U4136 (N_4136,N_3814,N_3857);
xnor U4137 (N_4137,N_3915,N_3984);
or U4138 (N_4138,N_3864,N_3839);
nand U4139 (N_4139,N_3813,N_3922);
or U4140 (N_4140,N_3868,N_3887);
xnor U4141 (N_4141,N_3886,N_3951);
xor U4142 (N_4142,N_3843,N_3897);
or U4143 (N_4143,N_3839,N_3818);
xor U4144 (N_4144,N_3900,N_3989);
nand U4145 (N_4145,N_3915,N_3904);
and U4146 (N_4146,N_3958,N_3840);
xnor U4147 (N_4147,N_3913,N_3833);
or U4148 (N_4148,N_3862,N_3834);
nand U4149 (N_4149,N_3846,N_3973);
or U4150 (N_4150,N_3844,N_3941);
or U4151 (N_4151,N_3908,N_3911);
nor U4152 (N_4152,N_3865,N_3931);
and U4153 (N_4153,N_3819,N_3912);
or U4154 (N_4154,N_3975,N_3935);
or U4155 (N_4155,N_3863,N_3997);
nor U4156 (N_4156,N_3859,N_3819);
xor U4157 (N_4157,N_3973,N_3975);
and U4158 (N_4158,N_3938,N_3834);
and U4159 (N_4159,N_3885,N_3803);
nand U4160 (N_4160,N_3890,N_3925);
nor U4161 (N_4161,N_3999,N_3899);
nor U4162 (N_4162,N_3884,N_3807);
and U4163 (N_4163,N_3824,N_3857);
or U4164 (N_4164,N_3943,N_3873);
nor U4165 (N_4165,N_3969,N_3927);
nand U4166 (N_4166,N_3963,N_3867);
nand U4167 (N_4167,N_3932,N_3924);
nor U4168 (N_4168,N_3923,N_3998);
or U4169 (N_4169,N_3803,N_3894);
nand U4170 (N_4170,N_3883,N_3894);
nand U4171 (N_4171,N_3952,N_3864);
nand U4172 (N_4172,N_3957,N_3959);
xnor U4173 (N_4173,N_3994,N_3807);
nor U4174 (N_4174,N_3841,N_3977);
and U4175 (N_4175,N_3863,N_3842);
or U4176 (N_4176,N_3852,N_3889);
and U4177 (N_4177,N_3919,N_3861);
nand U4178 (N_4178,N_3991,N_3947);
or U4179 (N_4179,N_3867,N_3899);
nor U4180 (N_4180,N_3875,N_3995);
xnor U4181 (N_4181,N_3807,N_3883);
nand U4182 (N_4182,N_3832,N_3876);
nor U4183 (N_4183,N_3809,N_3880);
or U4184 (N_4184,N_3873,N_3991);
nor U4185 (N_4185,N_3835,N_3902);
nand U4186 (N_4186,N_3810,N_3840);
and U4187 (N_4187,N_3887,N_3921);
nand U4188 (N_4188,N_3907,N_3903);
nor U4189 (N_4189,N_3823,N_3855);
xnor U4190 (N_4190,N_3884,N_3924);
nand U4191 (N_4191,N_3927,N_3942);
nand U4192 (N_4192,N_3841,N_3801);
nor U4193 (N_4193,N_3896,N_3965);
nor U4194 (N_4194,N_3936,N_3945);
nor U4195 (N_4195,N_3865,N_3877);
nand U4196 (N_4196,N_3962,N_3969);
xnor U4197 (N_4197,N_3918,N_3898);
nand U4198 (N_4198,N_3844,N_3961);
and U4199 (N_4199,N_3914,N_3953);
nand U4200 (N_4200,N_4129,N_4004);
or U4201 (N_4201,N_4183,N_4006);
xor U4202 (N_4202,N_4154,N_4116);
nor U4203 (N_4203,N_4167,N_4037);
or U4204 (N_4204,N_4185,N_4099);
xnor U4205 (N_4205,N_4094,N_4079);
or U4206 (N_4206,N_4070,N_4145);
and U4207 (N_4207,N_4127,N_4157);
or U4208 (N_4208,N_4069,N_4160);
or U4209 (N_4209,N_4056,N_4169);
nand U4210 (N_4210,N_4194,N_4189);
and U4211 (N_4211,N_4100,N_4149);
nor U4212 (N_4212,N_4098,N_4028);
nor U4213 (N_4213,N_4125,N_4151);
and U4214 (N_4214,N_4197,N_4140);
and U4215 (N_4215,N_4114,N_4104);
or U4216 (N_4216,N_4097,N_4150);
and U4217 (N_4217,N_4192,N_4077);
or U4218 (N_4218,N_4180,N_4193);
nor U4219 (N_4219,N_4175,N_4158);
and U4220 (N_4220,N_4075,N_4071);
xnor U4221 (N_4221,N_4113,N_4110);
or U4222 (N_4222,N_4041,N_4090);
and U4223 (N_4223,N_4044,N_4179);
nor U4224 (N_4224,N_4186,N_4024);
or U4225 (N_4225,N_4136,N_4184);
nand U4226 (N_4226,N_4188,N_4020);
or U4227 (N_4227,N_4091,N_4195);
and U4228 (N_4228,N_4173,N_4080);
nor U4229 (N_4229,N_4132,N_4134);
nand U4230 (N_4230,N_4139,N_4051);
nor U4231 (N_4231,N_4034,N_4081);
and U4232 (N_4232,N_4128,N_4187);
nand U4233 (N_4233,N_4049,N_4138);
or U4234 (N_4234,N_4121,N_4065);
nor U4235 (N_4235,N_4074,N_4066);
nand U4236 (N_4236,N_4115,N_4148);
xor U4237 (N_4237,N_4043,N_4111);
or U4238 (N_4238,N_4022,N_4038);
nand U4239 (N_4239,N_4102,N_4086);
xnor U4240 (N_4240,N_4085,N_4003);
and U4241 (N_4241,N_4096,N_4103);
or U4242 (N_4242,N_4163,N_4019);
and U4243 (N_4243,N_4053,N_4172);
nand U4244 (N_4244,N_4147,N_4182);
xor U4245 (N_4245,N_4068,N_4040);
nand U4246 (N_4246,N_4047,N_4010);
and U4247 (N_4247,N_4153,N_4118);
nor U4248 (N_4248,N_4124,N_4055);
nor U4249 (N_4249,N_4058,N_4048);
nor U4250 (N_4250,N_4108,N_4029);
or U4251 (N_4251,N_4120,N_4026);
nand U4252 (N_4252,N_4015,N_4067);
and U4253 (N_4253,N_4000,N_4165);
or U4254 (N_4254,N_4122,N_4162);
or U4255 (N_4255,N_4084,N_4072);
nor U4256 (N_4256,N_4057,N_4161);
or U4257 (N_4257,N_4119,N_4198);
or U4258 (N_4258,N_4107,N_4059);
and U4259 (N_4259,N_4046,N_4045);
nor U4260 (N_4260,N_4141,N_4076);
or U4261 (N_4261,N_4177,N_4143);
nand U4262 (N_4262,N_4061,N_4166);
nand U4263 (N_4263,N_4078,N_4033);
xnor U4264 (N_4264,N_4190,N_4036);
nor U4265 (N_4265,N_4021,N_4087);
or U4266 (N_4266,N_4027,N_4105);
or U4267 (N_4267,N_4133,N_4089);
xor U4268 (N_4268,N_4168,N_4191);
xnor U4269 (N_4269,N_4032,N_4176);
or U4270 (N_4270,N_4025,N_4106);
xnor U4271 (N_4271,N_4052,N_4093);
or U4272 (N_4272,N_4073,N_4013);
and U4273 (N_4273,N_4001,N_4171);
xnor U4274 (N_4274,N_4156,N_4060);
xnor U4275 (N_4275,N_4170,N_4088);
nand U4276 (N_4276,N_4063,N_4155);
nand U4277 (N_4277,N_4050,N_4109);
or U4278 (N_4278,N_4016,N_4199);
nor U4279 (N_4279,N_4137,N_4126);
nand U4280 (N_4280,N_4112,N_4007);
xor U4281 (N_4281,N_4130,N_4083);
and U4282 (N_4282,N_4117,N_4082);
nand U4283 (N_4283,N_4018,N_4002);
nor U4284 (N_4284,N_4164,N_4012);
nor U4285 (N_4285,N_4005,N_4131);
xor U4286 (N_4286,N_4196,N_4011);
nand U4287 (N_4287,N_4142,N_4144);
and U4288 (N_4288,N_4035,N_4178);
nor U4289 (N_4289,N_4054,N_4159);
or U4290 (N_4290,N_4101,N_4042);
and U4291 (N_4291,N_4030,N_4062);
and U4292 (N_4292,N_4095,N_4031);
and U4293 (N_4293,N_4017,N_4135);
and U4294 (N_4294,N_4092,N_4014);
nand U4295 (N_4295,N_4181,N_4123);
nand U4296 (N_4296,N_4023,N_4152);
or U4297 (N_4297,N_4008,N_4146);
and U4298 (N_4298,N_4064,N_4174);
or U4299 (N_4299,N_4039,N_4009);
nor U4300 (N_4300,N_4109,N_4093);
nand U4301 (N_4301,N_4094,N_4179);
and U4302 (N_4302,N_4094,N_4082);
and U4303 (N_4303,N_4030,N_4111);
or U4304 (N_4304,N_4184,N_4145);
xnor U4305 (N_4305,N_4082,N_4034);
xnor U4306 (N_4306,N_4063,N_4159);
nand U4307 (N_4307,N_4078,N_4096);
or U4308 (N_4308,N_4163,N_4016);
and U4309 (N_4309,N_4060,N_4035);
nand U4310 (N_4310,N_4031,N_4054);
nor U4311 (N_4311,N_4151,N_4019);
and U4312 (N_4312,N_4111,N_4104);
nand U4313 (N_4313,N_4120,N_4112);
and U4314 (N_4314,N_4002,N_4049);
nand U4315 (N_4315,N_4051,N_4021);
xnor U4316 (N_4316,N_4138,N_4164);
xnor U4317 (N_4317,N_4069,N_4165);
nor U4318 (N_4318,N_4112,N_4027);
nand U4319 (N_4319,N_4030,N_4053);
or U4320 (N_4320,N_4000,N_4056);
or U4321 (N_4321,N_4004,N_4184);
nor U4322 (N_4322,N_4099,N_4048);
or U4323 (N_4323,N_4113,N_4024);
and U4324 (N_4324,N_4059,N_4092);
nor U4325 (N_4325,N_4026,N_4114);
xor U4326 (N_4326,N_4132,N_4166);
nand U4327 (N_4327,N_4130,N_4107);
or U4328 (N_4328,N_4018,N_4192);
nor U4329 (N_4329,N_4009,N_4155);
xor U4330 (N_4330,N_4101,N_4038);
or U4331 (N_4331,N_4177,N_4093);
nor U4332 (N_4332,N_4079,N_4014);
nor U4333 (N_4333,N_4054,N_4000);
or U4334 (N_4334,N_4017,N_4059);
and U4335 (N_4335,N_4017,N_4167);
nand U4336 (N_4336,N_4089,N_4071);
and U4337 (N_4337,N_4082,N_4137);
or U4338 (N_4338,N_4192,N_4062);
and U4339 (N_4339,N_4130,N_4034);
or U4340 (N_4340,N_4177,N_4121);
or U4341 (N_4341,N_4057,N_4189);
nand U4342 (N_4342,N_4182,N_4194);
or U4343 (N_4343,N_4127,N_4187);
nand U4344 (N_4344,N_4028,N_4082);
xnor U4345 (N_4345,N_4008,N_4190);
and U4346 (N_4346,N_4180,N_4150);
xnor U4347 (N_4347,N_4108,N_4117);
or U4348 (N_4348,N_4003,N_4047);
nor U4349 (N_4349,N_4107,N_4110);
nor U4350 (N_4350,N_4123,N_4097);
and U4351 (N_4351,N_4009,N_4098);
xnor U4352 (N_4352,N_4049,N_4153);
nor U4353 (N_4353,N_4030,N_4126);
and U4354 (N_4354,N_4157,N_4047);
and U4355 (N_4355,N_4173,N_4192);
xnor U4356 (N_4356,N_4156,N_4123);
xor U4357 (N_4357,N_4067,N_4102);
and U4358 (N_4358,N_4008,N_4157);
nor U4359 (N_4359,N_4070,N_4149);
nor U4360 (N_4360,N_4105,N_4176);
and U4361 (N_4361,N_4177,N_4164);
nand U4362 (N_4362,N_4192,N_4162);
nor U4363 (N_4363,N_4185,N_4018);
and U4364 (N_4364,N_4034,N_4009);
or U4365 (N_4365,N_4003,N_4154);
nor U4366 (N_4366,N_4078,N_4044);
xnor U4367 (N_4367,N_4024,N_4179);
xor U4368 (N_4368,N_4182,N_4135);
and U4369 (N_4369,N_4016,N_4021);
and U4370 (N_4370,N_4120,N_4166);
and U4371 (N_4371,N_4184,N_4056);
xor U4372 (N_4372,N_4044,N_4151);
nor U4373 (N_4373,N_4019,N_4174);
nor U4374 (N_4374,N_4018,N_4179);
or U4375 (N_4375,N_4058,N_4015);
xor U4376 (N_4376,N_4089,N_4004);
xnor U4377 (N_4377,N_4008,N_4152);
or U4378 (N_4378,N_4192,N_4113);
or U4379 (N_4379,N_4134,N_4187);
and U4380 (N_4380,N_4031,N_4053);
nand U4381 (N_4381,N_4043,N_4001);
or U4382 (N_4382,N_4114,N_4143);
and U4383 (N_4383,N_4131,N_4187);
nor U4384 (N_4384,N_4124,N_4120);
xnor U4385 (N_4385,N_4164,N_4085);
nor U4386 (N_4386,N_4101,N_4024);
nor U4387 (N_4387,N_4177,N_4172);
xor U4388 (N_4388,N_4195,N_4047);
and U4389 (N_4389,N_4023,N_4070);
nand U4390 (N_4390,N_4054,N_4166);
xnor U4391 (N_4391,N_4131,N_4156);
nor U4392 (N_4392,N_4005,N_4120);
nor U4393 (N_4393,N_4113,N_4142);
and U4394 (N_4394,N_4188,N_4063);
and U4395 (N_4395,N_4145,N_4085);
and U4396 (N_4396,N_4050,N_4087);
nor U4397 (N_4397,N_4042,N_4117);
or U4398 (N_4398,N_4064,N_4051);
nand U4399 (N_4399,N_4192,N_4187);
xor U4400 (N_4400,N_4370,N_4365);
xnor U4401 (N_4401,N_4243,N_4266);
nor U4402 (N_4402,N_4241,N_4338);
nor U4403 (N_4403,N_4286,N_4357);
nor U4404 (N_4404,N_4358,N_4326);
nor U4405 (N_4405,N_4306,N_4354);
or U4406 (N_4406,N_4228,N_4232);
xnor U4407 (N_4407,N_4356,N_4274);
or U4408 (N_4408,N_4230,N_4353);
and U4409 (N_4409,N_4360,N_4296);
xor U4410 (N_4410,N_4307,N_4283);
nor U4411 (N_4411,N_4304,N_4214);
xnor U4412 (N_4412,N_4277,N_4205);
and U4413 (N_4413,N_4394,N_4219);
and U4414 (N_4414,N_4318,N_4250);
nand U4415 (N_4415,N_4227,N_4330);
nand U4416 (N_4416,N_4213,N_4217);
and U4417 (N_4417,N_4381,N_4239);
or U4418 (N_4418,N_4380,N_4313);
nand U4419 (N_4419,N_4280,N_4305);
nand U4420 (N_4420,N_4346,N_4324);
xor U4421 (N_4421,N_4351,N_4206);
nand U4422 (N_4422,N_4229,N_4233);
xor U4423 (N_4423,N_4308,N_4385);
nor U4424 (N_4424,N_4361,N_4235);
and U4425 (N_4425,N_4278,N_4222);
nand U4426 (N_4426,N_4387,N_4398);
nand U4427 (N_4427,N_4271,N_4234);
nor U4428 (N_4428,N_4345,N_4275);
nor U4429 (N_4429,N_4221,N_4236);
xor U4430 (N_4430,N_4389,N_4363);
and U4431 (N_4431,N_4382,N_4355);
xor U4432 (N_4432,N_4224,N_4281);
or U4433 (N_4433,N_4316,N_4253);
nand U4434 (N_4434,N_4334,N_4349);
xnor U4435 (N_4435,N_4264,N_4268);
nand U4436 (N_4436,N_4263,N_4270);
nor U4437 (N_4437,N_4362,N_4240);
nor U4438 (N_4438,N_4203,N_4320);
and U4439 (N_4439,N_4279,N_4367);
nor U4440 (N_4440,N_4294,N_4254);
xor U4441 (N_4441,N_4244,N_4285);
xnor U4442 (N_4442,N_4272,N_4300);
or U4443 (N_4443,N_4237,N_4395);
nor U4444 (N_4444,N_4210,N_4225);
nor U4445 (N_4445,N_4384,N_4276);
xor U4446 (N_4446,N_4379,N_4303);
nand U4447 (N_4447,N_4383,N_4238);
nand U4448 (N_4448,N_4332,N_4340);
or U4449 (N_4449,N_4317,N_4339);
nor U4450 (N_4450,N_4374,N_4377);
nand U4451 (N_4451,N_4267,N_4298);
nor U4452 (N_4452,N_4397,N_4226);
xor U4453 (N_4453,N_4329,N_4399);
xor U4454 (N_4454,N_4375,N_4328);
xor U4455 (N_4455,N_4297,N_4200);
xor U4456 (N_4456,N_4269,N_4341);
xor U4457 (N_4457,N_4388,N_4252);
nor U4458 (N_4458,N_4255,N_4315);
or U4459 (N_4459,N_4323,N_4299);
nor U4460 (N_4460,N_4212,N_4390);
or U4461 (N_4461,N_4314,N_4372);
nor U4462 (N_4462,N_4311,N_4260);
nand U4463 (N_4463,N_4261,N_4287);
nor U4464 (N_4464,N_4310,N_4215);
nand U4465 (N_4465,N_4218,N_4216);
and U4466 (N_4466,N_4378,N_4301);
xnor U4467 (N_4467,N_4208,N_4392);
and U4468 (N_4468,N_4333,N_4327);
and U4469 (N_4469,N_4242,N_4202);
nor U4470 (N_4470,N_4352,N_4325);
nand U4471 (N_4471,N_4248,N_4204);
and U4472 (N_4472,N_4246,N_4309);
and U4473 (N_4473,N_4376,N_4220);
nor U4474 (N_4474,N_4211,N_4288);
and U4475 (N_4475,N_4347,N_4350);
xor U4476 (N_4476,N_4247,N_4284);
nand U4477 (N_4477,N_4312,N_4291);
nand U4478 (N_4478,N_4386,N_4282);
or U4479 (N_4479,N_4335,N_4348);
and U4480 (N_4480,N_4259,N_4369);
xnor U4481 (N_4481,N_4231,N_4223);
nor U4482 (N_4482,N_4256,N_4265);
or U4483 (N_4483,N_4262,N_4373);
or U4484 (N_4484,N_4251,N_4249);
xor U4485 (N_4485,N_4336,N_4319);
xor U4486 (N_4486,N_4391,N_4368);
and U4487 (N_4487,N_4258,N_4302);
nor U4488 (N_4488,N_4344,N_4337);
xnor U4489 (N_4489,N_4290,N_4321);
nand U4490 (N_4490,N_4366,N_4396);
or U4491 (N_4491,N_4295,N_4342);
nor U4492 (N_4492,N_4207,N_4201);
nand U4493 (N_4493,N_4292,N_4371);
or U4494 (N_4494,N_4331,N_4273);
and U4495 (N_4495,N_4293,N_4359);
and U4496 (N_4496,N_4257,N_4364);
nand U4497 (N_4497,N_4343,N_4209);
xor U4498 (N_4498,N_4289,N_4245);
and U4499 (N_4499,N_4322,N_4393);
nor U4500 (N_4500,N_4395,N_4312);
or U4501 (N_4501,N_4208,N_4239);
and U4502 (N_4502,N_4299,N_4300);
nand U4503 (N_4503,N_4287,N_4307);
xnor U4504 (N_4504,N_4362,N_4241);
nor U4505 (N_4505,N_4243,N_4384);
and U4506 (N_4506,N_4258,N_4387);
xor U4507 (N_4507,N_4314,N_4336);
and U4508 (N_4508,N_4373,N_4385);
or U4509 (N_4509,N_4245,N_4217);
xor U4510 (N_4510,N_4271,N_4224);
nor U4511 (N_4511,N_4354,N_4247);
nor U4512 (N_4512,N_4234,N_4379);
nand U4513 (N_4513,N_4293,N_4252);
nor U4514 (N_4514,N_4368,N_4352);
xnor U4515 (N_4515,N_4209,N_4320);
and U4516 (N_4516,N_4298,N_4314);
nand U4517 (N_4517,N_4210,N_4223);
xor U4518 (N_4518,N_4311,N_4258);
nand U4519 (N_4519,N_4311,N_4302);
nor U4520 (N_4520,N_4321,N_4202);
and U4521 (N_4521,N_4283,N_4326);
or U4522 (N_4522,N_4388,N_4275);
nand U4523 (N_4523,N_4375,N_4278);
or U4524 (N_4524,N_4299,N_4318);
and U4525 (N_4525,N_4222,N_4391);
and U4526 (N_4526,N_4239,N_4288);
xnor U4527 (N_4527,N_4306,N_4292);
and U4528 (N_4528,N_4389,N_4395);
nand U4529 (N_4529,N_4255,N_4296);
or U4530 (N_4530,N_4228,N_4205);
and U4531 (N_4531,N_4267,N_4294);
or U4532 (N_4532,N_4273,N_4282);
nor U4533 (N_4533,N_4274,N_4230);
and U4534 (N_4534,N_4208,N_4379);
or U4535 (N_4535,N_4329,N_4210);
xnor U4536 (N_4536,N_4284,N_4252);
nand U4537 (N_4537,N_4339,N_4250);
xor U4538 (N_4538,N_4336,N_4375);
xnor U4539 (N_4539,N_4245,N_4329);
or U4540 (N_4540,N_4259,N_4234);
nand U4541 (N_4541,N_4264,N_4337);
xnor U4542 (N_4542,N_4276,N_4234);
or U4543 (N_4543,N_4327,N_4279);
or U4544 (N_4544,N_4366,N_4325);
nor U4545 (N_4545,N_4330,N_4339);
nor U4546 (N_4546,N_4379,N_4324);
or U4547 (N_4547,N_4225,N_4311);
xnor U4548 (N_4548,N_4343,N_4304);
or U4549 (N_4549,N_4246,N_4290);
and U4550 (N_4550,N_4294,N_4253);
nor U4551 (N_4551,N_4368,N_4234);
nand U4552 (N_4552,N_4257,N_4297);
and U4553 (N_4553,N_4223,N_4215);
or U4554 (N_4554,N_4364,N_4350);
nand U4555 (N_4555,N_4390,N_4267);
and U4556 (N_4556,N_4399,N_4352);
or U4557 (N_4557,N_4321,N_4338);
xor U4558 (N_4558,N_4335,N_4362);
or U4559 (N_4559,N_4239,N_4262);
nor U4560 (N_4560,N_4208,N_4381);
and U4561 (N_4561,N_4345,N_4363);
nand U4562 (N_4562,N_4384,N_4246);
and U4563 (N_4563,N_4318,N_4248);
nand U4564 (N_4564,N_4369,N_4285);
and U4565 (N_4565,N_4339,N_4320);
or U4566 (N_4566,N_4238,N_4333);
nor U4567 (N_4567,N_4218,N_4274);
nor U4568 (N_4568,N_4219,N_4310);
or U4569 (N_4569,N_4284,N_4262);
nand U4570 (N_4570,N_4283,N_4393);
xnor U4571 (N_4571,N_4217,N_4369);
and U4572 (N_4572,N_4302,N_4240);
xnor U4573 (N_4573,N_4319,N_4219);
nand U4574 (N_4574,N_4317,N_4215);
nand U4575 (N_4575,N_4226,N_4369);
xor U4576 (N_4576,N_4208,N_4302);
or U4577 (N_4577,N_4367,N_4324);
nand U4578 (N_4578,N_4357,N_4201);
nor U4579 (N_4579,N_4277,N_4268);
xnor U4580 (N_4580,N_4219,N_4226);
or U4581 (N_4581,N_4290,N_4221);
nor U4582 (N_4582,N_4346,N_4274);
xnor U4583 (N_4583,N_4389,N_4283);
nor U4584 (N_4584,N_4335,N_4200);
or U4585 (N_4585,N_4372,N_4320);
nor U4586 (N_4586,N_4297,N_4389);
xnor U4587 (N_4587,N_4337,N_4396);
or U4588 (N_4588,N_4301,N_4344);
xnor U4589 (N_4589,N_4347,N_4356);
nor U4590 (N_4590,N_4287,N_4269);
or U4591 (N_4591,N_4348,N_4277);
nand U4592 (N_4592,N_4367,N_4201);
and U4593 (N_4593,N_4237,N_4203);
nor U4594 (N_4594,N_4205,N_4368);
nand U4595 (N_4595,N_4280,N_4355);
nand U4596 (N_4596,N_4390,N_4247);
nand U4597 (N_4597,N_4316,N_4278);
nand U4598 (N_4598,N_4352,N_4247);
nor U4599 (N_4599,N_4328,N_4349);
or U4600 (N_4600,N_4474,N_4476);
or U4601 (N_4601,N_4407,N_4463);
nor U4602 (N_4602,N_4459,N_4576);
or U4603 (N_4603,N_4557,N_4580);
and U4604 (N_4604,N_4439,N_4428);
nor U4605 (N_4605,N_4539,N_4482);
nor U4606 (N_4606,N_4552,N_4418);
nand U4607 (N_4607,N_4414,N_4537);
nand U4608 (N_4608,N_4421,N_4560);
or U4609 (N_4609,N_4493,N_4487);
nor U4610 (N_4610,N_4511,N_4483);
nor U4611 (N_4611,N_4533,N_4462);
nor U4612 (N_4612,N_4598,N_4571);
nand U4613 (N_4613,N_4460,N_4410);
nand U4614 (N_4614,N_4412,N_4561);
xnor U4615 (N_4615,N_4570,N_4540);
or U4616 (N_4616,N_4440,N_4424);
xnor U4617 (N_4617,N_4575,N_4535);
nor U4618 (N_4618,N_4456,N_4534);
xnor U4619 (N_4619,N_4530,N_4595);
nor U4620 (N_4620,N_4492,N_4507);
nand U4621 (N_4621,N_4455,N_4422);
xnor U4622 (N_4622,N_4567,N_4505);
and U4623 (N_4623,N_4502,N_4510);
and U4624 (N_4624,N_4581,N_4568);
or U4625 (N_4625,N_4433,N_4472);
nand U4626 (N_4626,N_4520,N_4579);
and U4627 (N_4627,N_4402,N_4430);
nor U4628 (N_4628,N_4447,N_4548);
or U4629 (N_4629,N_4409,N_4469);
xnor U4630 (N_4630,N_4542,N_4411);
or U4631 (N_4631,N_4438,N_4431);
or U4632 (N_4632,N_4498,N_4450);
or U4633 (N_4633,N_4429,N_4513);
nor U4634 (N_4634,N_4521,N_4558);
or U4635 (N_4635,N_4585,N_4432);
and U4636 (N_4636,N_4522,N_4559);
and U4637 (N_4637,N_4536,N_4471);
nand U4638 (N_4638,N_4427,N_4484);
xor U4639 (N_4639,N_4566,N_4441);
nor U4640 (N_4640,N_4478,N_4479);
nor U4641 (N_4641,N_4490,N_4408);
xor U4642 (N_4642,N_4420,N_4413);
nand U4643 (N_4643,N_4517,N_4519);
nand U4644 (N_4644,N_4437,N_4443);
nand U4645 (N_4645,N_4596,N_4504);
or U4646 (N_4646,N_4594,N_4515);
nor U4647 (N_4647,N_4508,N_4445);
and U4648 (N_4648,N_4403,N_4400);
and U4649 (N_4649,N_4480,N_4562);
and U4650 (N_4650,N_4499,N_4587);
nand U4651 (N_4651,N_4494,N_4458);
nor U4652 (N_4652,N_4401,N_4582);
and U4653 (N_4653,N_4577,N_4541);
xnor U4654 (N_4654,N_4453,N_4491);
or U4655 (N_4655,N_4547,N_4436);
or U4656 (N_4656,N_4551,N_4564);
xnor U4657 (N_4657,N_4518,N_4470);
xor U4658 (N_4658,N_4496,N_4565);
or U4659 (N_4659,N_4554,N_4543);
xor U4660 (N_4660,N_4526,N_4444);
xnor U4661 (N_4661,N_4574,N_4415);
nor U4662 (N_4662,N_4528,N_4588);
and U4663 (N_4663,N_4544,N_4531);
nand U4664 (N_4664,N_4464,N_4452);
and U4665 (N_4665,N_4591,N_4473);
nor U4666 (N_4666,N_4523,N_4553);
nor U4667 (N_4667,N_4468,N_4516);
xnor U4668 (N_4668,N_4488,N_4524);
nand U4669 (N_4669,N_4572,N_4495);
or U4670 (N_4670,N_4417,N_4529);
or U4671 (N_4671,N_4477,N_4538);
nand U4672 (N_4672,N_4426,N_4593);
xor U4673 (N_4673,N_4556,N_4597);
xnor U4674 (N_4674,N_4563,N_4419);
nand U4675 (N_4675,N_4512,N_4405);
and U4676 (N_4676,N_4573,N_4532);
xnor U4677 (N_4677,N_4435,N_4461);
nand U4678 (N_4678,N_4466,N_4501);
nand U4679 (N_4679,N_4457,N_4509);
xor U4680 (N_4680,N_4586,N_4583);
nor U4681 (N_4681,N_4446,N_4525);
and U4682 (N_4682,N_4599,N_4448);
and U4683 (N_4683,N_4550,N_4584);
nand U4684 (N_4684,N_4569,N_4489);
nor U4685 (N_4685,N_4449,N_4506);
and U4686 (N_4686,N_4434,N_4590);
xnor U4687 (N_4687,N_4423,N_4465);
nor U4688 (N_4688,N_4404,N_4454);
nor U4689 (N_4689,N_4500,N_4545);
or U4690 (N_4690,N_4416,N_4406);
and U4691 (N_4691,N_4549,N_4475);
nor U4692 (N_4692,N_4527,N_4485);
nor U4693 (N_4693,N_4592,N_4589);
nor U4694 (N_4694,N_4442,N_4481);
xnor U4695 (N_4695,N_4578,N_4425);
xor U4696 (N_4696,N_4546,N_4514);
and U4697 (N_4697,N_4555,N_4497);
nor U4698 (N_4698,N_4486,N_4451);
and U4699 (N_4699,N_4503,N_4467);
nand U4700 (N_4700,N_4502,N_4507);
and U4701 (N_4701,N_4499,N_4420);
nand U4702 (N_4702,N_4489,N_4469);
nand U4703 (N_4703,N_4584,N_4551);
or U4704 (N_4704,N_4582,N_4439);
and U4705 (N_4705,N_4562,N_4507);
and U4706 (N_4706,N_4487,N_4458);
nand U4707 (N_4707,N_4568,N_4495);
xor U4708 (N_4708,N_4451,N_4477);
or U4709 (N_4709,N_4549,N_4522);
xor U4710 (N_4710,N_4564,N_4575);
nand U4711 (N_4711,N_4546,N_4457);
xnor U4712 (N_4712,N_4541,N_4528);
nor U4713 (N_4713,N_4431,N_4405);
or U4714 (N_4714,N_4546,N_4415);
and U4715 (N_4715,N_4422,N_4543);
nor U4716 (N_4716,N_4429,N_4542);
and U4717 (N_4717,N_4511,N_4525);
and U4718 (N_4718,N_4437,N_4538);
xor U4719 (N_4719,N_4492,N_4429);
or U4720 (N_4720,N_4425,N_4529);
nor U4721 (N_4721,N_4512,N_4455);
and U4722 (N_4722,N_4440,N_4429);
nand U4723 (N_4723,N_4473,N_4468);
and U4724 (N_4724,N_4457,N_4551);
nand U4725 (N_4725,N_4450,N_4406);
or U4726 (N_4726,N_4510,N_4466);
and U4727 (N_4727,N_4540,N_4400);
nand U4728 (N_4728,N_4473,N_4519);
xnor U4729 (N_4729,N_4520,N_4400);
nor U4730 (N_4730,N_4413,N_4453);
xnor U4731 (N_4731,N_4476,N_4498);
nand U4732 (N_4732,N_4535,N_4483);
nand U4733 (N_4733,N_4486,N_4434);
nor U4734 (N_4734,N_4574,N_4582);
xor U4735 (N_4735,N_4537,N_4513);
and U4736 (N_4736,N_4422,N_4563);
xnor U4737 (N_4737,N_4537,N_4481);
and U4738 (N_4738,N_4469,N_4467);
and U4739 (N_4739,N_4531,N_4598);
or U4740 (N_4740,N_4418,N_4558);
or U4741 (N_4741,N_4409,N_4523);
xnor U4742 (N_4742,N_4515,N_4524);
xnor U4743 (N_4743,N_4456,N_4459);
nand U4744 (N_4744,N_4564,N_4419);
and U4745 (N_4745,N_4409,N_4441);
and U4746 (N_4746,N_4529,N_4554);
or U4747 (N_4747,N_4521,N_4525);
and U4748 (N_4748,N_4440,N_4425);
or U4749 (N_4749,N_4453,N_4430);
and U4750 (N_4750,N_4513,N_4418);
nor U4751 (N_4751,N_4574,N_4446);
or U4752 (N_4752,N_4525,N_4578);
and U4753 (N_4753,N_4402,N_4400);
or U4754 (N_4754,N_4555,N_4568);
xnor U4755 (N_4755,N_4403,N_4464);
and U4756 (N_4756,N_4521,N_4421);
xnor U4757 (N_4757,N_4494,N_4506);
or U4758 (N_4758,N_4459,N_4430);
nor U4759 (N_4759,N_4530,N_4532);
nor U4760 (N_4760,N_4516,N_4511);
xor U4761 (N_4761,N_4543,N_4576);
nor U4762 (N_4762,N_4556,N_4568);
and U4763 (N_4763,N_4417,N_4479);
nor U4764 (N_4764,N_4496,N_4428);
nand U4765 (N_4765,N_4430,N_4418);
nor U4766 (N_4766,N_4577,N_4508);
or U4767 (N_4767,N_4402,N_4432);
or U4768 (N_4768,N_4542,N_4555);
and U4769 (N_4769,N_4553,N_4519);
xor U4770 (N_4770,N_4537,N_4413);
xor U4771 (N_4771,N_4406,N_4453);
and U4772 (N_4772,N_4497,N_4509);
or U4773 (N_4773,N_4578,N_4513);
nor U4774 (N_4774,N_4522,N_4468);
nor U4775 (N_4775,N_4462,N_4465);
xnor U4776 (N_4776,N_4457,N_4589);
and U4777 (N_4777,N_4424,N_4518);
and U4778 (N_4778,N_4409,N_4543);
and U4779 (N_4779,N_4517,N_4401);
and U4780 (N_4780,N_4596,N_4591);
or U4781 (N_4781,N_4489,N_4451);
or U4782 (N_4782,N_4413,N_4540);
nor U4783 (N_4783,N_4480,N_4463);
nand U4784 (N_4784,N_4433,N_4425);
nor U4785 (N_4785,N_4575,N_4453);
nand U4786 (N_4786,N_4414,N_4448);
xnor U4787 (N_4787,N_4408,N_4515);
and U4788 (N_4788,N_4545,N_4449);
nor U4789 (N_4789,N_4431,N_4554);
xor U4790 (N_4790,N_4496,N_4585);
and U4791 (N_4791,N_4478,N_4549);
nor U4792 (N_4792,N_4462,N_4511);
nand U4793 (N_4793,N_4523,N_4400);
xor U4794 (N_4794,N_4416,N_4455);
xnor U4795 (N_4795,N_4520,N_4483);
and U4796 (N_4796,N_4594,N_4503);
nand U4797 (N_4797,N_4525,N_4457);
nand U4798 (N_4798,N_4549,N_4438);
nand U4799 (N_4799,N_4492,N_4568);
xnor U4800 (N_4800,N_4615,N_4634);
and U4801 (N_4801,N_4704,N_4745);
nand U4802 (N_4802,N_4628,N_4609);
nand U4803 (N_4803,N_4719,N_4669);
and U4804 (N_4804,N_4630,N_4608);
or U4805 (N_4805,N_4759,N_4706);
or U4806 (N_4806,N_4671,N_4657);
xor U4807 (N_4807,N_4638,N_4649);
nor U4808 (N_4808,N_4784,N_4661);
and U4809 (N_4809,N_4764,N_4720);
xor U4810 (N_4810,N_4731,N_4748);
xnor U4811 (N_4811,N_4652,N_4667);
xnor U4812 (N_4812,N_4740,N_4767);
nor U4813 (N_4813,N_4697,N_4780);
and U4814 (N_4814,N_4774,N_4665);
or U4815 (N_4815,N_4680,N_4610);
or U4816 (N_4816,N_4741,N_4768);
or U4817 (N_4817,N_4729,N_4632);
nand U4818 (N_4818,N_4737,N_4646);
and U4819 (N_4819,N_4711,N_4633);
nor U4820 (N_4820,N_4676,N_4716);
xor U4821 (N_4821,N_4700,N_4755);
nor U4822 (N_4822,N_4692,N_4668);
nand U4823 (N_4823,N_4606,N_4637);
nor U4824 (N_4824,N_4777,N_4749);
and U4825 (N_4825,N_4756,N_4795);
nand U4826 (N_4826,N_4732,N_4611);
and U4827 (N_4827,N_4710,N_4738);
nor U4828 (N_4828,N_4799,N_4654);
and U4829 (N_4829,N_4771,N_4651);
and U4830 (N_4830,N_4666,N_4779);
nand U4831 (N_4831,N_4742,N_4778);
nand U4832 (N_4832,N_4757,N_4765);
xor U4833 (N_4833,N_4659,N_4708);
nand U4834 (N_4834,N_4790,N_4739);
xor U4835 (N_4835,N_4717,N_4673);
nor U4836 (N_4836,N_4624,N_4735);
or U4837 (N_4837,N_4715,N_4612);
xnor U4838 (N_4838,N_4734,N_4696);
or U4839 (N_4839,N_4725,N_4605);
or U4840 (N_4840,N_4678,N_4698);
nand U4841 (N_4841,N_4629,N_4641);
or U4842 (N_4842,N_4662,N_4644);
and U4843 (N_4843,N_4714,N_4766);
nand U4844 (N_4844,N_4601,N_4761);
and U4845 (N_4845,N_4685,N_4792);
nand U4846 (N_4846,N_4760,N_4702);
nor U4847 (N_4847,N_4619,N_4684);
nor U4848 (N_4848,N_4693,N_4603);
and U4849 (N_4849,N_4794,N_4726);
or U4850 (N_4850,N_4770,N_4683);
and U4851 (N_4851,N_4713,N_4650);
xor U4852 (N_4852,N_4688,N_4712);
xnor U4853 (N_4853,N_4751,N_4798);
nor U4854 (N_4854,N_4754,N_4769);
nand U4855 (N_4855,N_4635,N_4747);
nor U4856 (N_4856,N_4658,N_4721);
or U4857 (N_4857,N_4727,N_4627);
nand U4858 (N_4858,N_4783,N_4604);
and U4859 (N_4859,N_4736,N_4750);
xor U4860 (N_4860,N_4786,N_4622);
nand U4861 (N_4861,N_4643,N_4775);
or U4862 (N_4862,N_4655,N_4607);
nand U4863 (N_4863,N_4660,N_4631);
nand U4864 (N_4864,N_4656,N_4620);
nor U4865 (N_4865,N_4782,N_4724);
and U4866 (N_4866,N_4772,N_4733);
and U4867 (N_4867,N_4776,N_4625);
nand U4868 (N_4868,N_4743,N_4796);
or U4869 (N_4869,N_4753,N_4695);
xnor U4870 (N_4870,N_4648,N_4718);
and U4871 (N_4871,N_4752,N_4705);
xnor U4872 (N_4872,N_4707,N_4618);
and U4873 (N_4873,N_4763,N_4699);
xnor U4874 (N_4874,N_4600,N_4614);
and U4875 (N_4875,N_4787,N_4640);
nand U4876 (N_4876,N_4728,N_4788);
xnor U4877 (N_4877,N_4773,N_4789);
xnor U4878 (N_4878,N_4616,N_4691);
and U4879 (N_4879,N_4703,N_4709);
or U4880 (N_4880,N_4690,N_4617);
nand U4881 (N_4881,N_4687,N_4653);
and U4882 (N_4882,N_4613,N_4670);
nor U4883 (N_4883,N_4758,N_4672);
nor U4884 (N_4884,N_4647,N_4663);
nor U4885 (N_4885,N_4762,N_4723);
xor U4886 (N_4886,N_4694,N_4639);
or U4887 (N_4887,N_4701,N_4675);
nor U4888 (N_4888,N_4623,N_4797);
and U4889 (N_4889,N_4791,N_4785);
nor U4890 (N_4890,N_4626,N_4744);
nor U4891 (N_4891,N_4681,N_4679);
nor U4892 (N_4892,N_4602,N_4642);
xor U4893 (N_4893,N_4682,N_4621);
and U4894 (N_4894,N_4686,N_4664);
nand U4895 (N_4895,N_4689,N_4793);
or U4896 (N_4896,N_4636,N_4730);
nand U4897 (N_4897,N_4722,N_4781);
xor U4898 (N_4898,N_4674,N_4645);
and U4899 (N_4899,N_4677,N_4746);
xnor U4900 (N_4900,N_4789,N_4730);
or U4901 (N_4901,N_4624,N_4744);
nand U4902 (N_4902,N_4682,N_4656);
nand U4903 (N_4903,N_4780,N_4767);
and U4904 (N_4904,N_4749,N_4784);
nor U4905 (N_4905,N_4771,N_4783);
nand U4906 (N_4906,N_4750,N_4696);
nand U4907 (N_4907,N_4715,N_4689);
or U4908 (N_4908,N_4706,N_4612);
nand U4909 (N_4909,N_4676,N_4701);
xnor U4910 (N_4910,N_4760,N_4647);
or U4911 (N_4911,N_4628,N_4610);
or U4912 (N_4912,N_4616,N_4674);
nand U4913 (N_4913,N_4739,N_4715);
nor U4914 (N_4914,N_4791,N_4617);
nor U4915 (N_4915,N_4633,N_4642);
and U4916 (N_4916,N_4692,N_4786);
xor U4917 (N_4917,N_4700,N_4739);
or U4918 (N_4918,N_4657,N_4702);
xnor U4919 (N_4919,N_4717,N_4678);
nand U4920 (N_4920,N_4710,N_4742);
nor U4921 (N_4921,N_4731,N_4740);
and U4922 (N_4922,N_4752,N_4700);
nand U4923 (N_4923,N_4692,N_4647);
or U4924 (N_4924,N_4767,N_4710);
xor U4925 (N_4925,N_4679,N_4711);
and U4926 (N_4926,N_4620,N_4702);
nand U4927 (N_4927,N_4649,N_4746);
and U4928 (N_4928,N_4631,N_4719);
or U4929 (N_4929,N_4730,N_4751);
nand U4930 (N_4930,N_4690,N_4721);
and U4931 (N_4931,N_4616,N_4693);
xor U4932 (N_4932,N_4634,N_4732);
nand U4933 (N_4933,N_4673,N_4608);
and U4934 (N_4934,N_4770,N_4643);
and U4935 (N_4935,N_4740,N_4780);
nor U4936 (N_4936,N_4742,N_4730);
and U4937 (N_4937,N_4600,N_4797);
nor U4938 (N_4938,N_4676,N_4679);
nor U4939 (N_4939,N_4716,N_4785);
or U4940 (N_4940,N_4745,N_4691);
or U4941 (N_4941,N_4690,N_4747);
or U4942 (N_4942,N_4688,N_4795);
or U4943 (N_4943,N_4652,N_4770);
xor U4944 (N_4944,N_4676,N_4665);
xor U4945 (N_4945,N_4784,N_4657);
xor U4946 (N_4946,N_4602,N_4615);
nor U4947 (N_4947,N_4623,N_4761);
and U4948 (N_4948,N_4789,N_4725);
or U4949 (N_4949,N_4760,N_4660);
nand U4950 (N_4950,N_4684,N_4754);
or U4951 (N_4951,N_4615,N_4773);
or U4952 (N_4952,N_4799,N_4786);
xor U4953 (N_4953,N_4736,N_4779);
nand U4954 (N_4954,N_4779,N_4649);
xor U4955 (N_4955,N_4683,N_4693);
and U4956 (N_4956,N_4662,N_4752);
nor U4957 (N_4957,N_4702,N_4666);
xor U4958 (N_4958,N_4724,N_4760);
nor U4959 (N_4959,N_4785,N_4675);
xnor U4960 (N_4960,N_4777,N_4731);
or U4961 (N_4961,N_4789,N_4734);
or U4962 (N_4962,N_4716,N_4788);
xor U4963 (N_4963,N_4759,N_4687);
or U4964 (N_4964,N_4695,N_4681);
nand U4965 (N_4965,N_4648,N_4743);
or U4966 (N_4966,N_4652,N_4628);
xor U4967 (N_4967,N_4792,N_4673);
and U4968 (N_4968,N_4638,N_4725);
nand U4969 (N_4969,N_4638,N_4718);
nor U4970 (N_4970,N_4693,N_4726);
and U4971 (N_4971,N_4799,N_4735);
nor U4972 (N_4972,N_4647,N_4677);
nor U4973 (N_4973,N_4745,N_4625);
or U4974 (N_4974,N_4652,N_4674);
or U4975 (N_4975,N_4737,N_4794);
xnor U4976 (N_4976,N_4703,N_4614);
and U4977 (N_4977,N_4776,N_4799);
and U4978 (N_4978,N_4760,N_4734);
and U4979 (N_4979,N_4712,N_4642);
nand U4980 (N_4980,N_4753,N_4691);
or U4981 (N_4981,N_4735,N_4655);
and U4982 (N_4982,N_4650,N_4732);
and U4983 (N_4983,N_4767,N_4643);
and U4984 (N_4984,N_4674,N_4753);
and U4985 (N_4985,N_4681,N_4660);
xnor U4986 (N_4986,N_4776,N_4641);
nor U4987 (N_4987,N_4688,N_4621);
and U4988 (N_4988,N_4772,N_4775);
or U4989 (N_4989,N_4621,N_4668);
and U4990 (N_4990,N_4699,N_4771);
xnor U4991 (N_4991,N_4722,N_4791);
or U4992 (N_4992,N_4702,N_4601);
or U4993 (N_4993,N_4704,N_4614);
nand U4994 (N_4994,N_4630,N_4725);
nand U4995 (N_4995,N_4719,N_4701);
or U4996 (N_4996,N_4641,N_4788);
and U4997 (N_4997,N_4773,N_4709);
xor U4998 (N_4998,N_4684,N_4739);
and U4999 (N_4999,N_4765,N_4683);
or UO_0 (O_0,N_4800,N_4855);
nor UO_1 (O_1,N_4985,N_4958);
nand UO_2 (O_2,N_4953,N_4890);
and UO_3 (O_3,N_4825,N_4857);
or UO_4 (O_4,N_4870,N_4836);
and UO_5 (O_5,N_4976,N_4933);
xnor UO_6 (O_6,N_4990,N_4955);
or UO_7 (O_7,N_4871,N_4811);
xnor UO_8 (O_8,N_4878,N_4964);
or UO_9 (O_9,N_4898,N_4819);
nor UO_10 (O_10,N_4813,N_4892);
xor UO_11 (O_11,N_4803,N_4804);
xnor UO_12 (O_12,N_4856,N_4863);
or UO_13 (O_13,N_4928,N_4812);
or UO_14 (O_14,N_4806,N_4815);
nor UO_15 (O_15,N_4910,N_4989);
xor UO_16 (O_16,N_4826,N_4957);
nor UO_17 (O_17,N_4896,N_4822);
nand UO_18 (O_18,N_4943,N_4874);
xnor UO_19 (O_19,N_4846,N_4908);
nand UO_20 (O_20,N_4807,N_4835);
xor UO_21 (O_21,N_4986,N_4901);
xnor UO_22 (O_22,N_4997,N_4948);
nor UO_23 (O_23,N_4903,N_4899);
and UO_24 (O_24,N_4919,N_4994);
and UO_25 (O_25,N_4982,N_4951);
xnor UO_26 (O_26,N_4947,N_4984);
nor UO_27 (O_27,N_4946,N_4916);
xor UO_28 (O_28,N_4991,N_4816);
nor UO_29 (O_29,N_4918,N_4971);
nor UO_30 (O_30,N_4977,N_4817);
and UO_31 (O_31,N_4877,N_4830);
xnor UO_32 (O_32,N_4831,N_4861);
or UO_33 (O_33,N_4875,N_4904);
or UO_34 (O_34,N_4968,N_4956);
or UO_35 (O_35,N_4929,N_4920);
nor UO_36 (O_36,N_4897,N_4954);
xnor UO_37 (O_37,N_4839,N_4970);
or UO_38 (O_38,N_4973,N_4844);
nand UO_39 (O_39,N_4889,N_4848);
nor UO_40 (O_40,N_4880,N_4876);
or UO_41 (O_41,N_4832,N_4895);
nand UO_42 (O_42,N_4998,N_4860);
and UO_43 (O_43,N_4932,N_4814);
or UO_44 (O_44,N_4887,N_4917);
or UO_45 (O_45,N_4926,N_4969);
nor UO_46 (O_46,N_4938,N_4851);
xnor UO_47 (O_47,N_4885,N_4845);
xor UO_48 (O_48,N_4972,N_4801);
and UO_49 (O_49,N_4894,N_4859);
and UO_50 (O_50,N_4905,N_4865);
nand UO_51 (O_51,N_4999,N_4823);
and UO_52 (O_52,N_4967,N_4833);
nor UO_53 (O_53,N_4981,N_4843);
or UO_54 (O_54,N_4867,N_4907);
or UO_55 (O_55,N_4934,N_4940);
nand UO_56 (O_56,N_4808,N_4868);
and UO_57 (O_57,N_4837,N_4939);
nor UO_58 (O_58,N_4834,N_4937);
and UO_59 (O_59,N_4873,N_4941);
or UO_60 (O_60,N_4847,N_4979);
nor UO_61 (O_61,N_4911,N_4931);
nor UO_62 (O_62,N_4974,N_4862);
xnor UO_63 (O_63,N_4914,N_4802);
nor UO_64 (O_64,N_4962,N_4935);
or UO_65 (O_65,N_4820,N_4866);
or UO_66 (O_66,N_4995,N_4952);
nand UO_67 (O_67,N_4882,N_4827);
nor UO_68 (O_68,N_4992,N_4853);
and UO_69 (O_69,N_4944,N_4927);
or UO_70 (O_70,N_4987,N_4821);
and UO_71 (O_71,N_4988,N_4925);
nor UO_72 (O_72,N_4883,N_4913);
and UO_73 (O_73,N_4963,N_4886);
and UO_74 (O_74,N_4945,N_4965);
nor UO_75 (O_75,N_4950,N_4872);
nor UO_76 (O_76,N_4906,N_4915);
nand UO_77 (O_77,N_4852,N_4842);
xor UO_78 (O_78,N_4902,N_4960);
xor UO_79 (O_79,N_4818,N_4912);
and UO_80 (O_80,N_4881,N_4978);
nand UO_81 (O_81,N_4961,N_4921);
xnor UO_82 (O_82,N_4809,N_4923);
and UO_83 (O_83,N_4841,N_4858);
nand UO_84 (O_84,N_4924,N_4942);
nor UO_85 (O_85,N_4909,N_4930);
nand UO_86 (O_86,N_4949,N_4996);
and UO_87 (O_87,N_4840,N_4980);
or UO_88 (O_88,N_4884,N_4810);
xnor UO_89 (O_89,N_4993,N_4922);
nor UO_90 (O_90,N_4879,N_4975);
nor UO_91 (O_91,N_4829,N_4854);
nand UO_92 (O_92,N_4891,N_4864);
nand UO_93 (O_93,N_4936,N_4805);
or UO_94 (O_94,N_4838,N_4893);
nand UO_95 (O_95,N_4966,N_4869);
or UO_96 (O_96,N_4959,N_4983);
and UO_97 (O_97,N_4850,N_4900);
nand UO_98 (O_98,N_4888,N_4849);
xor UO_99 (O_99,N_4828,N_4824);
xor UO_100 (O_100,N_4887,N_4899);
nor UO_101 (O_101,N_4919,N_4833);
nor UO_102 (O_102,N_4877,N_4823);
xnor UO_103 (O_103,N_4878,N_4888);
xor UO_104 (O_104,N_4860,N_4936);
xnor UO_105 (O_105,N_4830,N_4990);
and UO_106 (O_106,N_4930,N_4828);
or UO_107 (O_107,N_4801,N_4955);
nand UO_108 (O_108,N_4805,N_4894);
and UO_109 (O_109,N_4999,N_4883);
nor UO_110 (O_110,N_4908,N_4999);
and UO_111 (O_111,N_4823,N_4838);
or UO_112 (O_112,N_4858,N_4951);
and UO_113 (O_113,N_4845,N_4977);
nand UO_114 (O_114,N_4962,N_4838);
nor UO_115 (O_115,N_4963,N_4951);
and UO_116 (O_116,N_4937,N_4992);
or UO_117 (O_117,N_4844,N_4954);
and UO_118 (O_118,N_4900,N_4987);
xnor UO_119 (O_119,N_4991,N_4948);
xor UO_120 (O_120,N_4835,N_4874);
xnor UO_121 (O_121,N_4989,N_4844);
and UO_122 (O_122,N_4845,N_4808);
and UO_123 (O_123,N_4816,N_4981);
nand UO_124 (O_124,N_4916,N_4811);
nor UO_125 (O_125,N_4840,N_4871);
xnor UO_126 (O_126,N_4876,N_4879);
nand UO_127 (O_127,N_4997,N_4876);
or UO_128 (O_128,N_4951,N_4863);
or UO_129 (O_129,N_4970,N_4866);
and UO_130 (O_130,N_4837,N_4956);
nand UO_131 (O_131,N_4867,N_4852);
xnor UO_132 (O_132,N_4947,N_4882);
or UO_133 (O_133,N_4878,N_4816);
nor UO_134 (O_134,N_4880,N_4993);
and UO_135 (O_135,N_4814,N_4961);
xor UO_136 (O_136,N_4816,N_4955);
or UO_137 (O_137,N_4854,N_4911);
and UO_138 (O_138,N_4983,N_4990);
and UO_139 (O_139,N_4993,N_4918);
nand UO_140 (O_140,N_4961,N_4824);
xor UO_141 (O_141,N_4924,N_4805);
xnor UO_142 (O_142,N_4984,N_4911);
nor UO_143 (O_143,N_4916,N_4931);
and UO_144 (O_144,N_4808,N_4828);
and UO_145 (O_145,N_4869,N_4854);
and UO_146 (O_146,N_4889,N_4832);
and UO_147 (O_147,N_4901,N_4957);
xnor UO_148 (O_148,N_4831,N_4904);
nor UO_149 (O_149,N_4903,N_4968);
nor UO_150 (O_150,N_4973,N_4903);
and UO_151 (O_151,N_4823,N_4831);
or UO_152 (O_152,N_4802,N_4898);
nand UO_153 (O_153,N_4973,N_4884);
nand UO_154 (O_154,N_4802,N_4866);
nand UO_155 (O_155,N_4906,N_4863);
nand UO_156 (O_156,N_4862,N_4938);
nand UO_157 (O_157,N_4818,N_4997);
or UO_158 (O_158,N_4821,N_4894);
xor UO_159 (O_159,N_4923,N_4830);
nand UO_160 (O_160,N_4874,N_4916);
xor UO_161 (O_161,N_4943,N_4956);
nor UO_162 (O_162,N_4902,N_4851);
or UO_163 (O_163,N_4835,N_4802);
or UO_164 (O_164,N_4974,N_4895);
nand UO_165 (O_165,N_4820,N_4892);
or UO_166 (O_166,N_4975,N_4997);
or UO_167 (O_167,N_4849,N_4864);
nor UO_168 (O_168,N_4876,N_4881);
and UO_169 (O_169,N_4971,N_4931);
nand UO_170 (O_170,N_4940,N_4969);
nand UO_171 (O_171,N_4920,N_4917);
xnor UO_172 (O_172,N_4938,N_4929);
and UO_173 (O_173,N_4908,N_4994);
nor UO_174 (O_174,N_4905,N_4837);
nand UO_175 (O_175,N_4893,N_4907);
and UO_176 (O_176,N_4949,N_4896);
xor UO_177 (O_177,N_4845,N_4838);
or UO_178 (O_178,N_4805,N_4947);
and UO_179 (O_179,N_4814,N_4984);
nor UO_180 (O_180,N_4940,N_4891);
nor UO_181 (O_181,N_4866,N_4922);
and UO_182 (O_182,N_4850,N_4905);
nor UO_183 (O_183,N_4834,N_4956);
nor UO_184 (O_184,N_4979,N_4993);
xor UO_185 (O_185,N_4826,N_4822);
and UO_186 (O_186,N_4913,N_4905);
or UO_187 (O_187,N_4988,N_4896);
and UO_188 (O_188,N_4914,N_4962);
and UO_189 (O_189,N_4887,N_4813);
nor UO_190 (O_190,N_4922,N_4843);
nor UO_191 (O_191,N_4828,N_4862);
nor UO_192 (O_192,N_4857,N_4867);
nor UO_193 (O_193,N_4803,N_4818);
and UO_194 (O_194,N_4892,N_4877);
or UO_195 (O_195,N_4841,N_4975);
nor UO_196 (O_196,N_4871,N_4972);
xor UO_197 (O_197,N_4858,N_4954);
nor UO_198 (O_198,N_4973,N_4830);
or UO_199 (O_199,N_4975,N_4877);
xnor UO_200 (O_200,N_4996,N_4821);
or UO_201 (O_201,N_4956,N_4858);
nor UO_202 (O_202,N_4843,N_4812);
or UO_203 (O_203,N_4929,N_4937);
or UO_204 (O_204,N_4920,N_4851);
nand UO_205 (O_205,N_4936,N_4930);
or UO_206 (O_206,N_4811,N_4867);
and UO_207 (O_207,N_4827,N_4822);
or UO_208 (O_208,N_4909,N_4960);
nand UO_209 (O_209,N_4871,N_4803);
nand UO_210 (O_210,N_4883,N_4893);
nor UO_211 (O_211,N_4823,N_4947);
or UO_212 (O_212,N_4934,N_4952);
nand UO_213 (O_213,N_4930,N_4906);
xor UO_214 (O_214,N_4942,N_4870);
and UO_215 (O_215,N_4904,N_4859);
nor UO_216 (O_216,N_4861,N_4912);
and UO_217 (O_217,N_4995,N_4815);
and UO_218 (O_218,N_4869,N_4956);
nand UO_219 (O_219,N_4817,N_4921);
and UO_220 (O_220,N_4833,N_4882);
nand UO_221 (O_221,N_4894,N_4888);
xor UO_222 (O_222,N_4909,N_4810);
or UO_223 (O_223,N_4814,N_4916);
or UO_224 (O_224,N_4941,N_4847);
nor UO_225 (O_225,N_4974,N_4934);
and UO_226 (O_226,N_4814,N_4911);
and UO_227 (O_227,N_4810,N_4982);
nand UO_228 (O_228,N_4997,N_4842);
nand UO_229 (O_229,N_4843,N_4996);
or UO_230 (O_230,N_4827,N_4902);
nand UO_231 (O_231,N_4953,N_4990);
nor UO_232 (O_232,N_4845,N_4933);
xnor UO_233 (O_233,N_4902,N_4964);
xnor UO_234 (O_234,N_4836,N_4835);
xnor UO_235 (O_235,N_4950,N_4873);
xor UO_236 (O_236,N_4837,N_4810);
nand UO_237 (O_237,N_4973,N_4927);
and UO_238 (O_238,N_4872,N_4862);
nand UO_239 (O_239,N_4949,N_4891);
xor UO_240 (O_240,N_4909,N_4873);
nand UO_241 (O_241,N_4960,N_4923);
nor UO_242 (O_242,N_4983,N_4914);
xor UO_243 (O_243,N_4840,N_4862);
xnor UO_244 (O_244,N_4913,N_4869);
nor UO_245 (O_245,N_4963,N_4869);
and UO_246 (O_246,N_4998,N_4912);
or UO_247 (O_247,N_4815,N_4970);
nor UO_248 (O_248,N_4998,N_4929);
nor UO_249 (O_249,N_4915,N_4925);
xor UO_250 (O_250,N_4845,N_4824);
and UO_251 (O_251,N_4977,N_4896);
nor UO_252 (O_252,N_4866,N_4999);
and UO_253 (O_253,N_4956,N_4931);
xor UO_254 (O_254,N_4863,N_4919);
and UO_255 (O_255,N_4881,N_4941);
nor UO_256 (O_256,N_4987,N_4928);
nand UO_257 (O_257,N_4850,N_4841);
nor UO_258 (O_258,N_4946,N_4872);
and UO_259 (O_259,N_4907,N_4946);
nand UO_260 (O_260,N_4963,N_4971);
or UO_261 (O_261,N_4950,N_4805);
xor UO_262 (O_262,N_4872,N_4987);
nand UO_263 (O_263,N_4874,N_4926);
xnor UO_264 (O_264,N_4892,N_4810);
nand UO_265 (O_265,N_4967,N_4870);
nand UO_266 (O_266,N_4806,N_4899);
nand UO_267 (O_267,N_4993,N_4832);
or UO_268 (O_268,N_4834,N_4969);
nor UO_269 (O_269,N_4968,N_4872);
xor UO_270 (O_270,N_4838,N_4932);
xor UO_271 (O_271,N_4868,N_4867);
or UO_272 (O_272,N_4892,N_4916);
nand UO_273 (O_273,N_4995,N_4900);
xor UO_274 (O_274,N_4939,N_4863);
nand UO_275 (O_275,N_4812,N_4883);
or UO_276 (O_276,N_4845,N_4937);
xor UO_277 (O_277,N_4916,N_4971);
nor UO_278 (O_278,N_4964,N_4894);
or UO_279 (O_279,N_4845,N_4926);
or UO_280 (O_280,N_4819,N_4822);
and UO_281 (O_281,N_4983,N_4803);
xor UO_282 (O_282,N_4983,N_4986);
xnor UO_283 (O_283,N_4936,N_4919);
nand UO_284 (O_284,N_4892,N_4969);
nor UO_285 (O_285,N_4927,N_4960);
xnor UO_286 (O_286,N_4881,N_4801);
nor UO_287 (O_287,N_4889,N_4981);
xor UO_288 (O_288,N_4985,N_4876);
xor UO_289 (O_289,N_4895,N_4901);
nand UO_290 (O_290,N_4880,N_4944);
xnor UO_291 (O_291,N_4974,N_4936);
nor UO_292 (O_292,N_4844,N_4978);
or UO_293 (O_293,N_4988,N_4943);
xnor UO_294 (O_294,N_4866,N_4875);
xnor UO_295 (O_295,N_4912,N_4960);
nor UO_296 (O_296,N_4841,N_4834);
nand UO_297 (O_297,N_4818,N_4978);
nor UO_298 (O_298,N_4857,N_4813);
nand UO_299 (O_299,N_4867,N_4893);
or UO_300 (O_300,N_4901,N_4937);
and UO_301 (O_301,N_4924,N_4824);
nand UO_302 (O_302,N_4914,N_4853);
or UO_303 (O_303,N_4877,N_4900);
or UO_304 (O_304,N_4990,N_4861);
nor UO_305 (O_305,N_4929,N_4926);
and UO_306 (O_306,N_4829,N_4938);
nand UO_307 (O_307,N_4805,N_4847);
nand UO_308 (O_308,N_4856,N_4841);
nor UO_309 (O_309,N_4874,N_4948);
or UO_310 (O_310,N_4947,N_4969);
and UO_311 (O_311,N_4903,N_4838);
nand UO_312 (O_312,N_4937,N_4951);
nand UO_313 (O_313,N_4973,N_4891);
or UO_314 (O_314,N_4857,N_4864);
nor UO_315 (O_315,N_4944,N_4872);
nand UO_316 (O_316,N_4917,N_4861);
and UO_317 (O_317,N_4932,N_4983);
nand UO_318 (O_318,N_4810,N_4819);
nand UO_319 (O_319,N_4947,N_4977);
nand UO_320 (O_320,N_4903,N_4900);
nor UO_321 (O_321,N_4972,N_4886);
xnor UO_322 (O_322,N_4920,N_4826);
nor UO_323 (O_323,N_4808,N_4802);
xor UO_324 (O_324,N_4871,N_4942);
and UO_325 (O_325,N_4800,N_4968);
nor UO_326 (O_326,N_4821,N_4924);
or UO_327 (O_327,N_4910,N_4946);
nor UO_328 (O_328,N_4944,N_4982);
and UO_329 (O_329,N_4981,N_4836);
xnor UO_330 (O_330,N_4815,N_4902);
nor UO_331 (O_331,N_4818,N_4910);
and UO_332 (O_332,N_4870,N_4895);
or UO_333 (O_333,N_4987,N_4801);
xnor UO_334 (O_334,N_4869,N_4948);
or UO_335 (O_335,N_4908,N_4888);
nand UO_336 (O_336,N_4838,N_4901);
or UO_337 (O_337,N_4889,N_4846);
or UO_338 (O_338,N_4809,N_4950);
xor UO_339 (O_339,N_4926,N_4925);
xor UO_340 (O_340,N_4992,N_4846);
nor UO_341 (O_341,N_4977,N_4914);
nor UO_342 (O_342,N_4893,N_4979);
nand UO_343 (O_343,N_4988,N_4830);
nor UO_344 (O_344,N_4835,N_4996);
or UO_345 (O_345,N_4810,N_4828);
nand UO_346 (O_346,N_4839,N_4946);
xor UO_347 (O_347,N_4966,N_4831);
or UO_348 (O_348,N_4983,N_4957);
nand UO_349 (O_349,N_4950,N_4947);
or UO_350 (O_350,N_4893,N_4937);
nor UO_351 (O_351,N_4927,N_4932);
and UO_352 (O_352,N_4803,N_4812);
nor UO_353 (O_353,N_4828,N_4873);
xor UO_354 (O_354,N_4827,N_4970);
nand UO_355 (O_355,N_4849,N_4959);
or UO_356 (O_356,N_4951,N_4902);
nor UO_357 (O_357,N_4880,N_4951);
and UO_358 (O_358,N_4964,N_4821);
and UO_359 (O_359,N_4959,N_4874);
nor UO_360 (O_360,N_4987,N_4947);
nor UO_361 (O_361,N_4817,N_4910);
and UO_362 (O_362,N_4816,N_4903);
xnor UO_363 (O_363,N_4825,N_4833);
nor UO_364 (O_364,N_4935,N_4944);
and UO_365 (O_365,N_4947,N_4836);
nand UO_366 (O_366,N_4968,N_4885);
and UO_367 (O_367,N_4985,N_4954);
and UO_368 (O_368,N_4884,N_4900);
or UO_369 (O_369,N_4831,N_4803);
and UO_370 (O_370,N_4991,N_4838);
and UO_371 (O_371,N_4854,N_4881);
nand UO_372 (O_372,N_4902,N_4836);
or UO_373 (O_373,N_4956,N_4812);
xnor UO_374 (O_374,N_4822,N_4977);
or UO_375 (O_375,N_4897,N_4857);
and UO_376 (O_376,N_4979,N_4917);
or UO_377 (O_377,N_4893,N_4863);
and UO_378 (O_378,N_4970,N_4998);
nor UO_379 (O_379,N_4807,N_4892);
xor UO_380 (O_380,N_4888,N_4825);
and UO_381 (O_381,N_4982,N_4805);
nand UO_382 (O_382,N_4974,N_4823);
xnor UO_383 (O_383,N_4920,N_4896);
and UO_384 (O_384,N_4959,N_4907);
nand UO_385 (O_385,N_4988,N_4891);
and UO_386 (O_386,N_4924,N_4888);
and UO_387 (O_387,N_4862,N_4845);
xor UO_388 (O_388,N_4886,N_4804);
or UO_389 (O_389,N_4910,N_4838);
xor UO_390 (O_390,N_4859,N_4819);
xnor UO_391 (O_391,N_4828,N_4843);
xnor UO_392 (O_392,N_4901,N_4922);
or UO_393 (O_393,N_4946,N_4804);
or UO_394 (O_394,N_4919,N_4853);
nor UO_395 (O_395,N_4846,N_4951);
nor UO_396 (O_396,N_4993,N_4932);
and UO_397 (O_397,N_4971,N_4838);
xor UO_398 (O_398,N_4902,N_4965);
nor UO_399 (O_399,N_4810,N_4871);
or UO_400 (O_400,N_4870,N_4915);
and UO_401 (O_401,N_4935,N_4991);
or UO_402 (O_402,N_4950,N_4875);
or UO_403 (O_403,N_4865,N_4838);
nor UO_404 (O_404,N_4916,N_4966);
and UO_405 (O_405,N_4926,N_4914);
or UO_406 (O_406,N_4801,N_4845);
and UO_407 (O_407,N_4962,N_4846);
or UO_408 (O_408,N_4867,N_4846);
xnor UO_409 (O_409,N_4800,N_4961);
nand UO_410 (O_410,N_4963,N_4950);
nor UO_411 (O_411,N_4907,N_4990);
and UO_412 (O_412,N_4909,N_4885);
or UO_413 (O_413,N_4932,N_4893);
nor UO_414 (O_414,N_4955,N_4831);
xnor UO_415 (O_415,N_4822,N_4805);
nand UO_416 (O_416,N_4957,N_4852);
xnor UO_417 (O_417,N_4928,N_4849);
and UO_418 (O_418,N_4925,N_4812);
or UO_419 (O_419,N_4871,N_4843);
nor UO_420 (O_420,N_4982,N_4857);
nor UO_421 (O_421,N_4993,N_4895);
xnor UO_422 (O_422,N_4896,N_4995);
nor UO_423 (O_423,N_4978,N_4973);
nand UO_424 (O_424,N_4899,N_4968);
xor UO_425 (O_425,N_4937,N_4892);
and UO_426 (O_426,N_4923,N_4840);
and UO_427 (O_427,N_4928,N_4872);
nor UO_428 (O_428,N_4963,N_4871);
xor UO_429 (O_429,N_4998,N_4868);
or UO_430 (O_430,N_4913,N_4977);
nor UO_431 (O_431,N_4999,N_4975);
nand UO_432 (O_432,N_4954,N_4833);
xor UO_433 (O_433,N_4984,N_4800);
xnor UO_434 (O_434,N_4844,N_4800);
or UO_435 (O_435,N_4846,N_4946);
xnor UO_436 (O_436,N_4927,N_4983);
nor UO_437 (O_437,N_4995,N_4808);
or UO_438 (O_438,N_4933,N_4871);
or UO_439 (O_439,N_4931,N_4941);
and UO_440 (O_440,N_4970,N_4973);
xor UO_441 (O_441,N_4855,N_4839);
nand UO_442 (O_442,N_4823,N_4933);
and UO_443 (O_443,N_4896,N_4843);
nor UO_444 (O_444,N_4880,N_4961);
xnor UO_445 (O_445,N_4927,N_4836);
nor UO_446 (O_446,N_4929,N_4984);
and UO_447 (O_447,N_4841,N_4905);
nand UO_448 (O_448,N_4982,N_4816);
nor UO_449 (O_449,N_4975,N_4820);
nand UO_450 (O_450,N_4911,N_4891);
or UO_451 (O_451,N_4902,N_4901);
and UO_452 (O_452,N_4904,N_4960);
nor UO_453 (O_453,N_4836,N_4871);
nand UO_454 (O_454,N_4923,N_4943);
xor UO_455 (O_455,N_4959,N_4911);
nand UO_456 (O_456,N_4844,N_4956);
or UO_457 (O_457,N_4966,N_4866);
and UO_458 (O_458,N_4827,N_4836);
and UO_459 (O_459,N_4906,N_4841);
xnor UO_460 (O_460,N_4838,N_4905);
nor UO_461 (O_461,N_4820,N_4985);
xor UO_462 (O_462,N_4847,N_4945);
and UO_463 (O_463,N_4919,N_4838);
nand UO_464 (O_464,N_4849,N_4858);
xnor UO_465 (O_465,N_4967,N_4995);
or UO_466 (O_466,N_4820,N_4898);
or UO_467 (O_467,N_4963,N_4968);
or UO_468 (O_468,N_4900,N_4983);
xnor UO_469 (O_469,N_4958,N_4817);
nor UO_470 (O_470,N_4860,N_4929);
and UO_471 (O_471,N_4828,N_4870);
xnor UO_472 (O_472,N_4826,N_4989);
xnor UO_473 (O_473,N_4865,N_4813);
or UO_474 (O_474,N_4856,N_4966);
and UO_475 (O_475,N_4903,N_4948);
and UO_476 (O_476,N_4912,N_4927);
or UO_477 (O_477,N_4916,N_4960);
nand UO_478 (O_478,N_4826,N_4927);
nand UO_479 (O_479,N_4820,N_4930);
or UO_480 (O_480,N_4900,N_4901);
or UO_481 (O_481,N_4939,N_4989);
nor UO_482 (O_482,N_4891,N_4933);
and UO_483 (O_483,N_4914,N_4894);
nor UO_484 (O_484,N_4808,N_4981);
and UO_485 (O_485,N_4849,N_4876);
nand UO_486 (O_486,N_4894,N_4827);
nor UO_487 (O_487,N_4801,N_4981);
or UO_488 (O_488,N_4964,N_4965);
nor UO_489 (O_489,N_4976,N_4833);
xor UO_490 (O_490,N_4983,N_4979);
or UO_491 (O_491,N_4801,N_4816);
nor UO_492 (O_492,N_4874,N_4831);
or UO_493 (O_493,N_4844,N_4889);
xnor UO_494 (O_494,N_4808,N_4877);
and UO_495 (O_495,N_4901,N_4949);
xor UO_496 (O_496,N_4800,N_4975);
or UO_497 (O_497,N_4948,N_4872);
xnor UO_498 (O_498,N_4927,N_4883);
xor UO_499 (O_499,N_4996,N_4887);
nand UO_500 (O_500,N_4876,N_4906);
nor UO_501 (O_501,N_4967,N_4897);
and UO_502 (O_502,N_4847,N_4970);
nor UO_503 (O_503,N_4966,N_4873);
or UO_504 (O_504,N_4828,N_4952);
and UO_505 (O_505,N_4826,N_4847);
nand UO_506 (O_506,N_4806,N_4891);
and UO_507 (O_507,N_4846,N_4973);
xor UO_508 (O_508,N_4922,N_4999);
or UO_509 (O_509,N_4906,N_4956);
or UO_510 (O_510,N_4826,N_4869);
nand UO_511 (O_511,N_4802,N_4833);
xor UO_512 (O_512,N_4924,N_4827);
nor UO_513 (O_513,N_4953,N_4954);
and UO_514 (O_514,N_4808,N_4895);
nand UO_515 (O_515,N_4981,N_4925);
nor UO_516 (O_516,N_4903,N_4828);
or UO_517 (O_517,N_4870,N_4939);
nor UO_518 (O_518,N_4801,N_4950);
and UO_519 (O_519,N_4998,N_4898);
and UO_520 (O_520,N_4846,N_4898);
or UO_521 (O_521,N_4985,N_4978);
and UO_522 (O_522,N_4973,N_4816);
xor UO_523 (O_523,N_4943,N_4876);
xnor UO_524 (O_524,N_4899,N_4812);
nand UO_525 (O_525,N_4825,N_4904);
nand UO_526 (O_526,N_4811,N_4983);
xor UO_527 (O_527,N_4913,N_4940);
or UO_528 (O_528,N_4823,N_4994);
nor UO_529 (O_529,N_4825,N_4896);
xnor UO_530 (O_530,N_4958,N_4879);
xnor UO_531 (O_531,N_4924,N_4965);
and UO_532 (O_532,N_4963,N_4936);
nand UO_533 (O_533,N_4952,N_4876);
or UO_534 (O_534,N_4940,N_4880);
or UO_535 (O_535,N_4998,N_4987);
nand UO_536 (O_536,N_4938,N_4947);
nand UO_537 (O_537,N_4991,N_4868);
xor UO_538 (O_538,N_4938,N_4839);
xnor UO_539 (O_539,N_4918,N_4999);
nor UO_540 (O_540,N_4891,N_4827);
nor UO_541 (O_541,N_4818,N_4961);
and UO_542 (O_542,N_4814,N_4888);
nand UO_543 (O_543,N_4966,N_4890);
nor UO_544 (O_544,N_4884,N_4941);
or UO_545 (O_545,N_4897,N_4883);
or UO_546 (O_546,N_4999,N_4942);
nor UO_547 (O_547,N_4836,N_4849);
or UO_548 (O_548,N_4884,N_4897);
or UO_549 (O_549,N_4900,N_4852);
and UO_550 (O_550,N_4895,N_4842);
xor UO_551 (O_551,N_4962,N_4858);
or UO_552 (O_552,N_4913,N_4861);
or UO_553 (O_553,N_4948,N_4839);
xor UO_554 (O_554,N_4907,N_4844);
nand UO_555 (O_555,N_4887,N_4911);
or UO_556 (O_556,N_4916,N_4887);
or UO_557 (O_557,N_4939,N_4971);
or UO_558 (O_558,N_4828,N_4888);
nand UO_559 (O_559,N_4970,N_4840);
and UO_560 (O_560,N_4919,N_4882);
nand UO_561 (O_561,N_4899,N_4997);
and UO_562 (O_562,N_4962,N_4997);
xnor UO_563 (O_563,N_4994,N_4998);
nor UO_564 (O_564,N_4832,N_4821);
nand UO_565 (O_565,N_4815,N_4978);
or UO_566 (O_566,N_4895,N_4891);
or UO_567 (O_567,N_4820,N_4814);
and UO_568 (O_568,N_4956,N_4828);
xor UO_569 (O_569,N_4905,N_4842);
nor UO_570 (O_570,N_4951,N_4916);
xor UO_571 (O_571,N_4833,N_4812);
xor UO_572 (O_572,N_4914,N_4960);
or UO_573 (O_573,N_4954,N_4878);
and UO_574 (O_574,N_4899,N_4873);
or UO_575 (O_575,N_4879,N_4829);
nand UO_576 (O_576,N_4949,N_4974);
nor UO_577 (O_577,N_4963,N_4911);
nand UO_578 (O_578,N_4839,N_4851);
nor UO_579 (O_579,N_4987,N_4879);
or UO_580 (O_580,N_4953,N_4874);
xnor UO_581 (O_581,N_4994,N_4819);
or UO_582 (O_582,N_4815,N_4886);
and UO_583 (O_583,N_4948,N_4868);
or UO_584 (O_584,N_4961,N_4933);
or UO_585 (O_585,N_4995,N_4821);
and UO_586 (O_586,N_4850,N_4990);
nand UO_587 (O_587,N_4907,N_4950);
nand UO_588 (O_588,N_4963,N_4825);
and UO_589 (O_589,N_4920,N_4844);
xor UO_590 (O_590,N_4913,N_4896);
nor UO_591 (O_591,N_4817,N_4843);
nand UO_592 (O_592,N_4810,N_4926);
nand UO_593 (O_593,N_4998,N_4984);
nor UO_594 (O_594,N_4845,N_4966);
nand UO_595 (O_595,N_4983,N_4903);
nor UO_596 (O_596,N_4985,N_4924);
and UO_597 (O_597,N_4951,N_4921);
xor UO_598 (O_598,N_4828,N_4960);
or UO_599 (O_599,N_4926,N_4974);
or UO_600 (O_600,N_4895,N_4821);
nand UO_601 (O_601,N_4954,N_4960);
nand UO_602 (O_602,N_4839,N_4950);
xor UO_603 (O_603,N_4991,N_4849);
or UO_604 (O_604,N_4956,N_4919);
or UO_605 (O_605,N_4922,N_4884);
nor UO_606 (O_606,N_4880,N_4905);
nor UO_607 (O_607,N_4926,N_4932);
xnor UO_608 (O_608,N_4894,N_4963);
nand UO_609 (O_609,N_4998,N_4801);
nor UO_610 (O_610,N_4844,N_4936);
nor UO_611 (O_611,N_4890,N_4822);
and UO_612 (O_612,N_4973,N_4980);
nor UO_613 (O_613,N_4963,N_4829);
or UO_614 (O_614,N_4934,N_4860);
and UO_615 (O_615,N_4808,N_4876);
or UO_616 (O_616,N_4918,N_4991);
nor UO_617 (O_617,N_4947,N_4801);
and UO_618 (O_618,N_4813,N_4920);
and UO_619 (O_619,N_4926,N_4904);
xor UO_620 (O_620,N_4811,N_4831);
nand UO_621 (O_621,N_4832,N_4991);
and UO_622 (O_622,N_4959,N_4880);
nor UO_623 (O_623,N_4946,N_4860);
nand UO_624 (O_624,N_4804,N_4916);
and UO_625 (O_625,N_4861,N_4875);
or UO_626 (O_626,N_4964,N_4837);
and UO_627 (O_627,N_4942,N_4963);
nor UO_628 (O_628,N_4943,N_4895);
nand UO_629 (O_629,N_4954,N_4921);
or UO_630 (O_630,N_4815,N_4901);
xnor UO_631 (O_631,N_4988,N_4948);
xor UO_632 (O_632,N_4941,N_4962);
and UO_633 (O_633,N_4923,N_4833);
nor UO_634 (O_634,N_4934,N_4806);
nor UO_635 (O_635,N_4905,N_4991);
and UO_636 (O_636,N_4873,N_4818);
or UO_637 (O_637,N_4975,N_4804);
nor UO_638 (O_638,N_4814,N_4818);
nand UO_639 (O_639,N_4890,N_4871);
nor UO_640 (O_640,N_4900,N_4811);
nor UO_641 (O_641,N_4864,N_4940);
nor UO_642 (O_642,N_4860,N_4809);
nand UO_643 (O_643,N_4884,N_4803);
and UO_644 (O_644,N_4968,N_4938);
nor UO_645 (O_645,N_4812,N_4907);
and UO_646 (O_646,N_4917,N_4873);
or UO_647 (O_647,N_4922,N_4965);
and UO_648 (O_648,N_4810,N_4941);
nor UO_649 (O_649,N_4868,N_4904);
nand UO_650 (O_650,N_4954,N_4855);
nor UO_651 (O_651,N_4942,N_4906);
xnor UO_652 (O_652,N_4905,N_4846);
or UO_653 (O_653,N_4872,N_4924);
nor UO_654 (O_654,N_4911,N_4872);
nand UO_655 (O_655,N_4961,N_4902);
nor UO_656 (O_656,N_4985,N_4909);
xnor UO_657 (O_657,N_4894,N_4813);
or UO_658 (O_658,N_4804,N_4885);
and UO_659 (O_659,N_4802,N_4969);
and UO_660 (O_660,N_4873,N_4959);
nand UO_661 (O_661,N_4916,N_4881);
nor UO_662 (O_662,N_4946,N_4958);
and UO_663 (O_663,N_4850,N_4833);
and UO_664 (O_664,N_4992,N_4807);
nor UO_665 (O_665,N_4888,N_4889);
nand UO_666 (O_666,N_4974,N_4800);
or UO_667 (O_667,N_4993,N_4994);
or UO_668 (O_668,N_4907,N_4960);
nand UO_669 (O_669,N_4974,N_4929);
nor UO_670 (O_670,N_4951,N_4914);
or UO_671 (O_671,N_4802,N_4801);
or UO_672 (O_672,N_4805,N_4983);
xnor UO_673 (O_673,N_4944,N_4920);
nor UO_674 (O_674,N_4851,N_4829);
xnor UO_675 (O_675,N_4935,N_4833);
nor UO_676 (O_676,N_4848,N_4994);
nor UO_677 (O_677,N_4959,N_4871);
nor UO_678 (O_678,N_4806,N_4804);
nand UO_679 (O_679,N_4880,N_4969);
nor UO_680 (O_680,N_4948,N_4863);
or UO_681 (O_681,N_4933,N_4985);
and UO_682 (O_682,N_4888,N_4906);
nor UO_683 (O_683,N_4982,N_4952);
nand UO_684 (O_684,N_4985,N_4926);
and UO_685 (O_685,N_4904,N_4915);
or UO_686 (O_686,N_4806,N_4937);
nor UO_687 (O_687,N_4807,N_4913);
or UO_688 (O_688,N_4937,N_4805);
and UO_689 (O_689,N_4964,N_4814);
nor UO_690 (O_690,N_4928,N_4903);
nor UO_691 (O_691,N_4977,N_4910);
nand UO_692 (O_692,N_4864,N_4905);
and UO_693 (O_693,N_4825,N_4848);
or UO_694 (O_694,N_4878,N_4915);
nor UO_695 (O_695,N_4959,N_4841);
xor UO_696 (O_696,N_4933,N_4901);
xor UO_697 (O_697,N_4833,N_4952);
nand UO_698 (O_698,N_4969,N_4954);
or UO_699 (O_699,N_4900,N_4813);
xor UO_700 (O_700,N_4911,N_4943);
xnor UO_701 (O_701,N_4933,N_4941);
nand UO_702 (O_702,N_4800,N_4834);
nand UO_703 (O_703,N_4953,N_4808);
nand UO_704 (O_704,N_4833,N_4804);
or UO_705 (O_705,N_4819,N_4856);
and UO_706 (O_706,N_4983,N_4958);
or UO_707 (O_707,N_4843,N_4957);
or UO_708 (O_708,N_4810,N_4984);
xnor UO_709 (O_709,N_4874,N_4951);
or UO_710 (O_710,N_4801,N_4889);
and UO_711 (O_711,N_4912,N_4991);
or UO_712 (O_712,N_4894,N_4949);
or UO_713 (O_713,N_4890,N_4977);
nor UO_714 (O_714,N_4907,N_4900);
or UO_715 (O_715,N_4921,N_4915);
nor UO_716 (O_716,N_4857,N_4972);
or UO_717 (O_717,N_4931,N_4979);
xnor UO_718 (O_718,N_4877,N_4984);
or UO_719 (O_719,N_4964,N_4833);
nor UO_720 (O_720,N_4992,N_4850);
nand UO_721 (O_721,N_4812,N_4875);
nand UO_722 (O_722,N_4899,N_4975);
nor UO_723 (O_723,N_4951,N_4820);
nand UO_724 (O_724,N_4864,N_4914);
xnor UO_725 (O_725,N_4818,N_4945);
nor UO_726 (O_726,N_4883,N_4898);
or UO_727 (O_727,N_4920,N_4940);
nand UO_728 (O_728,N_4922,N_4989);
nand UO_729 (O_729,N_4995,N_4992);
xnor UO_730 (O_730,N_4984,N_4969);
xor UO_731 (O_731,N_4926,N_4862);
nor UO_732 (O_732,N_4840,N_4886);
nor UO_733 (O_733,N_4950,N_4818);
nor UO_734 (O_734,N_4835,N_4869);
nand UO_735 (O_735,N_4899,N_4995);
nand UO_736 (O_736,N_4989,N_4934);
and UO_737 (O_737,N_4944,N_4916);
or UO_738 (O_738,N_4978,N_4837);
or UO_739 (O_739,N_4957,N_4927);
nor UO_740 (O_740,N_4895,N_4816);
and UO_741 (O_741,N_4934,N_4887);
nor UO_742 (O_742,N_4877,N_4908);
and UO_743 (O_743,N_4830,N_4947);
nor UO_744 (O_744,N_4913,N_4832);
and UO_745 (O_745,N_4853,N_4873);
nor UO_746 (O_746,N_4856,N_4846);
or UO_747 (O_747,N_4953,N_4888);
or UO_748 (O_748,N_4884,N_4886);
xnor UO_749 (O_749,N_4887,N_4940);
or UO_750 (O_750,N_4967,N_4993);
nand UO_751 (O_751,N_4808,N_4958);
xnor UO_752 (O_752,N_4815,N_4887);
nand UO_753 (O_753,N_4897,N_4997);
and UO_754 (O_754,N_4883,N_4830);
nand UO_755 (O_755,N_4993,N_4920);
or UO_756 (O_756,N_4906,N_4925);
and UO_757 (O_757,N_4880,N_4813);
nor UO_758 (O_758,N_4906,N_4978);
or UO_759 (O_759,N_4997,N_4894);
and UO_760 (O_760,N_4947,N_4852);
xnor UO_761 (O_761,N_4936,N_4889);
nand UO_762 (O_762,N_4888,N_4833);
or UO_763 (O_763,N_4856,N_4920);
and UO_764 (O_764,N_4988,N_4916);
nor UO_765 (O_765,N_4921,N_4850);
and UO_766 (O_766,N_4815,N_4954);
xnor UO_767 (O_767,N_4841,N_4810);
nand UO_768 (O_768,N_4982,N_4853);
xnor UO_769 (O_769,N_4970,N_4863);
and UO_770 (O_770,N_4961,N_4898);
nor UO_771 (O_771,N_4896,N_4827);
nor UO_772 (O_772,N_4801,N_4924);
nand UO_773 (O_773,N_4908,N_4836);
nand UO_774 (O_774,N_4935,N_4943);
xor UO_775 (O_775,N_4971,N_4874);
or UO_776 (O_776,N_4989,N_4974);
or UO_777 (O_777,N_4806,N_4938);
or UO_778 (O_778,N_4934,N_4878);
nor UO_779 (O_779,N_4962,N_4835);
xor UO_780 (O_780,N_4973,N_4958);
and UO_781 (O_781,N_4862,N_4899);
nand UO_782 (O_782,N_4963,N_4975);
or UO_783 (O_783,N_4924,N_4819);
xor UO_784 (O_784,N_4938,N_4982);
nor UO_785 (O_785,N_4854,N_4989);
nand UO_786 (O_786,N_4862,N_4950);
nor UO_787 (O_787,N_4974,N_4918);
nand UO_788 (O_788,N_4904,N_4869);
and UO_789 (O_789,N_4969,N_4993);
nand UO_790 (O_790,N_4866,N_4838);
nor UO_791 (O_791,N_4943,N_4886);
nor UO_792 (O_792,N_4895,N_4828);
nand UO_793 (O_793,N_4873,N_4944);
nand UO_794 (O_794,N_4815,N_4859);
nor UO_795 (O_795,N_4894,N_4916);
or UO_796 (O_796,N_4829,N_4868);
nor UO_797 (O_797,N_4853,N_4975);
or UO_798 (O_798,N_4871,N_4892);
and UO_799 (O_799,N_4872,N_4934);
nand UO_800 (O_800,N_4960,N_4870);
and UO_801 (O_801,N_4880,N_4985);
and UO_802 (O_802,N_4833,N_4931);
and UO_803 (O_803,N_4892,N_4906);
xnor UO_804 (O_804,N_4893,N_4927);
and UO_805 (O_805,N_4872,N_4937);
or UO_806 (O_806,N_4880,N_4971);
nor UO_807 (O_807,N_4891,N_4915);
nand UO_808 (O_808,N_4810,N_4961);
and UO_809 (O_809,N_4810,N_4867);
or UO_810 (O_810,N_4863,N_4935);
nand UO_811 (O_811,N_4849,N_4810);
nand UO_812 (O_812,N_4966,N_4885);
xor UO_813 (O_813,N_4873,N_4875);
nand UO_814 (O_814,N_4850,N_4861);
and UO_815 (O_815,N_4811,N_4837);
xnor UO_816 (O_816,N_4878,N_4921);
nor UO_817 (O_817,N_4820,N_4914);
or UO_818 (O_818,N_4829,N_4945);
xor UO_819 (O_819,N_4911,N_4940);
xor UO_820 (O_820,N_4823,N_4926);
nor UO_821 (O_821,N_4925,N_4972);
xor UO_822 (O_822,N_4805,N_4838);
nand UO_823 (O_823,N_4965,N_4876);
or UO_824 (O_824,N_4842,N_4961);
nand UO_825 (O_825,N_4964,N_4983);
or UO_826 (O_826,N_4837,N_4989);
and UO_827 (O_827,N_4980,N_4820);
or UO_828 (O_828,N_4977,N_4818);
nand UO_829 (O_829,N_4969,N_4858);
or UO_830 (O_830,N_4982,N_4813);
nand UO_831 (O_831,N_4982,N_4871);
and UO_832 (O_832,N_4853,N_4875);
nor UO_833 (O_833,N_4826,N_4930);
or UO_834 (O_834,N_4841,N_4955);
xnor UO_835 (O_835,N_4849,N_4985);
nor UO_836 (O_836,N_4913,N_4955);
or UO_837 (O_837,N_4939,N_4943);
nor UO_838 (O_838,N_4987,N_4855);
nor UO_839 (O_839,N_4894,N_4961);
and UO_840 (O_840,N_4838,N_4987);
nand UO_841 (O_841,N_4890,N_4800);
xor UO_842 (O_842,N_4986,N_4803);
nand UO_843 (O_843,N_4808,N_4804);
or UO_844 (O_844,N_4914,N_4996);
nor UO_845 (O_845,N_4928,N_4950);
nand UO_846 (O_846,N_4804,N_4964);
nor UO_847 (O_847,N_4833,N_4912);
nor UO_848 (O_848,N_4842,N_4998);
and UO_849 (O_849,N_4840,N_4898);
nor UO_850 (O_850,N_4861,N_4865);
nand UO_851 (O_851,N_4968,N_4969);
nor UO_852 (O_852,N_4816,N_4844);
or UO_853 (O_853,N_4821,N_4882);
or UO_854 (O_854,N_4844,N_4803);
xnor UO_855 (O_855,N_4822,N_4933);
or UO_856 (O_856,N_4836,N_4953);
nand UO_857 (O_857,N_4931,N_4947);
nor UO_858 (O_858,N_4943,N_4936);
or UO_859 (O_859,N_4995,N_4880);
xnor UO_860 (O_860,N_4953,N_4923);
or UO_861 (O_861,N_4847,N_4871);
xnor UO_862 (O_862,N_4818,N_4929);
xor UO_863 (O_863,N_4964,N_4871);
nand UO_864 (O_864,N_4924,N_4885);
nor UO_865 (O_865,N_4840,N_4872);
or UO_866 (O_866,N_4940,N_4929);
and UO_867 (O_867,N_4941,N_4892);
nand UO_868 (O_868,N_4877,N_4858);
or UO_869 (O_869,N_4995,N_4845);
xnor UO_870 (O_870,N_4830,N_4832);
and UO_871 (O_871,N_4818,N_4936);
and UO_872 (O_872,N_4947,N_4844);
and UO_873 (O_873,N_4996,N_4878);
nand UO_874 (O_874,N_4994,N_4944);
or UO_875 (O_875,N_4870,N_4929);
xor UO_876 (O_876,N_4857,N_4850);
or UO_877 (O_877,N_4841,N_4892);
nor UO_878 (O_878,N_4914,N_4994);
and UO_879 (O_879,N_4909,N_4856);
or UO_880 (O_880,N_4940,N_4829);
xnor UO_881 (O_881,N_4850,N_4864);
and UO_882 (O_882,N_4961,N_4816);
nand UO_883 (O_883,N_4809,N_4806);
xor UO_884 (O_884,N_4968,N_4990);
nor UO_885 (O_885,N_4902,N_4899);
nand UO_886 (O_886,N_4842,N_4803);
xnor UO_887 (O_887,N_4878,N_4887);
and UO_888 (O_888,N_4846,N_4887);
and UO_889 (O_889,N_4926,N_4989);
nor UO_890 (O_890,N_4910,N_4879);
nand UO_891 (O_891,N_4993,N_4983);
nor UO_892 (O_892,N_4969,N_4827);
and UO_893 (O_893,N_4890,N_4885);
nand UO_894 (O_894,N_4819,N_4989);
xor UO_895 (O_895,N_4836,N_4875);
nor UO_896 (O_896,N_4993,N_4823);
or UO_897 (O_897,N_4936,N_4965);
or UO_898 (O_898,N_4838,N_4840);
or UO_899 (O_899,N_4918,N_4977);
xnor UO_900 (O_900,N_4815,N_4837);
nand UO_901 (O_901,N_4829,N_4887);
or UO_902 (O_902,N_4808,N_4957);
and UO_903 (O_903,N_4800,N_4916);
xnor UO_904 (O_904,N_4950,N_4941);
or UO_905 (O_905,N_4993,N_4868);
or UO_906 (O_906,N_4845,N_4843);
xnor UO_907 (O_907,N_4821,N_4965);
nand UO_908 (O_908,N_4915,N_4875);
xnor UO_909 (O_909,N_4876,N_4837);
or UO_910 (O_910,N_4934,N_4997);
and UO_911 (O_911,N_4901,N_4989);
xnor UO_912 (O_912,N_4819,N_4884);
nand UO_913 (O_913,N_4873,N_4864);
nor UO_914 (O_914,N_4893,N_4940);
nor UO_915 (O_915,N_4911,N_4824);
and UO_916 (O_916,N_4804,N_4821);
nor UO_917 (O_917,N_4804,N_4892);
nand UO_918 (O_918,N_4872,N_4903);
nor UO_919 (O_919,N_4885,N_4842);
or UO_920 (O_920,N_4834,N_4989);
or UO_921 (O_921,N_4927,N_4830);
nor UO_922 (O_922,N_4885,N_4979);
xnor UO_923 (O_923,N_4818,N_4973);
xnor UO_924 (O_924,N_4813,N_4832);
nor UO_925 (O_925,N_4977,N_4815);
nand UO_926 (O_926,N_4959,N_4807);
or UO_927 (O_927,N_4992,N_4957);
xor UO_928 (O_928,N_4868,N_4801);
nand UO_929 (O_929,N_4892,N_4997);
nand UO_930 (O_930,N_4819,N_4932);
and UO_931 (O_931,N_4818,N_4884);
or UO_932 (O_932,N_4889,N_4818);
nand UO_933 (O_933,N_4865,N_4956);
and UO_934 (O_934,N_4871,N_4849);
nor UO_935 (O_935,N_4802,N_4941);
and UO_936 (O_936,N_4904,N_4866);
xnor UO_937 (O_937,N_4885,N_4940);
nor UO_938 (O_938,N_4820,N_4903);
xor UO_939 (O_939,N_4968,N_4947);
or UO_940 (O_940,N_4932,N_4877);
xor UO_941 (O_941,N_4975,N_4969);
nand UO_942 (O_942,N_4957,N_4989);
or UO_943 (O_943,N_4989,N_4903);
and UO_944 (O_944,N_4887,N_4903);
and UO_945 (O_945,N_4994,N_4913);
and UO_946 (O_946,N_4997,N_4817);
and UO_947 (O_947,N_4801,N_4942);
and UO_948 (O_948,N_4834,N_4957);
or UO_949 (O_949,N_4802,N_4968);
and UO_950 (O_950,N_4814,N_4831);
xnor UO_951 (O_951,N_4970,N_4832);
nand UO_952 (O_952,N_4819,N_4880);
and UO_953 (O_953,N_4970,N_4968);
nor UO_954 (O_954,N_4979,N_4839);
xnor UO_955 (O_955,N_4994,N_4906);
nor UO_956 (O_956,N_4856,N_4822);
xnor UO_957 (O_957,N_4965,N_4815);
xnor UO_958 (O_958,N_4988,N_4957);
nor UO_959 (O_959,N_4863,N_4800);
nand UO_960 (O_960,N_4885,N_4906);
nand UO_961 (O_961,N_4851,N_4826);
xnor UO_962 (O_962,N_4837,N_4992);
xor UO_963 (O_963,N_4907,N_4910);
or UO_964 (O_964,N_4908,N_4883);
and UO_965 (O_965,N_4825,N_4820);
xor UO_966 (O_966,N_4935,N_4820);
xor UO_967 (O_967,N_4943,N_4967);
and UO_968 (O_968,N_4949,N_4972);
and UO_969 (O_969,N_4986,N_4928);
and UO_970 (O_970,N_4952,N_4805);
nor UO_971 (O_971,N_4926,N_4987);
nand UO_972 (O_972,N_4835,N_4831);
nand UO_973 (O_973,N_4820,N_4896);
nand UO_974 (O_974,N_4810,N_4834);
or UO_975 (O_975,N_4839,N_4818);
nand UO_976 (O_976,N_4843,N_4919);
and UO_977 (O_977,N_4866,N_4930);
or UO_978 (O_978,N_4925,N_4965);
and UO_979 (O_979,N_4991,N_4829);
nor UO_980 (O_980,N_4959,N_4850);
and UO_981 (O_981,N_4930,N_4897);
and UO_982 (O_982,N_4945,N_4940);
nand UO_983 (O_983,N_4912,N_4968);
nand UO_984 (O_984,N_4837,N_4926);
or UO_985 (O_985,N_4883,N_4954);
or UO_986 (O_986,N_4982,N_4945);
and UO_987 (O_987,N_4914,N_4995);
xor UO_988 (O_988,N_4832,N_4845);
xor UO_989 (O_989,N_4875,N_4939);
nand UO_990 (O_990,N_4808,N_4811);
or UO_991 (O_991,N_4988,N_4964);
and UO_992 (O_992,N_4992,N_4816);
and UO_993 (O_993,N_4986,N_4973);
nand UO_994 (O_994,N_4905,N_4809);
or UO_995 (O_995,N_4872,N_4923);
nand UO_996 (O_996,N_4808,N_4809);
xnor UO_997 (O_997,N_4847,N_4858);
nor UO_998 (O_998,N_4923,N_4862);
xor UO_999 (O_999,N_4865,N_4955);
endmodule