module basic_2500_25000_3000_50_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_720,In_1740);
nor U1 (N_1,In_1031,In_2399);
nand U2 (N_2,In_1248,In_1602);
and U3 (N_3,In_523,In_2285);
nand U4 (N_4,In_675,In_1022);
nand U5 (N_5,In_297,In_585);
or U6 (N_6,In_837,In_1117);
nor U7 (N_7,In_71,In_373);
nor U8 (N_8,In_741,In_625);
xor U9 (N_9,In_2140,In_980);
and U10 (N_10,In_184,In_1392);
nor U11 (N_11,In_1129,In_1262);
and U12 (N_12,In_31,In_1891);
xnor U13 (N_13,In_2113,In_626);
and U14 (N_14,In_1410,In_1484);
or U15 (N_15,In_1178,In_77);
nor U16 (N_16,In_2169,In_1745);
nand U17 (N_17,In_426,In_1132);
nor U18 (N_18,In_367,In_2210);
xor U19 (N_19,In_598,In_1218);
nand U20 (N_20,In_1126,In_706);
or U21 (N_21,In_1863,In_145);
and U22 (N_22,In_589,In_167);
nor U23 (N_23,In_2281,In_1264);
nand U24 (N_24,In_2111,In_318);
nor U25 (N_25,In_560,In_2149);
nand U26 (N_26,In_2031,In_1186);
or U27 (N_27,In_707,In_1622);
xnor U28 (N_28,In_325,In_2306);
nor U29 (N_29,In_79,In_2312);
or U30 (N_30,In_1676,In_705);
and U31 (N_31,In_410,In_1454);
and U32 (N_32,In_271,In_1746);
and U33 (N_33,In_2311,In_228);
and U34 (N_34,In_1510,In_2290);
nand U35 (N_35,In_1439,In_2337);
nor U36 (N_36,In_1193,In_1690);
nand U37 (N_37,In_1697,In_833);
nor U38 (N_38,In_73,In_1504);
or U39 (N_39,In_1089,In_1919);
nand U40 (N_40,In_463,In_142);
nand U41 (N_41,In_248,In_2093);
xnor U42 (N_42,In_1878,In_402);
nand U43 (N_43,In_1652,In_2171);
nor U44 (N_44,In_173,In_1038);
xor U45 (N_45,In_1292,In_954);
nand U46 (N_46,In_28,In_179);
nor U47 (N_47,In_628,In_2436);
nor U48 (N_48,In_2372,In_836);
nor U49 (N_49,In_542,In_121);
and U50 (N_50,In_2294,In_1511);
nor U51 (N_51,In_199,In_59);
nand U52 (N_52,In_293,In_815);
nand U53 (N_53,In_1389,In_1271);
or U54 (N_54,In_634,In_1087);
and U55 (N_55,In_889,In_1340);
and U56 (N_56,In_1625,In_981);
xor U57 (N_57,In_2075,In_1060);
or U58 (N_58,In_52,In_1099);
or U59 (N_59,In_2099,In_490);
nor U60 (N_60,In_1704,In_290);
and U61 (N_61,In_1495,In_823);
or U62 (N_62,In_1643,In_2247);
nand U63 (N_63,In_1672,In_1836);
or U64 (N_64,In_340,In_2185);
xnor U65 (N_65,In_1378,In_2034);
and U66 (N_66,In_1150,In_1288);
and U67 (N_67,In_1486,In_2127);
or U68 (N_68,In_1924,In_635);
xor U69 (N_69,In_2167,In_372);
nand U70 (N_70,In_668,In_840);
and U71 (N_71,In_1276,In_1658);
or U72 (N_72,In_596,In_1073);
or U73 (N_73,In_1718,In_2462);
and U74 (N_74,In_26,In_1154);
nor U75 (N_75,In_1371,In_85);
or U76 (N_76,In_2023,In_657);
and U77 (N_77,In_245,In_1962);
xnor U78 (N_78,In_1237,In_1061);
or U79 (N_79,In_1959,In_264);
and U80 (N_80,In_216,In_256);
nand U81 (N_81,In_1110,In_2097);
or U82 (N_82,In_1015,In_1654);
nand U83 (N_83,In_1655,In_221);
nand U84 (N_84,In_2304,In_2042);
or U85 (N_85,In_619,In_1966);
and U86 (N_86,In_116,In_1147);
nand U87 (N_87,In_565,In_2349);
or U88 (N_88,In_362,In_496);
nor U89 (N_89,In_467,In_584);
or U90 (N_90,In_1930,In_270);
and U91 (N_91,In_2359,In_2451);
nor U92 (N_92,In_515,In_170);
nand U93 (N_93,In_1070,In_1685);
xnor U94 (N_94,In_1228,In_348);
xor U95 (N_95,In_384,In_855);
or U96 (N_96,In_2418,In_685);
and U97 (N_97,In_2371,In_1967);
nand U98 (N_98,In_1566,In_694);
nor U99 (N_99,In_2340,In_219);
nor U100 (N_100,In_1941,In_1720);
or U101 (N_101,In_1059,In_2427);
or U102 (N_102,In_2276,In_1161);
xor U103 (N_103,In_208,In_242);
nand U104 (N_104,In_1958,In_1463);
nor U105 (N_105,In_2239,In_1257);
nand U106 (N_106,In_739,In_1659);
nand U107 (N_107,In_2492,In_1816);
xor U108 (N_108,In_2231,In_842);
xnor U109 (N_109,In_725,In_1104);
nor U110 (N_110,In_2135,In_1997);
nand U111 (N_111,In_1423,In_189);
xor U112 (N_112,In_2412,In_235);
or U113 (N_113,In_273,In_1838);
nor U114 (N_114,In_2283,In_878);
nand U115 (N_115,In_1977,In_1425);
nor U116 (N_116,In_2491,In_1310);
and U117 (N_117,In_1028,In_234);
nor U118 (N_118,In_1713,In_1611);
nor U119 (N_119,In_1054,In_1435);
or U120 (N_120,In_447,In_1366);
and U121 (N_121,In_2036,In_1557);
nand U122 (N_122,In_385,In_2028);
xor U123 (N_123,In_950,In_1341);
nor U124 (N_124,In_1778,In_1192);
or U125 (N_125,In_1242,In_2490);
and U126 (N_126,In_202,In_1097);
and U127 (N_127,In_1174,In_1402);
and U128 (N_128,In_2019,In_1912);
or U129 (N_129,In_1553,In_289);
nor U130 (N_130,In_529,In_1456);
or U131 (N_131,In_2225,In_2048);
nand U132 (N_132,In_1567,In_727);
xor U133 (N_133,In_1046,In_538);
nor U134 (N_134,In_153,In_1585);
and U135 (N_135,In_1329,In_280);
or U136 (N_136,In_1005,In_737);
or U137 (N_137,In_1278,In_653);
nand U138 (N_138,In_757,In_1267);
nor U139 (N_139,In_2022,In_1837);
or U140 (N_140,In_2360,In_2182);
and U141 (N_141,In_1202,In_1814);
nor U142 (N_142,In_1295,In_343);
nand U143 (N_143,In_2029,In_590);
and U144 (N_144,In_1356,In_866);
nor U145 (N_145,In_1339,In_988);
or U146 (N_146,In_1898,In_2236);
or U147 (N_147,In_1164,In_14);
nor U148 (N_148,In_935,In_1461);
nand U149 (N_149,In_137,In_882);
and U150 (N_150,In_287,In_577);
xnor U151 (N_151,In_1416,In_1214);
or U152 (N_152,In_1010,In_2497);
or U153 (N_153,In_266,In_300);
nand U154 (N_154,In_1268,In_2237);
nand U155 (N_155,In_795,In_1524);
and U156 (N_156,In_647,In_1775);
nand U157 (N_157,In_1305,In_576);
nand U158 (N_158,In_22,In_1088);
or U159 (N_159,In_1342,In_311);
nor U160 (N_160,In_1398,In_2118);
nor U161 (N_161,In_1258,In_1064);
or U162 (N_162,In_6,In_2223);
xnor U163 (N_163,In_1650,In_226);
nand U164 (N_164,In_1732,In_409);
and U165 (N_165,In_1614,In_1063);
nand U166 (N_166,In_32,In_2055);
or U167 (N_167,In_1372,In_453);
nor U168 (N_168,In_1669,In_1594);
or U169 (N_169,In_1049,In_1335);
and U170 (N_170,In_1526,In_279);
xor U171 (N_171,In_620,In_1071);
xor U172 (N_172,In_66,In_1636);
nand U173 (N_173,In_2178,In_528);
and U174 (N_174,In_1448,In_2493);
nor U175 (N_175,In_2068,In_1568);
or U176 (N_176,In_916,In_554);
nor U177 (N_177,In_539,In_2385);
nor U178 (N_178,In_2197,In_2174);
or U179 (N_179,In_1610,In_2170);
nand U180 (N_180,In_2163,In_1715);
and U181 (N_181,In_667,In_1360);
and U182 (N_182,In_1621,In_1348);
nand U183 (N_183,In_860,In_295);
or U184 (N_184,In_1805,In_1647);
or U185 (N_185,In_799,In_717);
or U186 (N_186,In_1331,In_370);
and U187 (N_187,In_1794,In_1355);
nor U188 (N_188,In_1895,In_1586);
or U189 (N_189,In_2152,In_794);
nand U190 (N_190,In_830,In_2015);
nand U191 (N_191,In_1162,In_2448);
nor U192 (N_192,In_2046,In_1503);
and U193 (N_193,In_962,In_2381);
nand U194 (N_194,In_677,In_1918);
nand U195 (N_195,In_901,In_919);
nor U196 (N_196,In_1513,In_407);
nand U197 (N_197,In_1002,In_2063);
nand U198 (N_198,In_1333,In_819);
and U199 (N_199,In_2191,In_2187);
or U200 (N_200,In_704,In_659);
and U201 (N_201,In_1468,In_2350);
or U202 (N_202,In_1130,In_1179);
nand U203 (N_203,In_1896,In_39);
nor U204 (N_204,In_1469,In_485);
nor U205 (N_205,In_2,In_1365);
nand U206 (N_206,In_1656,In_1882);
nand U207 (N_207,In_1693,In_431);
nand U208 (N_208,In_1809,In_1582);
and U209 (N_209,In_2160,In_1082);
nand U210 (N_210,In_1668,In_1779);
nand U211 (N_211,In_973,In_1865);
nand U212 (N_212,In_908,In_2136);
nand U213 (N_213,In_2488,In_438);
nand U214 (N_214,In_2000,In_1216);
nand U215 (N_215,In_277,In_200);
and U216 (N_216,In_381,In_1892);
xnor U217 (N_217,In_387,In_2089);
nor U218 (N_218,In_1824,In_2221);
or U219 (N_219,In_1223,In_2059);
or U220 (N_220,In_133,In_1277);
nand U221 (N_221,In_1489,In_1969);
nor U222 (N_222,In_1180,In_2230);
nor U223 (N_223,In_650,In_884);
or U224 (N_224,In_2400,In_320);
nor U225 (N_225,In_29,In_1711);
and U226 (N_226,In_2030,In_1934);
or U227 (N_227,In_766,In_670);
nor U228 (N_228,In_1888,In_615);
and U229 (N_229,In_1897,In_1768);
or U230 (N_230,In_9,In_1408);
nor U231 (N_231,In_868,In_1079);
nor U232 (N_232,In_1281,In_826);
xor U233 (N_233,In_974,In_1134);
and U234 (N_234,In_1600,In_2278);
nand U235 (N_235,In_1637,In_2269);
nand U236 (N_236,In_12,In_990);
or U237 (N_237,In_427,In_1862);
or U238 (N_238,In_2486,In_2168);
nor U239 (N_239,In_1984,In_2369);
nor U240 (N_240,In_291,In_2244);
nor U241 (N_241,In_2282,In_2014);
nor U242 (N_242,In_20,In_2064);
xnor U243 (N_243,In_850,In_1235);
nor U244 (N_244,In_1675,In_1350);
nor U245 (N_245,In_1203,In_693);
nor U246 (N_246,In_1460,In_504);
xnor U247 (N_247,In_1671,In_939);
and U248 (N_248,In_1128,In_1793);
and U249 (N_249,In_1200,In_240);
nand U250 (N_250,In_1067,In_2235);
nand U251 (N_251,In_2379,In_592);
xnor U252 (N_252,In_1387,In_1390);
or U253 (N_253,In_441,In_905);
and U254 (N_254,In_721,In_1520);
or U255 (N_255,In_588,In_1995);
nand U256 (N_256,In_1290,In_2069);
or U257 (N_257,In_1803,In_1115);
and U258 (N_258,In_471,In_1472);
xnor U259 (N_259,In_1141,In_687);
and U260 (N_260,In_1245,In_1300);
or U261 (N_261,In_975,In_2474);
xnor U262 (N_262,In_2145,In_1095);
and U263 (N_263,In_1436,In_1210);
nand U264 (N_264,In_1666,In_825);
nor U265 (N_265,In_2038,In_1102);
xor U266 (N_266,In_817,In_586);
nor U267 (N_267,In_2256,In_1872);
and U268 (N_268,In_1549,In_672);
or U269 (N_269,In_686,In_449);
or U270 (N_270,In_107,In_437);
or U271 (N_271,In_1617,In_2375);
xor U272 (N_272,In_1558,In_70);
nor U273 (N_273,In_1797,In_2289);
or U274 (N_274,In_1572,In_1755);
nand U275 (N_275,In_1664,In_1197);
nand U276 (N_276,In_2130,In_209);
xor U277 (N_277,In_1120,In_2329);
nor U278 (N_278,In_1771,In_1956);
nand U279 (N_279,In_1287,In_1982);
and U280 (N_280,In_1999,In_928);
xnor U281 (N_281,In_703,In_992);
nand U282 (N_282,In_1113,In_123);
nor U283 (N_283,In_1404,In_1279);
xor U284 (N_284,In_1207,In_2408);
or U285 (N_285,In_1853,In_2142);
xnor U286 (N_286,In_229,In_2246);
nor U287 (N_287,In_1633,In_319);
or U288 (N_288,In_247,In_1873);
or U289 (N_289,In_1788,In_1808);
or U290 (N_290,In_152,In_2121);
or U291 (N_291,In_611,In_652);
nor U292 (N_292,In_1111,In_1595);
and U293 (N_293,In_618,In_811);
nor U294 (N_294,In_1639,In_1249);
xor U295 (N_295,In_37,In_357);
nand U296 (N_296,In_1762,In_644);
or U297 (N_297,In_1494,In_1532);
or U298 (N_298,In_193,In_783);
and U299 (N_299,In_2387,In_1748);
and U300 (N_300,In_1217,In_364);
or U301 (N_301,In_2206,In_2467);
and U302 (N_302,In_1151,In_952);
xnor U303 (N_303,In_654,In_10);
and U304 (N_304,In_1055,In_1584);
nand U305 (N_305,In_995,In_2403);
or U306 (N_306,In_690,In_1770);
and U307 (N_307,In_1050,In_1475);
nor U308 (N_308,In_1388,In_2287);
nor U309 (N_309,In_1972,In_972);
xor U310 (N_310,In_2214,In_1033);
nand U311 (N_311,In_932,In_108);
nor U312 (N_312,In_621,In_1880);
and U313 (N_313,In_2307,In_2021);
nand U314 (N_314,In_1869,In_1326);
or U315 (N_315,In_2266,In_1885);
or U316 (N_316,In_1407,In_24);
xnor U317 (N_317,In_812,In_1457);
nand U318 (N_318,In_1051,In_1138);
nor U319 (N_319,In_1514,In_947);
or U320 (N_320,In_1630,In_2386);
and U321 (N_321,In_669,In_1455);
nand U322 (N_322,In_2071,In_2241);
nor U323 (N_323,In_1726,In_1004);
nor U324 (N_324,In_2346,In_46);
nor U325 (N_325,In_1275,In_1975);
or U326 (N_326,In_2338,In_709);
nand U327 (N_327,In_1802,In_1026);
and U328 (N_328,In_413,In_1767);
or U329 (N_329,In_2261,In_261);
nor U330 (N_330,In_1688,In_651);
and U331 (N_331,In_1907,In_3);
or U332 (N_332,In_2298,In_1789);
or U333 (N_333,In_1399,In_1785);
or U334 (N_334,In_1725,In_788);
or U335 (N_335,In_1719,In_1904);
nor U336 (N_336,In_2079,In_1441);
nand U337 (N_337,In_570,In_1084);
xor U338 (N_338,In_314,In_284);
xor U339 (N_339,In_2006,In_400);
xnor U340 (N_340,In_870,In_689);
and U341 (N_341,In_742,In_2003);
and U342 (N_342,In_486,In_2487);
nor U343 (N_343,In_942,In_65);
nand U344 (N_344,In_1096,In_2199);
nand U345 (N_345,In_171,In_1618);
or U346 (N_346,In_1014,In_726);
xor U347 (N_347,In_904,In_1137);
or U348 (N_348,In_1027,In_1231);
nand U349 (N_349,In_894,In_2330);
nor U350 (N_350,In_1840,In_724);
xnor U351 (N_351,In_81,In_1260);
nand U352 (N_352,In_1478,In_2321);
nand U353 (N_353,In_2115,In_416);
or U354 (N_354,In_500,In_556);
nand U355 (N_355,In_88,In_521);
and U356 (N_356,In_1817,In_177);
or U357 (N_357,In_641,In_1000);
nor U358 (N_358,In_1800,In_1229);
and U359 (N_359,In_350,In_1774);
nor U360 (N_360,In_2056,In_2374);
nor U361 (N_361,In_2322,In_1306);
or U362 (N_362,In_1375,In_2499);
nand U363 (N_363,In_2459,In_30);
or U364 (N_364,In_94,In_637);
nand U365 (N_365,In_1763,In_312);
or U366 (N_366,In_802,In_925);
nand U367 (N_367,In_352,In_822);
or U368 (N_368,In_102,In_646);
or U369 (N_369,In_2481,In_1107);
nand U370 (N_370,In_1699,In_2429);
and U371 (N_371,In_2449,In_2188);
nand U372 (N_372,In_874,In_2423);
nand U373 (N_373,In_1199,In_2143);
nor U374 (N_374,In_2041,In_2421);
and U375 (N_375,In_524,In_391);
xor U376 (N_376,In_327,In_963);
nand U377 (N_377,In_537,In_1724);
or U378 (N_378,In_1533,In_1284);
and U379 (N_379,In_2392,In_2240);
nand U380 (N_380,In_545,In_610);
and U381 (N_381,In_2151,In_1782);
or U382 (N_382,In_425,In_867);
nand U383 (N_383,In_1381,In_1528);
or U384 (N_384,In_1981,In_1976);
xor U385 (N_385,In_2447,In_303);
nand U386 (N_386,In_1221,In_1393);
xnor U387 (N_387,In_2468,In_655);
nor U388 (N_388,In_1860,In_2378);
and U389 (N_389,In_1920,In_821);
nor U390 (N_390,In_1955,In_1634);
nand U391 (N_391,In_227,In_758);
nor U392 (N_392,In_233,In_23);
nand U393 (N_393,In_2013,In_286);
and U394 (N_394,In_483,In_1485);
nor U395 (N_395,In_665,In_2043);
nor U396 (N_396,In_1827,In_1722);
nand U397 (N_397,In_436,In_2284);
nand U398 (N_398,In_747,In_1025);
and U399 (N_399,In_1792,In_1498);
and U400 (N_400,In_1374,In_355);
nor U401 (N_401,In_2470,In_1406);
nor U402 (N_402,In_135,In_2413);
or U403 (N_403,In_1744,In_888);
nand U404 (N_404,In_1307,In_1612);
xor U405 (N_405,In_2415,In_1234);
and U406 (N_406,In_1090,In_13);
nor U407 (N_407,In_609,In_495);
nor U408 (N_408,In_1269,In_760);
or U409 (N_409,In_1246,In_2044);
xor U410 (N_410,In_2229,In_887);
nor U411 (N_411,In_1336,In_536);
and U412 (N_412,In_2137,In_1598);
xnor U413 (N_413,In_382,In_966);
nand U414 (N_414,In_429,In_144);
nand U415 (N_415,In_629,In_2450);
nand U416 (N_416,In_2331,In_337);
nor U417 (N_417,In_2125,In_875);
or U418 (N_418,In_423,In_921);
nor U419 (N_419,In_1285,In_2114);
or U420 (N_420,In_1522,In_1479);
nor U421 (N_421,In_1443,In_859);
nor U422 (N_422,In_2458,In_1509);
nand U423 (N_423,In_87,In_633);
or U424 (N_424,In_1094,In_946);
or U425 (N_425,In_1032,In_307);
nand U426 (N_426,In_1505,In_948);
or U427 (N_427,In_804,In_323);
or U428 (N_428,In_2299,In_702);
nor U429 (N_429,In_164,In_2495);
nand U430 (N_430,In_965,In_205);
nand U431 (N_431,In_787,In_328);
or U432 (N_432,In_1091,In_417);
and U433 (N_433,In_922,In_2325);
or U434 (N_434,In_1382,In_1023);
nor U435 (N_435,In_506,In_891);
or U436 (N_436,In_1707,In_1058);
and U437 (N_437,In_1916,In_2228);
nand U438 (N_438,In_844,In_474);
and U439 (N_439,In_2204,In_961);
xor U440 (N_440,In_2308,In_1327);
or U441 (N_441,In_1674,In_106);
nor U442 (N_442,In_930,In_1950);
or U443 (N_443,In_550,In_2184);
nor U444 (N_444,In_2207,In_1536);
xor U445 (N_445,In_2401,In_1649);
nor U446 (N_446,In_681,In_2345);
nand U447 (N_447,In_843,In_1158);
nor U448 (N_448,In_139,In_36);
or U449 (N_449,In_403,In_298);
and U450 (N_450,In_182,In_1487);
nor U451 (N_451,In_1114,In_743);
and U452 (N_452,In_956,In_767);
nor U453 (N_453,In_2116,In_2479);
nand U454 (N_454,In_604,In_322);
xnor U455 (N_455,In_1039,In_877);
nand U456 (N_456,In_2347,In_674);
and U457 (N_457,In_232,In_2402);
or U458 (N_458,In_2067,In_1261);
or U459 (N_459,In_1537,In_2291);
nor U460 (N_460,In_1444,In_748);
nor U461 (N_461,In_344,In_155);
nor U462 (N_462,In_2243,In_2242);
nand U463 (N_463,In_34,In_1351);
and U464 (N_464,In_1978,In_1282);
nor U465 (N_465,In_1580,In_593);
nor U466 (N_466,In_476,In_829);
nor U467 (N_467,In_8,In_1952);
and U468 (N_468,In_1189,In_1721);
nand U469 (N_469,In_838,In_1222);
or U470 (N_470,In_2198,In_1990);
or U471 (N_471,In_2159,In_648);
nor U472 (N_472,In_2002,In_1302);
xor U473 (N_473,In_1165,In_148);
xor U474 (N_474,In_489,In_1942);
xor U475 (N_475,In_432,In_2292);
and U476 (N_476,In_846,In_1893);
or U477 (N_477,In_365,In_1687);
or U478 (N_478,In_1974,In_873);
nor U479 (N_479,In_1561,In_522);
nand U480 (N_480,In_661,In_1299);
or U481 (N_481,In_1751,In_204);
nand U482 (N_482,In_149,In_1118);
and U483 (N_483,In_1272,In_912);
and U484 (N_484,In_605,In_19);
nor U485 (N_485,In_2265,In_374);
xnor U486 (N_486,In_1211,In_2257);
nand U487 (N_487,In_2303,In_239);
nor U488 (N_488,In_1450,In_1992);
nor U489 (N_489,In_1219,In_2323);
nand U490 (N_490,In_2262,In_161);
and U491 (N_491,In_2212,In_1317);
or U492 (N_492,In_2355,In_444);
nand U493 (N_493,In_442,In_701);
nand U494 (N_494,In_470,In_915);
nor U495 (N_495,In_1806,In_11);
or U496 (N_496,In_2132,In_1951);
nand U497 (N_497,In_110,In_2161);
or U498 (N_498,In_397,In_1101);
or U499 (N_499,In_2357,In_2264);
and U500 (N_500,In_1182,In_1212);
nand U501 (N_501,In_1550,In_1384);
and U502 (N_502,N_137,N_231);
and U503 (N_503,N_162,In_2407);
or U504 (N_504,In_2305,In_631);
or U505 (N_505,In_712,N_496);
and U506 (N_506,N_339,In_359);
nand U507 (N_507,N_109,N_311);
and U508 (N_508,N_29,In_259);
or U509 (N_509,N_244,In_2035);
nor U510 (N_510,In_746,In_722);
xor U511 (N_511,In_733,In_76);
or U512 (N_512,In_892,N_282);
nor U513 (N_513,In_2073,In_2092);
or U514 (N_514,In_510,N_482);
and U515 (N_515,In_1181,In_1359);
nand U516 (N_516,In_810,N_453);
nor U517 (N_517,In_2153,N_235);
and U518 (N_518,In_1964,In_1146);
and U519 (N_519,N_212,In_1620);
nor U520 (N_520,In_1742,In_1121);
or U521 (N_521,In_2367,N_74);
nor U522 (N_522,In_2267,In_2258);
nor U523 (N_523,In_377,In_2461);
nor U524 (N_524,In_310,In_2255);
nand U525 (N_525,N_326,N_99);
and U526 (N_526,In_1349,N_110);
nor U527 (N_527,N_467,In_1946);
or U528 (N_528,In_751,In_580);
xor U529 (N_529,In_1624,In_1850);
xor U530 (N_530,In_768,N_361);
and U531 (N_531,In_630,In_378);
and U532 (N_532,N_272,In_691);
or U533 (N_533,In_1481,N_366);
or U534 (N_534,In_25,In_1205);
and U535 (N_535,In_562,In_516);
nand U536 (N_536,In_1311,In_1108);
and U537 (N_537,N_301,In_390);
nor U538 (N_538,In_852,In_1270);
nand U539 (N_539,In_2016,In_236);
and U540 (N_540,In_885,In_159);
or U541 (N_541,In_91,In_1452);
or U542 (N_542,In_2081,In_1149);
and U543 (N_543,In_1700,In_1519);
nor U544 (N_544,In_1991,N_138);
nor U545 (N_545,N_489,N_225);
nand U546 (N_546,In_481,In_2117);
or U547 (N_547,In_1208,In_1286);
nand U548 (N_548,In_1608,In_1012);
nor U549 (N_549,In_540,In_1507);
nor U550 (N_550,In_2464,N_164);
nor U551 (N_551,In_1705,N_21);
nor U552 (N_552,In_40,In_1188);
and U553 (N_553,In_835,In_1220);
or U554 (N_554,In_190,In_1821);
nor U555 (N_555,In_1944,In_1933);
or U556 (N_556,In_223,N_377);
nand U557 (N_557,In_606,In_341);
nand U558 (N_558,In_587,N_125);
nor U559 (N_559,In_559,In_2384);
and U560 (N_560,In_1322,In_448);
nor U561 (N_561,N_146,In_250);
or U562 (N_562,In_197,In_98);
and U563 (N_563,In_617,In_1686);
nand U564 (N_564,In_1545,N_351);
and U565 (N_565,In_2353,In_1313);
nand U566 (N_566,N_347,In_1822);
and U567 (N_567,In_253,In_774);
and U568 (N_568,In_1823,In_1993);
nand U569 (N_569,In_957,In_2086);
and U570 (N_570,In_1665,In_1777);
nand U571 (N_571,N_411,In_2339);
nor U572 (N_572,In_130,In_2485);
and U573 (N_573,In_958,In_2332);
nor U574 (N_574,N_382,In_1753);
or U575 (N_575,In_1347,In_1852);
nor U576 (N_576,In_195,In_1960);
nor U577 (N_577,In_640,In_1689);
or U578 (N_578,In_96,In_2388);
or U579 (N_579,In_797,In_1616);
nand U580 (N_580,In_612,N_254);
and U581 (N_581,In_2405,In_1274);
nand U582 (N_582,In_2393,In_1851);
nand U583 (N_583,N_178,In_2344);
nor U584 (N_584,N_328,N_83);
nor U585 (N_585,N_462,In_1499);
nor U586 (N_586,In_174,In_1227);
xor U587 (N_587,In_2268,N_132);
xnor U588 (N_588,N_495,In_1380);
or U589 (N_589,In_1145,N_472);
and U590 (N_590,In_479,N_223);
nand U591 (N_591,In_968,In_2273);
nand U592 (N_592,In_1921,In_1125);
xnor U593 (N_593,In_2109,In_679);
and U594 (N_594,In_1900,In_1615);
and U595 (N_595,In_1515,In_1609);
nor U596 (N_596,In_1623,In_993);
nand U597 (N_597,In_469,In_2422);
or U598 (N_598,N_457,In_2324);
nor U599 (N_599,In_571,In_1925);
nand U600 (N_600,In_778,N_488);
nand U601 (N_601,In_740,In_1787);
nor U602 (N_602,In_2072,In_1170);
nand U603 (N_603,In_1994,In_696);
or U604 (N_604,In_175,In_2248);
and U605 (N_605,In_780,In_2453);
nand U606 (N_606,In_1529,In_666);
or U607 (N_607,In_2380,In_169);
nor U608 (N_608,N_243,In_1847);
nand U609 (N_609,In_2414,N_395);
xor U610 (N_610,In_1597,N_234);
nor U611 (N_611,In_752,In_1829);
nor U612 (N_612,In_132,In_1815);
xor U613 (N_613,In_2215,N_118);
nand U614 (N_614,In_366,In_1035);
and U615 (N_615,In_487,In_35);
and U616 (N_616,N_70,In_1948);
or U617 (N_617,In_1931,In_1963);
and U618 (N_618,N_207,In_55);
and U619 (N_619,In_944,In_1908);
xor U620 (N_620,N_88,N_232);
xnor U621 (N_621,In_1497,In_2120);
xor U622 (N_622,In_1702,N_475);
xor U623 (N_623,N_497,N_251);
and U624 (N_624,In_1646,N_155);
nor U625 (N_625,N_72,N_181);
nor U626 (N_626,In_158,N_278);
or U627 (N_627,N_102,N_421);
nand U628 (N_628,In_1488,In_1016);
nand U629 (N_629,In_67,In_1083);
or U630 (N_630,In_1954,In_194);
xnor U631 (N_631,In_104,In_2444);
nor U632 (N_632,In_602,In_2440);
nor U633 (N_633,In_1343,In_346);
nor U634 (N_634,In_2186,In_156);
or U635 (N_635,In_2219,In_1502);
xor U636 (N_636,N_376,N_403);
xor U637 (N_637,In_2105,In_1019);
or U638 (N_638,In_2439,N_370);
or U639 (N_639,In_1266,In_2226);
nand U640 (N_640,In_201,In_945);
nand U641 (N_641,N_481,In_1098);
or U642 (N_642,In_543,In_181);
nand U643 (N_643,N_152,In_484);
xnor U644 (N_644,In_1133,In_1660);
nor U645 (N_645,In_2314,In_770);
nand U646 (N_646,In_1419,N_424);
or U647 (N_647,In_533,N_43);
nand U648 (N_648,In_492,In_1081);
nor U649 (N_649,In_50,In_1731);
nor U650 (N_650,N_218,N_92);
nor U651 (N_651,N_237,In_1143);
nor U652 (N_652,In_399,In_2274);
and U653 (N_653,In_1801,In_1607);
nor U654 (N_654,N_480,In_1679);
nor U655 (N_655,N_156,N_38);
nor U656 (N_656,In_1560,N_194);
and U657 (N_657,In_404,In_2051);
and U658 (N_658,N_458,In_15);
nand U659 (N_659,In_781,In_512);
xor U660 (N_660,In_575,In_1048);
nand U661 (N_661,In_1581,In_1877);
nand U662 (N_662,In_600,N_362);
and U663 (N_663,In_2074,In_1103);
or U664 (N_664,N_327,In_1241);
and U665 (N_665,In_80,N_261);
xnor U666 (N_666,In_549,In_557);
xnor U667 (N_667,In_1571,N_294);
nand U668 (N_668,In_1759,N_193);
nand U669 (N_669,In_180,In_996);
or U670 (N_670,In_54,In_2196);
and U671 (N_671,In_714,In_2482);
or U672 (N_672,In_1338,In_154);
nand U673 (N_673,In_255,In_63);
or U674 (N_674,N_3,N_476);
and U675 (N_675,In_594,In_1011);
and U676 (N_676,In_1879,In_2173);
nor U677 (N_677,N_179,In_899);
and U678 (N_678,In_1176,In_1140);
or U679 (N_679,In_2363,In_1473);
nand U680 (N_680,In_363,In_74);
nor U681 (N_681,N_471,In_1739);
nor U682 (N_682,In_1303,In_597);
xnor U683 (N_683,N_36,In_986);
and U684 (N_684,In_452,N_290);
and U685 (N_685,In_841,In_926);
nand U686 (N_686,In_1804,In_534);
or U687 (N_687,In_2376,N_53);
or U688 (N_688,N_75,In_933);
nor U689 (N_689,N_324,In_1551);
nor U690 (N_690,In_2122,In_983);
nand U691 (N_691,In_1124,N_211);
or U692 (N_692,N_104,In_456);
nand U693 (N_693,In_1255,In_1044);
and U694 (N_694,In_309,In_1476);
and U695 (N_695,N_459,In_764);
and U696 (N_696,In_1345,In_1890);
xor U697 (N_697,In_338,In_90);
xnor U698 (N_698,In_1983,N_428);
or U699 (N_699,N_60,In_1163);
and U700 (N_700,N_203,In_1527);
or U701 (N_701,In_532,N_0);
or U702 (N_702,In_2404,In_1427);
or U703 (N_703,In_1727,N_460);
or U704 (N_704,In_2279,In_1265);
or U705 (N_705,N_49,In_1232);
nor U706 (N_706,N_18,In_663);
or U707 (N_707,In_715,In_1243);
and U708 (N_708,N_107,In_1166);
and U709 (N_709,In_1663,N_464);
or U710 (N_710,In_393,In_1587);
or U711 (N_711,In_383,In_1631);
or U712 (N_712,In_1238,In_2101);
or U713 (N_713,In_57,In_1516);
and U714 (N_714,In_698,In_2483);
or U715 (N_715,In_1324,In_115);
nand U716 (N_716,In_2334,N_337);
and U717 (N_717,In_1386,In_1155);
nor U718 (N_718,In_1849,N_95);
nor U719 (N_719,In_433,N_430);
or U720 (N_720,In_1889,In_2012);
nor U721 (N_721,In_1321,In_1492);
nand U722 (N_722,In_333,In_723);
xor U723 (N_723,In_971,In_2008);
nand U724 (N_724,In_977,N_112);
nand U725 (N_725,In_895,N_135);
and U726 (N_726,N_389,In_69);
or U727 (N_727,N_160,In_1909);
xnor U728 (N_728,In_1940,N_69);
nand U729 (N_729,N_50,In_1965);
and U730 (N_730,In_514,In_1854);
nand U731 (N_731,In_354,In_301);
or U732 (N_732,In_501,In_1304);
or U733 (N_733,N_438,N_305);
nand U734 (N_734,In_2466,In_424);
or U735 (N_735,N_58,In_520);
or U736 (N_736,N_283,N_293);
and U737 (N_737,In_2417,In_1449);
nand U738 (N_738,In_1541,N_423);
nand U739 (N_739,N_270,In_1191);
nor U740 (N_740,In_2455,In_269);
nor U741 (N_741,In_361,N_71);
nand U742 (N_742,In_48,In_527);
xor U743 (N_743,N_449,In_1483);
nand U744 (N_744,In_2217,In_2033);
and U745 (N_745,N_46,In_1783);
xnor U746 (N_746,In_2430,In_1986);
nand U747 (N_747,In_428,In_466);
or U748 (N_748,In_1694,N_418);
or U749 (N_749,N_6,In_1482);
nor U750 (N_750,N_285,In_1506);
xnor U751 (N_751,In_775,In_553);
or U752 (N_752,In_392,In_2496);
nor U753 (N_753,In_1501,N_4);
or U754 (N_754,In_1319,In_831);
or U755 (N_755,In_2394,N_260);
nand U756 (N_756,In_1412,In_955);
or U757 (N_757,In_530,In_305);
and U758 (N_758,N_226,In_358);
nand U759 (N_759,In_531,In_497);
or U760 (N_760,N_85,In_2213);
nand U761 (N_761,In_949,In_2150);
nor U762 (N_762,In_1065,In_2252);
and U763 (N_763,In_1825,In_1259);
and U764 (N_764,In_2045,N_62);
and U765 (N_765,In_1325,In_1644);
and U766 (N_766,In_1013,N_122);
and U767 (N_767,N_219,In_713);
and U768 (N_768,In_700,In_1438);
nor U769 (N_769,In_1206,N_175);
xnor U770 (N_770,In_334,In_517);
nor U771 (N_771,N_227,N_335);
nand U772 (N_772,In_166,N_47);
and U773 (N_773,In_1430,N_266);
nand U774 (N_774,In_1741,In_2205);
and U775 (N_775,In_2098,In_214);
nor U776 (N_776,N_350,N_490);
and U777 (N_777,In_813,In_1040);
nand U778 (N_778,In_1451,In_386);
nand U779 (N_779,In_1714,In_468);
xnor U780 (N_780,N_412,In_509);
and U781 (N_781,N_360,In_1169);
nand U782 (N_782,N_10,In_1641);
or U783 (N_783,In_1429,In_1037);
nand U784 (N_784,In_763,In_1760);
nor U785 (N_785,In_2434,In_480);
and U786 (N_786,N_343,In_272);
nand U787 (N_787,In_548,N_413);
and U788 (N_788,In_1021,In_1565);
or U789 (N_789,In_2475,N_291);
and U790 (N_790,In_60,In_561);
nor U791 (N_791,In_1196,In_1373);
or U792 (N_792,In_2437,In_246);
nor U793 (N_793,N_494,In_1968);
nand U794 (N_794,In_579,N_149);
nand U795 (N_795,N_279,In_1250);
or U796 (N_796,N_257,N_236);
or U797 (N_797,In_676,In_1605);
nand U798 (N_798,In_1517,In_849);
nand U799 (N_799,In_1552,In_692);
nor U800 (N_800,In_2432,N_348);
nand U801 (N_801,N_20,In_75);
nor U802 (N_802,In_574,In_1943);
nor U803 (N_803,In_1283,In_2358);
or U804 (N_804,N_499,In_2313);
nand U805 (N_805,N_113,In_2473);
xor U806 (N_806,N_470,In_342);
nand U807 (N_807,N_323,In_865);
nand U808 (N_808,In_931,In_907);
nand U809 (N_809,N_134,In_1296);
xor U810 (N_810,In_1923,N_142);
or U811 (N_811,In_1394,In_1947);
nand U812 (N_812,In_1396,In_789);
or U813 (N_813,In_909,In_206);
and U814 (N_814,In_756,In_964);
or U815 (N_815,N_280,In_1691);
nor U816 (N_816,In_541,In_738);
nand U817 (N_817,N_150,In_558);
or U818 (N_818,In_27,In_881);
nand U819 (N_819,In_118,In_2017);
or U820 (N_820,In_398,N_174);
and U821 (N_821,N_222,In_1183);
and U822 (N_822,In_2441,N_163);
or U823 (N_823,In_302,In_1883);
nand U824 (N_824,In_2001,In_1914);
nand U825 (N_825,In_879,In_454);
nor U826 (N_826,In_2083,In_2032);
or U827 (N_827,N_309,N_247);
nand U828 (N_828,In_2200,In_994);
and U829 (N_829,In_1330,N_435);
nand U830 (N_830,In_1471,In_1508);
or U831 (N_831,In_2465,N_268);
or U832 (N_832,In_2218,In_2175);
xnor U833 (N_833,In_736,In_2420);
or U834 (N_834,In_1297,In_2254);
and U835 (N_835,N_190,In_1420);
nor U836 (N_836,N_114,In_2395);
nor U837 (N_837,In_2335,In_2445);
and U838 (N_838,In_1701,In_1201);
xor U839 (N_839,In_1734,N_491);
and U840 (N_840,In_1034,N_123);
and U841 (N_841,In_505,In_238);
or U842 (N_842,In_1077,In_2094);
and U843 (N_843,In_1173,In_2201);
and U844 (N_844,In_656,N_451);
nand U845 (N_845,In_678,In_332);
nand U846 (N_846,N_319,N_84);
and U847 (N_847,N_307,N_82);
or U848 (N_848,In_2181,N_406);
nand U849 (N_849,In_1379,N_383);
nor U850 (N_850,N_444,In_645);
nor U851 (N_851,In_1209,In_188);
nor U852 (N_852,In_172,In_1928);
xnor U853 (N_853,In_1577,In_1627);
nand U854 (N_854,N_292,N_271);
nor U855 (N_855,N_252,In_900);
or U856 (N_856,In_2472,In_1953);
and U857 (N_857,N_240,In_176);
nor U858 (N_858,In_109,In_406);
nand U859 (N_859,In_987,In_914);
nand U860 (N_860,N_98,In_1766);
or U861 (N_861,In_56,In_616);
nand U862 (N_862,In_2253,In_1698);
or U863 (N_863,In_1328,In_997);
or U864 (N_864,N_2,In_929);
nand U865 (N_865,In_1579,In_160);
nand U866 (N_866,N_466,In_1555);
nor U867 (N_867,In_1100,N_169);
nand U868 (N_868,N_298,In_330);
or U869 (N_869,In_1020,In_1601);
and U870 (N_870,In_1085,In_1047);
and U871 (N_871,In_1546,N_454);
or U872 (N_872,In_2148,N_40);
nand U873 (N_873,In_1,N_365);
or U874 (N_874,N_191,In_1105);
and U875 (N_875,In_2194,In_1361);
or U876 (N_876,In_1810,N_57);
and U877 (N_877,In_1233,In_1651);
nor U878 (N_878,N_202,In_636);
or U879 (N_879,In_1431,In_2452);
xor U880 (N_880,In_1036,In_1198);
and U881 (N_881,N_213,N_461);
nor U882 (N_882,N_129,In_658);
xnor U883 (N_883,In_443,In_49);
nand U884 (N_884,In_1080,N_7);
or U885 (N_885,In_1403,In_2179);
xnor U886 (N_886,In_808,N_105);
nor U887 (N_887,In_1606,In_420);
or U888 (N_888,In_1142,In_759);
nor U889 (N_889,In_1291,In_72);
nand U890 (N_890,In_1225,In_1477);
xor U891 (N_891,In_178,In_1240);
nor U892 (N_892,In_276,N_16);
xor U893 (N_893,In_78,In_274);
and U894 (N_894,In_267,In_4);
or U895 (N_895,N_124,In_2476);
and U896 (N_896,N_385,In_1069);
nand U897 (N_897,N_204,In_2435);
nand U898 (N_898,In_459,N_422);
and U899 (N_899,In_412,In_1613);
xnor U900 (N_900,In_526,In_1353);
and U901 (N_901,In_818,In_1057);
and U902 (N_902,In_324,In_1906);
or U903 (N_903,N_269,In_1007);
nand U904 (N_904,In_688,In_2095);
xnor U905 (N_905,In_2352,In_1383);
nand U906 (N_906,In_2146,N_79);
nand U907 (N_907,N_145,In_1042);
nand U908 (N_908,In_624,In_1708);
xnor U909 (N_909,N_442,In_430);
nor U910 (N_910,N_14,In_112);
or U911 (N_911,In_511,N_111);
or U912 (N_912,In_664,In_1358);
and U913 (N_913,In_140,N_469);
nor U914 (N_914,In_1973,N_297);
nand U915 (N_915,In_1289,In_2124);
and U916 (N_916,In_2202,In_719);
nor U917 (N_917,In_2365,In_1543);
nand U918 (N_918,In_2007,In_2088);
and U919 (N_919,In_2164,In_136);
or U920 (N_920,In_2158,In_2061);
nor U921 (N_921,N_159,In_2477);
nand U922 (N_922,In_2020,In_1677);
and U923 (N_923,In_380,In_1831);
and U924 (N_924,N_437,In_729);
nand U925 (N_925,In_296,N_346);
nand U926 (N_926,N_183,In_784);
and U927 (N_927,In_2119,In_710);
nor U928 (N_928,N_277,In_2131);
xor U929 (N_929,In_2251,In_2233);
nand U930 (N_930,In_2070,N_117);
nor U931 (N_931,N_276,In_231);
or U932 (N_932,In_1599,N_331);
and U933 (N_933,In_591,In_2342);
nand U934 (N_934,In_89,In_1712);
or U935 (N_935,In_660,In_744);
or U936 (N_936,In_151,In_285);
and U937 (N_937,N_439,In_258);
nand U938 (N_938,In_1252,In_1445);
nor U939 (N_939,In_1569,In_845);
and U940 (N_940,In_1542,In_1866);
or U941 (N_941,N_434,In_1521);
and U942 (N_942,In_1160,N_59);
and U943 (N_943,In_2368,In_1682);
and U944 (N_944,In_1397,In_2126);
or U945 (N_945,N_315,In_2366);
nor U946 (N_946,In_1177,In_1913);
or U947 (N_947,In_16,In_100);
nor U948 (N_948,In_371,In_1078);
nand U949 (N_949,In_762,N_478);
nor U950 (N_950,N_168,In_1428);
and U951 (N_951,In_1703,In_854);
xor U952 (N_952,In_2260,In_1812);
nor U953 (N_953,In_779,N_167);
nand U954 (N_954,In_2416,N_255);
nand U955 (N_955,N_26,In_2377);
and U956 (N_956,In_2442,In_2049);
nor U957 (N_957,N_126,N_87);
nor U958 (N_958,In_886,In_1459);
and U959 (N_959,In_2356,In_750);
nor U960 (N_960,N_64,In_1418);
nand U961 (N_961,In_1131,In_525);
xor U962 (N_962,In_1540,In_2310);
or U963 (N_963,N_397,In_1761);
nor U964 (N_964,In_445,N_368);
nor U965 (N_965,In_2288,In_2300);
nor U966 (N_966,In_2383,In_349);
xnor U967 (N_967,In_786,In_2208);
nand U968 (N_968,In_2227,In_1405);
nor U969 (N_969,N_52,In_614);
or U970 (N_970,In_478,N_41);
xor U971 (N_971,In_765,In_1979);
nand U972 (N_972,N_425,In_1156);
nor U973 (N_973,In_880,N_304);
and U974 (N_974,In_1411,N_19);
nand U975 (N_975,In_1167,In_460);
or U976 (N_976,In_2220,In_1442);
or U977 (N_977,In_47,In_599);
nand U978 (N_978,N_61,In_1153);
and U979 (N_979,In_2027,In_1780);
nor U980 (N_980,In_1045,In_473);
nor U981 (N_981,In_168,In_2026);
or U982 (N_982,N_133,In_198);
xor U983 (N_983,In_212,In_1758);
and U984 (N_984,N_394,In_38);
or U985 (N_985,In_2156,In_1936);
nand U986 (N_986,N_456,In_1263);
and U987 (N_987,In_2155,N_372);
and U988 (N_988,In_1204,In_2084);
and U989 (N_989,In_572,In_1628);
nand U990 (N_990,In_213,In_1056);
and U991 (N_991,In_1716,In_2471);
xor U992 (N_992,In_1312,In_2060);
nor U993 (N_993,In_2460,N_208);
nand U994 (N_994,N_65,N_479);
and U995 (N_995,In_1743,In_1747);
xnor U996 (N_996,In_1518,N_352);
nand U997 (N_997,In_2054,In_435);
xor U998 (N_998,In_1662,N_9);
nand U999 (N_999,In_419,N_22);
nand U1000 (N_1000,N_740,N_386);
and U1001 (N_1001,N_97,N_448);
or U1002 (N_1002,In_1564,N_926);
xor U1003 (N_1003,In_2295,In_1440);
and U1004 (N_1004,In_2428,In_1368);
and U1005 (N_1005,N_344,N_743);
nand U1006 (N_1006,In_2052,In_861);
and U1007 (N_1007,In_451,N_500);
nor U1008 (N_1008,N_724,In_493);
or U1009 (N_1009,N_586,N_556);
nor U1010 (N_1010,N_948,N_539);
and U1011 (N_1011,In_989,N_680);
or U1012 (N_1012,N_721,N_568);
nand U1013 (N_1013,In_237,N_32);
nor U1014 (N_1014,N_120,N_686);
and U1015 (N_1015,N_958,In_2489);
and U1016 (N_1016,N_988,In_1523);
or U1017 (N_1017,N_843,In_967);
or U1018 (N_1018,In_1554,N_100);
xnor U1019 (N_1019,N_103,In_1692);
xor U1020 (N_1020,N_116,In_1813);
nor U1021 (N_1021,N_419,In_1570);
or U1022 (N_1022,N_465,N_674);
xor U1023 (N_1023,In_103,In_1680);
nand U1024 (N_1024,In_2478,In_940);
or U1025 (N_1025,N_230,N_836);
nor U1026 (N_1026,N_978,N_66);
or U1027 (N_1027,N_834,In_1846);
nor U1028 (N_1028,In_331,In_793);
nor U1029 (N_1029,In_1902,N_875);
nor U1030 (N_1030,In_824,N_601);
or U1031 (N_1031,N_527,In_547);
and U1032 (N_1032,N_144,In_1795);
nor U1033 (N_1033,N_563,N_310);
or U1034 (N_1034,N_596,In_1024);
and U1035 (N_1035,In_141,In_2058);
and U1036 (N_1036,In_394,N_514);
nor U1037 (N_1037,In_1168,N_287);
nand U1038 (N_1038,N_147,In_329);
xor U1039 (N_1039,In_2018,In_1127);
and U1040 (N_1040,N_391,N_776);
xor U1041 (N_1041,In_2104,N_822);
nand U1042 (N_1042,In_2154,In_896);
nand U1043 (N_1043,N_517,In_82);
nand U1044 (N_1044,N_443,N_771);
xor U1045 (N_1045,N_522,In_1172);
and U1046 (N_1046,In_2389,In_2316);
or U1047 (N_1047,N_340,In_1706);
nor U1048 (N_1048,In_150,N_486);
xnor U1049 (N_1049,In_498,In_2039);
and U1050 (N_1050,In_1834,N_387);
or U1051 (N_1051,N_729,In_44);
nor U1052 (N_1052,In_1735,In_2100);
nor U1053 (N_1053,In_1244,N_78);
xnor U1054 (N_1054,In_2362,N_275);
and U1055 (N_1055,In_1251,In_126);
and U1056 (N_1056,N_940,N_637);
nand U1057 (N_1057,N_807,In_1985);
nor U1058 (N_1058,N_374,N_508);
xor U1059 (N_1059,In_1480,In_2147);
or U1060 (N_1060,In_796,N_170);
nor U1061 (N_1061,N_265,In_53);
and U1062 (N_1062,In_2222,In_211);
nor U1063 (N_1063,N_610,N_862);
and U1064 (N_1064,N_989,In_2062);
nand U1065 (N_1065,N_758,N_599);
or U1066 (N_1066,In_1603,In_388);
or U1067 (N_1067,N_653,N_629);
nand U1068 (N_1068,In_1736,N_652);
and U1069 (N_1069,N_802,N_380);
nand U1070 (N_1070,N_784,In_1857);
nor U1071 (N_1071,In_2328,In_991);
nor U1072 (N_1072,In_2319,In_1332);
xnor U1073 (N_1073,In_2107,N_700);
and U1074 (N_1074,N_838,In_801);
or U1075 (N_1075,N_242,In_313);
nor U1076 (N_1076,N_668,In_777);
nand U1077 (N_1077,In_1346,N_584);
nand U1078 (N_1078,In_243,N_583);
or U1079 (N_1079,In_1917,N_349);
or U1080 (N_1080,In_257,In_1109);
xnor U1081 (N_1081,N_992,N_741);
and U1082 (N_1082,N_54,N_646);
or U1083 (N_1083,N_613,N_590);
and U1084 (N_1084,In_1556,N_728);
or U1085 (N_1085,In_379,In_809);
and U1086 (N_1086,N_999,N_927);
xor U1087 (N_1087,N_895,N_264);
and U1088 (N_1088,In_1987,In_1935);
or U1089 (N_1089,N_157,N_764);
xor U1090 (N_1090,N_224,In_1458);
nand U1091 (N_1091,N_216,In_1915);
nand U1092 (N_1092,N_955,In_1756);
or U1093 (N_1093,In_923,In_730);
or U1094 (N_1094,N_986,N_694);
or U1095 (N_1095,N_656,N_763);
and U1096 (N_1096,In_1213,N_742);
or U1097 (N_1097,In_51,N_679);
and U1098 (N_1098,In_1757,N_964);
nand U1099 (N_1099,N_1,N_587);
nand U1100 (N_1100,In_2108,In_422);
or U1101 (N_1101,In_1009,In_1548);
and U1102 (N_1102,N_712,N_687);
and U1103 (N_1103,N_115,N_650);
and U1104 (N_1104,In_1790,N_493);
nor U1105 (N_1105,N_15,N_249);
or U1106 (N_1106,In_2406,N_543);
or U1107 (N_1107,In_503,In_1575);
and U1108 (N_1108,In_1422,N_515);
nor U1109 (N_1109,In_1563,In_7);
or U1110 (N_1110,In_567,In_2096);
nor U1111 (N_1111,N_919,N_636);
or U1112 (N_1112,In_434,In_1224);
nor U1113 (N_1113,N_228,N_332);
or U1114 (N_1114,N_518,In_871);
nand U1115 (N_1115,N_663,N_195);
nand U1116 (N_1116,In_1638,N_855);
or U1117 (N_1117,N_312,N_336);
or U1118 (N_1118,N_820,In_1157);
and U1119 (N_1119,In_1709,In_294);
xnor U1120 (N_1120,N_367,N_956);
nand U1121 (N_1121,N_847,In_2189);
and U1122 (N_1122,In_95,In_1052);
and U1123 (N_1123,N_531,In_1512);
nor U1124 (N_1124,In_2327,In_2162);
nor U1125 (N_1125,N_993,In_1534);
nor U1126 (N_1126,In_1717,In_1253);
nand U1127 (N_1127,N_384,In_632);
or U1128 (N_1128,In_131,N_705);
or U1129 (N_1129,In_1635,In_910);
or U1130 (N_1130,N_373,In_623);
xor U1131 (N_1131,In_421,In_315);
nand U1132 (N_1132,N_585,In_513);
and U1133 (N_1133,In_551,In_292);
nand U1134 (N_1134,N_965,N_452);
nor U1135 (N_1135,In_2180,In_1629);
or U1136 (N_1136,In_1899,In_1971);
and U1137 (N_1137,In_832,In_1437);
nand U1138 (N_1138,In_937,In_1092);
nand U1139 (N_1139,In_1937,In_2382);
and U1140 (N_1140,In_1401,N_842);
nor U1141 (N_1141,In_1415,N_564);
nand U1142 (N_1142,N_791,In_639);
and U1143 (N_1143,N_794,In_564);
and U1144 (N_1144,N_198,N_987);
nand U1145 (N_1145,In_1573,N_617);
nor U1146 (N_1146,In_191,In_898);
and U1147 (N_1147,N_833,In_2438);
nor U1148 (N_1148,In_482,In_1074);
and U1149 (N_1149,N_562,In_1043);
or U1150 (N_1150,N_683,In_450);
xor U1151 (N_1151,N_852,N_766);
nand U1152 (N_1152,N_872,In_1786);
nor U1153 (N_1153,N_379,In_1194);
nor U1154 (N_1154,In_1842,N_809);
xnor U1155 (N_1155,N_405,N_513);
or U1156 (N_1156,N_253,In_1843);
or U1157 (N_1157,In_1750,In_1695);
nand U1158 (N_1158,N_554,N_849);
nor U1159 (N_1159,In_1493,In_827);
or U1160 (N_1160,In_1905,In_1500);
nand U1161 (N_1161,In_1819,In_1939);
or U1162 (N_1162,N_404,N_546);
nor U1163 (N_1163,N_672,N_34);
or U1164 (N_1164,N_189,In_2011);
nor U1165 (N_1165,In_336,N_248);
xor U1166 (N_1166,N_831,In_2193);
and U1167 (N_1167,N_426,In_1236);
or U1168 (N_1168,N_577,In_2396);
nand U1169 (N_1169,In_2297,In_1945);
and U1170 (N_1170,In_1645,N_187);
or U1171 (N_1171,In_2271,N_303);
or U1172 (N_1172,N_358,N_619);
and U1173 (N_1173,In_1344,In_2080);
and U1174 (N_1174,N_647,In_749);
xor U1175 (N_1175,In_1764,N_432);
nand U1176 (N_1176,N_567,N_560);
and U1177 (N_1177,N_258,In_1314);
or U1178 (N_1178,In_2195,In_461);
nor U1179 (N_1179,In_1465,In_465);
nand U1180 (N_1180,In_578,In_117);
and U1181 (N_1181,N_675,N_591);
or U1182 (N_1182,N_798,N_719);
and U1183 (N_1183,N_308,In_1592);
nor U1184 (N_1184,N_552,N_745);
and U1185 (N_1185,In_1773,In_83);
or U1186 (N_1186,N_979,In_1041);
nand U1187 (N_1187,N_976,In_2398);
nand U1188 (N_1188,In_1354,N_706);
xnor U1189 (N_1189,N_638,N_417);
xor U1190 (N_1190,In_1003,N_555);
xor U1191 (N_1191,N_941,N_805);
nand U1192 (N_1192,In_2301,N_876);
or U1193 (N_1193,In_2139,N_846);
nand U1194 (N_1194,In_673,In_138);
nor U1195 (N_1195,N_911,In_627);
nor U1196 (N_1196,In_1938,In_1776);
nor U1197 (N_1197,N_953,N_512);
or U1198 (N_1198,N_778,N_789);
nor U1199 (N_1199,In_769,N_982);
xnor U1200 (N_1200,In_475,In_288);
nor U1201 (N_1201,N_889,In_782);
nand U1202 (N_1202,In_1175,N_375);
nand U1203 (N_1203,N_594,N_684);
nand U1204 (N_1204,N_787,In_1316);
nor U1205 (N_1205,N_67,N_576);
or U1206 (N_1206,N_381,In_2232);
xnor U1207 (N_1207,In_1886,In_1447);
nor U1208 (N_1208,In_1596,In_275);
nor U1209 (N_1209,N_844,N_803);
nor U1210 (N_1210,In_125,N_906);
nor U1211 (N_1211,N_811,N_474);
and U1212 (N_1212,N_727,N_313);
and U1213 (N_1213,In_573,In_2457);
nor U1214 (N_1214,N_983,N_571);
and U1215 (N_1215,In_1106,In_369);
nor U1216 (N_1216,N_215,In_2005);
and U1217 (N_1217,In_1491,In_1593);
or U1218 (N_1218,N_779,N_813);
and U1219 (N_1219,In_943,N_643);
xnor U1220 (N_1220,In_2091,N_994);
or U1221 (N_1221,N_582,In_1075);
or U1222 (N_1222,N_734,N_892);
or U1223 (N_1223,N_628,In_1910);
and U1224 (N_1224,N_837,In_2431);
xor U1225 (N_1225,In_42,In_368);
nand U1226 (N_1226,N_288,In_941);
or U1227 (N_1227,N_607,N_511);
or U1228 (N_1228,In_984,In_970);
and U1229 (N_1229,N_267,N_51);
and U1230 (N_1230,In_2425,In_2203);
and U1231 (N_1231,In_2351,In_1929);
and U1232 (N_1232,In_1839,N_295);
or U1233 (N_1233,In_872,In_122);
nand U1234 (N_1234,N_655,In_1875);
nand U1235 (N_1235,N_93,In_2172);
nand U1236 (N_1236,In_1738,N_910);
nand U1237 (N_1237,In_2123,In_569);
nor U1238 (N_1238,In_613,In_680);
nand U1239 (N_1239,N_561,In_1867);
and U1240 (N_1240,In_1791,N_693);
or U1241 (N_1241,In_2224,N_540);
and U1242 (N_1242,N_781,In_356);
xnor U1243 (N_1243,In_1215,N_664);
nand U1244 (N_1244,In_642,N_73);
or U1245 (N_1245,In_953,N_429);
or U1246 (N_1246,In_263,In_1068);
nor U1247 (N_1247,In_396,N_657);
nand U1248 (N_1248,In_249,N_37);
nand U1249 (N_1249,N_783,N_286);
or U1250 (N_1250,N_905,In_1308);
and U1251 (N_1251,In_2037,In_1996);
nor U1252 (N_1252,In_1864,N_708);
nor U1253 (N_1253,In_1841,In_734);
xor U1254 (N_1254,N_130,In_316);
nand U1255 (N_1255,In_375,N_960);
nor U1256 (N_1256,N_681,N_357);
or U1257 (N_1257,N_185,In_405);
nor U1258 (N_1258,In_1171,In_192);
nand U1259 (N_1259,In_917,N_942);
and U1260 (N_1260,N_840,N_544);
or U1261 (N_1261,In_196,N_777);
or U1262 (N_1262,In_2433,In_1076);
nor U1263 (N_1263,N_874,N_492);
and U1264 (N_1264,N_732,N_881);
nand U1265 (N_1265,N_81,In_753);
or U1266 (N_1266,In_120,N_171);
nor U1267 (N_1267,In_1195,In_816);
nor U1268 (N_1268,In_682,N_615);
nand U1269 (N_1269,N_612,In_1723);
or U1270 (N_1270,N_559,N_990);
xnor U1271 (N_1271,In_0,In_1256);
or U1272 (N_1272,N_502,N_634);
nor U1273 (N_1273,N_866,In_2270);
xnor U1274 (N_1274,In_1377,In_1417);
or U1275 (N_1275,In_1657,In_251);
xor U1276 (N_1276,In_1826,In_439);
or U1277 (N_1277,N_897,N_334);
nor U1278 (N_1278,In_1811,N_934);
or U1279 (N_1279,In_1066,In_2286);
and U1280 (N_1280,N_931,In_1395);
xnor U1281 (N_1281,In_1247,In_2053);
and U1282 (N_1282,In_1642,N_551);
nand U1283 (N_1283,N_871,N_670);
nor U1284 (N_1284,N_35,N_642);
and U1285 (N_1285,N_440,In_924);
and U1286 (N_1286,N_468,In_1784);
nor U1287 (N_1287,N_427,N_765);
nand U1288 (N_1288,In_1871,N_832);
and U1289 (N_1289,N_96,In_218);
xnor U1290 (N_1290,In_1547,N_900);
xnor U1291 (N_1291,In_1932,In_1490);
nand U1292 (N_1292,N_962,N_715);
nor U1293 (N_1293,In_230,N_950);
nor U1294 (N_1294,N_633,N_436);
nor U1295 (N_1295,In_1626,In_207);
and U1296 (N_1296,N_245,In_2390);
nand U1297 (N_1297,In_1730,N_501);
nand U1298 (N_1298,In_607,N_322);
xor U1299 (N_1299,In_959,N_127);
nand U1300 (N_1300,In_807,In_508);
nor U1301 (N_1301,In_856,N_678);
and U1302 (N_1302,N_192,In_2106);
or U1303 (N_1303,In_772,N_302);
nor U1304 (N_1304,In_2480,N_143);
or U1305 (N_1305,In_165,In_847);
nand U1306 (N_1306,N_505,In_918);
nand U1307 (N_1307,N_42,In_1414);
nand U1308 (N_1308,N_761,N_767);
or U1309 (N_1309,In_776,In_2190);
nand U1310 (N_1310,N_817,N_648);
and U1311 (N_1311,In_1187,N_356);
or U1312 (N_1312,N_918,N_716);
and U1313 (N_1313,In_790,In_1799);
nand U1314 (N_1314,In_828,N_259);
xnor U1315 (N_1315,N_161,N_595);
nand U1316 (N_1316,N_209,In_268);
or U1317 (N_1317,N_883,N_536);
or U1318 (N_1318,N_148,N_593);
and U1319 (N_1319,N_790,N_980);
and U1320 (N_1320,N_720,N_616);
or U1321 (N_1321,N_547,In_1818);
nor U1322 (N_1322,N_446,In_1859);
nand U1323 (N_1323,In_2272,In_299);
nor U1324 (N_1324,In_252,N_68);
nand U1325 (N_1325,N_318,N_600);
nor U1326 (N_1326,In_1334,In_1927);
xnor U1327 (N_1327,In_2456,N_824);
xnor U1328 (N_1328,In_1619,In_1421);
xnor U1329 (N_1329,In_462,In_1884);
nand U1330 (N_1330,N_858,In_58);
nor U1331 (N_1331,In_1640,N_848);
nor U1332 (N_1332,N_153,In_1018);
or U1333 (N_1333,N_797,In_1673);
nor U1334 (N_1334,N_364,N_523);
nand U1335 (N_1335,In_814,N_701);
and U1336 (N_1336,N_48,N_973);
or U1337 (N_1337,In_1578,N_695);
nand U1338 (N_1338,N_826,In_1670);
and U1339 (N_1339,In_876,In_697);
or U1340 (N_1340,N_851,N_723);
or U1341 (N_1341,N_839,In_731);
and U1342 (N_1342,In_1391,In_1752);
xor U1343 (N_1343,N_775,N_507);
nand U1344 (N_1344,N_542,In_45);
and U1345 (N_1345,In_1008,N_136);
or U1346 (N_1346,In_353,N_341);
nand U1347 (N_1347,In_114,N_932);
nor U1348 (N_1348,In_308,N_525);
and U1349 (N_1349,In_1294,N_816);
or U1350 (N_1350,N_974,In_1737);
or U1351 (N_1351,N_572,N_498);
or U1352 (N_1352,N_354,N_27);
nor U1353 (N_1353,N_885,In_1832);
nand U1354 (N_1354,N_754,In_2010);
or U1355 (N_1355,N_682,In_43);
nor U1356 (N_1356,In_1830,N_378);
xnor U1357 (N_1357,N_333,In_1400);
and U1358 (N_1358,In_1796,In_1868);
and U1359 (N_1359,In_2354,N_273);
or U1360 (N_1360,N_954,N_604);
nor U1361 (N_1361,In_1881,N_5);
and U1362 (N_1362,N_902,N_710);
and U1363 (N_1363,N_575,N_923);
nor U1364 (N_1364,In_1072,In_2454);
nand U1365 (N_1365,N_861,N_904);
or U1366 (N_1366,In_1280,N_24);
nor U1367 (N_1367,In_339,In_1123);
nand U1368 (N_1368,In_414,In_1574);
nand U1369 (N_1369,In_1957,In_1184);
nor U1370 (N_1370,N_256,In_1861);
or U1371 (N_1371,N_524,In_1926);
xnor U1372 (N_1372,In_806,In_1772);
or U1373 (N_1373,In_1844,N_961);
xnor U1374 (N_1374,In_1998,N_952);
and U1375 (N_1375,In_2040,N_131);
nor U1376 (N_1376,In_1017,N_165);
and U1377 (N_1377,N_690,N_658);
and U1378 (N_1378,In_893,In_162);
nand U1379 (N_1379,In_1293,N_80);
and U1380 (N_1380,In_1848,N_399);
or U1381 (N_1381,In_1535,In_1901);
nand U1382 (N_1382,N_210,In_1544);
and U1383 (N_1383,In_897,N_11);
or U1384 (N_1384,N_939,N_602);
or U1385 (N_1385,In_906,In_622);
nand U1386 (N_1386,N_972,In_1190);
nand U1387 (N_1387,N_618,N_151);
nand U1388 (N_1388,In_2484,In_803);
xor U1389 (N_1389,N_532,N_935);
nor U1390 (N_1390,N_867,In_735);
nand U1391 (N_1391,N_408,In_99);
or U1392 (N_1392,In_472,N_274);
nand U1393 (N_1393,In_853,N_856);
nor U1394 (N_1394,N_450,In_1728);
and U1395 (N_1395,N_206,In_1434);
or U1396 (N_1396,N_859,In_2494);
or U1397 (N_1397,N_519,N_912);
or U1398 (N_1398,In_2141,In_2165);
nand U1399 (N_1399,N_641,N_56);
nand U1400 (N_1400,N_31,N_995);
nor U1401 (N_1401,In_858,N_317);
nand U1402 (N_1402,N_549,N_217);
nor U1403 (N_1403,In_911,In_1876);
xnor U1404 (N_1404,N_808,N_250);
and U1405 (N_1405,In_86,N_566);
and U1406 (N_1406,N_553,N_863);
and U1407 (N_1407,N_750,In_834);
and U1408 (N_1408,N_473,N_77);
or U1409 (N_1409,N_673,In_2411);
and U1410 (N_1410,In_1413,In_2078);
nor U1411 (N_1411,In_699,N_830);
nor U1412 (N_1412,In_101,In_1230);
xnor U1413 (N_1413,In_415,In_2102);
nand U1414 (N_1414,N_238,N_338);
and U1415 (N_1415,N_371,In_2443);
nor U1416 (N_1416,In_851,N_214);
nand U1417 (N_1417,In_1116,In_1139);
xnor U1418 (N_1418,In_716,N_550);
nand U1419 (N_1419,In_464,N_398);
xnor U1420 (N_1420,N_933,In_2103);
nand U1421 (N_1421,N_627,N_947);
nor U1422 (N_1422,N_692,N_548);
or U1423 (N_1423,N_76,N_484);
nand U1424 (N_1424,In_33,In_335);
xnor U1425 (N_1425,N_624,N_401);
nand U1426 (N_1426,N_951,N_857);
nand U1427 (N_1427,N_821,In_2259);
or U1428 (N_1428,In_982,N_483);
and U1429 (N_1429,N_485,N_321);
xor U1430 (N_1430,In_1576,In_1754);
nor U1431 (N_1431,N_284,N_908);
nor U1432 (N_1432,In_2333,N_773);
nand U1433 (N_1433,In_1362,In_864);
nand U1434 (N_1434,In_1474,In_1856);
and U1435 (N_1435,In_265,N_106);
nor U1436 (N_1436,N_685,N_815);
nand U1437 (N_1437,N_581,In_603);
nand U1438 (N_1438,In_568,In_2057);
nand U1439 (N_1439,N_186,In_638);
xnor U1440 (N_1440,N_534,N_891);
nand U1441 (N_1441,N_262,N_899);
and U1442 (N_1442,N_608,In_711);
and U1443 (N_1443,In_1254,N_25);
and U1444 (N_1444,In_2280,N_810);
or U1445 (N_1445,N_896,N_718);
nor U1446 (N_1446,N_199,N_611);
and U1447 (N_1447,In_1185,In_304);
or U1448 (N_1448,In_217,N_879);
xnor U1449 (N_1449,N_221,N_414);
xor U1450 (N_1450,In_326,N_711);
nor U1451 (N_1451,N_929,N_667);
or U1452 (N_1452,N_589,N_957);
nor U1453 (N_1453,N_239,In_68);
nand U1454 (N_1454,N_510,In_1988);
and U1455 (N_1455,In_21,In_2177);
xnor U1456 (N_1456,N_702,N_12);
and U1457 (N_1457,In_920,N_455);
nor U1458 (N_1458,N_966,In_820);
nand U1459 (N_1459,N_725,N_632);
or U1460 (N_1460,N_119,In_1667);
xnor U1461 (N_1461,In_491,N_263);
nor U1462 (N_1462,In_2302,In_2446);
xnor U1463 (N_1463,In_1239,N_785);
and U1464 (N_1464,In_1989,N_63);
nand U1465 (N_1465,In_1769,In_1318);
and U1466 (N_1466,N_806,N_937);
or U1467 (N_1467,N_55,In_985);
nand U1468 (N_1468,N_825,In_1590);
nor U1469 (N_1469,N_86,N_909);
and U1470 (N_1470,N_829,N_393);
and U1471 (N_1471,N_870,In_1858);
xor U1472 (N_1472,In_2318,In_862);
and U1473 (N_1473,N_369,In_2183);
nor U1474 (N_1474,N_128,N_353);
and U1475 (N_1475,In_2364,N_620);
nand U1476 (N_1476,In_203,N_565);
nor U1477 (N_1477,In_1781,N_845);
nand U1478 (N_1478,N_752,N_409);
or U1479 (N_1479,N_865,N_39);
or U1480 (N_1480,In_695,In_883);
xnor U1481 (N_1481,N_33,N_696);
nor U1482 (N_1482,In_262,In_282);
or U1483 (N_1483,In_800,In_1798);
or U1484 (N_1484,In_241,In_649);
and U1485 (N_1485,N_697,In_411);
and U1486 (N_1486,In_2277,In_1562);
xnor U1487 (N_1487,In_395,In_1298);
or U1488 (N_1488,N_182,N_689);
or U1489 (N_1489,In_1949,N_173);
or U1490 (N_1490,In_2320,N_869);
nand U1491 (N_1491,N_760,N_759);
or U1492 (N_1492,In_2469,In_1462);
nor U1493 (N_1493,N_17,In_754);
xnor U1494 (N_1494,In_2245,N_528);
nor U1495 (N_1495,N_850,In_2309);
nand U1496 (N_1496,N_28,N_996);
nand U1497 (N_1497,In_2211,In_1765);
or U1498 (N_1498,N_597,In_2176);
and U1499 (N_1499,N_184,In_1807);
or U1500 (N_1500,N_306,N_792);
nand U1501 (N_1501,N_1181,In_1367);
and U1502 (N_1502,N_916,In_581);
nor U1503 (N_1503,N_1240,N_1325);
nand U1504 (N_1504,N_1331,N_530);
xor U1505 (N_1505,N_44,In_1001);
or U1506 (N_1506,N_1061,N_698);
or U1507 (N_1507,N_1289,N_1366);
nor U1508 (N_1508,In_119,N_944);
nor U1509 (N_1509,N_854,In_1855);
and U1510 (N_1510,N_1047,In_902);
nor U1511 (N_1511,N_521,N_1390);
xnor U1512 (N_1512,N_1490,N_1424);
or U1513 (N_1513,N_1114,N_1017);
nor U1514 (N_1514,In_183,In_1470);
nand U1515 (N_1515,N_731,N_1297);
or U1516 (N_1516,N_1388,N_1479);
or U1517 (N_1517,N_177,N_289);
or U1518 (N_1518,N_1264,N_1391);
or U1519 (N_1519,N_1343,N_967);
nand U1520 (N_1520,In_771,N_1410);
xor U1521 (N_1521,In_2326,N_1445);
and U1522 (N_1522,N_1043,N_1276);
nor U1523 (N_1523,N_1427,N_296);
xor U1524 (N_1524,N_1131,N_1204);
nand U1525 (N_1525,N_1179,In_2087);
and U1526 (N_1526,N_755,N_749);
and U1527 (N_1527,In_1591,N_1356);
and U1528 (N_1528,N_1392,In_583);
nand U1529 (N_1529,N_1076,N_538);
and U1530 (N_1530,N_1214,In_1226);
and U1531 (N_1531,N_1444,N_1373);
nor U1532 (N_1532,N_1038,N_1109);
and U1533 (N_1533,In_1029,In_1369);
or U1534 (N_1534,N_1482,In_97);
xnor U1535 (N_1535,N_1067,N_780);
nand U1536 (N_1536,N_1273,N_1421);
and U1537 (N_1537,N_1160,N_1168);
nand U1538 (N_1538,N_1074,In_1409);
nand U1539 (N_1539,In_507,N_868);
or U1540 (N_1540,In_2315,N_665);
or U1541 (N_1541,N_1012,N_1124);
nand U1542 (N_1542,In_254,In_1357);
xnor U1543 (N_1543,N_314,N_886);
and U1544 (N_1544,N_1229,In_1030);
and U1545 (N_1545,N_1130,N_1357);
and U1546 (N_1546,N_1073,N_1227);
or U1547 (N_1547,N_943,N_1353);
nand U1548 (N_1548,N_1233,N_1494);
or U1549 (N_1549,In_938,N_1150);
nor U1550 (N_1550,N_415,N_1217);
and U1551 (N_1551,N_445,N_1174);
or U1552 (N_1552,In_1538,N_903);
nor U1553 (N_1553,N_1021,In_1678);
nor U1554 (N_1554,N_1161,N_1420);
xor U1555 (N_1555,N_666,N_1219);
nand U1556 (N_1556,N_659,N_1055);
xnor U1557 (N_1557,N_1122,N_1417);
nand U1558 (N_1558,N_981,N_1246);
or U1559 (N_1559,N_1381,In_2348);
or U1560 (N_1560,In_1112,In_1661);
nor U1561 (N_1561,N_1272,N_1468);
xor U1562 (N_1562,N_1423,N_1016);
xor U1563 (N_1563,N_1462,N_1039);
and U1564 (N_1564,N_1360,N_299);
nor U1565 (N_1565,N_1371,N_90);
or U1566 (N_1566,N_1441,In_2361);
and U1567 (N_1567,N_1393,N_1165);
or U1568 (N_1568,N_503,In_1653);
xor U1569 (N_1569,N_1163,N_799);
or U1570 (N_1570,N_1015,N_812);
nor U1571 (N_1571,N_558,N_1476);
and U1572 (N_1572,N_246,In_1453);
nand U1573 (N_1573,N_985,N_662);
and U1574 (N_1574,N_1389,In_61);
nand U1575 (N_1575,N_1025,N_1030);
nor U1576 (N_1576,N_1250,N_930);
or U1577 (N_1577,N_959,N_1042);
nand U1578 (N_1578,N_1457,N_1375);
nor U1579 (N_1579,In_1870,N_1265);
nand U1580 (N_1580,In_2424,N_101);
nand U1581 (N_1581,In_1604,N_1166);
nor U1582 (N_1582,N_1162,N_233);
or U1583 (N_1583,In_84,N_1148);
and U1584 (N_1584,N_1314,In_1683);
nand U1585 (N_1585,N_733,N_823);
or U1586 (N_1586,N_801,N_1268);
nand U1587 (N_1587,N_1094,In_1309);
nand U1588 (N_1588,In_1530,N_1285);
nand U1589 (N_1589,N_220,N_1075);
nor U1590 (N_1590,N_400,N_1492);
nand U1591 (N_1591,In_283,N_1127);
or U1592 (N_1592,In_2209,N_1434);
or U1593 (N_1593,N_1238,N_1339);
nand U1594 (N_1594,In_903,N_1121);
and U1595 (N_1595,N_579,N_1132);
nor U1596 (N_1596,In_1894,In_2296);
or U1597 (N_1597,In_519,N_1172);
nand U1598 (N_1598,N_1348,N_1173);
and U1599 (N_1599,In_458,In_785);
and U1600 (N_1600,N_1093,N_1129);
and U1601 (N_1601,N_860,N_1065);
nor U1602 (N_1602,N_325,N_688);
or U1603 (N_1603,N_176,N_1266);
and U1604 (N_1604,In_260,In_934);
nand U1605 (N_1605,N_1399,N_1102);
nor U1606 (N_1606,N_1470,N_1080);
nor U1607 (N_1607,In_2373,N_533);
xor U1608 (N_1608,In_662,N_1054);
nand U1609 (N_1609,In_1135,In_1062);
or U1610 (N_1610,In_2336,N_1472);
or U1611 (N_1611,N_717,In_347);
or U1612 (N_1612,N_1205,N_574);
nand U1613 (N_1613,In_2463,In_2144);
nor U1614 (N_1614,N_938,N_1011);
nand U1615 (N_1615,N_1275,In_111);
nor U1616 (N_1616,In_455,N_1278);
or U1617 (N_1617,N_1281,N_1310);
and U1618 (N_1618,N_671,N_1244);
and U1619 (N_1619,In_2112,N_1334);
nand U1620 (N_1620,N_949,In_608);
or U1621 (N_1621,N_1036,N_1257);
or U1622 (N_1622,N_1328,N_1247);
nand U1623 (N_1623,N_609,N_1137);
nor U1624 (N_1624,N_793,In_544);
and U1625 (N_1625,N_915,N_1253);
nor U1626 (N_1626,N_898,N_1005);
nand U1627 (N_1627,N_1270,In_1152);
and U1628 (N_1628,N_1008,N_172);
xnor U1629 (N_1629,N_1092,In_1887);
and U1630 (N_1630,In_1053,In_1588);
and U1631 (N_1631,N_1459,N_1083);
and U1632 (N_1632,N_1305,N_541);
nor U1633 (N_1633,N_1386,In_1352);
and U1634 (N_1634,N_747,N_1286);
or U1635 (N_1635,N_1403,N_1318);
nand U1636 (N_1636,N_1018,N_1026);
nor U1637 (N_1637,In_1681,N_1400);
nand U1638 (N_1638,N_1347,N_936);
and U1639 (N_1639,N_738,N_506);
and U1640 (N_1640,N_1406,N_1048);
nor U1641 (N_1641,In_2110,N_922);
nand U1642 (N_1642,In_1006,N_1213);
nor U1643 (N_1643,In_1632,In_671);
xnor U1644 (N_1644,N_1480,N_736);
or U1645 (N_1645,N_1136,In_2009);
and U1646 (N_1646,N_569,N_1464);
nand U1647 (N_1647,N_1224,In_1385);
or U1648 (N_1648,N_827,In_863);
nor U1649 (N_1649,In_951,In_2343);
xor U1650 (N_1650,N_573,N_463);
nor U1651 (N_1651,In_913,N_1226);
nor U1652 (N_1652,N_1133,N_1070);
nor U1653 (N_1653,N_707,In_732);
nand U1654 (N_1654,N_1396,N_1260);
or U1655 (N_1655,In_317,N_1117);
nor U1656 (N_1656,N_94,N_800);
nor U1657 (N_1657,N_1419,In_976);
and U1658 (N_1658,N_691,In_791);
nand U1659 (N_1659,N_1113,N_880);
or U1660 (N_1660,In_2192,N_1171);
nor U1661 (N_1661,N_1199,In_41);
or U1662 (N_1662,N_1319,N_1294);
or U1663 (N_1663,N_1426,N_1153);
nor U1664 (N_1664,In_2129,N_1118);
or U1665 (N_1665,N_1169,N_1157);
nand U1666 (N_1666,N_1290,N_1032);
nor U1667 (N_1667,N_744,In_643);
nor U1668 (N_1668,In_1301,N_316);
or U1669 (N_1669,In_2397,N_1465);
nor U1670 (N_1670,N_1194,N_1336);
and U1671 (N_1671,N_1338,In_683);
nor U1672 (N_1672,In_92,In_1589);
and U1673 (N_1673,N_1183,N_1354);
nand U1674 (N_1674,N_487,In_2391);
nand U1675 (N_1675,N_772,N_1301);
nor U1676 (N_1676,In_1376,N_1258);
nand U1677 (N_1677,N_1064,N_1033);
xnor U1678 (N_1678,N_1222,N_1323);
or U1679 (N_1679,N_1430,N_1442);
nand U1680 (N_1680,N_1218,In_134);
nand U1681 (N_1681,In_345,In_566);
nand U1682 (N_1682,N_1085,N_1359);
nand U1683 (N_1683,In_2128,N_1486);
and U1684 (N_1684,N_1197,N_23);
and U1685 (N_1685,In_857,N_1091);
and U1686 (N_1686,N_1287,N_1088);
xnor U1687 (N_1687,N_1378,N_1329);
nor U1688 (N_1688,N_1449,N_433);
and U1689 (N_1689,In_563,N_1300);
and U1690 (N_1690,N_977,In_1119);
nand U1691 (N_1691,N_1414,In_147);
and U1692 (N_1692,N_1372,In_2166);
nand U1693 (N_1693,N_1170,N_1466);
nor U1694 (N_1694,N_1164,N_1404);
nand U1695 (N_1695,N_1201,N_431);
and U1696 (N_1696,N_1198,N_1242);
or U1697 (N_1697,N_1180,N_1139);
or U1698 (N_1698,N_1200,N_1066);
or U1699 (N_1699,N_774,In_1835);
or U1700 (N_1700,N_1071,In_2498);
nand U1701 (N_1701,N_924,N_1436);
xnor U1702 (N_1702,N_1498,N_407);
or U1703 (N_1703,N_1023,N_1098);
nand U1704 (N_1704,In_1323,N_1195);
nor U1705 (N_1705,N_1340,N_201);
and U1706 (N_1706,N_639,N_1060);
xor U1707 (N_1707,N_606,N_1481);
nand U1708 (N_1708,N_1202,N_420);
or U1709 (N_1709,N_888,In_1820);
and U1710 (N_1710,N_1089,N_1437);
xnor U1711 (N_1711,N_158,In_792);
and U1712 (N_1712,N_1107,In_869);
and U1713 (N_1713,N_281,N_946);
nand U1714 (N_1714,N_726,N_1176);
and U1715 (N_1715,N_884,In_936);
and U1716 (N_1716,In_440,In_105);
and U1717 (N_1717,N_89,In_157);
or U1718 (N_1718,N_1283,N_1215);
and U1719 (N_1719,In_1136,N_1143);
xor U1720 (N_1720,N_1236,In_2157);
and U1721 (N_1721,N_1376,N_704);
nor U1722 (N_1722,In_1426,N_1463);
xor U1723 (N_1723,N_1077,N_1031);
or U1724 (N_1724,In_2085,N_1364);
or U1725 (N_1725,N_1370,N_907);
nor U1726 (N_1726,N_1046,N_8);
xnor U1727 (N_1727,N_1495,In_1370);
or U1728 (N_1728,N_1271,N_1259);
or U1729 (N_1729,N_1432,In_761);
and U1730 (N_1730,N_1304,N_1072);
nand U1731 (N_1731,N_1125,N_1374);
or U1732 (N_1732,In_1980,N_756);
nor U1733 (N_1733,N_570,N_703);
nor U1734 (N_1734,N_1138,N_1431);
and U1735 (N_1735,N_997,N_1411);
nor U1736 (N_1736,N_1177,N_526);
nand U1737 (N_1737,N_1096,N_1497);
nor U1738 (N_1738,N_1225,N_1159);
nor U1739 (N_1739,In_2216,N_1141);
nor U1740 (N_1740,N_1438,N_1435);
nand U1741 (N_1741,N_1081,N_1483);
nand U1742 (N_1742,N_1317,In_1466);
and U1743 (N_1743,In_848,N_1134);
nand U1744 (N_1744,N_1087,In_546);
and U1745 (N_1745,In_601,N_913);
xnor U1746 (N_1746,N_1001,In_186);
nor U1747 (N_1747,In_224,N_1450);
or U1748 (N_1748,In_185,N_1428);
and U1749 (N_1749,N_1221,N_537);
nor U1750 (N_1750,N_1346,N_1344);
nor U1751 (N_1751,N_1309,In_2082);
nor U1752 (N_1752,In_1424,N_416);
and U1753 (N_1753,N_769,N_1337);
and U1754 (N_1754,N_1341,N_1057);
and U1755 (N_1755,N_196,In_798);
or U1756 (N_1756,N_669,N_1175);
nand U1757 (N_1757,N_1298,In_2133);
nand U1758 (N_1758,In_1315,N_516);
nand U1759 (N_1759,N_392,N_1108);
xnor U1760 (N_1760,N_1440,N_166);
nor U1761 (N_1761,N_991,In_2076);
or U1762 (N_1762,In_1961,N_1100);
or U1763 (N_1763,N_1312,N_1135);
nor U1764 (N_1764,N_1156,In_1086);
or U1765 (N_1765,N_1115,In_728);
xnor U1766 (N_1766,N_677,In_127);
or U1767 (N_1767,N_1377,N_661);
or U1768 (N_1768,N_1333,In_2426);
or U1769 (N_1769,In_1337,In_2317);
nor U1770 (N_1770,In_17,N_1013);
and U1771 (N_1771,N_1368,N_1321);
nor U1772 (N_1772,N_1387,N_818);
nor U1773 (N_1773,N_739,N_1362);
or U1774 (N_1774,N_737,In_360);
xor U1775 (N_1775,N_1140,N_535);
xnor U1776 (N_1776,In_1531,N_1178);
nand U1777 (N_1777,N_592,In_839);
nand U1778 (N_1778,N_795,N_631);
nand U1779 (N_1779,In_62,N_1053);
nand U1780 (N_1780,N_1447,In_582);
nor U1781 (N_1781,N_1208,N_1052);
nand U1782 (N_1782,N_644,N_1320);
and U1783 (N_1783,N_746,In_2238);
and U1784 (N_1784,N_635,N_1473);
nand U1785 (N_1785,N_1296,N_410);
and U1786 (N_1786,N_963,N_1041);
nor U1787 (N_1787,N_1186,In_745);
nand U1788 (N_1788,N_545,In_278);
xor U1789 (N_1789,N_1184,N_1471);
and U1790 (N_1790,N_241,In_2066);
nor U1791 (N_1791,In_1525,N_1489);
nor U1792 (N_1792,N_1352,N_757);
or U1793 (N_1793,In_376,N_1101);
and U1794 (N_1794,N_1454,In_351);
nand U1795 (N_1795,In_2410,In_1464);
nor U1796 (N_1796,N_188,N_1349);
and U1797 (N_1797,N_388,N_1332);
xor U1798 (N_1798,N_396,N_504);
xnor U1799 (N_1799,N_853,N_925);
or U1800 (N_1800,N_1063,N_1147);
and U1801 (N_1801,N_614,N_649);
xnor U1802 (N_1802,N_1151,N_1413);
nand U1803 (N_1803,In_2250,N_1461);
and U1804 (N_1804,N_998,N_1196);
and U1805 (N_1805,N_205,N_1216);
nor U1806 (N_1806,N_108,N_1188);
or U1807 (N_1807,N_580,N_1282);
or U1808 (N_1808,N_1384,N_1451);
nand U1809 (N_1809,In_684,In_1874);
and U1810 (N_1810,N_1149,N_229);
and U1811 (N_1811,N_762,N_1330);
and U1812 (N_1812,N_320,N_1029);
nand U1813 (N_1813,N_873,N_1326);
or U1814 (N_1814,N_1496,N_1261);
nand U1815 (N_1815,In_129,N_1019);
or U1816 (N_1816,In_1903,N_1009);
or U1817 (N_1817,N_768,N_1220);
nand U1818 (N_1818,In_1559,N_1002);
nor U1819 (N_1819,N_441,N_782);
and U1820 (N_1820,In_1446,N_1382);
nand U1821 (N_1821,In_499,N_598);
nand U1822 (N_1822,N_1103,N_1439);
nor U1823 (N_1823,N_1119,N_1397);
nand U1824 (N_1824,N_660,N_1493);
nor U1825 (N_1825,In_2077,N_1485);
nor U1826 (N_1826,N_121,N_1004);
nor U1827 (N_1827,In_408,In_1733);
and U1828 (N_1828,In_502,N_894);
nand U1829 (N_1829,N_1086,N_1269);
and U1830 (N_1830,In_998,N_1256);
and U1831 (N_1831,N_1475,N_1154);
nor U1832 (N_1832,In_210,In_281);
or U1833 (N_1833,N_1237,In_2134);
nand U1834 (N_1834,N_402,N_1024);
nor U1835 (N_1835,In_960,In_1833);
and U1836 (N_1836,In_187,N_1104);
nor U1837 (N_1837,N_713,N_1034);
or U1838 (N_1838,N_1313,In_1467);
nand U1839 (N_1839,N_1288,N_1144);
and U1840 (N_1840,N_1235,N_1488);
xor U1841 (N_1841,In_1320,N_1499);
nand U1842 (N_1842,In_1432,In_2025);
or U1843 (N_1843,N_1418,N_1010);
and U1844 (N_1844,In_595,N_1241);
nand U1845 (N_1845,N_1245,N_329);
nand U1846 (N_1846,N_1409,In_143);
nand U1847 (N_1847,N_1267,In_2065);
or U1848 (N_1848,In_5,In_113);
and U1849 (N_1849,N_1453,N_901);
or U1850 (N_1850,N_1028,N_975);
or U1851 (N_1851,N_1279,N_1448);
xnor U1852 (N_1852,N_1316,N_140);
and U1853 (N_1853,N_45,N_945);
nor U1854 (N_1854,N_835,N_1090);
nand U1855 (N_1855,N_714,In_927);
nor U1856 (N_1856,In_999,N_1308);
xor U1857 (N_1857,In_1159,N_622);
or U1858 (N_1858,N_1307,N_1416);
and U1859 (N_1859,N_1000,N_1206);
nor U1860 (N_1860,N_1401,N_722);
xnor U1861 (N_1861,In_1363,N_1458);
and U1862 (N_1862,N_1491,N_1478);
or U1863 (N_1863,In_494,N_1128);
or U1864 (N_1864,N_1209,N_1355);
nor U1865 (N_1865,N_751,N_578);
and U1866 (N_1866,In_1093,N_1223);
nor U1867 (N_1867,N_1187,N_1099);
nor U1868 (N_1868,N_1110,In_222);
or U1869 (N_1869,In_1710,N_359);
nand U1870 (N_1870,N_300,In_1148);
or U1871 (N_1871,N_1097,N_1429);
nor U1872 (N_1872,N_1232,N_640);
and U1873 (N_1873,N_605,N_1003);
nor U1874 (N_1874,N_1014,In_418);
or U1875 (N_1875,N_1207,N_1105);
and U1876 (N_1876,In_2275,N_1210);
nor U1877 (N_1877,N_557,In_488);
xnor U1878 (N_1878,N_1079,N_154);
nor U1879 (N_1879,In_2234,N_676);
nor U1880 (N_1880,N_971,In_1696);
and U1881 (N_1881,N_621,In_718);
nor U1882 (N_1882,In_64,N_1456);
nor U1883 (N_1883,In_18,N_1212);
and U1884 (N_1884,N_804,N_1415);
nor U1885 (N_1885,N_917,N_882);
or U1886 (N_1886,N_1365,N_1040);
xor U1887 (N_1887,N_753,N_1189);
nor U1888 (N_1888,N_1255,N_1069);
nand U1889 (N_1889,N_625,N_748);
and U1890 (N_1890,N_1251,N_970);
nor U1891 (N_1891,N_1056,N_1243);
nor U1892 (N_1892,N_363,N_1082);
and U1893 (N_1893,N_1363,In_969);
nand U1894 (N_1894,N_1350,In_446);
nor U1895 (N_1895,N_1049,In_2370);
and U1896 (N_1896,N_623,N_921);
xnor U1897 (N_1897,N_1351,N_699);
and U1898 (N_1898,N_200,N_1050);
nor U1899 (N_1899,N_1078,N_969);
or U1900 (N_1900,In_225,In_477);
xnor U1901 (N_1901,In_1144,In_555);
xnor U1902 (N_1902,In_1122,N_529);
nor U1903 (N_1903,N_1292,N_91);
nand U1904 (N_1904,N_890,N_1185);
nor U1905 (N_1905,N_141,N_1191);
nor U1906 (N_1906,N_1477,N_796);
nand U1907 (N_1907,In_1729,N_709);
xor U1908 (N_1908,N_1303,N_1280);
nor U1909 (N_1909,N_1203,N_1422);
xnor U1910 (N_1910,In_1970,In_1648);
nand U1911 (N_1911,N_1395,N_1231);
and U1912 (N_1912,N_345,N_1367);
nor U1913 (N_1913,N_1302,N_1120);
and U1914 (N_1914,In_518,N_1412);
nand U1915 (N_1915,N_1380,N_139);
xor U1916 (N_1916,In_708,N_1345);
and U1917 (N_1917,In_2050,N_1284);
nor U1918 (N_1918,N_1192,N_1327);
and U1919 (N_1919,In_805,N_828);
nor U1920 (N_1920,N_1182,N_1123);
xnor U1921 (N_1921,In_2024,N_1433);
and U1922 (N_1922,In_215,In_2419);
and U1923 (N_1923,N_1254,N_1068);
and U1924 (N_1924,N_1277,In_2138);
or U1925 (N_1925,N_1487,N_1293);
and U1926 (N_1926,N_878,In_146);
nor U1927 (N_1927,N_654,N_180);
nor U1928 (N_1928,N_920,N_1051);
nand U1929 (N_1929,In_2249,N_1248);
nor U1930 (N_1930,N_1155,N_1455);
nor U1931 (N_1931,N_1324,In_1845);
nor U1932 (N_1932,In_552,N_477);
nor U1933 (N_1933,N_1383,N_509);
xnor U1934 (N_1934,N_355,N_1407);
nand U1935 (N_1935,N_1291,N_1425);
and U1936 (N_1936,N_588,N_1467);
xnor U1937 (N_1937,N_1484,N_447);
or U1938 (N_1938,In_1496,N_984);
nor U1939 (N_1939,N_1394,N_197);
and U1940 (N_1940,In_773,In_2090);
or U1941 (N_1941,N_788,N_1167);
or U1942 (N_1942,In_978,N_1446);
nand U1943 (N_1943,N_1045,N_928);
xor U1944 (N_1944,In_306,N_841);
or U1945 (N_1945,In_401,N_645);
and U1946 (N_1946,N_730,N_1249);
or U1947 (N_1947,N_1007,N_1369);
and U1948 (N_1948,In_1433,N_735);
nor U1949 (N_1949,N_1460,N_1262);
xnor U1950 (N_1950,N_1211,N_1385);
nand U1951 (N_1951,In_244,N_1274);
or U1952 (N_1952,N_1035,In_535);
or U1953 (N_1953,N_1469,N_1295);
and U1954 (N_1954,N_1322,N_1126);
and U1955 (N_1955,In_163,N_1408);
nor U1956 (N_1956,N_864,N_13);
nor U1957 (N_1957,In_1583,N_390);
xor U1958 (N_1958,N_1306,In_890);
or U1959 (N_1959,N_1361,N_893);
nor U1960 (N_1960,N_1402,In_1364);
nand U1961 (N_1961,In_2263,N_520);
nor U1962 (N_1962,N_630,N_1084);
and U1963 (N_1963,N_1379,In_128);
or U1964 (N_1964,N_1112,In_124);
and U1965 (N_1965,In_1273,N_1398);
or U1966 (N_1966,N_1239,In_321);
nand U1967 (N_1967,N_1342,N_1230);
or U1968 (N_1968,N_1474,N_1111);
nand U1969 (N_1969,N_1006,N_786);
xnor U1970 (N_1970,N_1252,N_1405);
and U1971 (N_1971,N_1234,In_2004);
xnor U1972 (N_1972,N_819,N_1263);
and U1973 (N_1973,In_1828,N_1315);
or U1974 (N_1974,N_887,N_1152);
nor U1975 (N_1975,N_1335,N_1452);
nor U1976 (N_1976,N_1027,N_1190);
nor U1977 (N_1977,In_979,N_1062);
or U1978 (N_1978,N_1145,In_755);
or U1979 (N_1979,In_2409,N_1146);
xnor U1980 (N_1980,In_2293,N_1228);
nor U1981 (N_1981,N_30,N_1193);
or U1982 (N_1982,In_389,N_1106);
and U1983 (N_1983,N_1058,N_1311);
nor U1984 (N_1984,N_342,In_1911);
or U1985 (N_1985,N_877,N_914);
and U1986 (N_1986,N_1158,In_93);
nor U1987 (N_1987,In_1922,N_1358);
or U1988 (N_1988,N_1116,N_1299);
xor U1989 (N_1989,N_330,N_626);
and U1990 (N_1990,In_457,N_968);
and U1991 (N_1991,N_814,N_1095);
nand U1992 (N_1992,In_1539,N_770);
xnor U1993 (N_1993,In_1749,N_1022);
nand U1994 (N_1994,N_603,N_651);
and U1995 (N_1995,N_1044,In_2047);
or U1996 (N_1996,N_1142,In_2341);
nor U1997 (N_1997,In_220,In_1684);
or U1998 (N_1998,N_1037,N_1059);
nand U1999 (N_1999,N_1020,N_1443);
nor U2000 (N_2000,N_1661,N_1644);
xor U2001 (N_2001,N_1600,N_1581);
nand U2002 (N_2002,N_1921,N_1586);
or U2003 (N_2003,N_1844,N_1977);
nand U2004 (N_2004,N_1668,N_1681);
xor U2005 (N_2005,N_1786,N_1673);
and U2006 (N_2006,N_1908,N_1788);
nor U2007 (N_2007,N_1958,N_1877);
and U2008 (N_2008,N_1553,N_1514);
nor U2009 (N_2009,N_1767,N_1851);
nor U2010 (N_2010,N_1738,N_1543);
nor U2011 (N_2011,N_1989,N_1963);
nand U2012 (N_2012,N_1974,N_1950);
and U2013 (N_2013,N_1972,N_1609);
nand U2014 (N_2014,N_1999,N_1973);
or U2015 (N_2015,N_1523,N_1933);
nor U2016 (N_2016,N_1755,N_1652);
or U2017 (N_2017,N_1593,N_1830);
nor U2018 (N_2018,N_1912,N_1854);
nor U2019 (N_2019,N_1682,N_1785);
nand U2020 (N_2020,N_1942,N_1686);
xor U2021 (N_2021,N_1747,N_1998);
nand U2022 (N_2022,N_1826,N_1855);
nand U2023 (N_2023,N_1874,N_1540);
xor U2024 (N_2024,N_1827,N_1640);
or U2025 (N_2025,N_1515,N_1743);
nor U2026 (N_2026,N_1551,N_1949);
and U2027 (N_2027,N_1872,N_1548);
nor U2028 (N_2028,N_1650,N_1825);
nor U2029 (N_2029,N_1662,N_1951);
or U2030 (N_2030,N_1726,N_1531);
and U2031 (N_2031,N_1649,N_1804);
or U2032 (N_2032,N_1533,N_1811);
or U2033 (N_2033,N_1539,N_1671);
or U2034 (N_2034,N_1565,N_1610);
and U2035 (N_2035,N_1544,N_1658);
xnor U2036 (N_2036,N_1653,N_1684);
xnor U2037 (N_2037,N_1805,N_1623);
and U2038 (N_2038,N_1672,N_1721);
nor U2039 (N_2039,N_1821,N_1742);
nor U2040 (N_2040,N_1729,N_1574);
nand U2041 (N_2041,N_1602,N_1667);
xnor U2042 (N_2042,N_1981,N_1841);
nand U2043 (N_2043,N_1637,N_1815);
xnor U2044 (N_2044,N_1535,N_1809);
nand U2045 (N_2045,N_1619,N_1643);
nand U2046 (N_2046,N_1787,N_1509);
nor U2047 (N_2047,N_1570,N_1969);
and U2048 (N_2048,N_1555,N_1895);
nor U2049 (N_2049,N_1597,N_1887);
nor U2050 (N_2050,N_1966,N_1703);
nor U2051 (N_2051,N_1964,N_1918);
or U2052 (N_2052,N_1939,N_1761);
or U2053 (N_2053,N_1994,N_1508);
nand U2054 (N_2054,N_1773,N_1792);
or U2055 (N_2055,N_1911,N_1756);
nor U2056 (N_2056,N_1913,N_1848);
and U2057 (N_2057,N_1707,N_1891);
nand U2058 (N_2058,N_1997,N_1930);
and U2059 (N_2059,N_1598,N_1875);
and U2060 (N_2060,N_1527,N_1893);
or U2061 (N_2061,N_1676,N_1807);
nand U2062 (N_2062,N_1639,N_1696);
and U2063 (N_2063,N_1698,N_1530);
or U2064 (N_2064,N_1611,N_1799);
and U2065 (N_2065,N_1559,N_1952);
xor U2066 (N_2066,N_1718,N_1915);
nor U2067 (N_2067,N_1724,N_1896);
and U2068 (N_2068,N_1968,N_1677);
nand U2069 (N_2069,N_1865,N_1594);
and U2070 (N_2070,N_1732,N_1769);
nand U2071 (N_2071,N_1599,N_1948);
xnor U2072 (N_2072,N_1711,N_1904);
and U2073 (N_2073,N_1754,N_1546);
nand U2074 (N_2074,N_1501,N_1596);
and U2075 (N_2075,N_1604,N_1660);
xnor U2076 (N_2076,N_1751,N_1585);
xor U2077 (N_2077,N_1556,N_1622);
and U2078 (N_2078,N_1513,N_1758);
nor U2079 (N_2079,N_1920,N_1664);
nand U2080 (N_2080,N_1840,N_1800);
and U2081 (N_2081,N_1847,N_1510);
nand U2082 (N_2082,N_1638,N_1987);
or U2083 (N_2083,N_1715,N_1860);
xor U2084 (N_2084,N_1730,N_1783);
nor U2085 (N_2085,N_1741,N_1834);
and U2086 (N_2086,N_1888,N_1823);
and U2087 (N_2087,N_1843,N_1562);
or U2088 (N_2088,N_1717,N_1691);
or U2089 (N_2089,N_1737,N_1621);
or U2090 (N_2090,N_1909,N_1852);
and U2091 (N_2091,N_1603,N_1897);
xnor U2092 (N_2092,N_1906,N_1704);
nand U2093 (N_2093,N_1947,N_1794);
nor U2094 (N_2094,N_1727,N_1745);
nand U2095 (N_2095,N_1654,N_1813);
nor U2096 (N_2096,N_1538,N_1694);
xor U2097 (N_2097,N_1608,N_1595);
or U2098 (N_2098,N_1503,N_1575);
xor U2099 (N_2099,N_1903,N_1505);
nor U2100 (N_2100,N_1746,N_1837);
nor U2101 (N_2101,N_1798,N_1749);
or U2102 (N_2102,N_1774,N_1629);
nand U2103 (N_2103,N_1763,N_1884);
nand U2104 (N_2104,N_1946,N_1701);
and U2105 (N_2105,N_1886,N_1863);
and U2106 (N_2106,N_1613,N_1725);
and U2107 (N_2107,N_1976,N_1905);
nand U2108 (N_2108,N_1615,N_1700);
nand U2109 (N_2109,N_1736,N_1557);
nor U2110 (N_2110,N_1914,N_1554);
nand U2111 (N_2111,N_1829,N_1666);
or U2112 (N_2112,N_1616,N_1552);
or U2113 (N_2113,N_1534,N_1831);
or U2114 (N_2114,N_1520,N_1642);
nand U2115 (N_2115,N_1902,N_1889);
nand U2116 (N_2116,N_1916,N_1795);
nand U2117 (N_2117,N_1541,N_1910);
nand U2118 (N_2118,N_1818,N_1858);
nor U2119 (N_2119,N_1614,N_1938);
nand U2120 (N_2120,N_1995,N_1766);
and U2121 (N_2121,N_1688,N_1960);
xor U2122 (N_2122,N_1606,N_1625);
nand U2123 (N_2123,N_1857,N_1564);
or U2124 (N_2124,N_1890,N_1945);
or U2125 (N_2125,N_1780,N_1648);
and U2126 (N_2126,N_1710,N_1862);
and U2127 (N_2127,N_1516,N_1771);
nor U2128 (N_2128,N_1706,N_1944);
or U2129 (N_2129,N_1528,N_1532);
nor U2130 (N_2130,N_1784,N_1669);
nor U2131 (N_2131,N_1776,N_1517);
and U2132 (N_2132,N_1789,N_1782);
and U2133 (N_2133,N_1733,N_1871);
nor U2134 (N_2134,N_1791,N_1983);
nor U2135 (N_2135,N_1985,N_1790);
and U2136 (N_2136,N_1931,N_1689);
nor U2137 (N_2137,N_1583,N_1859);
and U2138 (N_2138,N_1937,N_1683);
xor U2139 (N_2139,N_1744,N_1511);
nor U2140 (N_2140,N_1970,N_1752);
or U2141 (N_2141,N_1739,N_1940);
nand U2142 (N_2142,N_1880,N_1993);
and U2143 (N_2143,N_1521,N_1765);
nor U2144 (N_2144,N_1870,N_1612);
nand U2145 (N_2145,N_1592,N_1819);
and U2146 (N_2146,N_1748,N_1719);
and U2147 (N_2147,N_1569,N_1526);
nand U2148 (N_2148,N_1986,N_1576);
nor U2149 (N_2149,N_1971,N_1991);
and U2150 (N_2150,N_1646,N_1675);
or U2151 (N_2151,N_1797,N_1550);
nor U2152 (N_2152,N_1563,N_1632);
nor U2153 (N_2153,N_1839,N_1955);
or U2154 (N_2154,N_1647,N_1956);
and U2155 (N_2155,N_1892,N_1568);
xnor U2156 (N_2156,N_1656,N_1777);
and U2157 (N_2157,N_1967,N_1900);
or U2158 (N_2158,N_1731,N_1605);
nand U2159 (N_2159,N_1849,N_1779);
nand U2160 (N_2160,N_1584,N_1868);
xor U2161 (N_2161,N_1500,N_1927);
nand U2162 (N_2162,N_1984,N_1685);
and U2163 (N_2163,N_1722,N_1936);
xor U2164 (N_2164,N_1757,N_1728);
nand U2165 (N_2165,N_1567,N_1808);
or U2166 (N_2166,N_1926,N_1988);
nand U2167 (N_2167,N_1680,N_1867);
and U2168 (N_2168,N_1978,N_1573);
nand U2169 (N_2169,N_1941,N_1720);
and U2170 (N_2170,N_1735,N_1590);
nor U2171 (N_2171,N_1697,N_1547);
nor U2172 (N_2172,N_1845,N_1982);
or U2173 (N_2173,N_1634,N_1750);
nand U2174 (N_2174,N_1778,N_1641);
nand U2175 (N_2175,N_1624,N_1635);
or U2176 (N_2176,N_1572,N_1934);
nor U2177 (N_2177,N_1803,N_1655);
and U2178 (N_2178,N_1674,N_1522);
nor U2179 (N_2179,N_1992,N_1816);
and U2180 (N_2180,N_1580,N_1959);
or U2181 (N_2181,N_1762,N_1587);
nand U2182 (N_2182,N_1665,N_1558);
or U2183 (N_2183,N_1560,N_1836);
nand U2184 (N_2184,N_1607,N_1659);
xnor U2185 (N_2185,N_1549,N_1768);
or U2186 (N_2186,N_1820,N_1901);
and U2187 (N_2187,N_1702,N_1965);
and U2188 (N_2188,N_1536,N_1953);
or U2189 (N_2189,N_1705,N_1879);
xnor U2190 (N_2190,N_1627,N_1806);
nand U2191 (N_2191,N_1925,N_1631);
and U2192 (N_2192,N_1633,N_1824);
nor U2193 (N_2193,N_1861,N_1817);
and U2194 (N_2194,N_1759,N_1591);
or U2195 (N_2195,N_1853,N_1882);
xnor U2196 (N_2196,N_1917,N_1802);
and U2197 (N_2197,N_1740,N_1679);
or U2198 (N_2198,N_1626,N_1810);
and U2199 (N_2199,N_1923,N_1571);
xor U2200 (N_2200,N_1907,N_1801);
and U2201 (N_2201,N_1814,N_1876);
and U2202 (N_2202,N_1833,N_1924);
nand U2203 (N_2203,N_1502,N_1708);
or U2204 (N_2204,N_1692,N_1734);
nor U2205 (N_2205,N_1588,N_1690);
xor U2206 (N_2206,N_1699,N_1979);
nor U2207 (N_2207,N_1943,N_1772);
nor U2208 (N_2208,N_1695,N_1678);
and U2209 (N_2209,N_1663,N_1507);
nor U2210 (N_2210,N_1770,N_1620);
xor U2211 (N_2211,N_1618,N_1922);
xnor U2212 (N_2212,N_1812,N_1975);
nor U2213 (N_2213,N_1957,N_1504);
nor U2214 (N_2214,N_1822,N_1525);
or U2215 (N_2215,N_1578,N_1869);
nand U2216 (N_2216,N_1518,N_1670);
nor U2217 (N_2217,N_1873,N_1828);
and U2218 (N_2218,N_1566,N_1545);
or U2219 (N_2219,N_1561,N_1537);
nand U2220 (N_2220,N_1651,N_1506);
xnor U2221 (N_2221,N_1796,N_1935);
and U2222 (N_2222,N_1781,N_1645);
nor U2223 (N_2223,N_1885,N_1713);
or U2224 (N_2224,N_1716,N_1961);
or U2225 (N_2225,N_1932,N_1582);
or U2226 (N_2226,N_1846,N_1962);
or U2227 (N_2227,N_1577,N_1990);
or U2228 (N_2228,N_1894,N_1883);
xor U2229 (N_2229,N_1601,N_1838);
nand U2230 (N_2230,N_1709,N_1524);
or U2231 (N_2231,N_1775,N_1878);
or U2232 (N_2232,N_1793,N_1864);
or U2233 (N_2233,N_1881,N_1589);
or U2234 (N_2234,N_1723,N_1687);
nand U2235 (N_2235,N_1919,N_1519);
nand U2236 (N_2236,N_1712,N_1929);
or U2237 (N_2237,N_1542,N_1928);
nor U2238 (N_2238,N_1898,N_1764);
or U2239 (N_2239,N_1529,N_1856);
nor U2240 (N_2240,N_1714,N_1832);
nand U2241 (N_2241,N_1980,N_1996);
or U2242 (N_2242,N_1657,N_1617);
nand U2243 (N_2243,N_1899,N_1842);
xnor U2244 (N_2244,N_1835,N_1636);
and U2245 (N_2245,N_1512,N_1850);
nand U2246 (N_2246,N_1954,N_1630);
nor U2247 (N_2247,N_1866,N_1579);
nand U2248 (N_2248,N_1760,N_1693);
xor U2249 (N_2249,N_1628,N_1753);
and U2250 (N_2250,N_1820,N_1858);
nand U2251 (N_2251,N_1603,N_1780);
and U2252 (N_2252,N_1540,N_1951);
or U2253 (N_2253,N_1641,N_1616);
or U2254 (N_2254,N_1651,N_1892);
nand U2255 (N_2255,N_1734,N_1605);
nor U2256 (N_2256,N_1943,N_1680);
nor U2257 (N_2257,N_1548,N_1772);
and U2258 (N_2258,N_1820,N_1539);
and U2259 (N_2259,N_1509,N_1676);
and U2260 (N_2260,N_1951,N_1536);
nor U2261 (N_2261,N_1689,N_1996);
and U2262 (N_2262,N_1582,N_1757);
xnor U2263 (N_2263,N_1559,N_1921);
nor U2264 (N_2264,N_1604,N_1626);
xor U2265 (N_2265,N_1900,N_1934);
nor U2266 (N_2266,N_1732,N_1697);
nand U2267 (N_2267,N_1612,N_1969);
xnor U2268 (N_2268,N_1809,N_1672);
nor U2269 (N_2269,N_1745,N_1586);
nor U2270 (N_2270,N_1655,N_1690);
nand U2271 (N_2271,N_1671,N_1997);
nand U2272 (N_2272,N_1593,N_1534);
and U2273 (N_2273,N_1588,N_1838);
nor U2274 (N_2274,N_1647,N_1937);
nand U2275 (N_2275,N_1792,N_1945);
and U2276 (N_2276,N_1609,N_1981);
nor U2277 (N_2277,N_1900,N_1595);
or U2278 (N_2278,N_1602,N_1587);
or U2279 (N_2279,N_1754,N_1922);
nand U2280 (N_2280,N_1861,N_1957);
or U2281 (N_2281,N_1863,N_1685);
nor U2282 (N_2282,N_1692,N_1965);
and U2283 (N_2283,N_1530,N_1881);
nand U2284 (N_2284,N_1774,N_1737);
nand U2285 (N_2285,N_1684,N_1843);
or U2286 (N_2286,N_1521,N_1796);
nor U2287 (N_2287,N_1568,N_1939);
and U2288 (N_2288,N_1501,N_1923);
nor U2289 (N_2289,N_1527,N_1740);
or U2290 (N_2290,N_1962,N_1704);
nand U2291 (N_2291,N_1562,N_1951);
or U2292 (N_2292,N_1722,N_1643);
nor U2293 (N_2293,N_1802,N_1616);
and U2294 (N_2294,N_1532,N_1956);
nor U2295 (N_2295,N_1888,N_1669);
or U2296 (N_2296,N_1988,N_1909);
nand U2297 (N_2297,N_1714,N_1608);
nor U2298 (N_2298,N_1503,N_1552);
nor U2299 (N_2299,N_1731,N_1519);
and U2300 (N_2300,N_1834,N_1843);
and U2301 (N_2301,N_1983,N_1721);
nand U2302 (N_2302,N_1864,N_1884);
nand U2303 (N_2303,N_1506,N_1805);
nand U2304 (N_2304,N_1811,N_1591);
nand U2305 (N_2305,N_1953,N_1837);
and U2306 (N_2306,N_1861,N_1859);
nor U2307 (N_2307,N_1882,N_1942);
nor U2308 (N_2308,N_1692,N_1511);
nor U2309 (N_2309,N_1837,N_1668);
or U2310 (N_2310,N_1719,N_1760);
and U2311 (N_2311,N_1890,N_1624);
nor U2312 (N_2312,N_1911,N_1877);
nand U2313 (N_2313,N_1580,N_1906);
and U2314 (N_2314,N_1620,N_1928);
and U2315 (N_2315,N_1536,N_1967);
and U2316 (N_2316,N_1674,N_1510);
nand U2317 (N_2317,N_1899,N_1915);
and U2318 (N_2318,N_1883,N_1759);
nor U2319 (N_2319,N_1897,N_1857);
and U2320 (N_2320,N_1975,N_1995);
nor U2321 (N_2321,N_1782,N_1799);
nand U2322 (N_2322,N_1607,N_1557);
and U2323 (N_2323,N_1876,N_1508);
or U2324 (N_2324,N_1942,N_1944);
nor U2325 (N_2325,N_1768,N_1641);
nor U2326 (N_2326,N_1678,N_1921);
nand U2327 (N_2327,N_1742,N_1776);
or U2328 (N_2328,N_1759,N_1985);
or U2329 (N_2329,N_1917,N_1853);
or U2330 (N_2330,N_1895,N_1530);
nor U2331 (N_2331,N_1757,N_1797);
and U2332 (N_2332,N_1942,N_1501);
or U2333 (N_2333,N_1544,N_1566);
xor U2334 (N_2334,N_1559,N_1978);
and U2335 (N_2335,N_1650,N_1518);
and U2336 (N_2336,N_1903,N_1616);
or U2337 (N_2337,N_1647,N_1611);
and U2338 (N_2338,N_1533,N_1685);
nand U2339 (N_2339,N_1610,N_1910);
nor U2340 (N_2340,N_1634,N_1823);
nor U2341 (N_2341,N_1532,N_1694);
or U2342 (N_2342,N_1720,N_1844);
xor U2343 (N_2343,N_1987,N_1997);
nor U2344 (N_2344,N_1552,N_1991);
nor U2345 (N_2345,N_1937,N_1668);
and U2346 (N_2346,N_1687,N_1767);
nand U2347 (N_2347,N_1607,N_1792);
or U2348 (N_2348,N_1825,N_1681);
xor U2349 (N_2349,N_1976,N_1851);
nor U2350 (N_2350,N_1631,N_1950);
or U2351 (N_2351,N_1680,N_1995);
xnor U2352 (N_2352,N_1554,N_1885);
nand U2353 (N_2353,N_1968,N_1935);
xnor U2354 (N_2354,N_1811,N_1858);
nor U2355 (N_2355,N_1600,N_1974);
or U2356 (N_2356,N_1866,N_1945);
nor U2357 (N_2357,N_1579,N_1829);
xor U2358 (N_2358,N_1992,N_1521);
nor U2359 (N_2359,N_1723,N_1640);
nand U2360 (N_2360,N_1539,N_1509);
and U2361 (N_2361,N_1777,N_1725);
or U2362 (N_2362,N_1787,N_1608);
nor U2363 (N_2363,N_1732,N_1510);
nand U2364 (N_2364,N_1746,N_1761);
nor U2365 (N_2365,N_1670,N_1899);
and U2366 (N_2366,N_1730,N_1732);
nand U2367 (N_2367,N_1731,N_1667);
or U2368 (N_2368,N_1999,N_1786);
nand U2369 (N_2369,N_1877,N_1861);
xnor U2370 (N_2370,N_1653,N_1910);
xnor U2371 (N_2371,N_1834,N_1759);
nand U2372 (N_2372,N_1608,N_1848);
and U2373 (N_2373,N_1617,N_1537);
xor U2374 (N_2374,N_1544,N_1826);
or U2375 (N_2375,N_1637,N_1686);
xor U2376 (N_2376,N_1520,N_1995);
and U2377 (N_2377,N_1879,N_1865);
xor U2378 (N_2378,N_1747,N_1698);
nand U2379 (N_2379,N_1564,N_1614);
nor U2380 (N_2380,N_1898,N_1817);
nor U2381 (N_2381,N_1618,N_1566);
nor U2382 (N_2382,N_1515,N_1552);
nand U2383 (N_2383,N_1642,N_1838);
xor U2384 (N_2384,N_1545,N_1726);
or U2385 (N_2385,N_1603,N_1941);
nand U2386 (N_2386,N_1635,N_1520);
and U2387 (N_2387,N_1925,N_1986);
nand U2388 (N_2388,N_1543,N_1523);
nor U2389 (N_2389,N_1569,N_1508);
nor U2390 (N_2390,N_1889,N_1548);
nor U2391 (N_2391,N_1585,N_1503);
xor U2392 (N_2392,N_1524,N_1718);
nand U2393 (N_2393,N_1556,N_1584);
nand U2394 (N_2394,N_1962,N_1926);
or U2395 (N_2395,N_1771,N_1675);
xor U2396 (N_2396,N_1652,N_1570);
or U2397 (N_2397,N_1697,N_1955);
and U2398 (N_2398,N_1589,N_1861);
or U2399 (N_2399,N_1790,N_1704);
nand U2400 (N_2400,N_1737,N_1888);
or U2401 (N_2401,N_1541,N_1561);
nand U2402 (N_2402,N_1615,N_1565);
or U2403 (N_2403,N_1871,N_1724);
nor U2404 (N_2404,N_1707,N_1566);
nand U2405 (N_2405,N_1619,N_1801);
nor U2406 (N_2406,N_1789,N_1992);
nand U2407 (N_2407,N_1960,N_1913);
and U2408 (N_2408,N_1593,N_1846);
nor U2409 (N_2409,N_1651,N_1642);
nand U2410 (N_2410,N_1841,N_1893);
and U2411 (N_2411,N_1503,N_1508);
xnor U2412 (N_2412,N_1690,N_1570);
and U2413 (N_2413,N_1623,N_1881);
nor U2414 (N_2414,N_1559,N_1608);
or U2415 (N_2415,N_1967,N_1987);
nor U2416 (N_2416,N_1974,N_1860);
and U2417 (N_2417,N_1528,N_1762);
nand U2418 (N_2418,N_1806,N_1652);
and U2419 (N_2419,N_1867,N_1909);
and U2420 (N_2420,N_1743,N_1906);
or U2421 (N_2421,N_1867,N_1578);
nand U2422 (N_2422,N_1907,N_1553);
or U2423 (N_2423,N_1605,N_1602);
or U2424 (N_2424,N_1664,N_1834);
and U2425 (N_2425,N_1920,N_1621);
nand U2426 (N_2426,N_1672,N_1817);
nor U2427 (N_2427,N_1528,N_1803);
and U2428 (N_2428,N_1630,N_1616);
nand U2429 (N_2429,N_1752,N_1885);
or U2430 (N_2430,N_1538,N_1898);
xnor U2431 (N_2431,N_1538,N_1747);
and U2432 (N_2432,N_1605,N_1554);
nand U2433 (N_2433,N_1910,N_1792);
nand U2434 (N_2434,N_1767,N_1804);
or U2435 (N_2435,N_1771,N_1839);
and U2436 (N_2436,N_1608,N_1505);
and U2437 (N_2437,N_1730,N_1864);
nor U2438 (N_2438,N_1642,N_1595);
or U2439 (N_2439,N_1652,N_1669);
nor U2440 (N_2440,N_1729,N_1840);
nand U2441 (N_2441,N_1834,N_1936);
and U2442 (N_2442,N_1516,N_1714);
nand U2443 (N_2443,N_1619,N_1796);
nor U2444 (N_2444,N_1902,N_1717);
nor U2445 (N_2445,N_1861,N_1764);
or U2446 (N_2446,N_1741,N_1570);
nor U2447 (N_2447,N_1501,N_1591);
nand U2448 (N_2448,N_1995,N_1827);
or U2449 (N_2449,N_1840,N_1609);
nor U2450 (N_2450,N_1534,N_1974);
nand U2451 (N_2451,N_1696,N_1947);
or U2452 (N_2452,N_1591,N_1835);
or U2453 (N_2453,N_1587,N_1661);
nor U2454 (N_2454,N_1820,N_1735);
nor U2455 (N_2455,N_1553,N_1632);
nand U2456 (N_2456,N_1786,N_1853);
or U2457 (N_2457,N_1650,N_1679);
or U2458 (N_2458,N_1551,N_1842);
nor U2459 (N_2459,N_1765,N_1740);
nand U2460 (N_2460,N_1564,N_1938);
or U2461 (N_2461,N_1796,N_1520);
and U2462 (N_2462,N_1920,N_1834);
xor U2463 (N_2463,N_1795,N_1836);
nand U2464 (N_2464,N_1930,N_1848);
or U2465 (N_2465,N_1546,N_1507);
or U2466 (N_2466,N_1594,N_1906);
xor U2467 (N_2467,N_1524,N_1589);
and U2468 (N_2468,N_1618,N_1854);
nor U2469 (N_2469,N_1859,N_1846);
or U2470 (N_2470,N_1697,N_1535);
xnor U2471 (N_2471,N_1574,N_1792);
xor U2472 (N_2472,N_1764,N_1935);
nand U2473 (N_2473,N_1562,N_1762);
nor U2474 (N_2474,N_1605,N_1624);
and U2475 (N_2475,N_1782,N_1734);
or U2476 (N_2476,N_1508,N_1835);
or U2477 (N_2477,N_1592,N_1594);
nand U2478 (N_2478,N_1607,N_1520);
or U2479 (N_2479,N_1968,N_1885);
and U2480 (N_2480,N_1806,N_1755);
nand U2481 (N_2481,N_1957,N_1623);
nand U2482 (N_2482,N_1955,N_1706);
nor U2483 (N_2483,N_1560,N_1749);
or U2484 (N_2484,N_1643,N_1784);
and U2485 (N_2485,N_1944,N_1859);
nor U2486 (N_2486,N_1847,N_1949);
and U2487 (N_2487,N_1888,N_1537);
nand U2488 (N_2488,N_1955,N_1787);
xnor U2489 (N_2489,N_1810,N_1950);
or U2490 (N_2490,N_1551,N_1917);
nor U2491 (N_2491,N_1688,N_1824);
nor U2492 (N_2492,N_1608,N_1886);
xor U2493 (N_2493,N_1758,N_1725);
or U2494 (N_2494,N_1826,N_1561);
nor U2495 (N_2495,N_1818,N_1823);
and U2496 (N_2496,N_1665,N_1639);
xor U2497 (N_2497,N_1838,N_1830);
nor U2498 (N_2498,N_1562,N_1653);
and U2499 (N_2499,N_1927,N_1572);
or U2500 (N_2500,N_2164,N_2006);
nand U2501 (N_2501,N_2173,N_2382);
nor U2502 (N_2502,N_2187,N_2453);
or U2503 (N_2503,N_2032,N_2262);
and U2504 (N_2504,N_2348,N_2116);
or U2505 (N_2505,N_2364,N_2291);
and U2506 (N_2506,N_2148,N_2117);
nor U2507 (N_2507,N_2295,N_2473);
and U2508 (N_2508,N_2264,N_2228);
nand U2509 (N_2509,N_2410,N_2374);
nor U2510 (N_2510,N_2317,N_2195);
and U2511 (N_2511,N_2376,N_2122);
nand U2512 (N_2512,N_2071,N_2024);
nand U2513 (N_2513,N_2045,N_2238);
or U2514 (N_2514,N_2324,N_2476);
nand U2515 (N_2515,N_2466,N_2408);
or U2516 (N_2516,N_2460,N_2049);
nor U2517 (N_2517,N_2199,N_2176);
and U2518 (N_2518,N_2411,N_2151);
nor U2519 (N_2519,N_2048,N_2477);
nand U2520 (N_2520,N_2475,N_2258);
nor U2521 (N_2521,N_2146,N_2290);
and U2522 (N_2522,N_2426,N_2254);
or U2523 (N_2523,N_2125,N_2311);
nand U2524 (N_2524,N_2456,N_2085);
and U2525 (N_2525,N_2300,N_2177);
and U2526 (N_2526,N_2489,N_2380);
nand U2527 (N_2527,N_2040,N_2278);
nor U2528 (N_2528,N_2480,N_2096);
nand U2529 (N_2529,N_2183,N_2298);
nor U2530 (N_2530,N_2225,N_2230);
and U2531 (N_2531,N_2129,N_2232);
or U2532 (N_2532,N_2497,N_2201);
or U2533 (N_2533,N_2181,N_2345);
and U2534 (N_2534,N_2079,N_2197);
nand U2535 (N_2535,N_2434,N_2089);
nor U2536 (N_2536,N_2458,N_2236);
nor U2537 (N_2537,N_2144,N_2128);
or U2538 (N_2538,N_2483,N_2297);
or U2539 (N_2539,N_2482,N_2074);
or U2540 (N_2540,N_2373,N_2288);
nor U2541 (N_2541,N_2447,N_2438);
nand U2542 (N_2542,N_2240,N_2429);
and U2543 (N_2543,N_2108,N_2219);
nor U2544 (N_2544,N_2154,N_2479);
and U2545 (N_2545,N_2007,N_2166);
or U2546 (N_2546,N_2312,N_2461);
and U2547 (N_2547,N_2014,N_2267);
and U2548 (N_2548,N_2207,N_2033);
nand U2549 (N_2549,N_2051,N_2351);
xor U2550 (N_2550,N_2015,N_2491);
nand U2551 (N_2551,N_2140,N_2338);
or U2552 (N_2552,N_2104,N_2239);
or U2553 (N_2553,N_2004,N_2194);
and U2554 (N_2554,N_2444,N_2319);
xnor U2555 (N_2555,N_2145,N_2289);
or U2556 (N_2556,N_2180,N_2110);
or U2557 (N_2557,N_2242,N_2328);
or U2558 (N_2558,N_2066,N_2182);
nand U2559 (N_2559,N_2082,N_2214);
nand U2560 (N_2560,N_2155,N_2213);
nor U2561 (N_2561,N_2495,N_2088);
nor U2562 (N_2562,N_2494,N_2001);
or U2563 (N_2563,N_2406,N_2332);
and U2564 (N_2564,N_2440,N_2484);
or U2565 (N_2565,N_2087,N_2266);
and U2566 (N_2566,N_2205,N_2400);
or U2567 (N_2567,N_2398,N_2231);
or U2568 (N_2568,N_2170,N_2035);
or U2569 (N_2569,N_2292,N_2252);
nand U2570 (N_2570,N_2356,N_2042);
and U2571 (N_2571,N_2083,N_2283);
nand U2572 (N_2572,N_2314,N_2198);
nand U2573 (N_2573,N_2204,N_2243);
and U2574 (N_2574,N_2315,N_2130);
nand U2575 (N_2575,N_2309,N_2118);
or U2576 (N_2576,N_2255,N_2127);
nor U2577 (N_2577,N_2190,N_2404);
and U2578 (N_2578,N_2299,N_2249);
nand U2579 (N_2579,N_2422,N_2276);
and U2580 (N_2580,N_2123,N_2301);
or U2581 (N_2581,N_2184,N_2216);
and U2582 (N_2582,N_2103,N_2257);
or U2583 (N_2583,N_2244,N_2282);
nand U2584 (N_2584,N_2003,N_2462);
nor U2585 (N_2585,N_2072,N_2386);
nand U2586 (N_2586,N_2063,N_2346);
and U2587 (N_2587,N_2029,N_2133);
nand U2588 (N_2588,N_2080,N_2407);
nand U2589 (N_2589,N_2394,N_2392);
nor U2590 (N_2590,N_2367,N_2149);
nand U2591 (N_2591,N_2165,N_2174);
nor U2592 (N_2592,N_2158,N_2016);
or U2593 (N_2593,N_2384,N_2223);
xor U2594 (N_2594,N_2368,N_2416);
nor U2595 (N_2595,N_2284,N_2124);
nand U2596 (N_2596,N_2126,N_2270);
or U2597 (N_2597,N_2454,N_2058);
nor U2598 (N_2598,N_2038,N_2263);
nand U2599 (N_2599,N_2078,N_2469);
and U2600 (N_2600,N_2488,N_2415);
nor U2601 (N_2601,N_2353,N_2008);
and U2602 (N_2602,N_2340,N_2421);
nor U2603 (N_2603,N_2452,N_2136);
or U2604 (N_2604,N_2030,N_2269);
nand U2605 (N_2605,N_2344,N_2372);
nand U2606 (N_2606,N_2331,N_2409);
nor U2607 (N_2607,N_2305,N_2419);
or U2608 (N_2608,N_2457,N_2060);
or U2609 (N_2609,N_2451,N_2428);
or U2610 (N_2610,N_2112,N_2047);
and U2611 (N_2611,N_2009,N_2355);
nand U2612 (N_2612,N_2044,N_2385);
or U2613 (N_2613,N_2499,N_2342);
or U2614 (N_2614,N_2059,N_2043);
nor U2615 (N_2615,N_2221,N_2437);
nor U2616 (N_2616,N_2293,N_2381);
nand U2617 (N_2617,N_2468,N_2361);
nor U2618 (N_2618,N_2261,N_2339);
and U2619 (N_2619,N_2101,N_2478);
nand U2620 (N_2620,N_2463,N_2389);
nand U2621 (N_2621,N_2234,N_2152);
xor U2622 (N_2622,N_2253,N_2191);
and U2623 (N_2623,N_2193,N_2308);
and U2624 (N_2624,N_2241,N_2397);
or U2625 (N_2625,N_2106,N_2222);
and U2626 (N_2626,N_2196,N_2259);
and U2627 (N_2627,N_2435,N_2220);
and U2628 (N_2628,N_2304,N_2443);
nand U2629 (N_2629,N_2153,N_2189);
or U2630 (N_2630,N_2025,N_2286);
nand U2631 (N_2631,N_2011,N_2357);
nand U2632 (N_2632,N_2401,N_2012);
and U2633 (N_2633,N_2498,N_2465);
and U2634 (N_2634,N_2450,N_2327);
xnor U2635 (N_2635,N_2209,N_2274);
or U2636 (N_2636,N_2105,N_2280);
and U2637 (N_2637,N_2379,N_2020);
xnor U2638 (N_2638,N_2086,N_2065);
or U2639 (N_2639,N_2248,N_2455);
and U2640 (N_2640,N_2472,N_2141);
and U2641 (N_2641,N_2208,N_2203);
and U2642 (N_2642,N_2121,N_2098);
nand U2643 (N_2643,N_2251,N_2343);
nand U2644 (N_2644,N_2159,N_2211);
or U2645 (N_2645,N_2359,N_2417);
xor U2646 (N_2646,N_2431,N_2028);
nor U2647 (N_2647,N_2052,N_2387);
and U2648 (N_2648,N_2474,N_2002);
and U2649 (N_2649,N_2492,N_2057);
and U2650 (N_2650,N_2420,N_2202);
xnor U2651 (N_2651,N_2362,N_2320);
nor U2652 (N_2652,N_2306,N_2256);
nor U2653 (N_2653,N_2075,N_2336);
xnor U2654 (N_2654,N_2062,N_2206);
nor U2655 (N_2655,N_2427,N_2150);
nor U2656 (N_2656,N_2446,N_2172);
nand U2657 (N_2657,N_2493,N_2313);
nor U2658 (N_2658,N_2296,N_2081);
or U2659 (N_2659,N_2358,N_2247);
nand U2660 (N_2660,N_2388,N_2227);
nand U2661 (N_2661,N_2341,N_2084);
nand U2662 (N_2662,N_2390,N_2212);
nor U2663 (N_2663,N_2349,N_2056);
and U2664 (N_2664,N_2246,N_2114);
or U2665 (N_2665,N_2325,N_2160);
nand U2666 (N_2666,N_2281,N_2131);
nand U2667 (N_2667,N_2424,N_2200);
and U2668 (N_2668,N_2157,N_2099);
nor U2669 (N_2669,N_2217,N_2161);
nand U2670 (N_2670,N_2113,N_2470);
nor U2671 (N_2671,N_2448,N_2090);
xor U2672 (N_2672,N_2352,N_2186);
nand U2673 (N_2673,N_2277,N_2396);
nand U2674 (N_2674,N_2323,N_2371);
or U2675 (N_2675,N_2233,N_2021);
nor U2676 (N_2676,N_2226,N_2005);
xnor U2677 (N_2677,N_2097,N_2490);
nor U2678 (N_2678,N_2162,N_2070);
and U2679 (N_2679,N_2414,N_2142);
nor U2680 (N_2680,N_2360,N_2210);
and U2681 (N_2681,N_2055,N_2237);
nand U2682 (N_2682,N_2393,N_2445);
and U2683 (N_2683,N_2279,N_2481);
and U2684 (N_2684,N_2178,N_2464);
or U2685 (N_2685,N_2265,N_2436);
or U2686 (N_2686,N_2013,N_2046);
and U2687 (N_2687,N_2095,N_2039);
xor U2688 (N_2688,N_2111,N_2449);
nor U2689 (N_2689,N_2432,N_2412);
nand U2690 (N_2690,N_2287,N_2413);
and U2691 (N_2691,N_2037,N_2271);
and U2692 (N_2692,N_2350,N_2022);
nand U2693 (N_2693,N_2076,N_2459);
and U2694 (N_2694,N_2260,N_2303);
and U2695 (N_2695,N_2307,N_2496);
nor U2696 (N_2696,N_2215,N_2322);
nand U2697 (N_2697,N_2224,N_2363);
and U2698 (N_2698,N_2378,N_2017);
and U2699 (N_2699,N_2068,N_2041);
or U2700 (N_2700,N_2418,N_2018);
or U2701 (N_2701,N_2132,N_2143);
and U2702 (N_2702,N_2091,N_2405);
xnor U2703 (N_2703,N_2485,N_2334);
xor U2704 (N_2704,N_2139,N_2115);
and U2705 (N_2705,N_2235,N_2337);
and U2706 (N_2706,N_2391,N_2329);
nand U2707 (N_2707,N_2333,N_2192);
and U2708 (N_2708,N_2171,N_2441);
or U2709 (N_2709,N_2377,N_2107);
or U2710 (N_2710,N_2169,N_2423);
nor U2711 (N_2711,N_2369,N_2383);
and U2712 (N_2712,N_2486,N_2275);
nor U2713 (N_2713,N_2402,N_2294);
nor U2714 (N_2714,N_2010,N_2053);
and U2715 (N_2715,N_2250,N_2093);
nor U2716 (N_2716,N_2147,N_2302);
xnor U2717 (N_2717,N_2285,N_2326);
nand U2718 (N_2718,N_2268,N_2365);
nand U2719 (N_2719,N_2347,N_2069);
and U2720 (N_2720,N_2188,N_2138);
nor U2721 (N_2721,N_2433,N_2054);
nand U2722 (N_2722,N_2036,N_2467);
nor U2723 (N_2723,N_2094,N_2120);
nand U2724 (N_2724,N_2354,N_2442);
and U2725 (N_2725,N_2439,N_2077);
or U2726 (N_2726,N_2487,N_2370);
nand U2727 (N_2727,N_2471,N_2027);
nand U2728 (N_2728,N_2403,N_2034);
and U2729 (N_2729,N_2310,N_2067);
and U2730 (N_2730,N_2167,N_2061);
nand U2731 (N_2731,N_2318,N_2073);
or U2732 (N_2732,N_2273,N_2023);
nand U2733 (N_2733,N_2272,N_2330);
or U2734 (N_2734,N_2395,N_2000);
nor U2735 (N_2735,N_2119,N_2335);
and U2736 (N_2736,N_2175,N_2399);
or U2737 (N_2737,N_2026,N_2218);
and U2738 (N_2738,N_2316,N_2245);
nand U2739 (N_2739,N_2163,N_2179);
or U2740 (N_2740,N_2425,N_2019);
and U2741 (N_2741,N_2229,N_2100);
or U2742 (N_2742,N_2135,N_2064);
nor U2743 (N_2743,N_2092,N_2321);
nand U2744 (N_2744,N_2050,N_2156);
nand U2745 (N_2745,N_2137,N_2102);
nand U2746 (N_2746,N_2430,N_2375);
or U2747 (N_2747,N_2134,N_2109);
xnor U2748 (N_2748,N_2168,N_2031);
nor U2749 (N_2749,N_2185,N_2366);
nor U2750 (N_2750,N_2200,N_2458);
nand U2751 (N_2751,N_2098,N_2357);
nand U2752 (N_2752,N_2254,N_2260);
and U2753 (N_2753,N_2492,N_2010);
nand U2754 (N_2754,N_2492,N_2119);
nand U2755 (N_2755,N_2362,N_2296);
nand U2756 (N_2756,N_2022,N_2433);
and U2757 (N_2757,N_2046,N_2244);
or U2758 (N_2758,N_2233,N_2438);
or U2759 (N_2759,N_2294,N_2499);
and U2760 (N_2760,N_2473,N_2411);
or U2761 (N_2761,N_2328,N_2417);
or U2762 (N_2762,N_2353,N_2098);
or U2763 (N_2763,N_2336,N_2341);
xor U2764 (N_2764,N_2086,N_2344);
and U2765 (N_2765,N_2246,N_2037);
nand U2766 (N_2766,N_2156,N_2023);
nand U2767 (N_2767,N_2492,N_2273);
or U2768 (N_2768,N_2275,N_2439);
nand U2769 (N_2769,N_2385,N_2342);
nand U2770 (N_2770,N_2263,N_2183);
xor U2771 (N_2771,N_2309,N_2488);
and U2772 (N_2772,N_2381,N_2352);
xnor U2773 (N_2773,N_2480,N_2369);
nand U2774 (N_2774,N_2358,N_2465);
nor U2775 (N_2775,N_2414,N_2492);
nand U2776 (N_2776,N_2192,N_2325);
nor U2777 (N_2777,N_2176,N_2203);
or U2778 (N_2778,N_2300,N_2393);
or U2779 (N_2779,N_2290,N_2283);
nor U2780 (N_2780,N_2145,N_2293);
and U2781 (N_2781,N_2131,N_2396);
nor U2782 (N_2782,N_2467,N_2140);
xnor U2783 (N_2783,N_2270,N_2279);
and U2784 (N_2784,N_2311,N_2417);
xnor U2785 (N_2785,N_2358,N_2184);
or U2786 (N_2786,N_2112,N_2448);
nand U2787 (N_2787,N_2005,N_2432);
and U2788 (N_2788,N_2193,N_2125);
and U2789 (N_2789,N_2070,N_2442);
and U2790 (N_2790,N_2144,N_2194);
xor U2791 (N_2791,N_2497,N_2275);
nand U2792 (N_2792,N_2089,N_2361);
and U2793 (N_2793,N_2263,N_2339);
nor U2794 (N_2794,N_2303,N_2343);
or U2795 (N_2795,N_2325,N_2174);
or U2796 (N_2796,N_2255,N_2238);
nor U2797 (N_2797,N_2480,N_2234);
or U2798 (N_2798,N_2172,N_2235);
or U2799 (N_2799,N_2338,N_2414);
or U2800 (N_2800,N_2200,N_2496);
and U2801 (N_2801,N_2276,N_2147);
and U2802 (N_2802,N_2220,N_2349);
nor U2803 (N_2803,N_2138,N_2003);
xor U2804 (N_2804,N_2453,N_2450);
or U2805 (N_2805,N_2410,N_2167);
or U2806 (N_2806,N_2216,N_2350);
or U2807 (N_2807,N_2239,N_2281);
or U2808 (N_2808,N_2065,N_2257);
and U2809 (N_2809,N_2495,N_2207);
and U2810 (N_2810,N_2448,N_2492);
nand U2811 (N_2811,N_2220,N_2403);
or U2812 (N_2812,N_2090,N_2364);
xor U2813 (N_2813,N_2156,N_2315);
nand U2814 (N_2814,N_2354,N_2071);
nand U2815 (N_2815,N_2466,N_2305);
or U2816 (N_2816,N_2444,N_2032);
nand U2817 (N_2817,N_2369,N_2387);
and U2818 (N_2818,N_2062,N_2161);
and U2819 (N_2819,N_2336,N_2043);
and U2820 (N_2820,N_2200,N_2419);
or U2821 (N_2821,N_2300,N_2022);
nor U2822 (N_2822,N_2397,N_2040);
or U2823 (N_2823,N_2400,N_2313);
nor U2824 (N_2824,N_2113,N_2444);
nor U2825 (N_2825,N_2055,N_2409);
nand U2826 (N_2826,N_2248,N_2087);
nor U2827 (N_2827,N_2304,N_2021);
or U2828 (N_2828,N_2388,N_2284);
nor U2829 (N_2829,N_2131,N_2211);
nand U2830 (N_2830,N_2445,N_2084);
nor U2831 (N_2831,N_2126,N_2288);
nor U2832 (N_2832,N_2264,N_2176);
nor U2833 (N_2833,N_2165,N_2340);
or U2834 (N_2834,N_2470,N_2090);
or U2835 (N_2835,N_2267,N_2473);
nand U2836 (N_2836,N_2336,N_2212);
and U2837 (N_2837,N_2437,N_2496);
nor U2838 (N_2838,N_2221,N_2050);
nor U2839 (N_2839,N_2084,N_2294);
or U2840 (N_2840,N_2341,N_2246);
nand U2841 (N_2841,N_2313,N_2232);
and U2842 (N_2842,N_2213,N_2488);
nor U2843 (N_2843,N_2330,N_2154);
and U2844 (N_2844,N_2443,N_2378);
xnor U2845 (N_2845,N_2015,N_2230);
or U2846 (N_2846,N_2369,N_2304);
and U2847 (N_2847,N_2175,N_2429);
and U2848 (N_2848,N_2148,N_2210);
or U2849 (N_2849,N_2299,N_2379);
nor U2850 (N_2850,N_2172,N_2194);
nand U2851 (N_2851,N_2146,N_2071);
nor U2852 (N_2852,N_2093,N_2193);
nor U2853 (N_2853,N_2438,N_2269);
xnor U2854 (N_2854,N_2158,N_2090);
nor U2855 (N_2855,N_2143,N_2221);
nand U2856 (N_2856,N_2067,N_2313);
nand U2857 (N_2857,N_2118,N_2440);
nor U2858 (N_2858,N_2036,N_2251);
or U2859 (N_2859,N_2212,N_2061);
or U2860 (N_2860,N_2194,N_2497);
nor U2861 (N_2861,N_2436,N_2139);
and U2862 (N_2862,N_2223,N_2304);
and U2863 (N_2863,N_2011,N_2438);
and U2864 (N_2864,N_2119,N_2493);
nand U2865 (N_2865,N_2018,N_2064);
xnor U2866 (N_2866,N_2124,N_2446);
or U2867 (N_2867,N_2328,N_2061);
nor U2868 (N_2868,N_2304,N_2350);
and U2869 (N_2869,N_2477,N_2441);
or U2870 (N_2870,N_2145,N_2339);
nand U2871 (N_2871,N_2061,N_2321);
nor U2872 (N_2872,N_2442,N_2117);
xnor U2873 (N_2873,N_2321,N_2369);
nand U2874 (N_2874,N_2158,N_2357);
and U2875 (N_2875,N_2229,N_2464);
nand U2876 (N_2876,N_2025,N_2007);
nor U2877 (N_2877,N_2095,N_2142);
and U2878 (N_2878,N_2261,N_2359);
xnor U2879 (N_2879,N_2374,N_2205);
xnor U2880 (N_2880,N_2422,N_2167);
nor U2881 (N_2881,N_2268,N_2100);
xor U2882 (N_2882,N_2294,N_2040);
nor U2883 (N_2883,N_2047,N_2129);
xor U2884 (N_2884,N_2148,N_2084);
and U2885 (N_2885,N_2006,N_2335);
nand U2886 (N_2886,N_2339,N_2404);
and U2887 (N_2887,N_2078,N_2040);
xnor U2888 (N_2888,N_2414,N_2346);
nand U2889 (N_2889,N_2348,N_2431);
or U2890 (N_2890,N_2207,N_2187);
nor U2891 (N_2891,N_2145,N_2435);
nand U2892 (N_2892,N_2066,N_2355);
xnor U2893 (N_2893,N_2438,N_2189);
and U2894 (N_2894,N_2181,N_2330);
nor U2895 (N_2895,N_2086,N_2135);
or U2896 (N_2896,N_2119,N_2025);
nor U2897 (N_2897,N_2426,N_2265);
nand U2898 (N_2898,N_2338,N_2335);
or U2899 (N_2899,N_2326,N_2124);
nor U2900 (N_2900,N_2168,N_2422);
nand U2901 (N_2901,N_2042,N_2283);
or U2902 (N_2902,N_2366,N_2245);
nand U2903 (N_2903,N_2078,N_2071);
nand U2904 (N_2904,N_2323,N_2408);
nor U2905 (N_2905,N_2334,N_2299);
or U2906 (N_2906,N_2474,N_2362);
or U2907 (N_2907,N_2065,N_2095);
or U2908 (N_2908,N_2475,N_2345);
and U2909 (N_2909,N_2010,N_2094);
nor U2910 (N_2910,N_2400,N_2263);
or U2911 (N_2911,N_2041,N_2226);
nor U2912 (N_2912,N_2193,N_2406);
and U2913 (N_2913,N_2177,N_2081);
nand U2914 (N_2914,N_2247,N_2130);
nor U2915 (N_2915,N_2439,N_2196);
and U2916 (N_2916,N_2391,N_2106);
xnor U2917 (N_2917,N_2144,N_2089);
and U2918 (N_2918,N_2122,N_2319);
or U2919 (N_2919,N_2068,N_2321);
nand U2920 (N_2920,N_2326,N_2094);
and U2921 (N_2921,N_2183,N_2121);
or U2922 (N_2922,N_2113,N_2168);
or U2923 (N_2923,N_2157,N_2201);
and U2924 (N_2924,N_2320,N_2151);
or U2925 (N_2925,N_2451,N_2309);
nand U2926 (N_2926,N_2421,N_2452);
nand U2927 (N_2927,N_2059,N_2237);
nor U2928 (N_2928,N_2286,N_2156);
or U2929 (N_2929,N_2448,N_2312);
xor U2930 (N_2930,N_2137,N_2135);
nor U2931 (N_2931,N_2316,N_2238);
nand U2932 (N_2932,N_2310,N_2432);
nor U2933 (N_2933,N_2466,N_2021);
nand U2934 (N_2934,N_2452,N_2187);
nand U2935 (N_2935,N_2371,N_2235);
xnor U2936 (N_2936,N_2254,N_2126);
nand U2937 (N_2937,N_2075,N_2114);
xor U2938 (N_2938,N_2060,N_2005);
or U2939 (N_2939,N_2011,N_2171);
nand U2940 (N_2940,N_2404,N_2105);
nor U2941 (N_2941,N_2113,N_2446);
nor U2942 (N_2942,N_2266,N_2430);
nor U2943 (N_2943,N_2018,N_2310);
nand U2944 (N_2944,N_2325,N_2276);
or U2945 (N_2945,N_2438,N_2024);
and U2946 (N_2946,N_2151,N_2399);
and U2947 (N_2947,N_2391,N_2062);
nand U2948 (N_2948,N_2338,N_2126);
and U2949 (N_2949,N_2332,N_2493);
or U2950 (N_2950,N_2015,N_2381);
or U2951 (N_2951,N_2412,N_2158);
and U2952 (N_2952,N_2200,N_2320);
nand U2953 (N_2953,N_2224,N_2129);
and U2954 (N_2954,N_2068,N_2165);
and U2955 (N_2955,N_2414,N_2139);
nor U2956 (N_2956,N_2076,N_2424);
nand U2957 (N_2957,N_2079,N_2258);
nor U2958 (N_2958,N_2439,N_2412);
nor U2959 (N_2959,N_2166,N_2229);
nand U2960 (N_2960,N_2391,N_2456);
or U2961 (N_2961,N_2190,N_2370);
or U2962 (N_2962,N_2019,N_2053);
nand U2963 (N_2963,N_2099,N_2231);
nand U2964 (N_2964,N_2018,N_2331);
nor U2965 (N_2965,N_2378,N_2101);
or U2966 (N_2966,N_2105,N_2009);
and U2967 (N_2967,N_2074,N_2390);
or U2968 (N_2968,N_2280,N_2424);
xnor U2969 (N_2969,N_2203,N_2445);
and U2970 (N_2970,N_2400,N_2471);
nor U2971 (N_2971,N_2231,N_2026);
and U2972 (N_2972,N_2447,N_2244);
nand U2973 (N_2973,N_2310,N_2162);
nand U2974 (N_2974,N_2270,N_2070);
nand U2975 (N_2975,N_2432,N_2087);
nand U2976 (N_2976,N_2179,N_2030);
or U2977 (N_2977,N_2148,N_2011);
or U2978 (N_2978,N_2140,N_2395);
or U2979 (N_2979,N_2268,N_2368);
and U2980 (N_2980,N_2037,N_2156);
nand U2981 (N_2981,N_2498,N_2338);
nand U2982 (N_2982,N_2109,N_2220);
or U2983 (N_2983,N_2246,N_2018);
or U2984 (N_2984,N_2452,N_2474);
nor U2985 (N_2985,N_2170,N_2263);
nand U2986 (N_2986,N_2045,N_2460);
nand U2987 (N_2987,N_2341,N_2181);
and U2988 (N_2988,N_2093,N_2136);
nor U2989 (N_2989,N_2329,N_2457);
nor U2990 (N_2990,N_2154,N_2204);
and U2991 (N_2991,N_2419,N_2277);
xor U2992 (N_2992,N_2411,N_2337);
or U2993 (N_2993,N_2317,N_2407);
nor U2994 (N_2994,N_2458,N_2123);
or U2995 (N_2995,N_2278,N_2106);
or U2996 (N_2996,N_2013,N_2301);
nand U2997 (N_2997,N_2020,N_2378);
and U2998 (N_2998,N_2428,N_2087);
and U2999 (N_2999,N_2464,N_2355);
nor U3000 (N_3000,N_2523,N_2905);
nor U3001 (N_3001,N_2592,N_2960);
and U3002 (N_3002,N_2662,N_2886);
nand U3003 (N_3003,N_2907,N_2817);
nor U3004 (N_3004,N_2795,N_2947);
or U3005 (N_3005,N_2597,N_2675);
xnor U3006 (N_3006,N_2677,N_2882);
or U3007 (N_3007,N_2671,N_2839);
or U3008 (N_3008,N_2625,N_2536);
and U3009 (N_3009,N_2813,N_2652);
nand U3010 (N_3010,N_2678,N_2530);
nand U3011 (N_3011,N_2539,N_2922);
nand U3012 (N_3012,N_2520,N_2849);
nand U3013 (N_3013,N_2862,N_2572);
nand U3014 (N_3014,N_2582,N_2763);
or U3015 (N_3015,N_2807,N_2814);
nand U3016 (N_3016,N_2858,N_2878);
xnor U3017 (N_3017,N_2835,N_2921);
or U3018 (N_3018,N_2955,N_2904);
and U3019 (N_3019,N_2719,N_2594);
and U3020 (N_3020,N_2729,N_2571);
or U3021 (N_3021,N_2999,N_2647);
and U3022 (N_3022,N_2645,N_2506);
and U3023 (N_3023,N_2786,N_2900);
xor U3024 (N_3024,N_2838,N_2956);
or U3025 (N_3025,N_2965,N_2989);
xor U3026 (N_3026,N_2629,N_2889);
nand U3027 (N_3027,N_2575,N_2885);
xor U3028 (N_3028,N_2753,N_2828);
or U3029 (N_3029,N_2584,N_2747);
or U3030 (N_3030,N_2617,N_2770);
or U3031 (N_3031,N_2668,N_2957);
or U3032 (N_3032,N_2925,N_2613);
and U3033 (N_3033,N_2735,N_2961);
nor U3034 (N_3034,N_2994,N_2754);
and U3035 (N_3035,N_2550,N_2687);
or U3036 (N_3036,N_2816,N_2618);
and U3037 (N_3037,N_2896,N_2718);
nand U3038 (N_3038,N_2983,N_2864);
or U3039 (N_3039,N_2716,N_2610);
nor U3040 (N_3040,N_2940,N_2720);
xnor U3041 (N_3041,N_2758,N_2679);
nand U3042 (N_3042,N_2667,N_2837);
nor U3043 (N_3043,N_2593,N_2578);
and U3044 (N_3044,N_2590,N_2832);
or U3045 (N_3045,N_2627,N_2552);
or U3046 (N_3046,N_2636,N_2953);
or U3047 (N_3047,N_2829,N_2644);
or U3048 (N_3048,N_2676,N_2836);
nor U3049 (N_3049,N_2963,N_2910);
and U3050 (N_3050,N_2544,N_2628);
nor U3051 (N_3051,N_2902,N_2608);
nand U3052 (N_3052,N_2877,N_2982);
nand U3053 (N_3053,N_2693,N_2621);
nor U3054 (N_3054,N_2749,N_2833);
nor U3055 (N_3055,N_2852,N_2634);
nor U3056 (N_3056,N_2772,N_2917);
nand U3057 (N_3057,N_2505,N_2768);
nor U3058 (N_3058,N_2639,N_2726);
or U3059 (N_3059,N_2741,N_2551);
xnor U3060 (N_3060,N_2850,N_2527);
or U3061 (N_3061,N_2528,N_2525);
and U3062 (N_3062,N_2669,N_2611);
or U3063 (N_3063,N_2855,N_2640);
or U3064 (N_3064,N_2606,N_2650);
nand U3065 (N_3065,N_2579,N_2695);
nor U3066 (N_3066,N_2710,N_2898);
nand U3067 (N_3067,N_2932,N_2743);
nand U3068 (N_3068,N_2522,N_2901);
and U3069 (N_3069,N_2985,N_2823);
and U3070 (N_3070,N_2774,N_2993);
nand U3071 (N_3071,N_2563,N_2549);
or U3072 (N_3072,N_2865,N_2663);
nor U3073 (N_3073,N_2524,N_2631);
nand U3074 (N_3074,N_2673,N_2509);
and U3075 (N_3075,N_2703,N_2895);
nor U3076 (N_3076,N_2507,N_2767);
nand U3077 (N_3077,N_2612,N_2760);
nand U3078 (N_3078,N_2857,N_2622);
and U3079 (N_3079,N_2503,N_2851);
or U3080 (N_3080,N_2757,N_2958);
or U3081 (N_3081,N_2843,N_2806);
nor U3082 (N_3082,N_2946,N_2972);
nor U3083 (N_3083,N_2570,N_2574);
or U3084 (N_3084,N_2567,N_2756);
nand U3085 (N_3085,N_2598,N_2967);
and U3086 (N_3086,N_2822,N_2819);
nand U3087 (N_3087,N_2699,N_2740);
nand U3088 (N_3088,N_2542,N_2834);
and U3089 (N_3089,N_2804,N_2853);
or U3090 (N_3090,N_2547,N_2632);
nand U3091 (N_3091,N_2992,N_2808);
nor U3092 (N_3092,N_2721,N_2788);
or U3093 (N_3093,N_2709,N_2903);
and U3094 (N_3094,N_2688,N_2543);
nand U3095 (N_3095,N_2692,N_2927);
nor U3096 (N_3096,N_2746,N_2642);
xor U3097 (N_3097,N_2830,N_2979);
xnor U3098 (N_3098,N_2581,N_2971);
xor U3099 (N_3099,N_2970,N_2529);
xnor U3100 (N_3100,N_2751,N_2984);
xnor U3101 (N_3101,N_2775,N_2959);
or U3102 (N_3102,N_2931,N_2986);
nand U3103 (N_3103,N_2872,N_2769);
and U3104 (N_3104,N_2939,N_2897);
or U3105 (N_3105,N_2516,N_2653);
nand U3106 (N_3106,N_2587,N_2821);
nand U3107 (N_3107,N_2912,N_2704);
nor U3108 (N_3108,N_2748,N_2624);
nor U3109 (N_3109,N_2727,N_2514);
nand U3110 (N_3110,N_2890,N_2586);
nor U3111 (N_3111,N_2712,N_2920);
or U3112 (N_3112,N_2752,N_2661);
and U3113 (N_3113,N_2664,N_2777);
nand U3114 (N_3114,N_2540,N_2557);
nand U3115 (N_3115,N_2502,N_2654);
and U3116 (N_3116,N_2856,N_2919);
nor U3117 (N_3117,N_2738,N_2771);
and U3118 (N_3118,N_2537,N_2739);
nor U3119 (N_3119,N_2725,N_2684);
nor U3120 (N_3120,N_2964,N_2531);
or U3121 (N_3121,N_2519,N_2616);
nor U3122 (N_3122,N_2842,N_2831);
or U3123 (N_3123,N_2871,N_2981);
nand U3124 (N_3124,N_2556,N_2665);
nand U3125 (N_3125,N_2844,N_2873);
or U3126 (N_3126,N_2615,N_2708);
xor U3127 (N_3127,N_2690,N_2827);
nor U3128 (N_3128,N_2790,N_2724);
nor U3129 (N_3129,N_2635,N_2601);
and U3130 (N_3130,N_2685,N_2792);
and U3131 (N_3131,N_2996,N_2702);
or U3132 (N_3132,N_2680,N_2591);
or U3133 (N_3133,N_2561,N_2869);
or U3134 (N_3134,N_2534,N_2765);
xor U3135 (N_3135,N_2515,N_2697);
or U3136 (N_3136,N_2911,N_2784);
or U3137 (N_3137,N_2501,N_2553);
nor U3138 (N_3138,N_2780,N_2604);
nor U3139 (N_3139,N_2538,N_2915);
and U3140 (N_3140,N_2730,N_2863);
nand U3141 (N_3141,N_2934,N_2988);
nor U3142 (N_3142,N_2762,N_2585);
or U3143 (N_3143,N_2782,N_2643);
nand U3144 (N_3144,N_2785,N_2715);
nor U3145 (N_3145,N_2923,N_2626);
and U3146 (N_3146,N_2694,N_2545);
xor U3147 (N_3147,N_2793,N_2513);
or U3148 (N_3148,N_2870,N_2859);
xor U3149 (N_3149,N_2909,N_2825);
nor U3150 (N_3150,N_2605,N_2914);
or U3151 (N_3151,N_2766,N_2945);
or U3152 (N_3152,N_2944,N_2576);
nor U3153 (N_3153,N_2646,N_2681);
xnor U3154 (N_3154,N_2759,N_2995);
nand U3155 (N_3155,N_2805,N_2672);
or U3156 (N_3156,N_2781,N_2974);
and U3157 (N_3157,N_2734,N_2787);
and U3158 (N_3158,N_2799,N_2966);
nor U3159 (N_3159,N_2809,N_2638);
and U3160 (N_3160,N_2623,N_2991);
or U3161 (N_3161,N_2660,N_2564);
and U3162 (N_3162,N_2554,N_2783);
xor U3163 (N_3163,N_2926,N_2614);
and U3164 (N_3164,N_2811,N_2630);
nand U3165 (N_3165,N_2761,N_2742);
or U3166 (N_3166,N_2906,N_2800);
nand U3167 (N_3167,N_2848,N_2773);
or U3168 (N_3168,N_2731,N_2937);
or U3169 (N_3169,N_2568,N_2670);
nand U3170 (N_3170,N_2607,N_2930);
nand U3171 (N_3171,N_2541,N_2728);
or U3172 (N_3172,N_2950,N_2997);
xnor U3173 (N_3173,N_2875,N_2548);
xnor U3174 (N_3174,N_2512,N_2975);
nand U3175 (N_3175,N_2916,N_2560);
xnor U3176 (N_3176,N_2933,N_2508);
nand U3177 (N_3177,N_2948,N_2841);
nor U3178 (N_3178,N_2603,N_2893);
or U3179 (N_3179,N_2820,N_2689);
nand U3180 (N_3180,N_2533,N_2696);
or U3181 (N_3181,N_2854,N_2682);
and U3182 (N_3182,N_2517,N_2936);
xnor U3183 (N_3183,N_2691,N_2880);
and U3184 (N_3184,N_2973,N_2954);
xor U3185 (N_3185,N_2952,N_2504);
xor U3186 (N_3186,N_2745,N_2891);
nand U3187 (N_3187,N_2737,N_2573);
or U3188 (N_3188,N_2938,N_2619);
xor U3189 (N_3189,N_2659,N_2666);
and U3190 (N_3190,N_2649,N_2510);
xor U3191 (N_3191,N_2969,N_2845);
xor U3192 (N_3192,N_2881,N_2698);
nor U3193 (N_3193,N_2980,N_2764);
xnor U3194 (N_3194,N_2899,N_2779);
and U3195 (N_3195,N_2674,N_2532);
and U3196 (N_3196,N_2755,N_2818);
or U3197 (N_3197,N_2546,N_2589);
or U3198 (N_3198,N_2797,N_2648);
nand U3199 (N_3199,N_2651,N_2998);
xor U3200 (N_3200,N_2867,N_2658);
or U3201 (N_3201,N_2583,N_2892);
nand U3202 (N_3202,N_2723,N_2714);
and U3203 (N_3203,N_2620,N_2951);
nor U3204 (N_3204,N_2794,N_2978);
nor U3205 (N_3205,N_2713,N_2949);
or U3206 (N_3206,N_2599,N_2924);
and U3207 (N_3207,N_2987,N_2657);
nand U3208 (N_3208,N_2733,N_2596);
and U3209 (N_3209,N_2707,N_2796);
or U3210 (N_3210,N_2778,N_2812);
xnor U3211 (N_3211,N_2888,N_2883);
nand U3212 (N_3212,N_2580,N_2866);
and U3213 (N_3213,N_2801,N_2879);
and U3214 (N_3214,N_2511,N_2633);
or U3215 (N_3215,N_2750,N_2602);
nor U3216 (N_3216,N_2776,N_2609);
and U3217 (N_3217,N_2562,N_2683);
xnor U3218 (N_3218,N_2577,N_2706);
nor U3219 (N_3219,N_2810,N_2976);
nor U3220 (N_3220,N_2962,N_2518);
or U3221 (N_3221,N_2826,N_2791);
nand U3222 (N_3222,N_2705,N_2874);
or U3223 (N_3223,N_2555,N_2846);
nand U3224 (N_3224,N_2847,N_2935);
or U3225 (N_3225,N_2736,N_2928);
nor U3226 (N_3226,N_2526,N_2588);
nor U3227 (N_3227,N_2802,N_2701);
or U3228 (N_3228,N_2655,N_2894);
and U3229 (N_3229,N_2565,N_2913);
nand U3230 (N_3230,N_2968,N_2535);
or U3231 (N_3231,N_2521,N_2500);
nor U3232 (N_3232,N_2884,N_2824);
nor U3233 (N_3233,N_2840,N_2943);
or U3234 (N_3234,N_2798,N_2656);
nor U3235 (N_3235,N_2711,N_2637);
nor U3236 (N_3236,N_2941,N_2722);
or U3237 (N_3237,N_2566,N_2595);
and U3238 (N_3238,N_2929,N_2700);
nand U3239 (N_3239,N_2815,N_2559);
nor U3240 (N_3240,N_2732,N_2686);
and U3241 (N_3241,N_2918,N_2990);
nor U3242 (N_3242,N_2717,N_2744);
or U3243 (N_3243,N_2908,N_2641);
or U3244 (N_3244,N_2942,N_2558);
and U3245 (N_3245,N_2803,N_2977);
nand U3246 (N_3246,N_2860,N_2868);
or U3247 (N_3247,N_2569,N_2789);
or U3248 (N_3248,N_2887,N_2861);
or U3249 (N_3249,N_2600,N_2876);
or U3250 (N_3250,N_2805,N_2653);
nor U3251 (N_3251,N_2615,N_2922);
nor U3252 (N_3252,N_2857,N_2756);
and U3253 (N_3253,N_2791,N_2652);
and U3254 (N_3254,N_2587,N_2516);
or U3255 (N_3255,N_2936,N_2546);
and U3256 (N_3256,N_2574,N_2760);
or U3257 (N_3257,N_2511,N_2794);
or U3258 (N_3258,N_2645,N_2723);
xnor U3259 (N_3259,N_2685,N_2595);
nand U3260 (N_3260,N_2817,N_2744);
nand U3261 (N_3261,N_2632,N_2605);
or U3262 (N_3262,N_2961,N_2960);
xor U3263 (N_3263,N_2969,N_2576);
nand U3264 (N_3264,N_2846,N_2517);
or U3265 (N_3265,N_2677,N_2970);
and U3266 (N_3266,N_2525,N_2897);
and U3267 (N_3267,N_2958,N_2850);
nor U3268 (N_3268,N_2556,N_2740);
and U3269 (N_3269,N_2902,N_2803);
xnor U3270 (N_3270,N_2809,N_2938);
and U3271 (N_3271,N_2509,N_2662);
or U3272 (N_3272,N_2949,N_2645);
or U3273 (N_3273,N_2747,N_2934);
and U3274 (N_3274,N_2543,N_2758);
and U3275 (N_3275,N_2761,N_2534);
or U3276 (N_3276,N_2776,N_2687);
nor U3277 (N_3277,N_2697,N_2666);
nand U3278 (N_3278,N_2958,N_2881);
and U3279 (N_3279,N_2777,N_2670);
and U3280 (N_3280,N_2901,N_2926);
nand U3281 (N_3281,N_2692,N_2909);
and U3282 (N_3282,N_2809,N_2836);
and U3283 (N_3283,N_2850,N_2680);
or U3284 (N_3284,N_2532,N_2792);
nor U3285 (N_3285,N_2817,N_2952);
nor U3286 (N_3286,N_2699,N_2771);
or U3287 (N_3287,N_2865,N_2800);
and U3288 (N_3288,N_2763,N_2773);
nor U3289 (N_3289,N_2992,N_2723);
nand U3290 (N_3290,N_2783,N_2856);
or U3291 (N_3291,N_2807,N_2758);
nor U3292 (N_3292,N_2974,N_2561);
nand U3293 (N_3293,N_2846,N_2800);
nor U3294 (N_3294,N_2959,N_2835);
nor U3295 (N_3295,N_2548,N_2687);
and U3296 (N_3296,N_2680,N_2523);
or U3297 (N_3297,N_2570,N_2900);
or U3298 (N_3298,N_2943,N_2683);
xnor U3299 (N_3299,N_2613,N_2611);
nand U3300 (N_3300,N_2828,N_2953);
nor U3301 (N_3301,N_2635,N_2602);
nor U3302 (N_3302,N_2852,N_2684);
nand U3303 (N_3303,N_2902,N_2742);
nor U3304 (N_3304,N_2815,N_2817);
or U3305 (N_3305,N_2511,N_2914);
or U3306 (N_3306,N_2668,N_2716);
or U3307 (N_3307,N_2887,N_2671);
nand U3308 (N_3308,N_2617,N_2975);
or U3309 (N_3309,N_2868,N_2841);
nand U3310 (N_3310,N_2937,N_2778);
nor U3311 (N_3311,N_2586,N_2716);
and U3312 (N_3312,N_2523,N_2593);
nor U3313 (N_3313,N_2522,N_2890);
and U3314 (N_3314,N_2741,N_2995);
nand U3315 (N_3315,N_2920,N_2670);
nand U3316 (N_3316,N_2971,N_2606);
or U3317 (N_3317,N_2817,N_2888);
nor U3318 (N_3318,N_2599,N_2635);
and U3319 (N_3319,N_2985,N_2791);
nand U3320 (N_3320,N_2576,N_2649);
nand U3321 (N_3321,N_2507,N_2624);
nor U3322 (N_3322,N_2792,N_2660);
or U3323 (N_3323,N_2732,N_2608);
and U3324 (N_3324,N_2523,N_2690);
and U3325 (N_3325,N_2607,N_2674);
nand U3326 (N_3326,N_2720,N_2982);
nand U3327 (N_3327,N_2719,N_2532);
and U3328 (N_3328,N_2920,N_2864);
and U3329 (N_3329,N_2688,N_2840);
nor U3330 (N_3330,N_2791,N_2743);
nor U3331 (N_3331,N_2877,N_2902);
nand U3332 (N_3332,N_2556,N_2587);
nor U3333 (N_3333,N_2644,N_2852);
nor U3334 (N_3334,N_2765,N_2860);
or U3335 (N_3335,N_2946,N_2923);
nand U3336 (N_3336,N_2585,N_2706);
or U3337 (N_3337,N_2897,N_2777);
nand U3338 (N_3338,N_2801,N_2826);
nor U3339 (N_3339,N_2897,N_2661);
nand U3340 (N_3340,N_2893,N_2615);
nand U3341 (N_3341,N_2987,N_2563);
or U3342 (N_3342,N_2704,N_2646);
nor U3343 (N_3343,N_2674,N_2876);
and U3344 (N_3344,N_2956,N_2793);
xor U3345 (N_3345,N_2790,N_2711);
nand U3346 (N_3346,N_2968,N_2545);
xor U3347 (N_3347,N_2715,N_2675);
or U3348 (N_3348,N_2595,N_2738);
and U3349 (N_3349,N_2639,N_2875);
nand U3350 (N_3350,N_2523,N_2654);
nand U3351 (N_3351,N_2776,N_2642);
xnor U3352 (N_3352,N_2507,N_2872);
or U3353 (N_3353,N_2697,N_2651);
or U3354 (N_3354,N_2827,N_2970);
and U3355 (N_3355,N_2773,N_2679);
nor U3356 (N_3356,N_2792,N_2577);
nand U3357 (N_3357,N_2857,N_2959);
and U3358 (N_3358,N_2711,N_2550);
or U3359 (N_3359,N_2975,N_2884);
and U3360 (N_3360,N_2825,N_2706);
nand U3361 (N_3361,N_2598,N_2830);
and U3362 (N_3362,N_2574,N_2708);
nor U3363 (N_3363,N_2514,N_2828);
or U3364 (N_3364,N_2705,N_2729);
and U3365 (N_3365,N_2880,N_2874);
and U3366 (N_3366,N_2810,N_2515);
nand U3367 (N_3367,N_2727,N_2754);
nand U3368 (N_3368,N_2864,N_2666);
xor U3369 (N_3369,N_2720,N_2521);
nor U3370 (N_3370,N_2875,N_2536);
or U3371 (N_3371,N_2554,N_2503);
and U3372 (N_3372,N_2835,N_2663);
nor U3373 (N_3373,N_2905,N_2759);
nand U3374 (N_3374,N_2924,N_2827);
nand U3375 (N_3375,N_2691,N_2610);
xnor U3376 (N_3376,N_2694,N_2916);
nor U3377 (N_3377,N_2913,N_2523);
or U3378 (N_3378,N_2889,N_2512);
or U3379 (N_3379,N_2508,N_2849);
or U3380 (N_3380,N_2675,N_2535);
or U3381 (N_3381,N_2723,N_2904);
nor U3382 (N_3382,N_2858,N_2920);
xor U3383 (N_3383,N_2665,N_2876);
or U3384 (N_3384,N_2690,N_2881);
nand U3385 (N_3385,N_2698,N_2985);
nor U3386 (N_3386,N_2741,N_2742);
or U3387 (N_3387,N_2964,N_2991);
nor U3388 (N_3388,N_2502,N_2724);
nand U3389 (N_3389,N_2632,N_2623);
nand U3390 (N_3390,N_2504,N_2788);
nand U3391 (N_3391,N_2857,N_2618);
nor U3392 (N_3392,N_2980,N_2747);
nand U3393 (N_3393,N_2983,N_2917);
nand U3394 (N_3394,N_2628,N_2587);
nand U3395 (N_3395,N_2880,N_2773);
nor U3396 (N_3396,N_2708,N_2640);
nor U3397 (N_3397,N_2709,N_2994);
and U3398 (N_3398,N_2525,N_2601);
or U3399 (N_3399,N_2619,N_2658);
and U3400 (N_3400,N_2818,N_2756);
nand U3401 (N_3401,N_2535,N_2602);
and U3402 (N_3402,N_2767,N_2885);
nand U3403 (N_3403,N_2600,N_2625);
and U3404 (N_3404,N_2915,N_2736);
nand U3405 (N_3405,N_2873,N_2960);
or U3406 (N_3406,N_2525,N_2780);
and U3407 (N_3407,N_2929,N_2898);
nand U3408 (N_3408,N_2856,N_2934);
nor U3409 (N_3409,N_2505,N_2899);
and U3410 (N_3410,N_2933,N_2960);
xnor U3411 (N_3411,N_2672,N_2871);
xor U3412 (N_3412,N_2696,N_2808);
nand U3413 (N_3413,N_2993,N_2972);
nand U3414 (N_3414,N_2703,N_2649);
and U3415 (N_3415,N_2535,N_2670);
nand U3416 (N_3416,N_2699,N_2815);
nand U3417 (N_3417,N_2988,N_2618);
xnor U3418 (N_3418,N_2811,N_2524);
nor U3419 (N_3419,N_2947,N_2596);
nor U3420 (N_3420,N_2829,N_2688);
xor U3421 (N_3421,N_2599,N_2910);
or U3422 (N_3422,N_2612,N_2910);
nand U3423 (N_3423,N_2906,N_2803);
nor U3424 (N_3424,N_2675,N_2935);
xor U3425 (N_3425,N_2505,N_2827);
nor U3426 (N_3426,N_2715,N_2725);
nor U3427 (N_3427,N_2760,N_2672);
or U3428 (N_3428,N_2634,N_2811);
and U3429 (N_3429,N_2686,N_2708);
nor U3430 (N_3430,N_2815,N_2516);
xor U3431 (N_3431,N_2987,N_2736);
or U3432 (N_3432,N_2837,N_2947);
or U3433 (N_3433,N_2695,N_2979);
or U3434 (N_3434,N_2771,N_2912);
or U3435 (N_3435,N_2955,N_2737);
nor U3436 (N_3436,N_2700,N_2713);
and U3437 (N_3437,N_2784,N_2621);
xnor U3438 (N_3438,N_2602,N_2512);
and U3439 (N_3439,N_2663,N_2883);
and U3440 (N_3440,N_2615,N_2612);
xor U3441 (N_3441,N_2650,N_2946);
or U3442 (N_3442,N_2963,N_2760);
or U3443 (N_3443,N_2847,N_2623);
or U3444 (N_3444,N_2578,N_2540);
or U3445 (N_3445,N_2685,N_2999);
nor U3446 (N_3446,N_2638,N_2935);
nor U3447 (N_3447,N_2629,N_2706);
and U3448 (N_3448,N_2805,N_2940);
or U3449 (N_3449,N_2775,N_2721);
nor U3450 (N_3450,N_2970,N_2501);
nor U3451 (N_3451,N_2722,N_2988);
and U3452 (N_3452,N_2762,N_2722);
and U3453 (N_3453,N_2959,N_2771);
nand U3454 (N_3454,N_2601,N_2674);
nor U3455 (N_3455,N_2804,N_2581);
or U3456 (N_3456,N_2874,N_2872);
or U3457 (N_3457,N_2574,N_2723);
or U3458 (N_3458,N_2542,N_2545);
nand U3459 (N_3459,N_2730,N_2736);
and U3460 (N_3460,N_2553,N_2520);
and U3461 (N_3461,N_2867,N_2618);
and U3462 (N_3462,N_2637,N_2529);
nor U3463 (N_3463,N_2626,N_2895);
and U3464 (N_3464,N_2811,N_2652);
nor U3465 (N_3465,N_2819,N_2986);
or U3466 (N_3466,N_2756,N_2568);
or U3467 (N_3467,N_2672,N_2550);
nand U3468 (N_3468,N_2836,N_2581);
nand U3469 (N_3469,N_2584,N_2643);
nand U3470 (N_3470,N_2540,N_2895);
nand U3471 (N_3471,N_2571,N_2634);
nand U3472 (N_3472,N_2830,N_2681);
nand U3473 (N_3473,N_2984,N_2981);
or U3474 (N_3474,N_2985,N_2818);
nand U3475 (N_3475,N_2816,N_2924);
nor U3476 (N_3476,N_2554,N_2706);
or U3477 (N_3477,N_2909,N_2817);
nand U3478 (N_3478,N_2967,N_2721);
nor U3479 (N_3479,N_2882,N_2650);
or U3480 (N_3480,N_2562,N_2547);
or U3481 (N_3481,N_2699,N_2982);
nand U3482 (N_3482,N_2991,N_2817);
and U3483 (N_3483,N_2864,N_2978);
or U3484 (N_3484,N_2534,N_2807);
xnor U3485 (N_3485,N_2712,N_2650);
nor U3486 (N_3486,N_2950,N_2961);
or U3487 (N_3487,N_2818,N_2905);
and U3488 (N_3488,N_2645,N_2733);
or U3489 (N_3489,N_2685,N_2956);
or U3490 (N_3490,N_2692,N_2929);
nand U3491 (N_3491,N_2753,N_2961);
and U3492 (N_3492,N_2612,N_2603);
nand U3493 (N_3493,N_2935,N_2604);
nor U3494 (N_3494,N_2871,N_2702);
xor U3495 (N_3495,N_2868,N_2664);
nor U3496 (N_3496,N_2593,N_2612);
nand U3497 (N_3497,N_2560,N_2780);
and U3498 (N_3498,N_2858,N_2727);
nand U3499 (N_3499,N_2679,N_2970);
and U3500 (N_3500,N_3179,N_3399);
and U3501 (N_3501,N_3139,N_3053);
nor U3502 (N_3502,N_3287,N_3056);
or U3503 (N_3503,N_3403,N_3064);
and U3504 (N_3504,N_3119,N_3129);
xnor U3505 (N_3505,N_3061,N_3052);
xor U3506 (N_3506,N_3276,N_3166);
xnor U3507 (N_3507,N_3189,N_3217);
nor U3508 (N_3508,N_3341,N_3213);
nand U3509 (N_3509,N_3109,N_3377);
nor U3510 (N_3510,N_3333,N_3035);
and U3511 (N_3511,N_3021,N_3275);
and U3512 (N_3512,N_3418,N_3409);
or U3513 (N_3513,N_3019,N_3030);
xor U3514 (N_3514,N_3372,N_3088);
nand U3515 (N_3515,N_3340,N_3015);
nand U3516 (N_3516,N_3085,N_3290);
or U3517 (N_3517,N_3046,N_3337);
or U3518 (N_3518,N_3370,N_3439);
and U3519 (N_3519,N_3371,N_3176);
and U3520 (N_3520,N_3353,N_3142);
nand U3521 (N_3521,N_3181,N_3494);
and U3522 (N_3522,N_3448,N_3414);
or U3523 (N_3523,N_3241,N_3449);
nor U3524 (N_3524,N_3011,N_3442);
nand U3525 (N_3525,N_3288,N_3223);
nand U3526 (N_3526,N_3410,N_3062);
xnor U3527 (N_3527,N_3328,N_3134);
or U3528 (N_3528,N_3157,N_3146);
nand U3529 (N_3529,N_3274,N_3209);
and U3530 (N_3530,N_3206,N_3292);
nand U3531 (N_3531,N_3224,N_3164);
and U3532 (N_3532,N_3481,N_3091);
nand U3533 (N_3533,N_3248,N_3130);
or U3534 (N_3534,N_3155,N_3081);
nor U3535 (N_3535,N_3362,N_3249);
and U3536 (N_3536,N_3401,N_3231);
nand U3537 (N_3537,N_3354,N_3461);
and U3538 (N_3538,N_3092,N_3289);
nor U3539 (N_3539,N_3211,N_3296);
or U3540 (N_3540,N_3428,N_3280);
or U3541 (N_3541,N_3147,N_3295);
or U3542 (N_3542,N_3446,N_3283);
nand U3543 (N_3543,N_3273,N_3330);
nand U3544 (N_3544,N_3272,N_3349);
xnor U3545 (N_3545,N_3498,N_3205);
nand U3546 (N_3546,N_3323,N_3426);
nand U3547 (N_3547,N_3178,N_3282);
nor U3548 (N_3548,N_3200,N_3028);
nand U3549 (N_3549,N_3234,N_3201);
and U3550 (N_3550,N_3041,N_3121);
or U3551 (N_3551,N_3060,N_3188);
and U3552 (N_3552,N_3003,N_3012);
or U3553 (N_3553,N_3141,N_3090);
and U3554 (N_3554,N_3436,N_3383);
or U3555 (N_3555,N_3480,N_3154);
xnor U3556 (N_3556,N_3100,N_3363);
xnor U3557 (N_3557,N_3047,N_3450);
nor U3558 (N_3558,N_3116,N_3464);
nor U3559 (N_3559,N_3043,N_3360);
nand U3560 (N_3560,N_3271,N_3044);
nor U3561 (N_3561,N_3123,N_3084);
or U3562 (N_3562,N_3259,N_3322);
nor U3563 (N_3563,N_3350,N_3379);
nor U3564 (N_3564,N_3359,N_3455);
and U3565 (N_3565,N_3058,N_3468);
and U3566 (N_3566,N_3388,N_3482);
nor U3567 (N_3567,N_3315,N_3361);
nand U3568 (N_3568,N_3197,N_3261);
and U3569 (N_3569,N_3497,N_3059);
nand U3570 (N_3570,N_3055,N_3358);
nor U3571 (N_3571,N_3394,N_3396);
nand U3572 (N_3572,N_3438,N_3195);
or U3573 (N_3573,N_3304,N_3153);
and U3574 (N_3574,N_3489,N_3013);
and U3575 (N_3575,N_3402,N_3267);
or U3576 (N_3576,N_3242,N_3196);
nand U3577 (N_3577,N_3252,N_3472);
and U3578 (N_3578,N_3082,N_3392);
and U3579 (N_3579,N_3460,N_3148);
nor U3580 (N_3580,N_3108,N_3018);
nor U3581 (N_3581,N_3001,N_3318);
nand U3582 (N_3582,N_3485,N_3133);
nor U3583 (N_3583,N_3162,N_3111);
and U3584 (N_3584,N_3320,N_3079);
nor U3585 (N_3585,N_3313,N_3429);
or U3586 (N_3586,N_3457,N_3415);
and U3587 (N_3587,N_3413,N_3270);
nor U3588 (N_3588,N_3039,N_3484);
or U3589 (N_3589,N_3168,N_3086);
or U3590 (N_3590,N_3391,N_3306);
and U3591 (N_3591,N_3218,N_3294);
and U3592 (N_3592,N_3150,N_3346);
nor U3593 (N_3593,N_3260,N_3317);
and U3594 (N_3594,N_3034,N_3463);
nor U3595 (N_3595,N_3203,N_3279);
and U3596 (N_3596,N_3104,N_3066);
xor U3597 (N_3597,N_3040,N_3171);
or U3598 (N_3598,N_3348,N_3291);
and U3599 (N_3599,N_3338,N_3376);
nor U3600 (N_3600,N_3397,N_3452);
nor U3601 (N_3601,N_3487,N_3431);
nand U3602 (N_3602,N_3386,N_3471);
nand U3603 (N_3603,N_3327,N_3057);
or U3604 (N_3604,N_3037,N_3262);
nand U3605 (N_3605,N_3207,N_3006);
or U3606 (N_3606,N_3319,N_3278);
nor U3607 (N_3607,N_3281,N_3118);
nand U3608 (N_3608,N_3246,N_3299);
nand U3609 (N_3609,N_3405,N_3192);
xor U3610 (N_3610,N_3033,N_3398);
nand U3611 (N_3611,N_3238,N_3344);
nand U3612 (N_3612,N_3068,N_3311);
and U3613 (N_3613,N_3099,N_3264);
nor U3614 (N_3614,N_3182,N_3470);
and U3615 (N_3615,N_3172,N_3406);
xnor U3616 (N_3616,N_3444,N_3131);
nand U3617 (N_3617,N_3112,N_3000);
nand U3618 (N_3618,N_3007,N_3366);
nand U3619 (N_3619,N_3483,N_3173);
or U3620 (N_3620,N_3220,N_3054);
and U3621 (N_3621,N_3441,N_3072);
and U3622 (N_3622,N_3447,N_3478);
or U3623 (N_3623,N_3045,N_3076);
and U3624 (N_3624,N_3032,N_3493);
or U3625 (N_3625,N_3343,N_3375);
or U3626 (N_3626,N_3445,N_3297);
and U3627 (N_3627,N_3286,N_3073);
and U3628 (N_3628,N_3243,N_3352);
or U3629 (N_3629,N_3214,N_3114);
nor U3630 (N_3630,N_3204,N_3074);
nand U3631 (N_3631,N_3314,N_3198);
and U3632 (N_3632,N_3301,N_3244);
nor U3633 (N_3633,N_3016,N_3475);
or U3634 (N_3634,N_3474,N_3215);
and U3635 (N_3635,N_3456,N_3145);
or U3636 (N_3636,N_3325,N_3093);
or U3637 (N_3637,N_3151,N_3126);
nor U3638 (N_3638,N_3310,N_3219);
nor U3639 (N_3639,N_3095,N_3163);
nand U3640 (N_3640,N_3459,N_3412);
nand U3641 (N_3641,N_3347,N_3302);
and U3642 (N_3642,N_3422,N_3122);
xnor U3643 (N_3643,N_3185,N_3427);
or U3644 (N_3644,N_3269,N_3312);
nor U3645 (N_3645,N_3378,N_3423);
and U3646 (N_3646,N_3120,N_3331);
and U3647 (N_3647,N_3309,N_3335);
and U3648 (N_3648,N_3368,N_3228);
nand U3649 (N_3649,N_3125,N_3149);
nand U3650 (N_3650,N_3385,N_3124);
nand U3651 (N_3651,N_3477,N_3421);
nor U3652 (N_3652,N_3435,N_3174);
or U3653 (N_3653,N_3106,N_3369);
nor U3654 (N_3654,N_3127,N_3070);
nor U3655 (N_3655,N_3193,N_3050);
or U3656 (N_3656,N_3355,N_3365);
and U3657 (N_3657,N_3080,N_3138);
and U3658 (N_3658,N_3135,N_3321);
or U3659 (N_3659,N_3400,N_3143);
xor U3660 (N_3660,N_3115,N_3434);
nor U3661 (N_3661,N_3326,N_3165);
nor U3662 (N_3662,N_3184,N_3136);
or U3663 (N_3663,N_3454,N_3430);
nor U3664 (N_3664,N_3194,N_3334);
nor U3665 (N_3665,N_3107,N_3425);
and U3666 (N_3666,N_3373,N_3389);
nor U3667 (N_3667,N_3411,N_3424);
nand U3668 (N_3668,N_3177,N_3089);
nand U3669 (N_3669,N_3466,N_3258);
xor U3670 (N_3670,N_3458,N_3048);
xnor U3671 (N_3671,N_3437,N_3380);
nor U3672 (N_3672,N_3152,N_3117);
nor U3673 (N_3673,N_3020,N_3404);
and U3674 (N_3674,N_3324,N_3256);
or U3675 (N_3675,N_3268,N_3075);
nor U3676 (N_3676,N_3049,N_3105);
or U3677 (N_3677,N_3101,N_3005);
or U3678 (N_3678,N_3462,N_3381);
xor U3679 (N_3679,N_3029,N_3277);
nor U3680 (N_3680,N_3491,N_3357);
and U3681 (N_3681,N_3025,N_3308);
and U3682 (N_3682,N_3253,N_3251);
or U3683 (N_3683,N_3221,N_3071);
nor U3684 (N_3684,N_3156,N_3467);
nor U3685 (N_3685,N_3469,N_3009);
or U3686 (N_3686,N_3298,N_3160);
nor U3687 (N_3687,N_3307,N_3395);
and U3688 (N_3688,N_3096,N_3230);
or U3689 (N_3689,N_3180,N_3239);
nor U3690 (N_3690,N_3257,N_3202);
and U3691 (N_3691,N_3284,N_3097);
xor U3692 (N_3692,N_3247,N_3113);
xnor U3693 (N_3693,N_3233,N_3453);
nand U3694 (N_3694,N_3110,N_3199);
or U3695 (N_3695,N_3237,N_3067);
nor U3696 (N_3696,N_3103,N_3367);
or U3697 (N_3697,N_3190,N_3465);
or U3698 (N_3698,N_3022,N_3476);
or U3699 (N_3699,N_3473,N_3255);
or U3700 (N_3700,N_3137,N_3026);
nand U3701 (N_3701,N_3490,N_3488);
nand U3702 (N_3702,N_3140,N_3002);
nand U3703 (N_3703,N_3492,N_3300);
nand U3704 (N_3704,N_3208,N_3063);
nor U3705 (N_3705,N_3065,N_3042);
nor U3706 (N_3706,N_3144,N_3027);
or U3707 (N_3707,N_3186,N_3051);
nor U3708 (N_3708,N_3479,N_3038);
nand U3709 (N_3709,N_3408,N_3336);
nor U3710 (N_3710,N_3451,N_3102);
or U3711 (N_3711,N_3036,N_3159);
nand U3712 (N_3712,N_3024,N_3212);
nand U3713 (N_3713,N_3305,N_3175);
nand U3714 (N_3714,N_3332,N_3345);
nor U3715 (N_3715,N_3128,N_3031);
nor U3716 (N_3716,N_3351,N_3356);
nor U3717 (N_3717,N_3170,N_3390);
and U3718 (N_3718,N_3017,N_3285);
and U3719 (N_3719,N_3083,N_3132);
and U3720 (N_3720,N_3486,N_3014);
nand U3721 (N_3721,N_3316,N_3187);
xnor U3722 (N_3722,N_3495,N_3161);
or U3723 (N_3723,N_3227,N_3417);
or U3724 (N_3724,N_3419,N_3225);
and U3725 (N_3725,N_3078,N_3167);
nand U3726 (N_3726,N_3008,N_3499);
nor U3727 (N_3727,N_3004,N_3250);
and U3728 (N_3728,N_3094,N_3382);
or U3729 (N_3729,N_3420,N_3496);
or U3730 (N_3730,N_3443,N_3210);
nand U3731 (N_3731,N_3098,N_3263);
and U3732 (N_3732,N_3087,N_3393);
or U3733 (N_3733,N_3364,N_3235);
and U3734 (N_3734,N_3384,N_3240);
nor U3735 (N_3735,N_3432,N_3232);
nor U3736 (N_3736,N_3077,N_3329);
nor U3737 (N_3737,N_3433,N_3387);
or U3738 (N_3738,N_3339,N_3342);
and U3739 (N_3739,N_3158,N_3245);
and U3740 (N_3740,N_3416,N_3216);
nor U3741 (N_3741,N_3254,N_3265);
and U3742 (N_3742,N_3010,N_3191);
and U3743 (N_3743,N_3374,N_3183);
or U3744 (N_3744,N_3229,N_3293);
nand U3745 (N_3745,N_3266,N_3407);
and U3746 (N_3746,N_3069,N_3236);
and U3747 (N_3747,N_3169,N_3222);
nor U3748 (N_3748,N_3226,N_3303);
xnor U3749 (N_3749,N_3023,N_3440);
or U3750 (N_3750,N_3272,N_3079);
or U3751 (N_3751,N_3108,N_3378);
nor U3752 (N_3752,N_3162,N_3242);
nand U3753 (N_3753,N_3493,N_3209);
nor U3754 (N_3754,N_3003,N_3275);
or U3755 (N_3755,N_3107,N_3385);
nor U3756 (N_3756,N_3036,N_3269);
or U3757 (N_3757,N_3298,N_3063);
xnor U3758 (N_3758,N_3227,N_3421);
nor U3759 (N_3759,N_3449,N_3436);
nor U3760 (N_3760,N_3052,N_3420);
nand U3761 (N_3761,N_3050,N_3161);
or U3762 (N_3762,N_3392,N_3190);
or U3763 (N_3763,N_3030,N_3318);
xor U3764 (N_3764,N_3413,N_3447);
and U3765 (N_3765,N_3261,N_3195);
and U3766 (N_3766,N_3320,N_3282);
or U3767 (N_3767,N_3044,N_3487);
nand U3768 (N_3768,N_3207,N_3308);
and U3769 (N_3769,N_3425,N_3346);
nand U3770 (N_3770,N_3286,N_3038);
xor U3771 (N_3771,N_3123,N_3268);
nor U3772 (N_3772,N_3304,N_3432);
xor U3773 (N_3773,N_3386,N_3166);
and U3774 (N_3774,N_3114,N_3258);
nand U3775 (N_3775,N_3359,N_3218);
xnor U3776 (N_3776,N_3235,N_3412);
xor U3777 (N_3777,N_3330,N_3201);
or U3778 (N_3778,N_3252,N_3024);
xor U3779 (N_3779,N_3098,N_3146);
and U3780 (N_3780,N_3051,N_3393);
nand U3781 (N_3781,N_3037,N_3233);
or U3782 (N_3782,N_3198,N_3215);
nor U3783 (N_3783,N_3371,N_3437);
and U3784 (N_3784,N_3027,N_3488);
nor U3785 (N_3785,N_3251,N_3031);
nand U3786 (N_3786,N_3224,N_3339);
or U3787 (N_3787,N_3188,N_3409);
and U3788 (N_3788,N_3011,N_3417);
and U3789 (N_3789,N_3078,N_3405);
and U3790 (N_3790,N_3095,N_3459);
nor U3791 (N_3791,N_3283,N_3049);
nand U3792 (N_3792,N_3188,N_3468);
nor U3793 (N_3793,N_3369,N_3005);
nor U3794 (N_3794,N_3052,N_3360);
or U3795 (N_3795,N_3352,N_3178);
xor U3796 (N_3796,N_3425,N_3142);
xor U3797 (N_3797,N_3083,N_3189);
or U3798 (N_3798,N_3371,N_3332);
nor U3799 (N_3799,N_3120,N_3450);
or U3800 (N_3800,N_3487,N_3190);
nor U3801 (N_3801,N_3443,N_3017);
nand U3802 (N_3802,N_3041,N_3328);
or U3803 (N_3803,N_3030,N_3406);
and U3804 (N_3804,N_3072,N_3375);
or U3805 (N_3805,N_3240,N_3024);
and U3806 (N_3806,N_3040,N_3191);
and U3807 (N_3807,N_3488,N_3152);
nand U3808 (N_3808,N_3222,N_3191);
or U3809 (N_3809,N_3360,N_3335);
nand U3810 (N_3810,N_3162,N_3389);
nor U3811 (N_3811,N_3046,N_3419);
or U3812 (N_3812,N_3049,N_3037);
nand U3813 (N_3813,N_3126,N_3045);
nor U3814 (N_3814,N_3399,N_3292);
nor U3815 (N_3815,N_3321,N_3111);
or U3816 (N_3816,N_3285,N_3107);
or U3817 (N_3817,N_3002,N_3079);
nor U3818 (N_3818,N_3154,N_3011);
nand U3819 (N_3819,N_3245,N_3167);
or U3820 (N_3820,N_3366,N_3247);
nand U3821 (N_3821,N_3174,N_3070);
and U3822 (N_3822,N_3001,N_3315);
nand U3823 (N_3823,N_3411,N_3410);
and U3824 (N_3824,N_3329,N_3241);
and U3825 (N_3825,N_3341,N_3469);
and U3826 (N_3826,N_3365,N_3135);
nand U3827 (N_3827,N_3255,N_3311);
and U3828 (N_3828,N_3035,N_3289);
nand U3829 (N_3829,N_3234,N_3281);
nor U3830 (N_3830,N_3427,N_3191);
nand U3831 (N_3831,N_3066,N_3424);
and U3832 (N_3832,N_3165,N_3093);
or U3833 (N_3833,N_3090,N_3299);
xnor U3834 (N_3834,N_3238,N_3179);
and U3835 (N_3835,N_3074,N_3265);
nor U3836 (N_3836,N_3136,N_3314);
xor U3837 (N_3837,N_3034,N_3200);
or U3838 (N_3838,N_3262,N_3380);
nor U3839 (N_3839,N_3183,N_3432);
nand U3840 (N_3840,N_3098,N_3259);
nor U3841 (N_3841,N_3222,N_3430);
or U3842 (N_3842,N_3221,N_3006);
or U3843 (N_3843,N_3038,N_3231);
and U3844 (N_3844,N_3332,N_3394);
nor U3845 (N_3845,N_3285,N_3430);
and U3846 (N_3846,N_3140,N_3364);
nand U3847 (N_3847,N_3428,N_3117);
nor U3848 (N_3848,N_3196,N_3078);
xor U3849 (N_3849,N_3199,N_3177);
and U3850 (N_3850,N_3004,N_3340);
nand U3851 (N_3851,N_3438,N_3159);
and U3852 (N_3852,N_3435,N_3339);
or U3853 (N_3853,N_3322,N_3191);
and U3854 (N_3854,N_3490,N_3122);
nor U3855 (N_3855,N_3058,N_3404);
and U3856 (N_3856,N_3223,N_3253);
xnor U3857 (N_3857,N_3252,N_3370);
nor U3858 (N_3858,N_3336,N_3492);
nand U3859 (N_3859,N_3201,N_3320);
nand U3860 (N_3860,N_3432,N_3275);
or U3861 (N_3861,N_3354,N_3272);
or U3862 (N_3862,N_3330,N_3167);
nand U3863 (N_3863,N_3201,N_3232);
and U3864 (N_3864,N_3077,N_3148);
or U3865 (N_3865,N_3305,N_3049);
or U3866 (N_3866,N_3020,N_3495);
or U3867 (N_3867,N_3039,N_3177);
nand U3868 (N_3868,N_3144,N_3420);
nor U3869 (N_3869,N_3387,N_3050);
and U3870 (N_3870,N_3108,N_3286);
and U3871 (N_3871,N_3240,N_3386);
nand U3872 (N_3872,N_3255,N_3139);
nor U3873 (N_3873,N_3294,N_3182);
nand U3874 (N_3874,N_3249,N_3172);
or U3875 (N_3875,N_3333,N_3401);
or U3876 (N_3876,N_3211,N_3183);
nand U3877 (N_3877,N_3495,N_3162);
nor U3878 (N_3878,N_3201,N_3053);
nand U3879 (N_3879,N_3284,N_3081);
nand U3880 (N_3880,N_3055,N_3111);
and U3881 (N_3881,N_3428,N_3426);
nand U3882 (N_3882,N_3237,N_3330);
xor U3883 (N_3883,N_3339,N_3387);
nor U3884 (N_3884,N_3077,N_3416);
nand U3885 (N_3885,N_3122,N_3066);
and U3886 (N_3886,N_3465,N_3434);
nand U3887 (N_3887,N_3039,N_3368);
or U3888 (N_3888,N_3239,N_3200);
xnor U3889 (N_3889,N_3443,N_3478);
nor U3890 (N_3890,N_3238,N_3470);
nand U3891 (N_3891,N_3050,N_3008);
and U3892 (N_3892,N_3416,N_3305);
and U3893 (N_3893,N_3108,N_3395);
nor U3894 (N_3894,N_3199,N_3342);
and U3895 (N_3895,N_3027,N_3272);
nand U3896 (N_3896,N_3471,N_3464);
nor U3897 (N_3897,N_3385,N_3156);
and U3898 (N_3898,N_3123,N_3467);
nand U3899 (N_3899,N_3050,N_3096);
or U3900 (N_3900,N_3048,N_3443);
nand U3901 (N_3901,N_3348,N_3082);
nor U3902 (N_3902,N_3358,N_3054);
and U3903 (N_3903,N_3165,N_3401);
and U3904 (N_3904,N_3180,N_3278);
or U3905 (N_3905,N_3005,N_3392);
nor U3906 (N_3906,N_3123,N_3313);
nand U3907 (N_3907,N_3265,N_3421);
or U3908 (N_3908,N_3034,N_3465);
and U3909 (N_3909,N_3351,N_3237);
nand U3910 (N_3910,N_3183,N_3205);
or U3911 (N_3911,N_3056,N_3041);
nand U3912 (N_3912,N_3117,N_3100);
xnor U3913 (N_3913,N_3337,N_3468);
nand U3914 (N_3914,N_3278,N_3406);
and U3915 (N_3915,N_3291,N_3113);
nor U3916 (N_3916,N_3290,N_3262);
nand U3917 (N_3917,N_3344,N_3229);
nor U3918 (N_3918,N_3424,N_3128);
or U3919 (N_3919,N_3188,N_3252);
xnor U3920 (N_3920,N_3376,N_3048);
and U3921 (N_3921,N_3432,N_3063);
or U3922 (N_3922,N_3116,N_3304);
nand U3923 (N_3923,N_3036,N_3403);
or U3924 (N_3924,N_3168,N_3313);
and U3925 (N_3925,N_3164,N_3301);
nor U3926 (N_3926,N_3035,N_3232);
nor U3927 (N_3927,N_3388,N_3082);
xor U3928 (N_3928,N_3002,N_3345);
xnor U3929 (N_3929,N_3213,N_3315);
nor U3930 (N_3930,N_3233,N_3065);
and U3931 (N_3931,N_3433,N_3425);
nand U3932 (N_3932,N_3214,N_3496);
or U3933 (N_3933,N_3294,N_3044);
nand U3934 (N_3934,N_3185,N_3296);
nand U3935 (N_3935,N_3033,N_3042);
nor U3936 (N_3936,N_3439,N_3367);
or U3937 (N_3937,N_3017,N_3068);
nor U3938 (N_3938,N_3479,N_3124);
and U3939 (N_3939,N_3072,N_3487);
nor U3940 (N_3940,N_3245,N_3156);
nand U3941 (N_3941,N_3459,N_3027);
nor U3942 (N_3942,N_3351,N_3079);
nor U3943 (N_3943,N_3400,N_3037);
xnor U3944 (N_3944,N_3278,N_3389);
or U3945 (N_3945,N_3012,N_3457);
nor U3946 (N_3946,N_3285,N_3104);
nor U3947 (N_3947,N_3351,N_3342);
nand U3948 (N_3948,N_3037,N_3143);
xnor U3949 (N_3949,N_3018,N_3107);
nor U3950 (N_3950,N_3341,N_3043);
or U3951 (N_3951,N_3208,N_3019);
or U3952 (N_3952,N_3168,N_3451);
or U3953 (N_3953,N_3233,N_3361);
nand U3954 (N_3954,N_3289,N_3078);
and U3955 (N_3955,N_3414,N_3119);
xnor U3956 (N_3956,N_3126,N_3333);
and U3957 (N_3957,N_3466,N_3139);
and U3958 (N_3958,N_3250,N_3111);
or U3959 (N_3959,N_3116,N_3367);
nand U3960 (N_3960,N_3294,N_3479);
and U3961 (N_3961,N_3138,N_3110);
and U3962 (N_3962,N_3211,N_3356);
nor U3963 (N_3963,N_3111,N_3199);
nand U3964 (N_3964,N_3432,N_3417);
or U3965 (N_3965,N_3153,N_3031);
nand U3966 (N_3966,N_3412,N_3359);
xor U3967 (N_3967,N_3264,N_3027);
nor U3968 (N_3968,N_3169,N_3403);
nand U3969 (N_3969,N_3182,N_3302);
nand U3970 (N_3970,N_3172,N_3174);
xnor U3971 (N_3971,N_3024,N_3143);
and U3972 (N_3972,N_3485,N_3355);
and U3973 (N_3973,N_3083,N_3441);
and U3974 (N_3974,N_3293,N_3410);
or U3975 (N_3975,N_3252,N_3114);
nand U3976 (N_3976,N_3313,N_3476);
nand U3977 (N_3977,N_3285,N_3307);
and U3978 (N_3978,N_3203,N_3320);
xor U3979 (N_3979,N_3276,N_3149);
and U3980 (N_3980,N_3095,N_3108);
nand U3981 (N_3981,N_3407,N_3238);
nor U3982 (N_3982,N_3357,N_3069);
or U3983 (N_3983,N_3439,N_3340);
or U3984 (N_3984,N_3436,N_3318);
xnor U3985 (N_3985,N_3396,N_3035);
and U3986 (N_3986,N_3319,N_3449);
nor U3987 (N_3987,N_3090,N_3007);
xor U3988 (N_3988,N_3186,N_3002);
and U3989 (N_3989,N_3011,N_3036);
or U3990 (N_3990,N_3314,N_3025);
xnor U3991 (N_3991,N_3027,N_3022);
nor U3992 (N_3992,N_3017,N_3356);
nor U3993 (N_3993,N_3322,N_3391);
nor U3994 (N_3994,N_3267,N_3075);
or U3995 (N_3995,N_3154,N_3046);
and U3996 (N_3996,N_3299,N_3266);
nor U3997 (N_3997,N_3223,N_3216);
and U3998 (N_3998,N_3338,N_3070);
xor U3999 (N_3999,N_3015,N_3079);
xor U4000 (N_4000,N_3890,N_3547);
nor U4001 (N_4001,N_3705,N_3803);
nand U4002 (N_4002,N_3976,N_3557);
nor U4003 (N_4003,N_3985,N_3532);
nand U4004 (N_4004,N_3942,N_3970);
and U4005 (N_4005,N_3949,N_3741);
nand U4006 (N_4006,N_3542,N_3945);
nand U4007 (N_4007,N_3851,N_3700);
nor U4008 (N_4008,N_3875,N_3990);
nand U4009 (N_4009,N_3989,N_3702);
nand U4010 (N_4010,N_3939,N_3790);
xor U4011 (N_4011,N_3974,N_3601);
or U4012 (N_4012,N_3968,N_3716);
or U4013 (N_4013,N_3962,N_3513);
or U4014 (N_4014,N_3666,N_3841);
nor U4015 (N_4015,N_3564,N_3783);
nor U4016 (N_4016,N_3750,N_3895);
nor U4017 (N_4017,N_3820,N_3606);
or U4018 (N_4018,N_3578,N_3500);
xor U4019 (N_4019,N_3586,N_3948);
or U4020 (N_4020,N_3610,N_3929);
and U4021 (N_4021,N_3631,N_3537);
nand U4022 (N_4022,N_3793,N_3785);
nand U4023 (N_4023,N_3580,N_3863);
xor U4024 (N_4024,N_3650,N_3763);
and U4025 (N_4025,N_3726,N_3842);
and U4026 (N_4026,N_3769,N_3662);
nand U4027 (N_4027,N_3731,N_3552);
nor U4028 (N_4028,N_3972,N_3617);
or U4029 (N_4029,N_3922,N_3670);
nand U4030 (N_4030,N_3638,N_3663);
and U4031 (N_4031,N_3612,N_3888);
nor U4032 (N_4032,N_3519,N_3882);
or U4033 (N_4033,N_3923,N_3761);
nor U4034 (N_4034,N_3687,N_3739);
nand U4035 (N_4035,N_3987,N_3541);
nor U4036 (N_4036,N_3901,N_3717);
nand U4037 (N_4037,N_3577,N_3548);
and U4038 (N_4038,N_3986,N_3878);
and U4039 (N_4039,N_3819,N_3900);
xor U4040 (N_4040,N_3637,N_3646);
xnor U4041 (N_4041,N_3874,N_3518);
nor U4042 (N_4042,N_3908,N_3920);
and U4043 (N_4043,N_3680,N_3805);
nand U4044 (N_4044,N_3672,N_3517);
xor U4045 (N_4045,N_3921,N_3801);
nor U4046 (N_4046,N_3991,N_3816);
xor U4047 (N_4047,N_3529,N_3559);
and U4048 (N_4048,N_3679,N_3833);
nand U4049 (N_4049,N_3728,N_3583);
and U4050 (N_4050,N_3915,N_3897);
or U4051 (N_4051,N_3735,N_3864);
nor U4052 (N_4052,N_3540,N_3850);
or U4053 (N_4053,N_3659,N_3959);
and U4054 (N_4054,N_3524,N_3521);
nor U4055 (N_4055,N_3817,N_3597);
nand U4056 (N_4056,N_3853,N_3778);
nand U4057 (N_4057,N_3812,N_3550);
and U4058 (N_4058,N_3595,N_3749);
or U4059 (N_4059,N_3747,N_3993);
nor U4060 (N_4060,N_3604,N_3714);
xor U4061 (N_4061,N_3701,N_3957);
xor U4062 (N_4062,N_3737,N_3756);
nand U4063 (N_4063,N_3967,N_3574);
nand U4064 (N_4064,N_3998,N_3880);
nor U4065 (N_4065,N_3960,N_3907);
and U4066 (N_4066,N_3562,N_3773);
nand U4067 (N_4067,N_3914,N_3899);
or U4068 (N_4068,N_3782,N_3533);
or U4069 (N_4069,N_3682,N_3822);
or U4070 (N_4070,N_3905,N_3626);
or U4071 (N_4071,N_3732,N_3909);
and U4072 (N_4072,N_3876,N_3648);
xor U4073 (N_4073,N_3730,N_3535);
or U4074 (N_4074,N_3556,N_3706);
and U4075 (N_4075,N_3719,N_3544);
or U4076 (N_4076,N_3891,N_3947);
nor U4077 (N_4077,N_3683,N_3796);
and U4078 (N_4078,N_3613,N_3867);
nand U4079 (N_4079,N_3635,N_3599);
or U4080 (N_4080,N_3570,N_3752);
and U4081 (N_4081,N_3608,N_3757);
nand U4082 (N_4082,N_3733,N_3509);
nor U4083 (N_4083,N_3994,N_3800);
xnor U4084 (N_4084,N_3953,N_3893);
and U4085 (N_4085,N_3847,N_3636);
and U4086 (N_4086,N_3910,N_3966);
xor U4087 (N_4087,N_3924,N_3591);
nand U4088 (N_4088,N_3543,N_3568);
xor U4089 (N_4089,N_3775,N_3676);
nor U4090 (N_4090,N_3919,N_3804);
nor U4091 (N_4091,N_3653,N_3622);
or U4092 (N_4092,N_3585,N_3933);
xnor U4093 (N_4093,N_3871,N_3879);
nor U4094 (N_4094,N_3872,N_3545);
or U4095 (N_4095,N_3786,N_3697);
or U4096 (N_4096,N_3669,N_3588);
nor U4097 (N_4097,N_3955,N_3632);
and U4098 (N_4098,N_3710,N_3881);
or U4099 (N_4099,N_3896,N_3673);
nand U4100 (N_4100,N_3885,N_3992);
nor U4101 (N_4101,N_3536,N_3944);
nor U4102 (N_4102,N_3858,N_3977);
nand U4103 (N_4103,N_3639,N_3675);
nand U4104 (N_4104,N_3753,N_3645);
nor U4105 (N_4105,N_3627,N_3596);
nor U4106 (N_4106,N_3810,N_3937);
or U4107 (N_4107,N_3501,N_3649);
xnor U4108 (N_4108,N_3829,N_3551);
xnor U4109 (N_4109,N_3744,N_3983);
and U4110 (N_4110,N_3865,N_3678);
nor U4111 (N_4111,N_3625,N_3522);
nand U4112 (N_4112,N_3770,N_3852);
nand U4113 (N_4113,N_3502,N_3515);
or U4114 (N_4114,N_3788,N_3836);
nand U4115 (N_4115,N_3767,N_3765);
xor U4116 (N_4116,N_3898,N_3640);
nor U4117 (N_4117,N_3758,N_3877);
nor U4118 (N_4118,N_3712,N_3709);
nand U4119 (N_4119,N_3815,N_3724);
nand U4120 (N_4120,N_3651,N_3742);
or U4121 (N_4121,N_3759,N_3727);
and U4122 (N_4122,N_3904,N_3734);
nand U4123 (N_4123,N_3791,N_3722);
xnor U4124 (N_4124,N_3504,N_3546);
and U4125 (N_4125,N_3575,N_3861);
xnor U4126 (N_4126,N_3748,N_3889);
or U4127 (N_4127,N_3554,N_3707);
or U4128 (N_4128,N_3657,N_3615);
and U4129 (N_4129,N_3718,N_3859);
nand U4130 (N_4130,N_3661,N_3843);
xor U4131 (N_4131,N_3832,N_3979);
nor U4132 (N_4132,N_3658,N_3711);
or U4133 (N_4133,N_3723,N_3654);
nand U4134 (N_4134,N_3708,N_3931);
and U4135 (N_4135,N_3609,N_3930);
xor U4136 (N_4136,N_3799,N_3665);
nor U4137 (N_4137,N_3934,N_3981);
nand U4138 (N_4138,N_3507,N_3693);
nor U4139 (N_4139,N_3902,N_3961);
xnor U4140 (N_4140,N_3927,N_3621);
nand U4141 (N_4141,N_3980,N_3571);
nor U4142 (N_4142,N_3579,N_3698);
nand U4143 (N_4143,N_3779,N_3984);
xnor U4144 (N_4144,N_3720,N_3618);
nor U4145 (N_4145,N_3883,N_3956);
nor U4146 (N_4146,N_3794,N_3660);
and U4147 (N_4147,N_3592,N_3894);
xor U4148 (N_4148,N_3642,N_3837);
and U4149 (N_4149,N_3818,N_3685);
and U4150 (N_4150,N_3721,N_3764);
and U4151 (N_4151,N_3561,N_3906);
or U4152 (N_4152,N_3978,N_3534);
xnor U4153 (N_4153,N_3602,N_3982);
nor U4154 (N_4154,N_3807,N_3797);
and U4155 (N_4155,N_3652,N_3811);
nor U4156 (N_4156,N_3954,N_3538);
or U4157 (N_4157,N_3835,N_3674);
nor U4158 (N_4158,N_3743,N_3892);
nor U4159 (N_4159,N_3768,N_3780);
xor U4160 (N_4160,N_3520,N_3848);
xor U4161 (N_4161,N_3582,N_3809);
nand U4162 (N_4162,N_3826,N_3751);
xor U4163 (N_4163,N_3526,N_3576);
or U4164 (N_4164,N_3845,N_3691);
nand U4165 (N_4165,N_3656,N_3814);
or U4166 (N_4166,N_3624,N_3584);
or U4167 (N_4167,N_3681,N_3950);
and U4168 (N_4168,N_3629,N_3754);
nor U4169 (N_4169,N_3713,N_3928);
nand U4170 (N_4170,N_3846,N_3975);
nor U4171 (N_4171,N_3971,N_3995);
nor U4172 (N_4172,N_3725,N_3834);
and U4173 (N_4173,N_3516,N_3913);
nand U4174 (N_4174,N_3688,N_3593);
or U4175 (N_4175,N_3565,N_3553);
xnor U4176 (N_4176,N_3941,N_3792);
and U4177 (N_4177,N_3821,N_3911);
or U4178 (N_4178,N_3886,N_3999);
and U4179 (N_4179,N_3692,N_3849);
and U4180 (N_4180,N_3774,N_3917);
nand U4181 (N_4181,N_3772,N_3825);
or U4182 (N_4182,N_3997,N_3695);
and U4183 (N_4183,N_3798,N_3643);
xor U4184 (N_4184,N_3690,N_3795);
or U4185 (N_4185,N_3614,N_3938);
nand U4186 (N_4186,N_3808,N_3620);
nand U4187 (N_4187,N_3684,N_3789);
nand U4188 (N_4188,N_3527,N_3784);
and U4189 (N_4189,N_3539,N_3776);
or U4190 (N_4190,N_3619,N_3686);
nor U4191 (N_4191,N_3958,N_3943);
nor U4192 (N_4192,N_3855,N_3866);
or U4193 (N_4193,N_3838,N_3587);
xor U4194 (N_4194,N_3925,N_3762);
xnor U4195 (N_4195,N_3787,N_3703);
nor U4196 (N_4196,N_3508,N_3510);
and U4197 (N_4197,N_3926,N_3505);
nor U4198 (N_4198,N_3715,N_3667);
nand U4199 (N_4199,N_3860,N_3854);
or U4200 (N_4200,N_3831,N_3940);
nor U4201 (N_4201,N_3870,N_3932);
and U4202 (N_4202,N_3755,N_3525);
nor U4203 (N_4203,N_3589,N_3903);
nand U4204 (N_4204,N_3567,N_3696);
nor U4205 (N_4205,N_3647,N_3611);
or U4206 (N_4206,N_3569,N_3531);
nand U4207 (N_4207,N_3828,N_3655);
nor U4208 (N_4208,N_3844,N_3964);
nor U4209 (N_4209,N_3511,N_3530);
or U4210 (N_4210,N_3777,N_3868);
nand U4211 (N_4211,N_3628,N_3952);
or U4212 (N_4212,N_3887,N_3558);
and U4213 (N_4213,N_3664,N_3528);
and U4214 (N_4214,N_3605,N_3946);
nor U4215 (N_4215,N_3699,N_3689);
nor U4216 (N_4216,N_3988,N_3827);
nand U4217 (N_4217,N_3560,N_3549);
and U4218 (N_4218,N_3607,N_3671);
and U4219 (N_4219,N_3598,N_3503);
or U4220 (N_4220,N_3918,N_3641);
nor U4221 (N_4221,N_3839,N_3830);
nor U4222 (N_4222,N_3738,N_3506);
or U4223 (N_4223,N_3745,N_3996);
xnor U4224 (N_4224,N_3594,N_3823);
xnor U4225 (N_4225,N_3563,N_3704);
and U4226 (N_4226,N_3566,N_3824);
and U4227 (N_4227,N_3668,N_3634);
nor U4228 (N_4228,N_3581,N_3840);
nor U4229 (N_4229,N_3573,N_3590);
and U4230 (N_4230,N_3572,N_3760);
nand U4231 (N_4231,N_3916,N_3969);
nor U4232 (N_4232,N_3514,N_3771);
nand U4233 (N_4233,N_3633,N_3523);
nand U4234 (N_4234,N_3603,N_3630);
and U4235 (N_4235,N_3677,N_3736);
nand U4236 (N_4236,N_3806,N_3512);
and U4237 (N_4237,N_3936,N_3644);
nand U4238 (N_4238,N_3963,N_3729);
nand U4239 (N_4239,N_3746,N_3856);
and U4240 (N_4240,N_3766,N_3813);
or U4241 (N_4241,N_3740,N_3694);
or U4242 (N_4242,N_3973,N_3965);
and U4243 (N_4243,N_3862,N_3781);
nand U4244 (N_4244,N_3555,N_3802);
xor U4245 (N_4245,N_3623,N_3884);
nand U4246 (N_4246,N_3951,N_3873);
or U4247 (N_4247,N_3600,N_3935);
nand U4248 (N_4248,N_3616,N_3869);
nor U4249 (N_4249,N_3857,N_3912);
or U4250 (N_4250,N_3769,N_3823);
nor U4251 (N_4251,N_3732,N_3768);
nor U4252 (N_4252,N_3880,N_3644);
nand U4253 (N_4253,N_3614,N_3584);
and U4254 (N_4254,N_3878,N_3993);
nor U4255 (N_4255,N_3687,N_3710);
or U4256 (N_4256,N_3820,N_3722);
nand U4257 (N_4257,N_3553,N_3527);
or U4258 (N_4258,N_3706,N_3799);
or U4259 (N_4259,N_3919,N_3662);
and U4260 (N_4260,N_3855,N_3518);
nor U4261 (N_4261,N_3799,N_3932);
nor U4262 (N_4262,N_3709,N_3946);
nor U4263 (N_4263,N_3709,N_3752);
nand U4264 (N_4264,N_3587,N_3507);
nor U4265 (N_4265,N_3867,N_3961);
xnor U4266 (N_4266,N_3828,N_3725);
nand U4267 (N_4267,N_3924,N_3572);
nand U4268 (N_4268,N_3547,N_3532);
xor U4269 (N_4269,N_3558,N_3980);
xor U4270 (N_4270,N_3521,N_3706);
and U4271 (N_4271,N_3827,N_3899);
nor U4272 (N_4272,N_3644,N_3772);
nand U4273 (N_4273,N_3635,N_3532);
and U4274 (N_4274,N_3577,N_3987);
xnor U4275 (N_4275,N_3850,N_3579);
or U4276 (N_4276,N_3905,N_3734);
xor U4277 (N_4277,N_3797,N_3864);
nor U4278 (N_4278,N_3896,N_3698);
or U4279 (N_4279,N_3807,N_3667);
or U4280 (N_4280,N_3540,N_3974);
and U4281 (N_4281,N_3572,N_3900);
nor U4282 (N_4282,N_3628,N_3661);
and U4283 (N_4283,N_3553,N_3954);
and U4284 (N_4284,N_3774,N_3756);
xor U4285 (N_4285,N_3839,N_3747);
or U4286 (N_4286,N_3900,N_3978);
or U4287 (N_4287,N_3782,N_3994);
nand U4288 (N_4288,N_3944,N_3582);
nand U4289 (N_4289,N_3827,N_3971);
or U4290 (N_4290,N_3646,N_3588);
nand U4291 (N_4291,N_3993,N_3514);
and U4292 (N_4292,N_3634,N_3525);
nor U4293 (N_4293,N_3761,N_3514);
or U4294 (N_4294,N_3607,N_3739);
nor U4295 (N_4295,N_3669,N_3946);
or U4296 (N_4296,N_3772,N_3743);
or U4297 (N_4297,N_3702,N_3825);
xor U4298 (N_4298,N_3755,N_3869);
xor U4299 (N_4299,N_3697,N_3883);
xor U4300 (N_4300,N_3724,N_3966);
or U4301 (N_4301,N_3925,N_3642);
and U4302 (N_4302,N_3753,N_3525);
or U4303 (N_4303,N_3737,N_3551);
and U4304 (N_4304,N_3660,N_3758);
nor U4305 (N_4305,N_3694,N_3732);
and U4306 (N_4306,N_3630,N_3869);
xor U4307 (N_4307,N_3601,N_3500);
nand U4308 (N_4308,N_3674,N_3786);
and U4309 (N_4309,N_3515,N_3674);
or U4310 (N_4310,N_3960,N_3858);
nand U4311 (N_4311,N_3762,N_3742);
nand U4312 (N_4312,N_3744,N_3857);
or U4313 (N_4313,N_3858,N_3618);
xor U4314 (N_4314,N_3949,N_3512);
nand U4315 (N_4315,N_3633,N_3632);
and U4316 (N_4316,N_3611,N_3587);
nand U4317 (N_4317,N_3788,N_3908);
and U4318 (N_4318,N_3986,N_3911);
nor U4319 (N_4319,N_3706,N_3872);
or U4320 (N_4320,N_3825,N_3812);
xor U4321 (N_4321,N_3925,N_3676);
nand U4322 (N_4322,N_3838,N_3719);
or U4323 (N_4323,N_3702,N_3879);
and U4324 (N_4324,N_3988,N_3697);
or U4325 (N_4325,N_3843,N_3621);
or U4326 (N_4326,N_3629,N_3595);
and U4327 (N_4327,N_3950,N_3898);
xnor U4328 (N_4328,N_3555,N_3593);
nor U4329 (N_4329,N_3946,N_3932);
nor U4330 (N_4330,N_3596,N_3581);
and U4331 (N_4331,N_3809,N_3707);
or U4332 (N_4332,N_3665,N_3673);
nor U4333 (N_4333,N_3944,N_3566);
and U4334 (N_4334,N_3667,N_3681);
and U4335 (N_4335,N_3691,N_3639);
nor U4336 (N_4336,N_3953,N_3592);
or U4337 (N_4337,N_3737,N_3755);
or U4338 (N_4338,N_3745,N_3988);
nor U4339 (N_4339,N_3859,N_3649);
nor U4340 (N_4340,N_3529,N_3886);
nor U4341 (N_4341,N_3836,N_3597);
xor U4342 (N_4342,N_3751,N_3892);
nand U4343 (N_4343,N_3808,N_3507);
and U4344 (N_4344,N_3855,N_3655);
xor U4345 (N_4345,N_3850,N_3530);
nor U4346 (N_4346,N_3910,N_3764);
nand U4347 (N_4347,N_3864,N_3571);
nor U4348 (N_4348,N_3974,N_3716);
and U4349 (N_4349,N_3572,N_3948);
and U4350 (N_4350,N_3793,N_3535);
nor U4351 (N_4351,N_3679,N_3970);
and U4352 (N_4352,N_3933,N_3932);
or U4353 (N_4353,N_3679,N_3932);
and U4354 (N_4354,N_3973,N_3983);
or U4355 (N_4355,N_3524,N_3711);
or U4356 (N_4356,N_3994,N_3653);
or U4357 (N_4357,N_3819,N_3799);
and U4358 (N_4358,N_3583,N_3836);
or U4359 (N_4359,N_3589,N_3739);
nand U4360 (N_4360,N_3612,N_3676);
nand U4361 (N_4361,N_3862,N_3885);
nand U4362 (N_4362,N_3773,N_3592);
nor U4363 (N_4363,N_3889,N_3851);
nor U4364 (N_4364,N_3563,N_3999);
and U4365 (N_4365,N_3855,N_3805);
nor U4366 (N_4366,N_3532,N_3804);
nor U4367 (N_4367,N_3777,N_3901);
xor U4368 (N_4368,N_3616,N_3935);
or U4369 (N_4369,N_3862,N_3798);
and U4370 (N_4370,N_3922,N_3663);
nand U4371 (N_4371,N_3835,N_3748);
nand U4372 (N_4372,N_3588,N_3825);
nor U4373 (N_4373,N_3732,N_3639);
nand U4374 (N_4374,N_3503,N_3988);
and U4375 (N_4375,N_3848,N_3778);
and U4376 (N_4376,N_3763,N_3645);
xor U4377 (N_4377,N_3607,N_3630);
and U4378 (N_4378,N_3573,N_3952);
or U4379 (N_4379,N_3641,N_3688);
nor U4380 (N_4380,N_3710,N_3832);
nor U4381 (N_4381,N_3548,N_3708);
nor U4382 (N_4382,N_3755,N_3744);
nand U4383 (N_4383,N_3832,N_3708);
and U4384 (N_4384,N_3672,N_3704);
or U4385 (N_4385,N_3534,N_3637);
nor U4386 (N_4386,N_3584,N_3783);
or U4387 (N_4387,N_3657,N_3921);
or U4388 (N_4388,N_3978,N_3595);
and U4389 (N_4389,N_3919,N_3519);
and U4390 (N_4390,N_3849,N_3609);
or U4391 (N_4391,N_3860,N_3533);
nand U4392 (N_4392,N_3736,N_3631);
xor U4393 (N_4393,N_3803,N_3524);
nand U4394 (N_4394,N_3965,N_3709);
or U4395 (N_4395,N_3986,N_3779);
and U4396 (N_4396,N_3628,N_3970);
or U4397 (N_4397,N_3990,N_3998);
nor U4398 (N_4398,N_3516,N_3945);
or U4399 (N_4399,N_3710,N_3933);
nor U4400 (N_4400,N_3725,N_3567);
nand U4401 (N_4401,N_3714,N_3548);
and U4402 (N_4402,N_3644,N_3647);
and U4403 (N_4403,N_3586,N_3939);
and U4404 (N_4404,N_3735,N_3700);
nand U4405 (N_4405,N_3918,N_3607);
nor U4406 (N_4406,N_3541,N_3514);
or U4407 (N_4407,N_3873,N_3939);
nand U4408 (N_4408,N_3664,N_3544);
nor U4409 (N_4409,N_3810,N_3837);
nor U4410 (N_4410,N_3693,N_3669);
and U4411 (N_4411,N_3551,N_3980);
nand U4412 (N_4412,N_3680,N_3914);
nand U4413 (N_4413,N_3721,N_3754);
or U4414 (N_4414,N_3556,N_3527);
and U4415 (N_4415,N_3994,N_3592);
nand U4416 (N_4416,N_3576,N_3562);
and U4417 (N_4417,N_3939,N_3778);
nor U4418 (N_4418,N_3635,N_3523);
and U4419 (N_4419,N_3566,N_3618);
or U4420 (N_4420,N_3732,N_3670);
xnor U4421 (N_4421,N_3676,N_3532);
and U4422 (N_4422,N_3814,N_3557);
xnor U4423 (N_4423,N_3561,N_3631);
xnor U4424 (N_4424,N_3573,N_3831);
and U4425 (N_4425,N_3976,N_3752);
and U4426 (N_4426,N_3775,N_3796);
nor U4427 (N_4427,N_3918,N_3519);
nor U4428 (N_4428,N_3775,N_3800);
nand U4429 (N_4429,N_3650,N_3915);
nor U4430 (N_4430,N_3942,N_3960);
and U4431 (N_4431,N_3687,N_3658);
nand U4432 (N_4432,N_3573,N_3678);
nor U4433 (N_4433,N_3676,N_3935);
nand U4434 (N_4434,N_3883,N_3631);
nand U4435 (N_4435,N_3842,N_3884);
and U4436 (N_4436,N_3676,N_3552);
or U4437 (N_4437,N_3922,N_3566);
nand U4438 (N_4438,N_3971,N_3929);
nor U4439 (N_4439,N_3777,N_3523);
or U4440 (N_4440,N_3529,N_3883);
xnor U4441 (N_4441,N_3820,N_3690);
and U4442 (N_4442,N_3712,N_3568);
xnor U4443 (N_4443,N_3780,N_3503);
nor U4444 (N_4444,N_3909,N_3633);
nor U4445 (N_4445,N_3689,N_3831);
and U4446 (N_4446,N_3634,N_3913);
or U4447 (N_4447,N_3739,N_3972);
nand U4448 (N_4448,N_3736,N_3909);
xnor U4449 (N_4449,N_3927,N_3985);
nand U4450 (N_4450,N_3766,N_3651);
nor U4451 (N_4451,N_3837,N_3681);
or U4452 (N_4452,N_3505,N_3948);
xor U4453 (N_4453,N_3685,N_3968);
nand U4454 (N_4454,N_3748,N_3953);
nand U4455 (N_4455,N_3817,N_3508);
nor U4456 (N_4456,N_3720,N_3774);
nor U4457 (N_4457,N_3872,N_3633);
nand U4458 (N_4458,N_3619,N_3661);
nand U4459 (N_4459,N_3746,N_3575);
or U4460 (N_4460,N_3538,N_3644);
or U4461 (N_4461,N_3885,N_3657);
nand U4462 (N_4462,N_3709,N_3542);
and U4463 (N_4463,N_3892,N_3596);
or U4464 (N_4464,N_3615,N_3560);
nand U4465 (N_4465,N_3934,N_3747);
and U4466 (N_4466,N_3712,N_3984);
or U4467 (N_4467,N_3779,N_3817);
xnor U4468 (N_4468,N_3745,N_3811);
nor U4469 (N_4469,N_3992,N_3689);
nor U4470 (N_4470,N_3882,N_3570);
nand U4471 (N_4471,N_3770,N_3666);
nor U4472 (N_4472,N_3831,N_3548);
or U4473 (N_4473,N_3649,N_3534);
or U4474 (N_4474,N_3800,N_3873);
xnor U4475 (N_4475,N_3741,N_3743);
and U4476 (N_4476,N_3742,N_3995);
nand U4477 (N_4477,N_3711,N_3586);
and U4478 (N_4478,N_3777,N_3510);
nand U4479 (N_4479,N_3585,N_3580);
and U4480 (N_4480,N_3972,N_3940);
nor U4481 (N_4481,N_3659,N_3618);
and U4482 (N_4482,N_3976,N_3521);
xor U4483 (N_4483,N_3908,N_3566);
nand U4484 (N_4484,N_3923,N_3799);
nor U4485 (N_4485,N_3789,N_3920);
and U4486 (N_4486,N_3877,N_3562);
nand U4487 (N_4487,N_3947,N_3701);
or U4488 (N_4488,N_3640,N_3851);
and U4489 (N_4489,N_3545,N_3603);
and U4490 (N_4490,N_3867,N_3859);
nor U4491 (N_4491,N_3674,N_3871);
nor U4492 (N_4492,N_3937,N_3881);
nand U4493 (N_4493,N_3745,N_3971);
or U4494 (N_4494,N_3862,N_3954);
nor U4495 (N_4495,N_3852,N_3985);
nand U4496 (N_4496,N_3729,N_3519);
and U4497 (N_4497,N_3772,N_3827);
nand U4498 (N_4498,N_3685,N_3993);
or U4499 (N_4499,N_3636,N_3707);
or U4500 (N_4500,N_4236,N_4498);
nor U4501 (N_4501,N_4204,N_4464);
nand U4502 (N_4502,N_4069,N_4368);
or U4503 (N_4503,N_4011,N_4213);
nand U4504 (N_4504,N_4200,N_4243);
nand U4505 (N_4505,N_4296,N_4479);
or U4506 (N_4506,N_4333,N_4397);
or U4507 (N_4507,N_4427,N_4245);
xor U4508 (N_4508,N_4414,N_4266);
and U4509 (N_4509,N_4424,N_4343);
nor U4510 (N_4510,N_4127,N_4254);
nand U4511 (N_4511,N_4218,N_4417);
nor U4512 (N_4512,N_4340,N_4117);
or U4513 (N_4513,N_4138,N_4229);
or U4514 (N_4514,N_4446,N_4175);
nor U4515 (N_4515,N_4308,N_4348);
or U4516 (N_4516,N_4056,N_4119);
nor U4517 (N_4517,N_4231,N_4064);
nor U4518 (N_4518,N_4030,N_4357);
nor U4519 (N_4519,N_4210,N_4410);
or U4520 (N_4520,N_4303,N_4258);
xnor U4521 (N_4521,N_4451,N_4429);
nor U4522 (N_4522,N_4061,N_4361);
nand U4523 (N_4523,N_4112,N_4384);
nor U4524 (N_4524,N_4475,N_4339);
nor U4525 (N_4525,N_4194,N_4096);
or U4526 (N_4526,N_4047,N_4244);
nor U4527 (N_4527,N_4101,N_4201);
nand U4528 (N_4528,N_4419,N_4162);
nand U4529 (N_4529,N_4252,N_4079);
nand U4530 (N_4530,N_4174,N_4264);
and U4531 (N_4531,N_4330,N_4293);
and U4532 (N_4532,N_4452,N_4136);
and U4533 (N_4533,N_4376,N_4437);
nand U4534 (N_4534,N_4355,N_4025);
xnor U4535 (N_4535,N_4040,N_4081);
or U4536 (N_4536,N_4089,N_4251);
and U4537 (N_4537,N_4304,N_4416);
and U4538 (N_4538,N_4278,N_4404);
and U4539 (N_4539,N_4399,N_4386);
or U4540 (N_4540,N_4280,N_4421);
nand U4541 (N_4541,N_4019,N_4151);
or U4542 (N_4542,N_4327,N_4328);
and U4543 (N_4543,N_4158,N_4481);
or U4544 (N_4544,N_4347,N_4234);
and U4545 (N_4545,N_4318,N_4212);
nand U4546 (N_4546,N_4157,N_4380);
nand U4547 (N_4547,N_4302,N_4021);
nor U4548 (N_4548,N_4365,N_4499);
or U4549 (N_4549,N_4338,N_4431);
or U4550 (N_4550,N_4140,N_4250);
xor U4551 (N_4551,N_4354,N_4286);
or U4552 (N_4552,N_4493,N_4482);
nand U4553 (N_4553,N_4197,N_4209);
xor U4554 (N_4554,N_4179,N_4367);
nor U4555 (N_4555,N_4439,N_4316);
and U4556 (N_4556,N_4486,N_4160);
or U4557 (N_4557,N_4432,N_4092);
and U4558 (N_4558,N_4007,N_4467);
or U4559 (N_4559,N_4214,N_4279);
nor U4560 (N_4560,N_4014,N_4309);
nand U4561 (N_4561,N_4088,N_4045);
nor U4562 (N_4562,N_4087,N_4274);
nand U4563 (N_4563,N_4277,N_4120);
nand U4564 (N_4564,N_4332,N_4306);
nand U4565 (N_4565,N_4022,N_4379);
xor U4566 (N_4566,N_4297,N_4108);
nand U4567 (N_4567,N_4059,N_4460);
xnor U4568 (N_4568,N_4001,N_4063);
nor U4569 (N_4569,N_4484,N_4248);
or U4570 (N_4570,N_4456,N_4060);
nand U4571 (N_4571,N_4312,N_4448);
and U4572 (N_4572,N_4445,N_4066);
nor U4573 (N_4573,N_4177,N_4360);
and U4574 (N_4574,N_4294,N_4042);
or U4575 (N_4575,N_4391,N_4492);
xnor U4576 (N_4576,N_4033,N_4185);
or U4577 (N_4577,N_4137,N_4405);
and U4578 (N_4578,N_4170,N_4006);
xnor U4579 (N_4579,N_4104,N_4005);
xor U4580 (N_4580,N_4198,N_4093);
and U4581 (N_4581,N_4054,N_4097);
nor U4582 (N_4582,N_4496,N_4491);
or U4583 (N_4583,N_4166,N_4323);
nand U4584 (N_4584,N_4028,N_4106);
and U4585 (N_4585,N_4370,N_4270);
xor U4586 (N_4586,N_4390,N_4024);
nand U4587 (N_4587,N_4130,N_4366);
nand U4588 (N_4588,N_4186,N_4238);
xnor U4589 (N_4589,N_4053,N_4009);
or U4590 (N_4590,N_4271,N_4267);
xor U4591 (N_4591,N_4346,N_4122);
nor U4592 (N_4592,N_4462,N_4301);
nand U4593 (N_4593,N_4383,N_4159);
nor U4594 (N_4594,N_4415,N_4099);
and U4595 (N_4595,N_4283,N_4129);
xnor U4596 (N_4596,N_4242,N_4072);
nor U4597 (N_4597,N_4291,N_4351);
nor U4598 (N_4598,N_4016,N_4412);
nor U4599 (N_4599,N_4123,N_4110);
nand U4600 (N_4600,N_4259,N_4071);
nor U4601 (N_4601,N_4191,N_4461);
nand U4602 (N_4602,N_4468,N_4490);
xnor U4603 (N_4603,N_4165,N_4473);
xor U4604 (N_4604,N_4438,N_4409);
nor U4605 (N_4605,N_4241,N_4422);
nand U4606 (N_4606,N_4223,N_4337);
xor U4607 (N_4607,N_4457,N_4196);
and U4608 (N_4608,N_4288,N_4319);
nand U4609 (N_4609,N_4483,N_4034);
and U4610 (N_4610,N_4075,N_4115);
nor U4611 (N_4611,N_4239,N_4406);
or U4612 (N_4612,N_4026,N_4077);
and U4613 (N_4613,N_4444,N_4181);
nor U4614 (N_4614,N_4388,N_4008);
and U4615 (N_4615,N_4114,N_4336);
or U4616 (N_4616,N_4413,N_4341);
and U4617 (N_4617,N_4396,N_4334);
or U4618 (N_4618,N_4046,N_4113);
or U4619 (N_4619,N_4374,N_4272);
or U4620 (N_4620,N_4173,N_4225);
nor U4621 (N_4621,N_4135,N_4103);
nor U4622 (N_4622,N_4434,N_4168);
xor U4623 (N_4623,N_4472,N_4260);
nor U4624 (N_4624,N_4495,N_4377);
or U4625 (N_4625,N_4172,N_4356);
or U4626 (N_4626,N_4139,N_4287);
or U4627 (N_4627,N_4230,N_4176);
nor U4628 (N_4628,N_4070,N_4441);
or U4629 (N_4629,N_4335,N_4268);
or U4630 (N_4630,N_4344,N_4015);
or U4631 (N_4631,N_4211,N_4124);
or U4632 (N_4632,N_4039,N_4065);
nand U4633 (N_4633,N_4220,N_4382);
or U4634 (N_4634,N_4023,N_4048);
and U4635 (N_4635,N_4217,N_4420);
or U4636 (N_4636,N_4320,N_4480);
or U4637 (N_4637,N_4385,N_4400);
xnor U4638 (N_4638,N_4055,N_4305);
or U4639 (N_4639,N_4208,N_4222);
nor U4640 (N_4640,N_4202,N_4289);
nand U4641 (N_4641,N_4010,N_4269);
or U4642 (N_4642,N_4035,N_4311);
nor U4643 (N_4643,N_4276,N_4450);
and U4644 (N_4644,N_4128,N_4036);
and U4645 (N_4645,N_4371,N_4255);
and U4646 (N_4646,N_4310,N_4164);
xor U4647 (N_4647,N_4118,N_4192);
nand U4648 (N_4648,N_4183,N_4116);
nand U4649 (N_4649,N_4262,N_4362);
nor U4650 (N_4650,N_4156,N_4256);
nor U4651 (N_4651,N_4083,N_4322);
xor U4652 (N_4652,N_4050,N_4109);
nand U4653 (N_4653,N_4246,N_4433);
or U4654 (N_4654,N_4052,N_4029);
nor U4655 (N_4655,N_4263,N_4076);
and U4656 (N_4656,N_4349,N_4017);
nor U4657 (N_4657,N_4161,N_4000);
xnor U4658 (N_4658,N_4307,N_4426);
nor U4659 (N_4659,N_4418,N_4084);
and U4660 (N_4660,N_4085,N_4195);
xnor U4661 (N_4661,N_4369,N_4466);
or U4662 (N_4662,N_4375,N_4131);
and U4663 (N_4663,N_4193,N_4350);
nand U4664 (N_4664,N_4150,N_4411);
xor U4665 (N_4665,N_4068,N_4402);
or U4666 (N_4666,N_4363,N_4227);
or U4667 (N_4667,N_4455,N_4149);
nand U4668 (N_4668,N_4002,N_4216);
or U4669 (N_4669,N_4141,N_4342);
nand U4670 (N_4670,N_4265,N_4485);
and U4671 (N_4671,N_4273,N_4003);
nor U4672 (N_4672,N_4126,N_4121);
or U4673 (N_4673,N_4440,N_4474);
xnor U4674 (N_4674,N_4074,N_4031);
nor U4675 (N_4675,N_4378,N_4094);
nand U4676 (N_4676,N_4142,N_4465);
xor U4677 (N_4677,N_4423,N_4261);
nor U4678 (N_4678,N_4098,N_4476);
nand U4679 (N_4679,N_4314,N_4487);
and U4680 (N_4680,N_4295,N_4290);
nand U4681 (N_4681,N_4215,N_4169);
or U4682 (N_4682,N_4407,N_4020);
nor U4683 (N_4683,N_4292,N_4178);
or U4684 (N_4684,N_4073,N_4315);
nand U4685 (N_4685,N_4298,N_4107);
and U4686 (N_4686,N_4488,N_4373);
nor U4687 (N_4687,N_4027,N_4253);
nor U4688 (N_4688,N_4051,N_4032);
nor U4689 (N_4689,N_4326,N_4435);
nor U4690 (N_4690,N_4086,N_4043);
nand U4691 (N_4691,N_4387,N_4300);
xnor U4692 (N_4692,N_4228,N_4358);
and U4693 (N_4693,N_4247,N_4233);
or U4694 (N_4694,N_4313,N_4329);
and U4695 (N_4695,N_4147,N_4205);
and U4696 (N_4696,N_4062,N_4299);
xnor U4697 (N_4697,N_4189,N_4459);
or U4698 (N_4698,N_4470,N_4044);
nand U4699 (N_4699,N_4317,N_4240);
nor U4700 (N_4700,N_4359,N_4154);
nor U4701 (N_4701,N_4257,N_4067);
nand U4702 (N_4702,N_4408,N_4188);
or U4703 (N_4703,N_4389,N_4180);
nand U4704 (N_4704,N_4324,N_4478);
or U4705 (N_4705,N_4454,N_4443);
and U4706 (N_4706,N_4224,N_4232);
nor U4707 (N_4707,N_4012,N_4494);
xnor U4708 (N_4708,N_4038,N_4249);
xor U4709 (N_4709,N_4133,N_4425);
xnor U4710 (N_4710,N_4325,N_4235);
and U4711 (N_4711,N_4187,N_4497);
and U4712 (N_4712,N_4458,N_4226);
or U4713 (N_4713,N_4393,N_4144);
xor U4714 (N_4714,N_4285,N_4364);
nor U4715 (N_4715,N_4004,N_4403);
nand U4716 (N_4716,N_4281,N_4013);
nor U4717 (N_4717,N_4207,N_4155);
nand U4718 (N_4718,N_4447,N_4352);
nand U4719 (N_4719,N_4221,N_4398);
nor U4720 (N_4720,N_4163,N_4284);
or U4721 (N_4721,N_4353,N_4078);
nand U4722 (N_4722,N_4105,N_4469);
or U4723 (N_4723,N_4184,N_4381);
or U4724 (N_4724,N_4111,N_4102);
or U4725 (N_4725,N_4321,N_4082);
nand U4726 (N_4726,N_4430,N_4090);
and U4727 (N_4727,N_4132,N_4428);
nor U4728 (N_4728,N_4018,N_4152);
or U4729 (N_4729,N_4190,N_4057);
nor U4730 (N_4730,N_4146,N_4394);
or U4731 (N_4731,N_4219,N_4489);
nand U4732 (N_4732,N_4091,N_4041);
or U4733 (N_4733,N_4100,N_4171);
nand U4734 (N_4734,N_4275,N_4372);
or U4735 (N_4735,N_4182,N_4442);
nor U4736 (N_4736,N_4148,N_4153);
and U4737 (N_4737,N_4134,N_4095);
nor U4738 (N_4738,N_4449,N_4436);
nand U4739 (N_4739,N_4145,N_4477);
nor U4740 (N_4740,N_4167,N_4206);
nand U4741 (N_4741,N_4401,N_4199);
nor U4742 (N_4742,N_4331,N_4203);
nand U4743 (N_4743,N_4037,N_4395);
nor U4744 (N_4744,N_4143,N_4471);
and U4745 (N_4745,N_4058,N_4345);
and U4746 (N_4746,N_4237,N_4282);
or U4747 (N_4747,N_4125,N_4080);
nand U4748 (N_4748,N_4392,N_4453);
nor U4749 (N_4749,N_4049,N_4463);
or U4750 (N_4750,N_4004,N_4210);
nand U4751 (N_4751,N_4179,N_4294);
nand U4752 (N_4752,N_4390,N_4242);
nor U4753 (N_4753,N_4336,N_4108);
nand U4754 (N_4754,N_4205,N_4213);
or U4755 (N_4755,N_4126,N_4423);
nand U4756 (N_4756,N_4123,N_4496);
nand U4757 (N_4757,N_4324,N_4354);
nand U4758 (N_4758,N_4138,N_4145);
or U4759 (N_4759,N_4047,N_4277);
and U4760 (N_4760,N_4125,N_4496);
nand U4761 (N_4761,N_4463,N_4074);
nor U4762 (N_4762,N_4434,N_4356);
or U4763 (N_4763,N_4265,N_4461);
and U4764 (N_4764,N_4497,N_4015);
nand U4765 (N_4765,N_4433,N_4007);
nand U4766 (N_4766,N_4432,N_4143);
or U4767 (N_4767,N_4407,N_4090);
xnor U4768 (N_4768,N_4122,N_4384);
or U4769 (N_4769,N_4138,N_4473);
and U4770 (N_4770,N_4181,N_4022);
nand U4771 (N_4771,N_4256,N_4288);
and U4772 (N_4772,N_4266,N_4187);
and U4773 (N_4773,N_4223,N_4483);
nand U4774 (N_4774,N_4056,N_4421);
and U4775 (N_4775,N_4172,N_4166);
nor U4776 (N_4776,N_4280,N_4087);
and U4777 (N_4777,N_4160,N_4125);
xor U4778 (N_4778,N_4287,N_4027);
and U4779 (N_4779,N_4167,N_4268);
nor U4780 (N_4780,N_4271,N_4184);
xnor U4781 (N_4781,N_4194,N_4140);
nand U4782 (N_4782,N_4191,N_4280);
or U4783 (N_4783,N_4017,N_4121);
nand U4784 (N_4784,N_4385,N_4350);
xnor U4785 (N_4785,N_4066,N_4497);
xor U4786 (N_4786,N_4327,N_4261);
xor U4787 (N_4787,N_4287,N_4488);
and U4788 (N_4788,N_4054,N_4076);
and U4789 (N_4789,N_4099,N_4325);
nor U4790 (N_4790,N_4403,N_4117);
nand U4791 (N_4791,N_4153,N_4365);
or U4792 (N_4792,N_4218,N_4254);
or U4793 (N_4793,N_4473,N_4279);
xor U4794 (N_4794,N_4419,N_4111);
nor U4795 (N_4795,N_4189,N_4363);
nand U4796 (N_4796,N_4128,N_4460);
and U4797 (N_4797,N_4116,N_4496);
nand U4798 (N_4798,N_4357,N_4017);
nor U4799 (N_4799,N_4466,N_4215);
xor U4800 (N_4800,N_4072,N_4159);
nor U4801 (N_4801,N_4030,N_4234);
nand U4802 (N_4802,N_4232,N_4386);
nand U4803 (N_4803,N_4098,N_4241);
nand U4804 (N_4804,N_4030,N_4210);
nand U4805 (N_4805,N_4478,N_4177);
and U4806 (N_4806,N_4347,N_4350);
nor U4807 (N_4807,N_4359,N_4113);
nand U4808 (N_4808,N_4301,N_4349);
nor U4809 (N_4809,N_4496,N_4161);
and U4810 (N_4810,N_4314,N_4079);
nor U4811 (N_4811,N_4371,N_4282);
or U4812 (N_4812,N_4233,N_4463);
or U4813 (N_4813,N_4369,N_4353);
or U4814 (N_4814,N_4390,N_4159);
and U4815 (N_4815,N_4140,N_4323);
xnor U4816 (N_4816,N_4492,N_4428);
nand U4817 (N_4817,N_4068,N_4247);
or U4818 (N_4818,N_4398,N_4137);
nand U4819 (N_4819,N_4213,N_4176);
and U4820 (N_4820,N_4475,N_4130);
or U4821 (N_4821,N_4444,N_4459);
nand U4822 (N_4822,N_4452,N_4065);
and U4823 (N_4823,N_4011,N_4338);
or U4824 (N_4824,N_4126,N_4028);
nor U4825 (N_4825,N_4346,N_4482);
nand U4826 (N_4826,N_4111,N_4179);
or U4827 (N_4827,N_4391,N_4432);
or U4828 (N_4828,N_4290,N_4425);
nor U4829 (N_4829,N_4018,N_4127);
nor U4830 (N_4830,N_4236,N_4309);
or U4831 (N_4831,N_4445,N_4324);
and U4832 (N_4832,N_4215,N_4294);
nor U4833 (N_4833,N_4471,N_4266);
and U4834 (N_4834,N_4098,N_4274);
or U4835 (N_4835,N_4466,N_4186);
and U4836 (N_4836,N_4441,N_4476);
nor U4837 (N_4837,N_4043,N_4301);
or U4838 (N_4838,N_4399,N_4371);
nand U4839 (N_4839,N_4089,N_4091);
nand U4840 (N_4840,N_4079,N_4131);
xor U4841 (N_4841,N_4172,N_4261);
nor U4842 (N_4842,N_4302,N_4395);
nand U4843 (N_4843,N_4220,N_4457);
and U4844 (N_4844,N_4274,N_4282);
nor U4845 (N_4845,N_4192,N_4126);
and U4846 (N_4846,N_4211,N_4382);
and U4847 (N_4847,N_4281,N_4458);
or U4848 (N_4848,N_4332,N_4301);
and U4849 (N_4849,N_4327,N_4385);
or U4850 (N_4850,N_4064,N_4343);
xor U4851 (N_4851,N_4349,N_4129);
or U4852 (N_4852,N_4179,N_4194);
or U4853 (N_4853,N_4013,N_4359);
and U4854 (N_4854,N_4249,N_4000);
xor U4855 (N_4855,N_4068,N_4302);
or U4856 (N_4856,N_4116,N_4162);
and U4857 (N_4857,N_4363,N_4442);
nand U4858 (N_4858,N_4078,N_4030);
nand U4859 (N_4859,N_4436,N_4065);
nand U4860 (N_4860,N_4284,N_4291);
and U4861 (N_4861,N_4081,N_4137);
or U4862 (N_4862,N_4160,N_4336);
or U4863 (N_4863,N_4473,N_4054);
nand U4864 (N_4864,N_4029,N_4010);
nor U4865 (N_4865,N_4229,N_4443);
or U4866 (N_4866,N_4355,N_4089);
and U4867 (N_4867,N_4320,N_4074);
nand U4868 (N_4868,N_4466,N_4071);
or U4869 (N_4869,N_4161,N_4236);
nand U4870 (N_4870,N_4318,N_4031);
nand U4871 (N_4871,N_4176,N_4333);
and U4872 (N_4872,N_4180,N_4136);
nand U4873 (N_4873,N_4118,N_4041);
nand U4874 (N_4874,N_4181,N_4244);
nand U4875 (N_4875,N_4332,N_4374);
and U4876 (N_4876,N_4402,N_4203);
and U4877 (N_4877,N_4446,N_4083);
and U4878 (N_4878,N_4153,N_4156);
and U4879 (N_4879,N_4383,N_4414);
nand U4880 (N_4880,N_4267,N_4117);
and U4881 (N_4881,N_4138,N_4409);
and U4882 (N_4882,N_4496,N_4152);
or U4883 (N_4883,N_4371,N_4023);
or U4884 (N_4884,N_4145,N_4202);
and U4885 (N_4885,N_4345,N_4437);
nor U4886 (N_4886,N_4405,N_4017);
xor U4887 (N_4887,N_4369,N_4269);
or U4888 (N_4888,N_4124,N_4031);
and U4889 (N_4889,N_4056,N_4355);
nand U4890 (N_4890,N_4156,N_4351);
and U4891 (N_4891,N_4441,N_4392);
or U4892 (N_4892,N_4484,N_4188);
or U4893 (N_4893,N_4305,N_4129);
nor U4894 (N_4894,N_4357,N_4228);
or U4895 (N_4895,N_4048,N_4349);
nand U4896 (N_4896,N_4198,N_4499);
nor U4897 (N_4897,N_4114,N_4461);
nand U4898 (N_4898,N_4053,N_4477);
nor U4899 (N_4899,N_4332,N_4175);
and U4900 (N_4900,N_4318,N_4485);
xor U4901 (N_4901,N_4228,N_4189);
nand U4902 (N_4902,N_4143,N_4079);
or U4903 (N_4903,N_4041,N_4086);
nand U4904 (N_4904,N_4251,N_4241);
or U4905 (N_4905,N_4268,N_4336);
nand U4906 (N_4906,N_4106,N_4036);
or U4907 (N_4907,N_4116,N_4294);
xnor U4908 (N_4908,N_4275,N_4033);
nand U4909 (N_4909,N_4153,N_4212);
xor U4910 (N_4910,N_4130,N_4146);
and U4911 (N_4911,N_4362,N_4120);
or U4912 (N_4912,N_4127,N_4272);
nand U4913 (N_4913,N_4384,N_4172);
nor U4914 (N_4914,N_4204,N_4170);
nand U4915 (N_4915,N_4349,N_4401);
or U4916 (N_4916,N_4354,N_4108);
nor U4917 (N_4917,N_4356,N_4241);
nor U4918 (N_4918,N_4146,N_4496);
and U4919 (N_4919,N_4230,N_4418);
and U4920 (N_4920,N_4157,N_4340);
nand U4921 (N_4921,N_4002,N_4059);
nor U4922 (N_4922,N_4495,N_4257);
nand U4923 (N_4923,N_4020,N_4136);
nor U4924 (N_4924,N_4405,N_4276);
nor U4925 (N_4925,N_4442,N_4379);
or U4926 (N_4926,N_4355,N_4088);
nor U4927 (N_4927,N_4314,N_4051);
or U4928 (N_4928,N_4439,N_4458);
nor U4929 (N_4929,N_4362,N_4015);
nand U4930 (N_4930,N_4487,N_4133);
or U4931 (N_4931,N_4151,N_4242);
xor U4932 (N_4932,N_4192,N_4441);
and U4933 (N_4933,N_4346,N_4218);
nand U4934 (N_4934,N_4007,N_4314);
nand U4935 (N_4935,N_4353,N_4223);
nor U4936 (N_4936,N_4249,N_4302);
nand U4937 (N_4937,N_4270,N_4017);
nor U4938 (N_4938,N_4040,N_4181);
nand U4939 (N_4939,N_4034,N_4452);
or U4940 (N_4940,N_4336,N_4444);
nand U4941 (N_4941,N_4201,N_4470);
nand U4942 (N_4942,N_4339,N_4307);
or U4943 (N_4943,N_4454,N_4103);
and U4944 (N_4944,N_4338,N_4294);
nor U4945 (N_4945,N_4412,N_4105);
or U4946 (N_4946,N_4111,N_4355);
and U4947 (N_4947,N_4437,N_4155);
nor U4948 (N_4948,N_4431,N_4262);
or U4949 (N_4949,N_4460,N_4067);
nor U4950 (N_4950,N_4415,N_4290);
or U4951 (N_4951,N_4468,N_4238);
or U4952 (N_4952,N_4444,N_4410);
nor U4953 (N_4953,N_4464,N_4305);
nor U4954 (N_4954,N_4226,N_4076);
nor U4955 (N_4955,N_4166,N_4023);
xnor U4956 (N_4956,N_4359,N_4138);
xor U4957 (N_4957,N_4050,N_4403);
nor U4958 (N_4958,N_4296,N_4067);
and U4959 (N_4959,N_4442,N_4163);
nor U4960 (N_4960,N_4064,N_4191);
xnor U4961 (N_4961,N_4214,N_4176);
nand U4962 (N_4962,N_4183,N_4486);
or U4963 (N_4963,N_4351,N_4474);
or U4964 (N_4964,N_4468,N_4345);
or U4965 (N_4965,N_4336,N_4010);
and U4966 (N_4966,N_4251,N_4466);
xor U4967 (N_4967,N_4268,N_4055);
or U4968 (N_4968,N_4051,N_4493);
xor U4969 (N_4969,N_4409,N_4460);
or U4970 (N_4970,N_4144,N_4402);
and U4971 (N_4971,N_4105,N_4290);
nand U4972 (N_4972,N_4288,N_4295);
nand U4973 (N_4973,N_4340,N_4053);
nor U4974 (N_4974,N_4304,N_4340);
nor U4975 (N_4975,N_4241,N_4162);
or U4976 (N_4976,N_4384,N_4141);
and U4977 (N_4977,N_4042,N_4121);
or U4978 (N_4978,N_4078,N_4124);
nor U4979 (N_4979,N_4482,N_4004);
or U4980 (N_4980,N_4265,N_4373);
and U4981 (N_4981,N_4155,N_4154);
nand U4982 (N_4982,N_4234,N_4432);
and U4983 (N_4983,N_4266,N_4215);
xnor U4984 (N_4984,N_4017,N_4063);
xor U4985 (N_4985,N_4201,N_4317);
nand U4986 (N_4986,N_4241,N_4312);
nand U4987 (N_4987,N_4265,N_4336);
nand U4988 (N_4988,N_4302,N_4441);
nand U4989 (N_4989,N_4244,N_4420);
nand U4990 (N_4990,N_4280,N_4002);
and U4991 (N_4991,N_4133,N_4032);
nor U4992 (N_4992,N_4295,N_4421);
nor U4993 (N_4993,N_4275,N_4325);
and U4994 (N_4994,N_4308,N_4058);
nor U4995 (N_4995,N_4080,N_4384);
nor U4996 (N_4996,N_4208,N_4162);
and U4997 (N_4997,N_4292,N_4057);
or U4998 (N_4998,N_4439,N_4359);
nand U4999 (N_4999,N_4068,N_4363);
or U5000 (N_5000,N_4520,N_4673);
and U5001 (N_5001,N_4537,N_4879);
nor U5002 (N_5002,N_4581,N_4885);
or U5003 (N_5003,N_4941,N_4994);
or U5004 (N_5004,N_4844,N_4670);
or U5005 (N_5005,N_4672,N_4764);
and U5006 (N_5006,N_4899,N_4725);
nor U5007 (N_5007,N_4930,N_4731);
nand U5008 (N_5008,N_4538,N_4948);
nor U5009 (N_5009,N_4593,N_4977);
and U5010 (N_5010,N_4740,N_4522);
nand U5011 (N_5011,N_4821,N_4540);
xnor U5012 (N_5012,N_4727,N_4636);
nand U5013 (N_5013,N_4949,N_4648);
or U5014 (N_5014,N_4996,N_4788);
and U5015 (N_5015,N_4596,N_4738);
nor U5016 (N_5016,N_4528,N_4586);
or U5017 (N_5017,N_4660,N_4790);
or U5018 (N_5018,N_4912,N_4598);
nor U5019 (N_5019,N_4797,N_4810);
nor U5020 (N_5020,N_4524,N_4976);
and U5021 (N_5021,N_4779,N_4978);
and U5022 (N_5022,N_4862,N_4867);
or U5023 (N_5023,N_4804,N_4865);
xor U5024 (N_5024,N_4917,N_4756);
and U5025 (N_5025,N_4525,N_4892);
xnor U5026 (N_5026,N_4502,N_4795);
nand U5027 (N_5027,N_4608,N_4778);
and U5028 (N_5028,N_4572,N_4995);
or U5029 (N_5029,N_4989,N_4604);
and U5030 (N_5030,N_4927,N_4871);
or U5031 (N_5031,N_4551,N_4699);
nor U5032 (N_5032,N_4702,N_4816);
nand U5033 (N_5033,N_4814,N_4840);
nor U5034 (N_5034,N_4513,N_4590);
nand U5035 (N_5035,N_4801,N_4546);
and U5036 (N_5036,N_4591,N_4721);
or U5037 (N_5037,N_4761,N_4559);
or U5038 (N_5038,N_4896,N_4822);
or U5039 (N_5039,N_4951,N_4883);
xor U5040 (N_5040,N_4713,N_4835);
and U5041 (N_5041,N_4534,N_4645);
or U5042 (N_5042,N_4915,N_4594);
or U5043 (N_5043,N_4619,N_4923);
and U5044 (N_5044,N_4881,N_4985);
nor U5045 (N_5045,N_4858,N_4786);
nand U5046 (N_5046,N_4652,N_4580);
nand U5047 (N_5047,N_4578,N_4846);
nor U5048 (N_5048,N_4884,N_4588);
nor U5049 (N_5049,N_4857,N_4831);
and U5050 (N_5050,N_4733,N_4664);
nand U5051 (N_5051,N_4654,N_4806);
xnor U5052 (N_5052,N_4514,N_4919);
xor U5053 (N_5053,N_4511,N_4599);
or U5054 (N_5054,N_4837,N_4724);
xor U5055 (N_5055,N_4568,N_4753);
and U5056 (N_5056,N_4549,N_4613);
and U5057 (N_5057,N_4757,N_4911);
nand U5058 (N_5058,N_4722,N_4628);
or U5059 (N_5059,N_4841,N_4752);
or U5060 (N_5060,N_4880,N_4834);
or U5061 (N_5061,N_4970,N_4589);
or U5062 (N_5062,N_4610,N_4979);
or U5063 (N_5063,N_4928,N_4703);
nor U5064 (N_5064,N_4950,N_4820);
and U5065 (N_5065,N_4802,N_4798);
and U5066 (N_5066,N_4907,N_4886);
or U5067 (N_5067,N_4799,N_4662);
nand U5068 (N_5068,N_4633,N_4829);
xnor U5069 (N_5069,N_4629,N_4607);
nor U5070 (N_5070,N_4614,N_4624);
nand U5071 (N_5071,N_4621,N_4512);
or U5072 (N_5072,N_4770,N_4947);
and U5073 (N_5073,N_4620,N_4500);
or U5074 (N_5074,N_4640,N_4789);
nand U5075 (N_5075,N_4712,N_4584);
and U5076 (N_5076,N_4671,N_4611);
xor U5077 (N_5077,N_4973,N_4574);
nor U5078 (N_5078,N_4649,N_4940);
xor U5079 (N_5079,N_4582,N_4527);
or U5080 (N_5080,N_4560,N_4587);
nor U5081 (N_5081,N_4554,N_4931);
or U5082 (N_5082,N_4632,N_4683);
nor U5083 (N_5083,N_4811,N_4603);
and U5084 (N_5084,N_4987,N_4792);
nor U5085 (N_5085,N_4762,N_4661);
nor U5086 (N_5086,N_4622,N_4925);
or U5087 (N_5087,N_4895,N_4592);
and U5088 (N_5088,N_4818,N_4505);
xor U5089 (N_5089,N_4663,N_4533);
or U5090 (N_5090,N_4882,N_4914);
or U5091 (N_5091,N_4737,N_4746);
xnor U5092 (N_5092,N_4791,N_4817);
xnor U5093 (N_5093,N_4557,N_4877);
nand U5094 (N_5094,N_4743,N_4552);
nor U5095 (N_5095,N_4616,N_4718);
nand U5096 (N_5096,N_4609,N_4859);
nand U5097 (N_5097,N_4891,N_4894);
and U5098 (N_5098,N_4863,N_4965);
and U5099 (N_5099,N_4583,N_4576);
and U5100 (N_5100,N_4952,N_4523);
nand U5101 (N_5101,N_4787,N_4860);
or U5102 (N_5102,N_4675,N_4953);
nand U5103 (N_5103,N_4959,N_4769);
nor U5104 (N_5104,N_4984,N_4807);
nor U5105 (N_5105,N_4929,N_4676);
or U5106 (N_5106,N_4575,N_4605);
nand U5107 (N_5107,N_4689,N_4908);
or U5108 (N_5108,N_4966,N_4749);
or U5109 (N_5109,N_4601,N_4838);
nand U5110 (N_5110,N_4874,N_4680);
nand U5111 (N_5111,N_4830,N_4755);
nor U5112 (N_5112,N_4845,N_4937);
and U5113 (N_5113,N_4839,N_4750);
nand U5114 (N_5114,N_4700,N_4531);
nand U5115 (N_5115,N_4667,N_4626);
nand U5116 (N_5116,N_4707,N_4615);
or U5117 (N_5117,N_4665,N_4843);
nand U5118 (N_5118,N_4674,N_4847);
and U5119 (N_5119,N_4736,N_4999);
or U5120 (N_5120,N_4735,N_4944);
nor U5121 (N_5121,N_4720,N_4658);
or U5122 (N_5122,N_4964,N_4541);
nor U5123 (N_5123,N_4630,N_4530);
or U5124 (N_5124,N_4741,N_4759);
and U5125 (N_5125,N_4905,N_4766);
nand U5126 (N_5126,N_4517,N_4553);
xor U5127 (N_5127,N_4805,N_4955);
xor U5128 (N_5128,N_4852,N_4744);
nand U5129 (N_5129,N_4618,N_4641);
or U5130 (N_5130,N_4679,N_4783);
or U5131 (N_5131,N_4571,N_4967);
nor U5132 (N_5132,N_4714,N_4800);
and U5133 (N_5133,N_4569,N_4784);
and U5134 (N_5134,N_4920,N_4723);
xnor U5135 (N_5135,N_4861,N_4544);
and U5136 (N_5136,N_4813,N_4656);
nand U5137 (N_5137,N_4539,N_4849);
nor U5138 (N_5138,N_4958,N_4657);
xnor U5139 (N_5139,N_4754,N_4809);
and U5140 (N_5140,N_4600,N_4542);
and U5141 (N_5141,N_4774,N_4988);
nand U5142 (N_5142,N_4803,N_4545);
xnor U5143 (N_5143,N_4906,N_4748);
and U5144 (N_5144,N_4668,N_4824);
or U5145 (N_5145,N_4711,N_4701);
or U5146 (N_5146,N_4706,N_4926);
xor U5147 (N_5147,N_4682,N_4518);
nor U5148 (N_5148,N_4825,N_4691);
nand U5149 (N_5149,N_4781,N_4932);
or U5150 (N_5150,N_4564,N_4924);
nor U5151 (N_5151,N_4643,N_4828);
and U5152 (N_5152,N_4793,N_4634);
nand U5153 (N_5153,N_4776,N_4509);
nand U5154 (N_5154,N_4943,N_4921);
nand U5155 (N_5155,N_4901,N_4550);
or U5156 (N_5156,N_4773,N_4563);
xor U5157 (N_5157,N_4644,N_4902);
and U5158 (N_5158,N_4742,N_4510);
nand U5159 (N_5159,N_4728,N_4870);
xnor U5160 (N_5160,N_4638,N_4939);
and U5161 (N_5161,N_4697,N_4516);
xnor U5162 (N_5162,N_4515,N_4850);
xor U5163 (N_5163,N_4606,N_4957);
xor U5164 (N_5164,N_4916,N_4595);
and U5165 (N_5165,N_4782,N_4710);
nor U5166 (N_5166,N_4536,N_4688);
nor U5167 (N_5167,N_4526,N_4687);
nand U5168 (N_5168,N_4653,N_4956);
nor U5169 (N_5169,N_4692,N_4767);
nor U5170 (N_5170,N_4719,N_4819);
nor U5171 (N_5171,N_4888,N_4935);
nand U5172 (N_5172,N_4729,N_4686);
and U5173 (N_5173,N_4836,N_4684);
xnor U5174 (N_5174,N_4960,N_4565);
nor U5175 (N_5175,N_4936,N_4796);
xnor U5176 (N_5176,N_4969,N_4772);
nand U5177 (N_5177,N_4758,N_4981);
xnor U5178 (N_5178,N_4585,N_4982);
nand U5179 (N_5179,N_4543,N_4647);
nand U5180 (N_5180,N_4961,N_4659);
nand U5181 (N_5181,N_4826,N_4922);
and U5182 (N_5182,N_4780,N_4685);
nor U5183 (N_5183,N_4872,N_4579);
and U5184 (N_5184,N_4751,N_4875);
nand U5185 (N_5185,N_4763,N_4997);
nor U5186 (N_5186,N_4873,N_4681);
or U5187 (N_5187,N_4506,N_4558);
nor U5188 (N_5188,N_4887,N_4851);
nand U5189 (N_5189,N_4745,N_4693);
and U5190 (N_5190,N_4827,N_4716);
and U5191 (N_5191,N_4768,N_4876);
xnor U5192 (N_5192,N_4678,N_4808);
nand U5193 (N_5193,N_4785,N_4993);
or U5194 (N_5194,N_4890,N_4651);
or U5195 (N_5195,N_4991,N_4532);
nor U5196 (N_5196,N_4507,N_4739);
nor U5197 (N_5197,N_4573,N_4562);
or U5198 (N_5198,N_4698,N_4848);
xnor U5199 (N_5199,N_4567,N_4968);
or U5200 (N_5200,N_4503,N_4566);
or U5201 (N_5201,N_4962,N_4535);
or U5202 (N_5202,N_4529,N_4696);
nand U5203 (N_5203,N_4631,N_4519);
and U5204 (N_5204,N_4878,N_4864);
or U5205 (N_5205,N_4971,N_4732);
and U5206 (N_5206,N_4889,N_4909);
nand U5207 (N_5207,N_4655,N_4504);
or U5208 (N_5208,N_4717,N_4715);
nor U5209 (N_5209,N_4635,N_4646);
and U5210 (N_5210,N_4898,N_4547);
nand U5211 (N_5211,N_4910,N_4760);
and U5212 (N_5212,N_4556,N_4650);
nand U5213 (N_5213,N_4974,N_4866);
xor U5214 (N_5214,N_4856,N_4521);
nand U5215 (N_5215,N_4639,N_4708);
nor U5216 (N_5216,N_4855,N_4555);
or U5217 (N_5217,N_4998,N_4734);
and U5218 (N_5218,N_4868,N_4617);
nand U5219 (N_5219,N_4602,N_4669);
nand U5220 (N_5220,N_4854,N_4642);
nor U5221 (N_5221,N_4900,N_4869);
nor U5222 (N_5222,N_4934,N_4501);
nor U5223 (N_5223,N_4980,N_4815);
nand U5224 (N_5224,N_4986,N_4666);
and U5225 (N_5225,N_4983,N_4903);
or U5226 (N_5226,N_4777,N_4933);
or U5227 (N_5227,N_4942,N_4833);
nor U5228 (N_5228,N_4690,N_4775);
nand U5229 (N_5229,N_4508,N_4945);
and U5230 (N_5230,N_4597,N_4897);
and U5231 (N_5231,N_4637,N_4577);
or U5232 (N_5232,N_4694,N_4726);
and U5233 (N_5233,N_4704,N_4730);
or U5234 (N_5234,N_4842,N_4561);
nor U5235 (N_5235,N_4954,N_4705);
or U5236 (N_5236,N_4938,N_4990);
or U5237 (N_5237,N_4823,N_4832);
xor U5238 (N_5238,N_4946,N_4709);
or U5239 (N_5239,N_4963,N_4904);
or U5240 (N_5240,N_4893,N_4794);
or U5241 (N_5241,N_4913,N_4548);
nor U5242 (N_5242,N_4918,N_4677);
and U5243 (N_5243,N_4747,N_4975);
and U5244 (N_5244,N_4612,N_4812);
and U5245 (N_5245,N_4625,N_4853);
nand U5246 (N_5246,N_4992,N_4627);
nor U5247 (N_5247,N_4765,N_4771);
or U5248 (N_5248,N_4972,N_4695);
or U5249 (N_5249,N_4623,N_4570);
nand U5250 (N_5250,N_4788,N_4983);
or U5251 (N_5251,N_4987,N_4822);
nor U5252 (N_5252,N_4556,N_4819);
and U5253 (N_5253,N_4780,N_4572);
and U5254 (N_5254,N_4741,N_4925);
nand U5255 (N_5255,N_4682,N_4730);
and U5256 (N_5256,N_4533,N_4737);
nand U5257 (N_5257,N_4641,N_4807);
and U5258 (N_5258,N_4573,N_4926);
and U5259 (N_5259,N_4636,N_4939);
xor U5260 (N_5260,N_4728,N_4909);
xnor U5261 (N_5261,N_4562,N_4700);
nand U5262 (N_5262,N_4608,N_4805);
and U5263 (N_5263,N_4976,N_4783);
nand U5264 (N_5264,N_4681,N_4824);
and U5265 (N_5265,N_4631,N_4781);
xnor U5266 (N_5266,N_4791,N_4557);
or U5267 (N_5267,N_4509,N_4592);
nand U5268 (N_5268,N_4753,N_4717);
nor U5269 (N_5269,N_4985,N_4848);
or U5270 (N_5270,N_4682,N_4552);
and U5271 (N_5271,N_4854,N_4867);
or U5272 (N_5272,N_4584,N_4564);
nor U5273 (N_5273,N_4902,N_4688);
nand U5274 (N_5274,N_4678,N_4826);
nor U5275 (N_5275,N_4523,N_4846);
and U5276 (N_5276,N_4556,N_4713);
nor U5277 (N_5277,N_4966,N_4963);
xor U5278 (N_5278,N_4553,N_4611);
or U5279 (N_5279,N_4542,N_4932);
nor U5280 (N_5280,N_4864,N_4693);
or U5281 (N_5281,N_4681,N_4656);
or U5282 (N_5282,N_4754,N_4598);
or U5283 (N_5283,N_4571,N_4688);
nand U5284 (N_5284,N_4679,N_4728);
or U5285 (N_5285,N_4885,N_4944);
nor U5286 (N_5286,N_4797,N_4917);
nand U5287 (N_5287,N_4555,N_4620);
nand U5288 (N_5288,N_4651,N_4531);
nor U5289 (N_5289,N_4738,N_4503);
nand U5290 (N_5290,N_4859,N_4961);
nand U5291 (N_5291,N_4500,N_4534);
or U5292 (N_5292,N_4993,N_4613);
nand U5293 (N_5293,N_4934,N_4735);
nor U5294 (N_5294,N_4799,N_4557);
or U5295 (N_5295,N_4646,N_4661);
nor U5296 (N_5296,N_4568,N_4998);
nand U5297 (N_5297,N_4578,N_4883);
nor U5298 (N_5298,N_4755,N_4666);
nand U5299 (N_5299,N_4976,N_4583);
nand U5300 (N_5300,N_4664,N_4504);
nand U5301 (N_5301,N_4891,N_4783);
or U5302 (N_5302,N_4868,N_4776);
xor U5303 (N_5303,N_4991,N_4792);
or U5304 (N_5304,N_4753,N_4723);
nor U5305 (N_5305,N_4997,N_4643);
nand U5306 (N_5306,N_4721,N_4647);
or U5307 (N_5307,N_4645,N_4916);
or U5308 (N_5308,N_4935,N_4607);
nor U5309 (N_5309,N_4700,N_4836);
and U5310 (N_5310,N_4639,N_4665);
nor U5311 (N_5311,N_4790,N_4543);
nor U5312 (N_5312,N_4541,N_4873);
nand U5313 (N_5313,N_4799,N_4918);
nand U5314 (N_5314,N_4882,N_4586);
nand U5315 (N_5315,N_4522,N_4862);
or U5316 (N_5316,N_4749,N_4649);
and U5317 (N_5317,N_4869,N_4599);
nor U5318 (N_5318,N_4966,N_4833);
nand U5319 (N_5319,N_4827,N_4500);
nand U5320 (N_5320,N_4650,N_4663);
nor U5321 (N_5321,N_4883,N_4884);
and U5322 (N_5322,N_4893,N_4769);
and U5323 (N_5323,N_4543,N_4738);
nor U5324 (N_5324,N_4996,N_4514);
nand U5325 (N_5325,N_4825,N_4718);
nor U5326 (N_5326,N_4928,N_4628);
nor U5327 (N_5327,N_4958,N_4565);
or U5328 (N_5328,N_4904,N_4916);
or U5329 (N_5329,N_4822,N_4527);
nand U5330 (N_5330,N_4631,N_4979);
and U5331 (N_5331,N_4811,N_4732);
nand U5332 (N_5332,N_4716,N_4653);
nand U5333 (N_5333,N_4920,N_4687);
xor U5334 (N_5334,N_4775,N_4778);
nand U5335 (N_5335,N_4550,N_4860);
and U5336 (N_5336,N_4669,N_4500);
nand U5337 (N_5337,N_4545,N_4798);
xor U5338 (N_5338,N_4742,N_4565);
and U5339 (N_5339,N_4699,N_4836);
nor U5340 (N_5340,N_4503,N_4816);
nor U5341 (N_5341,N_4965,N_4508);
and U5342 (N_5342,N_4657,N_4844);
and U5343 (N_5343,N_4871,N_4743);
nand U5344 (N_5344,N_4818,N_4811);
or U5345 (N_5345,N_4541,N_4536);
nand U5346 (N_5346,N_4645,N_4504);
and U5347 (N_5347,N_4799,N_4741);
nand U5348 (N_5348,N_4637,N_4715);
xnor U5349 (N_5349,N_4746,N_4780);
nand U5350 (N_5350,N_4589,N_4757);
or U5351 (N_5351,N_4687,N_4976);
xnor U5352 (N_5352,N_4837,N_4876);
xnor U5353 (N_5353,N_4840,N_4509);
nor U5354 (N_5354,N_4914,N_4870);
or U5355 (N_5355,N_4866,N_4984);
nand U5356 (N_5356,N_4871,N_4947);
nor U5357 (N_5357,N_4576,N_4671);
or U5358 (N_5358,N_4535,N_4757);
nor U5359 (N_5359,N_4641,N_4653);
and U5360 (N_5360,N_4879,N_4701);
nor U5361 (N_5361,N_4882,N_4821);
xor U5362 (N_5362,N_4689,N_4636);
nand U5363 (N_5363,N_4931,N_4873);
nor U5364 (N_5364,N_4665,N_4764);
nor U5365 (N_5365,N_4526,N_4812);
and U5366 (N_5366,N_4623,N_4760);
or U5367 (N_5367,N_4911,N_4630);
or U5368 (N_5368,N_4968,N_4556);
nand U5369 (N_5369,N_4855,N_4540);
nand U5370 (N_5370,N_4763,N_4978);
and U5371 (N_5371,N_4910,N_4932);
and U5372 (N_5372,N_4998,N_4916);
or U5373 (N_5373,N_4721,N_4753);
or U5374 (N_5374,N_4976,N_4622);
nand U5375 (N_5375,N_4596,N_4796);
nand U5376 (N_5376,N_4932,N_4953);
or U5377 (N_5377,N_4910,N_4655);
nor U5378 (N_5378,N_4691,N_4628);
nor U5379 (N_5379,N_4678,N_4758);
and U5380 (N_5380,N_4822,N_4736);
nor U5381 (N_5381,N_4812,N_4631);
and U5382 (N_5382,N_4563,N_4996);
nand U5383 (N_5383,N_4905,N_4511);
and U5384 (N_5384,N_4590,N_4999);
nor U5385 (N_5385,N_4602,N_4949);
and U5386 (N_5386,N_4982,N_4553);
nor U5387 (N_5387,N_4677,N_4906);
and U5388 (N_5388,N_4531,N_4658);
and U5389 (N_5389,N_4962,N_4774);
nor U5390 (N_5390,N_4815,N_4587);
and U5391 (N_5391,N_4813,N_4589);
and U5392 (N_5392,N_4841,N_4791);
nor U5393 (N_5393,N_4962,N_4757);
and U5394 (N_5394,N_4649,N_4904);
or U5395 (N_5395,N_4700,N_4634);
xnor U5396 (N_5396,N_4542,N_4596);
nand U5397 (N_5397,N_4960,N_4831);
nor U5398 (N_5398,N_4974,N_4666);
nand U5399 (N_5399,N_4647,N_4909);
and U5400 (N_5400,N_4528,N_4895);
nor U5401 (N_5401,N_4943,N_4604);
and U5402 (N_5402,N_4587,N_4775);
nor U5403 (N_5403,N_4661,N_4819);
or U5404 (N_5404,N_4610,N_4578);
nand U5405 (N_5405,N_4620,N_4984);
and U5406 (N_5406,N_4792,N_4605);
and U5407 (N_5407,N_4987,N_4772);
or U5408 (N_5408,N_4661,N_4880);
nor U5409 (N_5409,N_4731,N_4742);
and U5410 (N_5410,N_4971,N_4656);
and U5411 (N_5411,N_4550,N_4738);
or U5412 (N_5412,N_4506,N_4586);
or U5413 (N_5413,N_4707,N_4649);
nor U5414 (N_5414,N_4733,N_4528);
nor U5415 (N_5415,N_4726,N_4916);
nand U5416 (N_5416,N_4754,N_4802);
or U5417 (N_5417,N_4810,N_4834);
or U5418 (N_5418,N_4692,N_4621);
or U5419 (N_5419,N_4636,N_4797);
nor U5420 (N_5420,N_4526,N_4689);
nand U5421 (N_5421,N_4584,N_4682);
nor U5422 (N_5422,N_4919,N_4649);
nor U5423 (N_5423,N_4890,N_4795);
xnor U5424 (N_5424,N_4581,N_4538);
or U5425 (N_5425,N_4896,N_4572);
or U5426 (N_5426,N_4612,N_4840);
nand U5427 (N_5427,N_4696,N_4553);
and U5428 (N_5428,N_4829,N_4524);
nand U5429 (N_5429,N_4941,N_4587);
nor U5430 (N_5430,N_4555,N_4522);
or U5431 (N_5431,N_4793,N_4767);
or U5432 (N_5432,N_4866,N_4724);
nor U5433 (N_5433,N_4945,N_4651);
xor U5434 (N_5434,N_4762,N_4989);
or U5435 (N_5435,N_4706,N_4581);
and U5436 (N_5436,N_4955,N_4884);
nand U5437 (N_5437,N_4674,N_4841);
or U5438 (N_5438,N_4883,N_4796);
xor U5439 (N_5439,N_4749,N_4977);
or U5440 (N_5440,N_4959,N_4575);
or U5441 (N_5441,N_4725,N_4724);
nor U5442 (N_5442,N_4936,N_4604);
nor U5443 (N_5443,N_4851,N_4675);
or U5444 (N_5444,N_4874,N_4692);
nand U5445 (N_5445,N_4633,N_4771);
or U5446 (N_5446,N_4677,N_4639);
nor U5447 (N_5447,N_4966,N_4746);
nand U5448 (N_5448,N_4875,N_4941);
or U5449 (N_5449,N_4752,N_4525);
nor U5450 (N_5450,N_4934,N_4943);
and U5451 (N_5451,N_4955,N_4579);
and U5452 (N_5452,N_4979,N_4541);
or U5453 (N_5453,N_4934,N_4634);
or U5454 (N_5454,N_4828,N_4531);
nand U5455 (N_5455,N_4521,N_4515);
or U5456 (N_5456,N_4919,N_4929);
and U5457 (N_5457,N_4918,N_4708);
and U5458 (N_5458,N_4828,N_4788);
nor U5459 (N_5459,N_4735,N_4730);
nor U5460 (N_5460,N_4906,N_4768);
nor U5461 (N_5461,N_4895,N_4882);
nand U5462 (N_5462,N_4823,N_4804);
and U5463 (N_5463,N_4806,N_4750);
and U5464 (N_5464,N_4728,N_4735);
nor U5465 (N_5465,N_4800,N_4750);
and U5466 (N_5466,N_4759,N_4693);
and U5467 (N_5467,N_4592,N_4873);
nand U5468 (N_5468,N_4750,N_4784);
nor U5469 (N_5469,N_4629,N_4580);
and U5470 (N_5470,N_4687,N_4794);
nand U5471 (N_5471,N_4894,N_4842);
xnor U5472 (N_5472,N_4552,N_4963);
or U5473 (N_5473,N_4634,N_4917);
and U5474 (N_5474,N_4896,N_4789);
nor U5475 (N_5475,N_4737,N_4729);
nand U5476 (N_5476,N_4991,N_4529);
and U5477 (N_5477,N_4904,N_4995);
or U5478 (N_5478,N_4705,N_4933);
nor U5479 (N_5479,N_4535,N_4740);
xnor U5480 (N_5480,N_4835,N_4585);
nand U5481 (N_5481,N_4547,N_4529);
nor U5482 (N_5482,N_4676,N_4870);
and U5483 (N_5483,N_4654,N_4811);
nor U5484 (N_5484,N_4955,N_4560);
nand U5485 (N_5485,N_4982,N_4924);
nand U5486 (N_5486,N_4809,N_4713);
nand U5487 (N_5487,N_4674,N_4814);
xnor U5488 (N_5488,N_4904,N_4712);
nor U5489 (N_5489,N_4606,N_4821);
nor U5490 (N_5490,N_4635,N_4985);
and U5491 (N_5491,N_4558,N_4500);
nand U5492 (N_5492,N_4515,N_4621);
nor U5493 (N_5493,N_4554,N_4796);
and U5494 (N_5494,N_4799,N_4697);
nor U5495 (N_5495,N_4511,N_4910);
nand U5496 (N_5496,N_4949,N_4631);
xnor U5497 (N_5497,N_4894,N_4930);
nand U5498 (N_5498,N_4807,N_4866);
nor U5499 (N_5499,N_4580,N_4854);
nand U5500 (N_5500,N_5386,N_5091);
xnor U5501 (N_5501,N_5052,N_5250);
and U5502 (N_5502,N_5181,N_5338);
or U5503 (N_5503,N_5140,N_5210);
nor U5504 (N_5504,N_5424,N_5170);
nor U5505 (N_5505,N_5272,N_5195);
nor U5506 (N_5506,N_5229,N_5293);
nor U5507 (N_5507,N_5261,N_5281);
xor U5508 (N_5508,N_5086,N_5473);
xnor U5509 (N_5509,N_5312,N_5233);
nand U5510 (N_5510,N_5037,N_5260);
xor U5511 (N_5511,N_5166,N_5454);
nand U5512 (N_5512,N_5378,N_5085);
and U5513 (N_5513,N_5374,N_5481);
or U5514 (N_5514,N_5194,N_5396);
and U5515 (N_5515,N_5249,N_5493);
nand U5516 (N_5516,N_5321,N_5299);
nor U5517 (N_5517,N_5452,N_5013);
and U5518 (N_5518,N_5259,N_5444);
or U5519 (N_5519,N_5044,N_5397);
nand U5520 (N_5520,N_5061,N_5377);
nand U5521 (N_5521,N_5235,N_5130);
and U5522 (N_5522,N_5209,N_5422);
nand U5523 (N_5523,N_5183,N_5006);
nor U5524 (N_5524,N_5110,N_5428);
xnor U5525 (N_5525,N_5141,N_5119);
or U5526 (N_5526,N_5198,N_5074);
nand U5527 (N_5527,N_5065,N_5277);
or U5528 (N_5528,N_5265,N_5201);
nor U5529 (N_5529,N_5484,N_5196);
or U5530 (N_5530,N_5108,N_5067);
or U5531 (N_5531,N_5418,N_5395);
or U5532 (N_5532,N_5350,N_5144);
and U5533 (N_5533,N_5020,N_5297);
and U5534 (N_5534,N_5150,N_5008);
xor U5535 (N_5535,N_5292,N_5326);
or U5536 (N_5536,N_5342,N_5003);
nor U5537 (N_5537,N_5335,N_5327);
or U5538 (N_5538,N_5398,N_5063);
nand U5539 (N_5539,N_5294,N_5227);
nor U5540 (N_5540,N_5171,N_5262);
nand U5541 (N_5541,N_5266,N_5200);
and U5542 (N_5542,N_5096,N_5245);
nand U5543 (N_5543,N_5392,N_5351);
and U5544 (N_5544,N_5113,N_5393);
xnor U5545 (N_5545,N_5451,N_5178);
nor U5546 (N_5546,N_5177,N_5291);
or U5547 (N_5547,N_5216,N_5236);
or U5548 (N_5548,N_5483,N_5426);
xor U5549 (N_5549,N_5363,N_5440);
or U5550 (N_5550,N_5267,N_5298);
or U5551 (N_5551,N_5151,N_5439);
or U5552 (N_5552,N_5107,N_5322);
nand U5553 (N_5553,N_5316,N_5295);
nand U5554 (N_5554,N_5358,N_5115);
or U5555 (N_5555,N_5190,N_5314);
nand U5556 (N_5556,N_5476,N_5399);
or U5557 (N_5557,N_5370,N_5328);
or U5558 (N_5558,N_5159,N_5051);
and U5559 (N_5559,N_5186,N_5224);
nor U5560 (N_5560,N_5076,N_5441);
nand U5561 (N_5561,N_5045,N_5274);
nand U5562 (N_5562,N_5134,N_5279);
and U5563 (N_5563,N_5301,N_5050);
or U5564 (N_5564,N_5005,N_5375);
and U5565 (N_5565,N_5032,N_5368);
and U5566 (N_5566,N_5099,N_5208);
or U5567 (N_5567,N_5055,N_5286);
and U5568 (N_5568,N_5491,N_5197);
xor U5569 (N_5569,N_5203,N_5359);
and U5570 (N_5570,N_5352,N_5495);
and U5571 (N_5571,N_5461,N_5019);
or U5572 (N_5572,N_5089,N_5361);
nand U5573 (N_5573,N_5340,N_5106);
and U5574 (N_5574,N_5367,N_5284);
and U5575 (N_5575,N_5163,N_5355);
or U5576 (N_5576,N_5143,N_5101);
or U5577 (N_5577,N_5460,N_5215);
xor U5578 (N_5578,N_5356,N_5102);
nand U5579 (N_5579,N_5191,N_5271);
nor U5580 (N_5580,N_5320,N_5456);
or U5581 (N_5581,N_5409,N_5357);
or U5582 (N_5582,N_5160,N_5057);
or U5583 (N_5583,N_5010,N_5218);
nand U5584 (N_5584,N_5238,N_5157);
nor U5585 (N_5585,N_5283,N_5349);
or U5586 (N_5586,N_5111,N_5251);
xor U5587 (N_5587,N_5420,N_5416);
xor U5588 (N_5588,N_5325,N_5148);
nor U5589 (N_5589,N_5225,N_5379);
and U5590 (N_5590,N_5289,N_5034);
or U5591 (N_5591,N_5394,N_5239);
xor U5592 (N_5592,N_5211,N_5025);
or U5593 (N_5593,N_5212,N_5470);
or U5594 (N_5594,N_5318,N_5332);
nor U5595 (N_5595,N_5475,N_5145);
nand U5596 (N_5596,N_5221,N_5288);
xnor U5597 (N_5597,N_5242,N_5385);
or U5598 (N_5598,N_5185,N_5078);
or U5599 (N_5599,N_5348,N_5339);
nor U5600 (N_5600,N_5463,N_5139);
and U5601 (N_5601,N_5009,N_5453);
nor U5602 (N_5602,N_5285,N_5254);
and U5603 (N_5603,N_5469,N_5124);
nor U5604 (N_5604,N_5169,N_5131);
nand U5605 (N_5605,N_5176,N_5064);
or U5606 (N_5606,N_5429,N_5031);
nand U5607 (N_5607,N_5499,N_5164);
nor U5608 (N_5608,N_5097,N_5287);
or U5609 (N_5609,N_5087,N_5280);
nand U5610 (N_5610,N_5012,N_5402);
and U5611 (N_5611,N_5069,N_5419);
xor U5612 (N_5612,N_5366,N_5468);
nor U5613 (N_5613,N_5466,N_5184);
nor U5614 (N_5614,N_5388,N_5095);
nor U5615 (N_5615,N_5205,N_5432);
or U5616 (N_5616,N_5474,N_5443);
and U5617 (N_5617,N_5334,N_5431);
xor U5618 (N_5618,N_5172,N_5448);
nand U5619 (N_5619,N_5090,N_5118);
and U5620 (N_5620,N_5192,N_5122);
nor U5621 (N_5621,N_5120,N_5018);
and U5622 (N_5622,N_5437,N_5058);
and U5623 (N_5623,N_5354,N_5180);
nor U5624 (N_5624,N_5498,N_5492);
nor U5625 (N_5625,N_5268,N_5077);
xor U5626 (N_5626,N_5270,N_5080);
nor U5627 (N_5627,N_5083,N_5415);
or U5628 (N_5628,N_5305,N_5438);
xor U5629 (N_5629,N_5389,N_5129);
and U5630 (N_5630,N_5026,N_5365);
nand U5631 (N_5631,N_5188,N_5158);
and U5632 (N_5632,N_5071,N_5347);
or U5633 (N_5633,N_5373,N_5059);
nor U5634 (N_5634,N_5165,N_5048);
nand U5635 (N_5635,N_5155,N_5489);
xnor U5636 (N_5636,N_5278,N_5362);
nand U5637 (N_5637,N_5060,N_5193);
or U5638 (N_5638,N_5391,N_5496);
nor U5639 (N_5639,N_5036,N_5258);
and U5640 (N_5640,N_5217,N_5040);
and U5641 (N_5641,N_5088,N_5412);
nor U5642 (N_5642,N_5346,N_5023);
or U5643 (N_5643,N_5345,N_5230);
or U5644 (N_5644,N_5387,N_5041);
or U5645 (N_5645,N_5081,N_5407);
and U5646 (N_5646,N_5455,N_5070);
or U5647 (N_5647,N_5282,N_5445);
xor U5648 (N_5648,N_5408,N_5263);
xor U5649 (N_5649,N_5175,N_5179);
and U5650 (N_5650,N_5100,N_5447);
xnor U5651 (N_5651,N_5331,N_5317);
and U5652 (N_5652,N_5147,N_5497);
nor U5653 (N_5653,N_5376,N_5187);
or U5654 (N_5654,N_5001,N_5042);
and U5655 (N_5655,N_5024,N_5433);
nor U5656 (N_5656,N_5204,N_5306);
nor U5657 (N_5657,N_5309,N_5182);
nor U5658 (N_5658,N_5202,N_5066);
and U5659 (N_5659,N_5311,N_5307);
or U5660 (N_5660,N_5223,N_5458);
and U5661 (N_5661,N_5465,N_5459);
xor U5662 (N_5662,N_5324,N_5146);
nand U5663 (N_5663,N_5341,N_5411);
nand U5664 (N_5664,N_5062,N_5472);
or U5665 (N_5665,N_5199,N_5093);
or U5666 (N_5666,N_5275,N_5132);
and U5667 (N_5667,N_5168,N_5053);
nor U5668 (N_5668,N_5343,N_5296);
nand U5669 (N_5669,N_5220,N_5329);
or U5670 (N_5670,N_5017,N_5478);
or U5671 (N_5671,N_5256,N_5353);
xor U5672 (N_5672,N_5380,N_5104);
and U5673 (N_5673,N_5021,N_5109);
nor U5674 (N_5674,N_5330,N_5384);
or U5675 (N_5675,N_5126,N_5068);
or U5676 (N_5676,N_5310,N_5153);
xor U5677 (N_5677,N_5257,N_5035);
nand U5678 (N_5678,N_5382,N_5105);
nand U5679 (N_5679,N_5406,N_5092);
or U5680 (N_5680,N_5033,N_5425);
nand U5681 (N_5681,N_5156,N_5390);
nor U5682 (N_5682,N_5127,N_5490);
nor U5683 (N_5683,N_5243,N_5253);
nor U5684 (N_5684,N_5421,N_5303);
nor U5685 (N_5685,N_5450,N_5047);
and U5686 (N_5686,N_5434,N_5414);
nand U5687 (N_5687,N_5308,N_5073);
nand U5688 (N_5688,N_5417,N_5174);
nor U5689 (N_5689,N_5477,N_5479);
or U5690 (N_5690,N_5046,N_5167);
nor U5691 (N_5691,N_5136,N_5049);
or U5692 (N_5692,N_5007,N_5462);
and U5693 (N_5693,N_5123,N_5371);
and U5694 (N_5694,N_5084,N_5116);
nor U5695 (N_5695,N_5121,N_5161);
nor U5696 (N_5696,N_5319,N_5446);
and U5697 (N_5697,N_5304,N_5098);
nor U5698 (N_5698,N_5467,N_5043);
or U5699 (N_5699,N_5149,N_5276);
nand U5700 (N_5700,N_5404,N_5457);
nand U5701 (N_5701,N_5228,N_5360);
nand U5702 (N_5702,N_5222,N_5079);
nand U5703 (N_5703,N_5400,N_5056);
and U5704 (N_5704,N_5436,N_5381);
nor U5705 (N_5705,N_5264,N_5369);
or U5706 (N_5706,N_5494,N_5435);
and U5707 (N_5707,N_5094,N_5219);
nor U5708 (N_5708,N_5449,N_5207);
or U5709 (N_5709,N_5240,N_5486);
or U5710 (N_5710,N_5162,N_5372);
or U5711 (N_5711,N_5244,N_5030);
and U5712 (N_5712,N_5237,N_5154);
nand U5713 (N_5713,N_5290,N_5427);
or U5714 (N_5714,N_5252,N_5214);
or U5715 (N_5715,N_5248,N_5075);
or U5716 (N_5716,N_5336,N_5430);
xnor U5717 (N_5717,N_5114,N_5082);
or U5718 (N_5718,N_5269,N_5054);
or U5719 (N_5719,N_5004,N_5273);
or U5720 (N_5720,N_5442,N_5300);
and U5721 (N_5721,N_5234,N_5038);
nor U5722 (N_5722,N_5028,N_5344);
and U5723 (N_5723,N_5471,N_5482);
nor U5724 (N_5724,N_5117,N_5173);
and U5725 (N_5725,N_5480,N_5206);
and U5726 (N_5726,N_5133,N_5383);
or U5727 (N_5727,N_5405,N_5423);
nand U5728 (N_5728,N_5112,N_5302);
nand U5729 (N_5729,N_5337,N_5000);
nand U5730 (N_5730,N_5464,N_5128);
and U5731 (N_5731,N_5015,N_5135);
and U5732 (N_5732,N_5039,N_5485);
or U5733 (N_5733,N_5488,N_5138);
nor U5734 (N_5734,N_5247,N_5027);
or U5735 (N_5735,N_5315,N_5011);
or U5736 (N_5736,N_5226,N_5014);
and U5737 (N_5737,N_5029,N_5323);
or U5738 (N_5738,N_5255,N_5016);
or U5739 (N_5739,N_5189,N_5333);
nor U5740 (N_5740,N_5241,N_5142);
and U5741 (N_5741,N_5002,N_5231);
and U5742 (N_5742,N_5232,N_5313);
and U5743 (N_5743,N_5413,N_5403);
nand U5744 (N_5744,N_5213,N_5364);
and U5745 (N_5745,N_5022,N_5152);
or U5746 (N_5746,N_5246,N_5103);
nand U5747 (N_5747,N_5401,N_5410);
or U5748 (N_5748,N_5125,N_5137);
nor U5749 (N_5749,N_5487,N_5072);
nand U5750 (N_5750,N_5015,N_5442);
or U5751 (N_5751,N_5303,N_5300);
nor U5752 (N_5752,N_5420,N_5352);
and U5753 (N_5753,N_5254,N_5400);
nand U5754 (N_5754,N_5392,N_5364);
nor U5755 (N_5755,N_5144,N_5300);
and U5756 (N_5756,N_5484,N_5008);
and U5757 (N_5757,N_5011,N_5037);
nand U5758 (N_5758,N_5193,N_5407);
nor U5759 (N_5759,N_5326,N_5196);
nor U5760 (N_5760,N_5196,N_5159);
or U5761 (N_5761,N_5142,N_5130);
and U5762 (N_5762,N_5455,N_5005);
nand U5763 (N_5763,N_5391,N_5381);
or U5764 (N_5764,N_5148,N_5270);
nand U5765 (N_5765,N_5348,N_5443);
nand U5766 (N_5766,N_5071,N_5210);
nand U5767 (N_5767,N_5477,N_5208);
nand U5768 (N_5768,N_5344,N_5416);
nor U5769 (N_5769,N_5418,N_5489);
or U5770 (N_5770,N_5134,N_5319);
xnor U5771 (N_5771,N_5165,N_5433);
or U5772 (N_5772,N_5074,N_5291);
or U5773 (N_5773,N_5268,N_5248);
and U5774 (N_5774,N_5399,N_5204);
and U5775 (N_5775,N_5066,N_5088);
or U5776 (N_5776,N_5210,N_5149);
xor U5777 (N_5777,N_5293,N_5483);
nor U5778 (N_5778,N_5112,N_5460);
nand U5779 (N_5779,N_5250,N_5152);
nor U5780 (N_5780,N_5331,N_5460);
or U5781 (N_5781,N_5339,N_5472);
xor U5782 (N_5782,N_5132,N_5371);
or U5783 (N_5783,N_5405,N_5252);
or U5784 (N_5784,N_5385,N_5164);
and U5785 (N_5785,N_5353,N_5342);
nor U5786 (N_5786,N_5179,N_5212);
nand U5787 (N_5787,N_5284,N_5237);
and U5788 (N_5788,N_5371,N_5296);
nor U5789 (N_5789,N_5419,N_5346);
nand U5790 (N_5790,N_5151,N_5391);
nor U5791 (N_5791,N_5013,N_5363);
and U5792 (N_5792,N_5046,N_5466);
and U5793 (N_5793,N_5368,N_5437);
or U5794 (N_5794,N_5247,N_5376);
and U5795 (N_5795,N_5225,N_5124);
and U5796 (N_5796,N_5497,N_5452);
nand U5797 (N_5797,N_5427,N_5309);
and U5798 (N_5798,N_5230,N_5472);
and U5799 (N_5799,N_5405,N_5469);
xor U5800 (N_5800,N_5154,N_5049);
and U5801 (N_5801,N_5355,N_5111);
and U5802 (N_5802,N_5182,N_5327);
and U5803 (N_5803,N_5046,N_5384);
nor U5804 (N_5804,N_5050,N_5128);
or U5805 (N_5805,N_5337,N_5241);
nor U5806 (N_5806,N_5002,N_5101);
and U5807 (N_5807,N_5445,N_5133);
nor U5808 (N_5808,N_5261,N_5493);
xor U5809 (N_5809,N_5482,N_5402);
or U5810 (N_5810,N_5339,N_5326);
nor U5811 (N_5811,N_5236,N_5040);
xor U5812 (N_5812,N_5477,N_5035);
nand U5813 (N_5813,N_5090,N_5007);
nor U5814 (N_5814,N_5247,N_5379);
or U5815 (N_5815,N_5480,N_5087);
nand U5816 (N_5816,N_5029,N_5053);
or U5817 (N_5817,N_5361,N_5418);
or U5818 (N_5818,N_5167,N_5271);
or U5819 (N_5819,N_5495,N_5368);
or U5820 (N_5820,N_5282,N_5456);
nor U5821 (N_5821,N_5133,N_5341);
and U5822 (N_5822,N_5243,N_5481);
or U5823 (N_5823,N_5262,N_5294);
nor U5824 (N_5824,N_5086,N_5060);
nand U5825 (N_5825,N_5288,N_5038);
nor U5826 (N_5826,N_5049,N_5272);
nor U5827 (N_5827,N_5278,N_5406);
and U5828 (N_5828,N_5095,N_5401);
nand U5829 (N_5829,N_5235,N_5258);
and U5830 (N_5830,N_5241,N_5125);
nand U5831 (N_5831,N_5391,N_5370);
nand U5832 (N_5832,N_5404,N_5015);
and U5833 (N_5833,N_5231,N_5339);
or U5834 (N_5834,N_5168,N_5255);
and U5835 (N_5835,N_5482,N_5411);
nand U5836 (N_5836,N_5301,N_5354);
nand U5837 (N_5837,N_5463,N_5331);
nand U5838 (N_5838,N_5060,N_5295);
nor U5839 (N_5839,N_5143,N_5026);
nor U5840 (N_5840,N_5075,N_5033);
nand U5841 (N_5841,N_5066,N_5080);
nor U5842 (N_5842,N_5447,N_5354);
nor U5843 (N_5843,N_5411,N_5199);
and U5844 (N_5844,N_5313,N_5155);
xor U5845 (N_5845,N_5369,N_5293);
or U5846 (N_5846,N_5455,N_5148);
nand U5847 (N_5847,N_5133,N_5173);
nand U5848 (N_5848,N_5237,N_5099);
and U5849 (N_5849,N_5026,N_5370);
nand U5850 (N_5850,N_5075,N_5080);
or U5851 (N_5851,N_5466,N_5150);
nor U5852 (N_5852,N_5096,N_5071);
or U5853 (N_5853,N_5460,N_5220);
or U5854 (N_5854,N_5128,N_5070);
nand U5855 (N_5855,N_5468,N_5333);
nand U5856 (N_5856,N_5071,N_5167);
nor U5857 (N_5857,N_5065,N_5295);
nand U5858 (N_5858,N_5382,N_5122);
nand U5859 (N_5859,N_5311,N_5213);
and U5860 (N_5860,N_5308,N_5469);
nand U5861 (N_5861,N_5384,N_5113);
nand U5862 (N_5862,N_5093,N_5423);
and U5863 (N_5863,N_5092,N_5036);
nor U5864 (N_5864,N_5480,N_5132);
nand U5865 (N_5865,N_5381,N_5348);
nor U5866 (N_5866,N_5281,N_5185);
or U5867 (N_5867,N_5048,N_5144);
or U5868 (N_5868,N_5037,N_5166);
or U5869 (N_5869,N_5205,N_5353);
xor U5870 (N_5870,N_5385,N_5153);
nor U5871 (N_5871,N_5287,N_5383);
or U5872 (N_5872,N_5354,N_5489);
and U5873 (N_5873,N_5465,N_5270);
and U5874 (N_5874,N_5198,N_5369);
nor U5875 (N_5875,N_5000,N_5186);
and U5876 (N_5876,N_5413,N_5261);
and U5877 (N_5877,N_5402,N_5445);
nor U5878 (N_5878,N_5474,N_5065);
nand U5879 (N_5879,N_5425,N_5305);
nor U5880 (N_5880,N_5271,N_5325);
nor U5881 (N_5881,N_5245,N_5041);
and U5882 (N_5882,N_5377,N_5002);
xor U5883 (N_5883,N_5317,N_5461);
xor U5884 (N_5884,N_5342,N_5116);
or U5885 (N_5885,N_5344,N_5056);
or U5886 (N_5886,N_5106,N_5235);
xnor U5887 (N_5887,N_5032,N_5080);
or U5888 (N_5888,N_5064,N_5294);
nand U5889 (N_5889,N_5323,N_5472);
and U5890 (N_5890,N_5263,N_5317);
or U5891 (N_5891,N_5084,N_5317);
or U5892 (N_5892,N_5210,N_5284);
nand U5893 (N_5893,N_5230,N_5174);
nand U5894 (N_5894,N_5072,N_5094);
or U5895 (N_5895,N_5175,N_5244);
and U5896 (N_5896,N_5132,N_5248);
or U5897 (N_5897,N_5296,N_5482);
nor U5898 (N_5898,N_5391,N_5404);
nand U5899 (N_5899,N_5343,N_5426);
or U5900 (N_5900,N_5308,N_5315);
and U5901 (N_5901,N_5353,N_5257);
nor U5902 (N_5902,N_5342,N_5489);
nor U5903 (N_5903,N_5421,N_5110);
or U5904 (N_5904,N_5268,N_5468);
nor U5905 (N_5905,N_5419,N_5333);
and U5906 (N_5906,N_5400,N_5353);
xnor U5907 (N_5907,N_5127,N_5393);
or U5908 (N_5908,N_5429,N_5455);
nand U5909 (N_5909,N_5074,N_5459);
or U5910 (N_5910,N_5206,N_5263);
nor U5911 (N_5911,N_5099,N_5140);
nand U5912 (N_5912,N_5453,N_5040);
nand U5913 (N_5913,N_5224,N_5446);
nand U5914 (N_5914,N_5061,N_5188);
nor U5915 (N_5915,N_5369,N_5494);
and U5916 (N_5916,N_5308,N_5355);
xor U5917 (N_5917,N_5179,N_5220);
and U5918 (N_5918,N_5235,N_5351);
nor U5919 (N_5919,N_5072,N_5062);
nand U5920 (N_5920,N_5177,N_5489);
and U5921 (N_5921,N_5262,N_5373);
and U5922 (N_5922,N_5093,N_5201);
or U5923 (N_5923,N_5062,N_5361);
and U5924 (N_5924,N_5360,N_5129);
or U5925 (N_5925,N_5283,N_5389);
or U5926 (N_5926,N_5158,N_5266);
and U5927 (N_5927,N_5294,N_5303);
and U5928 (N_5928,N_5487,N_5377);
or U5929 (N_5929,N_5165,N_5141);
or U5930 (N_5930,N_5000,N_5373);
and U5931 (N_5931,N_5208,N_5060);
xor U5932 (N_5932,N_5299,N_5298);
or U5933 (N_5933,N_5476,N_5030);
nand U5934 (N_5934,N_5409,N_5052);
nor U5935 (N_5935,N_5254,N_5472);
nor U5936 (N_5936,N_5416,N_5089);
nand U5937 (N_5937,N_5446,N_5399);
nand U5938 (N_5938,N_5224,N_5088);
nand U5939 (N_5939,N_5327,N_5427);
or U5940 (N_5940,N_5256,N_5407);
nor U5941 (N_5941,N_5438,N_5333);
nor U5942 (N_5942,N_5222,N_5228);
or U5943 (N_5943,N_5160,N_5341);
and U5944 (N_5944,N_5496,N_5041);
or U5945 (N_5945,N_5367,N_5262);
or U5946 (N_5946,N_5290,N_5443);
nand U5947 (N_5947,N_5363,N_5034);
nor U5948 (N_5948,N_5098,N_5458);
nand U5949 (N_5949,N_5024,N_5030);
nor U5950 (N_5950,N_5109,N_5094);
and U5951 (N_5951,N_5410,N_5304);
xor U5952 (N_5952,N_5100,N_5164);
nor U5953 (N_5953,N_5175,N_5328);
or U5954 (N_5954,N_5446,N_5429);
nand U5955 (N_5955,N_5011,N_5433);
xnor U5956 (N_5956,N_5196,N_5402);
nand U5957 (N_5957,N_5041,N_5204);
nor U5958 (N_5958,N_5158,N_5467);
xor U5959 (N_5959,N_5105,N_5122);
or U5960 (N_5960,N_5383,N_5027);
or U5961 (N_5961,N_5471,N_5473);
or U5962 (N_5962,N_5026,N_5302);
nor U5963 (N_5963,N_5457,N_5165);
nor U5964 (N_5964,N_5160,N_5108);
or U5965 (N_5965,N_5248,N_5023);
or U5966 (N_5966,N_5400,N_5445);
or U5967 (N_5967,N_5240,N_5393);
nand U5968 (N_5968,N_5281,N_5362);
or U5969 (N_5969,N_5309,N_5411);
xor U5970 (N_5970,N_5165,N_5495);
or U5971 (N_5971,N_5145,N_5414);
xor U5972 (N_5972,N_5161,N_5314);
nor U5973 (N_5973,N_5269,N_5379);
and U5974 (N_5974,N_5060,N_5228);
nand U5975 (N_5975,N_5010,N_5421);
and U5976 (N_5976,N_5197,N_5105);
nand U5977 (N_5977,N_5207,N_5456);
nand U5978 (N_5978,N_5141,N_5413);
nand U5979 (N_5979,N_5202,N_5087);
nor U5980 (N_5980,N_5316,N_5355);
nor U5981 (N_5981,N_5220,N_5199);
or U5982 (N_5982,N_5154,N_5404);
xor U5983 (N_5983,N_5208,N_5389);
and U5984 (N_5984,N_5048,N_5207);
nand U5985 (N_5985,N_5077,N_5224);
or U5986 (N_5986,N_5277,N_5032);
and U5987 (N_5987,N_5364,N_5388);
nand U5988 (N_5988,N_5106,N_5094);
xnor U5989 (N_5989,N_5025,N_5442);
nor U5990 (N_5990,N_5294,N_5174);
nand U5991 (N_5991,N_5024,N_5065);
nand U5992 (N_5992,N_5271,N_5051);
or U5993 (N_5993,N_5492,N_5434);
or U5994 (N_5994,N_5138,N_5484);
and U5995 (N_5995,N_5317,N_5479);
and U5996 (N_5996,N_5102,N_5001);
or U5997 (N_5997,N_5409,N_5189);
or U5998 (N_5998,N_5259,N_5343);
nor U5999 (N_5999,N_5486,N_5339);
and U6000 (N_6000,N_5679,N_5754);
and U6001 (N_6001,N_5635,N_5989);
nor U6002 (N_6002,N_5582,N_5820);
and U6003 (N_6003,N_5707,N_5940);
or U6004 (N_6004,N_5523,N_5658);
nor U6005 (N_6005,N_5792,N_5917);
nand U6006 (N_6006,N_5554,N_5779);
nor U6007 (N_6007,N_5963,N_5950);
xnor U6008 (N_6008,N_5734,N_5633);
and U6009 (N_6009,N_5529,N_5642);
and U6010 (N_6010,N_5544,N_5728);
nor U6011 (N_6011,N_5730,N_5619);
or U6012 (N_6012,N_5918,N_5849);
nand U6013 (N_6013,N_5915,N_5938);
nor U6014 (N_6014,N_5667,N_5946);
nand U6015 (N_6015,N_5861,N_5684);
nor U6016 (N_6016,N_5815,N_5751);
xnor U6017 (N_6017,N_5511,N_5678);
or U6018 (N_6018,N_5549,N_5829);
and U6019 (N_6019,N_5683,N_5741);
and U6020 (N_6020,N_5670,N_5931);
and U6021 (N_6021,N_5532,N_5524);
or U6022 (N_6022,N_5685,N_5726);
nand U6023 (N_6023,N_5793,N_5551);
nor U6024 (N_6024,N_5783,N_5747);
nor U6025 (N_6025,N_5876,N_5765);
and U6026 (N_6026,N_5797,N_5778);
and U6027 (N_6027,N_5837,N_5513);
nor U6028 (N_6028,N_5835,N_5641);
and U6029 (N_6029,N_5791,N_5817);
nand U6030 (N_6030,N_5941,N_5688);
and U6031 (N_6031,N_5697,N_5569);
nor U6032 (N_6032,N_5844,N_5882);
nand U6033 (N_6033,N_5603,N_5901);
or U6034 (N_6034,N_5905,N_5805);
xor U6035 (N_6035,N_5720,N_5789);
and U6036 (N_6036,N_5894,N_5659);
nand U6037 (N_6037,N_5690,N_5586);
and U6038 (N_6038,N_5864,N_5848);
nor U6039 (N_6039,N_5801,N_5859);
and U6040 (N_6040,N_5889,N_5957);
xor U6041 (N_6041,N_5903,N_5780);
or U6042 (N_6042,N_5863,N_5997);
and U6043 (N_6043,N_5893,N_5571);
nor U6044 (N_6044,N_5545,N_5872);
or U6045 (N_6045,N_5528,N_5722);
nand U6046 (N_6046,N_5890,N_5570);
and U6047 (N_6047,N_5561,N_5929);
nand U6048 (N_6048,N_5629,N_5852);
nor U6049 (N_6049,N_5883,N_5886);
or U6050 (N_6050,N_5921,N_5577);
and U6051 (N_6051,N_5972,N_5847);
xor U6052 (N_6052,N_5724,N_5613);
and U6053 (N_6053,N_5896,N_5624);
nand U6054 (N_6054,N_5669,N_5907);
xnor U6055 (N_6055,N_5846,N_5628);
nor U6056 (N_6056,N_5512,N_5742);
or U6057 (N_6057,N_5969,N_5655);
and U6058 (N_6058,N_5509,N_5737);
and U6059 (N_6059,N_5949,N_5622);
nor U6060 (N_6060,N_5911,N_5714);
nor U6061 (N_6061,N_5795,N_5839);
or U6062 (N_6062,N_5873,N_5943);
or U6063 (N_6063,N_5596,N_5716);
and U6064 (N_6064,N_5869,N_5536);
and U6065 (N_6065,N_5930,N_5701);
xnor U6066 (N_6066,N_5919,N_5588);
and U6067 (N_6067,N_5717,N_5825);
or U6068 (N_6068,N_5530,N_5761);
and U6069 (N_6069,N_5925,N_5804);
nand U6070 (N_6070,N_5712,N_5970);
or U6071 (N_6071,N_5926,N_5992);
nor U6072 (N_6072,N_5581,N_5660);
or U6073 (N_6073,N_5753,N_5502);
nor U6074 (N_6074,N_5508,N_5552);
and U6075 (N_6075,N_5991,N_5763);
nor U6076 (N_6076,N_5774,N_5843);
or U6077 (N_6077,N_5672,N_5968);
or U6078 (N_6078,N_5606,N_5636);
or U6079 (N_6079,N_5700,N_5776);
and U6080 (N_6080,N_5738,N_5773);
and U6081 (N_6081,N_5522,N_5695);
or U6082 (N_6082,N_5637,N_5934);
nand U6083 (N_6083,N_5782,N_5704);
nand U6084 (N_6084,N_5671,N_5924);
and U6085 (N_6085,N_5975,N_5654);
or U6086 (N_6086,N_5981,N_5923);
or U6087 (N_6087,N_5652,N_5759);
or U6088 (N_6088,N_5798,N_5572);
nand U6089 (N_6089,N_5750,N_5994);
or U6090 (N_6090,N_5945,N_5956);
xor U6091 (N_6091,N_5696,N_5814);
and U6092 (N_6092,N_5687,N_5944);
nand U6093 (N_6093,N_5760,N_5609);
nor U6094 (N_6094,N_5764,N_5996);
and U6095 (N_6095,N_5521,N_5816);
nor U6096 (N_6096,N_5645,N_5651);
and U6097 (N_6097,N_5807,N_5884);
or U6098 (N_6098,N_5600,N_5977);
and U6099 (N_6099,N_5546,N_5743);
nand U6100 (N_6100,N_5813,N_5576);
nand U6101 (N_6101,N_5518,N_5736);
nor U6102 (N_6102,N_5574,N_5653);
nand U6103 (N_6103,N_5727,N_5733);
or U6104 (N_6104,N_5965,N_5984);
or U6105 (N_6105,N_5526,N_5608);
or U6106 (N_6106,N_5649,N_5888);
nand U6107 (N_6107,N_5547,N_5838);
nand U6108 (N_6108,N_5604,N_5752);
nor U6109 (N_6109,N_5675,N_5575);
xnor U6110 (N_6110,N_5689,N_5506);
nand U6111 (N_6111,N_5897,N_5555);
and U6112 (N_6112,N_5702,N_5706);
nor U6113 (N_6113,N_5762,N_5694);
nor U6114 (N_6114,N_5673,N_5531);
nand U6115 (N_6115,N_5657,N_5812);
xnor U6116 (N_6116,N_5713,N_5592);
nor U6117 (N_6117,N_5982,N_5976);
or U6118 (N_6118,N_5955,N_5709);
nand U6119 (N_6119,N_5845,N_5858);
nor U6120 (N_6120,N_5824,N_5735);
nor U6121 (N_6121,N_5605,N_5537);
and U6122 (N_6122,N_5539,N_5595);
and U6123 (N_6123,N_5857,N_5935);
nand U6124 (N_6124,N_5880,N_5680);
or U6125 (N_6125,N_5729,N_5620);
or U6126 (N_6126,N_5607,N_5514);
or U6127 (N_6127,N_5556,N_5597);
or U6128 (N_6128,N_5818,N_5718);
and U6129 (N_6129,N_5585,N_5803);
nand U6130 (N_6130,N_5909,N_5987);
nand U6131 (N_6131,N_5922,N_5723);
nor U6132 (N_6132,N_5842,N_5860);
or U6133 (N_6133,N_5995,N_5507);
or U6134 (N_6134,N_5986,N_5715);
and U6135 (N_6135,N_5579,N_5627);
and U6136 (N_6136,N_5906,N_5661);
or U6137 (N_6137,N_5692,N_5932);
and U6138 (N_6138,N_5510,N_5802);
or U6139 (N_6139,N_5746,N_5564);
and U6140 (N_6140,N_5821,N_5646);
nand U6141 (N_6141,N_5594,N_5520);
nand U6142 (N_6142,N_5881,N_5568);
xnor U6143 (N_6143,N_5519,N_5623);
or U6144 (N_6144,N_5978,N_5503);
nor U6145 (N_6145,N_5535,N_5598);
and U6146 (N_6146,N_5904,N_5560);
or U6147 (N_6147,N_5999,N_5826);
nand U6148 (N_6148,N_5691,N_5617);
nor U6149 (N_6149,N_5983,N_5703);
nor U6150 (N_6150,N_5553,N_5565);
nor U6151 (N_6151,N_5912,N_5515);
or U6152 (N_6152,N_5583,N_5854);
and U6153 (N_6153,N_5501,N_5808);
nand U6154 (N_6154,N_5841,N_5740);
and U6155 (N_6155,N_5614,N_5666);
nand U6156 (N_6156,N_5942,N_5832);
and U6157 (N_6157,N_5631,N_5708);
nor U6158 (N_6158,N_5947,N_5809);
nor U6159 (N_6159,N_5504,N_5563);
and U6160 (N_6160,N_5767,N_5558);
and U6161 (N_6161,N_5542,N_5557);
and U6162 (N_6162,N_5664,N_5867);
or U6163 (N_6163,N_5732,N_5757);
or U6164 (N_6164,N_5541,N_5961);
nor U6165 (N_6165,N_5533,N_5819);
nor U6166 (N_6166,N_5634,N_5908);
xor U6167 (N_6167,N_5662,N_5775);
and U6168 (N_6168,N_5853,N_5862);
nand U6169 (N_6169,N_5621,N_5632);
nand U6170 (N_6170,N_5980,N_5875);
or U6171 (N_6171,N_5611,N_5806);
nand U6172 (N_6172,N_5916,N_5898);
nand U6173 (N_6173,N_5505,N_5612);
and U6174 (N_6174,N_5618,N_5705);
nand U6175 (N_6175,N_5674,N_5711);
and U6176 (N_6176,N_5587,N_5885);
nor U6177 (N_6177,N_5971,N_5985);
xor U6178 (N_6178,N_5840,N_5870);
and U6179 (N_6179,N_5874,N_5851);
or U6180 (N_6180,N_5786,N_5681);
nor U6181 (N_6181,N_5777,N_5788);
or U6182 (N_6182,N_5668,N_5865);
and U6183 (N_6183,N_5640,N_5974);
nand U6184 (N_6184,N_5534,N_5966);
nor U6185 (N_6185,N_5573,N_5951);
and U6186 (N_6186,N_5698,N_5787);
and U6187 (N_6187,N_5913,N_5630);
or U6188 (N_6188,N_5610,N_5756);
or U6189 (N_6189,N_5525,N_5686);
or U6190 (N_6190,N_5962,N_5626);
and U6191 (N_6191,N_5790,N_5602);
or U6192 (N_6192,N_5748,N_5952);
and U6193 (N_6193,N_5891,N_5566);
nand U6194 (N_6194,N_5771,N_5663);
xor U6195 (N_6195,N_5900,N_5914);
or U6196 (N_6196,N_5599,N_5936);
or U6197 (N_6197,N_5745,N_5892);
xnor U6198 (N_6198,N_5850,N_5644);
and U6199 (N_6199,N_5953,N_5866);
nand U6200 (N_6200,N_5638,N_5616);
xnor U6201 (N_6201,N_5538,N_5769);
nor U6202 (N_6202,N_5823,N_5580);
nand U6203 (N_6203,N_5739,N_5811);
or U6204 (N_6204,N_5540,N_5833);
or U6205 (N_6205,N_5967,N_5625);
or U6206 (N_6206,N_5948,N_5601);
or U6207 (N_6207,N_5770,N_5578);
nor U6208 (N_6208,N_5590,N_5682);
xor U6209 (N_6209,N_5768,N_5784);
or U6210 (N_6210,N_5593,N_5895);
or U6211 (N_6211,N_5822,N_5677);
xnor U6212 (N_6212,N_5719,N_5643);
xnor U6213 (N_6213,N_5927,N_5899);
nand U6214 (N_6214,N_5868,N_5993);
xnor U6215 (N_6215,N_5830,N_5828);
and U6216 (N_6216,N_5648,N_5517);
and U6217 (N_6217,N_5939,N_5647);
and U6218 (N_6218,N_5589,N_5877);
nor U6219 (N_6219,N_5785,N_5639);
xor U6220 (N_6220,N_5878,N_5794);
and U6221 (N_6221,N_5988,N_5699);
nand U6222 (N_6222,N_5998,N_5766);
nor U6223 (N_6223,N_5562,N_5920);
nor U6224 (N_6224,N_5749,N_5693);
or U6225 (N_6225,N_5500,N_5516);
and U6226 (N_6226,N_5928,N_5990);
nand U6227 (N_6227,N_5799,N_5960);
and U6228 (N_6228,N_5958,N_5710);
xnor U6229 (N_6229,N_5772,N_5656);
nand U6230 (N_6230,N_5959,N_5744);
nor U6231 (N_6231,N_5584,N_5721);
or U6232 (N_6232,N_5836,N_5591);
nor U6233 (N_6233,N_5781,N_5725);
xor U6234 (N_6234,N_5954,N_5856);
and U6235 (N_6235,N_5527,N_5973);
nand U6236 (N_6236,N_5887,N_5755);
or U6237 (N_6237,N_5615,N_5933);
nor U6238 (N_6238,N_5902,N_5543);
nor U6239 (N_6239,N_5550,N_5796);
or U6240 (N_6240,N_5676,N_5879);
nand U6241 (N_6241,N_5731,N_5665);
or U6242 (N_6242,N_5979,N_5831);
or U6243 (N_6243,N_5871,N_5800);
nor U6244 (N_6244,N_5937,N_5548);
nor U6245 (N_6245,N_5855,N_5834);
nor U6246 (N_6246,N_5910,N_5559);
and U6247 (N_6247,N_5758,N_5827);
and U6248 (N_6248,N_5964,N_5650);
and U6249 (N_6249,N_5810,N_5567);
xor U6250 (N_6250,N_5691,N_5911);
or U6251 (N_6251,N_5642,N_5709);
xnor U6252 (N_6252,N_5813,N_5918);
nor U6253 (N_6253,N_5525,N_5809);
nand U6254 (N_6254,N_5656,N_5557);
or U6255 (N_6255,N_5991,N_5955);
xnor U6256 (N_6256,N_5832,N_5545);
and U6257 (N_6257,N_5915,N_5552);
and U6258 (N_6258,N_5951,N_5738);
nand U6259 (N_6259,N_5814,N_5540);
and U6260 (N_6260,N_5762,N_5984);
or U6261 (N_6261,N_5641,N_5839);
or U6262 (N_6262,N_5882,N_5650);
xor U6263 (N_6263,N_5863,N_5946);
or U6264 (N_6264,N_5830,N_5909);
nor U6265 (N_6265,N_5599,N_5682);
nand U6266 (N_6266,N_5508,N_5749);
or U6267 (N_6267,N_5894,N_5765);
nand U6268 (N_6268,N_5501,N_5796);
or U6269 (N_6269,N_5742,N_5697);
nor U6270 (N_6270,N_5662,N_5770);
nand U6271 (N_6271,N_5996,N_5829);
nand U6272 (N_6272,N_5735,N_5909);
and U6273 (N_6273,N_5707,N_5705);
nor U6274 (N_6274,N_5890,N_5770);
nor U6275 (N_6275,N_5730,N_5639);
xnor U6276 (N_6276,N_5957,N_5799);
and U6277 (N_6277,N_5994,N_5858);
xnor U6278 (N_6278,N_5602,N_5652);
or U6279 (N_6279,N_5547,N_5875);
nand U6280 (N_6280,N_5684,N_5542);
xor U6281 (N_6281,N_5883,N_5506);
and U6282 (N_6282,N_5580,N_5682);
xor U6283 (N_6283,N_5995,N_5616);
and U6284 (N_6284,N_5995,N_5756);
xnor U6285 (N_6285,N_5694,N_5975);
or U6286 (N_6286,N_5711,N_5967);
or U6287 (N_6287,N_5581,N_5861);
and U6288 (N_6288,N_5583,N_5650);
nand U6289 (N_6289,N_5687,N_5619);
nor U6290 (N_6290,N_5531,N_5904);
nand U6291 (N_6291,N_5647,N_5769);
nand U6292 (N_6292,N_5557,N_5781);
and U6293 (N_6293,N_5937,N_5552);
or U6294 (N_6294,N_5874,N_5777);
and U6295 (N_6295,N_5957,N_5626);
nor U6296 (N_6296,N_5813,N_5746);
and U6297 (N_6297,N_5795,N_5886);
nand U6298 (N_6298,N_5629,N_5825);
nand U6299 (N_6299,N_5858,N_5744);
or U6300 (N_6300,N_5930,N_5559);
nand U6301 (N_6301,N_5565,N_5615);
nand U6302 (N_6302,N_5544,N_5743);
or U6303 (N_6303,N_5700,N_5746);
or U6304 (N_6304,N_5608,N_5866);
and U6305 (N_6305,N_5905,N_5939);
xnor U6306 (N_6306,N_5550,N_5951);
and U6307 (N_6307,N_5629,N_5875);
nor U6308 (N_6308,N_5743,N_5559);
xor U6309 (N_6309,N_5769,N_5829);
nand U6310 (N_6310,N_5653,N_5738);
nor U6311 (N_6311,N_5957,N_5951);
nor U6312 (N_6312,N_5605,N_5951);
and U6313 (N_6313,N_5720,N_5584);
or U6314 (N_6314,N_5936,N_5526);
or U6315 (N_6315,N_5550,N_5981);
and U6316 (N_6316,N_5965,N_5873);
or U6317 (N_6317,N_5760,N_5806);
or U6318 (N_6318,N_5779,N_5732);
or U6319 (N_6319,N_5750,N_5947);
nand U6320 (N_6320,N_5690,N_5699);
and U6321 (N_6321,N_5526,N_5517);
nand U6322 (N_6322,N_5585,N_5900);
nor U6323 (N_6323,N_5748,N_5574);
nand U6324 (N_6324,N_5912,N_5948);
nand U6325 (N_6325,N_5813,N_5588);
nor U6326 (N_6326,N_5529,N_5653);
xor U6327 (N_6327,N_5790,N_5963);
and U6328 (N_6328,N_5982,N_5952);
nor U6329 (N_6329,N_5673,N_5842);
nand U6330 (N_6330,N_5708,N_5904);
and U6331 (N_6331,N_5792,N_5822);
and U6332 (N_6332,N_5908,N_5685);
xnor U6333 (N_6333,N_5558,N_5626);
nand U6334 (N_6334,N_5790,N_5991);
nand U6335 (N_6335,N_5890,N_5780);
and U6336 (N_6336,N_5930,N_5608);
nor U6337 (N_6337,N_5882,N_5632);
or U6338 (N_6338,N_5673,N_5546);
nor U6339 (N_6339,N_5614,N_5721);
nand U6340 (N_6340,N_5861,N_5894);
nand U6341 (N_6341,N_5667,N_5576);
nand U6342 (N_6342,N_5966,N_5724);
nand U6343 (N_6343,N_5732,N_5783);
nand U6344 (N_6344,N_5737,N_5744);
nand U6345 (N_6345,N_5636,N_5581);
and U6346 (N_6346,N_5838,N_5683);
xor U6347 (N_6347,N_5612,N_5905);
xnor U6348 (N_6348,N_5570,N_5636);
xnor U6349 (N_6349,N_5801,N_5697);
and U6350 (N_6350,N_5820,N_5841);
nand U6351 (N_6351,N_5972,N_5662);
nor U6352 (N_6352,N_5638,N_5622);
nand U6353 (N_6353,N_5518,N_5511);
nand U6354 (N_6354,N_5980,N_5654);
nor U6355 (N_6355,N_5670,N_5838);
and U6356 (N_6356,N_5613,N_5940);
or U6357 (N_6357,N_5960,N_5985);
nand U6358 (N_6358,N_5584,N_5950);
nor U6359 (N_6359,N_5892,N_5613);
nand U6360 (N_6360,N_5749,N_5880);
nor U6361 (N_6361,N_5872,N_5777);
or U6362 (N_6362,N_5571,N_5805);
nor U6363 (N_6363,N_5766,N_5976);
or U6364 (N_6364,N_5544,N_5612);
or U6365 (N_6365,N_5642,N_5816);
or U6366 (N_6366,N_5839,N_5834);
xnor U6367 (N_6367,N_5687,N_5942);
nand U6368 (N_6368,N_5516,N_5611);
or U6369 (N_6369,N_5607,N_5710);
or U6370 (N_6370,N_5729,N_5954);
or U6371 (N_6371,N_5801,N_5763);
and U6372 (N_6372,N_5965,N_5950);
nor U6373 (N_6373,N_5847,N_5522);
and U6374 (N_6374,N_5753,N_5543);
and U6375 (N_6375,N_5768,N_5926);
and U6376 (N_6376,N_5835,N_5947);
nand U6377 (N_6377,N_5615,N_5898);
and U6378 (N_6378,N_5581,N_5681);
and U6379 (N_6379,N_5965,N_5538);
nor U6380 (N_6380,N_5977,N_5519);
nor U6381 (N_6381,N_5758,N_5974);
or U6382 (N_6382,N_5668,N_5916);
nor U6383 (N_6383,N_5509,N_5678);
nor U6384 (N_6384,N_5828,N_5563);
nand U6385 (N_6385,N_5818,N_5793);
nor U6386 (N_6386,N_5646,N_5969);
or U6387 (N_6387,N_5931,N_5623);
and U6388 (N_6388,N_5585,N_5990);
nand U6389 (N_6389,N_5911,N_5992);
nand U6390 (N_6390,N_5985,N_5794);
nor U6391 (N_6391,N_5979,N_5853);
nor U6392 (N_6392,N_5729,N_5900);
or U6393 (N_6393,N_5937,N_5702);
xnor U6394 (N_6394,N_5855,N_5952);
nand U6395 (N_6395,N_5837,N_5719);
nand U6396 (N_6396,N_5536,N_5836);
nor U6397 (N_6397,N_5773,N_5570);
nand U6398 (N_6398,N_5555,N_5572);
nand U6399 (N_6399,N_5841,N_5592);
and U6400 (N_6400,N_5992,N_5748);
and U6401 (N_6401,N_5908,N_5503);
or U6402 (N_6402,N_5670,N_5901);
or U6403 (N_6403,N_5605,N_5697);
or U6404 (N_6404,N_5644,N_5780);
nor U6405 (N_6405,N_5736,N_5866);
or U6406 (N_6406,N_5977,N_5553);
nand U6407 (N_6407,N_5923,N_5654);
and U6408 (N_6408,N_5970,N_5977);
and U6409 (N_6409,N_5670,N_5608);
or U6410 (N_6410,N_5712,N_5846);
xor U6411 (N_6411,N_5961,N_5603);
or U6412 (N_6412,N_5991,N_5997);
xnor U6413 (N_6413,N_5806,N_5711);
and U6414 (N_6414,N_5638,N_5885);
or U6415 (N_6415,N_5634,N_5625);
and U6416 (N_6416,N_5632,N_5837);
and U6417 (N_6417,N_5860,N_5713);
or U6418 (N_6418,N_5986,N_5569);
and U6419 (N_6419,N_5969,N_5626);
or U6420 (N_6420,N_5624,N_5881);
nor U6421 (N_6421,N_5883,N_5980);
or U6422 (N_6422,N_5927,N_5562);
and U6423 (N_6423,N_5913,N_5541);
or U6424 (N_6424,N_5904,N_5507);
xor U6425 (N_6425,N_5820,N_5618);
xnor U6426 (N_6426,N_5926,N_5996);
nor U6427 (N_6427,N_5585,N_5537);
nand U6428 (N_6428,N_5721,N_5672);
nor U6429 (N_6429,N_5844,N_5678);
or U6430 (N_6430,N_5696,N_5986);
or U6431 (N_6431,N_5841,N_5889);
and U6432 (N_6432,N_5822,N_5763);
and U6433 (N_6433,N_5758,N_5673);
nor U6434 (N_6434,N_5572,N_5629);
and U6435 (N_6435,N_5997,N_5556);
nand U6436 (N_6436,N_5872,N_5948);
nand U6437 (N_6437,N_5555,N_5800);
or U6438 (N_6438,N_5544,N_5516);
or U6439 (N_6439,N_5774,N_5934);
or U6440 (N_6440,N_5521,N_5733);
or U6441 (N_6441,N_5578,N_5582);
nor U6442 (N_6442,N_5606,N_5804);
nand U6443 (N_6443,N_5701,N_5786);
or U6444 (N_6444,N_5917,N_5679);
nand U6445 (N_6445,N_5787,N_5813);
nor U6446 (N_6446,N_5941,N_5712);
nor U6447 (N_6447,N_5664,N_5776);
nor U6448 (N_6448,N_5818,N_5578);
nor U6449 (N_6449,N_5503,N_5649);
nor U6450 (N_6450,N_5812,N_5979);
nand U6451 (N_6451,N_5870,N_5826);
nor U6452 (N_6452,N_5898,N_5827);
or U6453 (N_6453,N_5625,N_5806);
and U6454 (N_6454,N_5916,N_5769);
or U6455 (N_6455,N_5585,N_5941);
nand U6456 (N_6456,N_5756,N_5680);
nor U6457 (N_6457,N_5778,N_5793);
or U6458 (N_6458,N_5659,N_5892);
nand U6459 (N_6459,N_5779,N_5544);
nand U6460 (N_6460,N_5991,N_5915);
nand U6461 (N_6461,N_5943,N_5734);
or U6462 (N_6462,N_5958,N_5633);
nor U6463 (N_6463,N_5901,N_5804);
or U6464 (N_6464,N_5895,N_5849);
nand U6465 (N_6465,N_5798,N_5805);
and U6466 (N_6466,N_5710,N_5964);
nor U6467 (N_6467,N_5599,N_5976);
nor U6468 (N_6468,N_5569,N_5676);
xor U6469 (N_6469,N_5838,N_5998);
nand U6470 (N_6470,N_5826,N_5773);
xnor U6471 (N_6471,N_5875,N_5874);
or U6472 (N_6472,N_5780,N_5810);
nor U6473 (N_6473,N_5702,N_5559);
or U6474 (N_6474,N_5621,N_5550);
or U6475 (N_6475,N_5899,N_5776);
nand U6476 (N_6476,N_5636,N_5622);
or U6477 (N_6477,N_5962,N_5577);
nand U6478 (N_6478,N_5653,N_5566);
or U6479 (N_6479,N_5867,N_5868);
and U6480 (N_6480,N_5998,N_5993);
and U6481 (N_6481,N_5918,N_5816);
and U6482 (N_6482,N_5577,N_5630);
nor U6483 (N_6483,N_5692,N_5668);
nor U6484 (N_6484,N_5754,N_5636);
xor U6485 (N_6485,N_5864,N_5978);
nor U6486 (N_6486,N_5809,N_5794);
or U6487 (N_6487,N_5820,N_5725);
or U6488 (N_6488,N_5647,N_5767);
or U6489 (N_6489,N_5604,N_5827);
nor U6490 (N_6490,N_5745,N_5770);
nand U6491 (N_6491,N_5870,N_5983);
or U6492 (N_6492,N_5792,N_5531);
and U6493 (N_6493,N_5584,N_5710);
and U6494 (N_6494,N_5890,N_5601);
or U6495 (N_6495,N_5703,N_5641);
nand U6496 (N_6496,N_5584,N_5766);
and U6497 (N_6497,N_5627,N_5797);
and U6498 (N_6498,N_5770,N_5690);
and U6499 (N_6499,N_5779,N_5729);
nor U6500 (N_6500,N_6015,N_6017);
and U6501 (N_6501,N_6122,N_6477);
nand U6502 (N_6502,N_6319,N_6311);
nor U6503 (N_6503,N_6199,N_6298);
and U6504 (N_6504,N_6138,N_6348);
or U6505 (N_6505,N_6324,N_6023);
and U6506 (N_6506,N_6293,N_6337);
or U6507 (N_6507,N_6389,N_6192);
nor U6508 (N_6508,N_6271,N_6129);
nor U6509 (N_6509,N_6353,N_6277);
or U6510 (N_6510,N_6069,N_6259);
or U6511 (N_6511,N_6120,N_6180);
or U6512 (N_6512,N_6402,N_6176);
and U6513 (N_6513,N_6254,N_6279);
or U6514 (N_6514,N_6104,N_6431);
or U6515 (N_6515,N_6099,N_6457);
nor U6516 (N_6516,N_6411,N_6083);
nor U6517 (N_6517,N_6081,N_6397);
nand U6518 (N_6518,N_6189,N_6051);
and U6519 (N_6519,N_6170,N_6202);
nand U6520 (N_6520,N_6228,N_6361);
nand U6521 (N_6521,N_6339,N_6472);
or U6522 (N_6522,N_6035,N_6263);
nand U6523 (N_6523,N_6424,N_6173);
and U6524 (N_6524,N_6242,N_6384);
nor U6525 (N_6525,N_6148,N_6018);
nor U6526 (N_6526,N_6327,N_6103);
and U6527 (N_6527,N_6146,N_6299);
or U6528 (N_6528,N_6159,N_6095);
and U6529 (N_6529,N_6195,N_6485);
or U6530 (N_6530,N_6345,N_6190);
nor U6531 (N_6531,N_6031,N_6019);
and U6532 (N_6532,N_6282,N_6371);
nand U6533 (N_6533,N_6325,N_6467);
nor U6534 (N_6534,N_6445,N_6427);
nor U6535 (N_6535,N_6065,N_6399);
nor U6536 (N_6536,N_6128,N_6241);
and U6537 (N_6537,N_6047,N_6063);
nor U6538 (N_6538,N_6243,N_6010);
and U6539 (N_6539,N_6124,N_6370);
or U6540 (N_6540,N_6036,N_6125);
or U6541 (N_6541,N_6048,N_6064);
nor U6542 (N_6542,N_6200,N_6207);
or U6543 (N_6543,N_6471,N_6198);
nor U6544 (N_6544,N_6382,N_6067);
nand U6545 (N_6545,N_6330,N_6123);
nor U6546 (N_6546,N_6486,N_6256);
nor U6547 (N_6547,N_6493,N_6365);
xor U6548 (N_6548,N_6329,N_6496);
or U6549 (N_6549,N_6117,N_6340);
nor U6550 (N_6550,N_6367,N_6283);
nand U6551 (N_6551,N_6459,N_6084);
or U6552 (N_6552,N_6088,N_6321);
nand U6553 (N_6553,N_6196,N_6045);
xor U6554 (N_6554,N_6209,N_6106);
nand U6555 (N_6555,N_6026,N_6404);
nor U6556 (N_6556,N_6091,N_6461);
and U6557 (N_6557,N_6222,N_6420);
nor U6558 (N_6558,N_6226,N_6116);
nor U6559 (N_6559,N_6172,N_6188);
nand U6560 (N_6560,N_6488,N_6494);
and U6561 (N_6561,N_6470,N_6008);
nand U6562 (N_6562,N_6460,N_6272);
nor U6563 (N_6563,N_6113,N_6082);
nand U6564 (N_6564,N_6142,N_6149);
nand U6565 (N_6565,N_6257,N_6166);
nor U6566 (N_6566,N_6364,N_6027);
nand U6567 (N_6567,N_6037,N_6076);
or U6568 (N_6568,N_6267,N_6346);
and U6569 (N_6569,N_6309,N_6174);
nor U6570 (N_6570,N_6033,N_6294);
and U6571 (N_6571,N_6059,N_6347);
and U6572 (N_6572,N_6429,N_6251);
or U6573 (N_6573,N_6422,N_6139);
and U6574 (N_6574,N_6219,N_6187);
and U6575 (N_6575,N_6276,N_6287);
nand U6576 (N_6576,N_6167,N_6409);
and U6577 (N_6577,N_6246,N_6215);
and U6578 (N_6578,N_6410,N_6238);
nor U6579 (N_6579,N_6320,N_6318);
nand U6580 (N_6580,N_6469,N_6075);
nand U6581 (N_6581,N_6105,N_6000);
and U6582 (N_6582,N_6155,N_6157);
and U6583 (N_6583,N_6436,N_6145);
nand U6584 (N_6584,N_6073,N_6499);
nor U6585 (N_6585,N_6297,N_6323);
and U6586 (N_6586,N_6204,N_6233);
nor U6587 (N_6587,N_6093,N_6350);
and U6588 (N_6588,N_6206,N_6418);
nand U6589 (N_6589,N_6398,N_6316);
and U6590 (N_6590,N_6414,N_6401);
nand U6591 (N_6591,N_6230,N_6407);
and U6592 (N_6592,N_6406,N_6450);
or U6593 (N_6593,N_6131,N_6042);
or U6594 (N_6594,N_6086,N_6463);
nor U6595 (N_6595,N_6223,N_6498);
nand U6596 (N_6596,N_6295,N_6214);
or U6597 (N_6597,N_6349,N_6292);
nand U6598 (N_6598,N_6197,N_6400);
nor U6599 (N_6599,N_6383,N_6097);
nor U6600 (N_6600,N_6395,N_6220);
nor U6601 (N_6601,N_6437,N_6250);
nand U6602 (N_6602,N_6003,N_6273);
nor U6603 (N_6603,N_6335,N_6302);
or U6604 (N_6604,N_6090,N_6227);
nor U6605 (N_6605,N_6054,N_6355);
and U6606 (N_6606,N_6185,N_6338);
nor U6607 (N_6607,N_6344,N_6278);
nand U6608 (N_6608,N_6405,N_6438);
nand U6609 (N_6609,N_6009,N_6462);
nand U6610 (N_6610,N_6381,N_6343);
nor U6611 (N_6611,N_6164,N_6456);
or U6612 (N_6612,N_6072,N_6231);
and U6613 (N_6613,N_6213,N_6016);
and U6614 (N_6614,N_6160,N_6151);
or U6615 (N_6615,N_6248,N_6474);
nor U6616 (N_6616,N_6425,N_6432);
and U6617 (N_6617,N_6249,N_6171);
or U6618 (N_6618,N_6183,N_6495);
and U6619 (N_6619,N_6154,N_6265);
nor U6620 (N_6620,N_6479,N_6182);
nand U6621 (N_6621,N_6441,N_6134);
xnor U6622 (N_6622,N_6169,N_6130);
or U6623 (N_6623,N_6394,N_6115);
xor U6624 (N_6624,N_6179,N_6332);
nor U6625 (N_6625,N_6030,N_6034);
or U6626 (N_6626,N_6191,N_6264);
and U6627 (N_6627,N_6218,N_6062);
nand U6628 (N_6628,N_6217,N_6038);
nor U6629 (N_6629,N_6247,N_6268);
nor U6630 (N_6630,N_6181,N_6060);
nand U6631 (N_6631,N_6078,N_6061);
and U6632 (N_6632,N_6162,N_6216);
nand U6633 (N_6633,N_6177,N_6080);
nand U6634 (N_6634,N_6296,N_6101);
and U6635 (N_6635,N_6175,N_6433);
or U6636 (N_6636,N_6390,N_6464);
and U6637 (N_6637,N_6056,N_6290);
nor U6638 (N_6638,N_6133,N_6473);
nor U6639 (N_6639,N_6244,N_6396);
xnor U6640 (N_6640,N_6439,N_6270);
xor U6641 (N_6641,N_6412,N_6237);
nand U6642 (N_6642,N_6458,N_6252);
xnor U6643 (N_6643,N_6025,N_6303);
nand U6644 (N_6644,N_6109,N_6121);
nand U6645 (N_6645,N_6186,N_6225);
xnor U6646 (N_6646,N_6308,N_6356);
xor U6647 (N_6647,N_6255,N_6428);
xor U6648 (N_6648,N_6447,N_6032);
nor U6649 (N_6649,N_6194,N_6150);
and U6650 (N_6650,N_6449,N_6426);
or U6651 (N_6651,N_6313,N_6002);
nor U6652 (N_6652,N_6239,N_6111);
xor U6653 (N_6653,N_6141,N_6011);
or U6654 (N_6654,N_6451,N_6156);
and U6655 (N_6655,N_6068,N_6055);
or U6656 (N_6656,N_6322,N_6126);
or U6657 (N_6657,N_6480,N_6386);
and U6658 (N_6658,N_6261,N_6136);
nor U6659 (N_6659,N_6358,N_6184);
nand U6660 (N_6660,N_6430,N_6229);
nand U6661 (N_6661,N_6342,N_6004);
nor U6662 (N_6662,N_6341,N_6163);
nor U6663 (N_6663,N_6388,N_6286);
or U6664 (N_6664,N_6301,N_6285);
nand U6665 (N_6665,N_6387,N_6373);
nor U6666 (N_6666,N_6333,N_6366);
nor U6667 (N_6667,N_6481,N_6153);
nor U6668 (N_6668,N_6362,N_6391);
and U6669 (N_6669,N_6482,N_6201);
or U6670 (N_6670,N_6108,N_6442);
nand U6671 (N_6671,N_6107,N_6331);
nor U6672 (N_6672,N_6408,N_6168);
nand U6673 (N_6673,N_6492,N_6334);
and U6674 (N_6674,N_6094,N_6434);
nor U6675 (N_6675,N_6374,N_6284);
nor U6676 (N_6676,N_6098,N_6475);
nor U6677 (N_6677,N_6007,N_6363);
and U6678 (N_6678,N_6210,N_6092);
nand U6679 (N_6679,N_6260,N_6147);
or U6680 (N_6680,N_6315,N_6435);
nor U6681 (N_6681,N_6043,N_6288);
nor U6682 (N_6682,N_6127,N_6452);
nor U6683 (N_6683,N_6266,N_6379);
nor U6684 (N_6684,N_6497,N_6118);
nor U6685 (N_6685,N_6314,N_6360);
xor U6686 (N_6686,N_6253,N_6119);
nor U6687 (N_6687,N_6234,N_6484);
or U6688 (N_6688,N_6455,N_6211);
and U6689 (N_6689,N_6368,N_6300);
nand U6690 (N_6690,N_6014,N_6102);
nor U6691 (N_6691,N_6403,N_6205);
and U6692 (N_6692,N_6152,N_6417);
and U6693 (N_6693,N_6491,N_6375);
xnor U6694 (N_6694,N_6240,N_6328);
nand U6695 (N_6695,N_6012,N_6378);
xor U6696 (N_6696,N_6307,N_6245);
or U6697 (N_6697,N_6041,N_6232);
nor U6698 (N_6698,N_6193,N_6376);
or U6699 (N_6699,N_6236,N_6158);
nor U6700 (N_6700,N_6058,N_6085);
nand U6701 (N_6701,N_6212,N_6483);
and U6702 (N_6702,N_6203,N_6028);
or U6703 (N_6703,N_6454,N_6443);
nand U6704 (N_6704,N_6466,N_6306);
nand U6705 (N_6705,N_6066,N_6312);
and U6706 (N_6706,N_6005,N_6446);
or U6707 (N_6707,N_6110,N_6057);
nand U6708 (N_6708,N_6135,N_6413);
or U6709 (N_6709,N_6305,N_6453);
nor U6710 (N_6710,N_6114,N_6489);
and U6711 (N_6711,N_6112,N_6235);
and U6712 (N_6712,N_6224,N_6132);
nand U6713 (N_6713,N_6087,N_6274);
nand U6714 (N_6714,N_6100,N_6354);
nor U6715 (N_6715,N_6079,N_6258);
or U6716 (N_6716,N_6144,N_6074);
and U6717 (N_6717,N_6291,N_6029);
nand U6718 (N_6718,N_6165,N_6415);
and U6719 (N_6719,N_6221,N_6487);
and U6720 (N_6720,N_6369,N_6372);
nand U6721 (N_6721,N_6208,N_6001);
and U6722 (N_6722,N_6289,N_6269);
and U6723 (N_6723,N_6304,N_6444);
nor U6724 (N_6724,N_6049,N_6357);
nand U6725 (N_6725,N_6421,N_6021);
and U6726 (N_6726,N_6351,N_6281);
or U6727 (N_6727,N_6262,N_6020);
and U6728 (N_6728,N_6476,N_6052);
or U6729 (N_6729,N_6352,N_6140);
or U6730 (N_6730,N_6143,N_6416);
or U6731 (N_6731,N_6478,N_6022);
nand U6732 (N_6732,N_6137,N_6280);
and U6733 (N_6733,N_6419,N_6050);
nand U6734 (N_6734,N_6070,N_6465);
nor U6735 (N_6735,N_6440,N_6359);
or U6736 (N_6736,N_6044,N_6393);
nand U6737 (N_6737,N_6040,N_6377);
and U6738 (N_6738,N_6317,N_6071);
or U6739 (N_6739,N_6013,N_6024);
nor U6740 (N_6740,N_6006,N_6096);
nand U6741 (N_6741,N_6046,N_6448);
nand U6742 (N_6742,N_6039,N_6089);
nor U6743 (N_6743,N_6161,N_6423);
nor U6744 (N_6744,N_6178,N_6275);
and U6745 (N_6745,N_6336,N_6468);
and U6746 (N_6746,N_6490,N_6392);
and U6747 (N_6747,N_6077,N_6385);
nand U6748 (N_6748,N_6310,N_6053);
xnor U6749 (N_6749,N_6380,N_6326);
nand U6750 (N_6750,N_6212,N_6274);
xnor U6751 (N_6751,N_6154,N_6454);
or U6752 (N_6752,N_6403,N_6010);
nor U6753 (N_6753,N_6261,N_6151);
or U6754 (N_6754,N_6079,N_6451);
nor U6755 (N_6755,N_6212,N_6378);
or U6756 (N_6756,N_6144,N_6003);
nor U6757 (N_6757,N_6099,N_6391);
and U6758 (N_6758,N_6294,N_6461);
nand U6759 (N_6759,N_6338,N_6456);
and U6760 (N_6760,N_6478,N_6281);
xnor U6761 (N_6761,N_6365,N_6371);
and U6762 (N_6762,N_6021,N_6339);
or U6763 (N_6763,N_6144,N_6336);
nand U6764 (N_6764,N_6413,N_6376);
and U6765 (N_6765,N_6114,N_6144);
or U6766 (N_6766,N_6452,N_6383);
xnor U6767 (N_6767,N_6027,N_6281);
nand U6768 (N_6768,N_6056,N_6348);
nor U6769 (N_6769,N_6120,N_6401);
nor U6770 (N_6770,N_6225,N_6287);
and U6771 (N_6771,N_6456,N_6314);
xnor U6772 (N_6772,N_6144,N_6425);
and U6773 (N_6773,N_6188,N_6379);
or U6774 (N_6774,N_6290,N_6045);
or U6775 (N_6775,N_6043,N_6007);
nor U6776 (N_6776,N_6359,N_6076);
nor U6777 (N_6777,N_6150,N_6113);
nor U6778 (N_6778,N_6488,N_6329);
nand U6779 (N_6779,N_6225,N_6170);
and U6780 (N_6780,N_6243,N_6459);
and U6781 (N_6781,N_6090,N_6167);
and U6782 (N_6782,N_6296,N_6460);
or U6783 (N_6783,N_6334,N_6181);
nor U6784 (N_6784,N_6074,N_6130);
nor U6785 (N_6785,N_6421,N_6301);
nor U6786 (N_6786,N_6376,N_6104);
or U6787 (N_6787,N_6041,N_6133);
nor U6788 (N_6788,N_6228,N_6267);
nand U6789 (N_6789,N_6231,N_6103);
and U6790 (N_6790,N_6259,N_6023);
xnor U6791 (N_6791,N_6277,N_6116);
nand U6792 (N_6792,N_6081,N_6327);
xnor U6793 (N_6793,N_6447,N_6075);
xnor U6794 (N_6794,N_6383,N_6267);
nand U6795 (N_6795,N_6317,N_6034);
and U6796 (N_6796,N_6339,N_6225);
nor U6797 (N_6797,N_6469,N_6354);
nor U6798 (N_6798,N_6228,N_6368);
or U6799 (N_6799,N_6381,N_6092);
and U6800 (N_6800,N_6349,N_6307);
and U6801 (N_6801,N_6323,N_6129);
or U6802 (N_6802,N_6068,N_6112);
nand U6803 (N_6803,N_6235,N_6128);
and U6804 (N_6804,N_6317,N_6456);
xnor U6805 (N_6805,N_6497,N_6257);
nand U6806 (N_6806,N_6485,N_6351);
or U6807 (N_6807,N_6388,N_6010);
nor U6808 (N_6808,N_6470,N_6286);
xor U6809 (N_6809,N_6269,N_6412);
and U6810 (N_6810,N_6200,N_6430);
or U6811 (N_6811,N_6499,N_6480);
or U6812 (N_6812,N_6366,N_6354);
nand U6813 (N_6813,N_6020,N_6281);
or U6814 (N_6814,N_6361,N_6217);
and U6815 (N_6815,N_6349,N_6350);
nand U6816 (N_6816,N_6115,N_6013);
nor U6817 (N_6817,N_6312,N_6413);
nor U6818 (N_6818,N_6446,N_6394);
nand U6819 (N_6819,N_6433,N_6488);
and U6820 (N_6820,N_6302,N_6195);
nand U6821 (N_6821,N_6327,N_6074);
xnor U6822 (N_6822,N_6007,N_6296);
nand U6823 (N_6823,N_6218,N_6293);
and U6824 (N_6824,N_6087,N_6349);
or U6825 (N_6825,N_6213,N_6130);
or U6826 (N_6826,N_6291,N_6312);
and U6827 (N_6827,N_6398,N_6016);
and U6828 (N_6828,N_6445,N_6193);
or U6829 (N_6829,N_6158,N_6089);
or U6830 (N_6830,N_6373,N_6284);
and U6831 (N_6831,N_6229,N_6311);
and U6832 (N_6832,N_6488,N_6135);
nand U6833 (N_6833,N_6293,N_6129);
nand U6834 (N_6834,N_6332,N_6278);
and U6835 (N_6835,N_6342,N_6079);
nand U6836 (N_6836,N_6029,N_6396);
and U6837 (N_6837,N_6262,N_6113);
nand U6838 (N_6838,N_6300,N_6256);
nand U6839 (N_6839,N_6031,N_6355);
nor U6840 (N_6840,N_6129,N_6438);
nand U6841 (N_6841,N_6397,N_6346);
xor U6842 (N_6842,N_6095,N_6011);
nor U6843 (N_6843,N_6066,N_6272);
nor U6844 (N_6844,N_6201,N_6269);
and U6845 (N_6845,N_6381,N_6495);
xor U6846 (N_6846,N_6459,N_6206);
nor U6847 (N_6847,N_6387,N_6418);
or U6848 (N_6848,N_6372,N_6425);
nor U6849 (N_6849,N_6349,N_6166);
xnor U6850 (N_6850,N_6058,N_6032);
nor U6851 (N_6851,N_6070,N_6240);
or U6852 (N_6852,N_6288,N_6084);
xnor U6853 (N_6853,N_6316,N_6373);
xor U6854 (N_6854,N_6439,N_6008);
or U6855 (N_6855,N_6232,N_6450);
nand U6856 (N_6856,N_6046,N_6372);
and U6857 (N_6857,N_6097,N_6113);
xnor U6858 (N_6858,N_6100,N_6242);
nand U6859 (N_6859,N_6306,N_6308);
xnor U6860 (N_6860,N_6153,N_6284);
and U6861 (N_6861,N_6371,N_6097);
or U6862 (N_6862,N_6188,N_6021);
or U6863 (N_6863,N_6372,N_6348);
nand U6864 (N_6864,N_6192,N_6380);
and U6865 (N_6865,N_6390,N_6474);
and U6866 (N_6866,N_6157,N_6185);
nand U6867 (N_6867,N_6388,N_6099);
or U6868 (N_6868,N_6323,N_6065);
or U6869 (N_6869,N_6136,N_6140);
nand U6870 (N_6870,N_6172,N_6037);
nand U6871 (N_6871,N_6375,N_6032);
nand U6872 (N_6872,N_6295,N_6326);
nand U6873 (N_6873,N_6335,N_6260);
or U6874 (N_6874,N_6255,N_6365);
xnor U6875 (N_6875,N_6361,N_6085);
nor U6876 (N_6876,N_6056,N_6033);
nor U6877 (N_6877,N_6118,N_6138);
and U6878 (N_6878,N_6335,N_6331);
nor U6879 (N_6879,N_6429,N_6283);
xnor U6880 (N_6880,N_6480,N_6037);
nand U6881 (N_6881,N_6373,N_6313);
xnor U6882 (N_6882,N_6327,N_6087);
and U6883 (N_6883,N_6032,N_6160);
nor U6884 (N_6884,N_6288,N_6083);
nor U6885 (N_6885,N_6211,N_6183);
or U6886 (N_6886,N_6054,N_6498);
nand U6887 (N_6887,N_6348,N_6496);
and U6888 (N_6888,N_6462,N_6360);
and U6889 (N_6889,N_6158,N_6377);
and U6890 (N_6890,N_6371,N_6090);
or U6891 (N_6891,N_6272,N_6273);
nor U6892 (N_6892,N_6417,N_6279);
nand U6893 (N_6893,N_6245,N_6084);
nand U6894 (N_6894,N_6283,N_6306);
or U6895 (N_6895,N_6158,N_6173);
nand U6896 (N_6896,N_6402,N_6070);
or U6897 (N_6897,N_6235,N_6319);
or U6898 (N_6898,N_6102,N_6291);
xnor U6899 (N_6899,N_6460,N_6001);
xnor U6900 (N_6900,N_6061,N_6119);
nor U6901 (N_6901,N_6437,N_6225);
nand U6902 (N_6902,N_6024,N_6389);
and U6903 (N_6903,N_6429,N_6326);
nand U6904 (N_6904,N_6111,N_6331);
or U6905 (N_6905,N_6069,N_6271);
xor U6906 (N_6906,N_6449,N_6089);
and U6907 (N_6907,N_6304,N_6181);
nand U6908 (N_6908,N_6124,N_6123);
nand U6909 (N_6909,N_6211,N_6180);
or U6910 (N_6910,N_6305,N_6129);
or U6911 (N_6911,N_6426,N_6019);
and U6912 (N_6912,N_6142,N_6094);
and U6913 (N_6913,N_6375,N_6137);
nand U6914 (N_6914,N_6064,N_6418);
nor U6915 (N_6915,N_6361,N_6336);
nand U6916 (N_6916,N_6240,N_6309);
xnor U6917 (N_6917,N_6238,N_6327);
nor U6918 (N_6918,N_6475,N_6439);
and U6919 (N_6919,N_6305,N_6169);
nor U6920 (N_6920,N_6033,N_6096);
or U6921 (N_6921,N_6223,N_6413);
or U6922 (N_6922,N_6467,N_6214);
xor U6923 (N_6923,N_6342,N_6244);
and U6924 (N_6924,N_6122,N_6252);
nand U6925 (N_6925,N_6061,N_6002);
and U6926 (N_6926,N_6348,N_6420);
nor U6927 (N_6927,N_6384,N_6499);
and U6928 (N_6928,N_6139,N_6126);
nor U6929 (N_6929,N_6150,N_6247);
nand U6930 (N_6930,N_6470,N_6079);
or U6931 (N_6931,N_6088,N_6091);
nor U6932 (N_6932,N_6004,N_6345);
or U6933 (N_6933,N_6339,N_6213);
nor U6934 (N_6934,N_6187,N_6349);
and U6935 (N_6935,N_6120,N_6433);
or U6936 (N_6936,N_6489,N_6013);
nor U6937 (N_6937,N_6446,N_6051);
nand U6938 (N_6938,N_6269,N_6183);
xor U6939 (N_6939,N_6215,N_6134);
or U6940 (N_6940,N_6311,N_6184);
or U6941 (N_6941,N_6479,N_6275);
nand U6942 (N_6942,N_6091,N_6245);
xnor U6943 (N_6943,N_6233,N_6076);
and U6944 (N_6944,N_6254,N_6223);
nand U6945 (N_6945,N_6372,N_6403);
nor U6946 (N_6946,N_6163,N_6016);
nor U6947 (N_6947,N_6468,N_6399);
or U6948 (N_6948,N_6053,N_6092);
and U6949 (N_6949,N_6213,N_6195);
nor U6950 (N_6950,N_6054,N_6484);
and U6951 (N_6951,N_6029,N_6019);
nor U6952 (N_6952,N_6409,N_6164);
and U6953 (N_6953,N_6029,N_6431);
nand U6954 (N_6954,N_6086,N_6056);
or U6955 (N_6955,N_6045,N_6430);
and U6956 (N_6956,N_6276,N_6033);
xnor U6957 (N_6957,N_6089,N_6152);
or U6958 (N_6958,N_6424,N_6105);
xor U6959 (N_6959,N_6046,N_6234);
nand U6960 (N_6960,N_6210,N_6010);
nand U6961 (N_6961,N_6401,N_6475);
nor U6962 (N_6962,N_6128,N_6169);
and U6963 (N_6963,N_6235,N_6377);
nor U6964 (N_6964,N_6498,N_6366);
nor U6965 (N_6965,N_6059,N_6453);
nor U6966 (N_6966,N_6277,N_6239);
or U6967 (N_6967,N_6220,N_6010);
nand U6968 (N_6968,N_6155,N_6443);
nand U6969 (N_6969,N_6334,N_6021);
nand U6970 (N_6970,N_6172,N_6203);
or U6971 (N_6971,N_6262,N_6441);
and U6972 (N_6972,N_6030,N_6109);
nor U6973 (N_6973,N_6258,N_6177);
xnor U6974 (N_6974,N_6371,N_6464);
nand U6975 (N_6975,N_6255,N_6019);
and U6976 (N_6976,N_6495,N_6174);
nand U6977 (N_6977,N_6323,N_6417);
nor U6978 (N_6978,N_6275,N_6433);
nand U6979 (N_6979,N_6273,N_6253);
nor U6980 (N_6980,N_6204,N_6265);
nand U6981 (N_6981,N_6077,N_6177);
or U6982 (N_6982,N_6407,N_6431);
nand U6983 (N_6983,N_6325,N_6050);
nand U6984 (N_6984,N_6284,N_6348);
and U6985 (N_6985,N_6233,N_6349);
or U6986 (N_6986,N_6424,N_6298);
nand U6987 (N_6987,N_6172,N_6394);
or U6988 (N_6988,N_6475,N_6286);
and U6989 (N_6989,N_6167,N_6480);
nand U6990 (N_6990,N_6491,N_6419);
nor U6991 (N_6991,N_6242,N_6245);
nor U6992 (N_6992,N_6442,N_6008);
or U6993 (N_6993,N_6038,N_6036);
or U6994 (N_6994,N_6390,N_6070);
nor U6995 (N_6995,N_6421,N_6391);
and U6996 (N_6996,N_6335,N_6356);
nand U6997 (N_6997,N_6170,N_6067);
and U6998 (N_6998,N_6315,N_6073);
nand U6999 (N_6999,N_6017,N_6063);
or U7000 (N_7000,N_6771,N_6927);
xnor U7001 (N_7001,N_6722,N_6526);
and U7002 (N_7002,N_6732,N_6843);
and U7003 (N_7003,N_6877,N_6822);
or U7004 (N_7004,N_6667,N_6781);
and U7005 (N_7005,N_6511,N_6948);
nand U7006 (N_7006,N_6879,N_6565);
or U7007 (N_7007,N_6903,N_6514);
and U7008 (N_7008,N_6713,N_6718);
nand U7009 (N_7009,N_6500,N_6973);
and U7010 (N_7010,N_6640,N_6631);
or U7011 (N_7011,N_6795,N_6699);
or U7012 (N_7012,N_6712,N_6833);
nor U7013 (N_7013,N_6630,N_6842);
nor U7014 (N_7014,N_6706,N_6730);
or U7015 (N_7015,N_6900,N_6610);
xnor U7016 (N_7016,N_6536,N_6543);
nor U7017 (N_7017,N_6887,N_6996);
nand U7018 (N_7018,N_6673,N_6841);
or U7019 (N_7019,N_6666,N_6624);
and U7020 (N_7020,N_6837,N_6951);
and U7021 (N_7021,N_6937,N_6763);
nor U7022 (N_7022,N_6978,N_6683);
nor U7023 (N_7023,N_6794,N_6988);
and U7024 (N_7024,N_6603,N_6663);
nand U7025 (N_7025,N_6733,N_6827);
nor U7026 (N_7026,N_6995,N_6784);
nand U7027 (N_7027,N_6589,N_6648);
and U7028 (N_7028,N_6605,N_6654);
and U7029 (N_7029,N_6906,N_6510);
nand U7030 (N_7030,N_6588,N_6925);
nor U7031 (N_7031,N_6749,N_6670);
nor U7032 (N_7032,N_6919,N_6507);
and U7033 (N_7033,N_6846,N_6739);
nand U7034 (N_7034,N_6960,N_6793);
or U7035 (N_7035,N_6930,N_6556);
nand U7036 (N_7036,N_6518,N_6554);
and U7037 (N_7037,N_6936,N_6869);
or U7038 (N_7038,N_6862,N_6891);
or U7039 (N_7039,N_6899,N_6594);
nor U7040 (N_7040,N_6765,N_6885);
nor U7041 (N_7041,N_6724,N_6884);
nor U7042 (N_7042,N_6609,N_6987);
or U7043 (N_7043,N_6644,N_6786);
xor U7044 (N_7044,N_6551,N_6705);
nand U7045 (N_7045,N_6519,N_6883);
xnor U7046 (N_7046,N_6637,N_6621);
nand U7047 (N_7047,N_6611,N_6952);
nand U7048 (N_7048,N_6874,N_6503);
nand U7049 (N_7049,N_6704,N_6939);
or U7050 (N_7050,N_6620,N_6901);
nand U7051 (N_7051,N_6878,N_6791);
nand U7052 (N_7052,N_6632,N_6672);
xnor U7053 (N_7053,N_6715,N_6546);
nand U7054 (N_7054,N_6855,N_6854);
nor U7055 (N_7055,N_6954,N_6687);
and U7056 (N_7056,N_6780,N_6820);
and U7057 (N_7057,N_6623,N_6613);
nor U7058 (N_7058,N_6922,N_6686);
nand U7059 (N_7059,N_6591,N_6753);
nand U7060 (N_7060,N_6652,N_6680);
and U7061 (N_7061,N_6586,N_6950);
or U7062 (N_7062,N_6889,N_6559);
and U7063 (N_7063,N_6516,N_6831);
and U7064 (N_7064,N_6677,N_6612);
nor U7065 (N_7065,N_6545,N_6512);
and U7066 (N_7066,N_6804,N_6560);
nand U7067 (N_7067,N_6596,N_6671);
nor U7068 (N_7068,N_6964,N_6557);
nand U7069 (N_7069,N_6984,N_6721);
or U7070 (N_7070,N_6727,N_6701);
xor U7071 (N_7071,N_6608,N_6832);
nand U7072 (N_7072,N_6698,N_6576);
xnor U7073 (N_7073,N_6575,N_6912);
xnor U7074 (N_7074,N_6805,N_6916);
or U7075 (N_7075,N_6982,N_6897);
nand U7076 (N_7076,N_6505,N_6849);
or U7077 (N_7077,N_6751,N_6711);
or U7078 (N_7078,N_6634,N_6776);
and U7079 (N_7079,N_6639,N_6834);
or U7080 (N_7080,N_6895,N_6657);
and U7081 (N_7081,N_6726,N_6797);
nor U7082 (N_7082,N_6983,N_6653);
or U7083 (N_7083,N_6756,N_6907);
and U7084 (N_7084,N_6812,N_6898);
nor U7085 (N_7085,N_6650,N_6602);
and U7086 (N_7086,N_6920,N_6940);
and U7087 (N_7087,N_6892,N_6864);
or U7088 (N_7088,N_6537,N_6741);
and U7089 (N_7089,N_6583,N_6643);
or U7090 (N_7090,N_6770,N_6723);
nand U7091 (N_7091,N_6584,N_6803);
xnor U7092 (N_7092,N_6835,N_6953);
nand U7093 (N_7093,N_6913,N_6863);
and U7094 (N_7094,N_6959,N_6738);
nand U7095 (N_7095,N_6865,N_6761);
and U7096 (N_7096,N_6777,N_6798);
nor U7097 (N_7097,N_6572,N_6764);
nor U7098 (N_7098,N_6775,N_6994);
and U7099 (N_7099,N_6685,N_6946);
xnor U7100 (N_7100,N_6853,N_6923);
nor U7101 (N_7101,N_6998,N_6580);
nand U7102 (N_7102,N_6532,N_6905);
nand U7103 (N_7103,N_6789,N_6772);
or U7104 (N_7104,N_6689,N_6548);
and U7105 (N_7105,N_6720,N_6910);
and U7106 (N_7106,N_6755,N_6840);
and U7107 (N_7107,N_6601,N_6562);
and U7108 (N_7108,N_6915,N_6924);
nand U7109 (N_7109,N_6845,N_6989);
xor U7110 (N_7110,N_6993,N_6825);
and U7111 (N_7111,N_6675,N_6728);
or U7112 (N_7112,N_6968,N_6824);
and U7113 (N_7113,N_6540,N_6979);
nand U7114 (N_7114,N_6563,N_6676);
or U7115 (N_7115,N_6972,N_6760);
or U7116 (N_7116,N_6578,N_6719);
or U7117 (N_7117,N_6986,N_6649);
nand U7118 (N_7118,N_6808,N_6800);
nor U7119 (N_7119,N_6544,N_6867);
nand U7120 (N_7120,N_6528,N_6921);
xnor U7121 (N_7121,N_6607,N_6525);
or U7122 (N_7122,N_6681,N_6944);
nor U7123 (N_7123,N_6876,N_6541);
or U7124 (N_7124,N_6882,N_6933);
nor U7125 (N_7125,N_6547,N_6538);
nor U7126 (N_7126,N_6860,N_6646);
and U7127 (N_7127,N_6754,N_6521);
nor U7128 (N_7128,N_6758,N_6707);
nor U7129 (N_7129,N_6748,N_6714);
xnor U7130 (N_7130,N_6515,N_6896);
and U7131 (N_7131,N_6599,N_6617);
nor U7132 (N_7132,N_6660,N_6684);
or U7133 (N_7133,N_6848,N_6931);
or U7134 (N_7134,N_6830,N_6941);
and U7135 (N_7135,N_6622,N_6585);
and U7136 (N_7136,N_6809,N_6524);
nand U7137 (N_7137,N_6963,N_6504);
nand U7138 (N_7138,N_6980,N_6956);
or U7139 (N_7139,N_6629,N_6881);
and U7140 (N_7140,N_6935,N_6582);
and U7141 (N_7141,N_6625,N_6938);
xnor U7142 (N_7142,N_6796,N_6542);
and U7143 (N_7143,N_6813,N_6807);
or U7144 (N_7144,N_6806,N_6725);
or U7145 (N_7145,N_6592,N_6579);
or U7146 (N_7146,N_6947,N_6564);
nor U7147 (N_7147,N_6651,N_6971);
nand U7148 (N_7148,N_6774,N_6904);
and U7149 (N_7149,N_6549,N_6600);
and U7150 (N_7150,N_6506,N_6619);
nor U7151 (N_7151,N_6949,N_6945);
and U7152 (N_7152,N_6615,N_6970);
or U7153 (N_7153,N_6703,N_6742);
nand U7154 (N_7154,N_6688,N_6955);
xor U7155 (N_7155,N_6597,N_6523);
xnor U7156 (N_7156,N_6614,N_6908);
and U7157 (N_7157,N_6783,N_6981);
nand U7158 (N_7158,N_6735,N_6839);
and U7159 (N_7159,N_6561,N_6871);
nand U7160 (N_7160,N_6569,N_6766);
and U7161 (N_7161,N_6768,N_6858);
and U7162 (N_7162,N_6875,N_6550);
and U7163 (N_7163,N_6926,N_6692);
and U7164 (N_7164,N_6836,N_6659);
and U7165 (N_7165,N_6967,N_6759);
and U7166 (N_7166,N_6740,N_6785);
nand U7167 (N_7167,N_6792,N_6587);
or U7168 (N_7168,N_6818,N_6870);
nor U7169 (N_7169,N_6976,N_6581);
and U7170 (N_7170,N_6888,N_6917);
nand U7171 (N_7171,N_6838,N_6570);
nand U7172 (N_7172,N_6911,N_6509);
and U7173 (N_7173,N_6856,N_6520);
nor U7174 (N_7174,N_6873,N_6850);
xor U7175 (N_7175,N_6767,N_6731);
nand U7176 (N_7176,N_6778,N_6606);
and U7177 (N_7177,N_6574,N_6568);
nand U7178 (N_7178,N_6802,N_6501);
xor U7179 (N_7179,N_6716,N_6868);
or U7180 (N_7180,N_6969,N_6961);
nor U7181 (N_7181,N_6655,N_6943);
xnor U7182 (N_7182,N_6866,N_6508);
and U7183 (N_7183,N_6678,N_6664);
and U7184 (N_7184,N_6529,N_6577);
or U7185 (N_7185,N_6958,N_6788);
and U7186 (N_7186,N_6997,N_6992);
and U7187 (N_7187,N_6593,N_6799);
nand U7188 (N_7188,N_6890,N_6934);
nor U7189 (N_7189,N_6844,N_6750);
or U7190 (N_7190,N_6555,N_6618);
xnor U7191 (N_7191,N_6962,N_6902);
and U7192 (N_7192,N_6635,N_6928);
and U7193 (N_7193,N_6815,N_6914);
xnor U7194 (N_7194,N_6734,N_6513);
xnor U7195 (N_7195,N_6736,N_6880);
and U7196 (N_7196,N_6595,N_6814);
nand U7197 (N_7197,N_6893,N_6690);
nor U7198 (N_7198,N_6918,N_6744);
and U7199 (N_7199,N_6694,N_6700);
or U7200 (N_7200,N_6737,N_6787);
nand U7201 (N_7201,N_6656,N_6757);
nand U7202 (N_7202,N_6747,N_6645);
nor U7203 (N_7203,N_6762,N_6627);
xnor U7204 (N_7204,N_6985,N_6616);
or U7205 (N_7205,N_6826,N_6682);
or U7206 (N_7206,N_6782,N_6886);
and U7207 (N_7207,N_6991,N_6558);
nor U7208 (N_7208,N_6571,N_6567);
nor U7209 (N_7209,N_6823,N_6861);
or U7210 (N_7210,N_6533,N_6531);
and U7211 (N_7211,N_6790,N_6851);
or U7212 (N_7212,N_6932,N_6647);
nor U7213 (N_7213,N_6717,N_6965);
or U7214 (N_7214,N_6633,N_6909);
nor U7215 (N_7215,N_6668,N_6658);
nor U7216 (N_7216,N_6642,N_6810);
and U7217 (N_7217,N_6502,N_6828);
nor U7218 (N_7218,N_6817,N_6710);
nand U7219 (N_7219,N_6696,N_6852);
or U7220 (N_7220,N_6566,N_6527);
or U7221 (N_7221,N_6534,N_6821);
xor U7222 (N_7222,N_6708,N_6590);
nand U7223 (N_7223,N_6829,N_6957);
or U7224 (N_7224,N_6999,N_6819);
and U7225 (N_7225,N_6636,N_6894);
and U7226 (N_7226,N_6769,N_6779);
and U7227 (N_7227,N_6816,N_6872);
xor U7228 (N_7228,N_6517,N_6729);
or U7229 (N_7229,N_6535,N_6641);
nor U7230 (N_7230,N_6674,N_6553);
nor U7231 (N_7231,N_6966,N_6697);
or U7232 (N_7232,N_6626,N_6665);
and U7233 (N_7233,N_6628,N_6975);
nand U7234 (N_7234,N_6709,N_6604);
nand U7235 (N_7235,N_6801,N_6638);
xnor U7236 (N_7236,N_6811,N_6746);
or U7237 (N_7237,N_6679,N_6702);
nor U7238 (N_7238,N_6522,N_6929);
nand U7239 (N_7239,N_6743,N_6859);
and U7240 (N_7240,N_6773,N_6661);
or U7241 (N_7241,N_6695,N_6857);
nand U7242 (N_7242,N_6669,N_6990);
and U7243 (N_7243,N_6539,N_6691);
and U7244 (N_7244,N_6974,N_6752);
or U7245 (N_7245,N_6745,N_6847);
nand U7246 (N_7246,N_6573,N_6662);
and U7247 (N_7247,N_6693,N_6942);
or U7248 (N_7248,N_6977,N_6552);
or U7249 (N_7249,N_6530,N_6598);
nand U7250 (N_7250,N_6829,N_6714);
and U7251 (N_7251,N_6875,N_6824);
or U7252 (N_7252,N_6963,N_6940);
or U7253 (N_7253,N_6757,N_6848);
and U7254 (N_7254,N_6995,N_6881);
nor U7255 (N_7255,N_6618,N_6808);
or U7256 (N_7256,N_6819,N_6764);
nand U7257 (N_7257,N_6627,N_6523);
nand U7258 (N_7258,N_6909,N_6907);
and U7259 (N_7259,N_6674,N_6704);
xor U7260 (N_7260,N_6847,N_6508);
xnor U7261 (N_7261,N_6519,N_6534);
or U7262 (N_7262,N_6842,N_6973);
xor U7263 (N_7263,N_6816,N_6640);
and U7264 (N_7264,N_6748,N_6799);
nor U7265 (N_7265,N_6757,N_6875);
nand U7266 (N_7266,N_6507,N_6739);
nand U7267 (N_7267,N_6880,N_6664);
and U7268 (N_7268,N_6580,N_6820);
or U7269 (N_7269,N_6699,N_6593);
and U7270 (N_7270,N_6858,N_6502);
nand U7271 (N_7271,N_6722,N_6555);
nand U7272 (N_7272,N_6679,N_6516);
nand U7273 (N_7273,N_6523,N_6754);
nor U7274 (N_7274,N_6556,N_6792);
and U7275 (N_7275,N_6753,N_6821);
and U7276 (N_7276,N_6710,N_6806);
and U7277 (N_7277,N_6824,N_6752);
or U7278 (N_7278,N_6659,N_6974);
or U7279 (N_7279,N_6750,N_6617);
nor U7280 (N_7280,N_6953,N_6524);
nor U7281 (N_7281,N_6951,N_6516);
nor U7282 (N_7282,N_6789,N_6810);
nor U7283 (N_7283,N_6714,N_6626);
and U7284 (N_7284,N_6796,N_6901);
nand U7285 (N_7285,N_6553,N_6548);
nor U7286 (N_7286,N_6627,N_6632);
or U7287 (N_7287,N_6998,N_6881);
and U7288 (N_7288,N_6934,N_6505);
nor U7289 (N_7289,N_6663,N_6617);
xnor U7290 (N_7290,N_6697,N_6628);
and U7291 (N_7291,N_6910,N_6569);
and U7292 (N_7292,N_6507,N_6869);
and U7293 (N_7293,N_6614,N_6805);
nor U7294 (N_7294,N_6762,N_6976);
or U7295 (N_7295,N_6505,N_6595);
or U7296 (N_7296,N_6969,N_6625);
and U7297 (N_7297,N_6585,N_6537);
nor U7298 (N_7298,N_6777,N_6737);
or U7299 (N_7299,N_6959,N_6964);
and U7300 (N_7300,N_6807,N_6792);
nor U7301 (N_7301,N_6721,N_6594);
or U7302 (N_7302,N_6849,N_6682);
or U7303 (N_7303,N_6743,N_6546);
and U7304 (N_7304,N_6623,N_6881);
or U7305 (N_7305,N_6940,N_6954);
and U7306 (N_7306,N_6810,N_6726);
xor U7307 (N_7307,N_6744,N_6848);
xnor U7308 (N_7308,N_6513,N_6596);
or U7309 (N_7309,N_6844,N_6687);
xnor U7310 (N_7310,N_6885,N_6764);
and U7311 (N_7311,N_6528,N_6694);
and U7312 (N_7312,N_6741,N_6670);
xor U7313 (N_7313,N_6833,N_6906);
or U7314 (N_7314,N_6959,N_6520);
nor U7315 (N_7315,N_6833,N_6797);
nor U7316 (N_7316,N_6600,N_6763);
and U7317 (N_7317,N_6855,N_6683);
and U7318 (N_7318,N_6559,N_6827);
xor U7319 (N_7319,N_6727,N_6517);
or U7320 (N_7320,N_6984,N_6884);
or U7321 (N_7321,N_6859,N_6512);
nand U7322 (N_7322,N_6724,N_6807);
or U7323 (N_7323,N_6857,N_6504);
nand U7324 (N_7324,N_6560,N_6887);
nand U7325 (N_7325,N_6799,N_6587);
xor U7326 (N_7326,N_6662,N_6744);
and U7327 (N_7327,N_6705,N_6747);
nand U7328 (N_7328,N_6530,N_6779);
xor U7329 (N_7329,N_6790,N_6930);
and U7330 (N_7330,N_6634,N_6785);
nor U7331 (N_7331,N_6835,N_6587);
nor U7332 (N_7332,N_6502,N_6713);
nand U7333 (N_7333,N_6611,N_6719);
and U7334 (N_7334,N_6702,N_6984);
xor U7335 (N_7335,N_6542,N_6877);
nor U7336 (N_7336,N_6626,N_6757);
or U7337 (N_7337,N_6715,N_6527);
nand U7338 (N_7338,N_6627,N_6778);
nand U7339 (N_7339,N_6911,N_6969);
nand U7340 (N_7340,N_6517,N_6879);
nor U7341 (N_7341,N_6965,N_6938);
and U7342 (N_7342,N_6900,N_6798);
and U7343 (N_7343,N_6539,N_6574);
and U7344 (N_7344,N_6804,N_6598);
and U7345 (N_7345,N_6701,N_6756);
or U7346 (N_7346,N_6692,N_6579);
xnor U7347 (N_7347,N_6562,N_6644);
or U7348 (N_7348,N_6943,N_6945);
and U7349 (N_7349,N_6962,N_6573);
or U7350 (N_7350,N_6754,N_6965);
nor U7351 (N_7351,N_6830,N_6702);
and U7352 (N_7352,N_6917,N_6656);
and U7353 (N_7353,N_6724,N_6735);
nor U7354 (N_7354,N_6529,N_6899);
and U7355 (N_7355,N_6707,N_6621);
or U7356 (N_7356,N_6617,N_6837);
nand U7357 (N_7357,N_6740,N_6733);
and U7358 (N_7358,N_6801,N_6875);
xnor U7359 (N_7359,N_6880,N_6659);
nor U7360 (N_7360,N_6977,N_6984);
xor U7361 (N_7361,N_6602,N_6691);
or U7362 (N_7362,N_6506,N_6677);
and U7363 (N_7363,N_6600,N_6657);
xnor U7364 (N_7364,N_6717,N_6877);
xor U7365 (N_7365,N_6771,N_6677);
and U7366 (N_7366,N_6763,N_6813);
and U7367 (N_7367,N_6894,N_6771);
nand U7368 (N_7368,N_6912,N_6800);
and U7369 (N_7369,N_6644,N_6967);
nand U7370 (N_7370,N_6515,N_6963);
nand U7371 (N_7371,N_6774,N_6811);
nor U7372 (N_7372,N_6651,N_6981);
nand U7373 (N_7373,N_6758,N_6907);
nor U7374 (N_7374,N_6737,N_6628);
xor U7375 (N_7375,N_6958,N_6690);
and U7376 (N_7376,N_6901,N_6956);
and U7377 (N_7377,N_6974,N_6845);
xnor U7378 (N_7378,N_6796,N_6665);
or U7379 (N_7379,N_6686,N_6703);
nor U7380 (N_7380,N_6830,N_6976);
nor U7381 (N_7381,N_6851,N_6761);
xor U7382 (N_7382,N_6601,N_6936);
nor U7383 (N_7383,N_6730,N_6678);
nand U7384 (N_7384,N_6705,N_6781);
or U7385 (N_7385,N_6802,N_6573);
and U7386 (N_7386,N_6956,N_6623);
nand U7387 (N_7387,N_6863,N_6942);
nand U7388 (N_7388,N_6982,N_6736);
xnor U7389 (N_7389,N_6884,N_6862);
xnor U7390 (N_7390,N_6812,N_6615);
or U7391 (N_7391,N_6873,N_6809);
and U7392 (N_7392,N_6570,N_6928);
nand U7393 (N_7393,N_6626,N_6505);
nand U7394 (N_7394,N_6948,N_6861);
nand U7395 (N_7395,N_6821,N_6591);
nor U7396 (N_7396,N_6962,N_6646);
nor U7397 (N_7397,N_6822,N_6961);
and U7398 (N_7398,N_6588,N_6743);
nand U7399 (N_7399,N_6599,N_6990);
or U7400 (N_7400,N_6900,N_6754);
nor U7401 (N_7401,N_6935,N_6788);
or U7402 (N_7402,N_6989,N_6622);
or U7403 (N_7403,N_6506,N_6887);
nor U7404 (N_7404,N_6851,N_6922);
nor U7405 (N_7405,N_6850,N_6533);
xnor U7406 (N_7406,N_6719,N_6625);
nand U7407 (N_7407,N_6954,N_6567);
nand U7408 (N_7408,N_6739,N_6747);
or U7409 (N_7409,N_6563,N_6720);
xor U7410 (N_7410,N_6693,N_6930);
and U7411 (N_7411,N_6812,N_6918);
or U7412 (N_7412,N_6846,N_6566);
nor U7413 (N_7413,N_6672,N_6795);
or U7414 (N_7414,N_6955,N_6951);
nor U7415 (N_7415,N_6662,N_6835);
nor U7416 (N_7416,N_6515,N_6571);
nand U7417 (N_7417,N_6834,N_6584);
and U7418 (N_7418,N_6646,N_6727);
xor U7419 (N_7419,N_6923,N_6760);
and U7420 (N_7420,N_6882,N_6862);
xnor U7421 (N_7421,N_6548,N_6715);
nand U7422 (N_7422,N_6827,N_6757);
nand U7423 (N_7423,N_6918,N_6977);
nand U7424 (N_7424,N_6638,N_6814);
or U7425 (N_7425,N_6679,N_6593);
nor U7426 (N_7426,N_6724,N_6613);
or U7427 (N_7427,N_6855,N_6593);
nor U7428 (N_7428,N_6586,N_6615);
nand U7429 (N_7429,N_6904,N_6698);
or U7430 (N_7430,N_6810,N_6840);
and U7431 (N_7431,N_6660,N_6675);
nand U7432 (N_7432,N_6657,N_6894);
nand U7433 (N_7433,N_6864,N_6803);
or U7434 (N_7434,N_6836,N_6635);
xor U7435 (N_7435,N_6996,N_6828);
nor U7436 (N_7436,N_6630,N_6923);
or U7437 (N_7437,N_6645,N_6574);
xor U7438 (N_7438,N_6666,N_6595);
and U7439 (N_7439,N_6555,N_6713);
xnor U7440 (N_7440,N_6524,N_6897);
or U7441 (N_7441,N_6700,N_6678);
and U7442 (N_7442,N_6998,N_6596);
and U7443 (N_7443,N_6529,N_6875);
and U7444 (N_7444,N_6570,N_6808);
nand U7445 (N_7445,N_6520,N_6995);
nand U7446 (N_7446,N_6803,N_6624);
xnor U7447 (N_7447,N_6880,N_6965);
nand U7448 (N_7448,N_6596,N_6532);
or U7449 (N_7449,N_6691,N_6815);
nor U7450 (N_7450,N_6723,N_6749);
nand U7451 (N_7451,N_6667,N_6655);
or U7452 (N_7452,N_6797,N_6592);
nor U7453 (N_7453,N_6759,N_6874);
nand U7454 (N_7454,N_6870,N_6727);
or U7455 (N_7455,N_6752,N_6730);
nor U7456 (N_7456,N_6826,N_6753);
nor U7457 (N_7457,N_6655,N_6700);
nand U7458 (N_7458,N_6977,N_6523);
nand U7459 (N_7459,N_6954,N_6744);
nand U7460 (N_7460,N_6526,N_6691);
or U7461 (N_7461,N_6657,N_6870);
or U7462 (N_7462,N_6719,N_6977);
and U7463 (N_7463,N_6816,N_6501);
nor U7464 (N_7464,N_6525,N_6901);
and U7465 (N_7465,N_6799,N_6813);
or U7466 (N_7466,N_6994,N_6768);
nor U7467 (N_7467,N_6782,N_6991);
and U7468 (N_7468,N_6772,N_6847);
nand U7469 (N_7469,N_6542,N_6937);
nand U7470 (N_7470,N_6788,N_6682);
nor U7471 (N_7471,N_6503,N_6979);
nor U7472 (N_7472,N_6593,N_6947);
nand U7473 (N_7473,N_6674,N_6749);
and U7474 (N_7474,N_6540,N_6635);
nor U7475 (N_7475,N_6886,N_6942);
and U7476 (N_7476,N_6958,N_6727);
nand U7477 (N_7477,N_6622,N_6673);
and U7478 (N_7478,N_6708,N_6697);
or U7479 (N_7479,N_6905,N_6980);
nand U7480 (N_7480,N_6811,N_6815);
or U7481 (N_7481,N_6871,N_6914);
nand U7482 (N_7482,N_6511,N_6512);
or U7483 (N_7483,N_6940,N_6530);
and U7484 (N_7484,N_6848,N_6611);
xnor U7485 (N_7485,N_6671,N_6748);
nor U7486 (N_7486,N_6964,N_6609);
xnor U7487 (N_7487,N_6558,N_6919);
and U7488 (N_7488,N_6664,N_6627);
and U7489 (N_7489,N_6839,N_6886);
and U7490 (N_7490,N_6875,N_6910);
nand U7491 (N_7491,N_6917,N_6992);
nor U7492 (N_7492,N_6990,N_6642);
and U7493 (N_7493,N_6749,N_6505);
nor U7494 (N_7494,N_6929,N_6752);
nor U7495 (N_7495,N_6650,N_6606);
and U7496 (N_7496,N_6503,N_6835);
or U7497 (N_7497,N_6546,N_6643);
nor U7498 (N_7498,N_6635,N_6934);
or U7499 (N_7499,N_6533,N_6892);
or U7500 (N_7500,N_7108,N_7476);
or U7501 (N_7501,N_7171,N_7184);
or U7502 (N_7502,N_7407,N_7446);
xor U7503 (N_7503,N_7450,N_7136);
nand U7504 (N_7504,N_7102,N_7097);
or U7505 (N_7505,N_7137,N_7332);
nor U7506 (N_7506,N_7339,N_7485);
or U7507 (N_7507,N_7319,N_7314);
or U7508 (N_7508,N_7422,N_7261);
nand U7509 (N_7509,N_7372,N_7111);
and U7510 (N_7510,N_7281,N_7439);
nand U7511 (N_7511,N_7441,N_7321);
and U7512 (N_7512,N_7239,N_7061);
xnor U7513 (N_7513,N_7438,N_7241);
xor U7514 (N_7514,N_7382,N_7127);
and U7515 (N_7515,N_7164,N_7178);
and U7516 (N_7516,N_7435,N_7258);
nor U7517 (N_7517,N_7363,N_7226);
nor U7518 (N_7518,N_7249,N_7436);
and U7519 (N_7519,N_7140,N_7324);
or U7520 (N_7520,N_7199,N_7274);
or U7521 (N_7521,N_7381,N_7311);
and U7522 (N_7522,N_7055,N_7014);
nand U7523 (N_7523,N_7189,N_7267);
or U7524 (N_7524,N_7029,N_7046);
nor U7525 (N_7525,N_7196,N_7303);
nand U7526 (N_7526,N_7027,N_7473);
nand U7527 (N_7527,N_7343,N_7338);
nand U7528 (N_7528,N_7325,N_7491);
nor U7529 (N_7529,N_7119,N_7298);
and U7530 (N_7530,N_7038,N_7074);
xor U7531 (N_7531,N_7379,N_7421);
nand U7532 (N_7532,N_7086,N_7403);
nand U7533 (N_7533,N_7283,N_7291);
xor U7534 (N_7534,N_7366,N_7447);
nand U7535 (N_7535,N_7304,N_7415);
and U7536 (N_7536,N_7279,N_7115);
and U7537 (N_7537,N_7285,N_7188);
or U7538 (N_7538,N_7277,N_7440);
nand U7539 (N_7539,N_7091,N_7075);
and U7540 (N_7540,N_7329,N_7100);
nand U7541 (N_7541,N_7047,N_7272);
nand U7542 (N_7542,N_7158,N_7208);
nand U7543 (N_7543,N_7488,N_7008);
nor U7544 (N_7544,N_7357,N_7497);
and U7545 (N_7545,N_7054,N_7423);
xor U7546 (N_7546,N_7201,N_7263);
and U7547 (N_7547,N_7033,N_7180);
nand U7548 (N_7548,N_7289,N_7224);
or U7549 (N_7549,N_7093,N_7345);
nand U7550 (N_7550,N_7065,N_7044);
nand U7551 (N_7551,N_7235,N_7242);
nor U7552 (N_7552,N_7082,N_7323);
nor U7553 (N_7553,N_7313,N_7073);
nand U7554 (N_7554,N_7103,N_7430);
nor U7555 (N_7555,N_7286,N_7020);
and U7556 (N_7556,N_7309,N_7395);
nor U7557 (N_7557,N_7089,N_7149);
or U7558 (N_7558,N_7499,N_7072);
xnor U7559 (N_7559,N_7255,N_7348);
nand U7560 (N_7560,N_7223,N_7482);
nor U7561 (N_7561,N_7378,N_7232);
or U7562 (N_7562,N_7092,N_7260);
and U7563 (N_7563,N_7409,N_7009);
and U7564 (N_7564,N_7132,N_7269);
or U7565 (N_7565,N_7390,N_7138);
and U7566 (N_7566,N_7320,N_7041);
xnor U7567 (N_7567,N_7448,N_7204);
and U7568 (N_7568,N_7206,N_7344);
or U7569 (N_7569,N_7244,N_7191);
and U7570 (N_7570,N_7371,N_7248);
nand U7571 (N_7571,N_7406,N_7386);
nor U7572 (N_7572,N_7337,N_7259);
xnor U7573 (N_7573,N_7016,N_7211);
nor U7574 (N_7574,N_7152,N_7193);
nor U7575 (N_7575,N_7404,N_7150);
nand U7576 (N_7576,N_7394,N_7233);
nor U7577 (N_7577,N_7063,N_7183);
xnor U7578 (N_7578,N_7359,N_7481);
nor U7579 (N_7579,N_7017,N_7296);
and U7580 (N_7580,N_7351,N_7433);
xnor U7581 (N_7581,N_7388,N_7442);
or U7582 (N_7582,N_7494,N_7013);
and U7583 (N_7583,N_7402,N_7058);
nand U7584 (N_7584,N_7018,N_7419);
and U7585 (N_7585,N_7276,N_7453);
xnor U7586 (N_7586,N_7460,N_7498);
xnor U7587 (N_7587,N_7159,N_7397);
nand U7588 (N_7588,N_7399,N_7437);
or U7589 (N_7589,N_7443,N_7088);
and U7590 (N_7590,N_7462,N_7090);
or U7591 (N_7591,N_7236,N_7492);
or U7592 (N_7592,N_7374,N_7167);
or U7593 (N_7593,N_7221,N_7053);
nand U7594 (N_7594,N_7213,N_7237);
and U7595 (N_7595,N_7310,N_7445);
and U7596 (N_7596,N_7290,N_7114);
nand U7597 (N_7597,N_7326,N_7318);
and U7598 (N_7598,N_7257,N_7084);
nor U7599 (N_7599,N_7212,N_7000);
nor U7600 (N_7600,N_7078,N_7170);
or U7601 (N_7601,N_7389,N_7095);
nand U7602 (N_7602,N_7243,N_7302);
or U7603 (N_7603,N_7355,N_7262);
nand U7604 (N_7604,N_7360,N_7141);
nand U7605 (N_7605,N_7225,N_7124);
or U7606 (N_7606,N_7026,N_7240);
nor U7607 (N_7607,N_7327,N_7393);
or U7608 (N_7608,N_7021,N_7064);
xnor U7609 (N_7609,N_7375,N_7197);
and U7610 (N_7610,N_7117,N_7181);
and U7611 (N_7611,N_7340,N_7098);
or U7612 (N_7612,N_7135,N_7068);
nand U7613 (N_7613,N_7271,N_7299);
xor U7614 (N_7614,N_7315,N_7069);
nor U7615 (N_7615,N_7459,N_7007);
nor U7616 (N_7616,N_7347,N_7198);
nand U7617 (N_7617,N_7405,N_7294);
nand U7618 (N_7618,N_7330,N_7342);
nand U7619 (N_7619,N_7010,N_7083);
nand U7620 (N_7620,N_7173,N_7416);
nor U7621 (N_7621,N_7282,N_7101);
nand U7622 (N_7622,N_7216,N_7028);
xor U7623 (N_7623,N_7067,N_7085);
xor U7624 (N_7624,N_7050,N_7169);
or U7625 (N_7625,N_7478,N_7287);
and U7626 (N_7626,N_7032,N_7376);
nor U7627 (N_7627,N_7349,N_7365);
xnor U7628 (N_7628,N_7218,N_7024);
or U7629 (N_7629,N_7219,N_7099);
nor U7630 (N_7630,N_7128,N_7396);
or U7631 (N_7631,N_7011,N_7106);
or U7632 (N_7632,N_7229,N_7077);
or U7633 (N_7633,N_7306,N_7005);
nand U7634 (N_7634,N_7368,N_7134);
nand U7635 (N_7635,N_7387,N_7036);
or U7636 (N_7636,N_7483,N_7121);
or U7637 (N_7637,N_7070,N_7040);
nand U7638 (N_7638,N_7043,N_7454);
nor U7639 (N_7639,N_7495,N_7252);
or U7640 (N_7640,N_7080,N_7250);
and U7641 (N_7641,N_7457,N_7364);
nor U7642 (N_7642,N_7151,N_7391);
nand U7643 (N_7643,N_7493,N_7003);
or U7644 (N_7644,N_7015,N_7230);
xor U7645 (N_7645,N_7185,N_7350);
and U7646 (N_7646,N_7163,N_7479);
or U7647 (N_7647,N_7060,N_7203);
nand U7648 (N_7648,N_7358,N_7166);
or U7649 (N_7649,N_7175,N_7194);
nor U7650 (N_7650,N_7165,N_7207);
xnor U7651 (N_7651,N_7465,N_7186);
nand U7652 (N_7652,N_7179,N_7214);
nand U7653 (N_7653,N_7256,N_7023);
and U7654 (N_7654,N_7297,N_7292);
nor U7655 (N_7655,N_7035,N_7145);
and U7656 (N_7656,N_7467,N_7490);
and U7657 (N_7657,N_7056,N_7477);
nand U7658 (N_7658,N_7426,N_7126);
nand U7659 (N_7659,N_7489,N_7210);
or U7660 (N_7660,N_7107,N_7113);
nor U7661 (N_7661,N_7420,N_7238);
nor U7662 (N_7662,N_7373,N_7227);
nor U7663 (N_7663,N_7001,N_7187);
or U7664 (N_7664,N_7428,N_7112);
nor U7665 (N_7665,N_7051,N_7475);
nor U7666 (N_7666,N_7336,N_7066);
or U7667 (N_7667,N_7270,N_7461);
and U7668 (N_7668,N_7059,N_7417);
or U7669 (N_7669,N_7247,N_7300);
nand U7670 (N_7670,N_7392,N_7307);
and U7671 (N_7671,N_7168,N_7174);
or U7672 (N_7672,N_7317,N_7451);
nand U7673 (N_7673,N_7265,N_7254);
and U7674 (N_7674,N_7153,N_7192);
and U7675 (N_7675,N_7412,N_7228);
nor U7676 (N_7676,N_7331,N_7400);
nor U7677 (N_7677,N_7105,N_7120);
nor U7678 (N_7678,N_7104,N_7177);
and U7679 (N_7679,N_7215,N_7157);
nand U7680 (N_7680,N_7195,N_7470);
and U7681 (N_7681,N_7432,N_7352);
nand U7682 (N_7682,N_7251,N_7316);
nor U7683 (N_7683,N_7253,N_7039);
nor U7684 (N_7684,N_7062,N_7346);
nor U7685 (N_7685,N_7284,N_7472);
or U7686 (N_7686,N_7231,N_7334);
or U7687 (N_7687,N_7096,N_7322);
nand U7688 (N_7688,N_7487,N_7305);
nand U7689 (N_7689,N_7424,N_7019);
or U7690 (N_7690,N_7071,N_7474);
nor U7691 (N_7691,N_7484,N_7369);
nand U7692 (N_7692,N_7037,N_7385);
nor U7693 (N_7693,N_7148,N_7384);
or U7694 (N_7694,N_7048,N_7414);
and U7695 (N_7695,N_7246,N_7429);
xor U7696 (N_7696,N_7413,N_7308);
and U7697 (N_7697,N_7133,N_7129);
xor U7698 (N_7698,N_7456,N_7245);
and U7699 (N_7699,N_7411,N_7278);
or U7700 (N_7700,N_7004,N_7370);
xnor U7701 (N_7701,N_7034,N_7418);
nand U7702 (N_7702,N_7463,N_7444);
nor U7703 (N_7703,N_7362,N_7202);
nand U7704 (N_7704,N_7471,N_7116);
or U7705 (N_7705,N_7110,N_7361);
or U7706 (N_7706,N_7079,N_7268);
xor U7707 (N_7707,N_7486,N_7052);
nand U7708 (N_7708,N_7002,N_7209);
nand U7709 (N_7709,N_7190,N_7030);
nor U7710 (N_7710,N_7354,N_7353);
or U7711 (N_7711,N_7333,N_7022);
nor U7712 (N_7712,N_7087,N_7118);
and U7713 (N_7713,N_7328,N_7234);
xor U7714 (N_7714,N_7042,N_7131);
and U7715 (N_7715,N_7081,N_7160);
or U7716 (N_7716,N_7162,N_7288);
xor U7717 (N_7717,N_7094,N_7458);
nor U7718 (N_7718,N_7220,N_7301);
nand U7719 (N_7719,N_7464,N_7449);
nand U7720 (N_7720,N_7155,N_7312);
nand U7721 (N_7721,N_7295,N_7356);
xnor U7722 (N_7722,N_7266,N_7434);
and U7723 (N_7723,N_7156,N_7455);
xnor U7724 (N_7724,N_7200,N_7142);
nor U7725 (N_7725,N_7264,N_7293);
and U7726 (N_7726,N_7144,N_7383);
nor U7727 (N_7727,N_7154,N_7139);
nand U7728 (N_7728,N_7161,N_7380);
and U7729 (N_7729,N_7049,N_7275);
and U7730 (N_7730,N_7410,N_7452);
and U7731 (N_7731,N_7401,N_7377);
and U7732 (N_7732,N_7045,N_7147);
nor U7733 (N_7733,N_7335,N_7176);
nor U7734 (N_7734,N_7496,N_7480);
or U7735 (N_7735,N_7076,N_7280);
nor U7736 (N_7736,N_7006,N_7431);
and U7737 (N_7737,N_7057,N_7398);
nand U7738 (N_7738,N_7109,N_7468);
nand U7739 (N_7739,N_7222,N_7408);
or U7740 (N_7740,N_7182,N_7012);
nand U7741 (N_7741,N_7367,N_7205);
nand U7742 (N_7742,N_7123,N_7341);
nand U7743 (N_7743,N_7469,N_7125);
nand U7744 (N_7744,N_7425,N_7172);
or U7745 (N_7745,N_7122,N_7130);
nor U7746 (N_7746,N_7427,N_7217);
nand U7747 (N_7747,N_7273,N_7143);
nand U7748 (N_7748,N_7146,N_7031);
or U7749 (N_7749,N_7025,N_7466);
or U7750 (N_7750,N_7468,N_7366);
and U7751 (N_7751,N_7035,N_7305);
nor U7752 (N_7752,N_7232,N_7475);
or U7753 (N_7753,N_7290,N_7436);
nor U7754 (N_7754,N_7465,N_7389);
or U7755 (N_7755,N_7224,N_7056);
or U7756 (N_7756,N_7337,N_7189);
or U7757 (N_7757,N_7422,N_7227);
nor U7758 (N_7758,N_7028,N_7086);
nand U7759 (N_7759,N_7348,N_7256);
nand U7760 (N_7760,N_7470,N_7220);
nor U7761 (N_7761,N_7222,N_7209);
xnor U7762 (N_7762,N_7322,N_7272);
and U7763 (N_7763,N_7340,N_7157);
nor U7764 (N_7764,N_7239,N_7060);
nand U7765 (N_7765,N_7412,N_7211);
nand U7766 (N_7766,N_7250,N_7414);
nand U7767 (N_7767,N_7063,N_7325);
or U7768 (N_7768,N_7039,N_7356);
nor U7769 (N_7769,N_7123,N_7209);
or U7770 (N_7770,N_7183,N_7326);
nor U7771 (N_7771,N_7470,N_7131);
and U7772 (N_7772,N_7055,N_7313);
nor U7773 (N_7773,N_7147,N_7268);
nor U7774 (N_7774,N_7205,N_7233);
or U7775 (N_7775,N_7172,N_7118);
and U7776 (N_7776,N_7086,N_7097);
or U7777 (N_7777,N_7121,N_7220);
xor U7778 (N_7778,N_7134,N_7352);
nor U7779 (N_7779,N_7356,N_7026);
xor U7780 (N_7780,N_7060,N_7197);
or U7781 (N_7781,N_7029,N_7092);
nor U7782 (N_7782,N_7275,N_7174);
xnor U7783 (N_7783,N_7448,N_7403);
and U7784 (N_7784,N_7466,N_7417);
or U7785 (N_7785,N_7180,N_7341);
or U7786 (N_7786,N_7254,N_7266);
or U7787 (N_7787,N_7277,N_7137);
nor U7788 (N_7788,N_7399,N_7290);
nor U7789 (N_7789,N_7129,N_7017);
nor U7790 (N_7790,N_7435,N_7492);
nor U7791 (N_7791,N_7123,N_7114);
or U7792 (N_7792,N_7190,N_7390);
nor U7793 (N_7793,N_7455,N_7116);
nor U7794 (N_7794,N_7188,N_7210);
nand U7795 (N_7795,N_7350,N_7091);
or U7796 (N_7796,N_7048,N_7371);
xnor U7797 (N_7797,N_7358,N_7313);
nand U7798 (N_7798,N_7361,N_7413);
nand U7799 (N_7799,N_7490,N_7356);
or U7800 (N_7800,N_7390,N_7360);
xnor U7801 (N_7801,N_7182,N_7128);
and U7802 (N_7802,N_7023,N_7161);
and U7803 (N_7803,N_7144,N_7220);
xnor U7804 (N_7804,N_7328,N_7434);
and U7805 (N_7805,N_7074,N_7403);
or U7806 (N_7806,N_7113,N_7062);
or U7807 (N_7807,N_7428,N_7076);
nor U7808 (N_7808,N_7360,N_7447);
nand U7809 (N_7809,N_7029,N_7194);
nand U7810 (N_7810,N_7451,N_7070);
xor U7811 (N_7811,N_7030,N_7444);
nor U7812 (N_7812,N_7340,N_7456);
and U7813 (N_7813,N_7371,N_7105);
nor U7814 (N_7814,N_7406,N_7191);
nor U7815 (N_7815,N_7463,N_7135);
nand U7816 (N_7816,N_7477,N_7427);
or U7817 (N_7817,N_7275,N_7267);
xnor U7818 (N_7818,N_7243,N_7359);
nand U7819 (N_7819,N_7022,N_7329);
or U7820 (N_7820,N_7017,N_7267);
xor U7821 (N_7821,N_7260,N_7211);
nor U7822 (N_7822,N_7063,N_7413);
or U7823 (N_7823,N_7297,N_7461);
nand U7824 (N_7824,N_7348,N_7097);
nor U7825 (N_7825,N_7045,N_7078);
xnor U7826 (N_7826,N_7457,N_7328);
nand U7827 (N_7827,N_7225,N_7100);
or U7828 (N_7828,N_7251,N_7320);
nor U7829 (N_7829,N_7283,N_7398);
nand U7830 (N_7830,N_7365,N_7056);
nor U7831 (N_7831,N_7378,N_7390);
nand U7832 (N_7832,N_7302,N_7085);
and U7833 (N_7833,N_7013,N_7426);
nor U7834 (N_7834,N_7369,N_7348);
nand U7835 (N_7835,N_7240,N_7406);
nor U7836 (N_7836,N_7174,N_7165);
nor U7837 (N_7837,N_7359,N_7103);
and U7838 (N_7838,N_7037,N_7417);
nor U7839 (N_7839,N_7464,N_7040);
nand U7840 (N_7840,N_7317,N_7152);
nand U7841 (N_7841,N_7474,N_7124);
nand U7842 (N_7842,N_7030,N_7109);
nand U7843 (N_7843,N_7380,N_7133);
or U7844 (N_7844,N_7068,N_7319);
or U7845 (N_7845,N_7070,N_7467);
xnor U7846 (N_7846,N_7104,N_7486);
or U7847 (N_7847,N_7086,N_7138);
nand U7848 (N_7848,N_7489,N_7174);
nor U7849 (N_7849,N_7226,N_7464);
and U7850 (N_7850,N_7088,N_7149);
or U7851 (N_7851,N_7271,N_7480);
and U7852 (N_7852,N_7369,N_7156);
and U7853 (N_7853,N_7372,N_7168);
and U7854 (N_7854,N_7232,N_7420);
and U7855 (N_7855,N_7423,N_7122);
nor U7856 (N_7856,N_7321,N_7032);
nand U7857 (N_7857,N_7029,N_7411);
and U7858 (N_7858,N_7334,N_7227);
and U7859 (N_7859,N_7293,N_7140);
xnor U7860 (N_7860,N_7239,N_7230);
or U7861 (N_7861,N_7350,N_7157);
nor U7862 (N_7862,N_7439,N_7074);
xor U7863 (N_7863,N_7173,N_7427);
and U7864 (N_7864,N_7492,N_7464);
and U7865 (N_7865,N_7423,N_7155);
xnor U7866 (N_7866,N_7145,N_7089);
and U7867 (N_7867,N_7149,N_7061);
and U7868 (N_7868,N_7074,N_7333);
nor U7869 (N_7869,N_7117,N_7402);
or U7870 (N_7870,N_7051,N_7373);
or U7871 (N_7871,N_7294,N_7345);
nor U7872 (N_7872,N_7466,N_7278);
or U7873 (N_7873,N_7274,N_7248);
and U7874 (N_7874,N_7292,N_7134);
and U7875 (N_7875,N_7352,N_7064);
and U7876 (N_7876,N_7380,N_7353);
or U7877 (N_7877,N_7133,N_7461);
nor U7878 (N_7878,N_7426,N_7452);
nand U7879 (N_7879,N_7112,N_7047);
or U7880 (N_7880,N_7009,N_7172);
and U7881 (N_7881,N_7181,N_7299);
or U7882 (N_7882,N_7198,N_7284);
nand U7883 (N_7883,N_7097,N_7030);
or U7884 (N_7884,N_7014,N_7421);
and U7885 (N_7885,N_7432,N_7215);
nor U7886 (N_7886,N_7198,N_7449);
or U7887 (N_7887,N_7057,N_7029);
nand U7888 (N_7888,N_7057,N_7148);
nor U7889 (N_7889,N_7329,N_7499);
nor U7890 (N_7890,N_7355,N_7271);
or U7891 (N_7891,N_7119,N_7343);
and U7892 (N_7892,N_7078,N_7003);
and U7893 (N_7893,N_7153,N_7228);
nand U7894 (N_7894,N_7397,N_7065);
nand U7895 (N_7895,N_7248,N_7486);
nor U7896 (N_7896,N_7242,N_7069);
or U7897 (N_7897,N_7084,N_7337);
nand U7898 (N_7898,N_7096,N_7210);
and U7899 (N_7899,N_7498,N_7312);
and U7900 (N_7900,N_7290,N_7025);
and U7901 (N_7901,N_7312,N_7238);
and U7902 (N_7902,N_7267,N_7090);
or U7903 (N_7903,N_7086,N_7301);
nand U7904 (N_7904,N_7072,N_7276);
nand U7905 (N_7905,N_7256,N_7307);
nor U7906 (N_7906,N_7312,N_7288);
or U7907 (N_7907,N_7394,N_7260);
and U7908 (N_7908,N_7417,N_7027);
and U7909 (N_7909,N_7353,N_7288);
or U7910 (N_7910,N_7407,N_7359);
nor U7911 (N_7911,N_7294,N_7234);
nand U7912 (N_7912,N_7101,N_7458);
nand U7913 (N_7913,N_7451,N_7117);
nand U7914 (N_7914,N_7419,N_7327);
and U7915 (N_7915,N_7274,N_7431);
or U7916 (N_7916,N_7387,N_7245);
nand U7917 (N_7917,N_7464,N_7079);
nor U7918 (N_7918,N_7452,N_7106);
or U7919 (N_7919,N_7447,N_7333);
or U7920 (N_7920,N_7473,N_7433);
nand U7921 (N_7921,N_7175,N_7323);
and U7922 (N_7922,N_7211,N_7478);
nand U7923 (N_7923,N_7138,N_7495);
nor U7924 (N_7924,N_7074,N_7285);
nor U7925 (N_7925,N_7029,N_7258);
nand U7926 (N_7926,N_7048,N_7470);
nor U7927 (N_7927,N_7138,N_7267);
or U7928 (N_7928,N_7387,N_7364);
and U7929 (N_7929,N_7064,N_7136);
and U7930 (N_7930,N_7024,N_7313);
and U7931 (N_7931,N_7027,N_7085);
or U7932 (N_7932,N_7268,N_7254);
nand U7933 (N_7933,N_7038,N_7397);
nor U7934 (N_7934,N_7104,N_7455);
and U7935 (N_7935,N_7415,N_7474);
nor U7936 (N_7936,N_7063,N_7313);
nor U7937 (N_7937,N_7474,N_7309);
and U7938 (N_7938,N_7457,N_7275);
nand U7939 (N_7939,N_7096,N_7146);
nand U7940 (N_7940,N_7340,N_7291);
and U7941 (N_7941,N_7396,N_7397);
nor U7942 (N_7942,N_7004,N_7176);
and U7943 (N_7943,N_7118,N_7109);
xnor U7944 (N_7944,N_7167,N_7008);
and U7945 (N_7945,N_7092,N_7171);
and U7946 (N_7946,N_7243,N_7405);
nand U7947 (N_7947,N_7139,N_7028);
nand U7948 (N_7948,N_7184,N_7135);
nand U7949 (N_7949,N_7100,N_7497);
nand U7950 (N_7950,N_7419,N_7415);
or U7951 (N_7951,N_7424,N_7037);
nand U7952 (N_7952,N_7030,N_7027);
nand U7953 (N_7953,N_7339,N_7011);
nor U7954 (N_7954,N_7255,N_7455);
or U7955 (N_7955,N_7096,N_7052);
and U7956 (N_7956,N_7044,N_7299);
nor U7957 (N_7957,N_7141,N_7498);
and U7958 (N_7958,N_7082,N_7227);
xnor U7959 (N_7959,N_7020,N_7089);
nor U7960 (N_7960,N_7114,N_7098);
nor U7961 (N_7961,N_7326,N_7154);
nor U7962 (N_7962,N_7370,N_7312);
or U7963 (N_7963,N_7156,N_7319);
and U7964 (N_7964,N_7441,N_7175);
nand U7965 (N_7965,N_7245,N_7408);
nand U7966 (N_7966,N_7206,N_7350);
or U7967 (N_7967,N_7352,N_7268);
nor U7968 (N_7968,N_7327,N_7126);
nand U7969 (N_7969,N_7027,N_7013);
or U7970 (N_7970,N_7438,N_7154);
nor U7971 (N_7971,N_7499,N_7140);
or U7972 (N_7972,N_7131,N_7337);
nand U7973 (N_7973,N_7108,N_7330);
and U7974 (N_7974,N_7150,N_7425);
or U7975 (N_7975,N_7450,N_7351);
nor U7976 (N_7976,N_7313,N_7462);
and U7977 (N_7977,N_7028,N_7118);
nand U7978 (N_7978,N_7024,N_7427);
nor U7979 (N_7979,N_7415,N_7392);
nand U7980 (N_7980,N_7189,N_7116);
xnor U7981 (N_7981,N_7046,N_7370);
nor U7982 (N_7982,N_7230,N_7212);
nor U7983 (N_7983,N_7415,N_7173);
nand U7984 (N_7984,N_7367,N_7485);
nor U7985 (N_7985,N_7211,N_7415);
nand U7986 (N_7986,N_7268,N_7014);
or U7987 (N_7987,N_7400,N_7024);
nor U7988 (N_7988,N_7459,N_7036);
nor U7989 (N_7989,N_7173,N_7294);
xor U7990 (N_7990,N_7245,N_7125);
and U7991 (N_7991,N_7230,N_7351);
or U7992 (N_7992,N_7211,N_7039);
nor U7993 (N_7993,N_7482,N_7232);
nand U7994 (N_7994,N_7125,N_7360);
nand U7995 (N_7995,N_7091,N_7464);
xnor U7996 (N_7996,N_7147,N_7430);
or U7997 (N_7997,N_7102,N_7098);
nand U7998 (N_7998,N_7407,N_7189);
and U7999 (N_7999,N_7116,N_7064);
and U8000 (N_8000,N_7856,N_7541);
nand U8001 (N_8001,N_7651,N_7535);
nand U8002 (N_8002,N_7666,N_7654);
nand U8003 (N_8003,N_7890,N_7515);
nand U8004 (N_8004,N_7616,N_7552);
nor U8005 (N_8005,N_7915,N_7544);
and U8006 (N_8006,N_7585,N_7975);
nand U8007 (N_8007,N_7923,N_7985);
and U8008 (N_8008,N_7634,N_7600);
and U8009 (N_8009,N_7935,N_7982);
nor U8010 (N_8010,N_7657,N_7559);
or U8011 (N_8011,N_7653,N_7927);
nor U8012 (N_8012,N_7944,N_7547);
nor U8013 (N_8013,N_7939,N_7715);
or U8014 (N_8014,N_7551,N_7700);
and U8015 (N_8015,N_7797,N_7534);
nor U8016 (N_8016,N_7695,N_7542);
or U8017 (N_8017,N_7898,N_7553);
and U8018 (N_8018,N_7546,N_7829);
or U8019 (N_8019,N_7902,N_7726);
and U8020 (N_8020,N_7740,N_7998);
xor U8021 (N_8021,N_7967,N_7989);
nand U8022 (N_8022,N_7825,N_7721);
xor U8023 (N_8023,N_7576,N_7816);
and U8024 (N_8024,N_7995,N_7852);
or U8025 (N_8025,N_7684,N_7963);
nand U8026 (N_8026,N_7604,N_7947);
nand U8027 (N_8027,N_7808,N_7523);
or U8028 (N_8028,N_7500,N_7630);
and U8029 (N_8029,N_7512,N_7637);
and U8030 (N_8030,N_7997,N_7789);
and U8031 (N_8031,N_7878,N_7979);
nand U8032 (N_8032,N_7801,N_7660);
or U8033 (N_8033,N_7619,N_7556);
or U8034 (N_8034,N_7966,N_7781);
nor U8035 (N_8035,N_7577,N_7744);
and U8036 (N_8036,N_7569,N_7603);
nand U8037 (N_8037,N_7844,N_7804);
or U8038 (N_8038,N_7530,N_7655);
nor U8039 (N_8039,N_7873,N_7921);
and U8040 (N_8040,N_7893,N_7924);
or U8041 (N_8041,N_7988,N_7835);
and U8042 (N_8042,N_7599,N_7999);
xnor U8043 (N_8043,N_7882,N_7709);
nand U8044 (N_8044,N_7784,N_7658);
nand U8045 (N_8045,N_7888,N_7994);
and U8046 (N_8046,N_7627,N_7767);
nand U8047 (N_8047,N_7519,N_7503);
and U8048 (N_8048,N_7708,N_7764);
nand U8049 (N_8049,N_7734,N_7815);
nand U8050 (N_8050,N_7613,N_7570);
or U8051 (N_8051,N_7987,N_7800);
nand U8052 (N_8052,N_7824,N_7719);
nor U8053 (N_8053,N_7769,N_7615);
or U8054 (N_8054,N_7580,N_7645);
or U8055 (N_8055,N_7869,N_7795);
nor U8056 (N_8056,N_7957,N_7531);
nor U8057 (N_8057,N_7620,N_7920);
and U8058 (N_8058,N_7959,N_7713);
nand U8059 (N_8059,N_7518,N_7526);
nand U8060 (N_8060,N_7954,N_7656);
or U8061 (N_8061,N_7861,N_7639);
nor U8062 (N_8062,N_7511,N_7647);
nor U8063 (N_8063,N_7509,N_7748);
or U8064 (N_8064,N_7680,N_7943);
nand U8065 (N_8065,N_7848,N_7859);
and U8066 (N_8066,N_7590,N_7710);
nor U8067 (N_8067,N_7933,N_7607);
nor U8068 (N_8068,N_7635,N_7814);
xor U8069 (N_8069,N_7976,N_7786);
nand U8070 (N_8070,N_7909,N_7931);
nor U8071 (N_8071,N_7955,N_7727);
and U8072 (N_8072,N_7778,N_7894);
or U8073 (N_8073,N_7672,N_7840);
nor U8074 (N_8074,N_7817,N_7881);
nor U8075 (N_8075,N_7953,N_7971);
and U8076 (N_8076,N_7775,N_7728);
nor U8077 (N_8077,N_7807,N_7851);
or U8078 (N_8078,N_7904,N_7831);
nand U8079 (N_8079,N_7993,N_7629);
xor U8080 (N_8080,N_7794,N_7557);
or U8081 (N_8081,N_7846,N_7914);
and U8082 (N_8082,N_7796,N_7691);
nand U8083 (N_8083,N_7750,N_7618);
or U8084 (N_8084,N_7793,N_7932);
nor U8085 (N_8085,N_7593,N_7855);
or U8086 (N_8086,N_7688,N_7818);
nand U8087 (N_8087,N_7950,N_7761);
xnor U8088 (N_8088,N_7689,N_7510);
and U8089 (N_8089,N_7520,N_7641);
nor U8090 (N_8090,N_7929,N_7741);
nor U8091 (N_8091,N_7858,N_7925);
and U8092 (N_8092,N_7896,N_7571);
nand U8093 (N_8093,N_7774,N_7981);
nor U8094 (N_8094,N_7686,N_7663);
and U8095 (N_8095,N_7949,N_7501);
nand U8096 (N_8096,N_7903,N_7812);
or U8097 (N_8097,N_7757,N_7575);
nand U8098 (N_8098,N_7974,N_7675);
and U8099 (N_8099,N_7529,N_7780);
nor U8100 (N_8100,N_7847,N_7810);
or U8101 (N_8101,N_7703,N_7811);
or U8102 (N_8102,N_7598,N_7659);
and U8103 (N_8103,N_7839,N_7648);
and U8104 (N_8104,N_7564,N_7737);
xnor U8105 (N_8105,N_7681,N_7842);
nor U8106 (N_8106,N_7792,N_7673);
xor U8107 (N_8107,N_7883,N_7752);
xnor U8108 (N_8108,N_7961,N_7617);
or U8109 (N_8109,N_7555,N_7865);
and U8110 (N_8110,N_7813,N_7502);
nand U8111 (N_8111,N_7956,N_7732);
or U8112 (N_8112,N_7513,N_7828);
or U8113 (N_8113,N_7632,N_7517);
xor U8114 (N_8114,N_7803,N_7870);
nor U8115 (N_8115,N_7886,N_7910);
and U8116 (N_8116,N_7561,N_7572);
xor U8117 (N_8117,N_7631,N_7578);
or U8118 (N_8118,N_7574,N_7650);
nor U8119 (N_8119,N_7595,N_7738);
and U8120 (N_8120,N_7643,N_7678);
nor U8121 (N_8121,N_7514,N_7908);
nand U8122 (N_8122,N_7906,N_7749);
nor U8123 (N_8123,N_7567,N_7679);
xor U8124 (N_8124,N_7755,N_7687);
nor U8125 (N_8125,N_7917,N_7996);
or U8126 (N_8126,N_7505,N_7601);
nor U8127 (N_8127,N_7885,N_7760);
and U8128 (N_8128,N_7730,N_7916);
nor U8129 (N_8129,N_7614,N_7692);
nor U8130 (N_8130,N_7834,N_7562);
nor U8131 (N_8131,N_7753,N_7984);
and U8132 (N_8132,N_7581,N_7849);
nor U8133 (N_8133,N_7887,N_7897);
nand U8134 (N_8134,N_7969,N_7965);
and U8135 (N_8135,N_7573,N_7694);
nor U8136 (N_8136,N_7591,N_7621);
and U8137 (N_8137,N_7698,N_7946);
xor U8138 (N_8138,N_7725,N_7763);
xor U8139 (N_8139,N_7964,N_7986);
nand U8140 (N_8140,N_7714,N_7638);
nor U8141 (N_8141,N_7941,N_7758);
nor U8142 (N_8142,N_7992,N_7702);
nand U8143 (N_8143,N_7745,N_7754);
or U8144 (N_8144,N_7693,N_7733);
or U8145 (N_8145,N_7522,N_7788);
nand U8146 (N_8146,N_7646,N_7504);
nand U8147 (N_8147,N_7674,N_7587);
and U8148 (N_8148,N_7830,N_7685);
or U8149 (N_8149,N_7868,N_7864);
xnor U8150 (N_8150,N_7838,N_7605);
and U8151 (N_8151,N_7610,N_7798);
nor U8152 (N_8152,N_7696,N_7594);
xnor U8153 (N_8153,N_7945,N_7787);
nand U8154 (N_8154,N_7905,N_7528);
xnor U8155 (N_8155,N_7899,N_7867);
and U8156 (N_8156,N_7857,N_7771);
or U8157 (N_8157,N_7554,N_7579);
and U8158 (N_8158,N_7805,N_7806);
nand U8159 (N_8159,N_7712,N_7922);
nand U8160 (N_8160,N_7866,N_7589);
or U8161 (N_8161,N_7563,N_7705);
and U8162 (N_8162,N_7742,N_7799);
nor U8163 (N_8163,N_7623,N_7706);
nor U8164 (N_8164,N_7588,N_7913);
or U8165 (N_8165,N_7958,N_7662);
or U8166 (N_8166,N_7543,N_7900);
xnor U8167 (N_8167,N_7624,N_7602);
or U8168 (N_8168,N_7583,N_7586);
nand U8169 (N_8169,N_7550,N_7871);
and U8170 (N_8170,N_7676,N_7652);
nand U8171 (N_8171,N_7918,N_7756);
nor U8172 (N_8172,N_7677,N_7746);
and U8173 (N_8173,N_7565,N_7644);
or U8174 (N_8174,N_7545,N_7827);
nand U8175 (N_8175,N_7862,N_7895);
and U8176 (N_8176,N_7891,N_7991);
and U8177 (N_8177,N_7980,N_7736);
or U8178 (N_8178,N_7962,N_7960);
or U8179 (N_8179,N_7791,N_7699);
nand U8180 (N_8180,N_7779,N_7951);
nor U8181 (N_8181,N_7837,N_7875);
nor U8182 (N_8182,N_7854,N_7717);
nor U8183 (N_8183,N_7983,N_7880);
nor U8184 (N_8184,N_7516,N_7649);
nor U8185 (N_8185,N_7720,N_7919);
xnor U8186 (N_8186,N_7845,N_7671);
nor U8187 (N_8187,N_7524,N_7582);
nand U8188 (N_8188,N_7661,N_7665);
or U8189 (N_8189,N_7597,N_7821);
xnor U8190 (N_8190,N_7622,N_7836);
nand U8191 (N_8191,N_7701,N_7822);
nand U8192 (N_8192,N_7716,N_7697);
or U8193 (N_8193,N_7747,N_7860);
nor U8194 (N_8194,N_7762,N_7823);
nand U8195 (N_8195,N_7608,N_7548);
nand U8196 (N_8196,N_7783,N_7832);
nor U8197 (N_8197,N_7934,N_7874);
nand U8198 (N_8198,N_7843,N_7772);
nor U8199 (N_8199,N_7876,N_7536);
nand U8200 (N_8200,N_7759,N_7735);
xor U8201 (N_8201,N_7636,N_7668);
or U8202 (N_8202,N_7633,N_7612);
xor U8203 (N_8203,N_7642,N_7626);
nand U8204 (N_8204,N_7972,N_7532);
nand U8205 (N_8205,N_7533,N_7889);
and U8206 (N_8206,N_7977,N_7592);
and U8207 (N_8207,N_7667,N_7973);
nor U8208 (N_8208,N_7521,N_7729);
nor U8209 (N_8209,N_7948,N_7930);
and U8210 (N_8210,N_7768,N_7751);
nor U8211 (N_8211,N_7877,N_7863);
nand U8212 (N_8212,N_7926,N_7940);
nand U8213 (N_8213,N_7952,N_7978);
nor U8214 (N_8214,N_7892,N_7928);
or U8215 (N_8215,N_7879,N_7820);
nand U8216 (N_8216,N_7724,N_7539);
nand U8217 (N_8217,N_7942,N_7777);
or U8218 (N_8218,N_7682,N_7549);
and U8219 (N_8219,N_7731,N_7765);
nor U8220 (N_8220,N_7850,N_7790);
or U8221 (N_8221,N_7826,N_7776);
and U8222 (N_8222,N_7707,N_7782);
nor U8223 (N_8223,N_7872,N_7884);
and U8224 (N_8224,N_7901,N_7664);
and U8225 (N_8225,N_7584,N_7937);
nand U8226 (N_8226,N_7773,N_7938);
or U8227 (N_8227,N_7525,N_7640);
nor U8228 (N_8228,N_7690,N_7833);
nor U8229 (N_8229,N_7506,N_7560);
nand U8230 (N_8230,N_7670,N_7558);
and U8231 (N_8231,N_7508,N_7596);
nand U8232 (N_8232,N_7853,N_7718);
nor U8233 (N_8233,N_7907,N_7936);
and U8234 (N_8234,N_7609,N_7568);
nor U8235 (N_8235,N_7990,N_7770);
nor U8236 (N_8236,N_7970,N_7912);
xor U8237 (N_8237,N_7711,N_7628);
or U8238 (N_8238,N_7723,N_7802);
or U8239 (N_8239,N_7527,N_7739);
and U8240 (N_8240,N_7538,N_7683);
xor U8241 (N_8241,N_7606,N_7743);
nand U8242 (N_8242,N_7785,N_7809);
xor U8243 (N_8243,N_7537,N_7540);
and U8244 (N_8244,N_7704,N_7507);
and U8245 (N_8245,N_7625,N_7611);
and U8246 (N_8246,N_7911,N_7669);
and U8247 (N_8247,N_7722,N_7968);
nand U8248 (N_8248,N_7566,N_7819);
nand U8249 (N_8249,N_7766,N_7841);
xor U8250 (N_8250,N_7548,N_7773);
nor U8251 (N_8251,N_7929,N_7996);
or U8252 (N_8252,N_7642,N_7781);
nand U8253 (N_8253,N_7581,N_7830);
nand U8254 (N_8254,N_7688,N_7648);
or U8255 (N_8255,N_7711,N_7674);
and U8256 (N_8256,N_7805,N_7526);
and U8257 (N_8257,N_7530,N_7831);
and U8258 (N_8258,N_7919,N_7976);
or U8259 (N_8259,N_7677,N_7959);
and U8260 (N_8260,N_7988,N_7778);
nand U8261 (N_8261,N_7980,N_7526);
or U8262 (N_8262,N_7859,N_7988);
and U8263 (N_8263,N_7709,N_7528);
or U8264 (N_8264,N_7698,N_7738);
and U8265 (N_8265,N_7947,N_7939);
xor U8266 (N_8266,N_7803,N_7819);
nor U8267 (N_8267,N_7524,N_7622);
xnor U8268 (N_8268,N_7866,N_7786);
nand U8269 (N_8269,N_7727,N_7645);
nand U8270 (N_8270,N_7567,N_7624);
nand U8271 (N_8271,N_7510,N_7513);
and U8272 (N_8272,N_7676,N_7927);
or U8273 (N_8273,N_7765,N_7790);
and U8274 (N_8274,N_7529,N_7704);
xnor U8275 (N_8275,N_7515,N_7704);
nor U8276 (N_8276,N_7928,N_7505);
nand U8277 (N_8277,N_7755,N_7721);
nand U8278 (N_8278,N_7753,N_7641);
nor U8279 (N_8279,N_7983,N_7537);
and U8280 (N_8280,N_7843,N_7896);
or U8281 (N_8281,N_7567,N_7782);
xor U8282 (N_8282,N_7765,N_7916);
nor U8283 (N_8283,N_7986,N_7611);
or U8284 (N_8284,N_7524,N_7889);
nand U8285 (N_8285,N_7622,N_7719);
nor U8286 (N_8286,N_7782,N_7685);
nor U8287 (N_8287,N_7671,N_7842);
and U8288 (N_8288,N_7547,N_7740);
nor U8289 (N_8289,N_7714,N_7510);
and U8290 (N_8290,N_7954,N_7716);
xnor U8291 (N_8291,N_7948,N_7956);
xnor U8292 (N_8292,N_7991,N_7731);
nand U8293 (N_8293,N_7868,N_7928);
nand U8294 (N_8294,N_7956,N_7680);
or U8295 (N_8295,N_7839,N_7504);
nand U8296 (N_8296,N_7730,N_7851);
nand U8297 (N_8297,N_7852,N_7557);
nor U8298 (N_8298,N_7870,N_7706);
nor U8299 (N_8299,N_7763,N_7538);
nor U8300 (N_8300,N_7872,N_7714);
and U8301 (N_8301,N_7578,N_7962);
nand U8302 (N_8302,N_7531,N_7959);
or U8303 (N_8303,N_7835,N_7814);
nor U8304 (N_8304,N_7957,N_7578);
nor U8305 (N_8305,N_7900,N_7812);
or U8306 (N_8306,N_7696,N_7590);
xor U8307 (N_8307,N_7534,N_7807);
nor U8308 (N_8308,N_7991,N_7593);
and U8309 (N_8309,N_7693,N_7753);
nor U8310 (N_8310,N_7893,N_7841);
or U8311 (N_8311,N_7806,N_7692);
nor U8312 (N_8312,N_7883,N_7885);
and U8313 (N_8313,N_7732,N_7859);
xor U8314 (N_8314,N_7970,N_7835);
nor U8315 (N_8315,N_7591,N_7738);
or U8316 (N_8316,N_7938,N_7691);
and U8317 (N_8317,N_7649,N_7590);
or U8318 (N_8318,N_7882,N_7596);
nand U8319 (N_8319,N_7878,N_7634);
nor U8320 (N_8320,N_7650,N_7913);
nand U8321 (N_8321,N_7514,N_7782);
xor U8322 (N_8322,N_7570,N_7661);
nor U8323 (N_8323,N_7697,N_7511);
or U8324 (N_8324,N_7587,N_7889);
nand U8325 (N_8325,N_7728,N_7670);
nor U8326 (N_8326,N_7562,N_7522);
nor U8327 (N_8327,N_7909,N_7588);
nor U8328 (N_8328,N_7742,N_7854);
xor U8329 (N_8329,N_7689,N_7782);
or U8330 (N_8330,N_7951,N_7502);
and U8331 (N_8331,N_7639,N_7598);
nand U8332 (N_8332,N_7851,N_7582);
nand U8333 (N_8333,N_7635,N_7742);
or U8334 (N_8334,N_7588,N_7584);
xnor U8335 (N_8335,N_7800,N_7762);
and U8336 (N_8336,N_7997,N_7509);
and U8337 (N_8337,N_7618,N_7620);
and U8338 (N_8338,N_7588,N_7842);
and U8339 (N_8339,N_7900,N_7800);
nand U8340 (N_8340,N_7979,N_7989);
or U8341 (N_8341,N_7815,N_7771);
or U8342 (N_8342,N_7689,N_7595);
or U8343 (N_8343,N_7891,N_7736);
nand U8344 (N_8344,N_7816,N_7901);
or U8345 (N_8345,N_7870,N_7762);
nand U8346 (N_8346,N_7864,N_7928);
nand U8347 (N_8347,N_7739,N_7744);
nand U8348 (N_8348,N_7859,N_7685);
and U8349 (N_8349,N_7804,N_7509);
or U8350 (N_8350,N_7519,N_7550);
nor U8351 (N_8351,N_7775,N_7559);
or U8352 (N_8352,N_7800,N_7521);
and U8353 (N_8353,N_7509,N_7970);
nor U8354 (N_8354,N_7991,N_7652);
nor U8355 (N_8355,N_7813,N_7926);
nor U8356 (N_8356,N_7556,N_7949);
nand U8357 (N_8357,N_7854,N_7842);
nand U8358 (N_8358,N_7526,N_7851);
nand U8359 (N_8359,N_7873,N_7888);
nor U8360 (N_8360,N_7825,N_7749);
or U8361 (N_8361,N_7638,N_7502);
xor U8362 (N_8362,N_7646,N_7812);
nor U8363 (N_8363,N_7835,N_7686);
nand U8364 (N_8364,N_7762,N_7733);
or U8365 (N_8365,N_7650,N_7566);
nand U8366 (N_8366,N_7924,N_7921);
nor U8367 (N_8367,N_7858,N_7812);
nand U8368 (N_8368,N_7582,N_7680);
nand U8369 (N_8369,N_7896,N_7503);
nor U8370 (N_8370,N_7864,N_7555);
and U8371 (N_8371,N_7784,N_7712);
and U8372 (N_8372,N_7929,N_7820);
and U8373 (N_8373,N_7891,N_7669);
and U8374 (N_8374,N_7795,N_7604);
nor U8375 (N_8375,N_7759,N_7778);
and U8376 (N_8376,N_7699,N_7573);
or U8377 (N_8377,N_7826,N_7647);
or U8378 (N_8378,N_7533,N_7864);
or U8379 (N_8379,N_7876,N_7960);
xor U8380 (N_8380,N_7986,N_7837);
or U8381 (N_8381,N_7716,N_7624);
xnor U8382 (N_8382,N_7965,N_7720);
nor U8383 (N_8383,N_7958,N_7595);
and U8384 (N_8384,N_7723,N_7685);
or U8385 (N_8385,N_7566,N_7762);
and U8386 (N_8386,N_7867,N_7709);
xor U8387 (N_8387,N_7518,N_7994);
nor U8388 (N_8388,N_7550,N_7537);
nor U8389 (N_8389,N_7914,N_7998);
and U8390 (N_8390,N_7991,N_7864);
or U8391 (N_8391,N_7644,N_7743);
and U8392 (N_8392,N_7937,N_7908);
nand U8393 (N_8393,N_7608,N_7763);
nor U8394 (N_8394,N_7629,N_7842);
nor U8395 (N_8395,N_7622,N_7705);
nand U8396 (N_8396,N_7528,N_7771);
nand U8397 (N_8397,N_7871,N_7663);
nor U8398 (N_8398,N_7729,N_7768);
xor U8399 (N_8399,N_7861,N_7886);
and U8400 (N_8400,N_7974,N_7802);
xnor U8401 (N_8401,N_7539,N_7990);
and U8402 (N_8402,N_7580,N_7952);
xor U8403 (N_8403,N_7591,N_7759);
nor U8404 (N_8404,N_7817,N_7662);
or U8405 (N_8405,N_7806,N_7712);
nand U8406 (N_8406,N_7622,N_7538);
nand U8407 (N_8407,N_7833,N_7794);
and U8408 (N_8408,N_7759,N_7961);
nor U8409 (N_8409,N_7900,N_7860);
nand U8410 (N_8410,N_7919,N_7620);
nand U8411 (N_8411,N_7577,N_7513);
nand U8412 (N_8412,N_7576,N_7735);
nand U8413 (N_8413,N_7539,N_7663);
nor U8414 (N_8414,N_7816,N_7915);
nand U8415 (N_8415,N_7730,N_7833);
nor U8416 (N_8416,N_7720,N_7921);
and U8417 (N_8417,N_7732,N_7861);
nor U8418 (N_8418,N_7719,N_7697);
nor U8419 (N_8419,N_7535,N_7692);
nand U8420 (N_8420,N_7927,N_7784);
and U8421 (N_8421,N_7813,N_7671);
nor U8422 (N_8422,N_7895,N_7967);
and U8423 (N_8423,N_7987,N_7605);
or U8424 (N_8424,N_7781,N_7780);
and U8425 (N_8425,N_7600,N_7885);
or U8426 (N_8426,N_7607,N_7741);
or U8427 (N_8427,N_7976,N_7834);
or U8428 (N_8428,N_7821,N_7880);
and U8429 (N_8429,N_7727,N_7909);
nand U8430 (N_8430,N_7883,N_7834);
and U8431 (N_8431,N_7959,N_7867);
nor U8432 (N_8432,N_7848,N_7695);
nand U8433 (N_8433,N_7525,N_7825);
xnor U8434 (N_8434,N_7760,N_7979);
or U8435 (N_8435,N_7856,N_7570);
nor U8436 (N_8436,N_7652,N_7715);
or U8437 (N_8437,N_7542,N_7864);
nand U8438 (N_8438,N_7948,N_7524);
and U8439 (N_8439,N_7774,N_7740);
or U8440 (N_8440,N_7701,N_7621);
xnor U8441 (N_8441,N_7794,N_7572);
nor U8442 (N_8442,N_7658,N_7707);
nor U8443 (N_8443,N_7651,N_7992);
nand U8444 (N_8444,N_7509,N_7520);
xnor U8445 (N_8445,N_7754,N_7864);
nand U8446 (N_8446,N_7985,N_7828);
nor U8447 (N_8447,N_7785,N_7957);
or U8448 (N_8448,N_7797,N_7877);
nand U8449 (N_8449,N_7896,N_7502);
or U8450 (N_8450,N_7919,N_7515);
xnor U8451 (N_8451,N_7783,N_7511);
nand U8452 (N_8452,N_7787,N_7600);
nand U8453 (N_8453,N_7626,N_7763);
xnor U8454 (N_8454,N_7830,N_7934);
nand U8455 (N_8455,N_7892,N_7687);
and U8456 (N_8456,N_7884,N_7813);
xnor U8457 (N_8457,N_7500,N_7612);
and U8458 (N_8458,N_7986,N_7536);
nand U8459 (N_8459,N_7814,N_7915);
xnor U8460 (N_8460,N_7626,N_7595);
and U8461 (N_8461,N_7706,N_7905);
nor U8462 (N_8462,N_7651,N_7936);
xnor U8463 (N_8463,N_7568,N_7717);
or U8464 (N_8464,N_7925,N_7579);
and U8465 (N_8465,N_7597,N_7988);
or U8466 (N_8466,N_7654,N_7870);
nor U8467 (N_8467,N_7630,N_7975);
or U8468 (N_8468,N_7678,N_7784);
xnor U8469 (N_8469,N_7685,N_7558);
nor U8470 (N_8470,N_7571,N_7822);
nand U8471 (N_8471,N_7638,N_7558);
nor U8472 (N_8472,N_7615,N_7899);
nand U8473 (N_8473,N_7952,N_7759);
and U8474 (N_8474,N_7736,N_7515);
xor U8475 (N_8475,N_7711,N_7524);
nor U8476 (N_8476,N_7703,N_7626);
or U8477 (N_8477,N_7559,N_7525);
nand U8478 (N_8478,N_7940,N_7609);
or U8479 (N_8479,N_7871,N_7923);
or U8480 (N_8480,N_7768,N_7712);
or U8481 (N_8481,N_7575,N_7553);
nor U8482 (N_8482,N_7991,N_7676);
or U8483 (N_8483,N_7592,N_7522);
and U8484 (N_8484,N_7612,N_7814);
nor U8485 (N_8485,N_7679,N_7993);
and U8486 (N_8486,N_7846,N_7870);
or U8487 (N_8487,N_7759,N_7543);
and U8488 (N_8488,N_7574,N_7545);
or U8489 (N_8489,N_7901,N_7554);
or U8490 (N_8490,N_7797,N_7556);
or U8491 (N_8491,N_7650,N_7582);
or U8492 (N_8492,N_7583,N_7950);
nor U8493 (N_8493,N_7977,N_7697);
nand U8494 (N_8494,N_7867,N_7749);
xnor U8495 (N_8495,N_7661,N_7921);
nand U8496 (N_8496,N_7761,N_7548);
and U8497 (N_8497,N_7758,N_7835);
xnor U8498 (N_8498,N_7546,N_7752);
or U8499 (N_8499,N_7607,N_7951);
or U8500 (N_8500,N_8301,N_8490);
nand U8501 (N_8501,N_8299,N_8088);
xor U8502 (N_8502,N_8207,N_8430);
and U8503 (N_8503,N_8255,N_8108);
nand U8504 (N_8504,N_8069,N_8355);
nand U8505 (N_8505,N_8464,N_8244);
and U8506 (N_8506,N_8356,N_8466);
and U8507 (N_8507,N_8330,N_8358);
nor U8508 (N_8508,N_8087,N_8059);
xor U8509 (N_8509,N_8128,N_8304);
or U8510 (N_8510,N_8415,N_8376);
and U8511 (N_8511,N_8047,N_8392);
and U8512 (N_8512,N_8484,N_8313);
or U8513 (N_8513,N_8413,N_8257);
nand U8514 (N_8514,N_8414,N_8394);
nor U8515 (N_8515,N_8168,N_8188);
and U8516 (N_8516,N_8010,N_8460);
or U8517 (N_8517,N_8085,N_8037);
xnor U8518 (N_8518,N_8079,N_8176);
or U8519 (N_8519,N_8365,N_8288);
or U8520 (N_8520,N_8293,N_8223);
and U8521 (N_8521,N_8160,N_8316);
nor U8522 (N_8522,N_8473,N_8036);
nor U8523 (N_8523,N_8081,N_8434);
nand U8524 (N_8524,N_8116,N_8467);
or U8525 (N_8525,N_8431,N_8028);
and U8526 (N_8526,N_8171,N_8145);
or U8527 (N_8527,N_8399,N_8384);
nand U8528 (N_8528,N_8364,N_8478);
nor U8529 (N_8529,N_8461,N_8456);
or U8530 (N_8530,N_8311,N_8248);
xnor U8531 (N_8531,N_8155,N_8267);
xnor U8532 (N_8532,N_8105,N_8254);
and U8533 (N_8533,N_8300,N_8418);
nand U8534 (N_8534,N_8017,N_8396);
and U8535 (N_8535,N_8023,N_8095);
nand U8536 (N_8536,N_8219,N_8446);
and U8537 (N_8537,N_8089,N_8419);
xnor U8538 (N_8538,N_8498,N_8112);
nor U8539 (N_8539,N_8133,N_8055);
nor U8540 (N_8540,N_8408,N_8165);
nand U8541 (N_8541,N_8210,N_8329);
or U8542 (N_8542,N_8439,N_8317);
nor U8543 (N_8543,N_8063,N_8092);
nor U8544 (N_8544,N_8080,N_8091);
and U8545 (N_8545,N_8337,N_8336);
or U8546 (N_8546,N_8253,N_8127);
or U8547 (N_8547,N_8362,N_8237);
nand U8548 (N_8548,N_8049,N_8281);
nor U8549 (N_8549,N_8401,N_8177);
and U8550 (N_8550,N_8245,N_8457);
and U8551 (N_8551,N_8051,N_8472);
or U8552 (N_8552,N_8286,N_8346);
nand U8553 (N_8553,N_8012,N_8297);
nand U8554 (N_8554,N_8084,N_8178);
nor U8555 (N_8555,N_8287,N_8154);
and U8556 (N_8556,N_8027,N_8349);
xor U8557 (N_8557,N_8486,N_8305);
and U8558 (N_8558,N_8391,N_8339);
nand U8559 (N_8559,N_8251,N_8496);
xnor U8560 (N_8560,N_8277,N_8314);
nor U8561 (N_8561,N_8389,N_8363);
or U8562 (N_8562,N_8208,N_8372);
and U8563 (N_8563,N_8182,N_8249);
and U8564 (N_8564,N_8021,N_8334);
nand U8565 (N_8565,N_8147,N_8007);
nand U8566 (N_8566,N_8482,N_8427);
nand U8567 (N_8567,N_8064,N_8350);
xnor U8568 (N_8568,N_8322,N_8130);
xor U8569 (N_8569,N_8243,N_8068);
nand U8570 (N_8570,N_8416,N_8260);
or U8571 (N_8571,N_8453,N_8073);
xor U8572 (N_8572,N_8480,N_8435);
nor U8573 (N_8573,N_8371,N_8110);
or U8574 (N_8574,N_8443,N_8163);
and U8575 (N_8575,N_8175,N_8421);
or U8576 (N_8576,N_8377,N_8072);
or U8577 (N_8577,N_8270,N_8052);
nor U8578 (N_8578,N_8132,N_8106);
or U8579 (N_8579,N_8289,N_8444);
and U8580 (N_8580,N_8022,N_8184);
and U8581 (N_8581,N_8437,N_8221);
nand U8582 (N_8582,N_8169,N_8351);
and U8583 (N_8583,N_8200,N_8009);
or U8584 (N_8584,N_8098,N_8387);
and U8585 (N_8585,N_8016,N_8140);
nor U8586 (N_8586,N_8273,N_8048);
nand U8587 (N_8587,N_8279,N_8303);
or U8588 (N_8588,N_8438,N_8475);
and U8589 (N_8589,N_8426,N_8433);
and U8590 (N_8590,N_8468,N_8100);
nor U8591 (N_8591,N_8137,N_8046);
or U8592 (N_8592,N_8422,N_8240);
or U8593 (N_8593,N_8338,N_8264);
nand U8594 (N_8594,N_8216,N_8459);
nor U8595 (N_8595,N_8224,N_8451);
and U8596 (N_8596,N_8020,N_8343);
nor U8597 (N_8597,N_8226,N_8307);
or U8598 (N_8598,N_8462,N_8489);
nand U8599 (N_8599,N_8039,N_8152);
or U8600 (N_8600,N_8044,N_8463);
nand U8601 (N_8601,N_8381,N_8156);
xnor U8602 (N_8602,N_8143,N_8499);
and U8603 (N_8603,N_8231,N_8185);
and U8604 (N_8604,N_8125,N_8295);
xor U8605 (N_8605,N_8405,N_8378);
or U8606 (N_8606,N_8495,N_8187);
nand U8607 (N_8607,N_8388,N_8354);
nor U8608 (N_8608,N_8038,N_8053);
xnor U8609 (N_8609,N_8359,N_8344);
or U8610 (N_8610,N_8082,N_8164);
xnor U8611 (N_8611,N_8310,N_8386);
or U8612 (N_8612,N_8465,N_8144);
nand U8613 (N_8613,N_8192,N_8285);
and U8614 (N_8614,N_8335,N_8308);
and U8615 (N_8615,N_8050,N_8057);
and U8616 (N_8616,N_8246,N_8131);
or U8617 (N_8617,N_8026,N_8306);
or U8618 (N_8618,N_8390,N_8291);
or U8619 (N_8619,N_8442,N_8220);
nand U8620 (N_8620,N_8493,N_8385);
nor U8621 (N_8621,N_8455,N_8258);
nand U8622 (N_8622,N_8159,N_8294);
nand U8623 (N_8623,N_8280,N_8361);
nand U8624 (N_8624,N_8319,N_8271);
xor U8625 (N_8625,N_8158,N_8033);
nand U8626 (N_8626,N_8213,N_8202);
nor U8627 (N_8627,N_8101,N_8229);
xor U8628 (N_8628,N_8126,N_8205);
xor U8629 (N_8629,N_8031,N_8275);
or U8630 (N_8630,N_8167,N_8407);
and U8631 (N_8631,N_8352,N_8485);
xor U8632 (N_8632,N_8097,N_8129);
nor U8633 (N_8633,N_8374,N_8241);
and U8634 (N_8634,N_8206,N_8315);
nor U8635 (N_8635,N_8070,N_8077);
nor U8636 (N_8636,N_8061,N_8189);
or U8637 (N_8637,N_8170,N_8225);
nor U8638 (N_8638,N_8228,N_8491);
xor U8639 (N_8639,N_8488,N_8487);
nor U8640 (N_8640,N_8014,N_8261);
nor U8641 (N_8641,N_8006,N_8458);
xnor U8642 (N_8642,N_8321,N_8274);
or U8643 (N_8643,N_8099,N_8113);
and U8644 (N_8644,N_8449,N_8194);
or U8645 (N_8645,N_8368,N_8076);
and U8646 (N_8646,N_8290,N_8217);
or U8647 (N_8647,N_8004,N_8227);
and U8648 (N_8648,N_8492,N_8276);
and U8649 (N_8649,N_8429,N_8195);
and U8650 (N_8650,N_8262,N_8420);
nand U8651 (N_8651,N_8230,N_8001);
or U8652 (N_8652,N_8296,N_8436);
and U8653 (N_8653,N_8214,N_8424);
or U8654 (N_8654,N_8269,N_8157);
nor U8655 (N_8655,N_8284,N_8029);
nor U8656 (N_8656,N_8065,N_8215);
nor U8657 (N_8657,N_8066,N_8149);
or U8658 (N_8658,N_8323,N_8380);
or U8659 (N_8659,N_8441,N_8342);
or U8660 (N_8660,N_8403,N_8104);
and U8661 (N_8661,N_8043,N_8135);
nor U8662 (N_8662,N_8011,N_8440);
nor U8663 (N_8663,N_8234,N_8183);
or U8664 (N_8664,N_8432,N_8058);
and U8665 (N_8665,N_8201,N_8071);
nand U8666 (N_8666,N_8345,N_8114);
nor U8667 (N_8667,N_8327,N_8173);
or U8668 (N_8668,N_8370,N_8013);
nor U8669 (N_8669,N_8398,N_8186);
nand U8670 (N_8670,N_8174,N_8309);
nand U8671 (N_8671,N_8347,N_8259);
or U8672 (N_8672,N_8115,N_8369);
and U8673 (N_8673,N_8367,N_8268);
nand U8674 (N_8674,N_8139,N_8119);
nor U8675 (N_8675,N_8324,N_8136);
nor U8676 (N_8676,N_8332,N_8040);
nand U8677 (N_8677,N_8479,N_8483);
or U8678 (N_8678,N_8247,N_8180);
and U8679 (N_8679,N_8239,N_8161);
nor U8680 (N_8680,N_8124,N_8002);
or U8681 (N_8681,N_8041,N_8341);
nand U8682 (N_8682,N_8075,N_8162);
nand U8683 (N_8683,N_8193,N_8402);
and U8684 (N_8684,N_8411,N_8181);
nor U8685 (N_8685,N_8078,N_8410);
and U8686 (N_8686,N_8283,N_8000);
nand U8687 (N_8687,N_8109,N_8003);
nand U8688 (N_8688,N_8197,N_8425);
nand U8689 (N_8689,N_8302,N_8141);
or U8690 (N_8690,N_8242,N_8428);
and U8691 (N_8691,N_8117,N_8008);
nand U8692 (N_8692,N_8074,N_8054);
and U8693 (N_8693,N_8045,N_8111);
and U8694 (N_8694,N_8005,N_8400);
nand U8695 (N_8695,N_8320,N_8383);
xnor U8696 (N_8696,N_8042,N_8134);
nor U8697 (N_8697,N_8263,N_8266);
nor U8698 (N_8698,N_8094,N_8476);
and U8699 (N_8699,N_8477,N_8203);
nand U8700 (N_8700,N_8199,N_8015);
nor U8701 (N_8701,N_8179,N_8211);
nor U8702 (N_8702,N_8122,N_8024);
nand U8703 (N_8703,N_8233,N_8474);
xnor U8704 (N_8704,N_8357,N_8150);
xnor U8705 (N_8705,N_8340,N_8328);
nor U8706 (N_8706,N_8360,N_8373);
nand U8707 (N_8707,N_8107,N_8056);
and U8708 (N_8708,N_8412,N_8250);
nand U8709 (N_8709,N_8093,N_8404);
nand U8710 (N_8710,N_8025,N_8212);
and U8711 (N_8711,N_8103,N_8393);
nor U8712 (N_8712,N_8318,N_8382);
and U8713 (N_8713,N_8375,N_8138);
nand U8714 (N_8714,N_8417,N_8256);
nand U8715 (N_8715,N_8236,N_8123);
xor U8716 (N_8716,N_8292,N_8238);
xor U8717 (N_8717,N_8086,N_8153);
or U8718 (N_8718,N_8395,N_8450);
and U8719 (N_8719,N_8190,N_8232);
nor U8720 (N_8720,N_8298,N_8379);
and U8721 (N_8721,N_8034,N_8366);
nor U8722 (N_8722,N_8172,N_8196);
nand U8723 (N_8723,N_8454,N_8397);
nand U8724 (N_8724,N_8018,N_8198);
xnor U8725 (N_8725,N_8235,N_8445);
and U8726 (N_8726,N_8471,N_8032);
nand U8727 (N_8727,N_8209,N_8312);
nand U8728 (N_8728,N_8265,N_8326);
and U8729 (N_8729,N_8035,N_8121);
and U8730 (N_8730,N_8481,N_8148);
or U8731 (N_8731,N_8096,N_8406);
xor U8732 (N_8732,N_8409,N_8331);
nor U8733 (N_8733,N_8030,N_8278);
or U8734 (N_8734,N_8067,N_8083);
and U8735 (N_8735,N_8272,N_8494);
nand U8736 (N_8736,N_8353,N_8497);
or U8737 (N_8737,N_8282,N_8204);
xor U8738 (N_8738,N_8151,N_8102);
nand U8739 (N_8739,N_8452,N_8348);
or U8740 (N_8740,N_8090,N_8222);
xor U8741 (N_8741,N_8333,N_8019);
or U8742 (N_8742,N_8191,N_8218);
and U8743 (N_8743,N_8448,N_8447);
nand U8744 (N_8744,N_8142,N_8470);
nand U8745 (N_8745,N_8423,N_8118);
or U8746 (N_8746,N_8120,N_8146);
and U8747 (N_8747,N_8325,N_8166);
or U8748 (N_8748,N_8252,N_8062);
nand U8749 (N_8749,N_8060,N_8469);
and U8750 (N_8750,N_8196,N_8236);
nor U8751 (N_8751,N_8429,N_8111);
and U8752 (N_8752,N_8381,N_8286);
and U8753 (N_8753,N_8477,N_8204);
nand U8754 (N_8754,N_8361,N_8334);
and U8755 (N_8755,N_8499,N_8005);
nor U8756 (N_8756,N_8063,N_8025);
nor U8757 (N_8757,N_8080,N_8007);
nor U8758 (N_8758,N_8356,N_8250);
nand U8759 (N_8759,N_8061,N_8098);
nand U8760 (N_8760,N_8251,N_8183);
and U8761 (N_8761,N_8353,N_8339);
and U8762 (N_8762,N_8107,N_8093);
and U8763 (N_8763,N_8017,N_8332);
or U8764 (N_8764,N_8118,N_8429);
nand U8765 (N_8765,N_8169,N_8380);
nand U8766 (N_8766,N_8486,N_8283);
nand U8767 (N_8767,N_8476,N_8049);
xnor U8768 (N_8768,N_8355,N_8282);
nor U8769 (N_8769,N_8181,N_8124);
nor U8770 (N_8770,N_8088,N_8389);
nand U8771 (N_8771,N_8292,N_8030);
nor U8772 (N_8772,N_8337,N_8223);
and U8773 (N_8773,N_8063,N_8029);
nand U8774 (N_8774,N_8462,N_8480);
and U8775 (N_8775,N_8143,N_8223);
xor U8776 (N_8776,N_8460,N_8248);
or U8777 (N_8777,N_8423,N_8082);
xor U8778 (N_8778,N_8367,N_8254);
nand U8779 (N_8779,N_8464,N_8156);
nand U8780 (N_8780,N_8147,N_8487);
nand U8781 (N_8781,N_8191,N_8376);
or U8782 (N_8782,N_8447,N_8121);
nor U8783 (N_8783,N_8447,N_8092);
and U8784 (N_8784,N_8492,N_8346);
and U8785 (N_8785,N_8373,N_8420);
and U8786 (N_8786,N_8416,N_8061);
nor U8787 (N_8787,N_8463,N_8066);
and U8788 (N_8788,N_8284,N_8315);
nor U8789 (N_8789,N_8364,N_8144);
nand U8790 (N_8790,N_8371,N_8416);
xor U8791 (N_8791,N_8220,N_8119);
and U8792 (N_8792,N_8481,N_8387);
or U8793 (N_8793,N_8116,N_8061);
nor U8794 (N_8794,N_8185,N_8364);
or U8795 (N_8795,N_8207,N_8089);
nand U8796 (N_8796,N_8125,N_8065);
nand U8797 (N_8797,N_8219,N_8123);
nor U8798 (N_8798,N_8173,N_8313);
or U8799 (N_8799,N_8169,N_8128);
and U8800 (N_8800,N_8449,N_8115);
nor U8801 (N_8801,N_8178,N_8007);
and U8802 (N_8802,N_8000,N_8228);
or U8803 (N_8803,N_8162,N_8222);
or U8804 (N_8804,N_8430,N_8153);
and U8805 (N_8805,N_8313,N_8293);
nor U8806 (N_8806,N_8425,N_8083);
and U8807 (N_8807,N_8062,N_8186);
or U8808 (N_8808,N_8486,N_8115);
nor U8809 (N_8809,N_8106,N_8345);
or U8810 (N_8810,N_8438,N_8224);
nor U8811 (N_8811,N_8084,N_8394);
and U8812 (N_8812,N_8140,N_8403);
xnor U8813 (N_8813,N_8280,N_8215);
nor U8814 (N_8814,N_8460,N_8202);
nand U8815 (N_8815,N_8261,N_8191);
nor U8816 (N_8816,N_8386,N_8086);
and U8817 (N_8817,N_8094,N_8043);
nand U8818 (N_8818,N_8017,N_8335);
nand U8819 (N_8819,N_8109,N_8307);
or U8820 (N_8820,N_8080,N_8014);
and U8821 (N_8821,N_8232,N_8306);
or U8822 (N_8822,N_8086,N_8138);
xor U8823 (N_8823,N_8472,N_8168);
xnor U8824 (N_8824,N_8382,N_8281);
nand U8825 (N_8825,N_8003,N_8231);
or U8826 (N_8826,N_8143,N_8026);
nand U8827 (N_8827,N_8475,N_8465);
nand U8828 (N_8828,N_8065,N_8046);
nand U8829 (N_8829,N_8475,N_8479);
and U8830 (N_8830,N_8005,N_8474);
nand U8831 (N_8831,N_8028,N_8368);
nor U8832 (N_8832,N_8097,N_8058);
xnor U8833 (N_8833,N_8244,N_8406);
xnor U8834 (N_8834,N_8072,N_8473);
and U8835 (N_8835,N_8203,N_8079);
or U8836 (N_8836,N_8212,N_8274);
nand U8837 (N_8837,N_8014,N_8133);
nor U8838 (N_8838,N_8246,N_8437);
xnor U8839 (N_8839,N_8099,N_8320);
or U8840 (N_8840,N_8219,N_8032);
or U8841 (N_8841,N_8010,N_8315);
nor U8842 (N_8842,N_8363,N_8146);
nand U8843 (N_8843,N_8330,N_8099);
nand U8844 (N_8844,N_8258,N_8125);
and U8845 (N_8845,N_8308,N_8479);
or U8846 (N_8846,N_8324,N_8127);
xor U8847 (N_8847,N_8178,N_8203);
nand U8848 (N_8848,N_8369,N_8059);
and U8849 (N_8849,N_8141,N_8136);
or U8850 (N_8850,N_8055,N_8129);
and U8851 (N_8851,N_8469,N_8472);
or U8852 (N_8852,N_8432,N_8461);
nor U8853 (N_8853,N_8372,N_8382);
or U8854 (N_8854,N_8427,N_8030);
or U8855 (N_8855,N_8143,N_8171);
nand U8856 (N_8856,N_8100,N_8102);
nor U8857 (N_8857,N_8042,N_8132);
nor U8858 (N_8858,N_8382,N_8224);
nand U8859 (N_8859,N_8217,N_8252);
or U8860 (N_8860,N_8120,N_8187);
nand U8861 (N_8861,N_8158,N_8051);
or U8862 (N_8862,N_8409,N_8296);
and U8863 (N_8863,N_8315,N_8200);
nor U8864 (N_8864,N_8271,N_8116);
and U8865 (N_8865,N_8026,N_8494);
nor U8866 (N_8866,N_8278,N_8360);
and U8867 (N_8867,N_8050,N_8426);
nor U8868 (N_8868,N_8113,N_8390);
nand U8869 (N_8869,N_8392,N_8290);
nor U8870 (N_8870,N_8203,N_8117);
nand U8871 (N_8871,N_8069,N_8253);
or U8872 (N_8872,N_8437,N_8390);
nor U8873 (N_8873,N_8278,N_8210);
and U8874 (N_8874,N_8251,N_8256);
nand U8875 (N_8875,N_8256,N_8365);
nand U8876 (N_8876,N_8431,N_8052);
nand U8877 (N_8877,N_8208,N_8122);
nor U8878 (N_8878,N_8376,N_8119);
nand U8879 (N_8879,N_8230,N_8120);
nor U8880 (N_8880,N_8154,N_8050);
or U8881 (N_8881,N_8484,N_8419);
or U8882 (N_8882,N_8186,N_8276);
xnor U8883 (N_8883,N_8360,N_8018);
or U8884 (N_8884,N_8316,N_8238);
and U8885 (N_8885,N_8166,N_8020);
and U8886 (N_8886,N_8059,N_8229);
xor U8887 (N_8887,N_8216,N_8321);
nand U8888 (N_8888,N_8418,N_8255);
xnor U8889 (N_8889,N_8420,N_8157);
nand U8890 (N_8890,N_8347,N_8469);
or U8891 (N_8891,N_8201,N_8184);
nor U8892 (N_8892,N_8023,N_8203);
or U8893 (N_8893,N_8295,N_8206);
and U8894 (N_8894,N_8263,N_8390);
and U8895 (N_8895,N_8420,N_8018);
or U8896 (N_8896,N_8343,N_8422);
nor U8897 (N_8897,N_8402,N_8092);
nor U8898 (N_8898,N_8167,N_8079);
or U8899 (N_8899,N_8255,N_8376);
nor U8900 (N_8900,N_8173,N_8049);
nand U8901 (N_8901,N_8453,N_8273);
or U8902 (N_8902,N_8026,N_8201);
nor U8903 (N_8903,N_8365,N_8258);
and U8904 (N_8904,N_8443,N_8034);
and U8905 (N_8905,N_8353,N_8266);
or U8906 (N_8906,N_8003,N_8480);
nand U8907 (N_8907,N_8309,N_8161);
nand U8908 (N_8908,N_8372,N_8496);
nand U8909 (N_8909,N_8069,N_8403);
or U8910 (N_8910,N_8493,N_8043);
or U8911 (N_8911,N_8207,N_8107);
and U8912 (N_8912,N_8012,N_8306);
nor U8913 (N_8913,N_8112,N_8191);
nor U8914 (N_8914,N_8047,N_8395);
and U8915 (N_8915,N_8474,N_8265);
nor U8916 (N_8916,N_8028,N_8290);
nand U8917 (N_8917,N_8170,N_8427);
or U8918 (N_8918,N_8495,N_8251);
or U8919 (N_8919,N_8136,N_8378);
nor U8920 (N_8920,N_8278,N_8447);
nand U8921 (N_8921,N_8293,N_8037);
or U8922 (N_8922,N_8473,N_8188);
and U8923 (N_8923,N_8392,N_8108);
nor U8924 (N_8924,N_8130,N_8181);
or U8925 (N_8925,N_8185,N_8409);
and U8926 (N_8926,N_8163,N_8293);
or U8927 (N_8927,N_8362,N_8461);
nor U8928 (N_8928,N_8273,N_8389);
nand U8929 (N_8929,N_8436,N_8228);
and U8930 (N_8930,N_8088,N_8021);
nand U8931 (N_8931,N_8065,N_8414);
nor U8932 (N_8932,N_8067,N_8412);
xor U8933 (N_8933,N_8048,N_8246);
nand U8934 (N_8934,N_8469,N_8050);
nand U8935 (N_8935,N_8446,N_8248);
nand U8936 (N_8936,N_8355,N_8114);
nand U8937 (N_8937,N_8345,N_8479);
xor U8938 (N_8938,N_8068,N_8433);
xnor U8939 (N_8939,N_8278,N_8196);
or U8940 (N_8940,N_8454,N_8365);
nand U8941 (N_8941,N_8256,N_8211);
or U8942 (N_8942,N_8078,N_8191);
xor U8943 (N_8943,N_8133,N_8264);
xor U8944 (N_8944,N_8122,N_8337);
and U8945 (N_8945,N_8251,N_8053);
or U8946 (N_8946,N_8209,N_8071);
nor U8947 (N_8947,N_8080,N_8040);
nand U8948 (N_8948,N_8402,N_8418);
and U8949 (N_8949,N_8437,N_8180);
and U8950 (N_8950,N_8201,N_8194);
xnor U8951 (N_8951,N_8165,N_8325);
and U8952 (N_8952,N_8115,N_8059);
and U8953 (N_8953,N_8249,N_8012);
xor U8954 (N_8954,N_8124,N_8065);
nand U8955 (N_8955,N_8412,N_8044);
and U8956 (N_8956,N_8468,N_8107);
xor U8957 (N_8957,N_8266,N_8013);
nor U8958 (N_8958,N_8040,N_8111);
nor U8959 (N_8959,N_8107,N_8138);
and U8960 (N_8960,N_8031,N_8332);
or U8961 (N_8961,N_8012,N_8110);
xnor U8962 (N_8962,N_8315,N_8470);
nor U8963 (N_8963,N_8239,N_8300);
and U8964 (N_8964,N_8117,N_8018);
nand U8965 (N_8965,N_8423,N_8302);
and U8966 (N_8966,N_8084,N_8139);
or U8967 (N_8967,N_8046,N_8054);
nand U8968 (N_8968,N_8208,N_8263);
xnor U8969 (N_8969,N_8392,N_8315);
xnor U8970 (N_8970,N_8464,N_8136);
or U8971 (N_8971,N_8373,N_8323);
xnor U8972 (N_8972,N_8394,N_8426);
nand U8973 (N_8973,N_8257,N_8305);
or U8974 (N_8974,N_8427,N_8485);
or U8975 (N_8975,N_8245,N_8169);
nand U8976 (N_8976,N_8050,N_8088);
and U8977 (N_8977,N_8096,N_8211);
and U8978 (N_8978,N_8157,N_8363);
nand U8979 (N_8979,N_8227,N_8484);
and U8980 (N_8980,N_8274,N_8266);
or U8981 (N_8981,N_8414,N_8362);
xnor U8982 (N_8982,N_8444,N_8324);
or U8983 (N_8983,N_8323,N_8028);
nor U8984 (N_8984,N_8189,N_8079);
nor U8985 (N_8985,N_8414,N_8141);
or U8986 (N_8986,N_8081,N_8144);
nor U8987 (N_8987,N_8303,N_8495);
nand U8988 (N_8988,N_8052,N_8458);
nand U8989 (N_8989,N_8065,N_8101);
xnor U8990 (N_8990,N_8478,N_8249);
xor U8991 (N_8991,N_8412,N_8295);
and U8992 (N_8992,N_8198,N_8167);
nor U8993 (N_8993,N_8139,N_8461);
or U8994 (N_8994,N_8098,N_8124);
nor U8995 (N_8995,N_8396,N_8066);
nor U8996 (N_8996,N_8496,N_8436);
or U8997 (N_8997,N_8408,N_8299);
or U8998 (N_8998,N_8127,N_8252);
nor U8999 (N_8999,N_8223,N_8472);
nor U9000 (N_9000,N_8647,N_8888);
nand U9001 (N_9001,N_8953,N_8601);
and U9002 (N_9002,N_8924,N_8609);
and U9003 (N_9003,N_8939,N_8513);
nand U9004 (N_9004,N_8573,N_8827);
nand U9005 (N_9005,N_8949,N_8892);
nor U9006 (N_9006,N_8904,N_8944);
nand U9007 (N_9007,N_8731,N_8561);
nand U9008 (N_9008,N_8828,N_8659);
and U9009 (N_9009,N_8616,N_8652);
xnor U9010 (N_9010,N_8937,N_8841);
xnor U9011 (N_9011,N_8653,N_8893);
or U9012 (N_9012,N_8605,N_8726);
nor U9013 (N_9013,N_8711,N_8568);
and U9014 (N_9014,N_8803,N_8712);
nand U9015 (N_9015,N_8505,N_8899);
nand U9016 (N_9016,N_8762,N_8679);
nand U9017 (N_9017,N_8691,N_8639);
nand U9018 (N_9018,N_8940,N_8690);
and U9019 (N_9019,N_8859,N_8570);
or U9020 (N_9020,N_8694,N_8508);
nand U9021 (N_9021,N_8625,N_8540);
and U9022 (N_9022,N_8914,N_8770);
xor U9023 (N_9023,N_8825,N_8804);
xnor U9024 (N_9024,N_8510,N_8626);
nand U9025 (N_9025,N_8734,N_8722);
and U9026 (N_9026,N_8725,N_8507);
and U9027 (N_9027,N_8983,N_8778);
and U9028 (N_9028,N_8522,N_8801);
and U9029 (N_9029,N_8838,N_8754);
and U9030 (N_9030,N_8797,N_8836);
and U9031 (N_9031,N_8857,N_8539);
nor U9032 (N_9032,N_8771,N_8863);
or U9033 (N_9033,N_8799,N_8531);
nor U9034 (N_9034,N_8535,N_8602);
or U9035 (N_9035,N_8919,N_8648);
nor U9036 (N_9036,N_8945,N_8743);
or U9037 (N_9037,N_8528,N_8514);
nand U9038 (N_9038,N_8868,N_8824);
or U9039 (N_9039,N_8823,N_8707);
xnor U9040 (N_9040,N_8834,N_8637);
and U9041 (N_9041,N_8938,N_8879);
and U9042 (N_9042,N_8987,N_8680);
nand U9043 (N_9043,N_8670,N_8982);
or U9044 (N_9044,N_8622,N_8575);
nor U9045 (N_9045,N_8774,N_8555);
or U9046 (N_9046,N_8651,N_8643);
nor U9047 (N_9047,N_8809,N_8547);
or U9048 (N_9048,N_8693,N_8633);
and U9049 (N_9049,N_8736,N_8644);
xnor U9050 (N_9050,N_8994,N_8800);
nand U9051 (N_9051,N_8941,N_8884);
and U9052 (N_9052,N_8808,N_8960);
nor U9053 (N_9053,N_8735,N_8767);
or U9054 (N_9054,N_8727,N_8764);
or U9055 (N_9055,N_8959,N_8813);
xnor U9056 (N_9056,N_8607,N_8623);
or U9057 (N_9057,N_8847,N_8744);
xnor U9058 (N_9058,N_8966,N_8845);
nor U9059 (N_9059,N_8699,N_8550);
nor U9060 (N_9060,N_8970,N_8793);
or U9061 (N_9061,N_8990,N_8969);
and U9062 (N_9062,N_8759,N_8792);
nand U9063 (N_9063,N_8527,N_8501);
and U9064 (N_9064,N_8955,N_8586);
nor U9065 (N_9065,N_8566,N_8689);
or U9066 (N_9066,N_8806,N_8897);
and U9067 (N_9067,N_8781,N_8766);
or U9068 (N_9068,N_8965,N_8543);
and U9069 (N_9069,N_8738,N_8732);
xor U9070 (N_9070,N_8936,N_8850);
and U9071 (N_9071,N_8521,N_8851);
and U9072 (N_9072,N_8975,N_8589);
or U9073 (N_9073,N_8511,N_8701);
nand U9074 (N_9074,N_8934,N_8604);
and U9075 (N_9075,N_8822,N_8907);
nor U9076 (N_9076,N_8753,N_8819);
or U9077 (N_9077,N_8642,N_8783);
nor U9078 (N_9078,N_8532,N_8594);
or U9079 (N_9079,N_8921,N_8995);
nand U9080 (N_9080,N_8718,N_8925);
nand U9081 (N_9081,N_8668,N_8592);
and U9082 (N_9082,N_8746,N_8509);
xor U9083 (N_9083,N_8979,N_8794);
and U9084 (N_9084,N_8998,N_8871);
or U9085 (N_9085,N_8963,N_8911);
and U9086 (N_9086,N_8844,N_8667);
nand U9087 (N_9087,N_8603,N_8861);
and U9088 (N_9088,N_8910,N_8737);
or U9089 (N_9089,N_8577,N_8719);
and U9090 (N_9090,N_8745,N_8843);
and U9091 (N_9091,N_8943,N_8534);
xnor U9092 (N_9092,N_8752,N_8595);
nand U9093 (N_9093,N_8984,N_8525);
xnor U9094 (N_9094,N_8678,N_8660);
xor U9095 (N_9095,N_8624,N_8887);
nand U9096 (N_9096,N_8741,N_8830);
xnor U9097 (N_9097,N_8634,N_8903);
xnor U9098 (N_9098,N_8533,N_8923);
nand U9099 (N_9099,N_8567,N_8820);
nor U9100 (N_9100,N_8729,N_8890);
nand U9101 (N_9101,N_8777,N_8895);
or U9102 (N_9102,N_8549,N_8551);
or U9103 (N_9103,N_8583,N_8715);
nand U9104 (N_9104,N_8598,N_8536);
or U9105 (N_9105,N_8654,N_8523);
nor U9106 (N_9106,N_8906,N_8661);
nand U9107 (N_9107,N_8870,N_8512);
and U9108 (N_9108,N_8600,N_8790);
nand U9109 (N_9109,N_8858,N_8520);
and U9110 (N_9110,N_8645,N_8829);
and U9111 (N_9111,N_8537,N_8946);
nand U9112 (N_9112,N_8956,N_8541);
nor U9113 (N_9113,N_8872,N_8896);
nand U9114 (N_9114,N_8503,N_8628);
nor U9115 (N_9115,N_8916,N_8933);
nor U9116 (N_9116,N_8529,N_8742);
nand U9117 (N_9117,N_8957,N_8649);
and U9118 (N_9118,N_8913,N_8698);
nor U9119 (N_9119,N_8885,N_8524);
or U9120 (N_9120,N_8818,N_8991);
nand U9121 (N_9121,N_8951,N_8702);
nand U9122 (N_9122,N_8761,N_8849);
nand U9123 (N_9123,N_8671,N_8560);
nor U9124 (N_9124,N_8926,N_8565);
nor U9125 (N_9125,N_8557,N_8931);
nand U9126 (N_9126,N_8553,N_8807);
nand U9127 (N_9127,N_8684,N_8795);
or U9128 (N_9128,N_8848,N_8909);
nor U9129 (N_9129,N_8962,N_8610);
nor U9130 (N_9130,N_8562,N_8703);
xnor U9131 (N_9131,N_8612,N_8591);
nor U9132 (N_9132,N_8985,N_8814);
xor U9133 (N_9133,N_8901,N_8973);
and U9134 (N_9134,N_8915,N_8517);
and U9135 (N_9135,N_8657,N_8563);
and U9136 (N_9136,N_8717,N_8714);
nand U9137 (N_9137,N_8713,N_8996);
nor U9138 (N_9138,N_8831,N_8636);
nor U9139 (N_9139,N_8918,N_8786);
nand U9140 (N_9140,N_8988,N_8976);
nand U9141 (N_9141,N_8672,N_8878);
nor U9142 (N_9142,N_8611,N_8947);
and U9143 (N_9143,N_8687,N_8640);
or U9144 (N_9144,N_8784,N_8796);
nand U9145 (N_9145,N_8564,N_8968);
nand U9146 (N_9146,N_8620,N_8967);
nor U9147 (N_9147,N_8840,N_8812);
nand U9148 (N_9148,N_8578,N_8833);
nand U9149 (N_9149,N_8739,N_8789);
xnor U9150 (N_9150,N_8898,N_8614);
and U9151 (N_9151,N_8750,N_8758);
nor U9152 (N_9152,N_8723,N_8772);
xnor U9153 (N_9153,N_8826,N_8856);
and U9154 (N_9154,N_8697,N_8757);
or U9155 (N_9155,N_8972,N_8958);
nand U9156 (N_9156,N_8681,N_8842);
or U9157 (N_9157,N_8619,N_8632);
and U9158 (N_9158,N_8776,N_8902);
xnor U9159 (N_9159,N_8889,N_8695);
nor U9160 (N_9160,N_8730,N_8805);
and U9161 (N_9161,N_8621,N_8997);
or U9162 (N_9162,N_8655,N_8817);
xnor U9163 (N_9163,N_8705,N_8852);
xor U9164 (N_9164,N_8869,N_8710);
nand U9165 (N_9165,N_8948,N_8846);
nor U9166 (N_9166,N_8545,N_8815);
nand U9167 (N_9167,N_8558,N_8504);
nand U9168 (N_9168,N_8635,N_8688);
or U9169 (N_9169,N_8787,N_8666);
and U9170 (N_9170,N_8627,N_8608);
or U9171 (N_9171,N_8993,N_8894);
nor U9172 (N_9172,N_8585,N_8989);
nor U9173 (N_9173,N_8981,N_8816);
and U9174 (N_9174,N_8683,N_8971);
nand U9175 (N_9175,N_8708,N_8656);
nor U9176 (N_9176,N_8860,N_8999);
nor U9177 (N_9177,N_8552,N_8954);
or U9178 (N_9178,N_8516,N_8709);
and U9179 (N_9179,N_8704,N_8749);
or U9180 (N_9180,N_8986,N_8798);
and U9181 (N_9181,N_8917,N_8854);
nor U9182 (N_9182,N_8876,N_8728);
nand U9183 (N_9183,N_8821,N_8748);
and U9184 (N_9184,N_8500,N_8773);
or U9185 (N_9185,N_8542,N_8935);
nor U9186 (N_9186,N_8641,N_8782);
or U9187 (N_9187,N_8685,N_8733);
xor U9188 (N_9188,N_8839,N_8590);
and U9189 (N_9189,N_8631,N_8669);
or U9190 (N_9190,N_8700,N_8518);
and U9191 (N_9191,N_8961,N_8724);
or U9192 (N_9192,N_8617,N_8629);
nand U9193 (N_9193,N_8877,N_8571);
and U9194 (N_9194,N_8675,N_8587);
nor U9195 (N_9195,N_8886,N_8720);
nor U9196 (N_9196,N_8663,N_8810);
or U9197 (N_9197,N_8593,N_8883);
nand U9198 (N_9198,N_8665,N_8964);
xor U9199 (N_9199,N_8615,N_8788);
nand U9200 (N_9200,N_8584,N_8686);
and U9201 (N_9201,N_8875,N_8874);
and U9202 (N_9202,N_8952,N_8855);
or U9203 (N_9203,N_8928,N_8942);
or U9204 (N_9204,N_8802,N_8572);
nor U9205 (N_9205,N_8912,N_8662);
or U9206 (N_9206,N_8682,N_8646);
or U9207 (N_9207,N_8606,N_8867);
nand U9208 (N_9208,N_8905,N_8932);
and U9209 (N_9209,N_8526,N_8554);
or U9210 (N_9210,N_8599,N_8546);
and U9211 (N_9211,N_8574,N_8588);
or U9212 (N_9212,N_8548,N_8630);
nand U9213 (N_9213,N_8559,N_8880);
and U9214 (N_9214,N_8650,N_8763);
nor U9215 (N_9215,N_8747,N_8992);
nand U9216 (N_9216,N_8751,N_8920);
xnor U9217 (N_9217,N_8811,N_8922);
nor U9218 (N_9218,N_8696,N_8756);
or U9219 (N_9219,N_8908,N_8853);
nor U9220 (N_9220,N_8768,N_8556);
nand U9221 (N_9221,N_8581,N_8579);
nand U9222 (N_9222,N_8769,N_8974);
nand U9223 (N_9223,N_8676,N_8780);
nor U9224 (N_9224,N_8658,N_8674);
and U9225 (N_9225,N_8927,N_8502);
or U9226 (N_9226,N_8891,N_8864);
or U9227 (N_9227,N_8692,N_8862);
xor U9228 (N_9228,N_8835,N_8569);
or U9229 (N_9229,N_8506,N_8538);
nor U9230 (N_9230,N_8882,N_8597);
nand U9231 (N_9231,N_8832,N_8760);
or U9232 (N_9232,N_8765,N_8977);
xor U9233 (N_9233,N_8544,N_8618);
nor U9234 (N_9234,N_8580,N_8613);
and U9235 (N_9235,N_8596,N_8576);
xor U9236 (N_9236,N_8706,N_8673);
and U9237 (N_9237,N_8755,N_8980);
nor U9238 (N_9238,N_8775,N_8519);
or U9239 (N_9239,N_8930,N_8881);
and U9240 (N_9240,N_8785,N_8530);
nor U9241 (N_9241,N_8779,N_8716);
and U9242 (N_9242,N_8950,N_8515);
nand U9243 (N_9243,N_8929,N_8873);
xnor U9244 (N_9244,N_8582,N_8900);
or U9245 (N_9245,N_8791,N_8978);
nor U9246 (N_9246,N_8837,N_8865);
nand U9247 (N_9247,N_8740,N_8638);
xor U9248 (N_9248,N_8664,N_8721);
nand U9249 (N_9249,N_8866,N_8677);
nand U9250 (N_9250,N_8969,N_8997);
or U9251 (N_9251,N_8976,N_8813);
and U9252 (N_9252,N_8705,N_8576);
and U9253 (N_9253,N_8872,N_8866);
and U9254 (N_9254,N_8682,N_8640);
or U9255 (N_9255,N_8831,N_8826);
nand U9256 (N_9256,N_8575,N_8816);
or U9257 (N_9257,N_8654,N_8586);
and U9258 (N_9258,N_8859,N_8831);
nand U9259 (N_9259,N_8679,N_8577);
or U9260 (N_9260,N_8694,N_8996);
nor U9261 (N_9261,N_8952,N_8708);
nand U9262 (N_9262,N_8536,N_8902);
and U9263 (N_9263,N_8769,N_8685);
and U9264 (N_9264,N_8987,N_8749);
xor U9265 (N_9265,N_8784,N_8626);
and U9266 (N_9266,N_8568,N_8713);
nand U9267 (N_9267,N_8659,N_8724);
or U9268 (N_9268,N_8857,N_8504);
or U9269 (N_9269,N_8514,N_8572);
or U9270 (N_9270,N_8979,N_8506);
or U9271 (N_9271,N_8717,N_8948);
and U9272 (N_9272,N_8734,N_8875);
and U9273 (N_9273,N_8688,N_8578);
and U9274 (N_9274,N_8861,N_8747);
and U9275 (N_9275,N_8780,N_8629);
or U9276 (N_9276,N_8856,N_8895);
nor U9277 (N_9277,N_8731,N_8977);
nand U9278 (N_9278,N_8969,N_8799);
nand U9279 (N_9279,N_8539,N_8596);
nand U9280 (N_9280,N_8937,N_8918);
and U9281 (N_9281,N_8707,N_8662);
and U9282 (N_9282,N_8813,N_8693);
or U9283 (N_9283,N_8604,N_8888);
nand U9284 (N_9284,N_8745,N_8554);
nor U9285 (N_9285,N_8548,N_8718);
or U9286 (N_9286,N_8718,N_8526);
and U9287 (N_9287,N_8612,N_8888);
nand U9288 (N_9288,N_8759,N_8707);
nand U9289 (N_9289,N_8780,N_8687);
and U9290 (N_9290,N_8876,N_8791);
nand U9291 (N_9291,N_8510,N_8986);
nand U9292 (N_9292,N_8909,N_8628);
xnor U9293 (N_9293,N_8531,N_8681);
or U9294 (N_9294,N_8921,N_8827);
nand U9295 (N_9295,N_8601,N_8822);
nand U9296 (N_9296,N_8604,N_8753);
nor U9297 (N_9297,N_8600,N_8527);
nand U9298 (N_9298,N_8654,N_8712);
nand U9299 (N_9299,N_8977,N_8967);
or U9300 (N_9300,N_8625,N_8754);
and U9301 (N_9301,N_8571,N_8692);
or U9302 (N_9302,N_8915,N_8719);
nor U9303 (N_9303,N_8696,N_8752);
xor U9304 (N_9304,N_8893,N_8602);
and U9305 (N_9305,N_8682,N_8500);
xnor U9306 (N_9306,N_8857,N_8610);
or U9307 (N_9307,N_8512,N_8852);
and U9308 (N_9308,N_8693,N_8752);
nor U9309 (N_9309,N_8655,N_8551);
or U9310 (N_9310,N_8634,N_8757);
or U9311 (N_9311,N_8937,N_8987);
nand U9312 (N_9312,N_8526,N_8917);
nor U9313 (N_9313,N_8698,N_8824);
xor U9314 (N_9314,N_8601,N_8847);
nor U9315 (N_9315,N_8632,N_8516);
or U9316 (N_9316,N_8596,N_8826);
nand U9317 (N_9317,N_8745,N_8652);
nand U9318 (N_9318,N_8891,N_8704);
or U9319 (N_9319,N_8529,N_8704);
nand U9320 (N_9320,N_8664,N_8967);
or U9321 (N_9321,N_8616,N_8688);
and U9322 (N_9322,N_8608,N_8563);
nor U9323 (N_9323,N_8629,N_8674);
and U9324 (N_9324,N_8564,N_8572);
nand U9325 (N_9325,N_8586,N_8920);
or U9326 (N_9326,N_8688,N_8627);
nor U9327 (N_9327,N_8897,N_8970);
nor U9328 (N_9328,N_8930,N_8851);
nand U9329 (N_9329,N_8627,N_8603);
nand U9330 (N_9330,N_8942,N_8929);
nand U9331 (N_9331,N_8930,N_8853);
xor U9332 (N_9332,N_8573,N_8605);
and U9333 (N_9333,N_8905,N_8651);
xnor U9334 (N_9334,N_8619,N_8899);
and U9335 (N_9335,N_8890,N_8513);
nand U9336 (N_9336,N_8659,N_8857);
or U9337 (N_9337,N_8850,N_8684);
or U9338 (N_9338,N_8629,N_8737);
and U9339 (N_9339,N_8648,N_8954);
nor U9340 (N_9340,N_8957,N_8513);
nand U9341 (N_9341,N_8720,N_8628);
nor U9342 (N_9342,N_8643,N_8624);
and U9343 (N_9343,N_8859,N_8674);
and U9344 (N_9344,N_8853,N_8894);
or U9345 (N_9345,N_8563,N_8721);
and U9346 (N_9346,N_8506,N_8698);
and U9347 (N_9347,N_8707,N_8999);
xor U9348 (N_9348,N_8612,N_8729);
or U9349 (N_9349,N_8671,N_8543);
nor U9350 (N_9350,N_8685,N_8594);
or U9351 (N_9351,N_8505,N_8583);
and U9352 (N_9352,N_8981,N_8739);
nor U9353 (N_9353,N_8726,N_8677);
xor U9354 (N_9354,N_8822,N_8788);
and U9355 (N_9355,N_8866,N_8859);
and U9356 (N_9356,N_8584,N_8864);
nor U9357 (N_9357,N_8717,N_8843);
or U9358 (N_9358,N_8725,N_8518);
and U9359 (N_9359,N_8686,N_8564);
nor U9360 (N_9360,N_8823,N_8647);
nor U9361 (N_9361,N_8582,N_8769);
xor U9362 (N_9362,N_8951,N_8959);
nand U9363 (N_9363,N_8516,N_8648);
or U9364 (N_9364,N_8916,N_8783);
and U9365 (N_9365,N_8565,N_8854);
and U9366 (N_9366,N_8666,N_8784);
nor U9367 (N_9367,N_8551,N_8686);
or U9368 (N_9368,N_8921,N_8807);
nand U9369 (N_9369,N_8729,N_8525);
nand U9370 (N_9370,N_8931,N_8714);
or U9371 (N_9371,N_8618,N_8823);
or U9372 (N_9372,N_8995,N_8619);
or U9373 (N_9373,N_8748,N_8640);
nand U9374 (N_9374,N_8936,N_8931);
nor U9375 (N_9375,N_8982,N_8571);
and U9376 (N_9376,N_8635,N_8568);
nand U9377 (N_9377,N_8740,N_8883);
nor U9378 (N_9378,N_8883,N_8734);
xor U9379 (N_9379,N_8703,N_8598);
nor U9380 (N_9380,N_8626,N_8918);
nand U9381 (N_9381,N_8602,N_8650);
and U9382 (N_9382,N_8577,N_8559);
nand U9383 (N_9383,N_8650,N_8590);
xnor U9384 (N_9384,N_8685,N_8934);
or U9385 (N_9385,N_8607,N_8925);
and U9386 (N_9386,N_8529,N_8755);
and U9387 (N_9387,N_8697,N_8997);
xor U9388 (N_9388,N_8887,N_8954);
or U9389 (N_9389,N_8915,N_8972);
nor U9390 (N_9390,N_8875,N_8585);
xnor U9391 (N_9391,N_8608,N_8912);
nand U9392 (N_9392,N_8993,N_8626);
nor U9393 (N_9393,N_8571,N_8945);
or U9394 (N_9394,N_8574,N_8525);
nor U9395 (N_9395,N_8548,N_8555);
and U9396 (N_9396,N_8649,N_8653);
xnor U9397 (N_9397,N_8605,N_8743);
or U9398 (N_9398,N_8560,N_8995);
nand U9399 (N_9399,N_8832,N_8944);
nor U9400 (N_9400,N_8608,N_8661);
and U9401 (N_9401,N_8904,N_8713);
nand U9402 (N_9402,N_8544,N_8527);
nor U9403 (N_9403,N_8634,N_8670);
nand U9404 (N_9404,N_8558,N_8682);
xor U9405 (N_9405,N_8562,N_8520);
nor U9406 (N_9406,N_8611,N_8874);
and U9407 (N_9407,N_8681,N_8729);
and U9408 (N_9408,N_8543,N_8853);
or U9409 (N_9409,N_8927,N_8625);
or U9410 (N_9410,N_8660,N_8888);
or U9411 (N_9411,N_8881,N_8861);
and U9412 (N_9412,N_8874,N_8789);
and U9413 (N_9413,N_8570,N_8522);
xnor U9414 (N_9414,N_8686,N_8618);
nor U9415 (N_9415,N_8751,N_8942);
or U9416 (N_9416,N_8712,N_8653);
xnor U9417 (N_9417,N_8944,N_8815);
nand U9418 (N_9418,N_8971,N_8634);
and U9419 (N_9419,N_8511,N_8858);
and U9420 (N_9420,N_8637,N_8748);
nor U9421 (N_9421,N_8986,N_8874);
and U9422 (N_9422,N_8974,N_8594);
or U9423 (N_9423,N_8899,N_8706);
nand U9424 (N_9424,N_8948,N_8799);
or U9425 (N_9425,N_8925,N_8943);
nand U9426 (N_9426,N_8730,N_8654);
or U9427 (N_9427,N_8913,N_8881);
nor U9428 (N_9428,N_8785,N_8747);
nor U9429 (N_9429,N_8935,N_8826);
or U9430 (N_9430,N_8737,N_8924);
nor U9431 (N_9431,N_8981,N_8940);
nor U9432 (N_9432,N_8505,N_8921);
or U9433 (N_9433,N_8990,N_8515);
and U9434 (N_9434,N_8776,N_8642);
and U9435 (N_9435,N_8915,N_8706);
nand U9436 (N_9436,N_8931,N_8960);
nor U9437 (N_9437,N_8959,N_8904);
nor U9438 (N_9438,N_8835,N_8577);
or U9439 (N_9439,N_8765,N_8686);
nand U9440 (N_9440,N_8503,N_8735);
or U9441 (N_9441,N_8688,N_8587);
or U9442 (N_9442,N_8658,N_8514);
xnor U9443 (N_9443,N_8936,N_8704);
or U9444 (N_9444,N_8762,N_8862);
nor U9445 (N_9445,N_8955,N_8607);
and U9446 (N_9446,N_8735,N_8597);
or U9447 (N_9447,N_8604,N_8516);
and U9448 (N_9448,N_8810,N_8919);
nor U9449 (N_9449,N_8574,N_8626);
nand U9450 (N_9450,N_8827,N_8978);
nand U9451 (N_9451,N_8915,N_8795);
nor U9452 (N_9452,N_8684,N_8964);
or U9453 (N_9453,N_8771,N_8791);
or U9454 (N_9454,N_8886,N_8564);
nor U9455 (N_9455,N_8691,N_8657);
nand U9456 (N_9456,N_8829,N_8742);
nand U9457 (N_9457,N_8886,N_8935);
nor U9458 (N_9458,N_8624,N_8749);
nor U9459 (N_9459,N_8737,N_8921);
or U9460 (N_9460,N_8508,N_8861);
nand U9461 (N_9461,N_8904,N_8930);
nor U9462 (N_9462,N_8929,N_8978);
or U9463 (N_9463,N_8512,N_8949);
nor U9464 (N_9464,N_8626,N_8823);
and U9465 (N_9465,N_8590,N_8501);
and U9466 (N_9466,N_8989,N_8501);
and U9467 (N_9467,N_8741,N_8765);
nor U9468 (N_9468,N_8809,N_8864);
nand U9469 (N_9469,N_8980,N_8864);
nor U9470 (N_9470,N_8826,N_8956);
xor U9471 (N_9471,N_8799,N_8642);
or U9472 (N_9472,N_8719,N_8778);
or U9473 (N_9473,N_8639,N_8624);
or U9474 (N_9474,N_8855,N_8512);
or U9475 (N_9475,N_8849,N_8516);
nand U9476 (N_9476,N_8544,N_8685);
or U9477 (N_9477,N_8652,N_8937);
nand U9478 (N_9478,N_8751,N_8968);
or U9479 (N_9479,N_8829,N_8546);
and U9480 (N_9480,N_8699,N_8669);
and U9481 (N_9481,N_8817,N_8679);
nor U9482 (N_9482,N_8878,N_8953);
nand U9483 (N_9483,N_8638,N_8789);
nor U9484 (N_9484,N_8798,N_8765);
nand U9485 (N_9485,N_8959,N_8779);
nor U9486 (N_9486,N_8674,N_8526);
nand U9487 (N_9487,N_8865,N_8915);
xnor U9488 (N_9488,N_8783,N_8650);
and U9489 (N_9489,N_8731,N_8894);
or U9490 (N_9490,N_8741,N_8585);
nand U9491 (N_9491,N_8509,N_8782);
xor U9492 (N_9492,N_8969,N_8934);
nand U9493 (N_9493,N_8628,N_8666);
or U9494 (N_9494,N_8784,N_8746);
xnor U9495 (N_9495,N_8880,N_8641);
or U9496 (N_9496,N_8623,N_8958);
nor U9497 (N_9497,N_8853,N_8795);
or U9498 (N_9498,N_8625,N_8595);
or U9499 (N_9499,N_8941,N_8924);
nor U9500 (N_9500,N_9278,N_9114);
nand U9501 (N_9501,N_9410,N_9425);
nor U9502 (N_9502,N_9218,N_9246);
and U9503 (N_9503,N_9036,N_9302);
nor U9504 (N_9504,N_9186,N_9126);
or U9505 (N_9505,N_9123,N_9397);
or U9506 (N_9506,N_9001,N_9280);
or U9507 (N_9507,N_9212,N_9148);
or U9508 (N_9508,N_9402,N_9188);
or U9509 (N_9509,N_9442,N_9165);
and U9510 (N_9510,N_9020,N_9244);
nor U9511 (N_9511,N_9389,N_9092);
or U9512 (N_9512,N_9454,N_9324);
and U9513 (N_9513,N_9460,N_9136);
xor U9514 (N_9514,N_9417,N_9497);
xor U9515 (N_9515,N_9365,N_9271);
nor U9516 (N_9516,N_9264,N_9072);
nand U9517 (N_9517,N_9214,N_9448);
and U9518 (N_9518,N_9311,N_9469);
and U9519 (N_9519,N_9464,N_9489);
nor U9520 (N_9520,N_9172,N_9462);
nor U9521 (N_9521,N_9276,N_9336);
nand U9522 (N_9522,N_9354,N_9491);
nand U9523 (N_9523,N_9414,N_9069);
nor U9524 (N_9524,N_9376,N_9100);
nor U9525 (N_9525,N_9429,N_9248);
nand U9526 (N_9526,N_9117,N_9200);
nor U9527 (N_9527,N_9401,N_9315);
nand U9528 (N_9528,N_9164,N_9011);
or U9529 (N_9529,N_9317,N_9170);
nor U9530 (N_9530,N_9122,N_9438);
or U9531 (N_9531,N_9361,N_9344);
nor U9532 (N_9532,N_9427,N_9277);
nor U9533 (N_9533,N_9030,N_9059);
nand U9534 (N_9534,N_9211,N_9301);
and U9535 (N_9535,N_9289,N_9147);
or U9536 (N_9536,N_9213,N_9225);
and U9537 (N_9537,N_9192,N_9418);
or U9538 (N_9538,N_9499,N_9357);
nand U9539 (N_9539,N_9330,N_9140);
nand U9540 (N_9540,N_9199,N_9384);
or U9541 (N_9541,N_9099,N_9196);
nand U9542 (N_9542,N_9234,N_9028);
nor U9543 (N_9543,N_9159,N_9077);
and U9544 (N_9544,N_9257,N_9413);
or U9545 (N_9545,N_9025,N_9268);
and U9546 (N_9546,N_9203,N_9050);
nor U9547 (N_9547,N_9039,N_9431);
or U9548 (N_9548,N_9042,N_9013);
nor U9549 (N_9549,N_9457,N_9387);
and U9550 (N_9550,N_9000,N_9303);
nand U9551 (N_9551,N_9396,N_9370);
and U9552 (N_9552,N_9002,N_9133);
nor U9553 (N_9553,N_9073,N_9181);
nand U9554 (N_9554,N_9490,N_9441);
nor U9555 (N_9555,N_9012,N_9256);
and U9556 (N_9556,N_9209,N_9091);
nor U9557 (N_9557,N_9048,N_9374);
or U9558 (N_9558,N_9003,N_9157);
and U9559 (N_9559,N_9358,N_9131);
nand U9560 (N_9560,N_9052,N_9482);
nand U9561 (N_9561,N_9406,N_9338);
nor U9562 (N_9562,N_9076,N_9179);
nand U9563 (N_9563,N_9439,N_9296);
nor U9564 (N_9564,N_9216,N_9066);
and U9565 (N_9565,N_9379,N_9183);
xor U9566 (N_9566,N_9240,N_9421);
nor U9567 (N_9567,N_9107,N_9247);
nor U9568 (N_9568,N_9106,N_9177);
and U9569 (N_9569,N_9292,N_9024);
and U9570 (N_9570,N_9057,N_9382);
and U9571 (N_9571,N_9320,N_9022);
nand U9572 (N_9572,N_9120,N_9349);
and U9573 (N_9573,N_9445,N_9051);
or U9574 (N_9574,N_9436,N_9171);
or U9575 (N_9575,N_9056,N_9195);
nand U9576 (N_9576,N_9145,N_9153);
nand U9577 (N_9577,N_9037,N_9262);
nor U9578 (N_9578,N_9251,N_9005);
nor U9579 (N_9579,N_9254,N_9485);
nand U9580 (N_9580,N_9488,N_9486);
nand U9581 (N_9581,N_9156,N_9451);
nand U9582 (N_9582,N_9109,N_9346);
or U9583 (N_9583,N_9217,N_9093);
and U9584 (N_9584,N_9307,N_9061);
or U9585 (N_9585,N_9360,N_9393);
nand U9586 (N_9586,N_9258,N_9407);
nor U9587 (N_9587,N_9388,N_9327);
nand U9588 (N_9588,N_9064,N_9293);
xor U9589 (N_9589,N_9433,N_9071);
and U9590 (N_9590,N_9032,N_9049);
nand U9591 (N_9591,N_9353,N_9475);
or U9592 (N_9592,N_9450,N_9095);
and U9593 (N_9593,N_9252,N_9233);
nor U9594 (N_9594,N_9350,N_9129);
xor U9595 (N_9595,N_9190,N_9287);
nor U9596 (N_9596,N_9340,N_9121);
and U9597 (N_9597,N_9207,N_9381);
or U9598 (N_9598,N_9143,N_9021);
nand U9599 (N_9599,N_9308,N_9161);
and U9600 (N_9600,N_9331,N_9347);
or U9601 (N_9601,N_9204,N_9238);
xnor U9602 (N_9602,N_9038,N_9040);
nand U9603 (N_9603,N_9452,N_9415);
xnor U9604 (N_9604,N_9323,N_9363);
nor U9605 (N_9605,N_9079,N_9453);
nand U9606 (N_9606,N_9319,N_9239);
nor U9607 (N_9607,N_9409,N_9459);
xnor U9608 (N_9608,N_9151,N_9335);
or U9609 (N_9609,N_9149,N_9492);
nand U9610 (N_9610,N_9432,N_9480);
or U9611 (N_9611,N_9206,N_9297);
xor U9612 (N_9612,N_9437,N_9124);
and U9613 (N_9613,N_9312,N_9329);
nor U9614 (N_9614,N_9403,N_9286);
nor U9615 (N_9615,N_9108,N_9006);
or U9616 (N_9616,N_9428,N_9495);
or U9617 (N_9617,N_9102,N_9472);
xor U9618 (N_9618,N_9084,N_9424);
nand U9619 (N_9619,N_9259,N_9279);
xnor U9620 (N_9620,N_9377,N_9313);
and U9621 (N_9621,N_9010,N_9318);
and U9622 (N_9622,N_9112,N_9260);
and U9623 (N_9623,N_9477,N_9373);
and U9624 (N_9624,N_9456,N_9392);
nor U9625 (N_9625,N_9152,N_9103);
or U9626 (N_9626,N_9228,N_9231);
xnor U9627 (N_9627,N_9343,N_9070);
nor U9628 (N_9628,N_9111,N_9269);
or U9629 (N_9629,N_9355,N_9141);
or U9630 (N_9630,N_9339,N_9008);
or U9631 (N_9631,N_9332,N_9250);
or U9632 (N_9632,N_9368,N_9009);
and U9633 (N_9633,N_9322,N_9119);
nor U9634 (N_9634,N_9082,N_9283);
nor U9635 (N_9635,N_9198,N_9187);
nand U9636 (N_9636,N_9362,N_9162);
nand U9637 (N_9637,N_9202,N_9080);
or U9638 (N_9638,N_9185,N_9083);
nor U9639 (N_9639,N_9029,N_9173);
nand U9640 (N_9640,N_9235,N_9222);
and U9641 (N_9641,N_9169,N_9263);
nand U9642 (N_9642,N_9473,N_9175);
and U9643 (N_9643,N_9380,N_9449);
and U9644 (N_9644,N_9383,N_9096);
and U9645 (N_9645,N_9043,N_9325);
nor U9646 (N_9646,N_9180,N_9118);
and U9647 (N_9647,N_9422,N_9144);
and U9648 (N_9648,N_9134,N_9398);
nor U9649 (N_9649,N_9288,N_9366);
nand U9650 (N_9650,N_9054,N_9068);
or U9651 (N_9651,N_9087,N_9110);
or U9652 (N_9652,N_9137,N_9139);
nor U9653 (N_9653,N_9465,N_9337);
nand U9654 (N_9654,N_9146,N_9226);
or U9655 (N_9655,N_9385,N_9201);
or U9656 (N_9656,N_9018,N_9378);
or U9657 (N_9657,N_9310,N_9060);
nor U9658 (N_9658,N_9281,N_9017);
nand U9659 (N_9659,N_9270,N_9423);
nor U9660 (N_9660,N_9295,N_9394);
and U9661 (N_9661,N_9412,N_9466);
nor U9662 (N_9662,N_9487,N_9299);
xnor U9663 (N_9663,N_9285,N_9309);
and U9664 (N_9664,N_9046,N_9154);
or U9665 (N_9665,N_9227,N_9282);
and U9666 (N_9666,N_9342,N_9191);
nand U9667 (N_9667,N_9127,N_9430);
nand U9668 (N_9668,N_9341,N_9007);
or U9669 (N_9669,N_9168,N_9352);
xnor U9670 (N_9670,N_9399,N_9348);
nor U9671 (N_9671,N_9241,N_9088);
nand U9672 (N_9672,N_9027,N_9101);
nand U9673 (N_9673,N_9219,N_9035);
or U9674 (N_9674,N_9078,N_9266);
or U9675 (N_9675,N_9371,N_9434);
nor U9676 (N_9676,N_9483,N_9210);
or U9677 (N_9677,N_9019,N_9494);
nand U9678 (N_9678,N_9205,N_9130);
or U9679 (N_9679,N_9221,N_9390);
nand U9680 (N_9680,N_9160,N_9014);
nor U9681 (N_9681,N_9058,N_9305);
nor U9682 (N_9682,N_9224,N_9386);
xor U9683 (N_9683,N_9135,N_9443);
and U9684 (N_9684,N_9167,N_9408);
and U9685 (N_9685,N_9104,N_9455);
nor U9686 (N_9686,N_9125,N_9345);
nand U9687 (N_9687,N_9481,N_9463);
and U9688 (N_9688,N_9004,N_9208);
nand U9689 (N_9689,N_9420,N_9261);
nor U9690 (N_9690,N_9375,N_9031);
nand U9691 (N_9691,N_9498,N_9045);
nor U9692 (N_9692,N_9306,N_9416);
and U9693 (N_9693,N_9220,N_9215);
or U9694 (N_9694,N_9334,N_9496);
nand U9695 (N_9695,N_9075,N_9467);
nor U9696 (N_9696,N_9484,N_9237);
xnor U9697 (N_9697,N_9189,N_9367);
xnor U9698 (N_9698,N_9094,N_9034);
nand U9699 (N_9699,N_9446,N_9468);
and U9700 (N_9700,N_9391,N_9150);
and U9701 (N_9701,N_9253,N_9138);
or U9702 (N_9702,N_9435,N_9074);
and U9703 (N_9703,N_9193,N_9089);
and U9704 (N_9704,N_9314,N_9326);
nor U9705 (N_9705,N_9411,N_9194);
nor U9706 (N_9706,N_9369,N_9081);
nand U9707 (N_9707,N_9444,N_9275);
nand U9708 (N_9708,N_9098,N_9440);
and U9709 (N_9709,N_9458,N_9267);
and U9710 (N_9710,N_9113,N_9333);
xnor U9711 (N_9711,N_9232,N_9033);
xor U9712 (N_9712,N_9294,N_9236);
and U9713 (N_9713,N_9023,N_9166);
or U9714 (N_9714,N_9395,N_9359);
nor U9715 (N_9715,N_9163,N_9426);
xnor U9716 (N_9716,N_9223,N_9493);
and U9717 (N_9717,N_9041,N_9328);
and U9718 (N_9718,N_9016,N_9053);
nor U9719 (N_9719,N_9174,N_9085);
and U9720 (N_9720,N_9063,N_9321);
or U9721 (N_9721,N_9273,N_9298);
nor U9722 (N_9722,N_9116,N_9097);
nand U9723 (N_9723,N_9479,N_9478);
nand U9724 (N_9724,N_9055,N_9158);
nand U9725 (N_9725,N_9142,N_9067);
nand U9726 (N_9726,N_9128,N_9476);
or U9727 (N_9727,N_9356,N_9419);
nand U9728 (N_9728,N_9364,N_9265);
nor U9729 (N_9729,N_9155,N_9090);
nand U9730 (N_9730,N_9132,N_9176);
or U9731 (N_9731,N_9178,N_9230);
nor U9732 (N_9732,N_9351,N_9182);
or U9733 (N_9733,N_9229,N_9242);
or U9734 (N_9734,N_9461,N_9044);
xor U9735 (N_9735,N_9372,N_9300);
xnor U9736 (N_9736,N_9470,N_9105);
nand U9737 (N_9737,N_9447,N_9026);
nor U9738 (N_9738,N_9316,N_9249);
nor U9739 (N_9739,N_9474,N_9086);
or U9740 (N_9740,N_9015,N_9404);
and U9741 (N_9741,N_9274,N_9197);
or U9742 (N_9742,N_9184,N_9243);
and U9743 (N_9743,N_9284,N_9290);
nor U9744 (N_9744,N_9255,N_9272);
and U9745 (N_9745,N_9304,N_9400);
nor U9746 (N_9746,N_9065,N_9471);
and U9747 (N_9747,N_9047,N_9245);
or U9748 (N_9748,N_9062,N_9405);
nand U9749 (N_9749,N_9115,N_9291);
nand U9750 (N_9750,N_9177,N_9030);
nand U9751 (N_9751,N_9158,N_9035);
and U9752 (N_9752,N_9303,N_9134);
and U9753 (N_9753,N_9280,N_9356);
and U9754 (N_9754,N_9019,N_9149);
nand U9755 (N_9755,N_9435,N_9022);
or U9756 (N_9756,N_9248,N_9456);
and U9757 (N_9757,N_9499,N_9132);
nand U9758 (N_9758,N_9445,N_9094);
or U9759 (N_9759,N_9472,N_9319);
and U9760 (N_9760,N_9103,N_9385);
nor U9761 (N_9761,N_9109,N_9489);
or U9762 (N_9762,N_9117,N_9237);
or U9763 (N_9763,N_9458,N_9349);
nor U9764 (N_9764,N_9220,N_9048);
or U9765 (N_9765,N_9388,N_9342);
nor U9766 (N_9766,N_9490,N_9482);
or U9767 (N_9767,N_9157,N_9052);
nor U9768 (N_9768,N_9417,N_9065);
nor U9769 (N_9769,N_9340,N_9186);
xnor U9770 (N_9770,N_9154,N_9057);
xor U9771 (N_9771,N_9403,N_9126);
nor U9772 (N_9772,N_9011,N_9329);
nor U9773 (N_9773,N_9444,N_9356);
nand U9774 (N_9774,N_9199,N_9089);
or U9775 (N_9775,N_9449,N_9477);
or U9776 (N_9776,N_9082,N_9214);
nor U9777 (N_9777,N_9397,N_9432);
nand U9778 (N_9778,N_9176,N_9259);
nor U9779 (N_9779,N_9208,N_9204);
or U9780 (N_9780,N_9421,N_9159);
nand U9781 (N_9781,N_9135,N_9229);
nor U9782 (N_9782,N_9282,N_9054);
nand U9783 (N_9783,N_9418,N_9397);
and U9784 (N_9784,N_9395,N_9264);
or U9785 (N_9785,N_9363,N_9072);
and U9786 (N_9786,N_9258,N_9460);
nand U9787 (N_9787,N_9056,N_9069);
and U9788 (N_9788,N_9361,N_9338);
nor U9789 (N_9789,N_9353,N_9136);
nor U9790 (N_9790,N_9460,N_9230);
or U9791 (N_9791,N_9036,N_9064);
or U9792 (N_9792,N_9211,N_9467);
nor U9793 (N_9793,N_9393,N_9003);
or U9794 (N_9794,N_9028,N_9295);
or U9795 (N_9795,N_9422,N_9180);
or U9796 (N_9796,N_9295,N_9200);
nand U9797 (N_9797,N_9322,N_9445);
nor U9798 (N_9798,N_9149,N_9065);
and U9799 (N_9799,N_9463,N_9113);
nand U9800 (N_9800,N_9112,N_9290);
or U9801 (N_9801,N_9071,N_9236);
nand U9802 (N_9802,N_9203,N_9234);
or U9803 (N_9803,N_9301,N_9497);
xor U9804 (N_9804,N_9497,N_9356);
nor U9805 (N_9805,N_9166,N_9111);
xor U9806 (N_9806,N_9053,N_9250);
and U9807 (N_9807,N_9028,N_9394);
or U9808 (N_9808,N_9392,N_9236);
and U9809 (N_9809,N_9028,N_9443);
nor U9810 (N_9810,N_9499,N_9337);
or U9811 (N_9811,N_9307,N_9203);
and U9812 (N_9812,N_9498,N_9227);
or U9813 (N_9813,N_9014,N_9369);
nor U9814 (N_9814,N_9400,N_9469);
nand U9815 (N_9815,N_9075,N_9087);
or U9816 (N_9816,N_9021,N_9421);
nor U9817 (N_9817,N_9248,N_9329);
or U9818 (N_9818,N_9461,N_9255);
or U9819 (N_9819,N_9278,N_9468);
xor U9820 (N_9820,N_9249,N_9070);
nor U9821 (N_9821,N_9460,N_9284);
nor U9822 (N_9822,N_9028,N_9143);
or U9823 (N_9823,N_9362,N_9003);
nor U9824 (N_9824,N_9298,N_9152);
nand U9825 (N_9825,N_9308,N_9132);
nor U9826 (N_9826,N_9183,N_9191);
nand U9827 (N_9827,N_9214,N_9247);
nor U9828 (N_9828,N_9277,N_9152);
nor U9829 (N_9829,N_9140,N_9061);
nor U9830 (N_9830,N_9156,N_9216);
nand U9831 (N_9831,N_9468,N_9224);
and U9832 (N_9832,N_9148,N_9447);
nand U9833 (N_9833,N_9005,N_9001);
nor U9834 (N_9834,N_9362,N_9453);
xor U9835 (N_9835,N_9205,N_9399);
nor U9836 (N_9836,N_9013,N_9372);
or U9837 (N_9837,N_9106,N_9138);
nor U9838 (N_9838,N_9299,N_9476);
nand U9839 (N_9839,N_9356,N_9435);
or U9840 (N_9840,N_9089,N_9013);
nor U9841 (N_9841,N_9433,N_9414);
or U9842 (N_9842,N_9215,N_9410);
nand U9843 (N_9843,N_9336,N_9253);
and U9844 (N_9844,N_9186,N_9467);
nand U9845 (N_9845,N_9064,N_9487);
or U9846 (N_9846,N_9424,N_9279);
nand U9847 (N_9847,N_9181,N_9265);
or U9848 (N_9848,N_9165,N_9471);
or U9849 (N_9849,N_9310,N_9330);
and U9850 (N_9850,N_9126,N_9253);
nand U9851 (N_9851,N_9329,N_9405);
and U9852 (N_9852,N_9486,N_9458);
or U9853 (N_9853,N_9083,N_9001);
nor U9854 (N_9854,N_9090,N_9348);
nor U9855 (N_9855,N_9414,N_9195);
nor U9856 (N_9856,N_9115,N_9330);
nor U9857 (N_9857,N_9161,N_9198);
and U9858 (N_9858,N_9421,N_9487);
and U9859 (N_9859,N_9224,N_9399);
and U9860 (N_9860,N_9086,N_9454);
and U9861 (N_9861,N_9325,N_9385);
nor U9862 (N_9862,N_9127,N_9448);
or U9863 (N_9863,N_9462,N_9428);
and U9864 (N_9864,N_9263,N_9089);
nand U9865 (N_9865,N_9400,N_9336);
nor U9866 (N_9866,N_9060,N_9021);
xnor U9867 (N_9867,N_9413,N_9131);
nor U9868 (N_9868,N_9482,N_9412);
or U9869 (N_9869,N_9447,N_9340);
and U9870 (N_9870,N_9122,N_9232);
nor U9871 (N_9871,N_9307,N_9334);
or U9872 (N_9872,N_9174,N_9416);
nor U9873 (N_9873,N_9434,N_9233);
nand U9874 (N_9874,N_9359,N_9184);
nor U9875 (N_9875,N_9002,N_9394);
and U9876 (N_9876,N_9195,N_9261);
or U9877 (N_9877,N_9155,N_9356);
and U9878 (N_9878,N_9048,N_9093);
or U9879 (N_9879,N_9401,N_9025);
and U9880 (N_9880,N_9321,N_9286);
nor U9881 (N_9881,N_9125,N_9493);
xnor U9882 (N_9882,N_9439,N_9236);
xnor U9883 (N_9883,N_9055,N_9124);
nor U9884 (N_9884,N_9485,N_9134);
or U9885 (N_9885,N_9026,N_9334);
nand U9886 (N_9886,N_9261,N_9467);
and U9887 (N_9887,N_9288,N_9222);
or U9888 (N_9888,N_9467,N_9426);
nor U9889 (N_9889,N_9171,N_9472);
nor U9890 (N_9890,N_9042,N_9420);
and U9891 (N_9891,N_9354,N_9304);
nand U9892 (N_9892,N_9126,N_9172);
and U9893 (N_9893,N_9250,N_9086);
xor U9894 (N_9894,N_9351,N_9461);
nand U9895 (N_9895,N_9210,N_9278);
xor U9896 (N_9896,N_9488,N_9293);
and U9897 (N_9897,N_9354,N_9460);
and U9898 (N_9898,N_9204,N_9164);
nor U9899 (N_9899,N_9162,N_9321);
nand U9900 (N_9900,N_9053,N_9475);
xor U9901 (N_9901,N_9435,N_9157);
or U9902 (N_9902,N_9161,N_9096);
or U9903 (N_9903,N_9101,N_9403);
and U9904 (N_9904,N_9419,N_9311);
nand U9905 (N_9905,N_9438,N_9294);
nand U9906 (N_9906,N_9096,N_9030);
nand U9907 (N_9907,N_9396,N_9208);
xor U9908 (N_9908,N_9104,N_9421);
and U9909 (N_9909,N_9411,N_9096);
and U9910 (N_9910,N_9228,N_9336);
nand U9911 (N_9911,N_9058,N_9391);
and U9912 (N_9912,N_9308,N_9041);
or U9913 (N_9913,N_9287,N_9166);
nand U9914 (N_9914,N_9280,N_9018);
or U9915 (N_9915,N_9069,N_9271);
xnor U9916 (N_9916,N_9273,N_9201);
and U9917 (N_9917,N_9266,N_9020);
or U9918 (N_9918,N_9079,N_9187);
nand U9919 (N_9919,N_9217,N_9473);
nor U9920 (N_9920,N_9302,N_9423);
and U9921 (N_9921,N_9230,N_9268);
nand U9922 (N_9922,N_9185,N_9349);
and U9923 (N_9923,N_9235,N_9069);
xnor U9924 (N_9924,N_9012,N_9016);
and U9925 (N_9925,N_9003,N_9188);
xor U9926 (N_9926,N_9223,N_9014);
and U9927 (N_9927,N_9081,N_9041);
and U9928 (N_9928,N_9065,N_9382);
nor U9929 (N_9929,N_9207,N_9015);
and U9930 (N_9930,N_9027,N_9290);
nand U9931 (N_9931,N_9266,N_9215);
nand U9932 (N_9932,N_9298,N_9151);
and U9933 (N_9933,N_9497,N_9343);
nor U9934 (N_9934,N_9123,N_9245);
nor U9935 (N_9935,N_9320,N_9203);
or U9936 (N_9936,N_9343,N_9161);
nand U9937 (N_9937,N_9198,N_9185);
nor U9938 (N_9938,N_9038,N_9365);
xor U9939 (N_9939,N_9308,N_9253);
nor U9940 (N_9940,N_9467,N_9298);
and U9941 (N_9941,N_9269,N_9272);
or U9942 (N_9942,N_9243,N_9072);
nand U9943 (N_9943,N_9046,N_9453);
nand U9944 (N_9944,N_9292,N_9229);
nor U9945 (N_9945,N_9383,N_9128);
xnor U9946 (N_9946,N_9110,N_9161);
xor U9947 (N_9947,N_9403,N_9019);
or U9948 (N_9948,N_9377,N_9464);
nor U9949 (N_9949,N_9238,N_9279);
nor U9950 (N_9950,N_9085,N_9184);
nor U9951 (N_9951,N_9265,N_9283);
nor U9952 (N_9952,N_9301,N_9449);
nand U9953 (N_9953,N_9077,N_9154);
or U9954 (N_9954,N_9069,N_9244);
and U9955 (N_9955,N_9111,N_9114);
and U9956 (N_9956,N_9469,N_9306);
and U9957 (N_9957,N_9054,N_9364);
xnor U9958 (N_9958,N_9220,N_9280);
nor U9959 (N_9959,N_9156,N_9037);
and U9960 (N_9960,N_9027,N_9044);
and U9961 (N_9961,N_9272,N_9181);
or U9962 (N_9962,N_9395,N_9215);
nand U9963 (N_9963,N_9250,N_9166);
or U9964 (N_9964,N_9018,N_9129);
nand U9965 (N_9965,N_9076,N_9102);
and U9966 (N_9966,N_9110,N_9304);
or U9967 (N_9967,N_9347,N_9182);
nand U9968 (N_9968,N_9223,N_9478);
xnor U9969 (N_9969,N_9040,N_9312);
nand U9970 (N_9970,N_9111,N_9154);
nand U9971 (N_9971,N_9185,N_9078);
and U9972 (N_9972,N_9025,N_9244);
or U9973 (N_9973,N_9238,N_9414);
nand U9974 (N_9974,N_9322,N_9380);
or U9975 (N_9975,N_9378,N_9384);
or U9976 (N_9976,N_9322,N_9480);
nand U9977 (N_9977,N_9449,N_9288);
or U9978 (N_9978,N_9163,N_9454);
nand U9979 (N_9979,N_9439,N_9452);
nor U9980 (N_9980,N_9400,N_9294);
nor U9981 (N_9981,N_9322,N_9275);
and U9982 (N_9982,N_9368,N_9235);
and U9983 (N_9983,N_9016,N_9242);
or U9984 (N_9984,N_9418,N_9108);
nor U9985 (N_9985,N_9029,N_9393);
or U9986 (N_9986,N_9118,N_9210);
and U9987 (N_9987,N_9275,N_9143);
xor U9988 (N_9988,N_9134,N_9299);
nor U9989 (N_9989,N_9285,N_9162);
and U9990 (N_9990,N_9150,N_9194);
xnor U9991 (N_9991,N_9200,N_9356);
and U9992 (N_9992,N_9214,N_9251);
and U9993 (N_9993,N_9182,N_9251);
or U9994 (N_9994,N_9163,N_9018);
nand U9995 (N_9995,N_9443,N_9355);
xnor U9996 (N_9996,N_9329,N_9135);
nand U9997 (N_9997,N_9173,N_9245);
or U9998 (N_9998,N_9371,N_9012);
xor U9999 (N_9999,N_9156,N_9208);
xor U10000 (N_10000,N_9609,N_9874);
nor U10001 (N_10001,N_9978,N_9674);
or U10002 (N_10002,N_9859,N_9907);
and U10003 (N_10003,N_9543,N_9990);
nor U10004 (N_10004,N_9573,N_9505);
and U10005 (N_10005,N_9503,N_9793);
or U10006 (N_10006,N_9569,N_9718);
nor U10007 (N_10007,N_9871,N_9924);
or U10008 (N_10008,N_9676,N_9766);
nor U10009 (N_10009,N_9958,N_9646);
xor U10010 (N_10010,N_9783,N_9937);
nor U10011 (N_10011,N_9969,N_9513);
and U10012 (N_10012,N_9815,N_9555);
and U10013 (N_10013,N_9633,N_9743);
nand U10014 (N_10014,N_9568,N_9798);
or U10015 (N_10015,N_9515,N_9845);
nand U10016 (N_10016,N_9854,N_9911);
nor U10017 (N_10017,N_9868,N_9532);
and U10018 (N_10018,N_9946,N_9623);
or U10019 (N_10019,N_9919,N_9710);
nand U10020 (N_10020,N_9781,N_9677);
nor U10021 (N_10021,N_9920,N_9934);
nor U10022 (N_10022,N_9847,N_9707);
or U10023 (N_10023,N_9551,N_9735);
nor U10024 (N_10024,N_9620,N_9790);
nand U10025 (N_10025,N_9784,N_9604);
nand U10026 (N_10026,N_9891,N_9835);
and U10027 (N_10027,N_9510,N_9690);
nand U10028 (N_10028,N_9945,N_9948);
nor U10029 (N_10029,N_9703,N_9949);
nor U10030 (N_10030,N_9890,N_9849);
and U10031 (N_10031,N_9590,N_9522);
and U10032 (N_10032,N_9545,N_9720);
or U10033 (N_10033,N_9893,N_9819);
or U10034 (N_10034,N_9579,N_9561);
nor U10035 (N_10035,N_9827,N_9556);
and U10036 (N_10036,N_9776,N_9673);
nor U10037 (N_10037,N_9908,N_9968);
nand U10038 (N_10038,N_9980,N_9977);
nor U10039 (N_10039,N_9805,N_9615);
xnor U10040 (N_10040,N_9559,N_9898);
nand U10041 (N_10041,N_9747,N_9983);
nor U10042 (N_10042,N_9600,N_9836);
nor U10043 (N_10043,N_9638,N_9960);
and U10044 (N_10044,N_9933,N_9804);
and U10045 (N_10045,N_9918,N_9666);
nor U10046 (N_10046,N_9640,N_9962);
and U10047 (N_10047,N_9680,N_9509);
or U10048 (N_10048,N_9597,N_9668);
nand U10049 (N_10049,N_9756,N_9952);
or U10050 (N_10050,N_9996,N_9801);
nand U10051 (N_10051,N_9755,N_9731);
and U10052 (N_10052,N_9702,N_9560);
or U10053 (N_10053,N_9661,N_9758);
or U10054 (N_10054,N_9750,N_9669);
nand U10055 (N_10055,N_9976,N_9901);
and U10056 (N_10056,N_9809,N_9535);
nor U10057 (N_10057,N_9651,N_9670);
nor U10058 (N_10058,N_9991,N_9916);
nand U10059 (N_10059,N_9998,N_9672);
nand U10060 (N_10060,N_9923,N_9530);
or U10061 (N_10061,N_9899,N_9992);
nand U10062 (N_10062,N_9634,N_9955);
nand U10063 (N_10063,N_9981,N_9523);
xor U10064 (N_10064,N_9546,N_9812);
xnor U10065 (N_10065,N_9850,N_9824);
nand U10066 (N_10066,N_9709,N_9915);
and U10067 (N_10067,N_9917,N_9914);
nor U10068 (N_10068,N_9664,N_9502);
or U10069 (N_10069,N_9734,N_9950);
xnor U10070 (N_10070,N_9879,N_9741);
nor U10071 (N_10071,N_9571,N_9733);
nand U10072 (N_10072,N_9885,N_9764);
or U10073 (N_10073,N_9507,N_9662);
nor U10074 (N_10074,N_9882,N_9792);
nor U10075 (N_10075,N_9577,N_9873);
and U10076 (N_10076,N_9542,N_9653);
or U10077 (N_10077,N_9654,N_9880);
or U10078 (N_10078,N_9504,N_9944);
or U10079 (N_10079,N_9842,N_9831);
or U10080 (N_10080,N_9811,N_9925);
or U10081 (N_10081,N_9693,N_9697);
or U10082 (N_10082,N_9536,N_9829);
nand U10083 (N_10083,N_9994,N_9541);
nor U10084 (N_10084,N_9770,N_9681);
and U10085 (N_10085,N_9788,N_9726);
and U10086 (N_10086,N_9823,N_9947);
nor U10087 (N_10087,N_9685,N_9773);
or U10088 (N_10088,N_9956,N_9860);
nor U10089 (N_10089,N_9691,N_9951);
nand U10090 (N_10090,N_9594,N_9686);
and U10091 (N_10091,N_9926,N_9900);
nand U10092 (N_10092,N_9637,N_9699);
nor U10093 (N_10093,N_9759,N_9621);
or U10094 (N_10094,N_9822,N_9886);
nand U10095 (N_10095,N_9997,N_9730);
xor U10096 (N_10096,N_9524,N_9761);
and U10097 (N_10097,N_9554,N_9979);
or U10098 (N_10098,N_9993,N_9779);
nand U10099 (N_10099,N_9618,N_9807);
and U10100 (N_10100,N_9632,N_9749);
nand U10101 (N_10101,N_9563,N_9705);
or U10102 (N_10102,N_9768,N_9692);
xnor U10103 (N_10103,N_9663,N_9843);
nand U10104 (N_10104,N_9881,N_9675);
or U10105 (N_10105,N_9862,N_9598);
and U10106 (N_10106,N_9531,N_9762);
or U10107 (N_10107,N_9601,N_9953);
and U10108 (N_10108,N_9574,N_9625);
or U10109 (N_10109,N_9910,N_9712);
or U10110 (N_10110,N_9777,N_9639);
and U10111 (N_10111,N_9595,N_9570);
or U10112 (N_10112,N_9642,N_9866);
xor U10113 (N_10113,N_9902,N_9520);
nor U10114 (N_10114,N_9782,N_9533);
xnor U10115 (N_10115,N_9739,N_9737);
and U10116 (N_10116,N_9820,N_9723);
xor U10117 (N_10117,N_9665,N_9713);
xor U10118 (N_10118,N_9635,N_9856);
or U10119 (N_10119,N_9682,N_9678);
or U10120 (N_10120,N_9647,N_9557);
or U10121 (N_10121,N_9736,N_9817);
nor U10122 (N_10122,N_9722,N_9521);
or U10123 (N_10123,N_9791,N_9658);
nand U10124 (N_10124,N_9825,N_9789);
and U10125 (N_10125,N_9629,N_9772);
nor U10126 (N_10126,N_9622,N_9786);
nand U10127 (N_10127,N_9821,N_9644);
nor U10128 (N_10128,N_9580,N_9613);
xnor U10129 (N_10129,N_9857,N_9922);
nor U10130 (N_10130,N_9895,N_9905);
nor U10131 (N_10131,N_9909,N_9769);
nand U10132 (N_10132,N_9519,N_9855);
nor U10133 (N_10133,N_9548,N_9695);
nand U10134 (N_10134,N_9610,N_9514);
and U10135 (N_10135,N_9897,N_9775);
or U10136 (N_10136,N_9606,N_9566);
or U10137 (N_10137,N_9935,N_9869);
nand U10138 (N_10138,N_9887,N_9501);
and U10139 (N_10139,N_9974,N_9550);
nor U10140 (N_10140,N_9906,N_9921);
or U10141 (N_10141,N_9834,N_9913);
and U10142 (N_10142,N_9552,N_9975);
or U10143 (N_10143,N_9547,N_9785);
nand U10144 (N_10144,N_9567,N_9841);
or U10145 (N_10145,N_9527,N_9806);
nand U10146 (N_10146,N_9716,N_9701);
nor U10147 (N_10147,N_9752,N_9592);
and U10148 (N_10148,N_9837,N_9576);
nor U10149 (N_10149,N_9553,N_9867);
and U10150 (N_10150,N_9539,N_9534);
nor U10151 (N_10151,N_9982,N_9795);
xor U10152 (N_10152,N_9848,N_9989);
or U10153 (N_10153,N_9889,N_9748);
and U10154 (N_10154,N_9517,N_9813);
nand U10155 (N_10155,N_9689,N_9754);
nor U10156 (N_10156,N_9999,N_9591);
nor U10157 (N_10157,N_9603,N_9799);
nor U10158 (N_10158,N_9986,N_9802);
and U10159 (N_10159,N_9753,N_9888);
xor U10160 (N_10160,N_9954,N_9729);
nor U10161 (N_10161,N_9683,N_9537);
or U10162 (N_10162,N_9932,N_9896);
nand U10163 (N_10163,N_9744,N_9578);
or U10164 (N_10164,N_9616,N_9732);
nor U10165 (N_10165,N_9596,N_9648);
nand U10166 (N_10166,N_9608,N_9780);
nand U10167 (N_10167,N_9704,N_9738);
nand U10168 (N_10168,N_9605,N_9645);
or U10169 (N_10169,N_9544,N_9858);
nand U10170 (N_10170,N_9655,N_9833);
or U10171 (N_10171,N_9941,N_9963);
nor U10172 (N_10172,N_9828,N_9724);
and U10173 (N_10173,N_9714,N_9508);
or U10174 (N_10174,N_9984,N_9971);
or U10175 (N_10175,N_9787,N_9959);
nand U10176 (N_10176,N_9583,N_9771);
and U10177 (N_10177,N_9814,N_9582);
and U10178 (N_10178,N_9763,N_9586);
and U10179 (N_10179,N_9564,N_9745);
nor U10180 (N_10180,N_9558,N_9650);
nand U10181 (N_10181,N_9767,N_9972);
or U10182 (N_10182,N_9565,N_9853);
or U10183 (N_10183,N_9728,N_9538);
nor U10184 (N_10184,N_9757,N_9528);
nand U10185 (N_10185,N_9721,N_9904);
and U10186 (N_10186,N_9988,N_9800);
and U10187 (N_10187,N_9746,N_9684);
nor U10188 (N_10188,N_9864,N_9865);
nand U10189 (N_10189,N_9961,N_9816);
nor U10190 (N_10190,N_9725,N_9765);
and U10191 (N_10191,N_9927,N_9587);
or U10192 (N_10192,N_9870,N_9584);
and U10193 (N_10193,N_9656,N_9760);
nor U10194 (N_10194,N_9851,N_9774);
or U10195 (N_10195,N_9778,N_9830);
nor U10196 (N_10196,N_9940,N_9631);
or U10197 (N_10197,N_9516,N_9740);
or U10198 (N_10198,N_9985,N_9844);
or U10199 (N_10199,N_9627,N_9796);
or U10200 (N_10200,N_9742,N_9624);
nand U10201 (N_10201,N_9942,N_9832);
nor U10202 (N_10202,N_9943,N_9585);
nand U10203 (N_10203,N_9694,N_9876);
nand U10204 (N_10204,N_9839,N_9688);
nor U10205 (N_10205,N_9928,N_9549);
nor U10206 (N_10206,N_9652,N_9797);
nand U10207 (N_10207,N_9657,N_9929);
or U10208 (N_10208,N_9818,N_9589);
nor U10209 (N_10209,N_9711,N_9526);
or U10210 (N_10210,N_9727,N_9973);
and U10211 (N_10211,N_9679,N_9863);
xnor U10212 (N_10212,N_9826,N_9964);
nand U10213 (N_10213,N_9529,N_9698);
nand U10214 (N_10214,N_9619,N_9687);
or U10215 (N_10215,N_9614,N_9602);
and U10216 (N_10216,N_9803,N_9717);
nand U10217 (N_10217,N_9512,N_9612);
or U10218 (N_10218,N_9626,N_9967);
or U10219 (N_10219,N_9617,N_9930);
and U10220 (N_10220,N_9575,N_9794);
or U10221 (N_10221,N_9838,N_9810);
or U10222 (N_10222,N_9883,N_9995);
and U10223 (N_10223,N_9715,N_9706);
nand U10224 (N_10224,N_9877,N_9506);
nand U10225 (N_10225,N_9840,N_9846);
or U10226 (N_10226,N_9852,N_9518);
or U10227 (N_10227,N_9970,N_9872);
and U10228 (N_10228,N_9562,N_9708);
and U10229 (N_10229,N_9957,N_9659);
nand U10230 (N_10230,N_9611,N_9966);
or U10231 (N_10231,N_9938,N_9719);
or U10232 (N_10232,N_9808,N_9987);
nor U10233 (N_10233,N_9599,N_9660);
nor U10234 (N_10234,N_9939,N_9500);
or U10235 (N_10235,N_9931,N_9878);
and U10236 (N_10236,N_9525,N_9965);
or U10237 (N_10237,N_9667,N_9884);
nor U10238 (N_10238,N_9671,N_9903);
and U10239 (N_10239,N_9696,N_9540);
xnor U10240 (N_10240,N_9894,N_9511);
and U10241 (N_10241,N_9588,N_9636);
nand U10242 (N_10242,N_9861,N_9700);
nor U10243 (N_10243,N_9581,N_9875);
or U10244 (N_10244,N_9641,N_9649);
and U10245 (N_10245,N_9912,N_9751);
and U10246 (N_10246,N_9936,N_9630);
nor U10247 (N_10247,N_9572,N_9593);
or U10248 (N_10248,N_9628,N_9607);
or U10249 (N_10249,N_9643,N_9892);
and U10250 (N_10250,N_9845,N_9921);
and U10251 (N_10251,N_9938,N_9779);
and U10252 (N_10252,N_9709,N_9822);
nand U10253 (N_10253,N_9809,N_9504);
xor U10254 (N_10254,N_9829,N_9520);
nand U10255 (N_10255,N_9787,N_9518);
nor U10256 (N_10256,N_9643,N_9762);
xnor U10257 (N_10257,N_9778,N_9621);
nand U10258 (N_10258,N_9870,N_9947);
and U10259 (N_10259,N_9856,N_9812);
or U10260 (N_10260,N_9945,N_9633);
or U10261 (N_10261,N_9748,N_9854);
nand U10262 (N_10262,N_9840,N_9671);
nor U10263 (N_10263,N_9842,N_9883);
nand U10264 (N_10264,N_9950,N_9668);
nand U10265 (N_10265,N_9905,N_9860);
nand U10266 (N_10266,N_9942,N_9976);
and U10267 (N_10267,N_9604,N_9839);
nand U10268 (N_10268,N_9725,N_9926);
or U10269 (N_10269,N_9824,N_9614);
or U10270 (N_10270,N_9682,N_9747);
nor U10271 (N_10271,N_9993,N_9543);
nand U10272 (N_10272,N_9501,N_9549);
and U10273 (N_10273,N_9661,N_9933);
nand U10274 (N_10274,N_9638,N_9802);
nor U10275 (N_10275,N_9671,N_9905);
and U10276 (N_10276,N_9827,N_9548);
and U10277 (N_10277,N_9732,N_9746);
nor U10278 (N_10278,N_9717,N_9718);
or U10279 (N_10279,N_9564,N_9622);
and U10280 (N_10280,N_9682,N_9533);
and U10281 (N_10281,N_9997,N_9698);
or U10282 (N_10282,N_9745,N_9645);
nand U10283 (N_10283,N_9580,N_9738);
nand U10284 (N_10284,N_9564,N_9985);
or U10285 (N_10285,N_9554,N_9882);
or U10286 (N_10286,N_9734,N_9977);
or U10287 (N_10287,N_9745,N_9572);
or U10288 (N_10288,N_9925,N_9644);
and U10289 (N_10289,N_9675,N_9565);
nor U10290 (N_10290,N_9834,N_9590);
xnor U10291 (N_10291,N_9932,N_9842);
xor U10292 (N_10292,N_9995,N_9566);
and U10293 (N_10293,N_9627,N_9644);
nand U10294 (N_10294,N_9879,N_9504);
or U10295 (N_10295,N_9643,N_9716);
nand U10296 (N_10296,N_9549,N_9780);
xnor U10297 (N_10297,N_9740,N_9794);
nor U10298 (N_10298,N_9772,N_9579);
nand U10299 (N_10299,N_9639,N_9826);
nand U10300 (N_10300,N_9560,N_9799);
and U10301 (N_10301,N_9907,N_9512);
nor U10302 (N_10302,N_9948,N_9752);
and U10303 (N_10303,N_9837,N_9858);
and U10304 (N_10304,N_9645,N_9844);
nand U10305 (N_10305,N_9711,N_9927);
and U10306 (N_10306,N_9938,N_9531);
and U10307 (N_10307,N_9859,N_9683);
nand U10308 (N_10308,N_9511,N_9566);
nand U10309 (N_10309,N_9630,N_9995);
nor U10310 (N_10310,N_9530,N_9570);
or U10311 (N_10311,N_9772,N_9866);
nand U10312 (N_10312,N_9960,N_9595);
and U10313 (N_10313,N_9666,N_9713);
nand U10314 (N_10314,N_9967,N_9535);
xor U10315 (N_10315,N_9608,N_9963);
nor U10316 (N_10316,N_9918,N_9956);
xor U10317 (N_10317,N_9592,N_9575);
or U10318 (N_10318,N_9811,N_9698);
nand U10319 (N_10319,N_9532,N_9951);
nand U10320 (N_10320,N_9729,N_9826);
or U10321 (N_10321,N_9844,N_9874);
nor U10322 (N_10322,N_9949,N_9827);
nor U10323 (N_10323,N_9746,N_9587);
nand U10324 (N_10324,N_9769,N_9600);
nor U10325 (N_10325,N_9967,N_9598);
and U10326 (N_10326,N_9624,N_9617);
nor U10327 (N_10327,N_9719,N_9766);
nor U10328 (N_10328,N_9698,N_9845);
or U10329 (N_10329,N_9736,N_9868);
and U10330 (N_10330,N_9573,N_9970);
nand U10331 (N_10331,N_9574,N_9778);
nand U10332 (N_10332,N_9906,N_9853);
and U10333 (N_10333,N_9994,N_9551);
and U10334 (N_10334,N_9710,N_9672);
xnor U10335 (N_10335,N_9532,N_9735);
nand U10336 (N_10336,N_9956,N_9779);
xnor U10337 (N_10337,N_9849,N_9934);
nor U10338 (N_10338,N_9668,N_9657);
or U10339 (N_10339,N_9503,N_9922);
nand U10340 (N_10340,N_9531,N_9797);
nor U10341 (N_10341,N_9719,N_9777);
and U10342 (N_10342,N_9962,N_9807);
nand U10343 (N_10343,N_9613,N_9765);
nor U10344 (N_10344,N_9867,N_9650);
nor U10345 (N_10345,N_9941,N_9876);
nor U10346 (N_10346,N_9525,N_9822);
nand U10347 (N_10347,N_9535,N_9889);
and U10348 (N_10348,N_9723,N_9761);
and U10349 (N_10349,N_9578,N_9558);
or U10350 (N_10350,N_9570,N_9773);
nand U10351 (N_10351,N_9958,N_9680);
or U10352 (N_10352,N_9932,N_9887);
and U10353 (N_10353,N_9559,N_9981);
xor U10354 (N_10354,N_9983,N_9587);
nand U10355 (N_10355,N_9896,N_9745);
and U10356 (N_10356,N_9813,N_9975);
or U10357 (N_10357,N_9517,N_9947);
nor U10358 (N_10358,N_9987,N_9834);
nand U10359 (N_10359,N_9649,N_9595);
and U10360 (N_10360,N_9533,N_9620);
nand U10361 (N_10361,N_9712,N_9663);
or U10362 (N_10362,N_9968,N_9940);
nand U10363 (N_10363,N_9782,N_9973);
nand U10364 (N_10364,N_9792,N_9780);
nand U10365 (N_10365,N_9806,N_9827);
nor U10366 (N_10366,N_9791,N_9721);
and U10367 (N_10367,N_9573,N_9734);
or U10368 (N_10368,N_9736,N_9925);
xor U10369 (N_10369,N_9608,N_9839);
or U10370 (N_10370,N_9536,N_9868);
nand U10371 (N_10371,N_9799,N_9819);
nand U10372 (N_10372,N_9764,N_9731);
nor U10373 (N_10373,N_9990,N_9638);
xor U10374 (N_10374,N_9536,N_9599);
xnor U10375 (N_10375,N_9515,N_9864);
nand U10376 (N_10376,N_9695,N_9614);
and U10377 (N_10377,N_9987,N_9641);
nor U10378 (N_10378,N_9873,N_9951);
and U10379 (N_10379,N_9620,N_9695);
nand U10380 (N_10380,N_9779,N_9623);
nand U10381 (N_10381,N_9563,N_9616);
or U10382 (N_10382,N_9665,N_9958);
nand U10383 (N_10383,N_9971,N_9860);
nand U10384 (N_10384,N_9595,N_9974);
nand U10385 (N_10385,N_9784,N_9774);
nor U10386 (N_10386,N_9500,N_9813);
nor U10387 (N_10387,N_9521,N_9505);
or U10388 (N_10388,N_9540,N_9520);
nor U10389 (N_10389,N_9889,N_9532);
or U10390 (N_10390,N_9997,N_9616);
and U10391 (N_10391,N_9784,N_9766);
and U10392 (N_10392,N_9852,N_9808);
nand U10393 (N_10393,N_9935,N_9743);
or U10394 (N_10394,N_9640,N_9678);
and U10395 (N_10395,N_9963,N_9911);
nand U10396 (N_10396,N_9557,N_9842);
nand U10397 (N_10397,N_9870,N_9514);
xnor U10398 (N_10398,N_9603,N_9819);
or U10399 (N_10399,N_9859,N_9570);
nor U10400 (N_10400,N_9807,N_9775);
nand U10401 (N_10401,N_9755,N_9828);
xnor U10402 (N_10402,N_9520,N_9803);
xor U10403 (N_10403,N_9726,N_9613);
nor U10404 (N_10404,N_9902,N_9928);
nor U10405 (N_10405,N_9780,N_9512);
nor U10406 (N_10406,N_9995,N_9803);
nor U10407 (N_10407,N_9834,N_9859);
and U10408 (N_10408,N_9914,N_9616);
nand U10409 (N_10409,N_9991,N_9857);
nand U10410 (N_10410,N_9782,N_9858);
and U10411 (N_10411,N_9936,N_9538);
or U10412 (N_10412,N_9656,N_9954);
nand U10413 (N_10413,N_9841,N_9806);
and U10414 (N_10414,N_9799,N_9771);
nand U10415 (N_10415,N_9766,N_9874);
nand U10416 (N_10416,N_9929,N_9711);
nor U10417 (N_10417,N_9906,N_9612);
or U10418 (N_10418,N_9561,N_9680);
nor U10419 (N_10419,N_9524,N_9540);
nand U10420 (N_10420,N_9543,N_9720);
nor U10421 (N_10421,N_9727,N_9508);
nand U10422 (N_10422,N_9740,N_9772);
nand U10423 (N_10423,N_9501,N_9551);
or U10424 (N_10424,N_9508,N_9891);
nand U10425 (N_10425,N_9752,N_9643);
and U10426 (N_10426,N_9828,N_9843);
and U10427 (N_10427,N_9761,N_9638);
or U10428 (N_10428,N_9741,N_9885);
or U10429 (N_10429,N_9524,N_9991);
or U10430 (N_10430,N_9959,N_9594);
nor U10431 (N_10431,N_9683,N_9869);
xnor U10432 (N_10432,N_9843,N_9990);
nand U10433 (N_10433,N_9990,N_9816);
nand U10434 (N_10434,N_9754,N_9717);
or U10435 (N_10435,N_9590,N_9910);
nor U10436 (N_10436,N_9852,N_9578);
xor U10437 (N_10437,N_9751,N_9899);
xor U10438 (N_10438,N_9807,N_9662);
or U10439 (N_10439,N_9670,N_9981);
or U10440 (N_10440,N_9733,N_9507);
or U10441 (N_10441,N_9812,N_9977);
nand U10442 (N_10442,N_9889,N_9758);
nor U10443 (N_10443,N_9598,N_9998);
nor U10444 (N_10444,N_9791,N_9884);
or U10445 (N_10445,N_9868,N_9708);
or U10446 (N_10446,N_9606,N_9620);
or U10447 (N_10447,N_9962,N_9984);
or U10448 (N_10448,N_9831,N_9807);
nor U10449 (N_10449,N_9809,N_9679);
and U10450 (N_10450,N_9903,N_9927);
and U10451 (N_10451,N_9551,N_9620);
nor U10452 (N_10452,N_9664,N_9611);
or U10453 (N_10453,N_9791,N_9764);
nor U10454 (N_10454,N_9646,N_9742);
or U10455 (N_10455,N_9638,N_9819);
nor U10456 (N_10456,N_9834,N_9511);
nand U10457 (N_10457,N_9815,N_9517);
or U10458 (N_10458,N_9841,N_9681);
and U10459 (N_10459,N_9687,N_9792);
or U10460 (N_10460,N_9905,N_9501);
or U10461 (N_10461,N_9595,N_9650);
nor U10462 (N_10462,N_9983,N_9586);
and U10463 (N_10463,N_9879,N_9696);
and U10464 (N_10464,N_9530,N_9971);
nand U10465 (N_10465,N_9974,N_9626);
or U10466 (N_10466,N_9857,N_9977);
or U10467 (N_10467,N_9646,N_9782);
and U10468 (N_10468,N_9688,N_9844);
nor U10469 (N_10469,N_9945,N_9988);
xor U10470 (N_10470,N_9799,N_9997);
xor U10471 (N_10471,N_9543,N_9662);
nand U10472 (N_10472,N_9554,N_9731);
nor U10473 (N_10473,N_9712,N_9594);
xnor U10474 (N_10474,N_9881,N_9686);
and U10475 (N_10475,N_9608,N_9517);
or U10476 (N_10476,N_9829,N_9529);
nand U10477 (N_10477,N_9959,N_9944);
or U10478 (N_10478,N_9715,N_9763);
and U10479 (N_10479,N_9533,N_9959);
or U10480 (N_10480,N_9642,N_9820);
or U10481 (N_10481,N_9872,N_9783);
or U10482 (N_10482,N_9505,N_9823);
nand U10483 (N_10483,N_9628,N_9765);
nand U10484 (N_10484,N_9981,N_9775);
nand U10485 (N_10485,N_9942,N_9925);
xor U10486 (N_10486,N_9813,N_9883);
and U10487 (N_10487,N_9693,N_9571);
and U10488 (N_10488,N_9814,N_9968);
nand U10489 (N_10489,N_9880,N_9842);
nor U10490 (N_10490,N_9868,N_9607);
xor U10491 (N_10491,N_9990,N_9742);
and U10492 (N_10492,N_9713,N_9832);
and U10493 (N_10493,N_9899,N_9538);
and U10494 (N_10494,N_9931,N_9951);
xor U10495 (N_10495,N_9785,N_9815);
xnor U10496 (N_10496,N_9932,N_9890);
nor U10497 (N_10497,N_9538,N_9575);
or U10498 (N_10498,N_9772,N_9836);
or U10499 (N_10499,N_9865,N_9883);
nand U10500 (N_10500,N_10261,N_10037);
or U10501 (N_10501,N_10244,N_10157);
or U10502 (N_10502,N_10181,N_10375);
and U10503 (N_10503,N_10409,N_10014);
or U10504 (N_10504,N_10015,N_10373);
and U10505 (N_10505,N_10253,N_10263);
nand U10506 (N_10506,N_10092,N_10477);
and U10507 (N_10507,N_10210,N_10004);
nand U10508 (N_10508,N_10038,N_10208);
and U10509 (N_10509,N_10107,N_10403);
and U10510 (N_10510,N_10483,N_10449);
nor U10511 (N_10511,N_10492,N_10164);
nand U10512 (N_10512,N_10350,N_10182);
nand U10513 (N_10513,N_10448,N_10174);
nor U10514 (N_10514,N_10133,N_10006);
or U10515 (N_10515,N_10021,N_10200);
nor U10516 (N_10516,N_10335,N_10034);
and U10517 (N_10517,N_10411,N_10194);
nand U10518 (N_10518,N_10433,N_10463);
or U10519 (N_10519,N_10240,N_10281);
xnor U10520 (N_10520,N_10090,N_10159);
nand U10521 (N_10521,N_10291,N_10156);
nor U10522 (N_10522,N_10239,N_10029);
nor U10523 (N_10523,N_10176,N_10017);
nand U10524 (N_10524,N_10348,N_10255);
nand U10525 (N_10525,N_10051,N_10191);
and U10526 (N_10526,N_10259,N_10074);
xnor U10527 (N_10527,N_10079,N_10270);
xnor U10528 (N_10528,N_10457,N_10438);
nand U10529 (N_10529,N_10163,N_10356);
nand U10530 (N_10530,N_10179,N_10086);
and U10531 (N_10531,N_10394,N_10172);
and U10532 (N_10532,N_10072,N_10190);
nand U10533 (N_10533,N_10264,N_10301);
and U10534 (N_10534,N_10213,N_10115);
nand U10535 (N_10535,N_10130,N_10272);
nand U10536 (N_10536,N_10066,N_10258);
or U10537 (N_10537,N_10078,N_10286);
or U10538 (N_10538,N_10168,N_10305);
or U10539 (N_10539,N_10265,N_10040);
nor U10540 (N_10540,N_10376,N_10170);
nand U10541 (N_10541,N_10486,N_10318);
nor U10542 (N_10542,N_10118,N_10207);
and U10543 (N_10543,N_10032,N_10413);
nand U10544 (N_10544,N_10227,N_10439);
and U10545 (N_10545,N_10285,N_10494);
nand U10546 (N_10546,N_10059,N_10333);
or U10547 (N_10547,N_10219,N_10363);
xor U10548 (N_10548,N_10161,N_10322);
or U10549 (N_10549,N_10440,N_10251);
and U10550 (N_10550,N_10381,N_10497);
nand U10551 (N_10551,N_10472,N_10035);
nand U10552 (N_10552,N_10016,N_10343);
nand U10553 (N_10553,N_10382,N_10071);
and U10554 (N_10554,N_10248,N_10231);
and U10555 (N_10555,N_10186,N_10052);
nor U10556 (N_10556,N_10332,N_10150);
nand U10557 (N_10557,N_10204,N_10111);
and U10558 (N_10558,N_10142,N_10341);
and U10559 (N_10559,N_10018,N_10392);
nand U10560 (N_10560,N_10482,N_10456);
or U10561 (N_10561,N_10247,N_10279);
or U10562 (N_10562,N_10184,N_10027);
nand U10563 (N_10563,N_10033,N_10412);
nor U10564 (N_10564,N_10276,N_10422);
nand U10565 (N_10565,N_10103,N_10427);
nand U10566 (N_10566,N_10235,N_10093);
nand U10567 (N_10567,N_10102,N_10061);
xnor U10568 (N_10568,N_10464,N_10473);
or U10569 (N_10569,N_10479,N_10455);
nand U10570 (N_10570,N_10096,N_10269);
and U10571 (N_10571,N_10330,N_10387);
nand U10572 (N_10572,N_10154,N_10402);
nand U10573 (N_10573,N_10271,N_10222);
nand U10574 (N_10574,N_10368,N_10105);
nor U10575 (N_10575,N_10396,N_10389);
nor U10576 (N_10576,N_10432,N_10019);
xnor U10577 (N_10577,N_10081,N_10273);
or U10578 (N_10578,N_10198,N_10048);
nor U10579 (N_10579,N_10405,N_10178);
xor U10580 (N_10580,N_10050,N_10056);
or U10581 (N_10581,N_10012,N_10075);
xnor U10582 (N_10582,N_10446,N_10275);
nand U10583 (N_10583,N_10095,N_10094);
nor U10584 (N_10584,N_10311,N_10223);
xnor U10585 (N_10585,N_10408,N_10236);
xor U10586 (N_10586,N_10024,N_10380);
or U10587 (N_10587,N_10100,N_10212);
or U10588 (N_10588,N_10199,N_10119);
or U10589 (N_10589,N_10462,N_10460);
nand U10590 (N_10590,N_10484,N_10196);
nor U10591 (N_10591,N_10359,N_10496);
and U10592 (N_10592,N_10302,N_10453);
or U10593 (N_10593,N_10023,N_10042);
nand U10594 (N_10594,N_10237,N_10087);
nand U10595 (N_10595,N_10390,N_10209);
xor U10596 (N_10596,N_10310,N_10445);
xnor U10597 (N_10597,N_10011,N_10233);
or U10598 (N_10598,N_10076,N_10030);
and U10599 (N_10599,N_10287,N_10141);
nor U10600 (N_10600,N_10476,N_10431);
nor U10601 (N_10601,N_10088,N_10461);
nor U10602 (N_10602,N_10364,N_10321);
and U10603 (N_10603,N_10342,N_10481);
or U10604 (N_10604,N_10399,N_10124);
and U10605 (N_10605,N_10299,N_10465);
or U10606 (N_10606,N_10041,N_10160);
and U10607 (N_10607,N_10327,N_10139);
or U10608 (N_10608,N_10063,N_10282);
nand U10609 (N_10609,N_10358,N_10224);
or U10610 (N_10610,N_10151,N_10315);
nand U10611 (N_10611,N_10337,N_10135);
or U10612 (N_10612,N_10426,N_10188);
nand U10613 (N_10613,N_10371,N_10379);
xnor U10614 (N_10614,N_10314,N_10417);
and U10615 (N_10615,N_10468,N_10183);
nand U10616 (N_10616,N_10101,N_10128);
nand U10617 (N_10617,N_10296,N_10120);
nor U10618 (N_10618,N_10297,N_10067);
nand U10619 (N_10619,N_10158,N_10490);
nand U10620 (N_10620,N_10000,N_10429);
or U10621 (N_10621,N_10372,N_10498);
and U10622 (N_10622,N_10044,N_10425);
and U10623 (N_10623,N_10336,N_10127);
or U10624 (N_10624,N_10357,N_10054);
or U10625 (N_10625,N_10298,N_10008);
and U10626 (N_10626,N_10295,N_10386);
or U10627 (N_10627,N_10406,N_10121);
nor U10628 (N_10628,N_10062,N_10444);
or U10629 (N_10629,N_10442,N_10113);
nand U10630 (N_10630,N_10416,N_10126);
or U10631 (N_10631,N_10149,N_10189);
and U10632 (N_10632,N_10278,N_10435);
xnor U10633 (N_10633,N_10307,N_10117);
and U10634 (N_10634,N_10393,N_10122);
nor U10635 (N_10635,N_10424,N_10436);
or U10636 (N_10636,N_10192,N_10397);
nand U10637 (N_10637,N_10478,N_10137);
or U10638 (N_10638,N_10419,N_10098);
and U10639 (N_10639,N_10414,N_10331);
or U10640 (N_10640,N_10242,N_10277);
nand U10641 (N_10641,N_10060,N_10216);
or U10642 (N_10642,N_10138,N_10404);
or U10643 (N_10643,N_10312,N_10306);
and U10644 (N_10644,N_10131,N_10329);
nand U10645 (N_10645,N_10116,N_10171);
xnor U10646 (N_10646,N_10401,N_10423);
xor U10647 (N_10647,N_10441,N_10084);
nand U10648 (N_10648,N_10334,N_10153);
and U10649 (N_10649,N_10046,N_10064);
nor U10650 (N_10650,N_10474,N_10313);
and U10651 (N_10651,N_10352,N_10262);
xnor U10652 (N_10652,N_10268,N_10303);
and U10653 (N_10653,N_10220,N_10488);
nand U10654 (N_10654,N_10114,N_10089);
nand U10655 (N_10655,N_10215,N_10136);
nand U10656 (N_10656,N_10452,N_10443);
nand U10657 (N_10657,N_10290,N_10230);
nand U10658 (N_10658,N_10185,N_10099);
nand U10659 (N_10659,N_10288,N_10470);
nor U10660 (N_10660,N_10005,N_10053);
nor U10661 (N_10661,N_10328,N_10324);
nor U10662 (N_10662,N_10140,N_10245);
xor U10663 (N_10663,N_10058,N_10437);
and U10664 (N_10664,N_10001,N_10471);
nor U10665 (N_10665,N_10144,N_10069);
nand U10666 (N_10666,N_10274,N_10246);
nor U10667 (N_10667,N_10355,N_10266);
nor U10668 (N_10668,N_10447,N_10317);
nand U10669 (N_10669,N_10003,N_10395);
xor U10670 (N_10670,N_10203,N_10234);
nand U10671 (N_10671,N_10085,N_10284);
nand U10672 (N_10672,N_10345,N_10205);
nand U10673 (N_10673,N_10292,N_10323);
or U10674 (N_10674,N_10077,N_10145);
or U10675 (N_10675,N_10057,N_10031);
and U10676 (N_10676,N_10022,N_10028);
nor U10677 (N_10677,N_10489,N_10070);
and U10678 (N_10678,N_10112,N_10289);
and U10679 (N_10679,N_10354,N_10083);
nand U10680 (N_10680,N_10421,N_10206);
and U10681 (N_10681,N_10073,N_10211);
nor U10682 (N_10682,N_10214,N_10132);
nor U10683 (N_10683,N_10420,N_10434);
nor U10684 (N_10684,N_10459,N_10495);
nor U10685 (N_10685,N_10383,N_10361);
nand U10686 (N_10686,N_10045,N_10458);
or U10687 (N_10687,N_10026,N_10293);
or U10688 (N_10688,N_10047,N_10400);
nand U10689 (N_10689,N_10466,N_10043);
nand U10690 (N_10690,N_10377,N_10167);
or U10691 (N_10691,N_10049,N_10347);
and U10692 (N_10692,N_10475,N_10039);
or U10693 (N_10693,N_10097,N_10487);
nand U10694 (N_10694,N_10294,N_10002);
nand U10695 (N_10695,N_10110,N_10454);
or U10696 (N_10696,N_10080,N_10225);
nor U10697 (N_10697,N_10250,N_10106);
nand U10698 (N_10698,N_10491,N_10065);
or U10699 (N_10699,N_10148,N_10418);
nor U10700 (N_10700,N_10344,N_10316);
xor U10701 (N_10701,N_10013,N_10228);
nor U10702 (N_10702,N_10283,N_10351);
nand U10703 (N_10703,N_10369,N_10091);
or U10704 (N_10704,N_10415,N_10055);
nand U10705 (N_10705,N_10257,N_10195);
or U10706 (N_10706,N_10391,N_10353);
and U10707 (N_10707,N_10267,N_10143);
nand U10708 (N_10708,N_10256,N_10025);
or U10709 (N_10709,N_10147,N_10346);
or U10710 (N_10710,N_10485,N_10338);
or U10711 (N_10711,N_10134,N_10340);
nor U10712 (N_10712,N_10155,N_10428);
nor U10713 (N_10713,N_10365,N_10180);
nand U10714 (N_10714,N_10319,N_10374);
xor U10715 (N_10715,N_10010,N_10469);
nand U10716 (N_10716,N_10109,N_10173);
nor U10717 (N_10717,N_10202,N_10304);
nand U10718 (N_10718,N_10249,N_10349);
or U10719 (N_10719,N_10125,N_10229);
nand U10720 (N_10720,N_10398,N_10165);
and U10721 (N_10721,N_10187,N_10260);
xor U10722 (N_10722,N_10450,N_10036);
nor U10723 (N_10723,N_10238,N_10384);
nor U10724 (N_10724,N_10366,N_10326);
nand U10725 (N_10725,N_10221,N_10123);
nor U10726 (N_10726,N_10082,N_10241);
or U10727 (N_10727,N_10388,N_10360);
or U10728 (N_10728,N_10308,N_10104);
nor U10729 (N_10729,N_10020,N_10177);
and U10730 (N_10730,N_10152,N_10320);
nand U10731 (N_10731,N_10339,N_10309);
or U10732 (N_10732,N_10370,N_10362);
or U10733 (N_10733,N_10166,N_10280);
nor U10734 (N_10734,N_10108,N_10009);
nor U10735 (N_10735,N_10378,N_10367);
nor U10736 (N_10736,N_10243,N_10226);
or U10737 (N_10737,N_10197,N_10325);
and U10738 (N_10738,N_10169,N_10499);
and U10739 (N_10739,N_10068,N_10451);
nor U10740 (N_10740,N_10480,N_10300);
and U10741 (N_10741,N_10193,N_10385);
and U10742 (N_10742,N_10129,N_10467);
nor U10743 (N_10743,N_10252,N_10232);
nor U10744 (N_10744,N_10162,N_10254);
and U10745 (N_10745,N_10493,N_10175);
or U10746 (N_10746,N_10218,N_10146);
nor U10747 (N_10747,N_10201,N_10407);
or U10748 (N_10748,N_10410,N_10430);
or U10749 (N_10749,N_10007,N_10217);
nand U10750 (N_10750,N_10230,N_10292);
or U10751 (N_10751,N_10468,N_10403);
xor U10752 (N_10752,N_10279,N_10036);
or U10753 (N_10753,N_10386,N_10441);
or U10754 (N_10754,N_10449,N_10054);
or U10755 (N_10755,N_10073,N_10155);
or U10756 (N_10756,N_10149,N_10357);
nand U10757 (N_10757,N_10482,N_10214);
or U10758 (N_10758,N_10312,N_10372);
and U10759 (N_10759,N_10068,N_10030);
and U10760 (N_10760,N_10340,N_10099);
xnor U10761 (N_10761,N_10380,N_10033);
nand U10762 (N_10762,N_10482,N_10006);
and U10763 (N_10763,N_10068,N_10463);
and U10764 (N_10764,N_10023,N_10265);
nand U10765 (N_10765,N_10150,N_10096);
or U10766 (N_10766,N_10475,N_10089);
xnor U10767 (N_10767,N_10004,N_10271);
nor U10768 (N_10768,N_10497,N_10214);
nor U10769 (N_10769,N_10225,N_10159);
nor U10770 (N_10770,N_10447,N_10229);
or U10771 (N_10771,N_10224,N_10095);
and U10772 (N_10772,N_10383,N_10268);
nor U10773 (N_10773,N_10334,N_10381);
nand U10774 (N_10774,N_10338,N_10499);
and U10775 (N_10775,N_10264,N_10367);
or U10776 (N_10776,N_10391,N_10360);
nand U10777 (N_10777,N_10473,N_10395);
xor U10778 (N_10778,N_10157,N_10336);
or U10779 (N_10779,N_10124,N_10233);
or U10780 (N_10780,N_10469,N_10098);
or U10781 (N_10781,N_10212,N_10222);
and U10782 (N_10782,N_10283,N_10318);
or U10783 (N_10783,N_10059,N_10361);
and U10784 (N_10784,N_10171,N_10497);
nor U10785 (N_10785,N_10400,N_10467);
xnor U10786 (N_10786,N_10234,N_10180);
or U10787 (N_10787,N_10038,N_10062);
nor U10788 (N_10788,N_10016,N_10456);
and U10789 (N_10789,N_10338,N_10473);
nand U10790 (N_10790,N_10444,N_10460);
nor U10791 (N_10791,N_10226,N_10317);
nand U10792 (N_10792,N_10082,N_10441);
or U10793 (N_10793,N_10377,N_10141);
or U10794 (N_10794,N_10276,N_10368);
nand U10795 (N_10795,N_10096,N_10442);
nand U10796 (N_10796,N_10374,N_10266);
or U10797 (N_10797,N_10251,N_10082);
nor U10798 (N_10798,N_10053,N_10395);
nor U10799 (N_10799,N_10394,N_10150);
and U10800 (N_10800,N_10208,N_10026);
and U10801 (N_10801,N_10012,N_10234);
nor U10802 (N_10802,N_10103,N_10419);
or U10803 (N_10803,N_10086,N_10404);
nand U10804 (N_10804,N_10377,N_10283);
xor U10805 (N_10805,N_10186,N_10298);
or U10806 (N_10806,N_10089,N_10100);
xnor U10807 (N_10807,N_10454,N_10093);
nor U10808 (N_10808,N_10191,N_10336);
or U10809 (N_10809,N_10061,N_10063);
or U10810 (N_10810,N_10272,N_10134);
or U10811 (N_10811,N_10347,N_10419);
or U10812 (N_10812,N_10037,N_10004);
xnor U10813 (N_10813,N_10381,N_10402);
xnor U10814 (N_10814,N_10214,N_10136);
nor U10815 (N_10815,N_10373,N_10424);
nor U10816 (N_10816,N_10497,N_10164);
and U10817 (N_10817,N_10194,N_10068);
or U10818 (N_10818,N_10440,N_10448);
and U10819 (N_10819,N_10206,N_10070);
and U10820 (N_10820,N_10155,N_10109);
and U10821 (N_10821,N_10235,N_10462);
or U10822 (N_10822,N_10027,N_10223);
nand U10823 (N_10823,N_10490,N_10209);
nor U10824 (N_10824,N_10283,N_10053);
and U10825 (N_10825,N_10124,N_10025);
and U10826 (N_10826,N_10026,N_10373);
nor U10827 (N_10827,N_10063,N_10227);
nor U10828 (N_10828,N_10171,N_10247);
xnor U10829 (N_10829,N_10364,N_10429);
nor U10830 (N_10830,N_10048,N_10023);
nand U10831 (N_10831,N_10487,N_10204);
xor U10832 (N_10832,N_10419,N_10384);
nand U10833 (N_10833,N_10203,N_10362);
nand U10834 (N_10834,N_10261,N_10051);
nor U10835 (N_10835,N_10201,N_10062);
and U10836 (N_10836,N_10163,N_10373);
nor U10837 (N_10837,N_10475,N_10390);
nand U10838 (N_10838,N_10300,N_10243);
nand U10839 (N_10839,N_10354,N_10487);
and U10840 (N_10840,N_10434,N_10153);
or U10841 (N_10841,N_10234,N_10182);
xnor U10842 (N_10842,N_10305,N_10002);
nor U10843 (N_10843,N_10265,N_10064);
xnor U10844 (N_10844,N_10259,N_10078);
or U10845 (N_10845,N_10158,N_10389);
nor U10846 (N_10846,N_10156,N_10490);
nor U10847 (N_10847,N_10285,N_10430);
nor U10848 (N_10848,N_10206,N_10128);
and U10849 (N_10849,N_10061,N_10431);
nor U10850 (N_10850,N_10247,N_10278);
and U10851 (N_10851,N_10290,N_10434);
nor U10852 (N_10852,N_10461,N_10205);
nand U10853 (N_10853,N_10373,N_10346);
nand U10854 (N_10854,N_10445,N_10431);
and U10855 (N_10855,N_10488,N_10251);
or U10856 (N_10856,N_10299,N_10245);
and U10857 (N_10857,N_10222,N_10319);
xor U10858 (N_10858,N_10082,N_10173);
nor U10859 (N_10859,N_10290,N_10300);
and U10860 (N_10860,N_10385,N_10400);
nand U10861 (N_10861,N_10140,N_10125);
nor U10862 (N_10862,N_10309,N_10490);
xnor U10863 (N_10863,N_10378,N_10370);
or U10864 (N_10864,N_10258,N_10159);
nand U10865 (N_10865,N_10337,N_10191);
nand U10866 (N_10866,N_10047,N_10436);
or U10867 (N_10867,N_10456,N_10196);
nor U10868 (N_10868,N_10247,N_10465);
nor U10869 (N_10869,N_10258,N_10031);
nor U10870 (N_10870,N_10337,N_10078);
or U10871 (N_10871,N_10455,N_10488);
and U10872 (N_10872,N_10035,N_10309);
nand U10873 (N_10873,N_10182,N_10137);
xor U10874 (N_10874,N_10295,N_10312);
nand U10875 (N_10875,N_10056,N_10112);
and U10876 (N_10876,N_10241,N_10254);
nand U10877 (N_10877,N_10141,N_10112);
nand U10878 (N_10878,N_10449,N_10141);
xor U10879 (N_10879,N_10366,N_10404);
nor U10880 (N_10880,N_10409,N_10061);
and U10881 (N_10881,N_10100,N_10131);
nor U10882 (N_10882,N_10225,N_10199);
and U10883 (N_10883,N_10048,N_10292);
nand U10884 (N_10884,N_10306,N_10045);
nand U10885 (N_10885,N_10299,N_10208);
or U10886 (N_10886,N_10278,N_10130);
xnor U10887 (N_10887,N_10373,N_10190);
or U10888 (N_10888,N_10215,N_10244);
or U10889 (N_10889,N_10257,N_10128);
or U10890 (N_10890,N_10384,N_10000);
and U10891 (N_10891,N_10081,N_10142);
nor U10892 (N_10892,N_10254,N_10437);
or U10893 (N_10893,N_10307,N_10131);
nand U10894 (N_10894,N_10159,N_10119);
nand U10895 (N_10895,N_10482,N_10072);
xnor U10896 (N_10896,N_10386,N_10373);
nand U10897 (N_10897,N_10247,N_10495);
and U10898 (N_10898,N_10130,N_10489);
and U10899 (N_10899,N_10029,N_10173);
nand U10900 (N_10900,N_10464,N_10068);
or U10901 (N_10901,N_10256,N_10097);
nor U10902 (N_10902,N_10116,N_10312);
or U10903 (N_10903,N_10127,N_10072);
or U10904 (N_10904,N_10001,N_10052);
or U10905 (N_10905,N_10380,N_10009);
xnor U10906 (N_10906,N_10038,N_10410);
nor U10907 (N_10907,N_10209,N_10105);
nand U10908 (N_10908,N_10211,N_10329);
and U10909 (N_10909,N_10328,N_10023);
and U10910 (N_10910,N_10135,N_10062);
xnor U10911 (N_10911,N_10056,N_10216);
or U10912 (N_10912,N_10001,N_10475);
nand U10913 (N_10913,N_10017,N_10467);
nand U10914 (N_10914,N_10271,N_10202);
and U10915 (N_10915,N_10348,N_10151);
and U10916 (N_10916,N_10151,N_10243);
or U10917 (N_10917,N_10182,N_10470);
nand U10918 (N_10918,N_10050,N_10398);
nor U10919 (N_10919,N_10064,N_10201);
or U10920 (N_10920,N_10422,N_10491);
nand U10921 (N_10921,N_10277,N_10284);
nor U10922 (N_10922,N_10142,N_10492);
and U10923 (N_10923,N_10495,N_10105);
nand U10924 (N_10924,N_10132,N_10061);
and U10925 (N_10925,N_10005,N_10447);
or U10926 (N_10926,N_10422,N_10418);
nor U10927 (N_10927,N_10032,N_10342);
and U10928 (N_10928,N_10487,N_10043);
and U10929 (N_10929,N_10407,N_10094);
nand U10930 (N_10930,N_10190,N_10201);
xor U10931 (N_10931,N_10103,N_10278);
nand U10932 (N_10932,N_10265,N_10151);
nor U10933 (N_10933,N_10241,N_10264);
or U10934 (N_10934,N_10464,N_10446);
or U10935 (N_10935,N_10410,N_10004);
nand U10936 (N_10936,N_10336,N_10294);
xor U10937 (N_10937,N_10370,N_10135);
and U10938 (N_10938,N_10205,N_10231);
and U10939 (N_10939,N_10478,N_10220);
or U10940 (N_10940,N_10245,N_10221);
nor U10941 (N_10941,N_10393,N_10092);
or U10942 (N_10942,N_10212,N_10114);
nor U10943 (N_10943,N_10160,N_10120);
nand U10944 (N_10944,N_10308,N_10106);
and U10945 (N_10945,N_10127,N_10403);
nand U10946 (N_10946,N_10389,N_10277);
xnor U10947 (N_10947,N_10185,N_10333);
xor U10948 (N_10948,N_10214,N_10017);
and U10949 (N_10949,N_10325,N_10238);
nor U10950 (N_10950,N_10340,N_10365);
and U10951 (N_10951,N_10039,N_10376);
or U10952 (N_10952,N_10030,N_10227);
nand U10953 (N_10953,N_10422,N_10473);
and U10954 (N_10954,N_10038,N_10267);
nor U10955 (N_10955,N_10287,N_10046);
nor U10956 (N_10956,N_10331,N_10442);
and U10957 (N_10957,N_10119,N_10208);
and U10958 (N_10958,N_10321,N_10405);
and U10959 (N_10959,N_10411,N_10004);
nor U10960 (N_10960,N_10395,N_10251);
nor U10961 (N_10961,N_10397,N_10448);
nand U10962 (N_10962,N_10157,N_10315);
nor U10963 (N_10963,N_10472,N_10160);
nor U10964 (N_10964,N_10489,N_10394);
xor U10965 (N_10965,N_10210,N_10352);
and U10966 (N_10966,N_10413,N_10156);
or U10967 (N_10967,N_10355,N_10211);
nand U10968 (N_10968,N_10203,N_10005);
nand U10969 (N_10969,N_10228,N_10114);
nand U10970 (N_10970,N_10176,N_10481);
nand U10971 (N_10971,N_10051,N_10119);
xor U10972 (N_10972,N_10347,N_10143);
or U10973 (N_10973,N_10313,N_10116);
or U10974 (N_10974,N_10279,N_10319);
and U10975 (N_10975,N_10400,N_10332);
or U10976 (N_10976,N_10102,N_10119);
xnor U10977 (N_10977,N_10183,N_10302);
nand U10978 (N_10978,N_10246,N_10193);
nor U10979 (N_10979,N_10457,N_10316);
and U10980 (N_10980,N_10320,N_10148);
nand U10981 (N_10981,N_10050,N_10188);
nor U10982 (N_10982,N_10213,N_10465);
and U10983 (N_10983,N_10269,N_10183);
nand U10984 (N_10984,N_10478,N_10328);
nor U10985 (N_10985,N_10241,N_10452);
nor U10986 (N_10986,N_10281,N_10185);
nand U10987 (N_10987,N_10089,N_10367);
nor U10988 (N_10988,N_10027,N_10183);
nor U10989 (N_10989,N_10126,N_10381);
nor U10990 (N_10990,N_10031,N_10305);
xor U10991 (N_10991,N_10099,N_10361);
or U10992 (N_10992,N_10058,N_10453);
nand U10993 (N_10993,N_10314,N_10067);
nor U10994 (N_10994,N_10244,N_10453);
nor U10995 (N_10995,N_10466,N_10287);
nand U10996 (N_10996,N_10104,N_10005);
nor U10997 (N_10997,N_10365,N_10303);
nor U10998 (N_10998,N_10091,N_10477);
or U10999 (N_10999,N_10143,N_10084);
nand U11000 (N_11000,N_10625,N_10907);
nand U11001 (N_11001,N_10796,N_10866);
nor U11002 (N_11002,N_10867,N_10814);
and U11003 (N_11003,N_10777,N_10679);
xnor U11004 (N_11004,N_10649,N_10582);
nand U11005 (N_11005,N_10538,N_10652);
xnor U11006 (N_11006,N_10822,N_10514);
or U11007 (N_11007,N_10779,N_10503);
nand U11008 (N_11008,N_10977,N_10925);
nor U11009 (N_11009,N_10886,N_10921);
nor U11010 (N_11010,N_10601,N_10918);
and U11011 (N_11011,N_10697,N_10539);
nor U11012 (N_11012,N_10726,N_10882);
and U11013 (N_11013,N_10690,N_10781);
and U11014 (N_11014,N_10530,N_10888);
nor U11015 (N_11015,N_10761,N_10670);
and U11016 (N_11016,N_10745,N_10911);
or U11017 (N_11017,N_10688,N_10847);
and U11018 (N_11018,N_10710,N_10759);
and U11019 (N_11019,N_10946,N_10696);
and U11020 (N_11020,N_10893,N_10740);
nand U11021 (N_11021,N_10983,N_10634);
or U11022 (N_11022,N_10692,N_10685);
nor U11023 (N_11023,N_10535,N_10889);
xor U11024 (N_11024,N_10737,N_10532);
and U11025 (N_11025,N_10712,N_10956);
nand U11026 (N_11026,N_10899,N_10747);
or U11027 (N_11027,N_10780,N_10805);
or U11028 (N_11028,N_10678,N_10568);
or U11029 (N_11029,N_10676,N_10730);
and U11030 (N_11030,N_10868,N_10824);
nand U11031 (N_11031,N_10944,N_10701);
and U11032 (N_11032,N_10734,N_10638);
nand U11033 (N_11033,N_10661,N_10536);
and U11034 (N_11034,N_10607,N_10518);
or U11035 (N_11035,N_10579,N_10651);
nand U11036 (N_11036,N_10804,N_10926);
nand U11037 (N_11037,N_10577,N_10799);
and U11038 (N_11038,N_10757,N_10580);
or U11039 (N_11039,N_10520,N_10892);
and U11040 (N_11040,N_10978,N_10994);
nand U11041 (N_11041,N_10974,N_10985);
nand U11042 (N_11042,N_10686,N_10821);
nand U11043 (N_11043,N_10667,N_10820);
nor U11044 (N_11044,N_10852,N_10872);
or U11045 (N_11045,N_10954,N_10675);
nand U11046 (N_11046,N_10942,N_10961);
nor U11047 (N_11047,N_10873,N_10698);
xor U11048 (N_11048,N_10549,N_10750);
nand U11049 (N_11049,N_10680,N_10602);
nor U11050 (N_11050,N_10880,N_10809);
nand U11051 (N_11051,N_10849,N_10629);
or U11052 (N_11052,N_10548,N_10914);
xor U11053 (N_11053,N_10839,N_10639);
nand U11054 (N_11054,N_10844,N_10608);
or U11055 (N_11055,N_10603,N_10511);
nor U11056 (N_11056,N_10798,N_10795);
nand U11057 (N_11057,N_10711,N_10862);
nor U11058 (N_11058,N_10816,N_10566);
xor U11059 (N_11059,N_10550,N_10807);
nand U11060 (N_11060,N_10560,N_10534);
nor U11061 (N_11061,N_10771,N_10758);
nand U11062 (N_11062,N_10948,N_10653);
or U11063 (N_11063,N_10768,N_10641);
nand U11064 (N_11064,N_10883,N_10968);
nand U11065 (N_11065,N_10973,N_10562);
nand U11066 (N_11066,N_10962,N_10637);
nor U11067 (N_11067,N_10529,N_10501);
nand U11068 (N_11068,N_10903,N_10811);
or U11069 (N_11069,N_10797,N_10885);
nand U11070 (N_11070,N_10735,N_10500);
xor U11071 (N_11071,N_10995,N_10790);
and U11072 (N_11072,N_10674,N_10825);
or U11073 (N_11073,N_10552,N_10663);
and U11074 (N_11074,N_10785,N_10776);
nor U11075 (N_11075,N_10923,N_10632);
nand U11076 (N_11076,N_10664,N_10949);
or U11077 (N_11077,N_10997,N_10991);
nor U11078 (N_11078,N_10722,N_10935);
and U11079 (N_11079,N_10900,N_10633);
nor U11080 (N_11080,N_10871,N_10836);
nand U11081 (N_11081,N_10523,N_10570);
or U11082 (N_11082,N_10681,N_10982);
nor U11083 (N_11083,N_10967,N_10969);
nor U11084 (N_11084,N_10901,N_10541);
and U11085 (N_11085,N_10990,N_10837);
or U11086 (N_11086,N_10604,N_10794);
nor U11087 (N_11087,N_10905,N_10571);
nand U11088 (N_11088,N_10673,N_10908);
or U11089 (N_11089,N_10876,N_10666);
nor U11090 (N_11090,N_10590,N_10615);
or U11091 (N_11091,N_10960,N_10958);
and U11092 (N_11092,N_10829,N_10575);
or U11093 (N_11093,N_10806,N_10766);
and U11094 (N_11094,N_10741,N_10826);
and U11095 (N_11095,N_10861,N_10854);
xor U11096 (N_11096,N_10658,N_10955);
and U11097 (N_11097,N_10965,N_10507);
and U11098 (N_11098,N_10656,N_10999);
nor U11099 (N_11099,N_10537,N_10691);
and U11100 (N_11100,N_10522,N_10917);
nand U11101 (N_11101,N_10650,N_10619);
nor U11102 (N_11102,N_10706,N_10879);
xnor U11103 (N_11103,N_10792,N_10812);
nor U11104 (N_11104,N_10947,N_10838);
and U11105 (N_11105,N_10896,N_10753);
or U11106 (N_11106,N_10736,N_10988);
nand U11107 (N_11107,N_10662,N_10593);
or U11108 (N_11108,N_10751,N_10912);
or U11109 (N_11109,N_10598,N_10599);
nand U11110 (N_11110,N_10509,N_10930);
and U11111 (N_11111,N_10636,N_10906);
or U11112 (N_11112,N_10669,N_10895);
nor U11113 (N_11113,N_10544,N_10927);
nor U11114 (N_11114,N_10841,N_10578);
nand U11115 (N_11115,N_10922,N_10940);
and U11116 (N_11116,N_10966,N_10993);
and U11117 (N_11117,N_10996,N_10800);
or U11118 (N_11118,N_10937,N_10933);
or U11119 (N_11119,N_10920,N_10732);
nand U11120 (N_11120,N_10542,N_10739);
or U11121 (N_11121,N_10729,N_10916);
nand U11122 (N_11122,N_10936,N_10717);
or U11123 (N_11123,N_10764,N_10689);
nand U11124 (N_11124,N_10943,N_10823);
or U11125 (N_11125,N_10835,N_10772);
or U11126 (N_11126,N_10614,N_10787);
or U11127 (N_11127,N_10559,N_10733);
nand U11128 (N_11128,N_10668,N_10953);
nor U11129 (N_11129,N_10611,N_10760);
xor U11130 (N_11130,N_10831,N_10605);
xnor U11131 (N_11131,N_10724,N_10840);
nand U11132 (N_11132,N_10693,N_10517);
or U11133 (N_11133,N_10803,N_10533);
and U11134 (N_11134,N_10778,N_10600);
nor U11135 (N_11135,N_10924,N_10887);
and U11136 (N_11136,N_10624,N_10643);
nor U11137 (N_11137,N_10715,N_10521);
or U11138 (N_11138,N_10718,N_10524);
or U11139 (N_11139,N_10972,N_10526);
and U11140 (N_11140,N_10813,N_10786);
or U11141 (N_11141,N_10865,N_10815);
xnor U11142 (N_11142,N_10870,N_10709);
and U11143 (N_11143,N_10775,N_10738);
and U11144 (N_11144,N_10502,N_10556);
and U11145 (N_11145,N_10762,N_10702);
nand U11146 (N_11146,N_10703,N_10516);
and U11147 (N_11147,N_10657,N_10752);
or U11148 (N_11148,N_10585,N_10725);
nor U11149 (N_11149,N_10642,N_10595);
nor U11150 (N_11150,N_10897,N_10609);
or U11151 (N_11151,N_10976,N_10828);
and U11152 (N_11152,N_10583,N_10881);
nand U11153 (N_11153,N_10700,N_10720);
nor U11154 (N_11154,N_10510,N_10525);
and U11155 (N_11155,N_10856,N_10612);
nand U11156 (N_11156,N_10616,N_10606);
or U11157 (N_11157,N_10627,N_10553);
and U11158 (N_11158,N_10793,N_10596);
or U11159 (N_11159,N_10971,N_10891);
nand U11160 (N_11160,N_10843,N_10864);
nor U11161 (N_11161,N_10572,N_10731);
nor U11162 (N_11162,N_10540,N_10819);
xor U11163 (N_11163,N_10527,N_10555);
nand U11164 (N_11164,N_10992,N_10984);
xor U11165 (N_11165,N_10621,N_10986);
nand U11166 (N_11166,N_10950,N_10817);
nand U11167 (N_11167,N_10512,N_10830);
nand U11168 (N_11168,N_10694,N_10784);
nor U11169 (N_11169,N_10998,N_10554);
or U11170 (N_11170,N_10551,N_10853);
and U11171 (N_11171,N_10716,N_10743);
nor U11172 (N_11172,N_10569,N_10567);
and U11173 (N_11173,N_10928,N_10827);
or U11174 (N_11174,N_10513,N_10589);
nor U11175 (N_11175,N_10810,N_10902);
nor U11176 (N_11176,N_10573,N_10655);
xor U11177 (N_11177,N_10659,N_10874);
xor U11178 (N_11178,N_10845,N_10964);
nand U11179 (N_11179,N_10765,N_10719);
or U11180 (N_11180,N_10519,N_10644);
or U11181 (N_11181,N_10980,N_10576);
and U11182 (N_11182,N_10635,N_10646);
or U11183 (N_11183,N_10660,N_10695);
or U11184 (N_11184,N_10565,N_10707);
and U11185 (N_11185,N_10630,N_10851);
and U11186 (N_11186,N_10588,N_10774);
or U11187 (N_11187,N_10584,N_10699);
nand U11188 (N_11188,N_10528,N_10671);
and U11189 (N_11189,N_10788,N_10531);
or U11190 (N_11190,N_10875,N_10850);
nor U11191 (N_11191,N_10704,N_10989);
or U11192 (N_11192,N_10878,N_10756);
xor U11193 (N_11193,N_10763,N_10773);
or U11194 (N_11194,N_10848,N_10617);
or U11195 (N_11195,N_10504,N_10557);
and U11196 (N_11196,N_10834,N_10620);
and U11197 (N_11197,N_10963,N_10508);
or U11198 (N_11198,N_10648,N_10951);
nand U11199 (N_11199,N_10802,N_10975);
nor U11200 (N_11200,N_10808,N_10842);
nand U11201 (N_11201,N_10769,N_10919);
or U11202 (N_11202,N_10754,N_10592);
nand U11203 (N_11203,N_10505,N_10970);
or U11204 (N_11204,N_10684,N_10884);
nand U11205 (N_11205,N_10654,N_10945);
nor U11206 (N_11206,N_10913,N_10543);
and U11207 (N_11207,N_10742,N_10677);
and U11208 (N_11208,N_10506,N_10755);
or U11209 (N_11209,N_10770,N_10957);
nor U11210 (N_11210,N_10597,N_10858);
or U11211 (N_11211,N_10959,N_10591);
xor U11212 (N_11212,N_10727,N_10791);
nor U11213 (N_11213,N_10744,N_10587);
nor U11214 (N_11214,N_10748,N_10628);
xor U11215 (N_11215,N_10890,N_10941);
or U11216 (N_11216,N_10682,N_10938);
xnor U11217 (N_11217,N_10564,N_10613);
nand U11218 (N_11218,N_10855,N_10952);
nor U11219 (N_11219,N_10647,N_10610);
nand U11220 (N_11220,N_10515,N_10801);
nor U11221 (N_11221,N_10782,N_10909);
or U11222 (N_11222,N_10894,N_10563);
or U11223 (N_11223,N_10713,N_10987);
and U11224 (N_11224,N_10705,N_10846);
and U11225 (N_11225,N_10749,N_10640);
nor U11226 (N_11226,N_10546,N_10586);
nand U11227 (N_11227,N_10618,N_10939);
or U11228 (N_11228,N_10904,N_10687);
and U11229 (N_11229,N_10934,N_10746);
or U11230 (N_11230,N_10832,N_10929);
and U11231 (N_11231,N_10645,N_10721);
or U11232 (N_11232,N_10857,N_10932);
nand U11233 (N_11233,N_10574,N_10860);
nand U11234 (N_11234,N_10783,N_10818);
or U11235 (N_11235,N_10683,N_10558);
nor U11236 (N_11236,N_10931,N_10723);
and U11237 (N_11237,N_10915,N_10622);
and U11238 (N_11238,N_10979,N_10863);
nand U11239 (N_11239,N_10981,N_10547);
nand U11240 (N_11240,N_10714,N_10672);
and U11241 (N_11241,N_10898,N_10708);
nor U11242 (N_11242,N_10626,N_10631);
or U11243 (N_11243,N_10859,N_10833);
and U11244 (N_11244,N_10581,N_10869);
and U11245 (N_11245,N_10561,N_10789);
nand U11246 (N_11246,N_10665,N_10545);
nand U11247 (N_11247,N_10623,N_10910);
nand U11248 (N_11248,N_10767,N_10877);
and U11249 (N_11249,N_10728,N_10594);
nor U11250 (N_11250,N_10618,N_10874);
and U11251 (N_11251,N_10900,N_10949);
nor U11252 (N_11252,N_10722,N_10547);
nor U11253 (N_11253,N_10674,N_10556);
or U11254 (N_11254,N_10780,N_10585);
xor U11255 (N_11255,N_10746,N_10651);
nand U11256 (N_11256,N_10610,N_10756);
xor U11257 (N_11257,N_10629,N_10605);
nor U11258 (N_11258,N_10709,N_10575);
nand U11259 (N_11259,N_10970,N_10882);
or U11260 (N_11260,N_10597,N_10794);
and U11261 (N_11261,N_10960,N_10593);
nand U11262 (N_11262,N_10678,N_10878);
nand U11263 (N_11263,N_10724,N_10789);
and U11264 (N_11264,N_10716,N_10674);
and U11265 (N_11265,N_10619,N_10947);
or U11266 (N_11266,N_10780,N_10610);
nand U11267 (N_11267,N_10768,N_10728);
nand U11268 (N_11268,N_10706,N_10947);
nor U11269 (N_11269,N_10620,N_10841);
xnor U11270 (N_11270,N_10893,N_10661);
xor U11271 (N_11271,N_10726,N_10845);
nor U11272 (N_11272,N_10837,N_10580);
or U11273 (N_11273,N_10538,N_10536);
xor U11274 (N_11274,N_10968,N_10936);
or U11275 (N_11275,N_10996,N_10949);
or U11276 (N_11276,N_10686,N_10667);
xnor U11277 (N_11277,N_10648,N_10791);
and U11278 (N_11278,N_10595,N_10890);
nor U11279 (N_11279,N_10789,N_10785);
or U11280 (N_11280,N_10681,N_10612);
nand U11281 (N_11281,N_10848,N_10504);
and U11282 (N_11282,N_10906,N_10988);
nor U11283 (N_11283,N_10649,N_10611);
xnor U11284 (N_11284,N_10727,N_10558);
nor U11285 (N_11285,N_10830,N_10925);
or U11286 (N_11286,N_10697,N_10771);
or U11287 (N_11287,N_10901,N_10562);
nor U11288 (N_11288,N_10875,N_10992);
nor U11289 (N_11289,N_10776,N_10693);
nand U11290 (N_11290,N_10962,N_10686);
nand U11291 (N_11291,N_10546,N_10633);
and U11292 (N_11292,N_10533,N_10795);
and U11293 (N_11293,N_10502,N_10603);
nor U11294 (N_11294,N_10572,N_10743);
nor U11295 (N_11295,N_10876,N_10668);
or U11296 (N_11296,N_10740,N_10970);
nor U11297 (N_11297,N_10832,N_10562);
or U11298 (N_11298,N_10907,N_10769);
nor U11299 (N_11299,N_10662,N_10501);
nand U11300 (N_11300,N_10816,N_10502);
nand U11301 (N_11301,N_10786,N_10818);
nand U11302 (N_11302,N_10686,N_10793);
or U11303 (N_11303,N_10636,N_10677);
xor U11304 (N_11304,N_10507,N_10961);
nand U11305 (N_11305,N_10804,N_10835);
or U11306 (N_11306,N_10565,N_10544);
or U11307 (N_11307,N_10774,N_10687);
nor U11308 (N_11308,N_10771,N_10619);
nand U11309 (N_11309,N_10914,N_10739);
or U11310 (N_11310,N_10627,N_10763);
or U11311 (N_11311,N_10734,N_10772);
nor U11312 (N_11312,N_10794,N_10584);
nor U11313 (N_11313,N_10960,N_10990);
or U11314 (N_11314,N_10873,N_10547);
nor U11315 (N_11315,N_10742,N_10513);
and U11316 (N_11316,N_10948,N_10879);
or U11317 (N_11317,N_10556,N_10876);
nand U11318 (N_11318,N_10716,N_10856);
nand U11319 (N_11319,N_10543,N_10629);
nor U11320 (N_11320,N_10705,N_10703);
and U11321 (N_11321,N_10500,N_10606);
or U11322 (N_11322,N_10890,N_10961);
and U11323 (N_11323,N_10792,N_10927);
and U11324 (N_11324,N_10878,N_10542);
or U11325 (N_11325,N_10836,N_10669);
or U11326 (N_11326,N_10866,N_10544);
nor U11327 (N_11327,N_10641,N_10689);
or U11328 (N_11328,N_10848,N_10836);
or U11329 (N_11329,N_10639,N_10676);
nand U11330 (N_11330,N_10803,N_10715);
and U11331 (N_11331,N_10733,N_10845);
nand U11332 (N_11332,N_10621,N_10876);
and U11333 (N_11333,N_10614,N_10752);
or U11334 (N_11334,N_10631,N_10934);
nand U11335 (N_11335,N_10915,N_10938);
and U11336 (N_11336,N_10917,N_10742);
or U11337 (N_11337,N_10606,N_10761);
and U11338 (N_11338,N_10883,N_10755);
nor U11339 (N_11339,N_10565,N_10763);
and U11340 (N_11340,N_10760,N_10977);
and U11341 (N_11341,N_10589,N_10752);
nor U11342 (N_11342,N_10653,N_10981);
or U11343 (N_11343,N_10707,N_10799);
and U11344 (N_11344,N_10668,N_10788);
nor U11345 (N_11345,N_10584,N_10556);
or U11346 (N_11346,N_10979,N_10635);
nand U11347 (N_11347,N_10815,N_10975);
and U11348 (N_11348,N_10869,N_10654);
or U11349 (N_11349,N_10766,N_10954);
nor U11350 (N_11350,N_10682,N_10545);
and U11351 (N_11351,N_10963,N_10660);
or U11352 (N_11352,N_10992,N_10971);
nor U11353 (N_11353,N_10587,N_10932);
nor U11354 (N_11354,N_10910,N_10618);
or U11355 (N_11355,N_10648,N_10884);
or U11356 (N_11356,N_10834,N_10925);
or U11357 (N_11357,N_10527,N_10535);
nor U11358 (N_11358,N_10625,N_10801);
or U11359 (N_11359,N_10515,N_10608);
nand U11360 (N_11360,N_10971,N_10690);
nor U11361 (N_11361,N_10871,N_10898);
and U11362 (N_11362,N_10512,N_10655);
nand U11363 (N_11363,N_10887,N_10861);
or U11364 (N_11364,N_10645,N_10801);
xor U11365 (N_11365,N_10680,N_10964);
nand U11366 (N_11366,N_10749,N_10805);
xnor U11367 (N_11367,N_10574,N_10714);
or U11368 (N_11368,N_10798,N_10700);
nand U11369 (N_11369,N_10848,N_10701);
nor U11370 (N_11370,N_10537,N_10539);
and U11371 (N_11371,N_10990,N_10678);
xnor U11372 (N_11372,N_10585,N_10844);
nor U11373 (N_11373,N_10696,N_10577);
nor U11374 (N_11374,N_10758,N_10881);
nor U11375 (N_11375,N_10663,N_10872);
or U11376 (N_11376,N_10903,N_10627);
or U11377 (N_11377,N_10792,N_10595);
or U11378 (N_11378,N_10762,N_10522);
xor U11379 (N_11379,N_10706,N_10945);
nor U11380 (N_11380,N_10529,N_10848);
nor U11381 (N_11381,N_10897,N_10979);
nand U11382 (N_11382,N_10567,N_10556);
nor U11383 (N_11383,N_10644,N_10818);
nor U11384 (N_11384,N_10997,N_10964);
and U11385 (N_11385,N_10773,N_10745);
and U11386 (N_11386,N_10665,N_10916);
nor U11387 (N_11387,N_10938,N_10724);
nor U11388 (N_11388,N_10636,N_10731);
nor U11389 (N_11389,N_10850,N_10768);
and U11390 (N_11390,N_10845,N_10714);
xor U11391 (N_11391,N_10848,N_10941);
nor U11392 (N_11392,N_10984,N_10870);
or U11393 (N_11393,N_10570,N_10758);
nor U11394 (N_11394,N_10994,N_10589);
nor U11395 (N_11395,N_10708,N_10585);
and U11396 (N_11396,N_10760,N_10632);
nor U11397 (N_11397,N_10755,N_10565);
nor U11398 (N_11398,N_10761,N_10685);
nor U11399 (N_11399,N_10763,N_10690);
nand U11400 (N_11400,N_10887,N_10814);
and U11401 (N_11401,N_10765,N_10629);
and U11402 (N_11402,N_10799,N_10779);
xnor U11403 (N_11403,N_10795,N_10941);
and U11404 (N_11404,N_10759,N_10777);
nor U11405 (N_11405,N_10838,N_10861);
and U11406 (N_11406,N_10622,N_10611);
or U11407 (N_11407,N_10569,N_10942);
or U11408 (N_11408,N_10854,N_10763);
or U11409 (N_11409,N_10663,N_10755);
nand U11410 (N_11410,N_10561,N_10896);
and U11411 (N_11411,N_10915,N_10698);
nand U11412 (N_11412,N_10779,N_10985);
or U11413 (N_11413,N_10552,N_10931);
or U11414 (N_11414,N_10593,N_10604);
nor U11415 (N_11415,N_10616,N_10509);
or U11416 (N_11416,N_10881,N_10999);
or U11417 (N_11417,N_10820,N_10822);
and U11418 (N_11418,N_10947,N_10685);
xnor U11419 (N_11419,N_10911,N_10863);
or U11420 (N_11420,N_10828,N_10910);
and U11421 (N_11421,N_10765,N_10929);
nand U11422 (N_11422,N_10730,N_10673);
nand U11423 (N_11423,N_10685,N_10711);
or U11424 (N_11424,N_10741,N_10670);
nand U11425 (N_11425,N_10775,N_10799);
xor U11426 (N_11426,N_10865,N_10693);
and U11427 (N_11427,N_10864,N_10698);
nor U11428 (N_11428,N_10917,N_10932);
and U11429 (N_11429,N_10591,N_10917);
nand U11430 (N_11430,N_10524,N_10522);
nor U11431 (N_11431,N_10987,N_10635);
nor U11432 (N_11432,N_10922,N_10589);
nand U11433 (N_11433,N_10921,N_10977);
and U11434 (N_11434,N_10786,N_10829);
nand U11435 (N_11435,N_10830,N_10759);
or U11436 (N_11436,N_10699,N_10789);
nand U11437 (N_11437,N_10837,N_10883);
xnor U11438 (N_11438,N_10768,N_10642);
nor U11439 (N_11439,N_10947,N_10973);
nor U11440 (N_11440,N_10792,N_10929);
or U11441 (N_11441,N_10894,N_10941);
or U11442 (N_11442,N_10646,N_10612);
nand U11443 (N_11443,N_10958,N_10793);
nand U11444 (N_11444,N_10998,N_10795);
xnor U11445 (N_11445,N_10613,N_10954);
and U11446 (N_11446,N_10991,N_10905);
nand U11447 (N_11447,N_10516,N_10990);
or U11448 (N_11448,N_10973,N_10785);
nand U11449 (N_11449,N_10523,N_10640);
nand U11450 (N_11450,N_10896,N_10942);
and U11451 (N_11451,N_10854,N_10529);
and U11452 (N_11452,N_10836,N_10625);
and U11453 (N_11453,N_10890,N_10510);
or U11454 (N_11454,N_10884,N_10911);
or U11455 (N_11455,N_10885,N_10934);
xor U11456 (N_11456,N_10880,N_10907);
xnor U11457 (N_11457,N_10692,N_10781);
nand U11458 (N_11458,N_10796,N_10809);
or U11459 (N_11459,N_10998,N_10709);
nor U11460 (N_11460,N_10965,N_10969);
or U11461 (N_11461,N_10548,N_10950);
or U11462 (N_11462,N_10909,N_10664);
nor U11463 (N_11463,N_10740,N_10836);
nand U11464 (N_11464,N_10695,N_10958);
or U11465 (N_11465,N_10877,N_10782);
or U11466 (N_11466,N_10744,N_10867);
and U11467 (N_11467,N_10772,N_10964);
nor U11468 (N_11468,N_10687,N_10510);
nor U11469 (N_11469,N_10744,N_10608);
xor U11470 (N_11470,N_10616,N_10578);
nor U11471 (N_11471,N_10505,N_10562);
and U11472 (N_11472,N_10533,N_10874);
and U11473 (N_11473,N_10697,N_10518);
nand U11474 (N_11474,N_10594,N_10719);
xor U11475 (N_11475,N_10774,N_10896);
nor U11476 (N_11476,N_10634,N_10574);
and U11477 (N_11477,N_10795,N_10717);
nand U11478 (N_11478,N_10894,N_10583);
nand U11479 (N_11479,N_10747,N_10997);
nand U11480 (N_11480,N_10825,N_10831);
or U11481 (N_11481,N_10750,N_10554);
xnor U11482 (N_11482,N_10548,N_10814);
nand U11483 (N_11483,N_10975,N_10953);
and U11484 (N_11484,N_10582,N_10818);
nand U11485 (N_11485,N_10689,N_10805);
or U11486 (N_11486,N_10916,N_10759);
or U11487 (N_11487,N_10641,N_10502);
or U11488 (N_11488,N_10631,N_10597);
xor U11489 (N_11489,N_10903,N_10673);
and U11490 (N_11490,N_10775,N_10973);
xor U11491 (N_11491,N_10929,N_10984);
nand U11492 (N_11492,N_10692,N_10696);
nor U11493 (N_11493,N_10558,N_10581);
nor U11494 (N_11494,N_10517,N_10910);
nor U11495 (N_11495,N_10917,N_10579);
or U11496 (N_11496,N_10545,N_10953);
nor U11497 (N_11497,N_10604,N_10506);
nor U11498 (N_11498,N_10661,N_10558);
or U11499 (N_11499,N_10885,N_10919);
and U11500 (N_11500,N_11257,N_11017);
nor U11501 (N_11501,N_11157,N_11011);
nand U11502 (N_11502,N_11241,N_11062);
xor U11503 (N_11503,N_11283,N_11098);
xnor U11504 (N_11504,N_11326,N_11311);
and U11505 (N_11505,N_11380,N_11269);
or U11506 (N_11506,N_11091,N_11163);
nand U11507 (N_11507,N_11228,N_11023);
nor U11508 (N_11508,N_11175,N_11472);
nand U11509 (N_11509,N_11219,N_11295);
and U11510 (N_11510,N_11126,N_11347);
or U11511 (N_11511,N_11153,N_11189);
nor U11512 (N_11512,N_11349,N_11418);
nor U11513 (N_11513,N_11289,N_11460);
nand U11514 (N_11514,N_11248,N_11094);
or U11515 (N_11515,N_11089,N_11430);
nand U11516 (N_11516,N_11211,N_11376);
xor U11517 (N_11517,N_11379,N_11335);
and U11518 (N_11518,N_11333,N_11266);
nor U11519 (N_11519,N_11270,N_11281);
and U11520 (N_11520,N_11142,N_11398);
or U11521 (N_11521,N_11013,N_11217);
nand U11522 (N_11522,N_11093,N_11232);
nor U11523 (N_11523,N_11229,N_11396);
nand U11524 (N_11524,N_11144,N_11429);
or U11525 (N_11525,N_11192,N_11355);
nor U11526 (N_11526,N_11306,N_11156);
nand U11527 (N_11527,N_11360,N_11182);
or U11528 (N_11528,N_11403,N_11434);
and U11529 (N_11529,N_11246,N_11428);
nor U11530 (N_11530,N_11100,N_11127);
and U11531 (N_11531,N_11378,N_11179);
xor U11532 (N_11532,N_11481,N_11374);
nand U11533 (N_11533,N_11441,N_11484);
nor U11534 (N_11534,N_11329,N_11086);
xor U11535 (N_11535,N_11095,N_11286);
xnor U11536 (N_11536,N_11279,N_11332);
nand U11537 (N_11537,N_11168,N_11413);
or U11538 (N_11538,N_11421,N_11440);
nor U11539 (N_11539,N_11492,N_11452);
or U11540 (N_11540,N_11316,N_11302);
nand U11541 (N_11541,N_11363,N_11328);
xnor U11542 (N_11542,N_11214,N_11082);
and U11543 (N_11543,N_11358,N_11400);
xor U11544 (N_11544,N_11215,N_11446);
xnor U11545 (N_11545,N_11372,N_11467);
nand U11546 (N_11546,N_11384,N_11410);
nand U11547 (N_11547,N_11470,N_11046);
and U11548 (N_11548,N_11394,N_11395);
and U11549 (N_11549,N_11176,N_11435);
and U11550 (N_11550,N_11278,N_11498);
nor U11551 (N_11551,N_11310,N_11039);
nor U11552 (N_11552,N_11385,N_11244);
xnor U11553 (N_11553,N_11028,N_11317);
nor U11554 (N_11554,N_11019,N_11304);
or U11555 (N_11555,N_11321,N_11463);
and U11556 (N_11556,N_11407,N_11024);
nand U11557 (N_11557,N_11137,N_11292);
and U11558 (N_11558,N_11370,N_11053);
nand U11559 (N_11559,N_11212,N_11488);
nor U11560 (N_11560,N_11000,N_11366);
or U11561 (N_11561,N_11473,N_11030);
or U11562 (N_11562,N_11450,N_11088);
nand U11563 (N_11563,N_11108,N_11218);
and U11564 (N_11564,N_11060,N_11442);
nand U11565 (N_11565,N_11254,N_11064);
nand U11566 (N_11566,N_11164,N_11461);
or U11567 (N_11567,N_11287,N_11177);
nor U11568 (N_11568,N_11475,N_11107);
xor U11569 (N_11569,N_11027,N_11221);
xnor U11570 (N_11570,N_11008,N_11348);
nand U11571 (N_11571,N_11132,N_11495);
xor U11572 (N_11572,N_11154,N_11439);
xor U11573 (N_11573,N_11167,N_11146);
nand U11574 (N_11574,N_11051,N_11252);
or U11575 (N_11575,N_11392,N_11061);
nand U11576 (N_11576,N_11405,N_11387);
nand U11577 (N_11577,N_11462,N_11065);
and U11578 (N_11578,N_11105,N_11340);
and U11579 (N_11579,N_11052,N_11198);
nor U11580 (N_11580,N_11309,N_11298);
nand U11581 (N_11581,N_11256,N_11388);
and U11582 (N_11582,N_11101,N_11456);
nand U11583 (N_11583,N_11025,N_11466);
xnor U11584 (N_11584,N_11021,N_11250);
nor U11585 (N_11585,N_11477,N_11259);
xnor U11586 (N_11586,N_11102,N_11409);
and U11587 (N_11587,N_11206,N_11494);
or U11588 (N_11588,N_11300,N_11483);
xnor U11589 (N_11589,N_11097,N_11161);
xnor U11590 (N_11590,N_11263,N_11322);
or U11591 (N_11591,N_11239,N_11354);
and U11592 (N_11592,N_11031,N_11468);
and U11593 (N_11593,N_11282,N_11047);
and U11594 (N_11594,N_11114,N_11145);
and U11595 (N_11595,N_11227,N_11077);
nand U11596 (N_11596,N_11325,N_11247);
and U11597 (N_11597,N_11389,N_11341);
nor U11598 (N_11598,N_11303,N_11271);
nor U11599 (N_11599,N_11158,N_11345);
and U11600 (N_11600,N_11264,N_11399);
and U11601 (N_11601,N_11222,N_11201);
nand U11602 (N_11602,N_11152,N_11447);
nor U11603 (N_11603,N_11480,N_11180);
or U11604 (N_11604,N_11104,N_11045);
and U11605 (N_11605,N_11069,N_11103);
nand U11606 (N_11606,N_11131,N_11072);
and U11607 (N_11607,N_11408,N_11267);
nand U11608 (N_11608,N_11479,N_11453);
xnor U11609 (N_11609,N_11268,N_11207);
or U11610 (N_11610,N_11187,N_11369);
nand U11611 (N_11611,N_11174,N_11171);
or U11612 (N_11612,N_11169,N_11373);
nor U11613 (N_11613,N_11478,N_11210);
and U11614 (N_11614,N_11016,N_11487);
nor U11615 (N_11615,N_11141,N_11084);
or U11616 (N_11616,N_11070,N_11121);
and U11617 (N_11617,N_11136,N_11050);
or U11618 (N_11618,N_11299,N_11075);
nand U11619 (N_11619,N_11469,N_11411);
nor U11620 (N_11620,N_11401,N_11020);
nor U11621 (N_11621,N_11191,N_11296);
or U11622 (N_11622,N_11048,N_11438);
and U11623 (N_11623,N_11188,N_11415);
nand U11624 (N_11624,N_11004,N_11151);
nor U11625 (N_11625,N_11049,N_11033);
or U11626 (N_11626,N_11022,N_11116);
and U11627 (N_11627,N_11356,N_11386);
nand U11628 (N_11628,N_11111,N_11445);
nor U11629 (N_11629,N_11149,N_11068);
and U11630 (N_11630,N_11041,N_11476);
nand U11631 (N_11631,N_11249,N_11337);
or U11632 (N_11632,N_11138,N_11124);
and U11633 (N_11633,N_11087,N_11160);
nor U11634 (N_11634,N_11260,N_11391);
or U11635 (N_11635,N_11342,N_11390);
or U11636 (N_11636,N_11197,N_11006);
xnor U11637 (N_11637,N_11485,N_11242);
or U11638 (N_11638,N_11074,N_11275);
or U11639 (N_11639,N_11083,N_11314);
or U11640 (N_11640,N_11276,N_11417);
or U11641 (N_11641,N_11115,N_11085);
nand U11642 (N_11642,N_11120,N_11036);
xnor U11643 (N_11643,N_11420,N_11106);
and U11644 (N_11644,N_11220,N_11285);
nor U11645 (N_11645,N_11393,N_11251);
and U11646 (N_11646,N_11284,N_11007);
nand U11647 (N_11647,N_11262,N_11165);
nand U11648 (N_11648,N_11135,N_11181);
nor U11649 (N_11649,N_11080,N_11371);
nor U11650 (N_11650,N_11291,N_11324);
and U11651 (N_11651,N_11204,N_11213);
nand U11652 (N_11652,N_11336,N_11117);
nor U11653 (N_11653,N_11147,N_11067);
and U11654 (N_11654,N_11327,N_11338);
nor U11655 (N_11655,N_11003,N_11243);
nor U11656 (N_11656,N_11431,N_11464);
nand U11657 (N_11657,N_11190,N_11245);
nor U11658 (N_11658,N_11029,N_11140);
nand U11659 (N_11659,N_11044,N_11422);
nand U11660 (N_11660,N_11235,N_11056);
nand U11661 (N_11661,N_11294,N_11265);
nand U11662 (N_11662,N_11018,N_11493);
or U11663 (N_11663,N_11183,N_11313);
nor U11664 (N_11664,N_11362,N_11134);
or U11665 (N_11665,N_11320,N_11465);
nand U11666 (N_11666,N_11482,N_11357);
nand U11667 (N_11667,N_11226,N_11397);
and U11668 (N_11668,N_11312,N_11035);
xnor U11669 (N_11669,N_11377,N_11307);
or U11670 (N_11670,N_11150,N_11416);
or U11671 (N_11671,N_11381,N_11076);
or U11672 (N_11672,N_11375,N_11186);
nor U11673 (N_11673,N_11012,N_11034);
nand U11674 (N_11674,N_11489,N_11274);
and U11675 (N_11675,N_11425,N_11119);
nand U11676 (N_11676,N_11193,N_11330);
or U11677 (N_11677,N_11331,N_11293);
or U11678 (N_11678,N_11009,N_11352);
xnor U11679 (N_11679,N_11055,N_11208);
xor U11680 (N_11680,N_11129,N_11199);
nand U11681 (N_11681,N_11449,N_11353);
xnor U11682 (N_11682,N_11081,N_11491);
nand U11683 (N_11683,N_11471,N_11042);
nand U11684 (N_11684,N_11433,N_11280);
and U11685 (N_11685,N_11015,N_11110);
nor U11686 (N_11686,N_11092,N_11402);
and U11687 (N_11687,N_11184,N_11404);
nand U11688 (N_11688,N_11133,N_11113);
nand U11689 (N_11689,N_11159,N_11225);
nor U11690 (N_11690,N_11459,N_11490);
or U11691 (N_11691,N_11486,N_11202);
nor U11692 (N_11692,N_11436,N_11090);
nand U11693 (N_11693,N_11238,N_11364);
and U11694 (N_11694,N_11424,N_11178);
xor U11695 (N_11695,N_11172,N_11005);
and U11696 (N_11696,N_11231,N_11305);
nor U11697 (N_11697,N_11122,N_11237);
nor U11698 (N_11698,N_11130,N_11038);
nor U11699 (N_11699,N_11255,N_11315);
or U11700 (N_11700,N_11339,N_11162);
nand U11701 (N_11701,N_11230,N_11444);
nand U11702 (N_11702,N_11196,N_11002);
nand U11703 (N_11703,N_11155,N_11318);
or U11704 (N_11704,N_11059,N_11063);
xnor U11705 (N_11705,N_11451,N_11043);
nand U11706 (N_11706,N_11496,N_11234);
nand U11707 (N_11707,N_11079,N_11367);
and U11708 (N_11708,N_11143,N_11078);
xor U11709 (N_11709,N_11185,N_11412);
or U11710 (N_11710,N_11344,N_11323);
nor U11711 (N_11711,N_11437,N_11148);
nor U11712 (N_11712,N_11448,N_11361);
nand U11713 (N_11713,N_11258,N_11290);
and U11714 (N_11714,N_11073,N_11423);
or U11715 (N_11715,N_11195,N_11432);
or U11716 (N_11716,N_11301,N_11261);
nor U11717 (N_11717,N_11368,N_11288);
nor U11718 (N_11718,N_11426,N_11026);
and U11719 (N_11719,N_11359,N_11205);
nor U11720 (N_11720,N_11224,N_11058);
xnor U11721 (N_11721,N_11057,N_11071);
and U11722 (N_11722,N_11272,N_11365);
or U11723 (N_11723,N_11096,N_11099);
nor U11724 (N_11724,N_11499,N_11443);
and U11725 (N_11725,N_11014,N_11223);
or U11726 (N_11726,N_11170,N_11406);
and U11727 (N_11727,N_11040,N_11382);
nor U11728 (N_11728,N_11351,N_11455);
and U11729 (N_11729,N_11383,N_11203);
or U11730 (N_11730,N_11010,N_11236);
and U11731 (N_11731,N_11457,N_11112);
nand U11732 (N_11732,N_11497,N_11037);
nand U11733 (N_11733,N_11458,N_11216);
nand U11734 (N_11734,N_11123,N_11194);
nor U11735 (N_11735,N_11277,N_11209);
and U11736 (N_11736,N_11139,N_11297);
nor U11737 (N_11737,N_11253,N_11118);
and U11738 (N_11738,N_11414,N_11200);
nor U11739 (N_11739,N_11454,N_11273);
nand U11740 (N_11740,N_11427,N_11343);
nor U11741 (N_11741,N_11128,N_11419);
nor U11742 (N_11742,N_11054,N_11125);
nor U11743 (N_11743,N_11334,N_11240);
or U11744 (N_11744,N_11233,N_11109);
nand U11745 (N_11745,N_11001,N_11346);
nand U11746 (N_11746,N_11308,N_11166);
nor U11747 (N_11747,N_11066,N_11032);
nor U11748 (N_11748,N_11474,N_11173);
nand U11749 (N_11749,N_11319,N_11350);
and U11750 (N_11750,N_11422,N_11006);
and U11751 (N_11751,N_11231,N_11213);
xnor U11752 (N_11752,N_11358,N_11491);
nand U11753 (N_11753,N_11431,N_11286);
and U11754 (N_11754,N_11410,N_11304);
nand U11755 (N_11755,N_11298,N_11404);
and U11756 (N_11756,N_11457,N_11127);
xnor U11757 (N_11757,N_11460,N_11488);
nor U11758 (N_11758,N_11040,N_11432);
or U11759 (N_11759,N_11009,N_11058);
nor U11760 (N_11760,N_11343,N_11053);
xnor U11761 (N_11761,N_11214,N_11396);
nand U11762 (N_11762,N_11005,N_11158);
nor U11763 (N_11763,N_11150,N_11252);
nor U11764 (N_11764,N_11333,N_11069);
xor U11765 (N_11765,N_11127,N_11468);
nand U11766 (N_11766,N_11107,N_11428);
nand U11767 (N_11767,N_11043,N_11321);
nand U11768 (N_11768,N_11074,N_11111);
xor U11769 (N_11769,N_11135,N_11325);
nand U11770 (N_11770,N_11149,N_11407);
nand U11771 (N_11771,N_11271,N_11237);
nand U11772 (N_11772,N_11365,N_11057);
or U11773 (N_11773,N_11217,N_11181);
nand U11774 (N_11774,N_11110,N_11493);
nor U11775 (N_11775,N_11402,N_11058);
or U11776 (N_11776,N_11259,N_11102);
and U11777 (N_11777,N_11230,N_11308);
and U11778 (N_11778,N_11480,N_11377);
or U11779 (N_11779,N_11203,N_11461);
and U11780 (N_11780,N_11461,N_11113);
nand U11781 (N_11781,N_11253,N_11404);
and U11782 (N_11782,N_11280,N_11408);
or U11783 (N_11783,N_11349,N_11105);
xor U11784 (N_11784,N_11441,N_11101);
and U11785 (N_11785,N_11276,N_11065);
xor U11786 (N_11786,N_11322,N_11199);
and U11787 (N_11787,N_11048,N_11352);
nor U11788 (N_11788,N_11473,N_11334);
nor U11789 (N_11789,N_11166,N_11249);
xor U11790 (N_11790,N_11145,N_11472);
and U11791 (N_11791,N_11309,N_11466);
nand U11792 (N_11792,N_11489,N_11010);
nand U11793 (N_11793,N_11029,N_11422);
xor U11794 (N_11794,N_11331,N_11213);
nand U11795 (N_11795,N_11211,N_11390);
and U11796 (N_11796,N_11448,N_11280);
xor U11797 (N_11797,N_11479,N_11194);
nand U11798 (N_11798,N_11029,N_11074);
and U11799 (N_11799,N_11416,N_11007);
and U11800 (N_11800,N_11250,N_11042);
and U11801 (N_11801,N_11397,N_11477);
xnor U11802 (N_11802,N_11422,N_11291);
or U11803 (N_11803,N_11327,N_11215);
or U11804 (N_11804,N_11116,N_11390);
xor U11805 (N_11805,N_11125,N_11024);
or U11806 (N_11806,N_11164,N_11353);
nand U11807 (N_11807,N_11175,N_11234);
and U11808 (N_11808,N_11276,N_11057);
and U11809 (N_11809,N_11199,N_11417);
xnor U11810 (N_11810,N_11316,N_11220);
and U11811 (N_11811,N_11256,N_11442);
or U11812 (N_11812,N_11079,N_11160);
nand U11813 (N_11813,N_11426,N_11139);
xnor U11814 (N_11814,N_11446,N_11073);
xor U11815 (N_11815,N_11257,N_11182);
nor U11816 (N_11816,N_11068,N_11194);
nor U11817 (N_11817,N_11309,N_11018);
or U11818 (N_11818,N_11384,N_11077);
or U11819 (N_11819,N_11167,N_11224);
and U11820 (N_11820,N_11164,N_11240);
or U11821 (N_11821,N_11341,N_11361);
and U11822 (N_11822,N_11351,N_11168);
nor U11823 (N_11823,N_11106,N_11213);
xor U11824 (N_11824,N_11316,N_11332);
nand U11825 (N_11825,N_11349,N_11117);
or U11826 (N_11826,N_11068,N_11184);
or U11827 (N_11827,N_11490,N_11284);
nor U11828 (N_11828,N_11249,N_11347);
nand U11829 (N_11829,N_11124,N_11217);
or U11830 (N_11830,N_11251,N_11203);
nand U11831 (N_11831,N_11199,N_11165);
nand U11832 (N_11832,N_11313,N_11127);
and U11833 (N_11833,N_11393,N_11461);
xor U11834 (N_11834,N_11308,N_11364);
or U11835 (N_11835,N_11129,N_11489);
or U11836 (N_11836,N_11096,N_11491);
and U11837 (N_11837,N_11040,N_11221);
and U11838 (N_11838,N_11408,N_11153);
and U11839 (N_11839,N_11325,N_11102);
xnor U11840 (N_11840,N_11133,N_11163);
nand U11841 (N_11841,N_11360,N_11133);
nor U11842 (N_11842,N_11363,N_11452);
nor U11843 (N_11843,N_11042,N_11276);
nor U11844 (N_11844,N_11258,N_11448);
nand U11845 (N_11845,N_11247,N_11355);
nor U11846 (N_11846,N_11155,N_11372);
nand U11847 (N_11847,N_11095,N_11368);
nor U11848 (N_11848,N_11395,N_11325);
nor U11849 (N_11849,N_11474,N_11196);
or U11850 (N_11850,N_11457,N_11179);
nor U11851 (N_11851,N_11455,N_11150);
nor U11852 (N_11852,N_11415,N_11372);
nand U11853 (N_11853,N_11244,N_11149);
nor U11854 (N_11854,N_11427,N_11113);
nand U11855 (N_11855,N_11178,N_11251);
nand U11856 (N_11856,N_11465,N_11126);
or U11857 (N_11857,N_11082,N_11023);
or U11858 (N_11858,N_11264,N_11200);
and U11859 (N_11859,N_11367,N_11108);
nand U11860 (N_11860,N_11156,N_11403);
nand U11861 (N_11861,N_11402,N_11025);
or U11862 (N_11862,N_11049,N_11335);
nand U11863 (N_11863,N_11393,N_11422);
nor U11864 (N_11864,N_11429,N_11433);
and U11865 (N_11865,N_11277,N_11063);
xor U11866 (N_11866,N_11248,N_11466);
nand U11867 (N_11867,N_11302,N_11319);
nor U11868 (N_11868,N_11255,N_11180);
or U11869 (N_11869,N_11217,N_11467);
or U11870 (N_11870,N_11327,N_11321);
nand U11871 (N_11871,N_11393,N_11491);
nand U11872 (N_11872,N_11393,N_11011);
and U11873 (N_11873,N_11356,N_11166);
nor U11874 (N_11874,N_11022,N_11482);
nor U11875 (N_11875,N_11320,N_11093);
or U11876 (N_11876,N_11259,N_11071);
nor U11877 (N_11877,N_11178,N_11070);
and U11878 (N_11878,N_11013,N_11445);
nand U11879 (N_11879,N_11293,N_11114);
nand U11880 (N_11880,N_11122,N_11496);
nand U11881 (N_11881,N_11405,N_11334);
and U11882 (N_11882,N_11292,N_11471);
and U11883 (N_11883,N_11344,N_11177);
nand U11884 (N_11884,N_11427,N_11204);
nand U11885 (N_11885,N_11385,N_11460);
xnor U11886 (N_11886,N_11245,N_11376);
nor U11887 (N_11887,N_11280,N_11051);
or U11888 (N_11888,N_11312,N_11191);
and U11889 (N_11889,N_11353,N_11111);
nand U11890 (N_11890,N_11197,N_11432);
nand U11891 (N_11891,N_11380,N_11101);
nor U11892 (N_11892,N_11201,N_11244);
nor U11893 (N_11893,N_11068,N_11236);
or U11894 (N_11894,N_11205,N_11422);
or U11895 (N_11895,N_11124,N_11409);
nor U11896 (N_11896,N_11182,N_11407);
xor U11897 (N_11897,N_11268,N_11180);
and U11898 (N_11898,N_11040,N_11455);
nand U11899 (N_11899,N_11400,N_11013);
or U11900 (N_11900,N_11258,N_11438);
nor U11901 (N_11901,N_11176,N_11277);
and U11902 (N_11902,N_11376,N_11389);
and U11903 (N_11903,N_11348,N_11074);
nor U11904 (N_11904,N_11121,N_11158);
nand U11905 (N_11905,N_11490,N_11155);
and U11906 (N_11906,N_11218,N_11185);
xnor U11907 (N_11907,N_11239,N_11183);
and U11908 (N_11908,N_11006,N_11270);
nor U11909 (N_11909,N_11410,N_11358);
nand U11910 (N_11910,N_11160,N_11424);
or U11911 (N_11911,N_11025,N_11061);
and U11912 (N_11912,N_11377,N_11043);
or U11913 (N_11913,N_11326,N_11270);
and U11914 (N_11914,N_11311,N_11217);
and U11915 (N_11915,N_11186,N_11345);
xnor U11916 (N_11916,N_11421,N_11209);
nand U11917 (N_11917,N_11174,N_11463);
nor U11918 (N_11918,N_11007,N_11377);
and U11919 (N_11919,N_11398,N_11324);
or U11920 (N_11920,N_11169,N_11447);
and U11921 (N_11921,N_11242,N_11397);
and U11922 (N_11922,N_11341,N_11306);
xnor U11923 (N_11923,N_11377,N_11097);
nor U11924 (N_11924,N_11094,N_11007);
nand U11925 (N_11925,N_11044,N_11478);
or U11926 (N_11926,N_11469,N_11495);
and U11927 (N_11927,N_11063,N_11401);
nor U11928 (N_11928,N_11323,N_11310);
nand U11929 (N_11929,N_11316,N_11154);
and U11930 (N_11930,N_11481,N_11210);
or U11931 (N_11931,N_11474,N_11413);
nor U11932 (N_11932,N_11023,N_11078);
nor U11933 (N_11933,N_11245,N_11429);
xor U11934 (N_11934,N_11103,N_11341);
and U11935 (N_11935,N_11373,N_11027);
nor U11936 (N_11936,N_11357,N_11340);
nor U11937 (N_11937,N_11406,N_11447);
and U11938 (N_11938,N_11254,N_11329);
nor U11939 (N_11939,N_11387,N_11204);
or U11940 (N_11940,N_11048,N_11375);
or U11941 (N_11941,N_11028,N_11003);
xnor U11942 (N_11942,N_11347,N_11041);
or U11943 (N_11943,N_11412,N_11102);
nor U11944 (N_11944,N_11239,N_11335);
and U11945 (N_11945,N_11050,N_11392);
or U11946 (N_11946,N_11195,N_11460);
nor U11947 (N_11947,N_11477,N_11198);
and U11948 (N_11948,N_11019,N_11050);
nand U11949 (N_11949,N_11407,N_11164);
nor U11950 (N_11950,N_11251,N_11238);
and U11951 (N_11951,N_11317,N_11414);
nand U11952 (N_11952,N_11224,N_11466);
and U11953 (N_11953,N_11186,N_11360);
nand U11954 (N_11954,N_11092,N_11085);
xor U11955 (N_11955,N_11049,N_11090);
or U11956 (N_11956,N_11429,N_11462);
nor U11957 (N_11957,N_11117,N_11168);
nand U11958 (N_11958,N_11255,N_11338);
nor U11959 (N_11959,N_11182,N_11409);
or U11960 (N_11960,N_11199,N_11180);
nor U11961 (N_11961,N_11208,N_11426);
nand U11962 (N_11962,N_11059,N_11173);
and U11963 (N_11963,N_11430,N_11419);
or U11964 (N_11964,N_11251,N_11034);
or U11965 (N_11965,N_11498,N_11300);
xnor U11966 (N_11966,N_11048,N_11208);
nand U11967 (N_11967,N_11251,N_11320);
nand U11968 (N_11968,N_11389,N_11451);
xnor U11969 (N_11969,N_11160,N_11081);
nand U11970 (N_11970,N_11369,N_11071);
and U11971 (N_11971,N_11148,N_11103);
and U11972 (N_11972,N_11048,N_11004);
nand U11973 (N_11973,N_11111,N_11065);
or U11974 (N_11974,N_11118,N_11355);
and U11975 (N_11975,N_11046,N_11230);
nand U11976 (N_11976,N_11299,N_11431);
or U11977 (N_11977,N_11252,N_11296);
and U11978 (N_11978,N_11179,N_11344);
nand U11979 (N_11979,N_11298,N_11464);
and U11980 (N_11980,N_11263,N_11318);
and U11981 (N_11981,N_11234,N_11454);
nor U11982 (N_11982,N_11417,N_11311);
or U11983 (N_11983,N_11223,N_11359);
and U11984 (N_11984,N_11289,N_11462);
nor U11985 (N_11985,N_11157,N_11267);
nor U11986 (N_11986,N_11285,N_11483);
nand U11987 (N_11987,N_11451,N_11075);
nor U11988 (N_11988,N_11056,N_11188);
nand U11989 (N_11989,N_11270,N_11049);
or U11990 (N_11990,N_11353,N_11333);
and U11991 (N_11991,N_11002,N_11448);
nand U11992 (N_11992,N_11213,N_11345);
nand U11993 (N_11993,N_11171,N_11284);
and U11994 (N_11994,N_11093,N_11479);
and U11995 (N_11995,N_11266,N_11304);
and U11996 (N_11996,N_11282,N_11127);
or U11997 (N_11997,N_11279,N_11138);
nand U11998 (N_11998,N_11070,N_11265);
and U11999 (N_11999,N_11225,N_11434);
nor U12000 (N_12000,N_11712,N_11940);
nand U12001 (N_12001,N_11837,N_11830);
and U12002 (N_12002,N_11985,N_11887);
or U12003 (N_12003,N_11688,N_11708);
or U12004 (N_12004,N_11720,N_11973);
nand U12005 (N_12005,N_11654,N_11799);
nand U12006 (N_12006,N_11892,N_11538);
nand U12007 (N_12007,N_11714,N_11891);
and U12008 (N_12008,N_11789,N_11595);
or U12009 (N_12009,N_11513,N_11730);
or U12010 (N_12010,N_11767,N_11612);
and U12011 (N_12011,N_11813,N_11990);
or U12012 (N_12012,N_11858,N_11815);
nand U12013 (N_12013,N_11678,N_11782);
or U12014 (N_12014,N_11687,N_11844);
nand U12015 (N_12015,N_11849,N_11507);
or U12016 (N_12016,N_11845,N_11547);
nor U12017 (N_12017,N_11588,N_11929);
and U12018 (N_12018,N_11943,N_11855);
xor U12019 (N_12019,N_11899,N_11935);
or U12020 (N_12020,N_11853,N_11957);
nand U12021 (N_12021,N_11607,N_11975);
and U12022 (N_12022,N_11719,N_11821);
nand U12023 (N_12023,N_11555,N_11920);
xnor U12024 (N_12024,N_11976,N_11746);
and U12025 (N_12025,N_11805,N_11683);
nor U12026 (N_12026,N_11640,N_11979);
nor U12027 (N_12027,N_11885,N_11734);
nor U12028 (N_12028,N_11624,N_11890);
and U12029 (N_12029,N_11922,N_11982);
xnor U12030 (N_12030,N_11770,N_11515);
or U12031 (N_12031,N_11763,N_11584);
nand U12032 (N_12032,N_11748,N_11997);
or U12033 (N_12033,N_11665,N_11736);
and U12034 (N_12034,N_11505,N_11888);
nand U12035 (N_12035,N_11836,N_11702);
nor U12036 (N_12036,N_11857,N_11724);
nor U12037 (N_12037,N_11852,N_11539);
nor U12038 (N_12038,N_11949,N_11820);
xnor U12039 (N_12039,N_11895,N_11698);
and U12040 (N_12040,N_11671,N_11739);
nand U12041 (N_12041,N_11560,N_11741);
or U12042 (N_12042,N_11790,N_11953);
nor U12043 (N_12043,N_11727,N_11721);
and U12044 (N_12044,N_11601,N_11520);
nand U12045 (N_12045,N_11656,N_11930);
and U12046 (N_12046,N_11910,N_11946);
xnor U12047 (N_12047,N_11843,N_11627);
nand U12048 (N_12048,N_11901,N_11707);
or U12049 (N_12049,N_11585,N_11864);
or U12050 (N_12050,N_11598,N_11575);
nor U12051 (N_12051,N_11643,N_11919);
and U12052 (N_12052,N_11573,N_11699);
nand U12053 (N_12053,N_11916,N_11529);
or U12054 (N_12054,N_11868,N_11653);
nand U12055 (N_12055,N_11795,N_11851);
and U12056 (N_12056,N_11649,N_11765);
xnor U12057 (N_12057,N_11835,N_11609);
and U12058 (N_12058,N_11747,N_11711);
or U12059 (N_12059,N_11883,N_11915);
nand U12060 (N_12060,N_11806,N_11904);
xor U12061 (N_12061,N_11502,N_11618);
or U12062 (N_12062,N_11545,N_11784);
and U12063 (N_12063,N_11550,N_11684);
or U12064 (N_12064,N_11623,N_11797);
nand U12065 (N_12065,N_11523,N_11833);
and U12066 (N_12066,N_11589,N_11878);
nor U12067 (N_12067,N_11735,N_11576);
nand U12068 (N_12068,N_11673,N_11750);
nor U12069 (N_12069,N_11662,N_11625);
or U12070 (N_12070,N_11675,N_11691);
xnor U12071 (N_12071,N_11634,N_11956);
and U12072 (N_12072,N_11986,N_11993);
and U12073 (N_12073,N_11597,N_11717);
and U12074 (N_12074,N_11822,N_11798);
xnor U12075 (N_12075,N_11875,N_11945);
nor U12076 (N_12076,N_11840,N_11743);
xnor U12077 (N_12077,N_11593,N_11906);
or U12078 (N_12078,N_11559,N_11530);
nor U12079 (N_12079,N_11972,N_11674);
xor U12080 (N_12080,N_11621,N_11728);
nand U12081 (N_12081,N_11570,N_11599);
or U12082 (N_12082,N_11731,N_11670);
nor U12083 (N_12083,N_11508,N_11827);
nor U12084 (N_12084,N_11579,N_11948);
xnor U12085 (N_12085,N_11557,N_11944);
nand U12086 (N_12086,N_11517,N_11749);
nor U12087 (N_12087,N_11771,N_11603);
nor U12088 (N_12088,N_11859,N_11867);
nor U12089 (N_12089,N_11680,N_11518);
or U12090 (N_12090,N_11677,N_11974);
nand U12091 (N_12091,N_11549,N_11633);
or U12092 (N_12092,N_11686,N_11970);
and U12093 (N_12093,N_11808,N_11546);
xnor U12094 (N_12094,N_11817,N_11527);
and U12095 (N_12095,N_11889,N_11774);
nor U12096 (N_12096,N_11969,N_11810);
or U12097 (N_12097,N_11528,N_11966);
nand U12098 (N_12098,N_11936,N_11705);
and U12099 (N_12099,N_11984,N_11861);
and U12100 (N_12100,N_11777,N_11657);
nor U12101 (N_12101,N_11632,N_11586);
nor U12102 (N_12102,N_11617,N_11718);
and U12103 (N_12103,N_11902,N_11554);
and U12104 (N_12104,N_11882,N_11566);
xor U12105 (N_12105,N_11873,N_11532);
and U12106 (N_12106,N_11622,N_11918);
and U12107 (N_12107,N_11602,N_11773);
or U12108 (N_12108,N_11667,N_11682);
nor U12109 (N_12109,N_11534,N_11610);
nand U12110 (N_12110,N_11905,N_11998);
nand U12111 (N_12111,N_11783,N_11761);
and U12112 (N_12112,N_11960,N_11553);
nand U12113 (N_12113,N_11825,N_11577);
nor U12114 (N_12114,N_11694,N_11879);
nor U12115 (N_12115,N_11504,N_11860);
or U12116 (N_12116,N_11663,N_11543);
or U12117 (N_12117,N_11689,N_11819);
nand U12118 (N_12118,N_11596,N_11756);
nand U12119 (N_12119,N_11781,N_11600);
or U12120 (N_12120,N_11626,N_11792);
and U12121 (N_12121,N_11934,N_11939);
or U12122 (N_12122,N_11582,N_11655);
and U12123 (N_12123,N_11863,N_11569);
xor U12124 (N_12124,N_11893,N_11967);
or U12125 (N_12125,N_11572,N_11636);
nor U12126 (N_12126,N_11614,N_11876);
nand U12127 (N_12127,N_11881,N_11669);
nand U12128 (N_12128,N_11661,N_11704);
and U12129 (N_12129,N_11932,N_11506);
nor U12130 (N_12130,N_11531,N_11992);
xor U12131 (N_12131,N_11884,N_11759);
nand U12132 (N_12132,N_11787,N_11591);
nor U12133 (N_12133,N_11574,N_11824);
nor U12134 (N_12134,N_11762,N_11722);
or U12135 (N_12135,N_11668,N_11524);
and U12136 (N_12136,N_11514,N_11754);
and U12137 (N_12137,N_11696,N_11710);
or U12138 (N_12138,N_11897,N_11715);
nand U12139 (N_12139,N_11926,N_11594);
nand U12140 (N_12140,N_11793,N_11628);
nand U12141 (N_12141,N_11695,N_11796);
or U12142 (N_12142,N_11854,N_11651);
and U12143 (N_12143,N_11681,N_11877);
and U12144 (N_12144,N_11605,N_11676);
nor U12145 (N_12145,N_11914,N_11500);
nor U12146 (N_12146,N_11785,N_11788);
or U12147 (N_12147,N_11923,N_11801);
nor U12148 (N_12148,N_11959,N_11613);
xor U12149 (N_12149,N_11697,N_11764);
and U12150 (N_12150,N_11648,N_11729);
or U12151 (N_12151,N_11690,N_11869);
and U12152 (N_12152,N_11962,N_11733);
or U12153 (N_12153,N_11866,N_11757);
nand U12154 (N_12154,N_11666,N_11862);
nor U12155 (N_12155,N_11816,N_11841);
nand U12156 (N_12156,N_11658,N_11811);
xnor U12157 (N_12157,N_11896,N_11870);
and U12158 (N_12158,N_11629,N_11894);
and U12159 (N_12159,N_11900,N_11995);
nor U12160 (N_12160,N_11725,N_11871);
or U12161 (N_12161,N_11548,N_11556);
nand U12162 (N_12162,N_11700,N_11846);
and U12163 (N_12163,N_11941,N_11713);
and U12164 (N_12164,N_11692,N_11652);
or U12165 (N_12165,N_11786,N_11631);
and U12166 (N_12166,N_11512,N_11706);
nand U12167 (N_12167,N_11616,N_11672);
xor U12168 (N_12168,N_11950,N_11842);
or U12169 (N_12169,N_11907,N_11988);
and U12170 (N_12170,N_11753,N_11552);
nor U12171 (N_12171,N_11647,N_11563);
nor U12172 (N_12172,N_11758,N_11971);
nor U12173 (N_12173,N_11865,N_11642);
nor U12174 (N_12174,N_11650,N_11703);
nand U12175 (N_12175,N_11679,N_11768);
nor U12176 (N_12176,N_11778,N_11590);
or U12177 (N_12177,N_11780,N_11752);
nand U12178 (N_12178,N_11645,N_11947);
nor U12179 (N_12179,N_11525,N_11839);
or U12180 (N_12180,N_11537,N_11615);
and U12181 (N_12181,N_11581,N_11583);
nor U12182 (N_12182,N_11834,N_11903);
and U12183 (N_12183,N_11978,N_11503);
and U12184 (N_12184,N_11807,N_11968);
nor U12185 (N_12185,N_11536,N_11542);
and U12186 (N_12186,N_11567,N_11814);
and U12187 (N_12187,N_11937,N_11912);
nor U12188 (N_12188,N_11568,N_11608);
nand U12189 (N_12189,N_11541,N_11933);
xor U12190 (N_12190,N_11664,N_11991);
xor U12191 (N_12191,N_11938,N_11954);
and U12192 (N_12192,N_11755,N_11927);
nand U12193 (N_12193,N_11983,N_11921);
nand U12194 (N_12194,N_11744,N_11803);
nor U12195 (N_12195,N_11989,N_11535);
or U12196 (N_12196,N_11516,N_11802);
and U12197 (N_12197,N_11620,N_11809);
or U12198 (N_12198,N_11856,N_11587);
nor U12199 (N_12199,N_11886,N_11760);
nand U12200 (N_12200,N_11604,N_11977);
nor U12201 (N_12201,N_11776,N_11779);
xor U12202 (N_12202,N_11963,N_11660);
or U12203 (N_12203,N_11838,N_11994);
nor U12204 (N_12204,N_11925,N_11726);
and U12205 (N_12205,N_11928,N_11644);
or U12206 (N_12206,N_11880,N_11592);
or U12207 (N_12207,N_11908,N_11911);
nor U12208 (N_12208,N_11533,N_11742);
or U12209 (N_12209,N_11558,N_11641);
nand U12210 (N_12210,N_11521,N_11874);
nor U12211 (N_12211,N_11955,N_11723);
nand U12212 (N_12212,N_11522,N_11738);
or U12213 (N_12213,N_11740,N_11701);
nor U12214 (N_12214,N_11804,N_11829);
nor U12215 (N_12215,N_11800,N_11812);
nand U12216 (N_12216,N_11639,N_11909);
or U12217 (N_12217,N_11958,N_11511);
and U12218 (N_12218,N_11659,N_11818);
nor U12219 (N_12219,N_11980,N_11519);
nand U12220 (N_12220,N_11737,N_11850);
nor U12221 (N_12221,N_11999,N_11996);
or U12222 (N_12222,N_11917,N_11638);
and U12223 (N_12223,N_11606,N_11913);
and U12224 (N_12224,N_11580,N_11685);
nand U12225 (N_12225,N_11828,N_11872);
or U12226 (N_12226,N_11630,N_11564);
xor U12227 (N_12227,N_11823,N_11526);
nand U12228 (N_12228,N_11961,N_11551);
xnor U12229 (N_12229,N_11732,N_11766);
nand U12230 (N_12230,N_11716,N_11637);
or U12231 (N_12231,N_11561,N_11745);
and U12232 (N_12232,N_11693,N_11562);
nor U12233 (N_12233,N_11951,N_11964);
or U12234 (N_12234,N_11611,N_11571);
nand U12235 (N_12235,N_11565,N_11952);
nor U12236 (N_12236,N_11898,N_11509);
nand U12237 (N_12237,N_11831,N_11510);
and U12238 (N_12238,N_11981,N_11751);
nand U12239 (N_12239,N_11794,N_11646);
nor U12240 (N_12240,N_11832,N_11544);
nor U12241 (N_12241,N_11619,N_11791);
or U12242 (N_12242,N_11847,N_11931);
nor U12243 (N_12243,N_11965,N_11775);
nand U12244 (N_12244,N_11635,N_11924);
xnor U12245 (N_12245,N_11769,N_11826);
nor U12246 (N_12246,N_11987,N_11540);
nor U12247 (N_12247,N_11578,N_11772);
or U12248 (N_12248,N_11709,N_11501);
and U12249 (N_12249,N_11848,N_11942);
nand U12250 (N_12250,N_11629,N_11708);
nor U12251 (N_12251,N_11616,N_11615);
and U12252 (N_12252,N_11771,N_11913);
nor U12253 (N_12253,N_11853,N_11730);
or U12254 (N_12254,N_11929,N_11512);
or U12255 (N_12255,N_11580,N_11823);
or U12256 (N_12256,N_11530,N_11660);
or U12257 (N_12257,N_11607,N_11734);
nor U12258 (N_12258,N_11704,N_11509);
or U12259 (N_12259,N_11569,N_11543);
nand U12260 (N_12260,N_11531,N_11956);
and U12261 (N_12261,N_11761,N_11605);
or U12262 (N_12262,N_11886,N_11677);
xor U12263 (N_12263,N_11824,N_11589);
and U12264 (N_12264,N_11680,N_11576);
and U12265 (N_12265,N_11654,N_11717);
and U12266 (N_12266,N_11623,N_11851);
and U12267 (N_12267,N_11611,N_11902);
nand U12268 (N_12268,N_11708,N_11604);
nand U12269 (N_12269,N_11837,N_11639);
or U12270 (N_12270,N_11580,N_11534);
xnor U12271 (N_12271,N_11658,N_11629);
and U12272 (N_12272,N_11810,N_11908);
nor U12273 (N_12273,N_11619,N_11673);
xor U12274 (N_12274,N_11687,N_11777);
nor U12275 (N_12275,N_11743,N_11807);
and U12276 (N_12276,N_11579,N_11786);
and U12277 (N_12277,N_11882,N_11637);
or U12278 (N_12278,N_11718,N_11591);
nor U12279 (N_12279,N_11526,N_11916);
and U12280 (N_12280,N_11694,N_11918);
and U12281 (N_12281,N_11750,N_11571);
nand U12282 (N_12282,N_11601,N_11813);
and U12283 (N_12283,N_11683,N_11777);
nand U12284 (N_12284,N_11587,N_11506);
nor U12285 (N_12285,N_11986,N_11730);
or U12286 (N_12286,N_11817,N_11670);
nand U12287 (N_12287,N_11918,N_11873);
nor U12288 (N_12288,N_11612,N_11581);
nand U12289 (N_12289,N_11921,N_11503);
nor U12290 (N_12290,N_11990,N_11812);
xor U12291 (N_12291,N_11856,N_11739);
and U12292 (N_12292,N_11594,N_11954);
nand U12293 (N_12293,N_11978,N_11764);
nor U12294 (N_12294,N_11540,N_11839);
and U12295 (N_12295,N_11754,N_11852);
nor U12296 (N_12296,N_11745,N_11737);
nor U12297 (N_12297,N_11584,N_11959);
nand U12298 (N_12298,N_11862,N_11725);
nor U12299 (N_12299,N_11817,N_11740);
and U12300 (N_12300,N_11720,N_11630);
nand U12301 (N_12301,N_11806,N_11858);
nand U12302 (N_12302,N_11692,N_11603);
nor U12303 (N_12303,N_11635,N_11895);
and U12304 (N_12304,N_11961,N_11848);
nand U12305 (N_12305,N_11986,N_11529);
nor U12306 (N_12306,N_11849,N_11979);
nor U12307 (N_12307,N_11782,N_11653);
or U12308 (N_12308,N_11642,N_11901);
nor U12309 (N_12309,N_11570,N_11637);
or U12310 (N_12310,N_11939,N_11877);
nor U12311 (N_12311,N_11919,N_11668);
or U12312 (N_12312,N_11980,N_11908);
nor U12313 (N_12313,N_11780,N_11973);
xor U12314 (N_12314,N_11568,N_11961);
and U12315 (N_12315,N_11626,N_11744);
or U12316 (N_12316,N_11510,N_11651);
and U12317 (N_12317,N_11694,N_11561);
xor U12318 (N_12318,N_11885,N_11692);
nor U12319 (N_12319,N_11698,N_11658);
nand U12320 (N_12320,N_11531,N_11545);
nor U12321 (N_12321,N_11911,N_11537);
or U12322 (N_12322,N_11898,N_11822);
nand U12323 (N_12323,N_11916,N_11598);
or U12324 (N_12324,N_11707,N_11623);
and U12325 (N_12325,N_11589,N_11804);
or U12326 (N_12326,N_11560,N_11915);
nor U12327 (N_12327,N_11969,N_11652);
nand U12328 (N_12328,N_11810,N_11675);
or U12329 (N_12329,N_11513,N_11871);
or U12330 (N_12330,N_11770,N_11973);
and U12331 (N_12331,N_11991,N_11851);
or U12332 (N_12332,N_11877,N_11977);
nor U12333 (N_12333,N_11658,N_11649);
or U12334 (N_12334,N_11745,N_11712);
or U12335 (N_12335,N_11969,N_11577);
nand U12336 (N_12336,N_11527,N_11615);
or U12337 (N_12337,N_11538,N_11650);
or U12338 (N_12338,N_11731,N_11667);
nand U12339 (N_12339,N_11886,N_11985);
and U12340 (N_12340,N_11812,N_11769);
nor U12341 (N_12341,N_11508,N_11811);
or U12342 (N_12342,N_11956,N_11664);
and U12343 (N_12343,N_11868,N_11586);
nand U12344 (N_12344,N_11759,N_11873);
nand U12345 (N_12345,N_11539,N_11891);
or U12346 (N_12346,N_11771,N_11510);
nor U12347 (N_12347,N_11778,N_11668);
nand U12348 (N_12348,N_11888,N_11507);
nor U12349 (N_12349,N_11768,N_11583);
and U12350 (N_12350,N_11993,N_11617);
and U12351 (N_12351,N_11996,N_11986);
nand U12352 (N_12352,N_11534,N_11568);
and U12353 (N_12353,N_11611,N_11567);
and U12354 (N_12354,N_11804,N_11925);
or U12355 (N_12355,N_11691,N_11671);
and U12356 (N_12356,N_11698,N_11767);
and U12357 (N_12357,N_11742,N_11616);
and U12358 (N_12358,N_11507,N_11538);
nor U12359 (N_12359,N_11546,N_11575);
and U12360 (N_12360,N_11865,N_11635);
nor U12361 (N_12361,N_11676,N_11785);
xor U12362 (N_12362,N_11824,N_11615);
and U12363 (N_12363,N_11793,N_11676);
or U12364 (N_12364,N_11992,N_11513);
or U12365 (N_12365,N_11877,N_11686);
and U12366 (N_12366,N_11565,N_11770);
or U12367 (N_12367,N_11704,N_11722);
xnor U12368 (N_12368,N_11724,N_11918);
nand U12369 (N_12369,N_11923,N_11920);
or U12370 (N_12370,N_11689,N_11986);
and U12371 (N_12371,N_11535,N_11788);
and U12372 (N_12372,N_11706,N_11802);
nand U12373 (N_12373,N_11901,N_11961);
nor U12374 (N_12374,N_11836,N_11613);
and U12375 (N_12375,N_11764,N_11609);
xnor U12376 (N_12376,N_11668,N_11612);
and U12377 (N_12377,N_11806,N_11937);
and U12378 (N_12378,N_11730,N_11994);
and U12379 (N_12379,N_11958,N_11905);
or U12380 (N_12380,N_11820,N_11519);
nand U12381 (N_12381,N_11901,N_11951);
and U12382 (N_12382,N_11896,N_11781);
and U12383 (N_12383,N_11693,N_11984);
nor U12384 (N_12384,N_11837,N_11572);
or U12385 (N_12385,N_11564,N_11733);
nor U12386 (N_12386,N_11534,N_11549);
and U12387 (N_12387,N_11927,N_11564);
nand U12388 (N_12388,N_11623,N_11859);
and U12389 (N_12389,N_11870,N_11778);
and U12390 (N_12390,N_11798,N_11972);
or U12391 (N_12391,N_11594,N_11976);
and U12392 (N_12392,N_11821,N_11567);
or U12393 (N_12393,N_11932,N_11792);
nor U12394 (N_12394,N_11959,N_11508);
nand U12395 (N_12395,N_11961,N_11962);
nor U12396 (N_12396,N_11729,N_11609);
or U12397 (N_12397,N_11734,N_11618);
or U12398 (N_12398,N_11885,N_11510);
or U12399 (N_12399,N_11989,N_11595);
xnor U12400 (N_12400,N_11751,N_11740);
nand U12401 (N_12401,N_11611,N_11921);
or U12402 (N_12402,N_11749,N_11531);
nand U12403 (N_12403,N_11695,N_11974);
or U12404 (N_12404,N_11571,N_11922);
and U12405 (N_12405,N_11645,N_11983);
and U12406 (N_12406,N_11653,N_11729);
or U12407 (N_12407,N_11661,N_11625);
nand U12408 (N_12408,N_11615,N_11681);
or U12409 (N_12409,N_11619,N_11655);
nand U12410 (N_12410,N_11574,N_11808);
nand U12411 (N_12411,N_11722,N_11915);
or U12412 (N_12412,N_11521,N_11640);
or U12413 (N_12413,N_11718,N_11760);
nor U12414 (N_12414,N_11905,N_11809);
or U12415 (N_12415,N_11706,N_11549);
nor U12416 (N_12416,N_11649,N_11681);
nor U12417 (N_12417,N_11797,N_11718);
nor U12418 (N_12418,N_11893,N_11518);
nor U12419 (N_12419,N_11990,N_11510);
or U12420 (N_12420,N_11570,N_11641);
nand U12421 (N_12421,N_11667,N_11523);
or U12422 (N_12422,N_11508,N_11774);
nor U12423 (N_12423,N_11944,N_11905);
nand U12424 (N_12424,N_11822,N_11556);
or U12425 (N_12425,N_11512,N_11579);
nor U12426 (N_12426,N_11856,N_11943);
and U12427 (N_12427,N_11876,N_11927);
and U12428 (N_12428,N_11787,N_11815);
nand U12429 (N_12429,N_11512,N_11968);
nand U12430 (N_12430,N_11506,N_11502);
nand U12431 (N_12431,N_11567,N_11729);
and U12432 (N_12432,N_11562,N_11728);
and U12433 (N_12433,N_11520,N_11994);
nor U12434 (N_12434,N_11589,N_11516);
nor U12435 (N_12435,N_11875,N_11722);
nor U12436 (N_12436,N_11694,N_11989);
nor U12437 (N_12437,N_11725,N_11617);
xnor U12438 (N_12438,N_11920,N_11829);
nand U12439 (N_12439,N_11887,N_11546);
and U12440 (N_12440,N_11952,N_11625);
nand U12441 (N_12441,N_11989,N_11964);
nand U12442 (N_12442,N_11642,N_11655);
and U12443 (N_12443,N_11881,N_11555);
nand U12444 (N_12444,N_11989,N_11677);
nand U12445 (N_12445,N_11795,N_11776);
xnor U12446 (N_12446,N_11781,N_11548);
xnor U12447 (N_12447,N_11851,N_11606);
xnor U12448 (N_12448,N_11921,N_11689);
and U12449 (N_12449,N_11628,N_11863);
nor U12450 (N_12450,N_11910,N_11680);
xor U12451 (N_12451,N_11913,N_11672);
or U12452 (N_12452,N_11864,N_11639);
or U12453 (N_12453,N_11867,N_11810);
xnor U12454 (N_12454,N_11665,N_11655);
and U12455 (N_12455,N_11616,N_11830);
nor U12456 (N_12456,N_11817,N_11525);
nand U12457 (N_12457,N_11942,N_11609);
nand U12458 (N_12458,N_11835,N_11511);
and U12459 (N_12459,N_11964,N_11770);
nand U12460 (N_12460,N_11718,N_11709);
nand U12461 (N_12461,N_11637,N_11709);
or U12462 (N_12462,N_11892,N_11884);
or U12463 (N_12463,N_11841,N_11561);
nand U12464 (N_12464,N_11942,N_11631);
and U12465 (N_12465,N_11556,N_11800);
nand U12466 (N_12466,N_11689,N_11557);
and U12467 (N_12467,N_11886,N_11546);
or U12468 (N_12468,N_11850,N_11587);
and U12469 (N_12469,N_11552,N_11570);
and U12470 (N_12470,N_11869,N_11878);
nor U12471 (N_12471,N_11500,N_11888);
and U12472 (N_12472,N_11699,N_11972);
nor U12473 (N_12473,N_11728,N_11872);
nor U12474 (N_12474,N_11560,N_11572);
and U12475 (N_12475,N_11647,N_11861);
nor U12476 (N_12476,N_11655,N_11893);
and U12477 (N_12477,N_11851,N_11799);
xnor U12478 (N_12478,N_11677,N_11755);
or U12479 (N_12479,N_11964,N_11819);
and U12480 (N_12480,N_11771,N_11904);
nand U12481 (N_12481,N_11568,N_11807);
or U12482 (N_12482,N_11650,N_11742);
nor U12483 (N_12483,N_11898,N_11808);
or U12484 (N_12484,N_11584,N_11780);
and U12485 (N_12485,N_11677,N_11685);
xor U12486 (N_12486,N_11748,N_11803);
xor U12487 (N_12487,N_11673,N_11721);
or U12488 (N_12488,N_11593,N_11714);
nand U12489 (N_12489,N_11603,N_11700);
or U12490 (N_12490,N_11655,N_11565);
xnor U12491 (N_12491,N_11818,N_11943);
or U12492 (N_12492,N_11914,N_11891);
nand U12493 (N_12493,N_11969,N_11785);
nor U12494 (N_12494,N_11549,N_11605);
or U12495 (N_12495,N_11809,N_11848);
and U12496 (N_12496,N_11926,N_11661);
nand U12497 (N_12497,N_11692,N_11908);
nand U12498 (N_12498,N_11738,N_11950);
xor U12499 (N_12499,N_11714,N_11997);
and U12500 (N_12500,N_12000,N_12140);
and U12501 (N_12501,N_12312,N_12478);
and U12502 (N_12502,N_12320,N_12180);
nor U12503 (N_12503,N_12106,N_12104);
nor U12504 (N_12504,N_12326,N_12357);
nor U12505 (N_12505,N_12285,N_12255);
nand U12506 (N_12506,N_12491,N_12336);
or U12507 (N_12507,N_12277,N_12231);
nand U12508 (N_12508,N_12123,N_12243);
nand U12509 (N_12509,N_12211,N_12324);
nand U12510 (N_12510,N_12471,N_12012);
nor U12511 (N_12511,N_12168,N_12026);
and U12512 (N_12512,N_12011,N_12225);
nand U12513 (N_12513,N_12025,N_12189);
xor U12514 (N_12514,N_12114,N_12030);
or U12515 (N_12515,N_12193,N_12179);
or U12516 (N_12516,N_12328,N_12128);
and U12517 (N_12517,N_12110,N_12296);
or U12518 (N_12518,N_12341,N_12239);
nand U12519 (N_12519,N_12448,N_12349);
xnor U12520 (N_12520,N_12150,N_12160);
nor U12521 (N_12521,N_12437,N_12272);
xnor U12522 (N_12522,N_12356,N_12433);
xor U12523 (N_12523,N_12416,N_12032);
nand U12524 (N_12524,N_12379,N_12006);
or U12525 (N_12525,N_12236,N_12483);
and U12526 (N_12526,N_12352,N_12094);
nor U12527 (N_12527,N_12286,N_12013);
nand U12528 (N_12528,N_12283,N_12252);
nand U12529 (N_12529,N_12315,N_12474);
nand U12530 (N_12530,N_12139,N_12313);
and U12531 (N_12531,N_12181,N_12138);
nor U12532 (N_12532,N_12120,N_12171);
and U12533 (N_12533,N_12464,N_12308);
and U12534 (N_12534,N_12190,N_12216);
and U12535 (N_12535,N_12292,N_12327);
xnor U12536 (N_12536,N_12396,N_12268);
nand U12537 (N_12537,N_12438,N_12468);
or U12538 (N_12538,N_12257,N_12143);
nor U12539 (N_12539,N_12169,N_12302);
and U12540 (N_12540,N_12485,N_12348);
and U12541 (N_12541,N_12297,N_12037);
and U12542 (N_12542,N_12465,N_12333);
nand U12543 (N_12543,N_12183,N_12420);
or U12544 (N_12544,N_12119,N_12303);
and U12545 (N_12545,N_12295,N_12004);
nor U12546 (N_12546,N_12067,N_12423);
and U12547 (N_12547,N_12383,N_12487);
or U12548 (N_12548,N_12425,N_12126);
and U12549 (N_12549,N_12430,N_12362);
nand U12550 (N_12550,N_12080,N_12144);
nand U12551 (N_12551,N_12469,N_12056);
xor U12552 (N_12552,N_12184,N_12112);
or U12553 (N_12553,N_12164,N_12102);
nand U12554 (N_12554,N_12499,N_12061);
or U12555 (N_12555,N_12064,N_12460);
nor U12556 (N_12556,N_12365,N_12009);
and U12557 (N_12557,N_12251,N_12412);
nand U12558 (N_12558,N_12085,N_12335);
or U12559 (N_12559,N_12288,N_12463);
or U12560 (N_12560,N_12208,N_12316);
or U12561 (N_12561,N_12209,N_12141);
and U12562 (N_12562,N_12482,N_12087);
or U12563 (N_12563,N_12381,N_12219);
nand U12564 (N_12564,N_12230,N_12353);
xnor U12565 (N_12565,N_12175,N_12421);
and U12566 (N_12566,N_12446,N_12337);
or U12567 (N_12567,N_12311,N_12260);
or U12568 (N_12568,N_12456,N_12059);
nor U12569 (N_12569,N_12235,N_12279);
nor U12570 (N_12570,N_12426,N_12253);
nor U12571 (N_12571,N_12493,N_12237);
or U12572 (N_12572,N_12462,N_12165);
nor U12573 (N_12573,N_12151,N_12200);
nor U12574 (N_12574,N_12490,N_12125);
and U12575 (N_12575,N_12137,N_12476);
nor U12576 (N_12576,N_12449,N_12191);
nor U12577 (N_12577,N_12135,N_12173);
nor U12578 (N_12578,N_12095,N_12041);
and U12579 (N_12579,N_12192,N_12027);
nand U12580 (N_12580,N_12489,N_12355);
nor U12581 (N_12581,N_12305,N_12049);
and U12582 (N_12582,N_12254,N_12178);
nand U12583 (N_12583,N_12293,N_12452);
or U12584 (N_12584,N_12158,N_12222);
and U12585 (N_12585,N_12461,N_12334);
nor U12586 (N_12586,N_12401,N_12284);
nor U12587 (N_12587,N_12229,N_12280);
and U12588 (N_12588,N_12370,N_12220);
xor U12589 (N_12589,N_12132,N_12339);
xnor U12590 (N_12590,N_12016,N_12435);
nor U12591 (N_12591,N_12081,N_12246);
or U12592 (N_12592,N_12122,N_12318);
and U12593 (N_12593,N_12466,N_12345);
or U12594 (N_12594,N_12115,N_12459);
xnor U12595 (N_12595,N_12291,N_12176);
nor U12596 (N_12596,N_12270,N_12261);
or U12597 (N_12597,N_12198,N_12166);
or U12598 (N_12598,N_12325,N_12319);
and U12599 (N_12599,N_12071,N_12458);
xor U12600 (N_12600,N_12188,N_12263);
and U12601 (N_12601,N_12307,N_12215);
nor U12602 (N_12602,N_12098,N_12042);
nand U12603 (N_12603,N_12428,N_12258);
or U12604 (N_12604,N_12343,N_12149);
and U12605 (N_12605,N_12083,N_12107);
nor U12606 (N_12606,N_12274,N_12073);
nor U12607 (N_12607,N_12203,N_12360);
or U12608 (N_12608,N_12405,N_12177);
xor U12609 (N_12609,N_12155,N_12228);
nor U12610 (N_12610,N_12350,N_12124);
or U12611 (N_12611,N_12317,N_12391);
xor U12612 (N_12612,N_12245,N_12148);
or U12613 (N_12613,N_12267,N_12340);
and U12614 (N_12614,N_12033,N_12276);
and U12615 (N_12615,N_12494,N_12197);
nand U12616 (N_12616,N_12497,N_12029);
and U12617 (N_12617,N_12403,N_12024);
or U12618 (N_12618,N_12172,N_12413);
and U12619 (N_12619,N_12444,N_12127);
and U12620 (N_12620,N_12262,N_12060);
nor U12621 (N_12621,N_12019,N_12407);
and U12622 (N_12622,N_12048,N_12062);
nor U12623 (N_12623,N_12475,N_12035);
nor U12624 (N_12624,N_12118,N_12108);
and U12625 (N_12625,N_12068,N_12300);
nor U12626 (N_12626,N_12417,N_12408);
and U12627 (N_12627,N_12058,N_12218);
or U12628 (N_12628,N_12014,N_12450);
xor U12629 (N_12629,N_12418,N_12378);
nor U12630 (N_12630,N_12039,N_12306);
nor U12631 (N_12631,N_12020,N_12206);
nor U12632 (N_12632,N_12156,N_12358);
nand U12633 (N_12633,N_12109,N_12170);
nand U12634 (N_12634,N_12367,N_12445);
and U12635 (N_12635,N_12136,N_12199);
or U12636 (N_12636,N_12142,N_12113);
or U12637 (N_12637,N_12046,N_12447);
nor U12638 (N_12638,N_12034,N_12008);
and U12639 (N_12639,N_12131,N_12372);
or U12640 (N_12640,N_12082,N_12289);
or U12641 (N_12641,N_12099,N_12347);
nor U12642 (N_12642,N_12065,N_12051);
nor U12643 (N_12643,N_12375,N_12038);
or U12644 (N_12644,N_12031,N_12174);
nor U12645 (N_12645,N_12351,N_12159);
and U12646 (N_12646,N_12217,N_12153);
and U12647 (N_12647,N_12147,N_12233);
and U12648 (N_12648,N_12392,N_12117);
and U12649 (N_12649,N_12371,N_12227);
and U12650 (N_12650,N_12397,N_12201);
or U12651 (N_12651,N_12301,N_12278);
nand U12652 (N_12652,N_12384,N_12386);
and U12653 (N_12653,N_12338,N_12388);
nand U12654 (N_12654,N_12409,N_12380);
nor U12655 (N_12655,N_12439,N_12238);
nand U12656 (N_12656,N_12390,N_12436);
or U12657 (N_12657,N_12406,N_12097);
and U12658 (N_12658,N_12385,N_12361);
nand U12659 (N_12659,N_12086,N_12480);
xnor U12660 (N_12660,N_12167,N_12498);
nand U12661 (N_12661,N_12486,N_12047);
nand U12662 (N_12662,N_12434,N_12093);
nand U12663 (N_12663,N_12454,N_12373);
or U12664 (N_12664,N_12275,N_12299);
nand U12665 (N_12665,N_12273,N_12207);
nand U12666 (N_12666,N_12427,N_12111);
and U12667 (N_12667,N_12089,N_12074);
nor U12668 (N_12668,N_12072,N_12044);
nor U12669 (N_12669,N_12022,N_12023);
or U12670 (N_12670,N_12481,N_12269);
nor U12671 (N_12671,N_12134,N_12241);
nor U12672 (N_12672,N_12028,N_12146);
nor U12673 (N_12673,N_12100,N_12382);
or U12674 (N_12674,N_12212,N_12018);
nor U12675 (N_12675,N_12096,N_12399);
or U12676 (N_12676,N_12294,N_12005);
nand U12677 (N_12677,N_12342,N_12354);
and U12678 (N_12678,N_12457,N_12363);
nor U12679 (N_12679,N_12496,N_12232);
xor U12680 (N_12680,N_12344,N_12213);
nor U12681 (N_12681,N_12431,N_12271);
nor U12682 (N_12682,N_12078,N_12451);
nand U12683 (N_12683,N_12053,N_12331);
nand U12684 (N_12684,N_12321,N_12092);
nor U12685 (N_12685,N_12052,N_12376);
and U12686 (N_12686,N_12387,N_12453);
and U12687 (N_12687,N_12214,N_12057);
nand U12688 (N_12688,N_12369,N_12070);
or U12689 (N_12689,N_12411,N_12202);
nand U12690 (N_12690,N_12204,N_12130);
nand U12691 (N_12691,N_12003,N_12250);
nor U12692 (N_12692,N_12419,N_12414);
nor U12693 (N_12693,N_12374,N_12442);
and U12694 (N_12694,N_12393,N_12234);
nand U12695 (N_12695,N_12332,N_12040);
nand U12696 (N_12696,N_12145,N_12054);
nand U12697 (N_12697,N_12323,N_12079);
or U12698 (N_12698,N_12247,N_12398);
or U12699 (N_12699,N_12157,N_12162);
nor U12700 (N_12700,N_12259,N_12440);
xor U12701 (N_12701,N_12224,N_12121);
nor U12702 (N_12702,N_12256,N_12205);
or U12703 (N_12703,N_12455,N_12395);
or U12704 (N_12704,N_12248,N_12240);
nand U12705 (N_12705,N_12077,N_12484);
and U12706 (N_12706,N_12377,N_12163);
and U12707 (N_12707,N_12488,N_12364);
and U12708 (N_12708,N_12154,N_12330);
nor U12709 (N_12709,N_12021,N_12402);
or U12710 (N_12710,N_12043,N_12329);
nor U12711 (N_12711,N_12477,N_12010);
nor U12712 (N_12712,N_12105,N_12244);
or U12713 (N_12713,N_12015,N_12394);
and U12714 (N_12714,N_12185,N_12467);
and U12715 (N_12715,N_12088,N_12314);
and U12716 (N_12716,N_12322,N_12090);
or U12717 (N_12717,N_12410,N_12287);
and U12718 (N_12718,N_12422,N_12441);
nor U12719 (N_12719,N_12101,N_12346);
or U12720 (N_12720,N_12194,N_12069);
and U12721 (N_12721,N_12055,N_12007);
or U12722 (N_12722,N_12195,N_12187);
or U12723 (N_12723,N_12182,N_12495);
or U12724 (N_12724,N_12298,N_12429);
nor U12725 (N_12725,N_12264,N_12152);
nor U12726 (N_12726,N_12415,N_12186);
nor U12727 (N_12727,N_12492,N_12424);
xnor U12728 (N_12728,N_12368,N_12001);
and U12729 (N_12729,N_12036,N_12310);
xnor U12730 (N_12730,N_12066,N_12063);
xnor U12731 (N_12731,N_12443,N_12266);
xor U12732 (N_12732,N_12404,N_12133);
or U12733 (N_12733,N_12366,N_12075);
nor U12734 (N_12734,N_12076,N_12309);
or U12735 (N_12735,N_12282,N_12210);
or U12736 (N_12736,N_12226,N_12359);
and U12737 (N_12737,N_12400,N_12223);
or U12738 (N_12738,N_12281,N_12129);
or U12739 (N_12739,N_12045,N_12470);
or U12740 (N_12740,N_12084,N_12242);
or U12741 (N_12741,N_12221,N_12091);
nand U12742 (N_12742,N_12103,N_12304);
or U12743 (N_12743,N_12389,N_12050);
nor U12744 (N_12744,N_12196,N_12472);
nand U12745 (N_12745,N_12473,N_12290);
nor U12746 (N_12746,N_12479,N_12002);
and U12747 (N_12747,N_12017,N_12249);
nand U12748 (N_12748,N_12432,N_12116);
and U12749 (N_12749,N_12161,N_12265);
nand U12750 (N_12750,N_12142,N_12168);
nand U12751 (N_12751,N_12405,N_12096);
or U12752 (N_12752,N_12293,N_12408);
nand U12753 (N_12753,N_12417,N_12446);
xnor U12754 (N_12754,N_12453,N_12047);
nand U12755 (N_12755,N_12381,N_12062);
nand U12756 (N_12756,N_12356,N_12075);
nand U12757 (N_12757,N_12379,N_12044);
and U12758 (N_12758,N_12318,N_12391);
nand U12759 (N_12759,N_12060,N_12109);
and U12760 (N_12760,N_12326,N_12251);
xor U12761 (N_12761,N_12476,N_12306);
and U12762 (N_12762,N_12179,N_12207);
or U12763 (N_12763,N_12364,N_12300);
xor U12764 (N_12764,N_12407,N_12039);
and U12765 (N_12765,N_12381,N_12404);
or U12766 (N_12766,N_12114,N_12449);
and U12767 (N_12767,N_12390,N_12145);
xor U12768 (N_12768,N_12007,N_12397);
or U12769 (N_12769,N_12376,N_12476);
nor U12770 (N_12770,N_12244,N_12328);
xor U12771 (N_12771,N_12163,N_12383);
nand U12772 (N_12772,N_12085,N_12322);
or U12773 (N_12773,N_12068,N_12227);
and U12774 (N_12774,N_12069,N_12068);
nand U12775 (N_12775,N_12316,N_12426);
or U12776 (N_12776,N_12384,N_12375);
nand U12777 (N_12777,N_12040,N_12300);
nand U12778 (N_12778,N_12095,N_12051);
or U12779 (N_12779,N_12238,N_12412);
or U12780 (N_12780,N_12042,N_12346);
nand U12781 (N_12781,N_12143,N_12154);
nand U12782 (N_12782,N_12087,N_12263);
nor U12783 (N_12783,N_12227,N_12116);
and U12784 (N_12784,N_12095,N_12168);
or U12785 (N_12785,N_12310,N_12133);
nor U12786 (N_12786,N_12131,N_12134);
nor U12787 (N_12787,N_12215,N_12422);
xnor U12788 (N_12788,N_12451,N_12364);
nand U12789 (N_12789,N_12418,N_12454);
nand U12790 (N_12790,N_12416,N_12394);
nor U12791 (N_12791,N_12362,N_12023);
xor U12792 (N_12792,N_12127,N_12287);
and U12793 (N_12793,N_12012,N_12382);
or U12794 (N_12794,N_12340,N_12457);
or U12795 (N_12795,N_12001,N_12402);
nand U12796 (N_12796,N_12164,N_12456);
and U12797 (N_12797,N_12423,N_12433);
and U12798 (N_12798,N_12097,N_12430);
or U12799 (N_12799,N_12353,N_12331);
nor U12800 (N_12800,N_12051,N_12187);
nand U12801 (N_12801,N_12286,N_12193);
nor U12802 (N_12802,N_12045,N_12472);
nand U12803 (N_12803,N_12017,N_12222);
xnor U12804 (N_12804,N_12378,N_12363);
nor U12805 (N_12805,N_12314,N_12039);
or U12806 (N_12806,N_12160,N_12492);
nor U12807 (N_12807,N_12314,N_12496);
or U12808 (N_12808,N_12041,N_12112);
nand U12809 (N_12809,N_12072,N_12033);
nand U12810 (N_12810,N_12277,N_12369);
and U12811 (N_12811,N_12328,N_12309);
and U12812 (N_12812,N_12056,N_12353);
or U12813 (N_12813,N_12243,N_12081);
nor U12814 (N_12814,N_12441,N_12335);
and U12815 (N_12815,N_12347,N_12365);
xor U12816 (N_12816,N_12312,N_12043);
nor U12817 (N_12817,N_12139,N_12073);
nand U12818 (N_12818,N_12050,N_12348);
and U12819 (N_12819,N_12097,N_12235);
or U12820 (N_12820,N_12049,N_12399);
or U12821 (N_12821,N_12163,N_12124);
nand U12822 (N_12822,N_12011,N_12069);
and U12823 (N_12823,N_12320,N_12045);
xnor U12824 (N_12824,N_12053,N_12201);
or U12825 (N_12825,N_12494,N_12482);
and U12826 (N_12826,N_12030,N_12292);
or U12827 (N_12827,N_12072,N_12482);
nor U12828 (N_12828,N_12096,N_12336);
and U12829 (N_12829,N_12059,N_12340);
or U12830 (N_12830,N_12345,N_12444);
and U12831 (N_12831,N_12148,N_12475);
or U12832 (N_12832,N_12467,N_12408);
or U12833 (N_12833,N_12154,N_12389);
and U12834 (N_12834,N_12291,N_12236);
and U12835 (N_12835,N_12250,N_12127);
nor U12836 (N_12836,N_12167,N_12267);
nand U12837 (N_12837,N_12350,N_12364);
and U12838 (N_12838,N_12238,N_12107);
nor U12839 (N_12839,N_12463,N_12271);
and U12840 (N_12840,N_12118,N_12181);
xor U12841 (N_12841,N_12440,N_12143);
nand U12842 (N_12842,N_12052,N_12305);
or U12843 (N_12843,N_12491,N_12280);
or U12844 (N_12844,N_12064,N_12140);
and U12845 (N_12845,N_12312,N_12445);
and U12846 (N_12846,N_12259,N_12256);
nand U12847 (N_12847,N_12040,N_12290);
nor U12848 (N_12848,N_12173,N_12122);
or U12849 (N_12849,N_12497,N_12230);
and U12850 (N_12850,N_12336,N_12057);
or U12851 (N_12851,N_12176,N_12398);
and U12852 (N_12852,N_12299,N_12144);
xor U12853 (N_12853,N_12454,N_12029);
or U12854 (N_12854,N_12393,N_12191);
nor U12855 (N_12855,N_12385,N_12351);
and U12856 (N_12856,N_12297,N_12167);
and U12857 (N_12857,N_12231,N_12097);
nand U12858 (N_12858,N_12281,N_12061);
nand U12859 (N_12859,N_12197,N_12110);
or U12860 (N_12860,N_12068,N_12011);
nor U12861 (N_12861,N_12073,N_12280);
nor U12862 (N_12862,N_12299,N_12325);
xor U12863 (N_12863,N_12017,N_12111);
or U12864 (N_12864,N_12283,N_12022);
nand U12865 (N_12865,N_12195,N_12279);
or U12866 (N_12866,N_12371,N_12397);
nor U12867 (N_12867,N_12138,N_12226);
nand U12868 (N_12868,N_12114,N_12417);
nor U12869 (N_12869,N_12041,N_12306);
and U12870 (N_12870,N_12238,N_12358);
and U12871 (N_12871,N_12430,N_12195);
nand U12872 (N_12872,N_12098,N_12237);
xnor U12873 (N_12873,N_12477,N_12243);
nand U12874 (N_12874,N_12015,N_12175);
or U12875 (N_12875,N_12436,N_12065);
and U12876 (N_12876,N_12109,N_12449);
nand U12877 (N_12877,N_12093,N_12078);
nor U12878 (N_12878,N_12377,N_12195);
and U12879 (N_12879,N_12232,N_12212);
nand U12880 (N_12880,N_12225,N_12043);
or U12881 (N_12881,N_12023,N_12446);
nand U12882 (N_12882,N_12185,N_12238);
nand U12883 (N_12883,N_12176,N_12165);
nor U12884 (N_12884,N_12480,N_12441);
nor U12885 (N_12885,N_12044,N_12033);
nand U12886 (N_12886,N_12494,N_12351);
nor U12887 (N_12887,N_12141,N_12095);
or U12888 (N_12888,N_12326,N_12464);
or U12889 (N_12889,N_12218,N_12145);
and U12890 (N_12890,N_12020,N_12015);
and U12891 (N_12891,N_12493,N_12496);
or U12892 (N_12892,N_12465,N_12135);
nor U12893 (N_12893,N_12209,N_12145);
or U12894 (N_12894,N_12014,N_12131);
or U12895 (N_12895,N_12425,N_12355);
nor U12896 (N_12896,N_12276,N_12068);
or U12897 (N_12897,N_12058,N_12304);
nor U12898 (N_12898,N_12080,N_12025);
nor U12899 (N_12899,N_12311,N_12361);
nand U12900 (N_12900,N_12409,N_12273);
or U12901 (N_12901,N_12454,N_12442);
or U12902 (N_12902,N_12143,N_12141);
nand U12903 (N_12903,N_12459,N_12244);
nand U12904 (N_12904,N_12005,N_12109);
nor U12905 (N_12905,N_12235,N_12073);
nor U12906 (N_12906,N_12039,N_12189);
and U12907 (N_12907,N_12243,N_12201);
and U12908 (N_12908,N_12070,N_12351);
nand U12909 (N_12909,N_12255,N_12418);
and U12910 (N_12910,N_12364,N_12289);
or U12911 (N_12911,N_12353,N_12211);
and U12912 (N_12912,N_12346,N_12171);
xnor U12913 (N_12913,N_12241,N_12091);
nand U12914 (N_12914,N_12359,N_12176);
xor U12915 (N_12915,N_12288,N_12159);
nor U12916 (N_12916,N_12093,N_12211);
nand U12917 (N_12917,N_12073,N_12042);
and U12918 (N_12918,N_12113,N_12103);
and U12919 (N_12919,N_12061,N_12273);
and U12920 (N_12920,N_12009,N_12455);
or U12921 (N_12921,N_12124,N_12241);
nand U12922 (N_12922,N_12286,N_12182);
and U12923 (N_12923,N_12434,N_12270);
or U12924 (N_12924,N_12397,N_12115);
and U12925 (N_12925,N_12155,N_12321);
xor U12926 (N_12926,N_12171,N_12280);
nor U12927 (N_12927,N_12365,N_12263);
nor U12928 (N_12928,N_12267,N_12312);
or U12929 (N_12929,N_12235,N_12064);
and U12930 (N_12930,N_12301,N_12216);
xor U12931 (N_12931,N_12178,N_12145);
and U12932 (N_12932,N_12405,N_12247);
nor U12933 (N_12933,N_12277,N_12222);
nor U12934 (N_12934,N_12328,N_12195);
or U12935 (N_12935,N_12414,N_12116);
nor U12936 (N_12936,N_12118,N_12294);
or U12937 (N_12937,N_12078,N_12487);
nand U12938 (N_12938,N_12213,N_12011);
nor U12939 (N_12939,N_12471,N_12310);
and U12940 (N_12940,N_12079,N_12136);
and U12941 (N_12941,N_12075,N_12058);
nor U12942 (N_12942,N_12098,N_12435);
nand U12943 (N_12943,N_12009,N_12010);
nor U12944 (N_12944,N_12242,N_12111);
and U12945 (N_12945,N_12498,N_12126);
and U12946 (N_12946,N_12304,N_12139);
xor U12947 (N_12947,N_12310,N_12335);
or U12948 (N_12948,N_12495,N_12256);
xor U12949 (N_12949,N_12280,N_12139);
nor U12950 (N_12950,N_12413,N_12059);
and U12951 (N_12951,N_12392,N_12073);
nand U12952 (N_12952,N_12390,N_12234);
and U12953 (N_12953,N_12183,N_12499);
or U12954 (N_12954,N_12061,N_12020);
and U12955 (N_12955,N_12008,N_12149);
xnor U12956 (N_12956,N_12106,N_12295);
xnor U12957 (N_12957,N_12107,N_12411);
nand U12958 (N_12958,N_12276,N_12188);
or U12959 (N_12959,N_12259,N_12193);
nor U12960 (N_12960,N_12389,N_12319);
nor U12961 (N_12961,N_12415,N_12497);
or U12962 (N_12962,N_12318,N_12497);
nor U12963 (N_12963,N_12245,N_12143);
and U12964 (N_12964,N_12281,N_12047);
xnor U12965 (N_12965,N_12142,N_12334);
and U12966 (N_12966,N_12025,N_12421);
and U12967 (N_12967,N_12144,N_12294);
nand U12968 (N_12968,N_12193,N_12206);
or U12969 (N_12969,N_12042,N_12034);
or U12970 (N_12970,N_12420,N_12429);
or U12971 (N_12971,N_12327,N_12310);
xor U12972 (N_12972,N_12489,N_12266);
and U12973 (N_12973,N_12173,N_12106);
and U12974 (N_12974,N_12438,N_12138);
nor U12975 (N_12975,N_12044,N_12288);
xor U12976 (N_12976,N_12260,N_12331);
xor U12977 (N_12977,N_12248,N_12074);
or U12978 (N_12978,N_12214,N_12151);
nand U12979 (N_12979,N_12402,N_12020);
nand U12980 (N_12980,N_12223,N_12143);
nor U12981 (N_12981,N_12010,N_12359);
nor U12982 (N_12982,N_12382,N_12325);
xnor U12983 (N_12983,N_12442,N_12369);
or U12984 (N_12984,N_12315,N_12334);
nand U12985 (N_12985,N_12086,N_12123);
nand U12986 (N_12986,N_12226,N_12140);
xnor U12987 (N_12987,N_12154,N_12478);
or U12988 (N_12988,N_12343,N_12125);
nor U12989 (N_12989,N_12427,N_12094);
nor U12990 (N_12990,N_12415,N_12118);
nor U12991 (N_12991,N_12312,N_12026);
nor U12992 (N_12992,N_12185,N_12274);
nand U12993 (N_12993,N_12067,N_12397);
and U12994 (N_12994,N_12050,N_12034);
nand U12995 (N_12995,N_12137,N_12124);
nor U12996 (N_12996,N_12076,N_12193);
nand U12997 (N_12997,N_12103,N_12403);
nor U12998 (N_12998,N_12210,N_12021);
or U12999 (N_12999,N_12005,N_12404);
or U13000 (N_13000,N_12683,N_12625);
xnor U13001 (N_13001,N_12569,N_12973);
and U13002 (N_13002,N_12642,N_12589);
nand U13003 (N_13003,N_12972,N_12676);
nand U13004 (N_13004,N_12885,N_12701);
nand U13005 (N_13005,N_12700,N_12862);
and U13006 (N_13006,N_12922,N_12719);
xor U13007 (N_13007,N_12969,N_12735);
nor U13008 (N_13008,N_12587,N_12983);
nand U13009 (N_13009,N_12738,N_12779);
or U13010 (N_13010,N_12646,N_12889);
xor U13011 (N_13011,N_12825,N_12915);
nor U13012 (N_13012,N_12685,N_12696);
nor U13013 (N_13013,N_12766,N_12952);
nand U13014 (N_13014,N_12824,N_12596);
nand U13015 (N_13015,N_12560,N_12544);
nor U13016 (N_13016,N_12546,N_12871);
or U13017 (N_13017,N_12573,N_12925);
or U13018 (N_13018,N_12783,N_12511);
and U13019 (N_13019,N_12697,N_12883);
nand U13020 (N_13020,N_12718,N_12749);
and U13021 (N_13021,N_12599,N_12899);
nor U13022 (N_13022,N_12965,N_12895);
nand U13023 (N_13023,N_12561,N_12841);
and U13024 (N_13024,N_12665,N_12519);
nand U13025 (N_13025,N_12537,N_12687);
or U13026 (N_13026,N_12980,N_12928);
nand U13027 (N_13027,N_12624,N_12628);
nand U13028 (N_13028,N_12847,N_12612);
and U13029 (N_13029,N_12678,N_12880);
nor U13030 (N_13030,N_12814,N_12518);
nor U13031 (N_13031,N_12984,N_12887);
nand U13032 (N_13032,N_12706,N_12861);
xor U13033 (N_13033,N_12714,N_12745);
nor U13034 (N_13034,N_12954,N_12759);
or U13035 (N_13035,N_12660,N_12822);
and U13036 (N_13036,N_12635,N_12740);
nand U13037 (N_13037,N_12762,N_12727);
and U13038 (N_13038,N_12803,N_12852);
or U13039 (N_13039,N_12757,N_12831);
nor U13040 (N_13040,N_12939,N_12967);
nand U13041 (N_13041,N_12607,N_12975);
nor U13042 (N_13042,N_12555,N_12715);
nand U13043 (N_13043,N_12784,N_12842);
or U13044 (N_13044,N_12744,N_12594);
nand U13045 (N_13045,N_12894,N_12776);
and U13046 (N_13046,N_12901,N_12558);
xnor U13047 (N_13047,N_12731,N_12838);
and U13048 (N_13048,N_12898,N_12987);
nand U13049 (N_13049,N_12817,N_12750);
or U13050 (N_13050,N_12795,N_12811);
or U13051 (N_13051,N_12516,N_12668);
and U13052 (N_13052,N_12986,N_12963);
and U13053 (N_13053,N_12652,N_12637);
xor U13054 (N_13054,N_12548,N_12742);
or U13055 (N_13055,N_12720,N_12912);
nand U13056 (N_13056,N_12633,N_12802);
xnor U13057 (N_13057,N_12680,N_12746);
nor U13058 (N_13058,N_12846,N_12763);
or U13059 (N_13059,N_12961,N_12734);
nor U13060 (N_13060,N_12834,N_12931);
or U13061 (N_13061,N_12525,N_12992);
and U13062 (N_13062,N_12921,N_12869);
nand U13063 (N_13063,N_12835,N_12858);
nand U13064 (N_13064,N_12688,N_12579);
or U13065 (N_13065,N_12705,N_12760);
nor U13066 (N_13066,N_12608,N_12541);
and U13067 (N_13067,N_12998,N_12716);
nor U13068 (N_13068,N_12654,N_12995);
or U13069 (N_13069,N_12991,N_12593);
nand U13070 (N_13070,N_12551,N_12865);
nor U13071 (N_13071,N_12777,N_12845);
and U13072 (N_13072,N_12917,N_12989);
nand U13073 (N_13073,N_12513,N_12630);
and U13074 (N_13074,N_12606,N_12512);
and U13075 (N_13075,N_12591,N_12725);
or U13076 (N_13076,N_12753,N_12553);
or U13077 (N_13077,N_12819,N_12900);
nand U13078 (N_13078,N_12509,N_12528);
or U13079 (N_13079,N_12661,N_12855);
or U13080 (N_13080,N_12547,N_12966);
or U13081 (N_13081,N_12710,N_12780);
and U13082 (N_13082,N_12896,N_12545);
nand U13083 (N_13083,N_12684,N_12543);
nor U13084 (N_13084,N_12572,N_12810);
nand U13085 (N_13085,N_12857,N_12844);
nor U13086 (N_13086,N_12707,N_12532);
nand U13087 (N_13087,N_12786,N_12876);
or U13088 (N_13088,N_12761,N_12892);
and U13089 (N_13089,N_12631,N_12935);
or U13090 (N_13090,N_12911,N_12743);
nor U13091 (N_13091,N_12686,N_12667);
nand U13092 (N_13092,N_12897,N_12581);
nor U13093 (N_13093,N_12679,N_12778);
xor U13094 (N_13094,N_12657,N_12805);
nand U13095 (N_13095,N_12508,N_12626);
nand U13096 (N_13096,N_12829,N_12702);
or U13097 (N_13097,N_12976,N_12940);
or U13098 (N_13098,N_12658,N_12577);
nand U13099 (N_13099,N_12879,N_12774);
and U13100 (N_13100,N_12893,N_12874);
nor U13101 (N_13101,N_12588,N_12526);
or U13102 (N_13102,N_12693,N_12682);
nor U13103 (N_13103,N_12924,N_12755);
or U13104 (N_13104,N_12664,N_12632);
or U13105 (N_13105,N_12960,N_12517);
nor U13106 (N_13106,N_12908,N_12875);
nor U13107 (N_13107,N_12704,N_12971);
and U13108 (N_13108,N_12953,N_12767);
nor U13109 (N_13109,N_12501,N_12785);
or U13110 (N_13110,N_12914,N_12656);
nor U13111 (N_13111,N_12933,N_12938);
nor U13112 (N_13112,N_12616,N_12946);
nor U13113 (N_13113,N_12808,N_12634);
nor U13114 (N_13114,N_12691,N_12751);
nor U13115 (N_13115,N_12773,N_12775);
nand U13116 (N_13116,N_12799,N_12823);
and U13117 (N_13117,N_12698,N_12641);
and U13118 (N_13118,N_12789,N_12721);
nand U13119 (N_13119,N_12979,N_12993);
and U13120 (N_13120,N_12828,N_12540);
and U13121 (N_13121,N_12968,N_12574);
or U13122 (N_13122,N_12527,N_12671);
nor U13123 (N_13123,N_12836,N_12843);
and U13124 (N_13124,N_12945,N_12807);
nand U13125 (N_13125,N_12982,N_12524);
and U13126 (N_13126,N_12985,N_12709);
nor U13127 (N_13127,N_12730,N_12694);
and U13128 (N_13128,N_12563,N_12756);
nand U13129 (N_13129,N_12659,N_12595);
and U13130 (N_13130,N_12650,N_12813);
nand U13131 (N_13131,N_12891,N_12997);
nor U13132 (N_13132,N_12820,N_12601);
nand U13133 (N_13133,N_12653,N_12929);
or U13134 (N_13134,N_12673,N_12839);
xor U13135 (N_13135,N_12723,N_12506);
nor U13136 (N_13136,N_12959,N_12794);
and U13137 (N_13137,N_12765,N_12618);
xor U13138 (N_13138,N_12622,N_12796);
nor U13139 (N_13139,N_12739,N_12534);
nor U13140 (N_13140,N_12958,N_12964);
nor U13141 (N_13141,N_12539,N_12583);
and U13142 (N_13142,N_12977,N_12870);
or U13143 (N_13143,N_12833,N_12947);
nor U13144 (N_13144,N_12826,N_12941);
or U13145 (N_13145,N_12918,N_12830);
nor U13146 (N_13146,N_12978,N_12856);
and U13147 (N_13147,N_12884,N_12617);
or U13148 (N_13148,N_12726,N_12837);
and U13149 (N_13149,N_12535,N_12955);
nor U13150 (N_13150,N_12597,N_12800);
and U13151 (N_13151,N_12930,N_12866);
nor U13152 (N_13152,N_12565,N_12890);
nor U13153 (N_13153,N_12643,N_12638);
xor U13154 (N_13154,N_12598,N_12559);
nand U13155 (N_13155,N_12566,N_12913);
nor U13156 (N_13156,N_12717,N_12672);
and U13157 (N_13157,N_12620,N_12840);
nand U13158 (N_13158,N_12590,N_12926);
nand U13159 (N_13159,N_12951,N_12923);
or U13160 (N_13160,N_12957,N_12699);
or U13161 (N_13161,N_12562,N_12712);
or U13162 (N_13162,N_12550,N_12575);
and U13163 (N_13163,N_12904,N_12741);
nand U13164 (N_13164,N_12793,N_12907);
nand U13165 (N_13165,N_12651,N_12881);
nor U13166 (N_13166,N_12549,N_12722);
nor U13167 (N_13167,N_12797,N_12949);
or U13168 (N_13168,N_12640,N_12906);
nor U13169 (N_13169,N_12724,N_12956);
nor U13170 (N_13170,N_12747,N_12648);
and U13171 (N_13171,N_12703,N_12732);
or U13172 (N_13172,N_12586,N_12848);
or U13173 (N_13173,N_12663,N_12832);
nor U13174 (N_13174,N_12781,N_12737);
or U13175 (N_13175,N_12769,N_12804);
nor U13176 (N_13176,N_12859,N_12920);
xor U13177 (N_13177,N_12567,N_12950);
xnor U13178 (N_13178,N_12790,N_12554);
or U13179 (N_13179,N_12576,N_12981);
or U13180 (N_13180,N_12849,N_12645);
or U13181 (N_13181,N_12932,N_12568);
and U13182 (N_13182,N_12571,N_12728);
or U13183 (N_13183,N_12690,N_12729);
nor U13184 (N_13184,N_12999,N_12962);
nor U13185 (N_13185,N_12851,N_12936);
or U13186 (N_13186,N_12615,N_12613);
nand U13187 (N_13187,N_12521,N_12602);
nand U13188 (N_13188,N_12818,N_12937);
and U13189 (N_13189,N_12919,N_12570);
nand U13190 (N_13190,N_12812,N_12771);
and U13191 (N_13191,N_12504,N_12863);
or U13192 (N_13192,N_12788,N_12557);
and U13193 (N_13193,N_12806,N_12603);
nor U13194 (N_13194,N_12621,N_12604);
nand U13195 (N_13195,N_12644,N_12877);
xnor U13196 (N_13196,N_12882,N_12864);
nand U13197 (N_13197,N_12903,N_12655);
nand U13198 (N_13198,N_12600,N_12619);
nand U13199 (N_13199,N_12529,N_12662);
nand U13200 (N_13200,N_12868,N_12669);
or U13201 (N_13201,N_12860,N_12990);
or U13202 (N_13202,N_12614,N_12502);
or U13203 (N_13203,N_12639,N_12736);
xor U13204 (N_13204,N_12674,N_12533);
and U13205 (N_13205,N_12873,N_12522);
and U13206 (N_13206,N_12609,N_12666);
or U13207 (N_13207,N_12792,N_12636);
and U13208 (N_13208,N_12974,N_12787);
or U13209 (N_13209,N_12681,N_12994);
and U13210 (N_13210,N_12943,N_12605);
and U13211 (N_13211,N_12909,N_12768);
or U13212 (N_13212,N_12770,N_12520);
nand U13213 (N_13213,N_12507,N_12542);
nand U13214 (N_13214,N_12821,N_12627);
and U13215 (N_13215,N_12531,N_12503);
nor U13216 (N_13216,N_12692,N_12647);
nor U13217 (N_13217,N_12592,N_12552);
and U13218 (N_13218,N_12772,N_12505);
nand U13219 (N_13219,N_12910,N_12916);
and U13220 (N_13220,N_12611,N_12584);
and U13221 (N_13221,N_12629,N_12886);
or U13222 (N_13222,N_12582,N_12752);
and U13223 (N_13223,N_12695,N_12791);
xor U13224 (N_13224,N_12853,N_12970);
nand U13225 (N_13225,N_12530,N_12515);
or U13226 (N_13226,N_12610,N_12748);
and U13227 (N_13227,N_12670,N_12578);
nor U13228 (N_13228,N_12733,N_12996);
or U13229 (N_13229,N_12798,N_12623);
xor U13230 (N_13230,N_12689,N_12510);
nor U13231 (N_13231,N_12764,N_12988);
or U13232 (N_13232,N_12523,N_12872);
nand U13233 (N_13233,N_12564,N_12708);
or U13234 (N_13234,N_12927,N_12816);
nand U13235 (N_13235,N_12649,N_12942);
and U13236 (N_13236,N_12536,N_12934);
nand U13237 (N_13237,N_12850,N_12754);
and U13238 (N_13238,N_12677,N_12878);
and U13239 (N_13239,N_12711,N_12948);
or U13240 (N_13240,N_12801,N_12888);
nand U13241 (N_13241,N_12944,N_12902);
nand U13242 (N_13242,N_12854,N_12538);
nor U13243 (N_13243,N_12585,N_12809);
and U13244 (N_13244,N_12580,N_12905);
or U13245 (N_13245,N_12500,N_12514);
xor U13246 (N_13246,N_12827,N_12556);
xnor U13247 (N_13247,N_12867,N_12675);
and U13248 (N_13248,N_12758,N_12815);
or U13249 (N_13249,N_12782,N_12713);
and U13250 (N_13250,N_12919,N_12949);
nand U13251 (N_13251,N_12652,N_12586);
nand U13252 (N_13252,N_12741,N_12920);
and U13253 (N_13253,N_12587,N_12506);
nand U13254 (N_13254,N_12865,N_12787);
nand U13255 (N_13255,N_12622,N_12978);
nand U13256 (N_13256,N_12655,N_12976);
nand U13257 (N_13257,N_12602,N_12613);
nor U13258 (N_13258,N_12663,N_12724);
xor U13259 (N_13259,N_12699,N_12954);
or U13260 (N_13260,N_12860,N_12618);
xnor U13261 (N_13261,N_12613,N_12895);
xnor U13262 (N_13262,N_12933,N_12689);
or U13263 (N_13263,N_12837,N_12821);
nor U13264 (N_13264,N_12747,N_12566);
nor U13265 (N_13265,N_12744,N_12538);
and U13266 (N_13266,N_12621,N_12643);
nand U13267 (N_13267,N_12954,N_12659);
or U13268 (N_13268,N_12607,N_12644);
and U13269 (N_13269,N_12750,N_12552);
nor U13270 (N_13270,N_12583,N_12622);
and U13271 (N_13271,N_12508,N_12814);
nand U13272 (N_13272,N_12983,N_12822);
and U13273 (N_13273,N_12543,N_12729);
nand U13274 (N_13274,N_12761,N_12776);
nor U13275 (N_13275,N_12972,N_12943);
or U13276 (N_13276,N_12971,N_12843);
nor U13277 (N_13277,N_12848,N_12919);
nand U13278 (N_13278,N_12887,N_12641);
nor U13279 (N_13279,N_12561,N_12572);
and U13280 (N_13280,N_12922,N_12894);
and U13281 (N_13281,N_12683,N_12740);
nor U13282 (N_13282,N_12685,N_12730);
nand U13283 (N_13283,N_12874,N_12734);
and U13284 (N_13284,N_12512,N_12570);
xnor U13285 (N_13285,N_12774,N_12768);
and U13286 (N_13286,N_12899,N_12608);
nand U13287 (N_13287,N_12921,N_12870);
nand U13288 (N_13288,N_12575,N_12595);
or U13289 (N_13289,N_12971,N_12632);
nand U13290 (N_13290,N_12999,N_12679);
or U13291 (N_13291,N_12919,N_12619);
nand U13292 (N_13292,N_12967,N_12724);
nand U13293 (N_13293,N_12510,N_12860);
and U13294 (N_13294,N_12847,N_12839);
nor U13295 (N_13295,N_12873,N_12710);
nand U13296 (N_13296,N_12879,N_12730);
nor U13297 (N_13297,N_12786,N_12708);
and U13298 (N_13298,N_12972,N_12811);
nor U13299 (N_13299,N_12644,N_12672);
nand U13300 (N_13300,N_12633,N_12972);
and U13301 (N_13301,N_12901,N_12562);
xnor U13302 (N_13302,N_12952,N_12862);
nand U13303 (N_13303,N_12997,N_12900);
or U13304 (N_13304,N_12788,N_12732);
or U13305 (N_13305,N_12538,N_12615);
nor U13306 (N_13306,N_12682,N_12605);
nand U13307 (N_13307,N_12634,N_12966);
or U13308 (N_13308,N_12948,N_12990);
nor U13309 (N_13309,N_12621,N_12841);
and U13310 (N_13310,N_12885,N_12779);
or U13311 (N_13311,N_12820,N_12875);
and U13312 (N_13312,N_12733,N_12551);
and U13313 (N_13313,N_12688,N_12752);
nand U13314 (N_13314,N_12582,N_12564);
nor U13315 (N_13315,N_12664,N_12996);
nand U13316 (N_13316,N_12839,N_12857);
xor U13317 (N_13317,N_12790,N_12828);
or U13318 (N_13318,N_12843,N_12709);
or U13319 (N_13319,N_12568,N_12838);
nand U13320 (N_13320,N_12724,N_12996);
and U13321 (N_13321,N_12803,N_12534);
nand U13322 (N_13322,N_12763,N_12527);
xor U13323 (N_13323,N_12520,N_12645);
nor U13324 (N_13324,N_12806,N_12943);
or U13325 (N_13325,N_12962,N_12778);
or U13326 (N_13326,N_12649,N_12693);
or U13327 (N_13327,N_12508,N_12746);
nand U13328 (N_13328,N_12814,N_12668);
xnor U13329 (N_13329,N_12776,N_12962);
xor U13330 (N_13330,N_12966,N_12810);
nor U13331 (N_13331,N_12861,N_12588);
xor U13332 (N_13332,N_12833,N_12703);
or U13333 (N_13333,N_12674,N_12828);
and U13334 (N_13334,N_12521,N_12553);
nor U13335 (N_13335,N_12962,N_12756);
nand U13336 (N_13336,N_12973,N_12866);
and U13337 (N_13337,N_12906,N_12631);
xnor U13338 (N_13338,N_12943,N_12881);
and U13339 (N_13339,N_12815,N_12595);
and U13340 (N_13340,N_12711,N_12869);
or U13341 (N_13341,N_12881,N_12728);
nor U13342 (N_13342,N_12569,N_12579);
and U13343 (N_13343,N_12701,N_12608);
or U13344 (N_13344,N_12633,N_12843);
nand U13345 (N_13345,N_12599,N_12713);
nor U13346 (N_13346,N_12909,N_12918);
nor U13347 (N_13347,N_12748,N_12938);
nand U13348 (N_13348,N_12965,N_12627);
or U13349 (N_13349,N_12887,N_12665);
or U13350 (N_13350,N_12846,N_12518);
or U13351 (N_13351,N_12674,N_12635);
nor U13352 (N_13352,N_12905,N_12903);
nor U13353 (N_13353,N_12999,N_12883);
nand U13354 (N_13354,N_12869,N_12756);
nor U13355 (N_13355,N_12540,N_12675);
nor U13356 (N_13356,N_12598,N_12803);
nor U13357 (N_13357,N_12745,N_12944);
nor U13358 (N_13358,N_12968,N_12779);
nand U13359 (N_13359,N_12866,N_12594);
or U13360 (N_13360,N_12777,N_12614);
and U13361 (N_13361,N_12569,N_12650);
nand U13362 (N_13362,N_12647,N_12576);
nand U13363 (N_13363,N_12746,N_12896);
or U13364 (N_13364,N_12930,N_12513);
nand U13365 (N_13365,N_12819,N_12936);
nand U13366 (N_13366,N_12959,N_12714);
nor U13367 (N_13367,N_12541,N_12979);
xnor U13368 (N_13368,N_12696,N_12876);
nand U13369 (N_13369,N_12576,N_12859);
and U13370 (N_13370,N_12741,N_12730);
and U13371 (N_13371,N_12528,N_12943);
or U13372 (N_13372,N_12775,N_12587);
and U13373 (N_13373,N_12540,N_12981);
nor U13374 (N_13374,N_12970,N_12863);
and U13375 (N_13375,N_12622,N_12763);
nand U13376 (N_13376,N_12822,N_12655);
nor U13377 (N_13377,N_12953,N_12855);
nor U13378 (N_13378,N_12910,N_12965);
or U13379 (N_13379,N_12778,N_12521);
nor U13380 (N_13380,N_12894,N_12533);
nand U13381 (N_13381,N_12685,N_12999);
nor U13382 (N_13382,N_12881,N_12663);
nor U13383 (N_13383,N_12857,N_12583);
or U13384 (N_13384,N_12606,N_12889);
or U13385 (N_13385,N_12814,N_12682);
xnor U13386 (N_13386,N_12814,N_12531);
nor U13387 (N_13387,N_12738,N_12911);
nand U13388 (N_13388,N_12508,N_12815);
xnor U13389 (N_13389,N_12856,N_12898);
xor U13390 (N_13390,N_12999,N_12686);
nor U13391 (N_13391,N_12756,N_12992);
and U13392 (N_13392,N_12582,N_12901);
nand U13393 (N_13393,N_12799,N_12738);
or U13394 (N_13394,N_12788,N_12908);
nand U13395 (N_13395,N_12994,N_12784);
or U13396 (N_13396,N_12670,N_12825);
or U13397 (N_13397,N_12571,N_12628);
and U13398 (N_13398,N_12541,N_12592);
and U13399 (N_13399,N_12997,N_12963);
or U13400 (N_13400,N_12519,N_12979);
nor U13401 (N_13401,N_12744,N_12549);
nand U13402 (N_13402,N_12972,N_12857);
or U13403 (N_13403,N_12700,N_12539);
nand U13404 (N_13404,N_12935,N_12530);
and U13405 (N_13405,N_12683,N_12876);
nand U13406 (N_13406,N_12645,N_12705);
nor U13407 (N_13407,N_12942,N_12761);
or U13408 (N_13408,N_12838,N_12895);
nor U13409 (N_13409,N_12554,N_12897);
xnor U13410 (N_13410,N_12621,N_12542);
or U13411 (N_13411,N_12649,N_12786);
xnor U13412 (N_13412,N_12524,N_12744);
or U13413 (N_13413,N_12832,N_12920);
and U13414 (N_13414,N_12909,N_12941);
and U13415 (N_13415,N_12755,N_12865);
or U13416 (N_13416,N_12783,N_12813);
xnor U13417 (N_13417,N_12867,N_12816);
nor U13418 (N_13418,N_12741,N_12894);
nor U13419 (N_13419,N_12729,N_12583);
nor U13420 (N_13420,N_12781,N_12897);
and U13421 (N_13421,N_12617,N_12780);
or U13422 (N_13422,N_12568,N_12867);
nand U13423 (N_13423,N_12747,N_12576);
nor U13424 (N_13424,N_12709,N_12957);
or U13425 (N_13425,N_12888,N_12635);
or U13426 (N_13426,N_12634,N_12764);
or U13427 (N_13427,N_12819,N_12815);
and U13428 (N_13428,N_12870,N_12596);
nor U13429 (N_13429,N_12538,N_12735);
xor U13430 (N_13430,N_12598,N_12619);
xor U13431 (N_13431,N_12668,N_12849);
nor U13432 (N_13432,N_12766,N_12587);
or U13433 (N_13433,N_12932,N_12805);
or U13434 (N_13434,N_12621,N_12625);
and U13435 (N_13435,N_12602,N_12565);
nand U13436 (N_13436,N_12827,N_12692);
and U13437 (N_13437,N_12755,N_12653);
and U13438 (N_13438,N_12797,N_12674);
or U13439 (N_13439,N_12770,N_12754);
and U13440 (N_13440,N_12768,N_12996);
nor U13441 (N_13441,N_12501,N_12601);
xnor U13442 (N_13442,N_12951,N_12816);
nand U13443 (N_13443,N_12878,N_12669);
nor U13444 (N_13444,N_12978,N_12681);
or U13445 (N_13445,N_12846,N_12682);
nand U13446 (N_13446,N_12516,N_12964);
nor U13447 (N_13447,N_12630,N_12509);
or U13448 (N_13448,N_12997,N_12646);
nand U13449 (N_13449,N_12583,N_12681);
and U13450 (N_13450,N_12929,N_12831);
xor U13451 (N_13451,N_12913,N_12763);
or U13452 (N_13452,N_12796,N_12833);
and U13453 (N_13453,N_12836,N_12644);
xnor U13454 (N_13454,N_12585,N_12605);
and U13455 (N_13455,N_12889,N_12698);
nor U13456 (N_13456,N_12898,N_12508);
or U13457 (N_13457,N_12858,N_12521);
and U13458 (N_13458,N_12775,N_12847);
nor U13459 (N_13459,N_12655,N_12940);
and U13460 (N_13460,N_12538,N_12695);
or U13461 (N_13461,N_12993,N_12734);
nand U13462 (N_13462,N_12511,N_12558);
xnor U13463 (N_13463,N_12970,N_12809);
or U13464 (N_13464,N_12859,N_12946);
xor U13465 (N_13465,N_12843,N_12636);
or U13466 (N_13466,N_12694,N_12597);
and U13467 (N_13467,N_12740,N_12990);
nand U13468 (N_13468,N_12929,N_12623);
nor U13469 (N_13469,N_12967,N_12760);
nor U13470 (N_13470,N_12868,N_12856);
nand U13471 (N_13471,N_12598,N_12988);
nand U13472 (N_13472,N_12937,N_12545);
or U13473 (N_13473,N_12935,N_12980);
nand U13474 (N_13474,N_12782,N_12685);
or U13475 (N_13475,N_12744,N_12752);
and U13476 (N_13476,N_12712,N_12732);
nand U13477 (N_13477,N_12983,N_12566);
nand U13478 (N_13478,N_12819,N_12991);
or U13479 (N_13479,N_12862,N_12895);
xor U13480 (N_13480,N_12656,N_12785);
nand U13481 (N_13481,N_12526,N_12884);
or U13482 (N_13482,N_12635,N_12859);
and U13483 (N_13483,N_12559,N_12865);
or U13484 (N_13484,N_12514,N_12961);
xnor U13485 (N_13485,N_12532,N_12916);
or U13486 (N_13486,N_12736,N_12549);
and U13487 (N_13487,N_12592,N_12941);
or U13488 (N_13488,N_12938,N_12775);
or U13489 (N_13489,N_12898,N_12906);
nand U13490 (N_13490,N_12674,N_12715);
nor U13491 (N_13491,N_12555,N_12749);
or U13492 (N_13492,N_12991,N_12818);
or U13493 (N_13493,N_12601,N_12913);
or U13494 (N_13494,N_12580,N_12624);
xnor U13495 (N_13495,N_12807,N_12802);
and U13496 (N_13496,N_12580,N_12665);
nor U13497 (N_13497,N_12966,N_12805);
or U13498 (N_13498,N_12831,N_12565);
nor U13499 (N_13499,N_12896,N_12933);
or U13500 (N_13500,N_13320,N_13136);
or U13501 (N_13501,N_13310,N_13301);
xnor U13502 (N_13502,N_13210,N_13333);
nor U13503 (N_13503,N_13189,N_13040);
or U13504 (N_13504,N_13049,N_13240);
nor U13505 (N_13505,N_13271,N_13363);
nand U13506 (N_13506,N_13013,N_13241);
and U13507 (N_13507,N_13071,N_13024);
nand U13508 (N_13508,N_13453,N_13327);
xnor U13509 (N_13509,N_13304,N_13267);
nor U13510 (N_13510,N_13439,N_13361);
or U13511 (N_13511,N_13467,N_13403);
nand U13512 (N_13512,N_13044,N_13186);
xor U13513 (N_13513,N_13391,N_13041);
or U13514 (N_13514,N_13141,N_13209);
nand U13515 (N_13515,N_13171,N_13113);
or U13516 (N_13516,N_13314,N_13352);
or U13517 (N_13517,N_13160,N_13207);
and U13518 (N_13518,N_13367,N_13079);
and U13519 (N_13519,N_13112,N_13462);
nor U13520 (N_13520,N_13461,N_13018);
xor U13521 (N_13521,N_13337,N_13346);
and U13522 (N_13522,N_13266,N_13148);
or U13523 (N_13523,N_13120,N_13316);
and U13524 (N_13524,N_13022,N_13108);
and U13525 (N_13525,N_13036,N_13286);
or U13526 (N_13526,N_13475,N_13483);
or U13527 (N_13527,N_13368,N_13094);
or U13528 (N_13528,N_13381,N_13030);
and U13529 (N_13529,N_13255,N_13176);
and U13530 (N_13530,N_13116,N_13274);
and U13531 (N_13531,N_13139,N_13470);
and U13532 (N_13532,N_13052,N_13338);
nor U13533 (N_13533,N_13334,N_13124);
nor U13534 (N_13534,N_13308,N_13447);
nor U13535 (N_13535,N_13350,N_13109);
and U13536 (N_13536,N_13300,N_13206);
and U13537 (N_13537,N_13469,N_13114);
xnor U13538 (N_13538,N_13277,N_13054);
or U13539 (N_13539,N_13218,N_13174);
xor U13540 (N_13540,N_13395,N_13070);
or U13541 (N_13541,N_13004,N_13482);
and U13542 (N_13542,N_13331,N_13242);
xnor U13543 (N_13543,N_13134,N_13042);
and U13544 (N_13544,N_13053,N_13353);
and U13545 (N_13545,N_13480,N_13477);
or U13546 (N_13546,N_13418,N_13384);
nand U13547 (N_13547,N_13390,N_13043);
or U13548 (N_13548,N_13153,N_13227);
or U13549 (N_13549,N_13493,N_13322);
nand U13550 (N_13550,N_13211,N_13010);
nand U13551 (N_13551,N_13130,N_13085);
and U13552 (N_13552,N_13027,N_13101);
or U13553 (N_13553,N_13223,N_13358);
nand U13554 (N_13554,N_13437,N_13489);
nand U13555 (N_13555,N_13293,N_13057);
nor U13556 (N_13556,N_13061,N_13473);
xor U13557 (N_13557,N_13247,N_13138);
xor U13558 (N_13558,N_13398,N_13156);
or U13559 (N_13559,N_13422,N_13129);
xor U13560 (N_13560,N_13236,N_13448);
or U13561 (N_13561,N_13232,N_13200);
nor U13562 (N_13562,N_13180,N_13386);
xor U13563 (N_13563,N_13014,N_13115);
nand U13564 (N_13564,N_13295,N_13029);
nor U13565 (N_13565,N_13238,N_13283);
and U13566 (N_13566,N_13122,N_13377);
and U13567 (N_13567,N_13137,N_13262);
xnor U13568 (N_13568,N_13032,N_13360);
nand U13569 (N_13569,N_13144,N_13430);
xor U13570 (N_13570,N_13149,N_13111);
and U13571 (N_13571,N_13161,N_13201);
nor U13572 (N_13572,N_13259,N_13075);
xnor U13573 (N_13573,N_13167,N_13311);
and U13574 (N_13574,N_13035,N_13163);
or U13575 (N_13575,N_13154,N_13172);
nor U13576 (N_13576,N_13399,N_13400);
and U13577 (N_13577,N_13455,N_13369);
nand U13578 (N_13578,N_13324,N_13117);
nand U13579 (N_13579,N_13008,N_13038);
or U13580 (N_13580,N_13226,N_13062);
nor U13581 (N_13581,N_13012,N_13260);
and U13582 (N_13582,N_13328,N_13364);
or U13583 (N_13583,N_13047,N_13323);
nand U13584 (N_13584,N_13088,N_13292);
nor U13585 (N_13585,N_13181,N_13383);
and U13586 (N_13586,N_13050,N_13276);
nand U13587 (N_13587,N_13091,N_13365);
nor U13588 (N_13588,N_13246,N_13284);
nor U13589 (N_13589,N_13248,N_13429);
nand U13590 (N_13590,N_13414,N_13318);
or U13591 (N_13591,N_13471,N_13147);
and U13592 (N_13592,N_13285,N_13005);
and U13593 (N_13593,N_13374,N_13288);
and U13594 (N_13594,N_13179,N_13451);
xor U13595 (N_13595,N_13261,N_13023);
nand U13596 (N_13596,N_13060,N_13359);
nand U13597 (N_13597,N_13188,N_13495);
nor U13598 (N_13598,N_13028,N_13362);
and U13599 (N_13599,N_13278,N_13376);
and U13600 (N_13600,N_13289,N_13019);
or U13601 (N_13601,N_13491,N_13356);
nor U13602 (N_13602,N_13195,N_13099);
nor U13603 (N_13603,N_13048,N_13474);
and U13604 (N_13604,N_13411,N_13404);
nand U13605 (N_13605,N_13347,N_13162);
and U13606 (N_13606,N_13125,N_13494);
xnor U13607 (N_13607,N_13457,N_13002);
nand U13608 (N_13608,N_13279,N_13104);
xnor U13609 (N_13609,N_13196,N_13131);
and U13610 (N_13610,N_13045,N_13214);
or U13611 (N_13611,N_13031,N_13164);
and U13612 (N_13612,N_13083,N_13184);
or U13613 (N_13613,N_13069,N_13388);
nand U13614 (N_13614,N_13230,N_13066);
and U13615 (N_13615,N_13287,N_13326);
or U13616 (N_13616,N_13419,N_13312);
or U13617 (N_13617,N_13450,N_13348);
nor U13618 (N_13618,N_13212,N_13126);
or U13619 (N_13619,N_13275,N_13090);
and U13620 (N_13620,N_13098,N_13349);
xnor U13621 (N_13621,N_13265,N_13250);
or U13622 (N_13622,N_13434,N_13413);
xnor U13623 (N_13623,N_13145,N_13199);
or U13624 (N_13624,N_13344,N_13064);
nor U13625 (N_13625,N_13194,N_13315);
or U13626 (N_13626,N_13135,N_13401);
nor U13627 (N_13627,N_13441,N_13373);
nor U13628 (N_13628,N_13225,N_13281);
nor U13629 (N_13629,N_13375,N_13105);
nor U13630 (N_13630,N_13177,N_13272);
nor U13631 (N_13631,N_13192,N_13086);
nor U13632 (N_13632,N_13492,N_13110);
and U13633 (N_13633,N_13183,N_13170);
or U13634 (N_13634,N_13397,N_13372);
or U13635 (N_13635,N_13335,N_13249);
nand U13636 (N_13636,N_13329,N_13423);
nor U13637 (N_13637,N_13202,N_13121);
or U13638 (N_13638,N_13321,N_13151);
and U13639 (N_13639,N_13478,N_13243);
and U13640 (N_13640,N_13128,N_13325);
nand U13641 (N_13641,N_13444,N_13468);
nand U13642 (N_13642,N_13392,N_13234);
nor U13643 (N_13643,N_13082,N_13290);
nand U13644 (N_13644,N_13092,N_13056);
nor U13645 (N_13645,N_13305,N_13472);
nor U13646 (N_13646,N_13296,N_13175);
nor U13647 (N_13647,N_13393,N_13496);
xor U13648 (N_13648,N_13096,N_13222);
and U13649 (N_13649,N_13166,N_13100);
nor U13650 (N_13650,N_13197,N_13178);
nor U13651 (N_13651,N_13340,N_13157);
nand U13652 (N_13652,N_13432,N_13428);
and U13653 (N_13653,N_13476,N_13132);
nor U13654 (N_13654,N_13436,N_13059);
nand U13655 (N_13655,N_13417,N_13006);
or U13656 (N_13656,N_13396,N_13254);
nor U13657 (N_13657,N_13264,N_13332);
nand U13658 (N_13658,N_13158,N_13354);
nand U13659 (N_13659,N_13063,N_13465);
nor U13660 (N_13660,N_13466,N_13270);
or U13661 (N_13661,N_13421,N_13402);
or U13662 (N_13662,N_13306,N_13382);
and U13663 (N_13663,N_13345,N_13205);
nand U13664 (N_13664,N_13268,N_13068);
nand U13665 (N_13665,N_13009,N_13415);
xor U13666 (N_13666,N_13198,N_13309);
and U13667 (N_13667,N_13445,N_13011);
nor U13668 (N_13668,N_13438,N_13389);
nand U13669 (N_13669,N_13118,N_13370);
xnor U13670 (N_13670,N_13224,N_13142);
nand U13671 (N_13671,N_13371,N_13067);
nand U13672 (N_13672,N_13235,N_13256);
nor U13673 (N_13673,N_13420,N_13017);
nor U13674 (N_13674,N_13280,N_13425);
nor U13675 (N_13675,N_13037,N_13107);
nor U13676 (N_13676,N_13302,N_13237);
and U13677 (N_13677,N_13097,N_13217);
and U13678 (N_13678,N_13407,N_13229);
nor U13679 (N_13679,N_13410,N_13341);
and U13680 (N_13680,N_13409,N_13074);
and U13681 (N_13681,N_13203,N_13233);
or U13682 (N_13682,N_13193,N_13251);
xnor U13683 (N_13683,N_13095,N_13155);
and U13684 (N_13684,N_13351,N_13498);
nor U13685 (N_13685,N_13394,N_13025);
nor U13686 (N_13686,N_13343,N_13051);
or U13687 (N_13687,N_13077,N_13463);
nor U13688 (N_13688,N_13454,N_13431);
nor U13689 (N_13689,N_13385,N_13424);
nand U13690 (N_13690,N_13258,N_13412);
nand U13691 (N_13691,N_13357,N_13231);
or U13692 (N_13692,N_13106,N_13426);
nand U13693 (N_13693,N_13015,N_13252);
nor U13694 (N_13694,N_13299,N_13072);
nor U13695 (N_13695,N_13143,N_13140);
xnor U13696 (N_13696,N_13152,N_13076);
xor U13697 (N_13697,N_13055,N_13486);
nor U13698 (N_13698,N_13003,N_13294);
nor U13699 (N_13699,N_13215,N_13001);
and U13700 (N_13700,N_13446,N_13435);
nand U13701 (N_13701,N_13220,N_13216);
or U13702 (N_13702,N_13490,N_13168);
and U13703 (N_13703,N_13452,N_13078);
nor U13704 (N_13704,N_13464,N_13330);
xor U13705 (N_13705,N_13460,N_13016);
or U13706 (N_13706,N_13073,N_13146);
nor U13707 (N_13707,N_13481,N_13065);
xnor U13708 (N_13708,N_13440,N_13458);
and U13709 (N_13709,N_13133,N_13339);
nor U13710 (N_13710,N_13000,N_13405);
or U13711 (N_13711,N_13119,N_13366);
and U13712 (N_13712,N_13123,N_13007);
nand U13713 (N_13713,N_13303,N_13080);
or U13714 (N_13714,N_13456,N_13185);
nand U13715 (N_13715,N_13307,N_13182);
and U13716 (N_13716,N_13433,N_13187);
xor U13717 (N_13717,N_13169,N_13026);
xnor U13718 (N_13718,N_13034,N_13087);
or U13719 (N_13719,N_13449,N_13102);
xnor U13720 (N_13720,N_13282,N_13208);
and U13721 (N_13721,N_13190,N_13263);
and U13722 (N_13722,N_13273,N_13297);
or U13723 (N_13723,N_13253,N_13342);
nor U13724 (N_13724,N_13081,N_13103);
nor U13725 (N_13725,N_13150,N_13479);
nor U13726 (N_13726,N_13380,N_13269);
nor U13727 (N_13727,N_13443,N_13173);
nand U13728 (N_13728,N_13485,N_13089);
nand U13729 (N_13729,N_13387,N_13406);
xor U13730 (N_13730,N_13488,N_13416);
nand U13731 (N_13731,N_13499,N_13459);
nor U13732 (N_13732,N_13442,N_13221);
or U13733 (N_13733,N_13039,N_13228);
nor U13734 (N_13734,N_13165,N_13191);
xnor U13735 (N_13735,N_13020,N_13487);
or U13736 (N_13736,N_13245,N_13058);
or U13737 (N_13737,N_13127,N_13257);
xor U13738 (N_13738,N_13244,N_13291);
xnor U13739 (N_13739,N_13159,N_13046);
nand U13740 (N_13740,N_13084,N_13298);
and U13741 (N_13741,N_13497,N_13239);
nor U13742 (N_13742,N_13219,N_13378);
nor U13743 (N_13743,N_13408,N_13427);
nor U13744 (N_13744,N_13313,N_13319);
nand U13745 (N_13745,N_13379,N_13213);
or U13746 (N_13746,N_13093,N_13355);
and U13747 (N_13747,N_13033,N_13021);
nor U13748 (N_13748,N_13336,N_13317);
and U13749 (N_13749,N_13484,N_13204);
xnor U13750 (N_13750,N_13459,N_13054);
nor U13751 (N_13751,N_13260,N_13179);
nor U13752 (N_13752,N_13404,N_13430);
xnor U13753 (N_13753,N_13344,N_13289);
or U13754 (N_13754,N_13277,N_13431);
nor U13755 (N_13755,N_13409,N_13365);
and U13756 (N_13756,N_13425,N_13470);
or U13757 (N_13757,N_13070,N_13029);
xor U13758 (N_13758,N_13446,N_13101);
xor U13759 (N_13759,N_13261,N_13063);
or U13760 (N_13760,N_13156,N_13289);
and U13761 (N_13761,N_13206,N_13069);
nor U13762 (N_13762,N_13446,N_13434);
or U13763 (N_13763,N_13135,N_13093);
nor U13764 (N_13764,N_13307,N_13388);
or U13765 (N_13765,N_13248,N_13071);
nand U13766 (N_13766,N_13248,N_13153);
xnor U13767 (N_13767,N_13380,N_13015);
nor U13768 (N_13768,N_13447,N_13166);
nor U13769 (N_13769,N_13034,N_13208);
nand U13770 (N_13770,N_13353,N_13202);
or U13771 (N_13771,N_13308,N_13218);
nor U13772 (N_13772,N_13076,N_13494);
and U13773 (N_13773,N_13380,N_13045);
nor U13774 (N_13774,N_13397,N_13203);
or U13775 (N_13775,N_13412,N_13462);
and U13776 (N_13776,N_13180,N_13327);
nand U13777 (N_13777,N_13319,N_13392);
or U13778 (N_13778,N_13043,N_13360);
or U13779 (N_13779,N_13344,N_13477);
nand U13780 (N_13780,N_13327,N_13391);
or U13781 (N_13781,N_13467,N_13187);
or U13782 (N_13782,N_13380,N_13460);
nand U13783 (N_13783,N_13361,N_13016);
xnor U13784 (N_13784,N_13443,N_13490);
nand U13785 (N_13785,N_13480,N_13169);
nor U13786 (N_13786,N_13243,N_13409);
nand U13787 (N_13787,N_13352,N_13377);
or U13788 (N_13788,N_13035,N_13264);
xor U13789 (N_13789,N_13434,N_13204);
and U13790 (N_13790,N_13043,N_13465);
and U13791 (N_13791,N_13072,N_13122);
and U13792 (N_13792,N_13070,N_13257);
xnor U13793 (N_13793,N_13133,N_13370);
or U13794 (N_13794,N_13368,N_13462);
nand U13795 (N_13795,N_13176,N_13368);
nand U13796 (N_13796,N_13271,N_13047);
and U13797 (N_13797,N_13367,N_13301);
nand U13798 (N_13798,N_13314,N_13042);
or U13799 (N_13799,N_13204,N_13228);
and U13800 (N_13800,N_13413,N_13009);
nor U13801 (N_13801,N_13484,N_13288);
or U13802 (N_13802,N_13016,N_13424);
nor U13803 (N_13803,N_13473,N_13285);
nor U13804 (N_13804,N_13475,N_13485);
and U13805 (N_13805,N_13344,N_13459);
or U13806 (N_13806,N_13146,N_13496);
and U13807 (N_13807,N_13349,N_13387);
xnor U13808 (N_13808,N_13162,N_13069);
nor U13809 (N_13809,N_13188,N_13010);
or U13810 (N_13810,N_13468,N_13466);
or U13811 (N_13811,N_13360,N_13057);
xor U13812 (N_13812,N_13037,N_13427);
nor U13813 (N_13813,N_13296,N_13438);
nor U13814 (N_13814,N_13278,N_13313);
nand U13815 (N_13815,N_13331,N_13139);
or U13816 (N_13816,N_13497,N_13362);
and U13817 (N_13817,N_13262,N_13249);
or U13818 (N_13818,N_13210,N_13404);
or U13819 (N_13819,N_13429,N_13367);
or U13820 (N_13820,N_13109,N_13171);
or U13821 (N_13821,N_13252,N_13075);
nand U13822 (N_13822,N_13128,N_13039);
xor U13823 (N_13823,N_13352,N_13310);
or U13824 (N_13824,N_13437,N_13292);
nor U13825 (N_13825,N_13455,N_13054);
nand U13826 (N_13826,N_13241,N_13073);
and U13827 (N_13827,N_13250,N_13447);
nand U13828 (N_13828,N_13467,N_13138);
nand U13829 (N_13829,N_13034,N_13197);
or U13830 (N_13830,N_13109,N_13222);
or U13831 (N_13831,N_13431,N_13026);
nand U13832 (N_13832,N_13324,N_13098);
xor U13833 (N_13833,N_13122,N_13457);
nor U13834 (N_13834,N_13466,N_13318);
and U13835 (N_13835,N_13427,N_13039);
nand U13836 (N_13836,N_13306,N_13224);
and U13837 (N_13837,N_13107,N_13067);
and U13838 (N_13838,N_13174,N_13371);
nor U13839 (N_13839,N_13211,N_13351);
and U13840 (N_13840,N_13368,N_13097);
and U13841 (N_13841,N_13391,N_13383);
and U13842 (N_13842,N_13409,N_13334);
nand U13843 (N_13843,N_13452,N_13432);
nor U13844 (N_13844,N_13121,N_13337);
nand U13845 (N_13845,N_13060,N_13042);
nand U13846 (N_13846,N_13048,N_13084);
or U13847 (N_13847,N_13349,N_13388);
nand U13848 (N_13848,N_13048,N_13479);
nor U13849 (N_13849,N_13024,N_13205);
nand U13850 (N_13850,N_13416,N_13402);
and U13851 (N_13851,N_13103,N_13280);
xnor U13852 (N_13852,N_13107,N_13035);
or U13853 (N_13853,N_13131,N_13017);
nand U13854 (N_13854,N_13026,N_13313);
nor U13855 (N_13855,N_13167,N_13490);
or U13856 (N_13856,N_13104,N_13009);
and U13857 (N_13857,N_13324,N_13442);
nand U13858 (N_13858,N_13449,N_13385);
or U13859 (N_13859,N_13355,N_13441);
and U13860 (N_13860,N_13357,N_13207);
nand U13861 (N_13861,N_13380,N_13400);
or U13862 (N_13862,N_13495,N_13161);
nand U13863 (N_13863,N_13303,N_13480);
nor U13864 (N_13864,N_13163,N_13275);
or U13865 (N_13865,N_13003,N_13259);
or U13866 (N_13866,N_13270,N_13183);
nand U13867 (N_13867,N_13078,N_13067);
and U13868 (N_13868,N_13426,N_13354);
nor U13869 (N_13869,N_13276,N_13483);
or U13870 (N_13870,N_13128,N_13006);
and U13871 (N_13871,N_13489,N_13461);
or U13872 (N_13872,N_13021,N_13445);
or U13873 (N_13873,N_13043,N_13228);
and U13874 (N_13874,N_13047,N_13248);
nor U13875 (N_13875,N_13441,N_13345);
and U13876 (N_13876,N_13350,N_13193);
nor U13877 (N_13877,N_13151,N_13116);
nor U13878 (N_13878,N_13388,N_13247);
nor U13879 (N_13879,N_13076,N_13123);
or U13880 (N_13880,N_13455,N_13470);
or U13881 (N_13881,N_13463,N_13002);
nand U13882 (N_13882,N_13160,N_13141);
nor U13883 (N_13883,N_13156,N_13338);
and U13884 (N_13884,N_13077,N_13291);
or U13885 (N_13885,N_13315,N_13410);
nand U13886 (N_13886,N_13401,N_13337);
or U13887 (N_13887,N_13256,N_13461);
or U13888 (N_13888,N_13059,N_13049);
nor U13889 (N_13889,N_13022,N_13472);
nor U13890 (N_13890,N_13158,N_13308);
nor U13891 (N_13891,N_13331,N_13053);
nand U13892 (N_13892,N_13369,N_13340);
or U13893 (N_13893,N_13185,N_13204);
nor U13894 (N_13894,N_13116,N_13149);
nor U13895 (N_13895,N_13018,N_13278);
nand U13896 (N_13896,N_13259,N_13133);
and U13897 (N_13897,N_13091,N_13201);
or U13898 (N_13898,N_13213,N_13066);
or U13899 (N_13899,N_13392,N_13031);
nor U13900 (N_13900,N_13331,N_13175);
nand U13901 (N_13901,N_13249,N_13082);
or U13902 (N_13902,N_13249,N_13460);
or U13903 (N_13903,N_13061,N_13201);
nor U13904 (N_13904,N_13032,N_13123);
and U13905 (N_13905,N_13313,N_13092);
nand U13906 (N_13906,N_13412,N_13305);
or U13907 (N_13907,N_13234,N_13037);
or U13908 (N_13908,N_13230,N_13017);
nand U13909 (N_13909,N_13078,N_13100);
and U13910 (N_13910,N_13484,N_13393);
or U13911 (N_13911,N_13422,N_13317);
nor U13912 (N_13912,N_13108,N_13424);
nand U13913 (N_13913,N_13108,N_13204);
xnor U13914 (N_13914,N_13087,N_13159);
nand U13915 (N_13915,N_13374,N_13270);
nand U13916 (N_13916,N_13290,N_13090);
nor U13917 (N_13917,N_13010,N_13454);
and U13918 (N_13918,N_13377,N_13155);
nor U13919 (N_13919,N_13495,N_13430);
and U13920 (N_13920,N_13488,N_13083);
nand U13921 (N_13921,N_13296,N_13422);
and U13922 (N_13922,N_13041,N_13159);
nor U13923 (N_13923,N_13103,N_13267);
and U13924 (N_13924,N_13075,N_13418);
and U13925 (N_13925,N_13102,N_13412);
nor U13926 (N_13926,N_13351,N_13265);
nand U13927 (N_13927,N_13199,N_13109);
and U13928 (N_13928,N_13197,N_13419);
xnor U13929 (N_13929,N_13239,N_13446);
nor U13930 (N_13930,N_13496,N_13107);
and U13931 (N_13931,N_13410,N_13495);
nand U13932 (N_13932,N_13225,N_13476);
nand U13933 (N_13933,N_13427,N_13143);
and U13934 (N_13934,N_13495,N_13117);
nand U13935 (N_13935,N_13369,N_13439);
and U13936 (N_13936,N_13358,N_13004);
or U13937 (N_13937,N_13165,N_13012);
or U13938 (N_13938,N_13288,N_13345);
nand U13939 (N_13939,N_13456,N_13115);
nor U13940 (N_13940,N_13108,N_13417);
xnor U13941 (N_13941,N_13378,N_13431);
nand U13942 (N_13942,N_13219,N_13228);
or U13943 (N_13943,N_13260,N_13127);
nor U13944 (N_13944,N_13099,N_13276);
nor U13945 (N_13945,N_13233,N_13092);
nand U13946 (N_13946,N_13198,N_13155);
or U13947 (N_13947,N_13096,N_13178);
nand U13948 (N_13948,N_13114,N_13426);
or U13949 (N_13949,N_13228,N_13199);
xor U13950 (N_13950,N_13486,N_13129);
xnor U13951 (N_13951,N_13368,N_13146);
and U13952 (N_13952,N_13179,N_13482);
xnor U13953 (N_13953,N_13143,N_13030);
nand U13954 (N_13954,N_13473,N_13265);
nor U13955 (N_13955,N_13129,N_13380);
nand U13956 (N_13956,N_13251,N_13019);
nand U13957 (N_13957,N_13240,N_13401);
nand U13958 (N_13958,N_13173,N_13281);
nand U13959 (N_13959,N_13150,N_13072);
xnor U13960 (N_13960,N_13314,N_13010);
and U13961 (N_13961,N_13194,N_13496);
and U13962 (N_13962,N_13264,N_13376);
nand U13963 (N_13963,N_13373,N_13482);
and U13964 (N_13964,N_13483,N_13069);
or U13965 (N_13965,N_13382,N_13327);
nand U13966 (N_13966,N_13471,N_13463);
nor U13967 (N_13967,N_13391,N_13066);
nor U13968 (N_13968,N_13442,N_13288);
nand U13969 (N_13969,N_13041,N_13005);
nand U13970 (N_13970,N_13040,N_13375);
and U13971 (N_13971,N_13482,N_13386);
nand U13972 (N_13972,N_13452,N_13005);
or U13973 (N_13973,N_13005,N_13315);
nand U13974 (N_13974,N_13311,N_13220);
xor U13975 (N_13975,N_13256,N_13168);
or U13976 (N_13976,N_13145,N_13401);
nor U13977 (N_13977,N_13439,N_13263);
and U13978 (N_13978,N_13063,N_13116);
and U13979 (N_13979,N_13340,N_13153);
and U13980 (N_13980,N_13028,N_13250);
or U13981 (N_13981,N_13004,N_13041);
xnor U13982 (N_13982,N_13368,N_13216);
and U13983 (N_13983,N_13012,N_13413);
or U13984 (N_13984,N_13056,N_13390);
nand U13985 (N_13985,N_13432,N_13402);
nand U13986 (N_13986,N_13447,N_13356);
and U13987 (N_13987,N_13346,N_13013);
nor U13988 (N_13988,N_13213,N_13149);
nand U13989 (N_13989,N_13189,N_13231);
or U13990 (N_13990,N_13424,N_13357);
and U13991 (N_13991,N_13417,N_13335);
nand U13992 (N_13992,N_13322,N_13218);
and U13993 (N_13993,N_13310,N_13118);
nor U13994 (N_13994,N_13122,N_13155);
nor U13995 (N_13995,N_13233,N_13033);
nand U13996 (N_13996,N_13354,N_13417);
nor U13997 (N_13997,N_13374,N_13212);
and U13998 (N_13998,N_13426,N_13013);
nor U13999 (N_13999,N_13035,N_13386);
nand U14000 (N_14000,N_13931,N_13794);
or U14001 (N_14001,N_13973,N_13710);
or U14002 (N_14002,N_13533,N_13933);
nor U14003 (N_14003,N_13500,N_13965);
and U14004 (N_14004,N_13876,N_13513);
nand U14005 (N_14005,N_13668,N_13647);
and U14006 (N_14006,N_13755,N_13890);
and U14007 (N_14007,N_13634,N_13960);
and U14008 (N_14008,N_13840,N_13749);
or U14009 (N_14009,N_13773,N_13519);
nand U14010 (N_14010,N_13652,N_13686);
and U14011 (N_14011,N_13817,N_13692);
nor U14012 (N_14012,N_13587,N_13820);
or U14013 (N_14013,N_13545,N_13869);
or U14014 (N_14014,N_13664,N_13666);
and U14015 (N_14015,N_13530,N_13851);
nor U14016 (N_14016,N_13637,N_13827);
nand U14017 (N_14017,N_13517,N_13789);
and U14018 (N_14018,N_13752,N_13829);
or U14019 (N_14019,N_13910,N_13638);
nand U14020 (N_14020,N_13662,N_13640);
or U14021 (N_14021,N_13583,N_13909);
nand U14022 (N_14022,N_13774,N_13760);
xor U14023 (N_14023,N_13551,N_13783);
nor U14024 (N_14024,N_13724,N_13711);
or U14025 (N_14025,N_13705,N_13540);
nor U14026 (N_14026,N_13746,N_13858);
xnor U14027 (N_14027,N_13707,N_13725);
and U14028 (N_14028,N_13595,N_13957);
nor U14029 (N_14029,N_13942,N_13887);
and U14030 (N_14030,N_13850,N_13534);
nor U14031 (N_14031,N_13650,N_13733);
nand U14032 (N_14032,N_13782,N_13864);
or U14033 (N_14033,N_13722,N_13753);
nand U14034 (N_14034,N_13875,N_13883);
nand U14035 (N_14035,N_13572,N_13976);
nand U14036 (N_14036,N_13518,N_13983);
nand U14037 (N_14037,N_13510,N_13993);
and U14038 (N_14038,N_13508,N_13894);
and U14039 (N_14039,N_13970,N_13867);
or U14040 (N_14040,N_13826,N_13852);
or U14041 (N_14041,N_13588,N_13536);
nand U14042 (N_14042,N_13630,N_13712);
xor U14043 (N_14043,N_13527,N_13963);
nand U14044 (N_14044,N_13735,N_13905);
nand U14045 (N_14045,N_13861,N_13766);
or U14046 (N_14046,N_13882,N_13916);
and U14047 (N_14047,N_13521,N_13997);
nor U14048 (N_14048,N_13844,N_13667);
or U14049 (N_14049,N_13504,N_13609);
nor U14050 (N_14050,N_13619,N_13742);
nor U14051 (N_14051,N_13683,N_13635);
and U14052 (N_14052,N_13653,N_13512);
and U14053 (N_14053,N_13807,N_13915);
and U14054 (N_14054,N_13935,N_13843);
or U14055 (N_14055,N_13926,N_13924);
or U14056 (N_14056,N_13507,N_13694);
nand U14057 (N_14057,N_13586,N_13552);
and U14058 (N_14058,N_13661,N_13954);
nor U14059 (N_14059,N_13779,N_13633);
or U14060 (N_14060,N_13918,N_13862);
nor U14061 (N_14061,N_13900,N_13865);
nand U14062 (N_14062,N_13961,N_13772);
or U14063 (N_14063,N_13799,N_13870);
or U14064 (N_14064,N_13947,N_13855);
or U14065 (N_14065,N_13688,N_13987);
and U14066 (N_14066,N_13687,N_13901);
nor U14067 (N_14067,N_13522,N_13823);
or U14068 (N_14068,N_13571,N_13631);
nand U14069 (N_14069,N_13798,N_13800);
xor U14070 (N_14070,N_13599,N_13932);
xor U14071 (N_14071,N_13948,N_13695);
and U14072 (N_14072,N_13659,N_13984);
xor U14073 (N_14073,N_13863,N_13790);
nand U14074 (N_14074,N_13663,N_13685);
nand U14075 (N_14075,N_13832,N_13546);
nand U14076 (N_14076,N_13673,N_13816);
nand U14077 (N_14077,N_13645,N_13740);
nand U14078 (N_14078,N_13803,N_13505);
xnor U14079 (N_14079,N_13657,N_13582);
or U14080 (N_14080,N_13793,N_13729);
nand U14081 (N_14081,N_13718,N_13950);
nor U14082 (N_14082,N_13985,N_13743);
or U14083 (N_14083,N_13830,N_13660);
nor U14084 (N_14084,N_13547,N_13968);
and U14085 (N_14085,N_13515,N_13784);
nand U14086 (N_14086,N_13628,N_13568);
nor U14087 (N_14087,N_13770,N_13739);
nor U14088 (N_14088,N_13994,N_13592);
nor U14089 (N_14089,N_13842,N_13975);
nand U14090 (N_14090,N_13925,N_13560);
and U14091 (N_14091,N_13767,N_13538);
nor U14092 (N_14092,N_13971,N_13771);
nand U14093 (N_14093,N_13708,N_13516);
xnor U14094 (N_14094,N_13991,N_13777);
or U14095 (N_14095,N_13818,N_13612);
nand U14096 (N_14096,N_13921,N_13849);
and U14097 (N_14097,N_13643,N_13853);
nand U14098 (N_14098,N_13821,N_13556);
nand U14099 (N_14099,N_13693,N_13627);
or U14100 (N_14100,N_13966,N_13763);
nor U14101 (N_14101,N_13626,N_13780);
nand U14102 (N_14102,N_13728,N_13574);
nand U14103 (N_14103,N_13614,N_13952);
nand U14104 (N_14104,N_13651,N_13559);
or U14105 (N_14105,N_13689,N_13723);
and U14106 (N_14106,N_13956,N_13549);
nand U14107 (N_14107,N_13969,N_13613);
and U14108 (N_14108,N_13810,N_13778);
or U14109 (N_14109,N_13600,N_13715);
xnor U14110 (N_14110,N_13928,N_13745);
and U14111 (N_14111,N_13874,N_13822);
nand U14112 (N_14112,N_13691,N_13995);
nand U14113 (N_14113,N_13791,N_13848);
and U14114 (N_14114,N_13980,N_13529);
and U14115 (N_14115,N_13902,N_13854);
nand U14116 (N_14116,N_13509,N_13616);
and U14117 (N_14117,N_13597,N_13929);
and U14118 (N_14118,N_13611,N_13544);
and U14119 (N_14119,N_13681,N_13709);
xor U14120 (N_14120,N_13701,N_13736);
nor U14121 (N_14121,N_13744,N_13716);
nand U14122 (N_14122,N_13881,N_13506);
nor U14123 (N_14123,N_13603,N_13888);
nor U14124 (N_14124,N_13917,N_13636);
nand U14125 (N_14125,N_13781,N_13678);
nor U14126 (N_14126,N_13868,N_13676);
nor U14127 (N_14127,N_13554,N_13700);
or U14128 (N_14128,N_13589,N_13886);
or U14129 (N_14129,N_13892,N_13819);
nand U14130 (N_14130,N_13895,N_13584);
and U14131 (N_14131,N_13562,N_13656);
or U14132 (N_14132,N_13941,N_13804);
nor U14133 (N_14133,N_13542,N_13992);
nand U14134 (N_14134,N_13897,N_13805);
xor U14135 (N_14135,N_13986,N_13857);
nand U14136 (N_14136,N_13684,N_13788);
nand U14137 (N_14137,N_13675,N_13919);
or U14138 (N_14138,N_13741,N_13576);
and U14139 (N_14139,N_13776,N_13824);
or U14140 (N_14140,N_13768,N_13537);
and U14141 (N_14141,N_13503,N_13605);
and U14142 (N_14142,N_13525,N_13769);
and U14143 (N_14143,N_13696,N_13937);
or U14144 (N_14144,N_13904,N_13761);
and U14145 (N_14145,N_13811,N_13541);
nand U14146 (N_14146,N_13837,N_13623);
or U14147 (N_14147,N_13775,N_13801);
nor U14148 (N_14148,N_13615,N_13880);
or U14149 (N_14149,N_13978,N_13955);
nor U14150 (N_14150,N_13720,N_13502);
or U14151 (N_14151,N_13702,N_13945);
nand U14152 (N_14152,N_13879,N_13951);
nor U14153 (N_14153,N_13873,N_13658);
xnor U14154 (N_14154,N_13682,N_13737);
nor U14155 (N_14155,N_13714,N_13814);
nand U14156 (N_14156,N_13543,N_13856);
nand U14157 (N_14157,N_13558,N_13936);
or U14158 (N_14158,N_13699,N_13580);
nor U14159 (N_14159,N_13677,N_13938);
nor U14160 (N_14160,N_13912,N_13996);
nand U14161 (N_14161,N_13859,N_13730);
xor U14162 (N_14162,N_13646,N_13578);
or U14163 (N_14163,N_13573,N_13514);
or U14164 (N_14164,N_13569,N_13838);
or U14165 (N_14165,N_13898,N_13629);
nand U14166 (N_14166,N_13564,N_13557);
or U14167 (N_14167,N_13958,N_13553);
and U14168 (N_14168,N_13555,N_13672);
nor U14169 (N_14169,N_13639,N_13617);
and U14170 (N_14170,N_13786,N_13934);
nand U14171 (N_14171,N_13914,N_13885);
and U14172 (N_14172,N_13758,N_13899);
and U14173 (N_14173,N_13964,N_13998);
and U14174 (N_14174,N_13757,N_13602);
nor U14175 (N_14175,N_13579,N_13581);
or U14176 (N_14176,N_13526,N_13908);
nor U14177 (N_14177,N_13641,N_13893);
or U14178 (N_14178,N_13759,N_13999);
nor U14179 (N_14179,N_13665,N_13841);
or U14180 (N_14180,N_13732,N_13979);
and U14181 (N_14181,N_13812,N_13765);
nand U14182 (N_14182,N_13601,N_13949);
nor U14183 (N_14183,N_13642,N_13797);
nand U14184 (N_14184,N_13566,N_13726);
nand U14185 (N_14185,N_13836,N_13911);
or U14186 (N_14186,N_13698,N_13717);
xor U14187 (N_14187,N_13815,N_13520);
nand U14188 (N_14188,N_13977,N_13561);
nand U14189 (N_14189,N_13649,N_13532);
nor U14190 (N_14190,N_13577,N_13679);
nor U14191 (N_14191,N_13713,N_13787);
and U14192 (N_14192,N_13940,N_13825);
or U14193 (N_14193,N_13974,N_13808);
or U14194 (N_14194,N_13621,N_13671);
xor U14195 (N_14195,N_13511,N_13860);
nand U14196 (N_14196,N_13528,N_13754);
and U14197 (N_14197,N_13721,N_13884);
xnor U14198 (N_14198,N_13622,N_13891);
nand U14199 (N_14199,N_13930,N_13834);
nor U14200 (N_14200,N_13872,N_13644);
nand U14201 (N_14201,N_13943,N_13719);
xnor U14202 (N_14202,N_13704,N_13847);
xnor U14203 (N_14203,N_13795,N_13731);
nand U14204 (N_14204,N_13697,N_13846);
and U14205 (N_14205,N_13967,N_13990);
xnor U14206 (N_14206,N_13594,N_13590);
nor U14207 (N_14207,N_13906,N_13738);
xnor U14208 (N_14208,N_13624,N_13703);
nor U14209 (N_14209,N_13922,N_13748);
and U14210 (N_14210,N_13889,N_13607);
or U14211 (N_14211,N_13655,N_13806);
nand U14212 (N_14212,N_13654,N_13591);
nand U14213 (N_14213,N_13962,N_13751);
or U14214 (N_14214,N_13845,N_13871);
or U14215 (N_14215,N_13690,N_13792);
or U14216 (N_14216,N_13896,N_13648);
xnor U14217 (N_14217,N_13523,N_13944);
or U14218 (N_14218,N_13680,N_13608);
or U14219 (N_14219,N_13501,N_13946);
nand U14220 (N_14220,N_13548,N_13669);
nand U14221 (N_14221,N_13839,N_13972);
nor U14222 (N_14222,N_13734,N_13620);
nor U14223 (N_14223,N_13563,N_13550);
or U14224 (N_14224,N_13670,N_13632);
nor U14225 (N_14225,N_13706,N_13593);
xor U14226 (N_14226,N_13596,N_13567);
xor U14227 (N_14227,N_13939,N_13878);
and U14228 (N_14228,N_13828,N_13920);
nor U14229 (N_14229,N_13598,N_13927);
or U14230 (N_14230,N_13796,N_13565);
xor U14231 (N_14231,N_13535,N_13604);
or U14232 (N_14232,N_13524,N_13913);
and U14233 (N_14233,N_13585,N_13866);
nor U14234 (N_14234,N_13903,N_13809);
nor U14235 (N_14235,N_13674,N_13764);
or U14236 (N_14236,N_13923,N_13575);
or U14237 (N_14237,N_13833,N_13750);
and U14238 (N_14238,N_13606,N_13813);
and U14239 (N_14239,N_13531,N_13907);
or U14240 (N_14240,N_13570,N_13539);
or U14241 (N_14241,N_13981,N_13877);
or U14242 (N_14242,N_13610,N_13959);
and U14243 (N_14243,N_13727,N_13747);
or U14244 (N_14244,N_13618,N_13835);
nor U14245 (N_14245,N_13785,N_13756);
and U14246 (N_14246,N_13989,N_13802);
or U14247 (N_14247,N_13988,N_13831);
nand U14248 (N_14248,N_13953,N_13625);
nor U14249 (N_14249,N_13982,N_13762);
nand U14250 (N_14250,N_13619,N_13500);
nor U14251 (N_14251,N_13881,N_13864);
nand U14252 (N_14252,N_13730,N_13776);
or U14253 (N_14253,N_13768,N_13821);
and U14254 (N_14254,N_13938,N_13838);
or U14255 (N_14255,N_13847,N_13729);
xor U14256 (N_14256,N_13730,N_13773);
and U14257 (N_14257,N_13816,N_13967);
nor U14258 (N_14258,N_13783,N_13876);
or U14259 (N_14259,N_13976,N_13784);
xnor U14260 (N_14260,N_13900,N_13988);
and U14261 (N_14261,N_13646,N_13506);
nand U14262 (N_14262,N_13503,N_13736);
or U14263 (N_14263,N_13637,N_13530);
or U14264 (N_14264,N_13927,N_13879);
or U14265 (N_14265,N_13560,N_13963);
or U14266 (N_14266,N_13859,N_13631);
nand U14267 (N_14267,N_13951,N_13634);
nor U14268 (N_14268,N_13549,N_13806);
nor U14269 (N_14269,N_13773,N_13842);
nor U14270 (N_14270,N_13877,N_13753);
nor U14271 (N_14271,N_13545,N_13863);
nor U14272 (N_14272,N_13885,N_13602);
or U14273 (N_14273,N_13554,N_13568);
nor U14274 (N_14274,N_13525,N_13676);
xor U14275 (N_14275,N_13704,N_13731);
nor U14276 (N_14276,N_13558,N_13513);
or U14277 (N_14277,N_13883,N_13610);
or U14278 (N_14278,N_13539,N_13943);
nand U14279 (N_14279,N_13740,N_13652);
and U14280 (N_14280,N_13505,N_13912);
nor U14281 (N_14281,N_13798,N_13899);
nor U14282 (N_14282,N_13916,N_13926);
or U14283 (N_14283,N_13692,N_13722);
nor U14284 (N_14284,N_13656,N_13778);
or U14285 (N_14285,N_13719,N_13507);
and U14286 (N_14286,N_13693,N_13827);
or U14287 (N_14287,N_13873,N_13918);
and U14288 (N_14288,N_13568,N_13930);
nor U14289 (N_14289,N_13727,N_13854);
and U14290 (N_14290,N_13689,N_13704);
and U14291 (N_14291,N_13678,N_13572);
nand U14292 (N_14292,N_13551,N_13793);
and U14293 (N_14293,N_13590,N_13869);
nand U14294 (N_14294,N_13932,N_13533);
nor U14295 (N_14295,N_13671,N_13781);
or U14296 (N_14296,N_13673,N_13729);
nand U14297 (N_14297,N_13909,N_13931);
nand U14298 (N_14298,N_13985,N_13505);
xor U14299 (N_14299,N_13591,N_13753);
nand U14300 (N_14300,N_13862,N_13896);
or U14301 (N_14301,N_13920,N_13538);
xnor U14302 (N_14302,N_13900,N_13711);
nor U14303 (N_14303,N_13795,N_13814);
or U14304 (N_14304,N_13806,N_13913);
or U14305 (N_14305,N_13987,N_13792);
and U14306 (N_14306,N_13939,N_13778);
nand U14307 (N_14307,N_13716,N_13639);
nor U14308 (N_14308,N_13758,N_13908);
and U14309 (N_14309,N_13830,N_13846);
and U14310 (N_14310,N_13999,N_13692);
nand U14311 (N_14311,N_13578,N_13807);
and U14312 (N_14312,N_13907,N_13634);
and U14313 (N_14313,N_13712,N_13838);
or U14314 (N_14314,N_13538,N_13705);
nor U14315 (N_14315,N_13872,N_13854);
nand U14316 (N_14316,N_13518,N_13918);
nand U14317 (N_14317,N_13806,N_13531);
nor U14318 (N_14318,N_13750,N_13756);
nand U14319 (N_14319,N_13761,N_13994);
nor U14320 (N_14320,N_13810,N_13572);
nand U14321 (N_14321,N_13832,N_13915);
nor U14322 (N_14322,N_13864,N_13802);
or U14323 (N_14323,N_13965,N_13971);
nor U14324 (N_14324,N_13531,N_13734);
or U14325 (N_14325,N_13919,N_13737);
xnor U14326 (N_14326,N_13751,N_13884);
or U14327 (N_14327,N_13909,N_13668);
and U14328 (N_14328,N_13936,N_13863);
nand U14329 (N_14329,N_13986,N_13771);
nor U14330 (N_14330,N_13826,N_13683);
and U14331 (N_14331,N_13707,N_13848);
nand U14332 (N_14332,N_13578,N_13702);
nand U14333 (N_14333,N_13539,N_13886);
nand U14334 (N_14334,N_13710,N_13848);
nor U14335 (N_14335,N_13802,N_13566);
nand U14336 (N_14336,N_13835,N_13827);
nand U14337 (N_14337,N_13876,N_13930);
nor U14338 (N_14338,N_13588,N_13725);
nor U14339 (N_14339,N_13644,N_13623);
or U14340 (N_14340,N_13595,N_13716);
and U14341 (N_14341,N_13878,N_13907);
nor U14342 (N_14342,N_13511,N_13754);
nor U14343 (N_14343,N_13798,N_13886);
nand U14344 (N_14344,N_13925,N_13532);
or U14345 (N_14345,N_13982,N_13708);
or U14346 (N_14346,N_13653,N_13555);
nor U14347 (N_14347,N_13757,N_13584);
nand U14348 (N_14348,N_13802,N_13875);
or U14349 (N_14349,N_13733,N_13988);
and U14350 (N_14350,N_13959,N_13571);
xnor U14351 (N_14351,N_13594,N_13944);
or U14352 (N_14352,N_13723,N_13899);
nand U14353 (N_14353,N_13819,N_13993);
and U14354 (N_14354,N_13568,N_13895);
or U14355 (N_14355,N_13875,N_13719);
nor U14356 (N_14356,N_13806,N_13520);
and U14357 (N_14357,N_13643,N_13736);
nand U14358 (N_14358,N_13718,N_13590);
nand U14359 (N_14359,N_13942,N_13973);
or U14360 (N_14360,N_13502,N_13741);
and U14361 (N_14361,N_13501,N_13882);
nand U14362 (N_14362,N_13696,N_13877);
or U14363 (N_14363,N_13617,N_13957);
and U14364 (N_14364,N_13818,N_13687);
nand U14365 (N_14365,N_13766,N_13691);
nor U14366 (N_14366,N_13782,N_13554);
nor U14367 (N_14367,N_13601,N_13657);
and U14368 (N_14368,N_13840,N_13887);
nor U14369 (N_14369,N_13634,N_13744);
and U14370 (N_14370,N_13985,N_13641);
or U14371 (N_14371,N_13629,N_13679);
nor U14372 (N_14372,N_13988,N_13630);
or U14373 (N_14373,N_13855,N_13739);
nand U14374 (N_14374,N_13995,N_13635);
nand U14375 (N_14375,N_13798,N_13858);
or U14376 (N_14376,N_13820,N_13501);
and U14377 (N_14377,N_13662,N_13602);
and U14378 (N_14378,N_13803,N_13935);
and U14379 (N_14379,N_13627,N_13650);
and U14380 (N_14380,N_13958,N_13674);
and U14381 (N_14381,N_13624,N_13737);
and U14382 (N_14382,N_13689,N_13584);
nand U14383 (N_14383,N_13610,N_13549);
nor U14384 (N_14384,N_13615,N_13870);
nand U14385 (N_14385,N_13988,N_13617);
and U14386 (N_14386,N_13541,N_13823);
nor U14387 (N_14387,N_13890,N_13625);
or U14388 (N_14388,N_13635,N_13797);
nor U14389 (N_14389,N_13529,N_13542);
nor U14390 (N_14390,N_13781,N_13909);
or U14391 (N_14391,N_13875,N_13676);
and U14392 (N_14392,N_13582,N_13989);
nand U14393 (N_14393,N_13968,N_13590);
and U14394 (N_14394,N_13923,N_13921);
or U14395 (N_14395,N_13734,N_13997);
nand U14396 (N_14396,N_13710,N_13912);
nand U14397 (N_14397,N_13934,N_13548);
nor U14398 (N_14398,N_13708,N_13625);
or U14399 (N_14399,N_13890,N_13940);
xor U14400 (N_14400,N_13729,N_13539);
nand U14401 (N_14401,N_13797,N_13925);
xnor U14402 (N_14402,N_13626,N_13817);
nand U14403 (N_14403,N_13818,N_13789);
and U14404 (N_14404,N_13617,N_13558);
xor U14405 (N_14405,N_13883,N_13595);
nor U14406 (N_14406,N_13748,N_13745);
or U14407 (N_14407,N_13821,N_13875);
and U14408 (N_14408,N_13963,N_13573);
xor U14409 (N_14409,N_13653,N_13926);
or U14410 (N_14410,N_13845,N_13866);
nor U14411 (N_14411,N_13821,N_13847);
or U14412 (N_14412,N_13687,N_13598);
nor U14413 (N_14413,N_13825,N_13674);
and U14414 (N_14414,N_13686,N_13789);
nor U14415 (N_14415,N_13809,N_13639);
nand U14416 (N_14416,N_13991,N_13787);
nor U14417 (N_14417,N_13709,N_13745);
nand U14418 (N_14418,N_13858,N_13525);
xnor U14419 (N_14419,N_13640,N_13716);
or U14420 (N_14420,N_13833,N_13652);
nand U14421 (N_14421,N_13989,N_13624);
nand U14422 (N_14422,N_13918,N_13813);
nor U14423 (N_14423,N_13947,N_13732);
xor U14424 (N_14424,N_13565,N_13515);
xor U14425 (N_14425,N_13930,N_13747);
nor U14426 (N_14426,N_13779,N_13964);
nand U14427 (N_14427,N_13723,N_13890);
nor U14428 (N_14428,N_13754,N_13519);
xor U14429 (N_14429,N_13951,N_13739);
nor U14430 (N_14430,N_13749,N_13917);
nor U14431 (N_14431,N_13815,N_13714);
or U14432 (N_14432,N_13921,N_13591);
or U14433 (N_14433,N_13645,N_13504);
nand U14434 (N_14434,N_13528,N_13640);
or U14435 (N_14435,N_13983,N_13809);
nand U14436 (N_14436,N_13584,N_13740);
xnor U14437 (N_14437,N_13952,N_13993);
xor U14438 (N_14438,N_13943,N_13609);
nor U14439 (N_14439,N_13618,N_13622);
nor U14440 (N_14440,N_13711,N_13748);
and U14441 (N_14441,N_13512,N_13665);
xnor U14442 (N_14442,N_13921,N_13754);
nor U14443 (N_14443,N_13590,N_13997);
and U14444 (N_14444,N_13947,N_13895);
or U14445 (N_14445,N_13512,N_13889);
nor U14446 (N_14446,N_13854,N_13641);
and U14447 (N_14447,N_13579,N_13853);
and U14448 (N_14448,N_13952,N_13752);
or U14449 (N_14449,N_13660,N_13954);
and U14450 (N_14450,N_13836,N_13929);
and U14451 (N_14451,N_13526,N_13683);
and U14452 (N_14452,N_13574,N_13998);
or U14453 (N_14453,N_13859,N_13773);
xor U14454 (N_14454,N_13643,N_13683);
and U14455 (N_14455,N_13695,N_13655);
nand U14456 (N_14456,N_13890,N_13689);
and U14457 (N_14457,N_13641,N_13612);
or U14458 (N_14458,N_13733,N_13686);
and U14459 (N_14459,N_13670,N_13785);
and U14460 (N_14460,N_13719,N_13850);
nand U14461 (N_14461,N_13728,N_13821);
nand U14462 (N_14462,N_13842,N_13554);
nand U14463 (N_14463,N_13745,N_13660);
nand U14464 (N_14464,N_13975,N_13991);
nand U14465 (N_14465,N_13625,N_13815);
nor U14466 (N_14466,N_13879,N_13522);
xor U14467 (N_14467,N_13776,N_13713);
nor U14468 (N_14468,N_13523,N_13560);
nor U14469 (N_14469,N_13840,N_13525);
and U14470 (N_14470,N_13877,N_13502);
nand U14471 (N_14471,N_13524,N_13945);
or U14472 (N_14472,N_13740,N_13833);
or U14473 (N_14473,N_13971,N_13519);
xnor U14474 (N_14474,N_13801,N_13618);
or U14475 (N_14475,N_13903,N_13578);
or U14476 (N_14476,N_13597,N_13524);
or U14477 (N_14477,N_13854,N_13670);
nand U14478 (N_14478,N_13703,N_13925);
or U14479 (N_14479,N_13524,N_13933);
and U14480 (N_14480,N_13771,N_13762);
xor U14481 (N_14481,N_13816,N_13971);
nand U14482 (N_14482,N_13672,N_13755);
nor U14483 (N_14483,N_13796,N_13568);
and U14484 (N_14484,N_13543,N_13510);
nand U14485 (N_14485,N_13582,N_13906);
nor U14486 (N_14486,N_13911,N_13740);
nor U14487 (N_14487,N_13681,N_13842);
nor U14488 (N_14488,N_13846,N_13927);
nor U14489 (N_14489,N_13626,N_13709);
and U14490 (N_14490,N_13512,N_13533);
nand U14491 (N_14491,N_13783,N_13994);
or U14492 (N_14492,N_13660,N_13506);
nand U14493 (N_14493,N_13733,N_13508);
and U14494 (N_14494,N_13654,N_13556);
and U14495 (N_14495,N_13748,N_13956);
nand U14496 (N_14496,N_13580,N_13895);
or U14497 (N_14497,N_13570,N_13835);
nor U14498 (N_14498,N_13594,N_13543);
and U14499 (N_14499,N_13732,N_13708);
or U14500 (N_14500,N_14058,N_14353);
and U14501 (N_14501,N_14439,N_14088);
xor U14502 (N_14502,N_14382,N_14355);
and U14503 (N_14503,N_14024,N_14329);
nor U14504 (N_14504,N_14295,N_14260);
and U14505 (N_14505,N_14230,N_14362);
nand U14506 (N_14506,N_14471,N_14487);
and U14507 (N_14507,N_14434,N_14397);
nand U14508 (N_14508,N_14181,N_14436);
nor U14509 (N_14509,N_14299,N_14091);
xor U14510 (N_14510,N_14310,N_14048);
and U14511 (N_14511,N_14277,N_14428);
or U14512 (N_14512,N_14405,N_14121);
or U14513 (N_14513,N_14486,N_14477);
nand U14514 (N_14514,N_14367,N_14194);
and U14515 (N_14515,N_14422,N_14031);
or U14516 (N_14516,N_14231,N_14391);
and U14517 (N_14517,N_14330,N_14418);
or U14518 (N_14518,N_14416,N_14301);
xor U14519 (N_14519,N_14219,N_14496);
xnor U14520 (N_14520,N_14077,N_14119);
or U14521 (N_14521,N_14370,N_14460);
nand U14522 (N_14522,N_14432,N_14014);
or U14523 (N_14523,N_14317,N_14415);
or U14524 (N_14524,N_14149,N_14017);
nand U14525 (N_14525,N_14475,N_14417);
nand U14526 (N_14526,N_14093,N_14390);
or U14527 (N_14527,N_14221,N_14141);
and U14528 (N_14528,N_14045,N_14130);
nand U14529 (N_14529,N_14041,N_14163);
or U14530 (N_14530,N_14307,N_14117);
and U14531 (N_14531,N_14189,N_14257);
nor U14532 (N_14532,N_14003,N_14440);
and U14533 (N_14533,N_14204,N_14213);
and U14534 (N_14534,N_14006,N_14429);
xor U14535 (N_14535,N_14351,N_14228);
nand U14536 (N_14536,N_14446,N_14407);
nor U14537 (N_14537,N_14150,N_14450);
or U14538 (N_14538,N_14452,N_14065);
and U14539 (N_14539,N_14354,N_14347);
or U14540 (N_14540,N_14158,N_14344);
or U14541 (N_14541,N_14293,N_14110);
or U14542 (N_14542,N_14424,N_14318);
nand U14543 (N_14543,N_14379,N_14180);
nand U14544 (N_14544,N_14001,N_14314);
nand U14545 (N_14545,N_14075,N_14346);
nor U14546 (N_14546,N_14366,N_14489);
nor U14547 (N_14547,N_14171,N_14061);
xnor U14548 (N_14548,N_14143,N_14021);
and U14549 (N_14549,N_14223,N_14082);
and U14550 (N_14550,N_14335,N_14485);
and U14551 (N_14551,N_14078,N_14085);
nand U14552 (N_14552,N_14385,N_14215);
or U14553 (N_14553,N_14388,N_14381);
nor U14554 (N_14554,N_14499,N_14339);
nor U14555 (N_14555,N_14345,N_14466);
nor U14556 (N_14556,N_14195,N_14461);
or U14557 (N_14557,N_14177,N_14144);
nand U14558 (N_14558,N_14247,N_14242);
nand U14559 (N_14559,N_14152,N_14164);
or U14560 (N_14560,N_14095,N_14297);
nand U14561 (N_14561,N_14320,N_14057);
or U14562 (N_14562,N_14043,N_14029);
and U14563 (N_14563,N_14280,N_14020);
nor U14564 (N_14564,N_14127,N_14465);
nand U14565 (N_14565,N_14456,N_14115);
nor U14566 (N_14566,N_14350,N_14387);
or U14567 (N_14567,N_14254,N_14483);
or U14568 (N_14568,N_14401,N_14481);
or U14569 (N_14569,N_14212,N_14291);
nor U14570 (N_14570,N_14176,N_14265);
nand U14571 (N_14571,N_14101,N_14013);
nor U14572 (N_14572,N_14409,N_14298);
and U14573 (N_14573,N_14214,N_14140);
nor U14574 (N_14574,N_14285,N_14156);
nor U14575 (N_14575,N_14010,N_14454);
nor U14576 (N_14576,N_14455,N_14028);
nor U14577 (N_14577,N_14411,N_14125);
or U14578 (N_14578,N_14178,N_14210);
nand U14579 (N_14579,N_14060,N_14136);
xnor U14580 (N_14580,N_14448,N_14102);
nor U14581 (N_14581,N_14472,N_14296);
nand U14582 (N_14582,N_14403,N_14441);
nor U14583 (N_14583,N_14224,N_14090);
nor U14584 (N_14584,N_14071,N_14087);
nand U14585 (N_14585,N_14217,N_14201);
xnor U14586 (N_14586,N_14476,N_14209);
xnor U14587 (N_14587,N_14404,N_14459);
or U14588 (N_14588,N_14315,N_14137);
or U14589 (N_14589,N_14341,N_14161);
or U14590 (N_14590,N_14442,N_14395);
or U14591 (N_14591,N_14258,N_14283);
or U14592 (N_14592,N_14474,N_14490);
nor U14593 (N_14593,N_14286,N_14433);
nor U14594 (N_14594,N_14099,N_14222);
nor U14595 (N_14595,N_14106,N_14316);
nor U14596 (N_14596,N_14263,N_14063);
nor U14597 (N_14597,N_14270,N_14072);
nor U14598 (N_14598,N_14308,N_14216);
and U14599 (N_14599,N_14092,N_14208);
and U14600 (N_14600,N_14179,N_14288);
or U14601 (N_14601,N_14337,N_14049);
or U14602 (N_14602,N_14128,N_14174);
nor U14603 (N_14603,N_14444,N_14312);
nand U14604 (N_14604,N_14463,N_14226);
or U14605 (N_14605,N_14034,N_14253);
nor U14606 (N_14606,N_14100,N_14131);
or U14607 (N_14607,N_14113,N_14153);
nand U14608 (N_14608,N_14083,N_14042);
nand U14609 (N_14609,N_14064,N_14426);
xor U14610 (N_14610,N_14035,N_14000);
xnor U14611 (N_14611,N_14185,N_14166);
nand U14612 (N_14612,N_14427,N_14134);
nand U14613 (N_14613,N_14326,N_14451);
nand U14614 (N_14614,N_14290,N_14030);
nand U14615 (N_14615,N_14281,N_14142);
xnor U14616 (N_14616,N_14340,N_14044);
and U14617 (N_14617,N_14259,N_14437);
and U14618 (N_14618,N_14008,N_14386);
nor U14619 (N_14619,N_14357,N_14373);
or U14620 (N_14620,N_14334,N_14464);
or U14621 (N_14621,N_14383,N_14004);
nand U14622 (N_14622,N_14068,N_14300);
xnor U14623 (N_14623,N_14467,N_14108);
nor U14624 (N_14624,N_14053,N_14396);
nand U14625 (N_14625,N_14282,N_14272);
or U14626 (N_14626,N_14193,N_14038);
nand U14627 (N_14627,N_14022,N_14192);
or U14628 (N_14628,N_14393,N_14399);
or U14629 (N_14629,N_14449,N_14267);
or U14630 (N_14630,N_14132,N_14073);
nand U14631 (N_14631,N_14146,N_14089);
or U14632 (N_14632,N_14358,N_14438);
nor U14633 (N_14633,N_14250,N_14096);
nand U14634 (N_14634,N_14016,N_14245);
nor U14635 (N_14635,N_14323,N_14112);
nor U14636 (N_14636,N_14243,N_14311);
and U14637 (N_14637,N_14155,N_14187);
and U14638 (N_14638,N_14331,N_14468);
or U14639 (N_14639,N_14470,N_14107);
nor U14640 (N_14640,N_14074,N_14384);
nand U14641 (N_14641,N_14333,N_14015);
nand U14642 (N_14642,N_14248,N_14199);
or U14643 (N_14643,N_14328,N_14233);
nor U14644 (N_14644,N_14040,N_14162);
nor U14645 (N_14645,N_14484,N_14081);
and U14646 (N_14646,N_14462,N_14175);
and U14647 (N_14647,N_14046,N_14332);
xor U14648 (N_14648,N_14037,N_14349);
and U14649 (N_14649,N_14183,N_14343);
xor U14650 (N_14650,N_14148,N_14080);
nand U14651 (N_14651,N_14197,N_14431);
and U14652 (N_14652,N_14241,N_14012);
nor U14653 (N_14653,N_14145,N_14327);
or U14654 (N_14654,N_14457,N_14309);
nor U14655 (N_14655,N_14264,N_14443);
nand U14656 (N_14656,N_14190,N_14413);
nor U14657 (N_14657,N_14207,N_14066);
xnor U14658 (N_14658,N_14124,N_14206);
nand U14659 (N_14659,N_14419,N_14203);
and U14660 (N_14660,N_14005,N_14394);
or U14661 (N_14661,N_14410,N_14261);
nand U14662 (N_14662,N_14104,N_14139);
nor U14663 (N_14663,N_14160,N_14120);
or U14664 (N_14664,N_14033,N_14458);
or U14665 (N_14665,N_14109,N_14118);
xnor U14666 (N_14666,N_14122,N_14453);
and U14667 (N_14667,N_14002,N_14262);
nor U14668 (N_14668,N_14036,N_14322);
nand U14669 (N_14669,N_14009,N_14211);
nor U14670 (N_14670,N_14154,N_14196);
or U14671 (N_14671,N_14406,N_14062);
and U14672 (N_14672,N_14389,N_14011);
nand U14673 (N_14673,N_14306,N_14268);
or U14674 (N_14674,N_14239,N_14055);
nor U14675 (N_14675,N_14186,N_14236);
and U14676 (N_14676,N_14114,N_14287);
xor U14677 (N_14677,N_14244,N_14069);
or U14678 (N_14678,N_14498,N_14420);
xor U14679 (N_14679,N_14234,N_14138);
xnor U14680 (N_14680,N_14338,N_14374);
nor U14681 (N_14681,N_14421,N_14188);
nand U14682 (N_14682,N_14380,N_14492);
nor U14683 (N_14683,N_14086,N_14319);
nor U14684 (N_14684,N_14050,N_14056);
and U14685 (N_14685,N_14051,N_14054);
and U14686 (N_14686,N_14325,N_14359);
or U14687 (N_14687,N_14478,N_14479);
nor U14688 (N_14688,N_14047,N_14473);
nand U14689 (N_14689,N_14278,N_14157);
nand U14690 (N_14690,N_14365,N_14169);
nor U14691 (N_14691,N_14273,N_14289);
and U14692 (N_14692,N_14147,N_14067);
or U14693 (N_14693,N_14336,N_14123);
or U14694 (N_14694,N_14237,N_14172);
xor U14695 (N_14695,N_14302,N_14133);
nand U14696 (N_14696,N_14356,N_14469);
xnor U14697 (N_14697,N_14084,N_14402);
nor U14698 (N_14698,N_14304,N_14274);
or U14699 (N_14699,N_14220,N_14294);
nand U14700 (N_14700,N_14198,N_14129);
or U14701 (N_14701,N_14229,N_14023);
nand U14702 (N_14702,N_14491,N_14361);
nor U14703 (N_14703,N_14488,N_14376);
nor U14704 (N_14704,N_14255,N_14052);
nand U14705 (N_14705,N_14249,N_14240);
or U14706 (N_14706,N_14400,N_14360);
nor U14707 (N_14707,N_14430,N_14369);
nor U14708 (N_14708,N_14225,N_14218);
nand U14709 (N_14709,N_14105,N_14159);
or U14710 (N_14710,N_14173,N_14039);
nand U14711 (N_14711,N_14227,N_14266);
or U14712 (N_14712,N_14246,N_14126);
xor U14713 (N_14713,N_14342,N_14377);
nor U14714 (N_14714,N_14284,N_14375);
and U14715 (N_14715,N_14303,N_14372);
nand U14716 (N_14716,N_14425,N_14238);
or U14717 (N_14717,N_14276,N_14079);
nor U14718 (N_14718,N_14324,N_14497);
xor U14719 (N_14719,N_14447,N_14167);
or U14720 (N_14720,N_14363,N_14251);
nand U14721 (N_14721,N_14191,N_14007);
xor U14722 (N_14722,N_14200,N_14103);
or U14723 (N_14723,N_14482,N_14392);
nand U14724 (N_14724,N_14025,N_14271);
and U14725 (N_14725,N_14256,N_14116);
and U14726 (N_14726,N_14279,N_14070);
nand U14727 (N_14727,N_14445,N_14292);
and U14728 (N_14728,N_14494,N_14412);
nand U14729 (N_14729,N_14423,N_14027);
nand U14730 (N_14730,N_14165,N_14076);
nand U14731 (N_14731,N_14059,N_14252);
nand U14732 (N_14732,N_14098,N_14182);
or U14733 (N_14733,N_14032,N_14371);
nor U14734 (N_14734,N_14348,N_14019);
nand U14735 (N_14735,N_14364,N_14097);
nand U14736 (N_14736,N_14184,N_14151);
and U14737 (N_14737,N_14368,N_14094);
and U14738 (N_14738,N_14480,N_14269);
xnor U14739 (N_14739,N_14495,N_14493);
or U14740 (N_14740,N_14135,N_14232);
and U14741 (N_14741,N_14414,N_14168);
nand U14742 (N_14742,N_14235,N_14170);
and U14743 (N_14743,N_14408,N_14313);
nand U14744 (N_14744,N_14202,N_14205);
xor U14745 (N_14745,N_14111,N_14435);
or U14746 (N_14746,N_14305,N_14378);
nand U14747 (N_14747,N_14398,N_14026);
xnor U14748 (N_14748,N_14275,N_14018);
or U14749 (N_14749,N_14352,N_14321);
nand U14750 (N_14750,N_14464,N_14057);
and U14751 (N_14751,N_14414,N_14112);
or U14752 (N_14752,N_14247,N_14457);
nor U14753 (N_14753,N_14159,N_14252);
nor U14754 (N_14754,N_14020,N_14497);
or U14755 (N_14755,N_14171,N_14385);
or U14756 (N_14756,N_14466,N_14373);
nor U14757 (N_14757,N_14114,N_14007);
nand U14758 (N_14758,N_14058,N_14350);
nand U14759 (N_14759,N_14479,N_14084);
or U14760 (N_14760,N_14130,N_14316);
xnor U14761 (N_14761,N_14261,N_14136);
nor U14762 (N_14762,N_14171,N_14324);
and U14763 (N_14763,N_14329,N_14421);
or U14764 (N_14764,N_14200,N_14129);
and U14765 (N_14765,N_14042,N_14011);
xor U14766 (N_14766,N_14304,N_14365);
nor U14767 (N_14767,N_14300,N_14122);
or U14768 (N_14768,N_14339,N_14065);
nand U14769 (N_14769,N_14393,N_14309);
nor U14770 (N_14770,N_14083,N_14011);
or U14771 (N_14771,N_14136,N_14399);
and U14772 (N_14772,N_14116,N_14119);
nand U14773 (N_14773,N_14243,N_14310);
nand U14774 (N_14774,N_14295,N_14052);
nor U14775 (N_14775,N_14344,N_14435);
and U14776 (N_14776,N_14143,N_14264);
nor U14777 (N_14777,N_14269,N_14048);
nand U14778 (N_14778,N_14421,N_14005);
nor U14779 (N_14779,N_14236,N_14318);
xor U14780 (N_14780,N_14026,N_14422);
nand U14781 (N_14781,N_14381,N_14208);
nand U14782 (N_14782,N_14211,N_14453);
or U14783 (N_14783,N_14419,N_14136);
and U14784 (N_14784,N_14189,N_14285);
xor U14785 (N_14785,N_14122,N_14455);
or U14786 (N_14786,N_14350,N_14137);
xor U14787 (N_14787,N_14134,N_14442);
or U14788 (N_14788,N_14270,N_14318);
nand U14789 (N_14789,N_14458,N_14148);
xor U14790 (N_14790,N_14152,N_14461);
nand U14791 (N_14791,N_14168,N_14445);
nand U14792 (N_14792,N_14071,N_14425);
nor U14793 (N_14793,N_14193,N_14328);
nand U14794 (N_14794,N_14225,N_14216);
nor U14795 (N_14795,N_14081,N_14487);
and U14796 (N_14796,N_14119,N_14304);
or U14797 (N_14797,N_14435,N_14058);
or U14798 (N_14798,N_14361,N_14146);
xnor U14799 (N_14799,N_14001,N_14250);
nand U14800 (N_14800,N_14186,N_14281);
or U14801 (N_14801,N_14349,N_14498);
or U14802 (N_14802,N_14066,N_14123);
nor U14803 (N_14803,N_14415,N_14142);
and U14804 (N_14804,N_14474,N_14361);
nand U14805 (N_14805,N_14403,N_14260);
and U14806 (N_14806,N_14283,N_14132);
or U14807 (N_14807,N_14230,N_14140);
and U14808 (N_14808,N_14486,N_14276);
nand U14809 (N_14809,N_14344,N_14267);
and U14810 (N_14810,N_14062,N_14440);
nand U14811 (N_14811,N_14429,N_14027);
xnor U14812 (N_14812,N_14037,N_14088);
and U14813 (N_14813,N_14372,N_14154);
and U14814 (N_14814,N_14327,N_14334);
nor U14815 (N_14815,N_14216,N_14392);
or U14816 (N_14816,N_14360,N_14066);
nor U14817 (N_14817,N_14142,N_14258);
or U14818 (N_14818,N_14464,N_14459);
xnor U14819 (N_14819,N_14023,N_14176);
and U14820 (N_14820,N_14127,N_14112);
nand U14821 (N_14821,N_14435,N_14458);
xor U14822 (N_14822,N_14224,N_14485);
xor U14823 (N_14823,N_14349,N_14445);
xor U14824 (N_14824,N_14031,N_14213);
nand U14825 (N_14825,N_14247,N_14192);
and U14826 (N_14826,N_14035,N_14113);
and U14827 (N_14827,N_14378,N_14304);
and U14828 (N_14828,N_14025,N_14330);
and U14829 (N_14829,N_14013,N_14154);
nor U14830 (N_14830,N_14356,N_14489);
nand U14831 (N_14831,N_14282,N_14415);
and U14832 (N_14832,N_14328,N_14042);
nor U14833 (N_14833,N_14237,N_14431);
and U14834 (N_14834,N_14213,N_14371);
or U14835 (N_14835,N_14162,N_14322);
or U14836 (N_14836,N_14456,N_14102);
nor U14837 (N_14837,N_14257,N_14185);
nor U14838 (N_14838,N_14296,N_14245);
and U14839 (N_14839,N_14463,N_14347);
or U14840 (N_14840,N_14375,N_14430);
nand U14841 (N_14841,N_14280,N_14037);
nor U14842 (N_14842,N_14477,N_14119);
or U14843 (N_14843,N_14432,N_14322);
nand U14844 (N_14844,N_14387,N_14111);
and U14845 (N_14845,N_14331,N_14377);
nor U14846 (N_14846,N_14346,N_14419);
or U14847 (N_14847,N_14209,N_14147);
and U14848 (N_14848,N_14133,N_14267);
or U14849 (N_14849,N_14173,N_14130);
and U14850 (N_14850,N_14117,N_14212);
nor U14851 (N_14851,N_14487,N_14233);
nor U14852 (N_14852,N_14224,N_14051);
xor U14853 (N_14853,N_14263,N_14288);
and U14854 (N_14854,N_14434,N_14350);
nand U14855 (N_14855,N_14046,N_14040);
or U14856 (N_14856,N_14148,N_14012);
nand U14857 (N_14857,N_14449,N_14448);
nor U14858 (N_14858,N_14147,N_14334);
and U14859 (N_14859,N_14274,N_14039);
nand U14860 (N_14860,N_14071,N_14070);
nor U14861 (N_14861,N_14425,N_14138);
or U14862 (N_14862,N_14428,N_14298);
nor U14863 (N_14863,N_14443,N_14143);
or U14864 (N_14864,N_14059,N_14020);
and U14865 (N_14865,N_14419,N_14314);
xnor U14866 (N_14866,N_14306,N_14025);
or U14867 (N_14867,N_14493,N_14205);
or U14868 (N_14868,N_14002,N_14361);
nand U14869 (N_14869,N_14339,N_14125);
nor U14870 (N_14870,N_14413,N_14007);
xor U14871 (N_14871,N_14079,N_14476);
nand U14872 (N_14872,N_14215,N_14287);
or U14873 (N_14873,N_14484,N_14430);
nand U14874 (N_14874,N_14176,N_14444);
nor U14875 (N_14875,N_14124,N_14078);
and U14876 (N_14876,N_14077,N_14198);
nor U14877 (N_14877,N_14289,N_14105);
and U14878 (N_14878,N_14186,N_14453);
or U14879 (N_14879,N_14066,N_14471);
nand U14880 (N_14880,N_14214,N_14350);
xnor U14881 (N_14881,N_14421,N_14291);
or U14882 (N_14882,N_14240,N_14416);
and U14883 (N_14883,N_14123,N_14483);
or U14884 (N_14884,N_14197,N_14412);
or U14885 (N_14885,N_14180,N_14053);
nand U14886 (N_14886,N_14073,N_14154);
and U14887 (N_14887,N_14192,N_14154);
nor U14888 (N_14888,N_14050,N_14209);
nor U14889 (N_14889,N_14218,N_14347);
nand U14890 (N_14890,N_14259,N_14066);
xnor U14891 (N_14891,N_14201,N_14121);
and U14892 (N_14892,N_14007,N_14002);
nor U14893 (N_14893,N_14016,N_14425);
or U14894 (N_14894,N_14420,N_14233);
or U14895 (N_14895,N_14454,N_14422);
and U14896 (N_14896,N_14214,N_14161);
and U14897 (N_14897,N_14077,N_14011);
xor U14898 (N_14898,N_14411,N_14262);
or U14899 (N_14899,N_14080,N_14414);
nand U14900 (N_14900,N_14305,N_14358);
and U14901 (N_14901,N_14455,N_14214);
and U14902 (N_14902,N_14198,N_14147);
nand U14903 (N_14903,N_14060,N_14476);
nor U14904 (N_14904,N_14097,N_14050);
xnor U14905 (N_14905,N_14344,N_14277);
nor U14906 (N_14906,N_14048,N_14282);
nand U14907 (N_14907,N_14324,N_14081);
nor U14908 (N_14908,N_14473,N_14418);
xnor U14909 (N_14909,N_14431,N_14182);
and U14910 (N_14910,N_14084,N_14092);
or U14911 (N_14911,N_14098,N_14092);
nor U14912 (N_14912,N_14492,N_14165);
and U14913 (N_14913,N_14307,N_14100);
nand U14914 (N_14914,N_14411,N_14297);
nand U14915 (N_14915,N_14439,N_14221);
xor U14916 (N_14916,N_14263,N_14485);
nor U14917 (N_14917,N_14231,N_14374);
and U14918 (N_14918,N_14122,N_14429);
and U14919 (N_14919,N_14380,N_14034);
or U14920 (N_14920,N_14334,N_14196);
xor U14921 (N_14921,N_14262,N_14080);
nand U14922 (N_14922,N_14274,N_14313);
nor U14923 (N_14923,N_14446,N_14005);
nor U14924 (N_14924,N_14351,N_14245);
nand U14925 (N_14925,N_14493,N_14374);
nor U14926 (N_14926,N_14009,N_14432);
or U14927 (N_14927,N_14407,N_14209);
nand U14928 (N_14928,N_14057,N_14195);
or U14929 (N_14929,N_14008,N_14116);
or U14930 (N_14930,N_14419,N_14044);
nand U14931 (N_14931,N_14037,N_14176);
or U14932 (N_14932,N_14284,N_14061);
xnor U14933 (N_14933,N_14072,N_14491);
xor U14934 (N_14934,N_14385,N_14487);
and U14935 (N_14935,N_14338,N_14261);
or U14936 (N_14936,N_14256,N_14481);
nor U14937 (N_14937,N_14318,N_14438);
and U14938 (N_14938,N_14388,N_14476);
or U14939 (N_14939,N_14496,N_14308);
or U14940 (N_14940,N_14460,N_14108);
xnor U14941 (N_14941,N_14389,N_14316);
and U14942 (N_14942,N_14108,N_14218);
nand U14943 (N_14943,N_14393,N_14352);
and U14944 (N_14944,N_14139,N_14260);
and U14945 (N_14945,N_14239,N_14118);
xnor U14946 (N_14946,N_14445,N_14096);
and U14947 (N_14947,N_14103,N_14474);
or U14948 (N_14948,N_14326,N_14019);
or U14949 (N_14949,N_14389,N_14449);
or U14950 (N_14950,N_14457,N_14216);
and U14951 (N_14951,N_14332,N_14377);
nand U14952 (N_14952,N_14205,N_14244);
or U14953 (N_14953,N_14078,N_14297);
nand U14954 (N_14954,N_14351,N_14445);
or U14955 (N_14955,N_14425,N_14291);
and U14956 (N_14956,N_14300,N_14041);
nand U14957 (N_14957,N_14273,N_14252);
and U14958 (N_14958,N_14348,N_14308);
xor U14959 (N_14959,N_14123,N_14392);
or U14960 (N_14960,N_14353,N_14068);
nand U14961 (N_14961,N_14266,N_14455);
xor U14962 (N_14962,N_14103,N_14296);
or U14963 (N_14963,N_14460,N_14126);
nor U14964 (N_14964,N_14496,N_14258);
and U14965 (N_14965,N_14465,N_14053);
nand U14966 (N_14966,N_14306,N_14145);
nor U14967 (N_14967,N_14271,N_14209);
or U14968 (N_14968,N_14007,N_14131);
nand U14969 (N_14969,N_14225,N_14425);
nand U14970 (N_14970,N_14160,N_14068);
or U14971 (N_14971,N_14408,N_14084);
nand U14972 (N_14972,N_14158,N_14428);
and U14973 (N_14973,N_14256,N_14002);
and U14974 (N_14974,N_14012,N_14231);
xor U14975 (N_14975,N_14092,N_14172);
nor U14976 (N_14976,N_14009,N_14460);
and U14977 (N_14977,N_14336,N_14389);
xnor U14978 (N_14978,N_14057,N_14467);
or U14979 (N_14979,N_14105,N_14176);
nand U14980 (N_14980,N_14349,N_14267);
or U14981 (N_14981,N_14058,N_14129);
or U14982 (N_14982,N_14192,N_14472);
nand U14983 (N_14983,N_14340,N_14307);
and U14984 (N_14984,N_14213,N_14321);
nor U14985 (N_14985,N_14469,N_14179);
nand U14986 (N_14986,N_14097,N_14184);
and U14987 (N_14987,N_14397,N_14459);
nor U14988 (N_14988,N_14111,N_14127);
and U14989 (N_14989,N_14456,N_14169);
and U14990 (N_14990,N_14032,N_14496);
and U14991 (N_14991,N_14093,N_14431);
nor U14992 (N_14992,N_14028,N_14295);
xnor U14993 (N_14993,N_14354,N_14269);
and U14994 (N_14994,N_14026,N_14403);
or U14995 (N_14995,N_14045,N_14018);
nand U14996 (N_14996,N_14212,N_14414);
nand U14997 (N_14997,N_14002,N_14079);
nand U14998 (N_14998,N_14400,N_14016);
and U14999 (N_14999,N_14468,N_14312);
nand U15000 (N_15000,N_14606,N_14716);
nor U15001 (N_15001,N_14643,N_14763);
or U15002 (N_15002,N_14565,N_14732);
or U15003 (N_15003,N_14779,N_14795);
nor U15004 (N_15004,N_14739,N_14512);
nor U15005 (N_15005,N_14642,N_14540);
nand U15006 (N_15006,N_14586,N_14638);
nor U15007 (N_15007,N_14912,N_14721);
nand U15008 (N_15008,N_14743,N_14740);
nand U15009 (N_15009,N_14841,N_14979);
nor U15010 (N_15010,N_14943,N_14682);
and U15011 (N_15011,N_14817,N_14977);
nand U15012 (N_15012,N_14530,N_14972);
nand U15013 (N_15013,N_14574,N_14834);
nor U15014 (N_15014,N_14759,N_14526);
and U15015 (N_15015,N_14703,N_14805);
xor U15016 (N_15016,N_14927,N_14899);
xor U15017 (N_15017,N_14630,N_14553);
nor U15018 (N_15018,N_14714,N_14903);
nand U15019 (N_15019,N_14864,N_14515);
nor U15020 (N_15020,N_14902,N_14810);
nand U15021 (N_15021,N_14722,N_14564);
nor U15022 (N_15022,N_14889,N_14860);
and U15023 (N_15023,N_14713,N_14788);
or U15024 (N_15024,N_14980,N_14873);
or U15025 (N_15025,N_14723,N_14745);
nor U15026 (N_15026,N_14556,N_14915);
and U15027 (N_15027,N_14949,N_14663);
or U15028 (N_15028,N_14659,N_14560);
and U15029 (N_15029,N_14568,N_14958);
nor U15030 (N_15030,N_14547,N_14942);
nand U15031 (N_15031,N_14991,N_14803);
or U15032 (N_15032,N_14572,N_14602);
nand U15033 (N_15033,N_14896,N_14617);
nor U15034 (N_15034,N_14907,N_14531);
or U15035 (N_15035,N_14822,N_14744);
and U15036 (N_15036,N_14888,N_14988);
or U15037 (N_15037,N_14761,N_14625);
or U15038 (N_15038,N_14809,N_14830);
xor U15039 (N_15039,N_14708,N_14725);
and U15040 (N_15040,N_14550,N_14711);
nor U15041 (N_15041,N_14557,N_14571);
nand U15042 (N_15042,N_14598,N_14673);
and U15043 (N_15043,N_14612,N_14506);
or U15044 (N_15044,N_14882,N_14777);
or U15045 (N_15045,N_14534,N_14885);
and U15046 (N_15046,N_14683,N_14909);
and U15047 (N_15047,N_14866,N_14825);
and U15048 (N_15048,N_14906,N_14733);
nor U15049 (N_15049,N_14842,N_14691);
and U15050 (N_15050,N_14575,N_14939);
nor U15051 (N_15051,N_14604,N_14601);
nand U15052 (N_15052,N_14814,N_14762);
or U15053 (N_15053,N_14868,N_14946);
nor U15054 (N_15054,N_14964,N_14827);
and U15055 (N_15055,N_14687,N_14752);
nand U15056 (N_15056,N_14766,N_14554);
and U15057 (N_15057,N_14799,N_14595);
nand U15058 (N_15058,N_14605,N_14951);
or U15059 (N_15059,N_14693,N_14548);
and U15060 (N_15060,N_14781,N_14987);
and U15061 (N_15061,N_14583,N_14774);
nand U15062 (N_15062,N_14941,N_14507);
nand U15063 (N_15063,N_14924,N_14812);
nand U15064 (N_15064,N_14837,N_14971);
or U15065 (N_15065,N_14621,N_14751);
or U15066 (N_15066,N_14956,N_14597);
nand U15067 (N_15067,N_14710,N_14544);
nor U15068 (N_15068,N_14816,N_14932);
nor U15069 (N_15069,N_14986,N_14930);
and U15070 (N_15070,N_14831,N_14858);
or U15071 (N_15071,N_14627,N_14633);
or U15072 (N_15072,N_14776,N_14995);
and U15073 (N_15073,N_14773,N_14729);
and U15074 (N_15074,N_14563,N_14847);
nor U15075 (N_15075,N_14892,N_14967);
or U15076 (N_15076,N_14501,N_14819);
nand U15077 (N_15077,N_14874,N_14843);
nand U15078 (N_15078,N_14828,N_14854);
nand U15079 (N_15079,N_14724,N_14615);
and U15080 (N_15080,N_14654,N_14698);
nand U15081 (N_15081,N_14665,N_14566);
nand U15082 (N_15082,N_14981,N_14537);
and U15083 (N_15083,N_14562,N_14832);
and U15084 (N_15084,N_14916,N_14666);
xnor U15085 (N_15085,N_14500,N_14973);
or U15086 (N_15086,N_14801,N_14694);
nor U15087 (N_15087,N_14599,N_14804);
or U15088 (N_15088,N_14976,N_14985);
nor U15089 (N_15089,N_14686,N_14636);
nor U15090 (N_15090,N_14808,N_14855);
nor U15091 (N_15091,N_14840,N_14504);
nor U15092 (N_15092,N_14950,N_14662);
or U15093 (N_15093,N_14883,N_14518);
or U15094 (N_15094,N_14718,N_14639);
or U15095 (N_15095,N_14671,N_14993);
nor U15096 (N_15096,N_14959,N_14990);
nor U15097 (N_15097,N_14582,N_14620);
or U15098 (N_15098,N_14905,N_14755);
or U15099 (N_15099,N_14791,N_14960);
and U15100 (N_15100,N_14645,N_14919);
nor U15101 (N_15101,N_14589,N_14806);
xnor U15102 (N_15102,N_14997,N_14697);
or U15103 (N_15103,N_14726,N_14839);
or U15104 (N_15104,N_14975,N_14727);
or U15105 (N_15105,N_14719,N_14994);
nand U15106 (N_15106,N_14525,N_14661);
nand U15107 (N_15107,N_14535,N_14921);
and U15108 (N_15108,N_14770,N_14516);
or U15109 (N_15109,N_14579,N_14992);
nand U15110 (N_15110,N_14670,N_14747);
nor U15111 (N_15111,N_14690,N_14737);
nand U15112 (N_15112,N_14528,N_14712);
nand U15113 (N_15113,N_14646,N_14879);
nand U15114 (N_15114,N_14624,N_14846);
nor U15115 (N_15115,N_14541,N_14901);
or U15116 (N_15116,N_14920,N_14651);
or U15117 (N_15117,N_14877,N_14677);
nand U15118 (N_15118,N_14783,N_14539);
nor U15119 (N_15119,N_14641,N_14862);
nor U15120 (N_15120,N_14758,N_14767);
and U15121 (N_15121,N_14514,N_14730);
nor U15122 (N_15122,N_14836,N_14517);
nor U15123 (N_15123,N_14632,N_14585);
and U15124 (N_15124,N_14533,N_14933);
nor U15125 (N_15125,N_14771,N_14911);
and U15126 (N_15126,N_14945,N_14989);
and U15127 (N_15127,N_14861,N_14780);
or U15128 (N_15128,N_14728,N_14684);
nor U15129 (N_15129,N_14765,N_14925);
nor U15130 (N_15130,N_14853,N_14692);
nor U15131 (N_15131,N_14948,N_14884);
and U15132 (N_15132,N_14735,N_14798);
or U15133 (N_15133,N_14970,N_14587);
nor U15134 (N_15134,N_14567,N_14616);
nor U15135 (N_15135,N_14851,N_14521);
and U15136 (N_15136,N_14891,N_14978);
nand U15137 (N_15137,N_14520,N_14944);
and U15138 (N_15138,N_14870,N_14821);
nor U15139 (N_15139,N_14826,N_14707);
and U15140 (N_15140,N_14596,N_14982);
xor U15141 (N_15141,N_14818,N_14593);
xor U15142 (N_15142,N_14961,N_14505);
nor U15143 (N_15143,N_14838,N_14576);
and U15144 (N_15144,N_14570,N_14910);
and U15145 (N_15145,N_14772,N_14775);
and U15146 (N_15146,N_14820,N_14764);
and U15147 (N_15147,N_14797,N_14931);
nor U15148 (N_15148,N_14503,N_14867);
nor U15149 (N_15149,N_14529,N_14536);
or U15150 (N_15150,N_14894,N_14569);
and U15151 (N_15151,N_14705,N_14588);
nor U15152 (N_15152,N_14918,N_14913);
and U15153 (N_15153,N_14917,N_14935);
and U15154 (N_15154,N_14688,N_14709);
nand U15155 (N_15155,N_14701,N_14699);
nor U15156 (N_15156,N_14786,N_14667);
or U15157 (N_15157,N_14753,N_14619);
or U15158 (N_15158,N_14513,N_14937);
and U15159 (N_15159,N_14637,N_14790);
xor U15160 (N_15160,N_14502,N_14549);
and U15161 (N_15161,N_14509,N_14706);
nand U15162 (N_15162,N_14760,N_14897);
nor U15163 (N_15163,N_14965,N_14650);
nor U15164 (N_15164,N_14929,N_14890);
or U15165 (N_15165,N_14787,N_14757);
and U15166 (N_15166,N_14573,N_14750);
nand U15167 (N_15167,N_14756,N_14908);
and U15168 (N_15168,N_14702,N_14700);
nor U15169 (N_15169,N_14734,N_14609);
nor U15170 (N_15170,N_14784,N_14849);
nand U15171 (N_15171,N_14695,N_14631);
or U15172 (N_15172,N_14947,N_14656);
nor U15173 (N_15173,N_14893,N_14669);
nor U15174 (N_15174,N_14923,N_14789);
or U15175 (N_15175,N_14648,N_14845);
or U15176 (N_15176,N_14524,N_14928);
and U15177 (N_15177,N_14922,N_14658);
nand U15178 (N_15178,N_14672,N_14934);
nand U15179 (N_15179,N_14738,N_14895);
nand U15180 (N_15180,N_14510,N_14800);
xor U15181 (N_15181,N_14741,N_14628);
and U15182 (N_15182,N_14998,N_14966);
and U15183 (N_15183,N_14996,N_14559);
nor U15184 (N_15184,N_14792,N_14865);
nand U15185 (N_15185,N_14607,N_14963);
nor U15186 (N_15186,N_14898,N_14634);
nand U15187 (N_15187,N_14731,N_14717);
nor U15188 (N_15188,N_14655,N_14626);
and U15189 (N_15189,N_14749,N_14871);
nor U15190 (N_15190,N_14668,N_14881);
nand U15191 (N_15191,N_14657,N_14720);
or U15192 (N_15192,N_14848,N_14875);
and U15193 (N_15193,N_14685,N_14835);
nand U15194 (N_15194,N_14580,N_14594);
nand U15195 (N_15195,N_14676,N_14578);
nor U15196 (N_15196,N_14952,N_14545);
or U15197 (N_15197,N_14940,N_14696);
and U15198 (N_15198,N_14785,N_14532);
xnor U15199 (N_15199,N_14542,N_14968);
nand U15200 (N_15200,N_14768,N_14647);
or U15201 (N_15201,N_14983,N_14527);
nor U15202 (N_15202,N_14660,N_14622);
nor U15203 (N_15203,N_14778,N_14823);
nand U15204 (N_15204,N_14844,N_14522);
and U15205 (N_15205,N_14603,N_14863);
nand U15206 (N_15206,N_14926,N_14813);
or U15207 (N_15207,N_14618,N_14704);
xnor U15208 (N_15208,N_14955,N_14523);
nand U15209 (N_15209,N_14546,N_14736);
xor U15210 (N_15210,N_14904,N_14807);
nor U15211 (N_15211,N_14974,N_14581);
nand U15212 (N_15212,N_14856,N_14815);
and U15213 (N_15213,N_14824,N_14623);
nor U15214 (N_15214,N_14561,N_14878);
nand U15215 (N_15215,N_14962,N_14600);
and U15216 (N_15216,N_14610,N_14802);
or U15217 (N_15217,N_14558,N_14614);
and U15218 (N_15218,N_14664,N_14590);
or U15219 (N_15219,N_14900,N_14679);
or U15220 (N_15220,N_14829,N_14519);
and U15221 (N_15221,N_14936,N_14850);
or U15222 (N_15222,N_14689,N_14511);
nor U15223 (N_15223,N_14644,N_14914);
or U15224 (N_15224,N_14833,N_14754);
or U15225 (N_15225,N_14592,N_14591);
or U15226 (N_15226,N_14794,N_14859);
or U15227 (N_15227,N_14635,N_14551);
or U15228 (N_15228,N_14640,N_14675);
nand U15229 (N_15229,N_14811,N_14653);
nand U15230 (N_15230,N_14938,N_14613);
and U15231 (N_15231,N_14742,N_14555);
nor U15232 (N_15232,N_14680,N_14674);
or U15233 (N_15233,N_14629,N_14999);
xor U15234 (N_15234,N_14611,N_14584);
nor U15235 (N_15235,N_14857,N_14543);
nor U15236 (N_15236,N_14954,N_14984);
and U15237 (N_15237,N_14852,N_14796);
nor U15238 (N_15238,N_14969,N_14769);
nor U15239 (N_15239,N_14876,N_14608);
nor U15240 (N_15240,N_14681,N_14577);
or U15241 (N_15241,N_14887,N_14508);
and U15242 (N_15242,N_14649,N_14957);
and U15243 (N_15243,N_14715,N_14652);
nand U15244 (N_15244,N_14746,N_14953);
and U15245 (N_15245,N_14552,N_14869);
or U15246 (N_15246,N_14748,N_14678);
and U15247 (N_15247,N_14538,N_14886);
nor U15248 (N_15248,N_14872,N_14782);
xnor U15249 (N_15249,N_14880,N_14793);
nor U15250 (N_15250,N_14922,N_14700);
nor U15251 (N_15251,N_14875,N_14561);
and U15252 (N_15252,N_14703,N_14821);
or U15253 (N_15253,N_14634,N_14869);
nand U15254 (N_15254,N_14794,N_14606);
and U15255 (N_15255,N_14615,N_14585);
nand U15256 (N_15256,N_14877,N_14502);
nand U15257 (N_15257,N_14615,N_14871);
or U15258 (N_15258,N_14967,N_14681);
or U15259 (N_15259,N_14879,N_14840);
or U15260 (N_15260,N_14556,N_14648);
and U15261 (N_15261,N_14677,N_14941);
nand U15262 (N_15262,N_14633,N_14904);
nor U15263 (N_15263,N_14990,N_14814);
or U15264 (N_15264,N_14939,N_14790);
and U15265 (N_15265,N_14794,N_14759);
nor U15266 (N_15266,N_14725,N_14606);
and U15267 (N_15267,N_14779,N_14657);
or U15268 (N_15268,N_14536,N_14821);
or U15269 (N_15269,N_14964,N_14545);
nor U15270 (N_15270,N_14682,N_14975);
nor U15271 (N_15271,N_14853,N_14606);
nor U15272 (N_15272,N_14596,N_14922);
and U15273 (N_15273,N_14954,N_14698);
or U15274 (N_15274,N_14749,N_14589);
and U15275 (N_15275,N_14503,N_14623);
or U15276 (N_15276,N_14763,N_14889);
nor U15277 (N_15277,N_14586,N_14804);
nand U15278 (N_15278,N_14718,N_14742);
nor U15279 (N_15279,N_14951,N_14920);
nand U15280 (N_15280,N_14553,N_14682);
nor U15281 (N_15281,N_14604,N_14773);
nor U15282 (N_15282,N_14728,N_14742);
nor U15283 (N_15283,N_14595,N_14920);
xnor U15284 (N_15284,N_14507,N_14708);
nand U15285 (N_15285,N_14993,N_14546);
nand U15286 (N_15286,N_14755,N_14528);
xor U15287 (N_15287,N_14833,N_14987);
nand U15288 (N_15288,N_14992,N_14623);
and U15289 (N_15289,N_14968,N_14596);
nand U15290 (N_15290,N_14685,N_14680);
nor U15291 (N_15291,N_14568,N_14509);
nand U15292 (N_15292,N_14724,N_14660);
nand U15293 (N_15293,N_14762,N_14676);
nand U15294 (N_15294,N_14832,N_14648);
nor U15295 (N_15295,N_14550,N_14812);
or U15296 (N_15296,N_14928,N_14940);
nand U15297 (N_15297,N_14835,N_14566);
or U15298 (N_15298,N_14940,N_14865);
and U15299 (N_15299,N_14622,N_14862);
nor U15300 (N_15300,N_14858,N_14689);
nand U15301 (N_15301,N_14798,N_14922);
or U15302 (N_15302,N_14755,N_14562);
or U15303 (N_15303,N_14672,N_14787);
nor U15304 (N_15304,N_14795,N_14514);
nor U15305 (N_15305,N_14638,N_14672);
nand U15306 (N_15306,N_14806,N_14593);
nor U15307 (N_15307,N_14617,N_14626);
nor U15308 (N_15308,N_14817,N_14803);
or U15309 (N_15309,N_14528,N_14502);
or U15310 (N_15310,N_14868,N_14610);
and U15311 (N_15311,N_14642,N_14519);
nor U15312 (N_15312,N_14819,N_14956);
or U15313 (N_15313,N_14521,N_14515);
nand U15314 (N_15314,N_14893,N_14861);
or U15315 (N_15315,N_14931,N_14849);
or U15316 (N_15316,N_14593,N_14975);
or U15317 (N_15317,N_14527,N_14525);
nand U15318 (N_15318,N_14640,N_14739);
nor U15319 (N_15319,N_14990,N_14982);
or U15320 (N_15320,N_14807,N_14611);
or U15321 (N_15321,N_14724,N_14503);
nor U15322 (N_15322,N_14615,N_14888);
nand U15323 (N_15323,N_14532,N_14884);
and U15324 (N_15324,N_14609,N_14929);
nor U15325 (N_15325,N_14561,N_14927);
nor U15326 (N_15326,N_14556,N_14923);
or U15327 (N_15327,N_14964,N_14537);
and U15328 (N_15328,N_14924,N_14907);
nand U15329 (N_15329,N_14638,N_14905);
nand U15330 (N_15330,N_14509,N_14596);
nor U15331 (N_15331,N_14867,N_14818);
nor U15332 (N_15332,N_14524,N_14557);
nor U15333 (N_15333,N_14754,N_14982);
nand U15334 (N_15334,N_14518,N_14787);
nand U15335 (N_15335,N_14570,N_14535);
and U15336 (N_15336,N_14960,N_14789);
and U15337 (N_15337,N_14972,N_14584);
or U15338 (N_15338,N_14682,N_14839);
and U15339 (N_15339,N_14836,N_14965);
and U15340 (N_15340,N_14808,N_14776);
nor U15341 (N_15341,N_14670,N_14715);
or U15342 (N_15342,N_14974,N_14973);
nor U15343 (N_15343,N_14946,N_14943);
or U15344 (N_15344,N_14614,N_14576);
xnor U15345 (N_15345,N_14990,N_14797);
nand U15346 (N_15346,N_14815,N_14775);
nand U15347 (N_15347,N_14655,N_14566);
and U15348 (N_15348,N_14605,N_14762);
nor U15349 (N_15349,N_14601,N_14961);
xor U15350 (N_15350,N_14937,N_14618);
and U15351 (N_15351,N_14715,N_14576);
or U15352 (N_15352,N_14617,N_14589);
or U15353 (N_15353,N_14562,N_14649);
or U15354 (N_15354,N_14708,N_14859);
and U15355 (N_15355,N_14624,N_14941);
nand U15356 (N_15356,N_14502,N_14980);
or U15357 (N_15357,N_14956,N_14667);
nor U15358 (N_15358,N_14928,N_14528);
nand U15359 (N_15359,N_14990,N_14992);
nand U15360 (N_15360,N_14729,N_14569);
or U15361 (N_15361,N_14579,N_14786);
and U15362 (N_15362,N_14997,N_14735);
nor U15363 (N_15363,N_14859,N_14743);
nand U15364 (N_15364,N_14756,N_14599);
and U15365 (N_15365,N_14792,N_14782);
nor U15366 (N_15366,N_14981,N_14996);
or U15367 (N_15367,N_14980,N_14886);
or U15368 (N_15368,N_14606,N_14786);
and U15369 (N_15369,N_14848,N_14817);
nor U15370 (N_15370,N_14849,N_14912);
xnor U15371 (N_15371,N_14761,N_14785);
nand U15372 (N_15372,N_14855,N_14769);
nor U15373 (N_15373,N_14538,N_14602);
and U15374 (N_15374,N_14681,N_14653);
nand U15375 (N_15375,N_14984,N_14663);
xor U15376 (N_15376,N_14764,N_14754);
xor U15377 (N_15377,N_14969,N_14988);
or U15378 (N_15378,N_14831,N_14748);
and U15379 (N_15379,N_14659,N_14613);
and U15380 (N_15380,N_14599,N_14657);
or U15381 (N_15381,N_14878,N_14865);
nor U15382 (N_15382,N_14768,N_14907);
nand U15383 (N_15383,N_14625,N_14938);
or U15384 (N_15384,N_14981,N_14902);
and U15385 (N_15385,N_14518,N_14834);
and U15386 (N_15386,N_14770,N_14514);
or U15387 (N_15387,N_14994,N_14805);
and U15388 (N_15388,N_14838,N_14563);
nand U15389 (N_15389,N_14733,N_14763);
nor U15390 (N_15390,N_14533,N_14730);
xor U15391 (N_15391,N_14832,N_14919);
nand U15392 (N_15392,N_14834,N_14794);
and U15393 (N_15393,N_14790,N_14559);
nor U15394 (N_15394,N_14919,N_14813);
nor U15395 (N_15395,N_14902,N_14793);
nand U15396 (N_15396,N_14931,N_14667);
or U15397 (N_15397,N_14876,N_14940);
nand U15398 (N_15398,N_14837,N_14968);
nor U15399 (N_15399,N_14851,N_14849);
nor U15400 (N_15400,N_14822,N_14753);
nand U15401 (N_15401,N_14816,N_14585);
or U15402 (N_15402,N_14821,N_14962);
and U15403 (N_15403,N_14792,N_14749);
or U15404 (N_15404,N_14815,N_14702);
or U15405 (N_15405,N_14938,N_14560);
xnor U15406 (N_15406,N_14677,N_14828);
and U15407 (N_15407,N_14843,N_14719);
nor U15408 (N_15408,N_14595,N_14731);
nor U15409 (N_15409,N_14556,N_14778);
or U15410 (N_15410,N_14788,N_14515);
nor U15411 (N_15411,N_14521,N_14957);
nor U15412 (N_15412,N_14941,N_14687);
or U15413 (N_15413,N_14602,N_14582);
nand U15414 (N_15414,N_14931,N_14621);
nand U15415 (N_15415,N_14988,N_14789);
nor U15416 (N_15416,N_14846,N_14762);
or U15417 (N_15417,N_14932,N_14561);
nand U15418 (N_15418,N_14740,N_14915);
nor U15419 (N_15419,N_14521,N_14770);
nor U15420 (N_15420,N_14732,N_14951);
nor U15421 (N_15421,N_14715,N_14559);
nand U15422 (N_15422,N_14808,N_14864);
nor U15423 (N_15423,N_14811,N_14820);
or U15424 (N_15424,N_14520,N_14837);
nand U15425 (N_15425,N_14544,N_14564);
nor U15426 (N_15426,N_14857,N_14867);
or U15427 (N_15427,N_14554,N_14581);
xnor U15428 (N_15428,N_14756,N_14846);
xor U15429 (N_15429,N_14881,N_14928);
nor U15430 (N_15430,N_14532,N_14724);
xor U15431 (N_15431,N_14797,N_14710);
and U15432 (N_15432,N_14657,N_14848);
nor U15433 (N_15433,N_14566,N_14703);
or U15434 (N_15434,N_14680,N_14837);
xor U15435 (N_15435,N_14754,N_14948);
nor U15436 (N_15436,N_14842,N_14677);
xnor U15437 (N_15437,N_14645,N_14760);
nand U15438 (N_15438,N_14594,N_14624);
nand U15439 (N_15439,N_14996,N_14636);
nand U15440 (N_15440,N_14841,N_14940);
nand U15441 (N_15441,N_14834,N_14859);
or U15442 (N_15442,N_14837,N_14572);
nand U15443 (N_15443,N_14621,N_14787);
or U15444 (N_15444,N_14942,N_14578);
nor U15445 (N_15445,N_14552,N_14850);
xor U15446 (N_15446,N_14712,N_14633);
and U15447 (N_15447,N_14557,N_14634);
and U15448 (N_15448,N_14600,N_14847);
nand U15449 (N_15449,N_14683,N_14857);
xor U15450 (N_15450,N_14568,N_14681);
xnor U15451 (N_15451,N_14764,N_14749);
or U15452 (N_15452,N_14860,N_14817);
or U15453 (N_15453,N_14852,N_14994);
or U15454 (N_15454,N_14790,N_14510);
and U15455 (N_15455,N_14842,N_14980);
xnor U15456 (N_15456,N_14841,N_14637);
and U15457 (N_15457,N_14578,N_14963);
and U15458 (N_15458,N_14784,N_14654);
nand U15459 (N_15459,N_14650,N_14840);
nand U15460 (N_15460,N_14853,N_14742);
and U15461 (N_15461,N_14568,N_14823);
nor U15462 (N_15462,N_14891,N_14549);
xnor U15463 (N_15463,N_14828,N_14728);
nand U15464 (N_15464,N_14529,N_14999);
nand U15465 (N_15465,N_14930,N_14922);
or U15466 (N_15466,N_14961,N_14985);
nand U15467 (N_15467,N_14966,N_14835);
and U15468 (N_15468,N_14509,N_14939);
and U15469 (N_15469,N_14503,N_14575);
or U15470 (N_15470,N_14940,N_14736);
nor U15471 (N_15471,N_14762,N_14827);
nand U15472 (N_15472,N_14609,N_14769);
nor U15473 (N_15473,N_14923,N_14908);
or U15474 (N_15474,N_14733,N_14597);
nor U15475 (N_15475,N_14873,N_14845);
xor U15476 (N_15476,N_14826,N_14562);
xor U15477 (N_15477,N_14780,N_14748);
and U15478 (N_15478,N_14759,N_14757);
nor U15479 (N_15479,N_14711,N_14697);
or U15480 (N_15480,N_14572,N_14502);
or U15481 (N_15481,N_14929,N_14531);
nand U15482 (N_15482,N_14869,N_14947);
or U15483 (N_15483,N_14524,N_14746);
and U15484 (N_15484,N_14813,N_14931);
and U15485 (N_15485,N_14885,N_14576);
or U15486 (N_15486,N_14934,N_14628);
or U15487 (N_15487,N_14797,N_14524);
and U15488 (N_15488,N_14541,N_14862);
or U15489 (N_15489,N_14709,N_14848);
or U15490 (N_15490,N_14932,N_14799);
nor U15491 (N_15491,N_14979,N_14980);
or U15492 (N_15492,N_14593,N_14658);
xor U15493 (N_15493,N_14523,N_14647);
and U15494 (N_15494,N_14696,N_14571);
nand U15495 (N_15495,N_14621,N_14677);
nand U15496 (N_15496,N_14933,N_14982);
or U15497 (N_15497,N_14972,N_14522);
nor U15498 (N_15498,N_14962,N_14893);
nand U15499 (N_15499,N_14797,N_14789);
nand U15500 (N_15500,N_15132,N_15161);
and U15501 (N_15501,N_15299,N_15203);
nand U15502 (N_15502,N_15468,N_15276);
nor U15503 (N_15503,N_15439,N_15070);
nor U15504 (N_15504,N_15195,N_15490);
nand U15505 (N_15505,N_15366,N_15165);
and U15506 (N_15506,N_15228,N_15213);
xor U15507 (N_15507,N_15475,N_15217);
or U15508 (N_15508,N_15360,N_15336);
and U15509 (N_15509,N_15303,N_15013);
xor U15510 (N_15510,N_15495,N_15214);
or U15511 (N_15511,N_15335,N_15477);
nor U15512 (N_15512,N_15371,N_15291);
or U15513 (N_15513,N_15334,N_15412);
or U15514 (N_15514,N_15038,N_15145);
xnor U15515 (N_15515,N_15426,N_15316);
and U15516 (N_15516,N_15176,N_15315);
xor U15517 (N_15517,N_15040,N_15295);
or U15518 (N_15518,N_15088,N_15318);
or U15519 (N_15519,N_15319,N_15355);
or U15520 (N_15520,N_15033,N_15251);
or U15521 (N_15521,N_15249,N_15440);
nand U15522 (N_15522,N_15274,N_15041);
nor U15523 (N_15523,N_15449,N_15459);
nor U15524 (N_15524,N_15167,N_15090);
nand U15525 (N_15525,N_15447,N_15288);
or U15526 (N_15526,N_15436,N_15317);
or U15527 (N_15527,N_15256,N_15285);
or U15528 (N_15528,N_15372,N_15064);
nor U15529 (N_15529,N_15455,N_15441);
nor U15530 (N_15530,N_15446,N_15473);
or U15531 (N_15531,N_15066,N_15414);
and U15532 (N_15532,N_15438,N_15113);
and U15533 (N_15533,N_15278,N_15400);
or U15534 (N_15534,N_15125,N_15222);
or U15535 (N_15535,N_15102,N_15467);
nor U15536 (N_15536,N_15045,N_15065);
nor U15537 (N_15537,N_15420,N_15312);
nor U15538 (N_15538,N_15331,N_15374);
nand U15539 (N_15539,N_15068,N_15133);
nand U15540 (N_15540,N_15362,N_15351);
and U15541 (N_15541,N_15164,N_15304);
nand U15542 (N_15542,N_15245,N_15286);
nor U15543 (N_15543,N_15155,N_15107);
and U15544 (N_15544,N_15175,N_15456);
or U15545 (N_15545,N_15399,N_15275);
or U15546 (N_15546,N_15387,N_15021);
or U15547 (N_15547,N_15442,N_15271);
and U15548 (N_15548,N_15212,N_15154);
nor U15549 (N_15549,N_15152,N_15158);
and U15550 (N_15550,N_15320,N_15062);
nor U15551 (N_15551,N_15029,N_15270);
or U15552 (N_15552,N_15389,N_15402);
or U15553 (N_15553,N_15224,N_15418);
nor U15554 (N_15554,N_15476,N_15244);
nor U15555 (N_15555,N_15466,N_15103);
nor U15556 (N_15556,N_15488,N_15487);
nor U15557 (N_15557,N_15483,N_15147);
xor U15558 (N_15558,N_15119,N_15173);
or U15559 (N_15559,N_15169,N_15131);
or U15560 (N_15560,N_15457,N_15392);
and U15561 (N_15561,N_15445,N_15301);
and U15562 (N_15562,N_15443,N_15397);
and U15563 (N_15563,N_15017,N_15398);
nor U15564 (N_15564,N_15142,N_15308);
nand U15565 (N_15565,N_15246,N_15128);
nand U15566 (N_15566,N_15054,N_15280);
or U15567 (N_15567,N_15451,N_15265);
or U15568 (N_15568,N_15464,N_15298);
and U15569 (N_15569,N_15363,N_15353);
and U15570 (N_15570,N_15434,N_15369);
nor U15571 (N_15571,N_15309,N_15236);
or U15572 (N_15572,N_15327,N_15004);
or U15573 (N_15573,N_15094,N_15344);
xnor U15574 (N_15574,N_15492,N_15404);
nor U15575 (N_15575,N_15302,N_15432);
nor U15576 (N_15576,N_15461,N_15043);
and U15577 (N_15577,N_15072,N_15221);
or U15578 (N_15578,N_15210,N_15453);
nand U15579 (N_15579,N_15215,N_15061);
nor U15580 (N_15580,N_15078,N_15310);
nand U15581 (N_15581,N_15023,N_15261);
nand U15582 (N_15582,N_15338,N_15325);
nand U15583 (N_15583,N_15020,N_15383);
nor U15584 (N_15584,N_15011,N_15435);
and U15585 (N_15585,N_15307,N_15352);
xnor U15586 (N_15586,N_15000,N_15294);
nand U15587 (N_15587,N_15156,N_15471);
or U15588 (N_15588,N_15124,N_15110);
nor U15589 (N_15589,N_15139,N_15148);
nor U15590 (N_15590,N_15071,N_15016);
nor U15591 (N_15591,N_15187,N_15284);
or U15592 (N_15592,N_15200,N_15034);
xnor U15593 (N_15593,N_15342,N_15401);
or U15594 (N_15594,N_15347,N_15207);
and U15595 (N_15595,N_15185,N_15204);
nor U15596 (N_15596,N_15123,N_15141);
xor U15597 (N_15597,N_15146,N_15485);
nand U15598 (N_15598,N_15364,N_15267);
or U15599 (N_15599,N_15452,N_15377);
nand U15600 (N_15600,N_15259,N_15001);
nand U15601 (N_15601,N_15015,N_15235);
nor U15602 (N_15602,N_15114,N_15462);
and U15603 (N_15603,N_15037,N_15117);
nand U15604 (N_15604,N_15425,N_15243);
nand U15605 (N_15605,N_15381,N_15049);
nor U15606 (N_15606,N_15170,N_15223);
and U15607 (N_15607,N_15480,N_15350);
nor U15608 (N_15608,N_15093,N_15100);
and U15609 (N_15609,N_15465,N_15277);
and U15610 (N_15610,N_15266,N_15340);
nand U15611 (N_15611,N_15112,N_15499);
or U15612 (N_15612,N_15050,N_15287);
nor U15613 (N_15613,N_15039,N_15463);
and U15614 (N_15614,N_15230,N_15391);
nand U15615 (N_15615,N_15348,N_15370);
nand U15616 (N_15616,N_15012,N_15422);
nor U15617 (N_15617,N_15297,N_15419);
or U15618 (N_15618,N_15082,N_15162);
or U15619 (N_15619,N_15053,N_15375);
or U15620 (N_15620,N_15014,N_15130);
nand U15621 (N_15621,N_15378,N_15010);
and U15622 (N_15622,N_15460,N_15120);
and U15623 (N_15623,N_15218,N_15448);
xor U15624 (N_15624,N_15240,N_15163);
or U15625 (N_15625,N_15356,N_15408);
or U15626 (N_15626,N_15421,N_15205);
or U15627 (N_15627,N_15086,N_15498);
nand U15628 (N_15628,N_15314,N_15354);
or U15629 (N_15629,N_15191,N_15493);
nor U15630 (N_15630,N_15368,N_15181);
xor U15631 (N_15631,N_15027,N_15046);
nand U15632 (N_15632,N_15178,N_15345);
or U15633 (N_15633,N_15386,N_15388);
or U15634 (N_15634,N_15024,N_15239);
or U15635 (N_15635,N_15056,N_15198);
or U15636 (N_15636,N_15144,N_15211);
nand U15637 (N_15637,N_15326,N_15036);
or U15638 (N_15638,N_15450,N_15143);
nor U15639 (N_15639,N_15127,N_15116);
xor U15640 (N_15640,N_15136,N_15006);
and U15641 (N_15641,N_15098,N_15115);
or U15642 (N_15642,N_15379,N_15192);
nor U15643 (N_15643,N_15233,N_15196);
or U15644 (N_15644,N_15324,N_15407);
or U15645 (N_15645,N_15341,N_15097);
or U15646 (N_15646,N_15232,N_15415);
or U15647 (N_15647,N_15253,N_15394);
or U15648 (N_15648,N_15227,N_15486);
and U15649 (N_15649,N_15026,N_15199);
xor U15650 (N_15650,N_15365,N_15052);
or U15651 (N_15651,N_15151,N_15323);
nor U15652 (N_15652,N_15279,N_15108);
and U15653 (N_15653,N_15393,N_15427);
and U15654 (N_15654,N_15484,N_15497);
xor U15655 (N_15655,N_15454,N_15060);
nand U15656 (N_15656,N_15157,N_15329);
nand U15657 (N_15657,N_15423,N_15059);
or U15658 (N_15658,N_15359,N_15332);
or U15659 (N_15659,N_15126,N_15376);
xor U15660 (N_15660,N_15106,N_15409);
or U15661 (N_15661,N_15349,N_15208);
and U15662 (N_15662,N_15373,N_15343);
nor U15663 (N_15663,N_15197,N_15109);
or U15664 (N_15664,N_15219,N_15009);
nor U15665 (N_15665,N_15346,N_15382);
or U15666 (N_15666,N_15283,N_15067);
and U15667 (N_15667,N_15403,N_15247);
and U15668 (N_15668,N_15289,N_15075);
or U15669 (N_15669,N_15395,N_15002);
nand U15670 (N_15670,N_15008,N_15361);
or U15671 (N_15671,N_15481,N_15472);
nand U15672 (N_15672,N_15242,N_15380);
nand U15673 (N_15673,N_15444,N_15272);
or U15674 (N_15674,N_15296,N_15140);
nor U15675 (N_15675,N_15051,N_15031);
and U15676 (N_15676,N_15339,N_15225);
or U15677 (N_15677,N_15081,N_15413);
and U15678 (N_15678,N_15311,N_15135);
nor U15679 (N_15679,N_15428,N_15069);
or U15680 (N_15680,N_15105,N_15092);
nand U15681 (N_15681,N_15258,N_15030);
and U15682 (N_15682,N_15216,N_15085);
or U15683 (N_15683,N_15206,N_15474);
nand U15684 (N_15684,N_15188,N_15183);
nand U15685 (N_15685,N_15087,N_15405);
nor U15686 (N_15686,N_15057,N_15171);
nor U15687 (N_15687,N_15255,N_15293);
or U15688 (N_15688,N_15194,N_15305);
or U15689 (N_15689,N_15313,N_15149);
nand U15690 (N_15690,N_15250,N_15469);
nor U15691 (N_15691,N_15264,N_15055);
and U15692 (N_15692,N_15063,N_15025);
nand U15693 (N_15693,N_15073,N_15084);
nor U15694 (N_15694,N_15234,N_15269);
nand U15695 (N_15695,N_15410,N_15074);
and U15696 (N_15696,N_15478,N_15189);
and U15697 (N_15697,N_15238,N_15411);
and U15698 (N_15698,N_15077,N_15416);
nand U15699 (N_15699,N_15138,N_15166);
nand U15700 (N_15700,N_15384,N_15035);
nor U15701 (N_15701,N_15179,N_15281);
and U15702 (N_15702,N_15032,N_15385);
and U15703 (N_15703,N_15172,N_15328);
xor U15704 (N_15704,N_15470,N_15091);
or U15705 (N_15705,N_15430,N_15058);
or U15706 (N_15706,N_15083,N_15458);
nand U15707 (N_15707,N_15160,N_15186);
nand U15708 (N_15708,N_15177,N_15231);
nor U15709 (N_15709,N_15337,N_15491);
nand U15710 (N_15710,N_15202,N_15321);
and U15711 (N_15711,N_15431,N_15229);
nand U15712 (N_15712,N_15417,N_15079);
xnor U15713 (N_15713,N_15424,N_15209);
and U15714 (N_15714,N_15080,N_15153);
and U15715 (N_15715,N_15095,N_15019);
nor U15716 (N_15716,N_15122,N_15494);
or U15717 (N_15717,N_15159,N_15190);
xnor U15718 (N_15718,N_15273,N_15300);
or U15719 (N_15719,N_15322,N_15096);
and U15720 (N_15720,N_15252,N_15201);
nor U15721 (N_15721,N_15099,N_15101);
and U15722 (N_15722,N_15260,N_15005);
nor U15723 (N_15723,N_15184,N_15263);
xnor U15724 (N_15724,N_15357,N_15134);
nand U15725 (N_15725,N_15121,N_15429);
nor U15726 (N_15726,N_15168,N_15174);
or U15727 (N_15727,N_15433,N_15262);
nor U15728 (N_15728,N_15237,N_15268);
xor U15729 (N_15729,N_15282,N_15390);
and U15730 (N_15730,N_15129,N_15048);
and U15731 (N_15731,N_15118,N_15290);
xor U15732 (N_15732,N_15226,N_15104);
nor U15733 (N_15733,N_15479,N_15111);
and U15734 (N_15734,N_15076,N_15496);
nand U15735 (N_15735,N_15330,N_15358);
nand U15736 (N_15736,N_15137,N_15180);
or U15737 (N_15737,N_15007,N_15089);
and U15738 (N_15738,N_15220,N_15292);
nor U15739 (N_15739,N_15150,N_15367);
and U15740 (N_15740,N_15042,N_15241);
xor U15741 (N_15741,N_15028,N_15437);
and U15742 (N_15742,N_15018,N_15003);
or U15743 (N_15743,N_15489,N_15193);
xnor U15744 (N_15744,N_15044,N_15333);
and U15745 (N_15745,N_15047,N_15396);
nand U15746 (N_15746,N_15257,N_15254);
nand U15747 (N_15747,N_15022,N_15306);
nor U15748 (N_15748,N_15406,N_15482);
xnor U15749 (N_15749,N_15182,N_15248);
nand U15750 (N_15750,N_15262,N_15468);
nor U15751 (N_15751,N_15486,N_15301);
nand U15752 (N_15752,N_15326,N_15398);
and U15753 (N_15753,N_15110,N_15389);
and U15754 (N_15754,N_15426,N_15238);
xor U15755 (N_15755,N_15118,N_15435);
nor U15756 (N_15756,N_15410,N_15313);
and U15757 (N_15757,N_15213,N_15141);
and U15758 (N_15758,N_15028,N_15152);
nand U15759 (N_15759,N_15431,N_15370);
xnor U15760 (N_15760,N_15324,N_15211);
nand U15761 (N_15761,N_15108,N_15240);
nor U15762 (N_15762,N_15128,N_15353);
and U15763 (N_15763,N_15301,N_15059);
and U15764 (N_15764,N_15332,N_15144);
nand U15765 (N_15765,N_15438,N_15332);
nand U15766 (N_15766,N_15266,N_15071);
xor U15767 (N_15767,N_15413,N_15276);
or U15768 (N_15768,N_15255,N_15449);
or U15769 (N_15769,N_15125,N_15049);
nand U15770 (N_15770,N_15363,N_15235);
nor U15771 (N_15771,N_15315,N_15294);
and U15772 (N_15772,N_15131,N_15069);
and U15773 (N_15773,N_15367,N_15479);
nand U15774 (N_15774,N_15377,N_15297);
and U15775 (N_15775,N_15405,N_15040);
nand U15776 (N_15776,N_15273,N_15461);
nand U15777 (N_15777,N_15442,N_15023);
nor U15778 (N_15778,N_15496,N_15396);
or U15779 (N_15779,N_15119,N_15121);
and U15780 (N_15780,N_15048,N_15244);
nand U15781 (N_15781,N_15451,N_15096);
nand U15782 (N_15782,N_15357,N_15440);
and U15783 (N_15783,N_15098,N_15013);
xnor U15784 (N_15784,N_15374,N_15161);
and U15785 (N_15785,N_15350,N_15455);
or U15786 (N_15786,N_15075,N_15390);
nor U15787 (N_15787,N_15451,N_15086);
nor U15788 (N_15788,N_15087,N_15457);
nor U15789 (N_15789,N_15366,N_15446);
or U15790 (N_15790,N_15036,N_15111);
and U15791 (N_15791,N_15435,N_15347);
xnor U15792 (N_15792,N_15213,N_15244);
nand U15793 (N_15793,N_15002,N_15213);
xor U15794 (N_15794,N_15468,N_15013);
xor U15795 (N_15795,N_15385,N_15057);
nand U15796 (N_15796,N_15319,N_15044);
nand U15797 (N_15797,N_15069,N_15444);
nand U15798 (N_15798,N_15255,N_15466);
xnor U15799 (N_15799,N_15064,N_15169);
nor U15800 (N_15800,N_15193,N_15468);
nand U15801 (N_15801,N_15294,N_15245);
nor U15802 (N_15802,N_15248,N_15359);
and U15803 (N_15803,N_15337,N_15250);
nor U15804 (N_15804,N_15279,N_15250);
nand U15805 (N_15805,N_15301,N_15485);
or U15806 (N_15806,N_15164,N_15443);
nand U15807 (N_15807,N_15099,N_15242);
or U15808 (N_15808,N_15194,N_15009);
nand U15809 (N_15809,N_15020,N_15118);
or U15810 (N_15810,N_15470,N_15274);
xor U15811 (N_15811,N_15092,N_15268);
and U15812 (N_15812,N_15313,N_15481);
nand U15813 (N_15813,N_15200,N_15202);
nand U15814 (N_15814,N_15110,N_15191);
or U15815 (N_15815,N_15297,N_15208);
or U15816 (N_15816,N_15021,N_15214);
nor U15817 (N_15817,N_15470,N_15108);
or U15818 (N_15818,N_15240,N_15336);
nor U15819 (N_15819,N_15276,N_15193);
nand U15820 (N_15820,N_15403,N_15168);
xnor U15821 (N_15821,N_15253,N_15176);
and U15822 (N_15822,N_15437,N_15237);
nand U15823 (N_15823,N_15251,N_15423);
nand U15824 (N_15824,N_15463,N_15270);
or U15825 (N_15825,N_15105,N_15073);
nand U15826 (N_15826,N_15437,N_15289);
xor U15827 (N_15827,N_15462,N_15277);
nand U15828 (N_15828,N_15468,N_15347);
nand U15829 (N_15829,N_15123,N_15291);
nor U15830 (N_15830,N_15408,N_15271);
xnor U15831 (N_15831,N_15074,N_15434);
nand U15832 (N_15832,N_15192,N_15155);
nand U15833 (N_15833,N_15154,N_15075);
and U15834 (N_15834,N_15172,N_15250);
nand U15835 (N_15835,N_15331,N_15266);
nor U15836 (N_15836,N_15002,N_15375);
or U15837 (N_15837,N_15398,N_15169);
nand U15838 (N_15838,N_15187,N_15173);
nor U15839 (N_15839,N_15031,N_15070);
and U15840 (N_15840,N_15290,N_15372);
or U15841 (N_15841,N_15001,N_15140);
or U15842 (N_15842,N_15198,N_15341);
xor U15843 (N_15843,N_15409,N_15261);
xor U15844 (N_15844,N_15292,N_15117);
nor U15845 (N_15845,N_15141,N_15017);
and U15846 (N_15846,N_15131,N_15136);
nor U15847 (N_15847,N_15205,N_15222);
and U15848 (N_15848,N_15008,N_15484);
or U15849 (N_15849,N_15120,N_15393);
and U15850 (N_15850,N_15271,N_15288);
xnor U15851 (N_15851,N_15371,N_15286);
and U15852 (N_15852,N_15197,N_15078);
nand U15853 (N_15853,N_15373,N_15251);
nor U15854 (N_15854,N_15001,N_15460);
or U15855 (N_15855,N_15110,N_15112);
or U15856 (N_15856,N_15061,N_15268);
or U15857 (N_15857,N_15359,N_15239);
nor U15858 (N_15858,N_15454,N_15144);
nor U15859 (N_15859,N_15410,N_15368);
xnor U15860 (N_15860,N_15354,N_15128);
nor U15861 (N_15861,N_15317,N_15427);
and U15862 (N_15862,N_15348,N_15444);
and U15863 (N_15863,N_15062,N_15486);
nor U15864 (N_15864,N_15395,N_15171);
nand U15865 (N_15865,N_15485,N_15110);
nand U15866 (N_15866,N_15367,N_15361);
or U15867 (N_15867,N_15252,N_15164);
nor U15868 (N_15868,N_15141,N_15167);
nand U15869 (N_15869,N_15119,N_15332);
or U15870 (N_15870,N_15107,N_15275);
or U15871 (N_15871,N_15454,N_15282);
or U15872 (N_15872,N_15225,N_15368);
xor U15873 (N_15873,N_15340,N_15230);
nor U15874 (N_15874,N_15225,N_15168);
or U15875 (N_15875,N_15343,N_15145);
or U15876 (N_15876,N_15066,N_15247);
nand U15877 (N_15877,N_15015,N_15323);
and U15878 (N_15878,N_15231,N_15356);
nor U15879 (N_15879,N_15071,N_15229);
nand U15880 (N_15880,N_15011,N_15474);
and U15881 (N_15881,N_15089,N_15165);
xnor U15882 (N_15882,N_15363,N_15104);
nor U15883 (N_15883,N_15483,N_15408);
nand U15884 (N_15884,N_15067,N_15285);
nor U15885 (N_15885,N_15138,N_15073);
and U15886 (N_15886,N_15065,N_15274);
and U15887 (N_15887,N_15270,N_15085);
nand U15888 (N_15888,N_15071,N_15434);
nand U15889 (N_15889,N_15401,N_15409);
nand U15890 (N_15890,N_15212,N_15462);
nor U15891 (N_15891,N_15175,N_15004);
nand U15892 (N_15892,N_15040,N_15485);
nand U15893 (N_15893,N_15023,N_15453);
nand U15894 (N_15894,N_15330,N_15105);
or U15895 (N_15895,N_15360,N_15230);
nand U15896 (N_15896,N_15235,N_15161);
nand U15897 (N_15897,N_15472,N_15159);
xor U15898 (N_15898,N_15000,N_15251);
nor U15899 (N_15899,N_15458,N_15121);
or U15900 (N_15900,N_15207,N_15064);
or U15901 (N_15901,N_15057,N_15479);
nand U15902 (N_15902,N_15489,N_15299);
and U15903 (N_15903,N_15319,N_15281);
and U15904 (N_15904,N_15024,N_15141);
nand U15905 (N_15905,N_15017,N_15336);
or U15906 (N_15906,N_15458,N_15369);
xnor U15907 (N_15907,N_15220,N_15235);
nor U15908 (N_15908,N_15436,N_15023);
xnor U15909 (N_15909,N_15128,N_15231);
or U15910 (N_15910,N_15246,N_15069);
and U15911 (N_15911,N_15338,N_15152);
and U15912 (N_15912,N_15086,N_15396);
or U15913 (N_15913,N_15378,N_15399);
and U15914 (N_15914,N_15247,N_15074);
or U15915 (N_15915,N_15227,N_15264);
nand U15916 (N_15916,N_15011,N_15476);
and U15917 (N_15917,N_15256,N_15396);
or U15918 (N_15918,N_15463,N_15236);
or U15919 (N_15919,N_15140,N_15183);
nand U15920 (N_15920,N_15135,N_15373);
nor U15921 (N_15921,N_15242,N_15483);
nand U15922 (N_15922,N_15008,N_15471);
nand U15923 (N_15923,N_15340,N_15086);
and U15924 (N_15924,N_15053,N_15157);
or U15925 (N_15925,N_15174,N_15219);
or U15926 (N_15926,N_15379,N_15198);
and U15927 (N_15927,N_15149,N_15025);
nand U15928 (N_15928,N_15291,N_15409);
nand U15929 (N_15929,N_15101,N_15413);
nand U15930 (N_15930,N_15472,N_15304);
and U15931 (N_15931,N_15280,N_15139);
nand U15932 (N_15932,N_15139,N_15021);
xor U15933 (N_15933,N_15039,N_15440);
nand U15934 (N_15934,N_15148,N_15384);
or U15935 (N_15935,N_15320,N_15364);
nand U15936 (N_15936,N_15112,N_15018);
and U15937 (N_15937,N_15226,N_15076);
or U15938 (N_15938,N_15323,N_15373);
or U15939 (N_15939,N_15279,N_15243);
nand U15940 (N_15940,N_15180,N_15220);
nand U15941 (N_15941,N_15063,N_15050);
nor U15942 (N_15942,N_15457,N_15222);
nand U15943 (N_15943,N_15208,N_15326);
and U15944 (N_15944,N_15003,N_15460);
nand U15945 (N_15945,N_15092,N_15148);
nand U15946 (N_15946,N_15298,N_15078);
and U15947 (N_15947,N_15298,N_15228);
nand U15948 (N_15948,N_15439,N_15137);
nor U15949 (N_15949,N_15043,N_15072);
and U15950 (N_15950,N_15258,N_15014);
or U15951 (N_15951,N_15143,N_15087);
or U15952 (N_15952,N_15131,N_15250);
and U15953 (N_15953,N_15182,N_15369);
or U15954 (N_15954,N_15431,N_15263);
nor U15955 (N_15955,N_15142,N_15117);
and U15956 (N_15956,N_15323,N_15241);
or U15957 (N_15957,N_15149,N_15240);
or U15958 (N_15958,N_15302,N_15196);
xnor U15959 (N_15959,N_15418,N_15378);
nor U15960 (N_15960,N_15283,N_15114);
nand U15961 (N_15961,N_15229,N_15419);
nor U15962 (N_15962,N_15474,N_15018);
nor U15963 (N_15963,N_15002,N_15108);
nand U15964 (N_15964,N_15158,N_15130);
xnor U15965 (N_15965,N_15030,N_15117);
nand U15966 (N_15966,N_15131,N_15409);
or U15967 (N_15967,N_15188,N_15100);
nor U15968 (N_15968,N_15114,N_15192);
or U15969 (N_15969,N_15231,N_15443);
and U15970 (N_15970,N_15421,N_15215);
nand U15971 (N_15971,N_15333,N_15236);
or U15972 (N_15972,N_15353,N_15204);
nor U15973 (N_15973,N_15498,N_15209);
and U15974 (N_15974,N_15358,N_15069);
nor U15975 (N_15975,N_15008,N_15104);
nand U15976 (N_15976,N_15395,N_15435);
or U15977 (N_15977,N_15234,N_15015);
and U15978 (N_15978,N_15090,N_15351);
xnor U15979 (N_15979,N_15374,N_15438);
xor U15980 (N_15980,N_15386,N_15465);
nand U15981 (N_15981,N_15046,N_15364);
and U15982 (N_15982,N_15037,N_15108);
nor U15983 (N_15983,N_15204,N_15137);
nor U15984 (N_15984,N_15043,N_15209);
nor U15985 (N_15985,N_15363,N_15236);
nor U15986 (N_15986,N_15214,N_15287);
nand U15987 (N_15987,N_15329,N_15100);
nand U15988 (N_15988,N_15020,N_15146);
and U15989 (N_15989,N_15353,N_15346);
nor U15990 (N_15990,N_15162,N_15348);
nand U15991 (N_15991,N_15030,N_15044);
xnor U15992 (N_15992,N_15324,N_15104);
or U15993 (N_15993,N_15041,N_15229);
nand U15994 (N_15994,N_15108,N_15066);
nand U15995 (N_15995,N_15438,N_15390);
nor U15996 (N_15996,N_15141,N_15042);
and U15997 (N_15997,N_15289,N_15140);
and U15998 (N_15998,N_15019,N_15384);
xor U15999 (N_15999,N_15467,N_15430);
nor U16000 (N_16000,N_15647,N_15913);
or U16001 (N_16001,N_15739,N_15535);
or U16002 (N_16002,N_15598,N_15650);
xnor U16003 (N_16003,N_15893,N_15867);
xnor U16004 (N_16004,N_15555,N_15736);
nand U16005 (N_16005,N_15824,N_15670);
nand U16006 (N_16006,N_15511,N_15892);
and U16007 (N_16007,N_15671,N_15741);
or U16008 (N_16008,N_15789,N_15928);
or U16009 (N_16009,N_15742,N_15768);
or U16010 (N_16010,N_15515,N_15680);
nor U16011 (N_16011,N_15596,N_15641);
nor U16012 (N_16012,N_15600,N_15534);
nor U16013 (N_16013,N_15510,N_15926);
or U16014 (N_16014,N_15805,N_15947);
xnor U16015 (N_16015,N_15801,N_15646);
or U16016 (N_16016,N_15716,N_15575);
or U16017 (N_16017,N_15514,N_15621);
and U16018 (N_16018,N_15862,N_15669);
nand U16019 (N_16019,N_15725,N_15830);
or U16020 (N_16020,N_15744,N_15677);
or U16021 (N_16021,N_15577,N_15727);
and U16022 (N_16022,N_15502,N_15729);
nand U16023 (N_16023,N_15775,N_15886);
or U16024 (N_16024,N_15539,N_15977);
nor U16025 (N_16025,N_15948,N_15910);
and U16026 (N_16026,N_15975,N_15642);
and U16027 (N_16027,N_15780,N_15936);
and U16028 (N_16028,N_15664,N_15961);
xnor U16029 (N_16029,N_15553,N_15818);
and U16030 (N_16030,N_15749,N_15964);
xnor U16031 (N_16031,N_15812,N_15632);
nor U16032 (N_16032,N_15651,N_15732);
and U16033 (N_16033,N_15663,N_15603);
and U16034 (N_16034,N_15792,N_15526);
or U16035 (N_16035,N_15513,N_15687);
nor U16036 (N_16036,N_15631,N_15797);
and U16037 (N_16037,N_15639,N_15622);
or U16038 (N_16038,N_15833,N_15943);
nor U16039 (N_16039,N_15579,N_15836);
or U16040 (N_16040,N_15740,N_15815);
nand U16041 (N_16041,N_15724,N_15564);
nor U16042 (N_16042,N_15710,N_15831);
nor U16043 (N_16043,N_15745,N_15626);
or U16044 (N_16044,N_15887,N_15751);
nor U16045 (N_16045,N_15849,N_15601);
nor U16046 (N_16046,N_15552,N_15547);
nand U16047 (N_16047,N_15912,N_15630);
nand U16048 (N_16048,N_15860,N_15512);
nand U16049 (N_16049,N_15619,N_15755);
nor U16050 (N_16050,N_15994,N_15814);
nand U16051 (N_16051,N_15854,N_15690);
nand U16052 (N_16052,N_15519,N_15707);
or U16053 (N_16053,N_15859,N_15907);
xnor U16054 (N_16054,N_15866,N_15802);
and U16055 (N_16055,N_15712,N_15784);
and U16056 (N_16056,N_15652,N_15640);
nor U16057 (N_16057,N_15923,N_15655);
nor U16058 (N_16058,N_15999,N_15604);
and U16059 (N_16059,N_15997,N_15902);
nor U16060 (N_16060,N_15672,N_15599);
nor U16061 (N_16061,N_15982,N_15843);
nand U16062 (N_16062,N_15696,N_15826);
xnor U16063 (N_16063,N_15901,N_15549);
xnor U16064 (N_16064,N_15605,N_15819);
nand U16065 (N_16065,N_15609,N_15827);
or U16066 (N_16066,N_15572,N_15798);
nand U16067 (N_16067,N_15897,N_15558);
nor U16068 (N_16068,N_15846,N_15582);
and U16069 (N_16069,N_15532,N_15697);
xor U16070 (N_16070,N_15571,N_15538);
nor U16071 (N_16071,N_15618,N_15816);
and U16072 (N_16072,N_15813,N_15635);
and U16073 (N_16073,N_15656,N_15654);
nor U16074 (N_16074,N_15828,N_15963);
nor U16075 (N_16075,N_15971,N_15962);
nand U16076 (N_16076,N_15611,N_15995);
and U16077 (N_16077,N_15684,N_15734);
and U16078 (N_16078,N_15911,N_15983);
nor U16079 (N_16079,N_15884,N_15730);
nor U16080 (N_16080,N_15883,N_15844);
and U16081 (N_16081,N_15726,N_15638);
nor U16082 (N_16082,N_15706,N_15541);
or U16083 (N_16083,N_15820,N_15771);
and U16084 (N_16084,N_15597,N_15972);
or U16085 (N_16085,N_15533,N_15675);
or U16086 (N_16086,N_15855,N_15842);
or U16087 (N_16087,N_15701,N_15984);
and U16088 (N_16088,N_15550,N_15737);
nor U16089 (N_16089,N_15998,N_15607);
or U16090 (N_16090,N_15950,N_15914);
and U16091 (N_16091,N_15834,N_15803);
nor U16092 (N_16092,N_15864,N_15505);
xor U16093 (N_16093,N_15665,N_15590);
xnor U16094 (N_16094,N_15685,N_15688);
nor U16095 (N_16095,N_15958,N_15960);
or U16096 (N_16096,N_15880,N_15625);
nor U16097 (N_16097,N_15700,N_15856);
and U16098 (N_16098,N_15698,N_15979);
or U16099 (N_16099,N_15874,N_15628);
nand U16100 (N_16100,N_15569,N_15714);
or U16101 (N_16101,N_15536,N_15557);
or U16102 (N_16102,N_15903,N_15996);
nor U16103 (N_16103,N_15989,N_15785);
xnor U16104 (N_16104,N_15981,N_15986);
nand U16105 (N_16105,N_15882,N_15787);
and U16106 (N_16106,N_15674,N_15758);
or U16107 (N_16107,N_15681,N_15545);
and U16108 (N_16108,N_15929,N_15861);
xor U16109 (N_16109,N_15668,N_15506);
nor U16110 (N_16110,N_15602,N_15643);
and U16111 (N_16111,N_15917,N_15645);
xnor U16112 (N_16112,N_15660,N_15937);
or U16113 (N_16113,N_15835,N_15786);
or U16114 (N_16114,N_15992,N_15817);
and U16115 (N_16115,N_15543,N_15870);
nand U16116 (N_16116,N_15863,N_15587);
nor U16117 (N_16117,N_15774,N_15586);
nand U16118 (N_16118,N_15591,N_15916);
and U16119 (N_16119,N_15537,N_15548);
nor U16120 (N_16120,N_15779,N_15847);
nor U16121 (N_16121,N_15795,N_15560);
and U16122 (N_16122,N_15561,N_15759);
or U16123 (N_16123,N_15872,N_15578);
nor U16124 (N_16124,N_15869,N_15829);
xnor U16125 (N_16125,N_15918,N_15951);
nand U16126 (N_16126,N_15889,N_15679);
nand U16127 (N_16127,N_15851,N_15702);
nor U16128 (N_16128,N_15973,N_15501);
or U16129 (N_16129,N_15503,N_15898);
and U16130 (N_16130,N_15633,N_15781);
and U16131 (N_16131,N_15959,N_15920);
nor U16132 (N_16132,N_15517,N_15704);
and U16133 (N_16133,N_15508,N_15765);
nand U16134 (N_16134,N_15764,N_15763);
nor U16135 (N_16135,N_15676,N_15877);
and U16136 (N_16136,N_15772,N_15809);
nand U16137 (N_16137,N_15615,N_15556);
and U16138 (N_16138,N_15875,N_15769);
nand U16139 (N_16139,N_15623,N_15673);
nor U16140 (N_16140,N_15988,N_15617);
nand U16141 (N_16141,N_15717,N_15594);
and U16142 (N_16142,N_15715,N_15757);
and U16143 (N_16143,N_15993,N_15927);
xor U16144 (N_16144,N_15858,N_15531);
nor U16145 (N_16145,N_15791,N_15566);
nor U16146 (N_16146,N_15832,N_15748);
xnor U16147 (N_16147,N_15529,N_15906);
and U16148 (N_16148,N_15807,N_15967);
nor U16149 (N_16149,N_15581,N_15788);
nor U16150 (N_16150,N_15709,N_15689);
xnor U16151 (N_16151,N_15990,N_15796);
and U16152 (N_16152,N_15551,N_15793);
nand U16153 (N_16153,N_15661,N_15778);
xor U16154 (N_16154,N_15921,N_15747);
nor U16155 (N_16155,N_15713,N_15987);
nand U16156 (N_16156,N_15974,N_15991);
or U16157 (N_16157,N_15752,N_15970);
and U16158 (N_16158,N_15653,N_15939);
and U16159 (N_16159,N_15507,N_15624);
nor U16160 (N_16160,N_15894,N_15546);
nand U16161 (N_16161,N_15904,N_15799);
and U16162 (N_16162,N_15940,N_15530);
nor U16163 (N_16163,N_15935,N_15562);
or U16164 (N_16164,N_15754,N_15636);
and U16165 (N_16165,N_15705,N_15794);
or U16166 (N_16166,N_15522,N_15840);
nand U16167 (N_16167,N_15808,N_15949);
and U16168 (N_16168,N_15592,N_15678);
nand U16169 (N_16169,N_15509,N_15930);
nor U16170 (N_16170,N_15612,N_15648);
nand U16171 (N_16171,N_15852,N_15899);
nand U16172 (N_16172,N_15876,N_15719);
nor U16173 (N_16173,N_15733,N_15580);
xnor U16174 (N_16174,N_15574,N_15738);
nand U16175 (N_16175,N_15881,N_15666);
nor U16176 (N_16176,N_15504,N_15576);
and U16177 (N_16177,N_15720,N_15563);
and U16178 (N_16178,N_15955,N_15924);
nor U16179 (N_16179,N_15516,N_15608);
nor U16180 (N_16180,N_15746,N_15845);
xor U16181 (N_16181,N_15693,N_15976);
and U16182 (N_16182,N_15878,N_15838);
or U16183 (N_16183,N_15777,N_15966);
xnor U16184 (N_16184,N_15938,N_15699);
and U16185 (N_16185,N_15782,N_15770);
nor U16186 (N_16186,N_15885,N_15968);
or U16187 (N_16187,N_15957,N_15521);
and U16188 (N_16188,N_15821,N_15853);
and U16189 (N_16189,N_15567,N_15637);
nor U16190 (N_16190,N_15879,N_15570);
or U16191 (N_16191,N_15905,N_15583);
nor U16192 (N_16192,N_15554,N_15629);
xnor U16193 (N_16193,N_15692,N_15800);
and U16194 (N_16194,N_15934,N_15761);
nand U16195 (N_16195,N_15750,N_15614);
xnor U16196 (N_16196,N_15723,N_15783);
or U16197 (N_16197,N_15890,N_15978);
or U16198 (N_16198,N_15822,N_15841);
nand U16199 (N_16199,N_15985,N_15888);
nand U16200 (N_16200,N_15954,N_15695);
nor U16201 (N_16201,N_15544,N_15520);
or U16202 (N_16202,N_15965,N_15756);
nand U16203 (N_16203,N_15891,N_15525);
and U16204 (N_16204,N_15953,N_15873);
xor U16205 (N_16205,N_15682,N_15871);
and U16206 (N_16206,N_15518,N_15944);
or U16207 (N_16207,N_15839,N_15634);
or U16208 (N_16208,N_15523,N_15811);
xor U16209 (N_16209,N_15909,N_15735);
nand U16210 (N_16210,N_15711,N_15919);
xnor U16211 (N_16211,N_15848,N_15559);
nor U16212 (N_16212,N_15925,N_15718);
nor U16213 (N_16213,N_15776,N_15790);
and U16214 (N_16214,N_15667,N_15932);
nor U16215 (N_16215,N_15500,N_15610);
nand U16216 (N_16216,N_15931,N_15766);
nand U16217 (N_16217,N_15657,N_15568);
and U16218 (N_16218,N_15694,N_15895);
and U16219 (N_16219,N_15980,N_15627);
and U16220 (N_16220,N_15806,N_15760);
nor U16221 (N_16221,N_15528,N_15952);
nor U16222 (N_16222,N_15573,N_15767);
and U16223 (N_16223,N_15946,N_15850);
nand U16224 (N_16224,N_15900,N_15896);
nor U16225 (N_16225,N_15728,N_15644);
or U16226 (N_16226,N_15584,N_15933);
or U16227 (N_16227,N_15908,N_15595);
nand U16228 (N_16228,N_15773,N_15585);
xor U16229 (N_16229,N_15804,N_15588);
or U16230 (N_16230,N_15731,N_15542);
xnor U16231 (N_16231,N_15942,N_15722);
nor U16232 (N_16232,N_15691,N_15606);
or U16233 (N_16233,N_15762,N_15683);
nor U16234 (N_16234,N_15658,N_15945);
nor U16235 (N_16235,N_15915,N_15753);
nor U16236 (N_16236,N_15721,N_15956);
xor U16237 (N_16237,N_15565,N_15837);
and U16238 (N_16238,N_15810,N_15662);
or U16239 (N_16239,N_15708,N_15613);
xnor U16240 (N_16240,N_15703,N_15941);
nor U16241 (N_16241,N_15686,N_15593);
xnor U16242 (N_16242,N_15868,N_15649);
nor U16243 (N_16243,N_15922,N_15659);
nand U16244 (N_16244,N_15540,N_15524);
or U16245 (N_16245,N_15743,N_15616);
or U16246 (N_16246,N_15823,N_15825);
and U16247 (N_16247,N_15969,N_15620);
and U16248 (N_16248,N_15589,N_15527);
xnor U16249 (N_16249,N_15857,N_15865);
and U16250 (N_16250,N_15743,N_15796);
nand U16251 (N_16251,N_15667,N_15596);
xnor U16252 (N_16252,N_15946,N_15649);
nor U16253 (N_16253,N_15849,N_15881);
nand U16254 (N_16254,N_15637,N_15650);
or U16255 (N_16255,N_15966,N_15961);
and U16256 (N_16256,N_15814,N_15899);
nor U16257 (N_16257,N_15517,N_15614);
and U16258 (N_16258,N_15796,N_15839);
and U16259 (N_16259,N_15776,N_15575);
or U16260 (N_16260,N_15534,N_15719);
nor U16261 (N_16261,N_15962,N_15951);
or U16262 (N_16262,N_15780,N_15751);
nor U16263 (N_16263,N_15699,N_15713);
and U16264 (N_16264,N_15769,N_15616);
nand U16265 (N_16265,N_15814,N_15750);
and U16266 (N_16266,N_15651,N_15667);
xnor U16267 (N_16267,N_15887,N_15906);
nor U16268 (N_16268,N_15555,N_15787);
xnor U16269 (N_16269,N_15771,N_15815);
or U16270 (N_16270,N_15651,N_15746);
xor U16271 (N_16271,N_15781,N_15891);
nor U16272 (N_16272,N_15885,N_15987);
and U16273 (N_16273,N_15958,N_15849);
xor U16274 (N_16274,N_15964,N_15769);
nand U16275 (N_16275,N_15589,N_15620);
nor U16276 (N_16276,N_15707,N_15831);
nor U16277 (N_16277,N_15986,N_15660);
and U16278 (N_16278,N_15930,N_15640);
nand U16279 (N_16279,N_15679,N_15575);
or U16280 (N_16280,N_15990,N_15542);
nor U16281 (N_16281,N_15774,N_15769);
xor U16282 (N_16282,N_15664,N_15526);
nor U16283 (N_16283,N_15800,N_15888);
nand U16284 (N_16284,N_15647,N_15896);
and U16285 (N_16285,N_15733,N_15979);
or U16286 (N_16286,N_15994,N_15788);
xor U16287 (N_16287,N_15513,N_15937);
and U16288 (N_16288,N_15548,N_15933);
nand U16289 (N_16289,N_15502,N_15954);
nand U16290 (N_16290,N_15576,N_15620);
xor U16291 (N_16291,N_15535,N_15848);
nor U16292 (N_16292,N_15514,N_15648);
nand U16293 (N_16293,N_15872,N_15625);
nand U16294 (N_16294,N_15569,N_15955);
xnor U16295 (N_16295,N_15878,N_15716);
xor U16296 (N_16296,N_15572,N_15685);
nor U16297 (N_16297,N_15524,N_15857);
nor U16298 (N_16298,N_15692,N_15866);
or U16299 (N_16299,N_15666,N_15701);
or U16300 (N_16300,N_15519,N_15796);
and U16301 (N_16301,N_15663,N_15802);
nand U16302 (N_16302,N_15664,N_15747);
nand U16303 (N_16303,N_15867,N_15918);
nand U16304 (N_16304,N_15811,N_15857);
nand U16305 (N_16305,N_15809,N_15511);
and U16306 (N_16306,N_15652,N_15726);
nand U16307 (N_16307,N_15786,N_15628);
nor U16308 (N_16308,N_15539,N_15859);
and U16309 (N_16309,N_15752,N_15555);
xor U16310 (N_16310,N_15580,N_15941);
and U16311 (N_16311,N_15665,N_15981);
and U16312 (N_16312,N_15734,N_15953);
nor U16313 (N_16313,N_15949,N_15541);
nor U16314 (N_16314,N_15870,N_15876);
and U16315 (N_16315,N_15751,N_15595);
xor U16316 (N_16316,N_15505,N_15879);
nor U16317 (N_16317,N_15862,N_15735);
nor U16318 (N_16318,N_15550,N_15935);
or U16319 (N_16319,N_15981,N_15967);
nor U16320 (N_16320,N_15971,N_15709);
or U16321 (N_16321,N_15545,N_15893);
and U16322 (N_16322,N_15625,N_15701);
or U16323 (N_16323,N_15678,N_15662);
nor U16324 (N_16324,N_15572,N_15844);
and U16325 (N_16325,N_15794,N_15950);
or U16326 (N_16326,N_15555,N_15633);
and U16327 (N_16327,N_15616,N_15992);
nor U16328 (N_16328,N_15963,N_15796);
or U16329 (N_16329,N_15541,N_15708);
nand U16330 (N_16330,N_15990,N_15815);
and U16331 (N_16331,N_15509,N_15924);
and U16332 (N_16332,N_15868,N_15862);
or U16333 (N_16333,N_15516,N_15989);
and U16334 (N_16334,N_15944,N_15719);
xnor U16335 (N_16335,N_15946,N_15762);
and U16336 (N_16336,N_15771,N_15802);
or U16337 (N_16337,N_15963,N_15635);
and U16338 (N_16338,N_15820,N_15935);
xor U16339 (N_16339,N_15615,N_15667);
or U16340 (N_16340,N_15568,N_15729);
or U16341 (N_16341,N_15502,N_15949);
nor U16342 (N_16342,N_15793,N_15761);
nand U16343 (N_16343,N_15772,N_15587);
nor U16344 (N_16344,N_15956,N_15799);
nand U16345 (N_16345,N_15871,N_15556);
nor U16346 (N_16346,N_15918,N_15621);
nor U16347 (N_16347,N_15894,N_15830);
and U16348 (N_16348,N_15909,N_15636);
or U16349 (N_16349,N_15734,N_15652);
or U16350 (N_16350,N_15796,N_15585);
nand U16351 (N_16351,N_15910,N_15880);
xor U16352 (N_16352,N_15860,N_15949);
or U16353 (N_16353,N_15507,N_15929);
xnor U16354 (N_16354,N_15926,N_15641);
nor U16355 (N_16355,N_15706,N_15835);
and U16356 (N_16356,N_15505,N_15983);
or U16357 (N_16357,N_15502,N_15841);
nand U16358 (N_16358,N_15969,N_15672);
or U16359 (N_16359,N_15591,N_15710);
and U16360 (N_16360,N_15754,N_15776);
and U16361 (N_16361,N_15564,N_15900);
nand U16362 (N_16362,N_15663,N_15506);
or U16363 (N_16363,N_15632,N_15564);
nand U16364 (N_16364,N_15776,N_15802);
and U16365 (N_16365,N_15897,N_15609);
and U16366 (N_16366,N_15957,N_15855);
nor U16367 (N_16367,N_15583,N_15553);
and U16368 (N_16368,N_15964,N_15574);
and U16369 (N_16369,N_15518,N_15896);
and U16370 (N_16370,N_15728,N_15870);
nor U16371 (N_16371,N_15703,N_15919);
or U16372 (N_16372,N_15508,N_15805);
nor U16373 (N_16373,N_15598,N_15628);
or U16374 (N_16374,N_15951,N_15944);
nand U16375 (N_16375,N_15509,N_15627);
nand U16376 (N_16376,N_15676,N_15511);
nor U16377 (N_16377,N_15665,N_15856);
xor U16378 (N_16378,N_15795,N_15827);
and U16379 (N_16379,N_15998,N_15695);
xor U16380 (N_16380,N_15891,N_15945);
nor U16381 (N_16381,N_15648,N_15917);
nand U16382 (N_16382,N_15966,N_15676);
and U16383 (N_16383,N_15647,N_15667);
or U16384 (N_16384,N_15853,N_15538);
xor U16385 (N_16385,N_15648,N_15810);
and U16386 (N_16386,N_15581,N_15745);
nand U16387 (N_16387,N_15877,N_15974);
and U16388 (N_16388,N_15875,N_15716);
xnor U16389 (N_16389,N_15624,N_15656);
nand U16390 (N_16390,N_15564,N_15526);
nor U16391 (N_16391,N_15902,N_15790);
nor U16392 (N_16392,N_15936,N_15731);
nor U16393 (N_16393,N_15633,N_15944);
and U16394 (N_16394,N_15678,N_15706);
and U16395 (N_16395,N_15685,N_15765);
nand U16396 (N_16396,N_15619,N_15824);
nand U16397 (N_16397,N_15742,N_15646);
nand U16398 (N_16398,N_15620,N_15839);
and U16399 (N_16399,N_15797,N_15821);
nand U16400 (N_16400,N_15994,N_15583);
nor U16401 (N_16401,N_15741,N_15854);
or U16402 (N_16402,N_15994,N_15948);
or U16403 (N_16403,N_15849,N_15698);
or U16404 (N_16404,N_15653,N_15969);
nor U16405 (N_16405,N_15560,N_15638);
nor U16406 (N_16406,N_15583,N_15719);
and U16407 (N_16407,N_15937,N_15913);
nor U16408 (N_16408,N_15555,N_15552);
and U16409 (N_16409,N_15577,N_15784);
nand U16410 (N_16410,N_15747,N_15833);
or U16411 (N_16411,N_15593,N_15671);
and U16412 (N_16412,N_15930,N_15794);
nor U16413 (N_16413,N_15630,N_15980);
or U16414 (N_16414,N_15703,N_15552);
or U16415 (N_16415,N_15738,N_15905);
nor U16416 (N_16416,N_15599,N_15527);
nand U16417 (N_16417,N_15771,N_15616);
or U16418 (N_16418,N_15910,N_15737);
xnor U16419 (N_16419,N_15916,N_15860);
and U16420 (N_16420,N_15748,N_15741);
and U16421 (N_16421,N_15785,N_15640);
or U16422 (N_16422,N_15838,N_15526);
nor U16423 (N_16423,N_15629,N_15617);
nor U16424 (N_16424,N_15975,N_15886);
nor U16425 (N_16425,N_15611,N_15520);
or U16426 (N_16426,N_15854,N_15864);
and U16427 (N_16427,N_15500,N_15623);
and U16428 (N_16428,N_15586,N_15523);
nor U16429 (N_16429,N_15870,N_15679);
and U16430 (N_16430,N_15803,N_15850);
nor U16431 (N_16431,N_15517,N_15748);
xnor U16432 (N_16432,N_15575,N_15806);
and U16433 (N_16433,N_15656,N_15546);
nor U16434 (N_16434,N_15719,N_15546);
nand U16435 (N_16435,N_15517,N_15950);
nor U16436 (N_16436,N_15529,N_15799);
nand U16437 (N_16437,N_15601,N_15653);
xor U16438 (N_16438,N_15931,N_15663);
nand U16439 (N_16439,N_15668,N_15648);
or U16440 (N_16440,N_15528,N_15857);
nand U16441 (N_16441,N_15670,N_15543);
nor U16442 (N_16442,N_15943,N_15962);
and U16443 (N_16443,N_15794,N_15810);
nand U16444 (N_16444,N_15898,N_15749);
nor U16445 (N_16445,N_15959,N_15960);
nor U16446 (N_16446,N_15541,N_15656);
and U16447 (N_16447,N_15841,N_15546);
nand U16448 (N_16448,N_15708,N_15980);
nor U16449 (N_16449,N_15599,N_15792);
or U16450 (N_16450,N_15941,N_15573);
nand U16451 (N_16451,N_15904,N_15647);
and U16452 (N_16452,N_15801,N_15816);
nor U16453 (N_16453,N_15544,N_15542);
nor U16454 (N_16454,N_15522,N_15560);
nor U16455 (N_16455,N_15979,N_15829);
and U16456 (N_16456,N_15720,N_15759);
and U16457 (N_16457,N_15864,N_15535);
nor U16458 (N_16458,N_15729,N_15826);
or U16459 (N_16459,N_15549,N_15614);
and U16460 (N_16460,N_15775,N_15898);
nor U16461 (N_16461,N_15895,N_15738);
and U16462 (N_16462,N_15516,N_15868);
nand U16463 (N_16463,N_15935,N_15882);
and U16464 (N_16464,N_15725,N_15899);
nand U16465 (N_16465,N_15501,N_15649);
nor U16466 (N_16466,N_15895,N_15522);
xnor U16467 (N_16467,N_15847,N_15558);
or U16468 (N_16468,N_15869,N_15637);
nor U16469 (N_16469,N_15750,N_15916);
nor U16470 (N_16470,N_15518,N_15619);
xnor U16471 (N_16471,N_15811,N_15797);
xor U16472 (N_16472,N_15586,N_15761);
nor U16473 (N_16473,N_15901,N_15978);
nand U16474 (N_16474,N_15607,N_15856);
nor U16475 (N_16475,N_15820,N_15814);
nand U16476 (N_16476,N_15865,N_15807);
and U16477 (N_16477,N_15899,N_15885);
and U16478 (N_16478,N_15794,N_15718);
nand U16479 (N_16479,N_15792,N_15700);
nand U16480 (N_16480,N_15521,N_15955);
nor U16481 (N_16481,N_15897,N_15956);
and U16482 (N_16482,N_15654,N_15946);
nand U16483 (N_16483,N_15823,N_15697);
nor U16484 (N_16484,N_15719,N_15618);
nor U16485 (N_16485,N_15839,N_15880);
or U16486 (N_16486,N_15988,N_15904);
and U16487 (N_16487,N_15607,N_15776);
xor U16488 (N_16488,N_15752,N_15664);
nand U16489 (N_16489,N_15966,N_15553);
and U16490 (N_16490,N_15776,N_15642);
or U16491 (N_16491,N_15740,N_15507);
nand U16492 (N_16492,N_15588,N_15992);
or U16493 (N_16493,N_15654,N_15593);
and U16494 (N_16494,N_15586,N_15577);
nand U16495 (N_16495,N_15569,N_15603);
nor U16496 (N_16496,N_15520,N_15523);
nor U16497 (N_16497,N_15596,N_15519);
and U16498 (N_16498,N_15516,N_15567);
xnor U16499 (N_16499,N_15874,N_15932);
or U16500 (N_16500,N_16361,N_16349);
nor U16501 (N_16501,N_16156,N_16254);
nand U16502 (N_16502,N_16238,N_16046);
nor U16503 (N_16503,N_16108,N_16200);
nand U16504 (N_16504,N_16430,N_16436);
nor U16505 (N_16505,N_16373,N_16129);
or U16506 (N_16506,N_16490,N_16325);
nand U16507 (N_16507,N_16179,N_16287);
xor U16508 (N_16508,N_16012,N_16122);
or U16509 (N_16509,N_16149,N_16450);
and U16510 (N_16510,N_16198,N_16441);
nand U16511 (N_16511,N_16498,N_16398);
or U16512 (N_16512,N_16479,N_16295);
or U16513 (N_16513,N_16334,N_16404);
nor U16514 (N_16514,N_16084,N_16275);
and U16515 (N_16515,N_16085,N_16352);
or U16516 (N_16516,N_16312,N_16458);
or U16517 (N_16517,N_16071,N_16069);
nand U16518 (N_16518,N_16204,N_16185);
and U16519 (N_16519,N_16375,N_16004);
nand U16520 (N_16520,N_16453,N_16386);
nand U16521 (N_16521,N_16078,N_16030);
and U16522 (N_16522,N_16270,N_16428);
nor U16523 (N_16523,N_16273,N_16460);
or U16524 (N_16524,N_16035,N_16292);
nand U16525 (N_16525,N_16408,N_16443);
nand U16526 (N_16526,N_16143,N_16043);
nor U16527 (N_16527,N_16187,N_16444);
nor U16528 (N_16528,N_16029,N_16212);
and U16529 (N_16529,N_16387,N_16374);
xor U16530 (N_16530,N_16128,N_16332);
or U16531 (N_16531,N_16065,N_16094);
and U16532 (N_16532,N_16345,N_16484);
or U16533 (N_16533,N_16383,N_16159);
nor U16534 (N_16534,N_16233,N_16305);
or U16535 (N_16535,N_16499,N_16471);
or U16536 (N_16536,N_16378,N_16298);
and U16537 (N_16537,N_16344,N_16465);
nor U16538 (N_16538,N_16054,N_16291);
nor U16539 (N_16539,N_16322,N_16337);
or U16540 (N_16540,N_16017,N_16231);
nand U16541 (N_16541,N_16440,N_16262);
xnor U16542 (N_16542,N_16308,N_16303);
or U16543 (N_16543,N_16388,N_16381);
or U16544 (N_16544,N_16124,N_16183);
or U16545 (N_16545,N_16409,N_16492);
xnor U16546 (N_16546,N_16496,N_16193);
xnor U16547 (N_16547,N_16488,N_16468);
xnor U16548 (N_16548,N_16152,N_16057);
or U16549 (N_16549,N_16144,N_16497);
and U16550 (N_16550,N_16219,N_16127);
and U16551 (N_16551,N_16354,N_16318);
nand U16552 (N_16552,N_16396,N_16363);
and U16553 (N_16553,N_16105,N_16220);
nor U16554 (N_16554,N_16058,N_16269);
or U16555 (N_16555,N_16136,N_16358);
nand U16556 (N_16556,N_16203,N_16037);
or U16557 (N_16557,N_16131,N_16045);
and U16558 (N_16558,N_16245,N_16316);
xor U16559 (N_16559,N_16125,N_16210);
nand U16560 (N_16560,N_16264,N_16080);
xnor U16561 (N_16561,N_16376,N_16330);
and U16562 (N_16562,N_16118,N_16424);
and U16563 (N_16563,N_16423,N_16459);
nor U16564 (N_16564,N_16306,N_16066);
and U16565 (N_16565,N_16215,N_16456);
nand U16566 (N_16566,N_16402,N_16008);
xnor U16567 (N_16567,N_16195,N_16117);
and U16568 (N_16568,N_16031,N_16184);
nand U16569 (N_16569,N_16181,N_16082);
and U16570 (N_16570,N_16447,N_16163);
nor U16571 (N_16571,N_16324,N_16164);
and U16572 (N_16572,N_16432,N_16229);
or U16573 (N_16573,N_16250,N_16106);
nor U16574 (N_16574,N_16205,N_16107);
and U16575 (N_16575,N_16469,N_16294);
nor U16576 (N_16576,N_16293,N_16304);
nor U16577 (N_16577,N_16491,N_16445);
nand U16578 (N_16578,N_16257,N_16024);
and U16579 (N_16579,N_16281,N_16434);
nor U16580 (N_16580,N_16135,N_16138);
nor U16581 (N_16581,N_16145,N_16414);
nor U16582 (N_16582,N_16147,N_16323);
nor U16583 (N_16583,N_16253,N_16272);
or U16584 (N_16584,N_16333,N_16000);
xor U16585 (N_16585,N_16161,N_16222);
and U16586 (N_16586,N_16360,N_16486);
nand U16587 (N_16587,N_16403,N_16463);
and U16588 (N_16588,N_16148,N_16422);
nor U16589 (N_16589,N_16277,N_16236);
and U16590 (N_16590,N_16096,N_16346);
nor U16591 (N_16591,N_16480,N_16327);
or U16592 (N_16592,N_16002,N_16251);
nand U16593 (N_16593,N_16049,N_16418);
nand U16594 (N_16594,N_16494,N_16232);
nor U16595 (N_16595,N_16064,N_16177);
nand U16596 (N_16596,N_16213,N_16466);
nor U16597 (N_16597,N_16151,N_16188);
or U16598 (N_16598,N_16223,N_16495);
nor U16599 (N_16599,N_16086,N_16347);
or U16600 (N_16600,N_16299,N_16001);
xor U16601 (N_16601,N_16199,N_16100);
xnor U16602 (N_16602,N_16025,N_16070);
nor U16603 (N_16603,N_16095,N_16393);
and U16604 (N_16604,N_16237,N_16015);
nand U16605 (N_16605,N_16371,N_16252);
or U16606 (N_16606,N_16493,N_16379);
nand U16607 (N_16607,N_16289,N_16112);
or U16608 (N_16608,N_16353,N_16052);
or U16609 (N_16609,N_16313,N_16470);
or U16610 (N_16610,N_16258,N_16178);
nor U16611 (N_16611,N_16259,N_16307);
nor U16612 (N_16612,N_16076,N_16014);
nor U16613 (N_16613,N_16315,N_16317);
and U16614 (N_16614,N_16048,N_16420);
and U16615 (N_16615,N_16462,N_16176);
nand U16616 (N_16616,N_16266,N_16362);
nand U16617 (N_16617,N_16477,N_16101);
xnor U16618 (N_16618,N_16067,N_16074);
nor U16619 (N_16619,N_16090,N_16310);
nand U16620 (N_16620,N_16335,N_16256);
nor U16621 (N_16621,N_16399,N_16032);
or U16622 (N_16622,N_16126,N_16435);
or U16623 (N_16623,N_16239,N_16454);
nor U16624 (N_16624,N_16206,N_16150);
and U16625 (N_16625,N_16201,N_16230);
or U16626 (N_16626,N_16091,N_16120);
or U16627 (N_16627,N_16429,N_16370);
and U16628 (N_16628,N_16023,N_16365);
nand U16629 (N_16629,N_16320,N_16225);
nand U16630 (N_16630,N_16140,N_16167);
and U16631 (N_16631,N_16234,N_16007);
xor U16632 (N_16632,N_16467,N_16134);
nor U16633 (N_16633,N_16060,N_16482);
or U16634 (N_16634,N_16075,N_16242);
and U16635 (N_16635,N_16036,N_16366);
and U16636 (N_16636,N_16226,N_16413);
or U16637 (N_16637,N_16350,N_16359);
nor U16638 (N_16638,N_16146,N_16377);
and U16639 (N_16639,N_16214,N_16157);
and U16640 (N_16640,N_16174,N_16412);
xnor U16641 (N_16641,N_16415,N_16392);
nand U16642 (N_16642,N_16355,N_16077);
nor U16643 (N_16643,N_16050,N_16020);
nand U16644 (N_16644,N_16166,N_16472);
and U16645 (N_16645,N_16265,N_16191);
nand U16646 (N_16646,N_16040,N_16218);
xor U16647 (N_16647,N_16489,N_16426);
nand U16648 (N_16648,N_16416,N_16087);
nand U16649 (N_16649,N_16243,N_16019);
and U16650 (N_16650,N_16457,N_16142);
nor U16651 (N_16651,N_16110,N_16247);
or U16652 (N_16652,N_16442,N_16263);
or U16653 (N_16653,N_16286,N_16338);
and U16654 (N_16654,N_16451,N_16194);
and U16655 (N_16655,N_16246,N_16133);
nand U16656 (N_16656,N_16068,N_16329);
or U16657 (N_16657,N_16439,N_16385);
nand U16658 (N_16658,N_16227,N_16328);
nand U16659 (N_16659,N_16154,N_16475);
xnor U16660 (N_16660,N_16059,N_16321);
or U16661 (N_16661,N_16417,N_16170);
or U16662 (N_16662,N_16348,N_16446);
or U16663 (N_16663,N_16190,N_16153);
and U16664 (N_16664,N_16208,N_16209);
nor U16665 (N_16665,N_16400,N_16056);
xor U16666 (N_16666,N_16182,N_16102);
xnor U16667 (N_16667,N_16063,N_16421);
and U16668 (N_16668,N_16003,N_16088);
and U16669 (N_16669,N_16038,N_16285);
nor U16670 (N_16670,N_16217,N_16476);
nand U16671 (N_16671,N_16072,N_16260);
nand U16672 (N_16672,N_16478,N_16397);
nand U16673 (N_16673,N_16041,N_16016);
or U16674 (N_16674,N_16175,N_16005);
nand U16675 (N_16675,N_16311,N_16437);
and U16676 (N_16676,N_16314,N_16279);
nor U16677 (N_16677,N_16033,N_16158);
or U16678 (N_16678,N_16039,N_16121);
or U16679 (N_16679,N_16274,N_16389);
nor U16680 (N_16680,N_16172,N_16483);
and U16681 (N_16681,N_16301,N_16160);
and U16682 (N_16682,N_16255,N_16427);
nand U16683 (N_16683,N_16228,N_16180);
or U16684 (N_16684,N_16047,N_16391);
nand U16685 (N_16685,N_16006,N_16367);
and U16686 (N_16686,N_16013,N_16197);
and U16687 (N_16687,N_16487,N_16173);
nand U16688 (N_16688,N_16109,N_16248);
nor U16689 (N_16689,N_16189,N_16368);
nor U16690 (N_16690,N_16425,N_16132);
and U16691 (N_16691,N_16485,N_16419);
xor U16692 (N_16692,N_16452,N_16081);
nand U16693 (N_16693,N_16438,N_16051);
xnor U16694 (N_16694,N_16202,N_16342);
nor U16695 (N_16695,N_16042,N_16319);
and U16696 (N_16696,N_16116,N_16244);
and U16697 (N_16697,N_16114,N_16284);
or U16698 (N_16698,N_16027,N_16062);
nor U16699 (N_16699,N_16384,N_16382);
nor U16700 (N_16700,N_16390,N_16267);
or U16701 (N_16701,N_16331,N_16162);
xor U16702 (N_16702,N_16302,N_16288);
nor U16703 (N_16703,N_16123,N_16290);
or U16704 (N_16704,N_16249,N_16364);
or U16705 (N_16705,N_16103,N_16448);
and U16706 (N_16706,N_16073,N_16407);
or U16707 (N_16707,N_16224,N_16473);
nor U16708 (N_16708,N_16211,N_16336);
nand U16709 (N_16709,N_16079,N_16139);
and U16710 (N_16710,N_16431,N_16296);
or U16711 (N_16711,N_16028,N_16235);
or U16712 (N_16712,N_16241,N_16169);
nor U16713 (N_16713,N_16406,N_16034);
or U16714 (N_16714,N_16021,N_16083);
nand U16715 (N_16715,N_16221,N_16089);
nor U16716 (N_16716,N_16411,N_16009);
nand U16717 (N_16717,N_16401,N_16481);
and U16718 (N_16718,N_16341,N_16092);
nor U16719 (N_16719,N_16171,N_16395);
and U16720 (N_16720,N_16111,N_16297);
nor U16721 (N_16721,N_16168,N_16155);
and U16722 (N_16722,N_16280,N_16394);
xor U16723 (N_16723,N_16119,N_16449);
nor U16724 (N_16724,N_16115,N_16278);
nor U16725 (N_16725,N_16011,N_16268);
nand U16726 (N_16726,N_16018,N_16369);
xnor U16727 (N_16727,N_16271,N_16104);
nand U16728 (N_16728,N_16455,N_16061);
xnor U16729 (N_16729,N_16405,N_16340);
nor U16730 (N_16730,N_16165,N_16461);
and U16731 (N_16731,N_16357,N_16309);
or U16732 (N_16732,N_16216,N_16196);
nand U16733 (N_16733,N_16380,N_16026);
xnor U16734 (N_16734,N_16130,N_16351);
nand U16735 (N_16735,N_16113,N_16240);
and U16736 (N_16736,N_16276,N_16326);
xor U16737 (N_16737,N_16474,N_16433);
nand U16738 (N_16738,N_16339,N_16099);
nand U16739 (N_16739,N_16098,N_16186);
and U16740 (N_16740,N_16053,N_16282);
and U16741 (N_16741,N_16343,N_16300);
and U16742 (N_16742,N_16261,N_16044);
and U16743 (N_16743,N_16192,N_16010);
and U16744 (N_16744,N_16464,N_16207);
or U16745 (N_16745,N_16097,N_16283);
and U16746 (N_16746,N_16410,N_16356);
or U16747 (N_16747,N_16022,N_16141);
nand U16748 (N_16748,N_16372,N_16093);
nor U16749 (N_16749,N_16055,N_16137);
or U16750 (N_16750,N_16091,N_16469);
nor U16751 (N_16751,N_16284,N_16182);
nand U16752 (N_16752,N_16389,N_16103);
or U16753 (N_16753,N_16209,N_16380);
nor U16754 (N_16754,N_16173,N_16293);
or U16755 (N_16755,N_16300,N_16290);
and U16756 (N_16756,N_16345,N_16265);
and U16757 (N_16757,N_16161,N_16443);
and U16758 (N_16758,N_16414,N_16241);
or U16759 (N_16759,N_16220,N_16372);
nor U16760 (N_16760,N_16154,N_16353);
nor U16761 (N_16761,N_16250,N_16472);
or U16762 (N_16762,N_16335,N_16061);
nand U16763 (N_16763,N_16457,N_16106);
or U16764 (N_16764,N_16476,N_16112);
nor U16765 (N_16765,N_16179,N_16345);
or U16766 (N_16766,N_16478,N_16451);
nand U16767 (N_16767,N_16209,N_16367);
nor U16768 (N_16768,N_16470,N_16100);
and U16769 (N_16769,N_16043,N_16034);
nand U16770 (N_16770,N_16312,N_16022);
nor U16771 (N_16771,N_16111,N_16084);
nor U16772 (N_16772,N_16200,N_16252);
nand U16773 (N_16773,N_16348,N_16164);
nor U16774 (N_16774,N_16480,N_16264);
nor U16775 (N_16775,N_16218,N_16025);
xnor U16776 (N_16776,N_16351,N_16435);
or U16777 (N_16777,N_16021,N_16133);
or U16778 (N_16778,N_16230,N_16216);
and U16779 (N_16779,N_16466,N_16037);
or U16780 (N_16780,N_16060,N_16439);
and U16781 (N_16781,N_16432,N_16078);
nand U16782 (N_16782,N_16195,N_16431);
or U16783 (N_16783,N_16004,N_16114);
and U16784 (N_16784,N_16005,N_16296);
xor U16785 (N_16785,N_16150,N_16182);
xnor U16786 (N_16786,N_16050,N_16026);
or U16787 (N_16787,N_16040,N_16108);
and U16788 (N_16788,N_16096,N_16495);
nor U16789 (N_16789,N_16050,N_16209);
and U16790 (N_16790,N_16091,N_16355);
nand U16791 (N_16791,N_16423,N_16210);
and U16792 (N_16792,N_16020,N_16492);
nand U16793 (N_16793,N_16390,N_16421);
and U16794 (N_16794,N_16356,N_16480);
nand U16795 (N_16795,N_16385,N_16045);
or U16796 (N_16796,N_16020,N_16450);
nand U16797 (N_16797,N_16384,N_16448);
nand U16798 (N_16798,N_16364,N_16346);
and U16799 (N_16799,N_16176,N_16374);
and U16800 (N_16800,N_16402,N_16496);
nor U16801 (N_16801,N_16385,N_16323);
nand U16802 (N_16802,N_16088,N_16480);
or U16803 (N_16803,N_16001,N_16167);
and U16804 (N_16804,N_16462,N_16037);
xnor U16805 (N_16805,N_16472,N_16174);
nor U16806 (N_16806,N_16193,N_16404);
and U16807 (N_16807,N_16015,N_16170);
nand U16808 (N_16808,N_16128,N_16189);
nand U16809 (N_16809,N_16283,N_16355);
and U16810 (N_16810,N_16008,N_16104);
and U16811 (N_16811,N_16295,N_16366);
nor U16812 (N_16812,N_16094,N_16348);
and U16813 (N_16813,N_16340,N_16216);
nand U16814 (N_16814,N_16105,N_16333);
and U16815 (N_16815,N_16357,N_16336);
and U16816 (N_16816,N_16334,N_16463);
nor U16817 (N_16817,N_16134,N_16094);
nand U16818 (N_16818,N_16323,N_16133);
nor U16819 (N_16819,N_16234,N_16477);
and U16820 (N_16820,N_16478,N_16202);
or U16821 (N_16821,N_16159,N_16219);
and U16822 (N_16822,N_16424,N_16416);
nor U16823 (N_16823,N_16224,N_16423);
nand U16824 (N_16824,N_16272,N_16292);
nand U16825 (N_16825,N_16189,N_16305);
nor U16826 (N_16826,N_16090,N_16225);
nor U16827 (N_16827,N_16450,N_16308);
nand U16828 (N_16828,N_16055,N_16487);
or U16829 (N_16829,N_16193,N_16311);
xor U16830 (N_16830,N_16246,N_16030);
or U16831 (N_16831,N_16330,N_16249);
and U16832 (N_16832,N_16350,N_16152);
and U16833 (N_16833,N_16281,N_16064);
and U16834 (N_16834,N_16086,N_16445);
or U16835 (N_16835,N_16068,N_16022);
nand U16836 (N_16836,N_16054,N_16454);
xnor U16837 (N_16837,N_16184,N_16213);
or U16838 (N_16838,N_16086,N_16013);
and U16839 (N_16839,N_16351,N_16340);
nor U16840 (N_16840,N_16190,N_16267);
xnor U16841 (N_16841,N_16100,N_16037);
nor U16842 (N_16842,N_16110,N_16213);
or U16843 (N_16843,N_16250,N_16001);
xnor U16844 (N_16844,N_16166,N_16270);
and U16845 (N_16845,N_16451,N_16252);
or U16846 (N_16846,N_16284,N_16149);
xor U16847 (N_16847,N_16411,N_16123);
nor U16848 (N_16848,N_16418,N_16486);
nand U16849 (N_16849,N_16112,N_16279);
or U16850 (N_16850,N_16376,N_16049);
and U16851 (N_16851,N_16144,N_16130);
or U16852 (N_16852,N_16395,N_16253);
nor U16853 (N_16853,N_16044,N_16413);
or U16854 (N_16854,N_16439,N_16430);
or U16855 (N_16855,N_16374,N_16241);
nor U16856 (N_16856,N_16339,N_16429);
or U16857 (N_16857,N_16161,N_16006);
nor U16858 (N_16858,N_16458,N_16257);
nor U16859 (N_16859,N_16015,N_16406);
and U16860 (N_16860,N_16415,N_16153);
or U16861 (N_16861,N_16211,N_16236);
xnor U16862 (N_16862,N_16178,N_16158);
nor U16863 (N_16863,N_16284,N_16202);
nand U16864 (N_16864,N_16222,N_16466);
or U16865 (N_16865,N_16154,N_16021);
nand U16866 (N_16866,N_16038,N_16359);
and U16867 (N_16867,N_16002,N_16433);
nand U16868 (N_16868,N_16183,N_16268);
nand U16869 (N_16869,N_16102,N_16418);
xnor U16870 (N_16870,N_16120,N_16471);
and U16871 (N_16871,N_16092,N_16255);
and U16872 (N_16872,N_16308,N_16113);
or U16873 (N_16873,N_16124,N_16300);
nor U16874 (N_16874,N_16440,N_16240);
or U16875 (N_16875,N_16231,N_16489);
nor U16876 (N_16876,N_16076,N_16463);
and U16877 (N_16877,N_16191,N_16122);
nand U16878 (N_16878,N_16463,N_16089);
nand U16879 (N_16879,N_16016,N_16369);
nor U16880 (N_16880,N_16349,N_16383);
or U16881 (N_16881,N_16334,N_16035);
nor U16882 (N_16882,N_16161,N_16404);
or U16883 (N_16883,N_16423,N_16036);
nor U16884 (N_16884,N_16351,N_16287);
or U16885 (N_16885,N_16157,N_16112);
xor U16886 (N_16886,N_16344,N_16481);
or U16887 (N_16887,N_16236,N_16117);
and U16888 (N_16888,N_16257,N_16297);
nor U16889 (N_16889,N_16034,N_16324);
and U16890 (N_16890,N_16246,N_16470);
nor U16891 (N_16891,N_16367,N_16003);
nand U16892 (N_16892,N_16224,N_16383);
nor U16893 (N_16893,N_16333,N_16227);
or U16894 (N_16894,N_16072,N_16024);
and U16895 (N_16895,N_16160,N_16186);
or U16896 (N_16896,N_16388,N_16359);
and U16897 (N_16897,N_16287,N_16192);
nand U16898 (N_16898,N_16089,N_16169);
and U16899 (N_16899,N_16368,N_16474);
nor U16900 (N_16900,N_16157,N_16140);
xnor U16901 (N_16901,N_16285,N_16264);
nor U16902 (N_16902,N_16380,N_16227);
and U16903 (N_16903,N_16048,N_16262);
or U16904 (N_16904,N_16381,N_16193);
or U16905 (N_16905,N_16025,N_16360);
and U16906 (N_16906,N_16489,N_16187);
nor U16907 (N_16907,N_16323,N_16495);
nor U16908 (N_16908,N_16057,N_16035);
or U16909 (N_16909,N_16283,N_16192);
or U16910 (N_16910,N_16403,N_16279);
nor U16911 (N_16911,N_16088,N_16308);
nor U16912 (N_16912,N_16449,N_16208);
xnor U16913 (N_16913,N_16270,N_16305);
xor U16914 (N_16914,N_16215,N_16439);
and U16915 (N_16915,N_16308,N_16390);
nand U16916 (N_16916,N_16003,N_16267);
and U16917 (N_16917,N_16429,N_16226);
nor U16918 (N_16918,N_16304,N_16468);
nor U16919 (N_16919,N_16041,N_16464);
nand U16920 (N_16920,N_16075,N_16026);
nand U16921 (N_16921,N_16449,N_16267);
and U16922 (N_16922,N_16115,N_16441);
nand U16923 (N_16923,N_16063,N_16066);
or U16924 (N_16924,N_16012,N_16280);
and U16925 (N_16925,N_16123,N_16410);
xor U16926 (N_16926,N_16136,N_16150);
or U16927 (N_16927,N_16106,N_16013);
and U16928 (N_16928,N_16297,N_16230);
and U16929 (N_16929,N_16172,N_16247);
or U16930 (N_16930,N_16399,N_16174);
nor U16931 (N_16931,N_16079,N_16369);
and U16932 (N_16932,N_16092,N_16304);
nand U16933 (N_16933,N_16178,N_16031);
nor U16934 (N_16934,N_16308,N_16236);
or U16935 (N_16935,N_16333,N_16045);
or U16936 (N_16936,N_16105,N_16041);
nor U16937 (N_16937,N_16095,N_16236);
and U16938 (N_16938,N_16318,N_16282);
and U16939 (N_16939,N_16086,N_16071);
and U16940 (N_16940,N_16335,N_16270);
nor U16941 (N_16941,N_16495,N_16229);
nor U16942 (N_16942,N_16460,N_16318);
xnor U16943 (N_16943,N_16412,N_16277);
nand U16944 (N_16944,N_16198,N_16467);
or U16945 (N_16945,N_16434,N_16141);
and U16946 (N_16946,N_16433,N_16165);
nand U16947 (N_16947,N_16169,N_16449);
xor U16948 (N_16948,N_16488,N_16048);
nand U16949 (N_16949,N_16026,N_16177);
or U16950 (N_16950,N_16150,N_16219);
nor U16951 (N_16951,N_16162,N_16428);
and U16952 (N_16952,N_16107,N_16046);
nand U16953 (N_16953,N_16431,N_16102);
nand U16954 (N_16954,N_16423,N_16029);
nand U16955 (N_16955,N_16150,N_16147);
nand U16956 (N_16956,N_16326,N_16229);
or U16957 (N_16957,N_16344,N_16052);
nand U16958 (N_16958,N_16015,N_16342);
xnor U16959 (N_16959,N_16107,N_16133);
nor U16960 (N_16960,N_16259,N_16349);
xnor U16961 (N_16961,N_16311,N_16272);
nor U16962 (N_16962,N_16081,N_16067);
nand U16963 (N_16963,N_16154,N_16426);
and U16964 (N_16964,N_16378,N_16242);
and U16965 (N_16965,N_16117,N_16252);
nand U16966 (N_16966,N_16489,N_16163);
nor U16967 (N_16967,N_16352,N_16357);
or U16968 (N_16968,N_16381,N_16237);
nand U16969 (N_16969,N_16400,N_16449);
nand U16970 (N_16970,N_16172,N_16056);
and U16971 (N_16971,N_16036,N_16353);
or U16972 (N_16972,N_16407,N_16252);
nor U16973 (N_16973,N_16154,N_16255);
and U16974 (N_16974,N_16495,N_16082);
or U16975 (N_16975,N_16421,N_16296);
and U16976 (N_16976,N_16096,N_16113);
and U16977 (N_16977,N_16448,N_16263);
nand U16978 (N_16978,N_16250,N_16276);
and U16979 (N_16979,N_16221,N_16385);
nand U16980 (N_16980,N_16036,N_16336);
and U16981 (N_16981,N_16022,N_16408);
nor U16982 (N_16982,N_16396,N_16323);
nand U16983 (N_16983,N_16110,N_16317);
and U16984 (N_16984,N_16244,N_16282);
or U16985 (N_16985,N_16320,N_16423);
nand U16986 (N_16986,N_16036,N_16317);
or U16987 (N_16987,N_16046,N_16475);
and U16988 (N_16988,N_16482,N_16242);
or U16989 (N_16989,N_16451,N_16246);
nand U16990 (N_16990,N_16115,N_16411);
or U16991 (N_16991,N_16374,N_16147);
or U16992 (N_16992,N_16095,N_16185);
or U16993 (N_16993,N_16393,N_16260);
and U16994 (N_16994,N_16338,N_16112);
and U16995 (N_16995,N_16437,N_16219);
or U16996 (N_16996,N_16203,N_16485);
nand U16997 (N_16997,N_16084,N_16471);
and U16998 (N_16998,N_16326,N_16126);
and U16999 (N_16999,N_16015,N_16344);
and U17000 (N_17000,N_16574,N_16643);
nand U17001 (N_17001,N_16908,N_16992);
and U17002 (N_17002,N_16617,N_16584);
nor U17003 (N_17003,N_16951,N_16701);
or U17004 (N_17004,N_16579,N_16962);
and U17005 (N_17005,N_16652,N_16732);
xor U17006 (N_17006,N_16630,N_16664);
nor U17007 (N_17007,N_16957,N_16684);
and U17008 (N_17008,N_16720,N_16937);
xor U17009 (N_17009,N_16911,N_16677);
nand U17010 (N_17010,N_16641,N_16818);
nand U17011 (N_17011,N_16853,N_16946);
nor U17012 (N_17012,N_16873,N_16581);
nor U17013 (N_17013,N_16777,N_16921);
nor U17014 (N_17014,N_16578,N_16882);
and U17015 (N_17015,N_16721,N_16916);
xnor U17016 (N_17016,N_16835,N_16536);
xnor U17017 (N_17017,N_16567,N_16688);
nand U17018 (N_17018,N_16839,N_16788);
or U17019 (N_17019,N_16546,N_16909);
or U17020 (N_17020,N_16815,N_16650);
or U17021 (N_17021,N_16986,N_16770);
or U17022 (N_17022,N_16849,N_16583);
nor U17023 (N_17023,N_16504,N_16562);
nand U17024 (N_17024,N_16527,N_16586);
nand U17025 (N_17025,N_16859,N_16513);
nand U17026 (N_17026,N_16742,N_16978);
or U17027 (N_17027,N_16990,N_16791);
nand U17028 (N_17028,N_16865,N_16629);
nor U17029 (N_17029,N_16863,N_16890);
nor U17030 (N_17030,N_16825,N_16885);
nand U17031 (N_17031,N_16861,N_16717);
or U17032 (N_17032,N_16902,N_16556);
or U17033 (N_17033,N_16670,N_16539);
nor U17034 (N_17034,N_16712,N_16592);
nand U17035 (N_17035,N_16622,N_16699);
nor U17036 (N_17036,N_16797,N_16984);
and U17037 (N_17037,N_16858,N_16786);
or U17038 (N_17038,N_16662,N_16910);
or U17039 (N_17039,N_16893,N_16730);
xnor U17040 (N_17040,N_16750,N_16820);
nand U17041 (N_17041,N_16692,N_16700);
nand U17042 (N_17042,N_16549,N_16972);
xnor U17043 (N_17043,N_16781,N_16804);
and U17044 (N_17044,N_16837,N_16529);
and U17045 (N_17045,N_16522,N_16644);
nor U17046 (N_17046,N_16512,N_16794);
and U17047 (N_17047,N_16552,N_16526);
nor U17048 (N_17048,N_16875,N_16942);
or U17049 (N_17049,N_16572,N_16686);
nor U17050 (N_17050,N_16704,N_16758);
or U17051 (N_17051,N_16760,N_16649);
xor U17052 (N_17052,N_16570,N_16761);
nor U17053 (N_17053,N_16591,N_16842);
nor U17054 (N_17054,N_16678,N_16520);
xor U17055 (N_17055,N_16880,N_16614);
or U17056 (N_17056,N_16506,N_16599);
or U17057 (N_17057,N_16856,N_16999);
nor U17058 (N_17058,N_16975,N_16639);
or U17059 (N_17059,N_16889,N_16940);
nand U17060 (N_17060,N_16564,N_16703);
xor U17061 (N_17061,N_16654,N_16553);
nor U17062 (N_17062,N_16779,N_16737);
and U17063 (N_17063,N_16780,N_16667);
nand U17064 (N_17064,N_16618,N_16879);
nor U17065 (N_17065,N_16531,N_16941);
nor U17066 (N_17066,N_16577,N_16658);
and U17067 (N_17067,N_16901,N_16679);
nand U17068 (N_17068,N_16613,N_16636);
or U17069 (N_17069,N_16741,N_16870);
xor U17070 (N_17070,N_16881,N_16965);
or U17071 (N_17071,N_16759,N_16896);
nand U17072 (N_17072,N_16841,N_16573);
nand U17073 (N_17073,N_16651,N_16917);
nor U17074 (N_17074,N_16582,N_16855);
or U17075 (N_17075,N_16558,N_16868);
xnor U17076 (N_17076,N_16982,N_16607);
and U17077 (N_17077,N_16929,N_16874);
nor U17078 (N_17078,N_16866,N_16697);
nor U17079 (N_17079,N_16616,N_16799);
nand U17080 (N_17080,N_16603,N_16521);
nand U17081 (N_17081,N_16894,N_16631);
nor U17082 (N_17082,N_16734,N_16566);
or U17083 (N_17083,N_16598,N_16869);
nand U17084 (N_17084,N_16843,N_16587);
nor U17085 (N_17085,N_16805,N_16571);
xor U17086 (N_17086,N_16682,N_16695);
nand U17087 (N_17087,N_16974,N_16938);
and U17088 (N_17088,N_16718,N_16764);
xnor U17089 (N_17089,N_16936,N_16518);
xor U17090 (N_17090,N_16647,N_16877);
nor U17091 (N_17091,N_16500,N_16844);
nor U17092 (N_17092,N_16762,N_16983);
nor U17093 (N_17093,N_16906,N_16806);
and U17094 (N_17094,N_16748,N_16585);
nand U17095 (N_17095,N_16976,N_16733);
nand U17096 (N_17096,N_16511,N_16887);
nand U17097 (N_17097,N_16540,N_16959);
and U17098 (N_17098,N_16627,N_16969);
and U17099 (N_17099,N_16722,N_16826);
and U17100 (N_17100,N_16787,N_16538);
nand U17101 (N_17101,N_16600,N_16687);
or U17102 (N_17102,N_16832,N_16535);
and U17103 (N_17103,N_16604,N_16508);
nor U17104 (N_17104,N_16809,N_16694);
and U17105 (N_17105,N_16681,N_16862);
xnor U17106 (N_17106,N_16775,N_16778);
nor U17107 (N_17107,N_16763,N_16774);
nor U17108 (N_17108,N_16810,N_16743);
nor U17109 (N_17109,N_16950,N_16514);
or U17110 (N_17110,N_16561,N_16812);
nor U17111 (N_17111,N_16707,N_16637);
nand U17112 (N_17112,N_16793,N_16903);
and U17113 (N_17113,N_16996,N_16857);
and U17114 (N_17114,N_16830,N_16751);
nor U17115 (N_17115,N_16635,N_16925);
or U17116 (N_17116,N_16998,N_16659);
nor U17117 (N_17117,N_16533,N_16728);
and U17118 (N_17118,N_16821,N_16831);
nand U17119 (N_17119,N_16723,N_16968);
nor U17120 (N_17120,N_16785,N_16668);
or U17121 (N_17121,N_16516,N_16789);
nor U17122 (N_17122,N_16543,N_16752);
and U17123 (N_17123,N_16755,N_16698);
xnor U17124 (N_17124,N_16833,N_16933);
nand U17125 (N_17125,N_16665,N_16705);
and U17126 (N_17126,N_16502,N_16899);
and U17127 (N_17127,N_16930,N_16727);
nor U17128 (N_17128,N_16559,N_16550);
and U17129 (N_17129,N_16987,N_16551);
xor U17130 (N_17130,N_16919,N_16634);
and U17131 (N_17131,N_16729,N_16845);
nand U17132 (N_17132,N_16935,N_16801);
nor U17133 (N_17133,N_16803,N_16971);
xor U17134 (N_17134,N_16886,N_16746);
nand U17135 (N_17135,N_16609,N_16864);
nor U17136 (N_17136,N_16671,N_16981);
nand U17137 (N_17137,N_16878,N_16757);
nand U17138 (N_17138,N_16666,N_16534);
and U17139 (N_17139,N_16589,N_16847);
xnor U17140 (N_17140,N_16883,N_16924);
and U17141 (N_17141,N_16738,N_16931);
nand U17142 (N_17142,N_16768,N_16872);
nor U17143 (N_17143,N_16822,N_16606);
or U17144 (N_17144,N_16994,N_16947);
or U17145 (N_17145,N_16792,N_16615);
and U17146 (N_17146,N_16740,N_16673);
nor U17147 (N_17147,N_16685,N_16653);
xnor U17148 (N_17148,N_16624,N_16580);
nor U17149 (N_17149,N_16854,N_16747);
or U17150 (N_17150,N_16690,N_16939);
or U17151 (N_17151,N_16913,N_16530);
or U17152 (N_17152,N_16544,N_16515);
nor U17153 (N_17153,N_16541,N_16918);
and U17154 (N_17154,N_16555,N_16696);
nor U17155 (N_17155,N_16744,N_16807);
nor U17156 (N_17156,N_16731,N_16714);
nand U17157 (N_17157,N_16611,N_16726);
nand U17158 (N_17158,N_16846,N_16871);
or U17159 (N_17159,N_16706,N_16927);
nor U17160 (N_17160,N_16575,N_16776);
xnor U17161 (N_17161,N_16588,N_16963);
nor U17162 (N_17162,N_16510,N_16554);
or U17163 (N_17163,N_16828,N_16713);
or U17164 (N_17164,N_16568,N_16767);
and U17165 (N_17165,N_16642,N_16949);
or U17166 (N_17166,N_16923,N_16612);
or U17167 (N_17167,N_16798,N_16638);
and U17168 (N_17168,N_16771,N_16766);
and U17169 (N_17169,N_16988,N_16897);
or U17170 (N_17170,N_16905,N_16632);
and U17171 (N_17171,N_16663,N_16952);
or U17172 (N_17172,N_16509,N_16547);
nand U17173 (N_17173,N_16557,N_16898);
nand U17174 (N_17174,N_16989,N_16716);
nor U17175 (N_17175,N_16724,N_16576);
xor U17176 (N_17176,N_16814,N_16829);
and U17177 (N_17177,N_16503,N_16710);
xor U17178 (N_17178,N_16953,N_16605);
and U17179 (N_17179,N_16517,N_16657);
nor U17180 (N_17180,N_16790,N_16985);
and U17181 (N_17181,N_16895,N_16958);
nor U17182 (N_17182,N_16676,N_16997);
nor U17183 (N_17183,N_16850,N_16528);
xor U17184 (N_17184,N_16954,N_16628);
and U17185 (N_17185,N_16765,N_16593);
nand U17186 (N_17186,N_16523,N_16620);
xnor U17187 (N_17187,N_16802,N_16595);
and U17188 (N_17188,N_16915,N_16800);
nor U17189 (N_17189,N_16795,N_16524);
nor U17190 (N_17190,N_16633,N_16934);
nand U17191 (N_17191,N_16914,N_16623);
or U17192 (N_17192,N_16660,N_16966);
or U17193 (N_17193,N_16827,N_16689);
and U17194 (N_17194,N_16545,N_16955);
nand U17195 (N_17195,N_16819,N_16594);
and U17196 (N_17196,N_16860,N_16693);
or U17197 (N_17197,N_16784,N_16876);
nand U17198 (N_17198,N_16739,N_16680);
and U17199 (N_17199,N_16888,N_16501);
nor U17200 (N_17200,N_16922,N_16736);
or U17201 (N_17201,N_16813,N_16796);
and U17202 (N_17202,N_16754,N_16960);
or U17203 (N_17203,N_16610,N_16773);
nor U17204 (N_17204,N_16756,N_16912);
or U17205 (N_17205,N_16772,N_16725);
xnor U17206 (N_17206,N_16597,N_16948);
or U17207 (N_17207,N_16596,N_16749);
and U17208 (N_17208,N_16943,N_16851);
or U17209 (N_17209,N_16719,N_16945);
nand U17210 (N_17210,N_16840,N_16602);
nand U17211 (N_17211,N_16816,N_16537);
nor U17212 (N_17212,N_16979,N_16621);
or U17213 (N_17213,N_16808,N_16565);
nand U17214 (N_17214,N_16560,N_16519);
nor U17215 (N_17215,N_16926,N_16656);
nand U17216 (N_17216,N_16735,N_16892);
nand U17217 (N_17217,N_16824,N_16675);
xnor U17218 (N_17218,N_16884,N_16995);
nor U17219 (N_17219,N_16891,N_16970);
and U17220 (N_17220,N_16548,N_16977);
and U17221 (N_17221,N_16542,N_16532);
nand U17222 (N_17222,N_16928,N_16900);
and U17223 (N_17223,N_16932,N_16980);
or U17224 (N_17224,N_16944,N_16753);
nand U17225 (N_17225,N_16646,N_16625);
and U17226 (N_17226,N_16745,N_16811);
xnor U17227 (N_17227,N_16907,N_16848);
nor U17228 (N_17228,N_16674,N_16683);
or U17229 (N_17229,N_16645,N_16967);
and U17230 (N_17230,N_16590,N_16702);
or U17231 (N_17231,N_16956,N_16601);
nand U17232 (N_17232,N_16507,N_16782);
nor U17233 (N_17233,N_16708,N_16711);
and U17234 (N_17234,N_16619,N_16608);
nand U17235 (N_17235,N_16973,N_16505);
nand U17236 (N_17236,N_16661,N_16834);
nand U17237 (N_17237,N_16655,N_16783);
or U17238 (N_17238,N_16823,N_16715);
and U17239 (N_17239,N_16525,N_16817);
nand U17240 (N_17240,N_16648,N_16920);
nor U17241 (N_17241,N_16964,N_16640);
nor U17242 (N_17242,N_16836,N_16691);
xnor U17243 (N_17243,N_16867,N_16838);
xor U17244 (N_17244,N_16993,N_16672);
nor U17245 (N_17245,N_16769,N_16904);
or U17246 (N_17246,N_16626,N_16669);
nor U17247 (N_17247,N_16569,N_16961);
nand U17248 (N_17248,N_16709,N_16563);
and U17249 (N_17249,N_16991,N_16852);
or U17250 (N_17250,N_16574,N_16634);
nor U17251 (N_17251,N_16762,N_16611);
xor U17252 (N_17252,N_16801,N_16691);
or U17253 (N_17253,N_16572,N_16673);
and U17254 (N_17254,N_16885,N_16925);
nor U17255 (N_17255,N_16885,N_16631);
nor U17256 (N_17256,N_16829,N_16908);
xor U17257 (N_17257,N_16640,N_16519);
nor U17258 (N_17258,N_16706,N_16797);
and U17259 (N_17259,N_16575,N_16723);
nand U17260 (N_17260,N_16659,N_16823);
and U17261 (N_17261,N_16827,N_16825);
xor U17262 (N_17262,N_16573,N_16936);
or U17263 (N_17263,N_16992,N_16902);
nor U17264 (N_17264,N_16645,N_16834);
or U17265 (N_17265,N_16707,N_16995);
nand U17266 (N_17266,N_16949,N_16971);
and U17267 (N_17267,N_16627,N_16528);
nor U17268 (N_17268,N_16865,N_16947);
nand U17269 (N_17269,N_16501,N_16853);
or U17270 (N_17270,N_16914,N_16875);
nand U17271 (N_17271,N_16744,N_16641);
nand U17272 (N_17272,N_16989,N_16810);
and U17273 (N_17273,N_16608,N_16819);
nor U17274 (N_17274,N_16716,N_16849);
and U17275 (N_17275,N_16633,N_16896);
nor U17276 (N_17276,N_16742,N_16656);
nor U17277 (N_17277,N_16941,N_16572);
nand U17278 (N_17278,N_16987,N_16750);
nand U17279 (N_17279,N_16996,N_16618);
nand U17280 (N_17280,N_16623,N_16787);
nand U17281 (N_17281,N_16957,N_16813);
nor U17282 (N_17282,N_16808,N_16677);
nor U17283 (N_17283,N_16704,N_16969);
xnor U17284 (N_17284,N_16797,N_16808);
nor U17285 (N_17285,N_16878,N_16711);
nor U17286 (N_17286,N_16812,N_16912);
nand U17287 (N_17287,N_16950,N_16588);
nor U17288 (N_17288,N_16912,N_16571);
nand U17289 (N_17289,N_16940,N_16742);
nand U17290 (N_17290,N_16723,N_16639);
and U17291 (N_17291,N_16852,N_16503);
nor U17292 (N_17292,N_16758,N_16508);
nor U17293 (N_17293,N_16863,N_16691);
or U17294 (N_17294,N_16801,N_16989);
or U17295 (N_17295,N_16521,N_16653);
nor U17296 (N_17296,N_16982,N_16972);
or U17297 (N_17297,N_16690,N_16837);
xor U17298 (N_17298,N_16900,N_16558);
and U17299 (N_17299,N_16924,N_16657);
or U17300 (N_17300,N_16637,N_16685);
nor U17301 (N_17301,N_16633,N_16966);
nand U17302 (N_17302,N_16958,N_16503);
and U17303 (N_17303,N_16926,N_16672);
nand U17304 (N_17304,N_16806,N_16615);
nor U17305 (N_17305,N_16813,N_16788);
and U17306 (N_17306,N_16527,N_16574);
xnor U17307 (N_17307,N_16604,N_16854);
nand U17308 (N_17308,N_16632,N_16825);
nor U17309 (N_17309,N_16504,N_16914);
or U17310 (N_17310,N_16673,N_16772);
xor U17311 (N_17311,N_16831,N_16826);
or U17312 (N_17312,N_16647,N_16613);
nor U17313 (N_17313,N_16861,N_16841);
and U17314 (N_17314,N_16972,N_16846);
nand U17315 (N_17315,N_16568,N_16739);
and U17316 (N_17316,N_16861,N_16710);
or U17317 (N_17317,N_16879,N_16885);
nor U17318 (N_17318,N_16653,N_16939);
nor U17319 (N_17319,N_16654,N_16836);
nor U17320 (N_17320,N_16733,N_16993);
and U17321 (N_17321,N_16886,N_16859);
nand U17322 (N_17322,N_16530,N_16740);
and U17323 (N_17323,N_16770,N_16729);
xnor U17324 (N_17324,N_16777,N_16782);
and U17325 (N_17325,N_16593,N_16835);
nand U17326 (N_17326,N_16744,N_16800);
and U17327 (N_17327,N_16982,N_16653);
and U17328 (N_17328,N_16566,N_16613);
nor U17329 (N_17329,N_16746,N_16944);
and U17330 (N_17330,N_16533,N_16688);
and U17331 (N_17331,N_16957,N_16763);
nand U17332 (N_17332,N_16555,N_16801);
or U17333 (N_17333,N_16516,N_16910);
or U17334 (N_17334,N_16702,N_16739);
and U17335 (N_17335,N_16823,N_16981);
and U17336 (N_17336,N_16685,N_16813);
or U17337 (N_17337,N_16993,N_16772);
nor U17338 (N_17338,N_16505,N_16670);
nand U17339 (N_17339,N_16528,N_16744);
xnor U17340 (N_17340,N_16727,N_16739);
nor U17341 (N_17341,N_16900,N_16903);
or U17342 (N_17342,N_16512,N_16575);
or U17343 (N_17343,N_16633,N_16798);
or U17344 (N_17344,N_16902,N_16502);
or U17345 (N_17345,N_16901,N_16987);
or U17346 (N_17346,N_16545,N_16884);
nand U17347 (N_17347,N_16675,N_16828);
and U17348 (N_17348,N_16583,N_16864);
and U17349 (N_17349,N_16824,N_16782);
nor U17350 (N_17350,N_16947,N_16771);
nor U17351 (N_17351,N_16916,N_16660);
xor U17352 (N_17352,N_16677,N_16981);
nor U17353 (N_17353,N_16684,N_16945);
xor U17354 (N_17354,N_16537,N_16834);
or U17355 (N_17355,N_16877,N_16590);
and U17356 (N_17356,N_16621,N_16976);
nand U17357 (N_17357,N_16783,N_16767);
and U17358 (N_17358,N_16619,N_16815);
or U17359 (N_17359,N_16813,N_16758);
and U17360 (N_17360,N_16510,N_16961);
nor U17361 (N_17361,N_16787,N_16594);
or U17362 (N_17362,N_16956,N_16588);
and U17363 (N_17363,N_16984,N_16511);
nor U17364 (N_17364,N_16599,N_16616);
nand U17365 (N_17365,N_16681,N_16869);
nor U17366 (N_17366,N_16900,N_16925);
or U17367 (N_17367,N_16718,N_16501);
and U17368 (N_17368,N_16929,N_16968);
nor U17369 (N_17369,N_16626,N_16926);
or U17370 (N_17370,N_16840,N_16927);
and U17371 (N_17371,N_16690,N_16838);
nand U17372 (N_17372,N_16860,N_16799);
nand U17373 (N_17373,N_16977,N_16573);
nand U17374 (N_17374,N_16854,N_16662);
and U17375 (N_17375,N_16712,N_16932);
nor U17376 (N_17376,N_16910,N_16779);
nand U17377 (N_17377,N_16819,N_16947);
nand U17378 (N_17378,N_16872,N_16790);
and U17379 (N_17379,N_16691,N_16994);
and U17380 (N_17380,N_16993,N_16604);
xor U17381 (N_17381,N_16834,N_16923);
or U17382 (N_17382,N_16702,N_16941);
xor U17383 (N_17383,N_16834,N_16525);
or U17384 (N_17384,N_16533,N_16607);
nor U17385 (N_17385,N_16579,N_16592);
nor U17386 (N_17386,N_16893,N_16958);
or U17387 (N_17387,N_16865,N_16517);
or U17388 (N_17388,N_16876,N_16914);
or U17389 (N_17389,N_16911,N_16630);
nor U17390 (N_17390,N_16790,N_16637);
and U17391 (N_17391,N_16683,N_16731);
or U17392 (N_17392,N_16634,N_16810);
or U17393 (N_17393,N_16959,N_16664);
nand U17394 (N_17394,N_16859,N_16511);
and U17395 (N_17395,N_16890,N_16719);
nor U17396 (N_17396,N_16593,N_16742);
or U17397 (N_17397,N_16886,N_16957);
nand U17398 (N_17398,N_16781,N_16979);
nor U17399 (N_17399,N_16997,N_16843);
nor U17400 (N_17400,N_16902,N_16730);
nor U17401 (N_17401,N_16553,N_16870);
or U17402 (N_17402,N_16560,N_16874);
nand U17403 (N_17403,N_16960,N_16669);
nor U17404 (N_17404,N_16563,N_16891);
nand U17405 (N_17405,N_16739,N_16655);
or U17406 (N_17406,N_16655,N_16701);
nor U17407 (N_17407,N_16964,N_16605);
nand U17408 (N_17408,N_16962,N_16824);
and U17409 (N_17409,N_16935,N_16822);
and U17410 (N_17410,N_16781,N_16986);
and U17411 (N_17411,N_16611,N_16801);
xnor U17412 (N_17412,N_16586,N_16694);
or U17413 (N_17413,N_16951,N_16771);
and U17414 (N_17414,N_16990,N_16908);
or U17415 (N_17415,N_16775,N_16559);
nand U17416 (N_17416,N_16602,N_16782);
nand U17417 (N_17417,N_16556,N_16993);
or U17418 (N_17418,N_16796,N_16877);
nor U17419 (N_17419,N_16576,N_16526);
nor U17420 (N_17420,N_16727,N_16802);
nor U17421 (N_17421,N_16783,N_16614);
or U17422 (N_17422,N_16831,N_16899);
or U17423 (N_17423,N_16779,N_16726);
nand U17424 (N_17424,N_16801,N_16584);
nor U17425 (N_17425,N_16529,N_16606);
nand U17426 (N_17426,N_16916,N_16612);
nand U17427 (N_17427,N_16729,N_16924);
nor U17428 (N_17428,N_16956,N_16732);
nor U17429 (N_17429,N_16610,N_16939);
and U17430 (N_17430,N_16522,N_16931);
and U17431 (N_17431,N_16977,N_16559);
nor U17432 (N_17432,N_16856,N_16838);
nor U17433 (N_17433,N_16725,N_16508);
or U17434 (N_17434,N_16893,N_16667);
nand U17435 (N_17435,N_16904,N_16529);
nor U17436 (N_17436,N_16556,N_16602);
nor U17437 (N_17437,N_16541,N_16505);
nor U17438 (N_17438,N_16546,N_16855);
nor U17439 (N_17439,N_16672,N_16664);
nand U17440 (N_17440,N_16903,N_16869);
nand U17441 (N_17441,N_16553,N_16731);
and U17442 (N_17442,N_16798,N_16772);
and U17443 (N_17443,N_16661,N_16877);
and U17444 (N_17444,N_16581,N_16660);
xor U17445 (N_17445,N_16617,N_16595);
and U17446 (N_17446,N_16608,N_16866);
or U17447 (N_17447,N_16904,N_16526);
nor U17448 (N_17448,N_16704,N_16843);
or U17449 (N_17449,N_16922,N_16592);
or U17450 (N_17450,N_16823,N_16943);
nor U17451 (N_17451,N_16518,N_16623);
nand U17452 (N_17452,N_16650,N_16918);
or U17453 (N_17453,N_16545,N_16918);
nand U17454 (N_17454,N_16600,N_16583);
or U17455 (N_17455,N_16943,N_16921);
nand U17456 (N_17456,N_16749,N_16902);
or U17457 (N_17457,N_16830,N_16626);
and U17458 (N_17458,N_16742,N_16797);
and U17459 (N_17459,N_16543,N_16764);
nand U17460 (N_17460,N_16833,N_16500);
and U17461 (N_17461,N_16577,N_16692);
or U17462 (N_17462,N_16901,N_16974);
nand U17463 (N_17463,N_16749,N_16558);
nor U17464 (N_17464,N_16565,N_16938);
xor U17465 (N_17465,N_16625,N_16864);
nor U17466 (N_17466,N_16992,N_16594);
or U17467 (N_17467,N_16599,N_16785);
nor U17468 (N_17468,N_16675,N_16687);
nor U17469 (N_17469,N_16676,N_16518);
nand U17470 (N_17470,N_16992,N_16773);
and U17471 (N_17471,N_16719,N_16934);
or U17472 (N_17472,N_16892,N_16982);
and U17473 (N_17473,N_16691,N_16653);
and U17474 (N_17474,N_16700,N_16766);
and U17475 (N_17475,N_16649,N_16842);
and U17476 (N_17476,N_16612,N_16516);
or U17477 (N_17477,N_16669,N_16601);
nor U17478 (N_17478,N_16568,N_16853);
and U17479 (N_17479,N_16839,N_16762);
and U17480 (N_17480,N_16628,N_16585);
and U17481 (N_17481,N_16812,N_16537);
nor U17482 (N_17482,N_16939,N_16968);
or U17483 (N_17483,N_16551,N_16934);
nand U17484 (N_17484,N_16674,N_16607);
nand U17485 (N_17485,N_16740,N_16855);
nor U17486 (N_17486,N_16592,N_16678);
nand U17487 (N_17487,N_16879,N_16547);
and U17488 (N_17488,N_16818,N_16802);
nand U17489 (N_17489,N_16898,N_16784);
nor U17490 (N_17490,N_16749,N_16500);
nor U17491 (N_17491,N_16524,N_16844);
nor U17492 (N_17492,N_16574,N_16801);
xnor U17493 (N_17493,N_16842,N_16577);
or U17494 (N_17494,N_16824,N_16763);
and U17495 (N_17495,N_16717,N_16578);
nor U17496 (N_17496,N_16586,N_16674);
nor U17497 (N_17497,N_16625,N_16640);
and U17498 (N_17498,N_16807,N_16534);
or U17499 (N_17499,N_16850,N_16764);
and U17500 (N_17500,N_17229,N_17282);
or U17501 (N_17501,N_17340,N_17001);
or U17502 (N_17502,N_17106,N_17151);
or U17503 (N_17503,N_17235,N_17327);
or U17504 (N_17504,N_17101,N_17481);
nor U17505 (N_17505,N_17209,N_17195);
or U17506 (N_17506,N_17414,N_17048);
nand U17507 (N_17507,N_17354,N_17245);
or U17508 (N_17508,N_17255,N_17356);
nor U17509 (N_17509,N_17444,N_17382);
and U17510 (N_17510,N_17247,N_17013);
nor U17511 (N_17511,N_17049,N_17482);
nand U17512 (N_17512,N_17141,N_17443);
xor U17513 (N_17513,N_17097,N_17402);
nor U17514 (N_17514,N_17188,N_17092);
or U17515 (N_17515,N_17430,N_17012);
or U17516 (N_17516,N_17294,N_17258);
and U17517 (N_17517,N_17221,N_17308);
or U17518 (N_17518,N_17336,N_17051);
nor U17519 (N_17519,N_17373,N_17187);
and U17520 (N_17520,N_17387,N_17031);
nor U17521 (N_17521,N_17413,N_17446);
nor U17522 (N_17522,N_17149,N_17194);
and U17523 (N_17523,N_17253,N_17234);
xnor U17524 (N_17524,N_17041,N_17330);
xnor U17525 (N_17525,N_17244,N_17168);
nand U17526 (N_17526,N_17071,N_17409);
and U17527 (N_17527,N_17456,N_17321);
and U17528 (N_17528,N_17000,N_17355);
nand U17529 (N_17529,N_17096,N_17262);
or U17530 (N_17530,N_17197,N_17098);
and U17531 (N_17531,N_17448,N_17326);
and U17532 (N_17532,N_17062,N_17124);
or U17533 (N_17533,N_17046,N_17167);
nand U17534 (N_17534,N_17475,N_17017);
nor U17535 (N_17535,N_17399,N_17289);
and U17536 (N_17536,N_17192,N_17349);
nand U17537 (N_17537,N_17045,N_17054);
or U17538 (N_17538,N_17014,N_17395);
xor U17539 (N_17539,N_17180,N_17135);
nand U17540 (N_17540,N_17074,N_17237);
or U17541 (N_17541,N_17385,N_17155);
or U17542 (N_17542,N_17021,N_17496);
and U17543 (N_17543,N_17199,N_17346);
xor U17544 (N_17544,N_17086,N_17064);
and U17545 (N_17545,N_17019,N_17468);
nor U17546 (N_17546,N_17206,N_17302);
or U17547 (N_17547,N_17470,N_17478);
and U17548 (N_17548,N_17408,N_17236);
and U17549 (N_17549,N_17488,N_17486);
nand U17550 (N_17550,N_17281,N_17497);
or U17551 (N_17551,N_17028,N_17100);
nor U17552 (N_17552,N_17052,N_17334);
and U17553 (N_17553,N_17069,N_17147);
nor U17554 (N_17554,N_17251,N_17285);
nor U17555 (N_17555,N_17227,N_17304);
nand U17556 (N_17556,N_17161,N_17472);
nor U17557 (N_17557,N_17146,N_17118);
or U17558 (N_17558,N_17034,N_17176);
nor U17559 (N_17559,N_17172,N_17437);
or U17560 (N_17560,N_17498,N_17133);
nor U17561 (N_17561,N_17317,N_17166);
or U17562 (N_17562,N_17136,N_17309);
xnor U17563 (N_17563,N_17239,N_17094);
and U17564 (N_17564,N_17451,N_17366);
or U17565 (N_17565,N_17174,N_17431);
nand U17566 (N_17566,N_17427,N_17440);
and U17567 (N_17567,N_17314,N_17162);
nand U17568 (N_17568,N_17002,N_17128);
xnor U17569 (N_17569,N_17277,N_17307);
or U17570 (N_17570,N_17053,N_17068);
and U17571 (N_17571,N_17248,N_17464);
and U17572 (N_17572,N_17156,N_17339);
nand U17573 (N_17573,N_17193,N_17202);
and U17574 (N_17574,N_17404,N_17150);
nor U17575 (N_17575,N_17113,N_17479);
or U17576 (N_17576,N_17060,N_17087);
xor U17577 (N_17577,N_17441,N_17127);
or U17578 (N_17578,N_17471,N_17445);
or U17579 (N_17579,N_17350,N_17211);
and U17580 (N_17580,N_17463,N_17333);
or U17581 (N_17581,N_17272,N_17186);
or U17582 (N_17582,N_17424,N_17119);
nor U17583 (N_17583,N_17175,N_17061);
nor U17584 (N_17584,N_17417,N_17400);
nand U17585 (N_17585,N_17210,N_17439);
or U17586 (N_17586,N_17114,N_17015);
xor U17587 (N_17587,N_17191,N_17035);
and U17588 (N_17588,N_17325,N_17261);
and U17589 (N_17589,N_17213,N_17422);
nor U17590 (N_17590,N_17341,N_17215);
and U17591 (N_17591,N_17222,N_17225);
or U17592 (N_17592,N_17429,N_17485);
nor U17593 (N_17593,N_17072,N_17415);
and U17594 (N_17594,N_17280,N_17489);
or U17595 (N_17595,N_17286,N_17303);
nand U17596 (N_17596,N_17364,N_17025);
xnor U17597 (N_17597,N_17453,N_17105);
and U17598 (N_17598,N_17393,N_17335);
nand U17599 (N_17599,N_17059,N_17425);
xnor U17600 (N_17600,N_17203,N_17063);
nor U17601 (N_17601,N_17284,N_17365);
nor U17602 (N_17602,N_17142,N_17143);
and U17603 (N_17603,N_17338,N_17200);
and U17604 (N_17604,N_17005,N_17290);
nand U17605 (N_17605,N_17216,N_17270);
or U17606 (N_17606,N_17416,N_17291);
and U17607 (N_17607,N_17140,N_17158);
nor U17608 (N_17608,N_17426,N_17265);
xor U17609 (N_17609,N_17065,N_17165);
and U17610 (N_17610,N_17018,N_17138);
nand U17611 (N_17611,N_17102,N_17358);
or U17612 (N_17612,N_17466,N_17360);
or U17613 (N_17613,N_17132,N_17075);
or U17614 (N_17614,N_17287,N_17322);
nor U17615 (N_17615,N_17331,N_17357);
and U17616 (N_17616,N_17306,N_17348);
nor U17617 (N_17617,N_17389,N_17438);
nand U17618 (N_17618,N_17420,N_17205);
nand U17619 (N_17619,N_17368,N_17010);
or U17620 (N_17620,N_17103,N_17397);
or U17621 (N_17621,N_17020,N_17076);
nor U17622 (N_17622,N_17109,N_17108);
or U17623 (N_17623,N_17337,N_17465);
or U17624 (N_17624,N_17469,N_17264);
and U17625 (N_17625,N_17288,N_17487);
and U17626 (N_17626,N_17233,N_17042);
or U17627 (N_17627,N_17079,N_17372);
nand U17628 (N_17628,N_17173,N_17342);
and U17629 (N_17629,N_17148,N_17003);
nand U17630 (N_17630,N_17240,N_17371);
nand U17631 (N_17631,N_17329,N_17266);
or U17632 (N_17632,N_17169,N_17131);
or U17633 (N_17633,N_17104,N_17467);
nand U17634 (N_17634,N_17091,N_17243);
xor U17635 (N_17635,N_17083,N_17328);
nor U17636 (N_17636,N_17219,N_17401);
nor U17637 (N_17637,N_17170,N_17311);
nand U17638 (N_17638,N_17116,N_17037);
or U17639 (N_17639,N_17057,N_17082);
nor U17640 (N_17640,N_17353,N_17207);
xnor U17641 (N_17641,N_17318,N_17381);
nor U17642 (N_17642,N_17230,N_17492);
nand U17643 (N_17643,N_17436,N_17078);
and U17644 (N_17644,N_17198,N_17386);
nand U17645 (N_17645,N_17345,N_17295);
nand U17646 (N_17646,N_17405,N_17231);
nand U17647 (N_17647,N_17184,N_17299);
and U17648 (N_17648,N_17305,N_17218);
nand U17649 (N_17649,N_17190,N_17499);
nand U17650 (N_17650,N_17275,N_17370);
xnor U17651 (N_17651,N_17178,N_17374);
and U17652 (N_17652,N_17145,N_17055);
nor U17653 (N_17653,N_17183,N_17455);
nand U17654 (N_17654,N_17319,N_17112);
and U17655 (N_17655,N_17279,N_17312);
nor U17656 (N_17656,N_17004,N_17458);
xnor U17657 (N_17657,N_17232,N_17073);
nand U17658 (N_17658,N_17375,N_17406);
and U17659 (N_17659,N_17457,N_17434);
and U17660 (N_17660,N_17367,N_17412);
nand U17661 (N_17661,N_17477,N_17423);
nand U17662 (N_17662,N_17208,N_17214);
nor U17663 (N_17663,N_17450,N_17352);
and U17664 (N_17664,N_17171,N_17452);
nand U17665 (N_17665,N_17257,N_17139);
or U17666 (N_17666,N_17377,N_17058);
nand U17667 (N_17667,N_17007,N_17315);
nor U17668 (N_17668,N_17196,N_17241);
xor U17669 (N_17669,N_17181,N_17316);
nor U17670 (N_17670,N_17454,N_17081);
nor U17671 (N_17671,N_17369,N_17220);
nor U17672 (N_17672,N_17029,N_17276);
and U17673 (N_17673,N_17421,N_17050);
xnor U17674 (N_17674,N_17152,N_17310);
nor U17675 (N_17675,N_17296,N_17269);
nand U17676 (N_17676,N_17023,N_17398);
and U17677 (N_17677,N_17493,N_17332);
nor U17678 (N_17678,N_17107,N_17077);
or U17679 (N_17679,N_17410,N_17343);
nor U17680 (N_17680,N_17204,N_17473);
or U17681 (N_17681,N_17223,N_17238);
nor U17682 (N_17682,N_17024,N_17449);
xor U17683 (N_17683,N_17088,N_17383);
nand U17684 (N_17684,N_17320,N_17495);
nand U17685 (N_17685,N_17164,N_17297);
nor U17686 (N_17686,N_17484,N_17278);
xnor U17687 (N_17687,N_17126,N_17144);
nor U17688 (N_17688,N_17130,N_17163);
and U17689 (N_17689,N_17324,N_17036);
nand U17690 (N_17690,N_17388,N_17435);
nor U17691 (N_17691,N_17390,N_17267);
nand U17692 (N_17692,N_17047,N_17418);
nor U17693 (N_17693,N_17376,N_17380);
nor U17694 (N_17694,N_17379,N_17407);
or U17695 (N_17695,N_17252,N_17110);
nand U17696 (N_17696,N_17044,N_17259);
nand U17697 (N_17697,N_17032,N_17268);
and U17698 (N_17698,N_17474,N_17384);
nand U17699 (N_17699,N_17351,N_17403);
and U17700 (N_17700,N_17117,N_17300);
and U17701 (N_17701,N_17459,N_17298);
and U17702 (N_17702,N_17033,N_17494);
nand U17703 (N_17703,N_17084,N_17125);
and U17704 (N_17704,N_17263,N_17122);
xor U17705 (N_17705,N_17392,N_17123);
xor U17706 (N_17706,N_17011,N_17056);
nor U17707 (N_17707,N_17189,N_17038);
and U17708 (N_17708,N_17153,N_17447);
and U17709 (N_17709,N_17362,N_17480);
and U17710 (N_17710,N_17301,N_17027);
and U17711 (N_17711,N_17157,N_17428);
nand U17712 (N_17712,N_17040,N_17160);
nand U17713 (N_17713,N_17432,N_17120);
or U17714 (N_17714,N_17090,N_17391);
nor U17715 (N_17715,N_17228,N_17217);
or U17716 (N_17716,N_17111,N_17030);
nand U17717 (N_17717,N_17080,N_17129);
and U17718 (N_17718,N_17121,N_17022);
and U17719 (N_17719,N_17185,N_17066);
nand U17720 (N_17720,N_17095,N_17246);
nand U17721 (N_17721,N_17067,N_17043);
nand U17722 (N_17722,N_17201,N_17292);
or U17723 (N_17723,N_17271,N_17085);
nor U17724 (N_17724,N_17254,N_17260);
or U17725 (N_17725,N_17115,N_17009);
nand U17726 (N_17726,N_17347,N_17226);
nor U17727 (N_17727,N_17483,N_17323);
or U17728 (N_17728,N_17159,N_17224);
and U17729 (N_17729,N_17274,N_17293);
and U17730 (N_17730,N_17442,N_17460);
nor U17731 (N_17731,N_17250,N_17490);
nor U17732 (N_17732,N_17179,N_17008);
or U17733 (N_17733,N_17344,N_17433);
xnor U17734 (N_17734,N_17089,N_17462);
and U17735 (N_17735,N_17154,N_17137);
and U17736 (N_17736,N_17378,N_17396);
nand U17737 (N_17737,N_17016,N_17491);
or U17738 (N_17738,N_17070,N_17026);
nand U17739 (N_17739,N_17461,N_17273);
or U17740 (N_17740,N_17411,N_17256);
or U17741 (N_17741,N_17361,N_17359);
and U17742 (N_17742,N_17134,N_17093);
nand U17743 (N_17743,N_17212,N_17242);
nor U17744 (N_17744,N_17177,N_17099);
nor U17745 (N_17745,N_17419,N_17039);
nor U17746 (N_17746,N_17313,N_17283);
or U17747 (N_17747,N_17249,N_17182);
nor U17748 (N_17748,N_17363,N_17394);
nand U17749 (N_17749,N_17476,N_17006);
nand U17750 (N_17750,N_17129,N_17479);
nor U17751 (N_17751,N_17484,N_17229);
nor U17752 (N_17752,N_17036,N_17434);
nor U17753 (N_17753,N_17415,N_17148);
or U17754 (N_17754,N_17320,N_17312);
nand U17755 (N_17755,N_17118,N_17200);
xor U17756 (N_17756,N_17238,N_17115);
and U17757 (N_17757,N_17045,N_17433);
nor U17758 (N_17758,N_17058,N_17197);
xor U17759 (N_17759,N_17085,N_17091);
or U17760 (N_17760,N_17450,N_17205);
nor U17761 (N_17761,N_17222,N_17426);
and U17762 (N_17762,N_17059,N_17146);
or U17763 (N_17763,N_17454,N_17399);
and U17764 (N_17764,N_17462,N_17058);
and U17765 (N_17765,N_17423,N_17088);
xnor U17766 (N_17766,N_17372,N_17380);
nand U17767 (N_17767,N_17077,N_17006);
and U17768 (N_17768,N_17013,N_17005);
nor U17769 (N_17769,N_17053,N_17092);
nand U17770 (N_17770,N_17492,N_17079);
and U17771 (N_17771,N_17258,N_17309);
or U17772 (N_17772,N_17304,N_17422);
nand U17773 (N_17773,N_17391,N_17252);
and U17774 (N_17774,N_17206,N_17445);
nand U17775 (N_17775,N_17404,N_17359);
and U17776 (N_17776,N_17179,N_17446);
or U17777 (N_17777,N_17367,N_17446);
and U17778 (N_17778,N_17122,N_17374);
xnor U17779 (N_17779,N_17476,N_17265);
and U17780 (N_17780,N_17277,N_17168);
and U17781 (N_17781,N_17369,N_17447);
nor U17782 (N_17782,N_17211,N_17418);
and U17783 (N_17783,N_17412,N_17341);
nor U17784 (N_17784,N_17147,N_17226);
and U17785 (N_17785,N_17429,N_17436);
and U17786 (N_17786,N_17135,N_17243);
nand U17787 (N_17787,N_17085,N_17391);
nor U17788 (N_17788,N_17135,N_17225);
xor U17789 (N_17789,N_17071,N_17192);
nand U17790 (N_17790,N_17402,N_17050);
nand U17791 (N_17791,N_17086,N_17000);
or U17792 (N_17792,N_17306,N_17196);
or U17793 (N_17793,N_17325,N_17370);
nor U17794 (N_17794,N_17384,N_17391);
nand U17795 (N_17795,N_17353,N_17177);
nand U17796 (N_17796,N_17271,N_17016);
or U17797 (N_17797,N_17372,N_17014);
nor U17798 (N_17798,N_17467,N_17462);
nor U17799 (N_17799,N_17046,N_17021);
and U17800 (N_17800,N_17412,N_17053);
nand U17801 (N_17801,N_17413,N_17062);
nand U17802 (N_17802,N_17346,N_17109);
or U17803 (N_17803,N_17276,N_17330);
or U17804 (N_17804,N_17023,N_17129);
or U17805 (N_17805,N_17496,N_17197);
nor U17806 (N_17806,N_17410,N_17415);
nor U17807 (N_17807,N_17390,N_17227);
nand U17808 (N_17808,N_17135,N_17211);
xnor U17809 (N_17809,N_17108,N_17469);
or U17810 (N_17810,N_17376,N_17276);
nand U17811 (N_17811,N_17483,N_17275);
nand U17812 (N_17812,N_17439,N_17380);
nor U17813 (N_17813,N_17474,N_17299);
and U17814 (N_17814,N_17360,N_17497);
nor U17815 (N_17815,N_17100,N_17217);
nor U17816 (N_17816,N_17497,N_17332);
or U17817 (N_17817,N_17188,N_17218);
or U17818 (N_17818,N_17114,N_17156);
nand U17819 (N_17819,N_17260,N_17285);
nor U17820 (N_17820,N_17054,N_17111);
nand U17821 (N_17821,N_17436,N_17065);
nor U17822 (N_17822,N_17173,N_17157);
nor U17823 (N_17823,N_17391,N_17103);
and U17824 (N_17824,N_17331,N_17052);
nand U17825 (N_17825,N_17042,N_17083);
nor U17826 (N_17826,N_17306,N_17431);
nand U17827 (N_17827,N_17180,N_17386);
nand U17828 (N_17828,N_17222,N_17279);
or U17829 (N_17829,N_17497,N_17358);
xnor U17830 (N_17830,N_17109,N_17318);
and U17831 (N_17831,N_17074,N_17147);
or U17832 (N_17832,N_17306,N_17201);
nor U17833 (N_17833,N_17072,N_17410);
or U17834 (N_17834,N_17336,N_17398);
or U17835 (N_17835,N_17321,N_17373);
nor U17836 (N_17836,N_17271,N_17249);
xor U17837 (N_17837,N_17132,N_17466);
and U17838 (N_17838,N_17359,N_17235);
and U17839 (N_17839,N_17459,N_17416);
and U17840 (N_17840,N_17469,N_17217);
nor U17841 (N_17841,N_17470,N_17209);
and U17842 (N_17842,N_17366,N_17402);
nor U17843 (N_17843,N_17227,N_17216);
nand U17844 (N_17844,N_17068,N_17103);
nor U17845 (N_17845,N_17047,N_17491);
and U17846 (N_17846,N_17234,N_17208);
xor U17847 (N_17847,N_17400,N_17185);
nand U17848 (N_17848,N_17423,N_17385);
nand U17849 (N_17849,N_17185,N_17284);
nor U17850 (N_17850,N_17184,N_17498);
xor U17851 (N_17851,N_17364,N_17339);
and U17852 (N_17852,N_17210,N_17302);
nor U17853 (N_17853,N_17253,N_17108);
nor U17854 (N_17854,N_17298,N_17125);
nor U17855 (N_17855,N_17436,N_17082);
and U17856 (N_17856,N_17100,N_17141);
and U17857 (N_17857,N_17481,N_17204);
and U17858 (N_17858,N_17402,N_17414);
nor U17859 (N_17859,N_17351,N_17130);
nand U17860 (N_17860,N_17090,N_17125);
nor U17861 (N_17861,N_17485,N_17400);
or U17862 (N_17862,N_17376,N_17184);
nor U17863 (N_17863,N_17139,N_17280);
nor U17864 (N_17864,N_17244,N_17475);
and U17865 (N_17865,N_17397,N_17224);
or U17866 (N_17866,N_17049,N_17222);
and U17867 (N_17867,N_17364,N_17144);
or U17868 (N_17868,N_17013,N_17125);
nand U17869 (N_17869,N_17449,N_17041);
or U17870 (N_17870,N_17182,N_17434);
xnor U17871 (N_17871,N_17003,N_17039);
nor U17872 (N_17872,N_17365,N_17160);
nand U17873 (N_17873,N_17077,N_17349);
nor U17874 (N_17874,N_17131,N_17130);
nor U17875 (N_17875,N_17408,N_17189);
or U17876 (N_17876,N_17324,N_17253);
and U17877 (N_17877,N_17394,N_17328);
or U17878 (N_17878,N_17009,N_17000);
nand U17879 (N_17879,N_17231,N_17272);
xor U17880 (N_17880,N_17227,N_17376);
and U17881 (N_17881,N_17007,N_17444);
and U17882 (N_17882,N_17444,N_17142);
and U17883 (N_17883,N_17158,N_17075);
and U17884 (N_17884,N_17067,N_17310);
or U17885 (N_17885,N_17181,N_17466);
nand U17886 (N_17886,N_17394,N_17285);
nor U17887 (N_17887,N_17058,N_17030);
nand U17888 (N_17888,N_17034,N_17084);
xnor U17889 (N_17889,N_17399,N_17365);
nand U17890 (N_17890,N_17431,N_17309);
or U17891 (N_17891,N_17334,N_17107);
or U17892 (N_17892,N_17285,N_17051);
nor U17893 (N_17893,N_17211,N_17017);
nand U17894 (N_17894,N_17327,N_17462);
and U17895 (N_17895,N_17015,N_17438);
xor U17896 (N_17896,N_17226,N_17154);
or U17897 (N_17897,N_17273,N_17124);
nand U17898 (N_17898,N_17037,N_17365);
nor U17899 (N_17899,N_17377,N_17492);
nand U17900 (N_17900,N_17350,N_17046);
nor U17901 (N_17901,N_17170,N_17372);
and U17902 (N_17902,N_17147,N_17148);
and U17903 (N_17903,N_17179,N_17427);
or U17904 (N_17904,N_17309,N_17314);
xor U17905 (N_17905,N_17155,N_17065);
nand U17906 (N_17906,N_17180,N_17384);
nor U17907 (N_17907,N_17226,N_17202);
or U17908 (N_17908,N_17469,N_17402);
and U17909 (N_17909,N_17493,N_17430);
and U17910 (N_17910,N_17405,N_17099);
nor U17911 (N_17911,N_17301,N_17405);
nand U17912 (N_17912,N_17160,N_17298);
nand U17913 (N_17913,N_17101,N_17488);
nor U17914 (N_17914,N_17450,N_17395);
and U17915 (N_17915,N_17350,N_17467);
nor U17916 (N_17916,N_17319,N_17028);
nor U17917 (N_17917,N_17060,N_17203);
nor U17918 (N_17918,N_17268,N_17381);
and U17919 (N_17919,N_17008,N_17028);
and U17920 (N_17920,N_17182,N_17153);
and U17921 (N_17921,N_17018,N_17422);
nor U17922 (N_17922,N_17280,N_17420);
nand U17923 (N_17923,N_17206,N_17392);
and U17924 (N_17924,N_17383,N_17074);
or U17925 (N_17925,N_17045,N_17001);
nand U17926 (N_17926,N_17230,N_17250);
nor U17927 (N_17927,N_17051,N_17313);
or U17928 (N_17928,N_17097,N_17228);
xnor U17929 (N_17929,N_17308,N_17439);
nor U17930 (N_17930,N_17360,N_17317);
xor U17931 (N_17931,N_17487,N_17292);
or U17932 (N_17932,N_17084,N_17481);
nand U17933 (N_17933,N_17458,N_17091);
nor U17934 (N_17934,N_17036,N_17250);
nand U17935 (N_17935,N_17169,N_17179);
and U17936 (N_17936,N_17361,N_17418);
nand U17937 (N_17937,N_17189,N_17204);
or U17938 (N_17938,N_17369,N_17495);
and U17939 (N_17939,N_17019,N_17466);
nand U17940 (N_17940,N_17026,N_17325);
nor U17941 (N_17941,N_17250,N_17470);
nor U17942 (N_17942,N_17040,N_17343);
and U17943 (N_17943,N_17207,N_17321);
and U17944 (N_17944,N_17129,N_17218);
xnor U17945 (N_17945,N_17270,N_17480);
and U17946 (N_17946,N_17155,N_17011);
and U17947 (N_17947,N_17151,N_17456);
and U17948 (N_17948,N_17423,N_17076);
nor U17949 (N_17949,N_17444,N_17133);
nand U17950 (N_17950,N_17045,N_17094);
or U17951 (N_17951,N_17372,N_17382);
nand U17952 (N_17952,N_17012,N_17000);
or U17953 (N_17953,N_17335,N_17089);
xor U17954 (N_17954,N_17309,N_17225);
and U17955 (N_17955,N_17218,N_17296);
and U17956 (N_17956,N_17368,N_17450);
nand U17957 (N_17957,N_17058,N_17128);
or U17958 (N_17958,N_17490,N_17061);
or U17959 (N_17959,N_17179,N_17473);
nand U17960 (N_17960,N_17489,N_17413);
nand U17961 (N_17961,N_17193,N_17015);
nor U17962 (N_17962,N_17037,N_17341);
nor U17963 (N_17963,N_17353,N_17226);
xnor U17964 (N_17964,N_17342,N_17065);
and U17965 (N_17965,N_17432,N_17495);
xor U17966 (N_17966,N_17297,N_17232);
or U17967 (N_17967,N_17053,N_17492);
and U17968 (N_17968,N_17035,N_17102);
and U17969 (N_17969,N_17276,N_17289);
or U17970 (N_17970,N_17062,N_17201);
nand U17971 (N_17971,N_17431,N_17334);
xnor U17972 (N_17972,N_17260,N_17037);
or U17973 (N_17973,N_17131,N_17070);
nor U17974 (N_17974,N_17482,N_17471);
and U17975 (N_17975,N_17370,N_17383);
or U17976 (N_17976,N_17407,N_17496);
xnor U17977 (N_17977,N_17029,N_17234);
or U17978 (N_17978,N_17247,N_17341);
and U17979 (N_17979,N_17235,N_17345);
nand U17980 (N_17980,N_17429,N_17418);
xor U17981 (N_17981,N_17219,N_17159);
nand U17982 (N_17982,N_17013,N_17006);
or U17983 (N_17983,N_17440,N_17085);
xor U17984 (N_17984,N_17104,N_17239);
xnor U17985 (N_17985,N_17265,N_17349);
or U17986 (N_17986,N_17454,N_17326);
nor U17987 (N_17987,N_17040,N_17177);
or U17988 (N_17988,N_17209,N_17203);
and U17989 (N_17989,N_17145,N_17305);
or U17990 (N_17990,N_17122,N_17202);
xnor U17991 (N_17991,N_17169,N_17375);
and U17992 (N_17992,N_17357,N_17100);
and U17993 (N_17993,N_17271,N_17241);
xnor U17994 (N_17994,N_17466,N_17177);
nand U17995 (N_17995,N_17117,N_17017);
nand U17996 (N_17996,N_17164,N_17073);
nand U17997 (N_17997,N_17195,N_17342);
xor U17998 (N_17998,N_17150,N_17468);
or U17999 (N_17999,N_17228,N_17114);
xnor U18000 (N_18000,N_17528,N_17681);
xnor U18001 (N_18001,N_17522,N_17586);
and U18002 (N_18002,N_17782,N_17870);
and U18003 (N_18003,N_17701,N_17737);
and U18004 (N_18004,N_17729,N_17665);
nor U18005 (N_18005,N_17839,N_17962);
nor U18006 (N_18006,N_17874,N_17551);
or U18007 (N_18007,N_17695,N_17976);
and U18008 (N_18008,N_17602,N_17856);
nor U18009 (N_18009,N_17584,N_17595);
or U18010 (N_18010,N_17974,N_17670);
nand U18011 (N_18011,N_17575,N_17654);
nor U18012 (N_18012,N_17802,N_17863);
and U18013 (N_18013,N_17535,N_17912);
nand U18014 (N_18014,N_17752,N_17953);
nand U18015 (N_18015,N_17588,N_17941);
nand U18016 (N_18016,N_17574,N_17753);
xnor U18017 (N_18017,N_17795,N_17609);
xor U18018 (N_18018,N_17950,N_17655);
or U18019 (N_18019,N_17608,N_17997);
nand U18020 (N_18020,N_17909,N_17790);
nor U18021 (N_18021,N_17508,N_17754);
nand U18022 (N_18022,N_17559,N_17973);
and U18023 (N_18023,N_17623,N_17774);
or U18024 (N_18024,N_17809,N_17759);
nor U18025 (N_18025,N_17614,N_17893);
nand U18026 (N_18026,N_17514,N_17859);
and U18027 (N_18027,N_17851,N_17642);
nand U18028 (N_18028,N_17924,N_17986);
and U18029 (N_18029,N_17748,N_17747);
or U18030 (N_18030,N_17844,N_17880);
nand U18031 (N_18031,N_17589,N_17547);
nand U18032 (N_18032,N_17662,N_17980);
and U18033 (N_18033,N_17762,N_17597);
and U18034 (N_18034,N_17627,N_17557);
nand U18035 (N_18035,N_17920,N_17938);
and U18036 (N_18036,N_17587,N_17702);
or U18037 (N_18037,N_17720,N_17860);
or U18038 (N_18038,N_17883,N_17657);
xnor U18039 (N_18039,N_17675,N_17686);
and U18040 (N_18040,N_17612,N_17668);
and U18041 (N_18041,N_17576,N_17871);
or U18042 (N_18042,N_17733,N_17847);
nand U18043 (N_18043,N_17850,N_17968);
nor U18044 (N_18044,N_17821,N_17591);
and U18045 (N_18045,N_17827,N_17961);
and U18046 (N_18046,N_17635,N_17512);
and U18047 (N_18047,N_17780,N_17788);
xnor U18048 (N_18048,N_17823,N_17676);
nand U18049 (N_18049,N_17836,N_17845);
nand U18050 (N_18050,N_17598,N_17704);
nor U18051 (N_18051,N_17690,N_17817);
and U18052 (N_18052,N_17825,N_17699);
or U18053 (N_18053,N_17711,N_17682);
or U18054 (N_18054,N_17855,N_17915);
and U18055 (N_18055,N_17777,N_17698);
nor U18056 (N_18056,N_17914,N_17792);
nand U18057 (N_18057,N_17877,N_17800);
and U18058 (N_18058,N_17913,N_17744);
nand U18059 (N_18059,N_17515,N_17735);
nand U18060 (N_18060,N_17793,N_17542);
and U18061 (N_18061,N_17583,N_17843);
nor U18062 (N_18062,N_17873,N_17904);
and U18063 (N_18063,N_17803,N_17728);
and U18064 (N_18064,N_17911,N_17977);
nor U18065 (N_18065,N_17537,N_17771);
nor U18066 (N_18066,N_17978,N_17837);
and U18067 (N_18067,N_17956,N_17981);
nor U18068 (N_18068,N_17760,N_17633);
and U18069 (N_18069,N_17523,N_17710);
nand U18070 (N_18070,N_17922,N_17745);
or U18071 (N_18071,N_17969,N_17677);
nor U18072 (N_18072,N_17556,N_17683);
or U18073 (N_18073,N_17765,N_17822);
nand U18074 (N_18074,N_17524,N_17776);
and U18075 (N_18075,N_17755,N_17819);
nor U18076 (N_18076,N_17810,N_17879);
and U18077 (N_18077,N_17831,N_17562);
and U18078 (N_18078,N_17884,N_17910);
or U18079 (N_18079,N_17533,N_17707);
nor U18080 (N_18080,N_17585,N_17580);
nand U18081 (N_18081,N_17526,N_17749);
nor U18082 (N_18082,N_17518,N_17621);
and U18083 (N_18083,N_17814,N_17541);
nand U18084 (N_18084,N_17853,N_17693);
and U18085 (N_18085,N_17996,N_17740);
nand U18086 (N_18086,N_17527,N_17954);
xnor U18087 (N_18087,N_17797,N_17544);
nor U18088 (N_18088,N_17942,N_17935);
and U18089 (N_18089,N_17897,N_17939);
or U18090 (N_18090,N_17875,N_17769);
xor U18091 (N_18091,N_17966,N_17645);
nand U18092 (N_18092,N_17649,N_17592);
and U18093 (N_18093,N_17715,N_17948);
nor U18094 (N_18094,N_17507,N_17743);
and U18095 (N_18095,N_17898,N_17687);
nand U18096 (N_18096,N_17739,N_17947);
nand U18097 (N_18097,N_17640,N_17620);
nor U18098 (N_18098,N_17727,N_17896);
nor U18099 (N_18099,N_17931,N_17830);
and U18100 (N_18100,N_17804,N_17503);
nand U18101 (N_18101,N_17929,N_17990);
or U18102 (N_18102,N_17918,N_17758);
nand U18103 (N_18103,N_17519,N_17786);
nor U18104 (N_18104,N_17638,N_17594);
nand U18105 (N_18105,N_17680,N_17987);
nor U18106 (N_18106,N_17553,N_17960);
xor U18107 (N_18107,N_17555,N_17626);
xnor U18108 (N_18108,N_17878,N_17779);
and U18109 (N_18109,N_17516,N_17561);
and U18110 (N_18110,N_17500,N_17796);
and U18111 (N_18111,N_17549,N_17824);
and U18112 (N_18112,N_17894,N_17805);
and U18113 (N_18113,N_17998,N_17509);
nor U18114 (N_18114,N_17854,N_17852);
and U18115 (N_18115,N_17732,N_17937);
nand U18116 (N_18116,N_17659,N_17599);
nor U18117 (N_18117,N_17919,N_17653);
and U18118 (N_18118,N_17502,N_17988);
xor U18119 (N_18119,N_17892,N_17573);
nor U18120 (N_18120,N_17866,N_17572);
and U18121 (N_18121,N_17926,N_17949);
nand U18122 (N_18122,N_17766,N_17634);
nor U18123 (N_18123,N_17724,N_17846);
and U18124 (N_18124,N_17579,N_17603);
nand U18125 (N_18125,N_17770,N_17921);
or U18126 (N_18126,N_17833,N_17965);
or U18127 (N_18127,N_17504,N_17857);
nand U18128 (N_18128,N_17558,N_17881);
and U18129 (N_18129,N_17708,N_17905);
nand U18130 (N_18130,N_17505,N_17959);
or U18131 (N_18131,N_17826,N_17889);
and U18132 (N_18132,N_17607,N_17664);
or U18133 (N_18133,N_17652,N_17784);
nor U18134 (N_18134,N_17582,N_17781);
nand U18135 (N_18135,N_17807,N_17991);
or U18136 (N_18136,N_17725,N_17722);
nor U18137 (N_18137,N_17958,N_17577);
or U18138 (N_18138,N_17689,N_17726);
and U18139 (N_18139,N_17798,N_17811);
nor U18140 (N_18140,N_17813,N_17818);
nor U18141 (N_18141,N_17712,N_17964);
or U18142 (N_18142,N_17650,N_17674);
or U18143 (N_18143,N_17861,N_17713);
xor U18144 (N_18144,N_17778,N_17511);
nand U18145 (N_18145,N_17775,N_17936);
or U18146 (N_18146,N_17692,N_17546);
xnor U18147 (N_18147,N_17746,N_17940);
nor U18148 (N_18148,N_17899,N_17791);
nor U18149 (N_18149,N_17705,N_17773);
nor U18150 (N_18150,N_17995,N_17646);
or U18151 (N_18151,N_17891,N_17761);
and U18152 (N_18152,N_17691,N_17887);
nor U18153 (N_18153,N_17764,N_17841);
or U18154 (N_18154,N_17679,N_17631);
and U18155 (N_18155,N_17536,N_17628);
nor U18156 (N_18156,N_17714,N_17916);
and U18157 (N_18157,N_17566,N_17742);
nor U18158 (N_18158,N_17787,N_17751);
and U18159 (N_18159,N_17678,N_17605);
nor U18160 (N_18160,N_17581,N_17928);
nor U18161 (N_18161,N_17719,N_17886);
nor U18162 (N_18162,N_17967,N_17858);
nand U18163 (N_18163,N_17907,N_17756);
and U18164 (N_18164,N_17625,N_17906);
or U18165 (N_18165,N_17658,N_17994);
nor U18166 (N_18166,N_17815,N_17517);
or U18167 (N_18167,N_17501,N_17783);
and U18168 (N_18168,N_17694,N_17848);
and U18169 (N_18169,N_17540,N_17944);
or U18170 (N_18170,N_17552,N_17569);
xor U18171 (N_18171,N_17864,N_17917);
or U18172 (N_18172,N_17616,N_17721);
nor U18173 (N_18173,N_17606,N_17930);
nor U18174 (N_18174,N_17736,N_17543);
xnor U18175 (N_18175,N_17900,N_17660);
nand U18176 (N_18176,N_17666,N_17510);
nor U18177 (N_18177,N_17868,N_17521);
nand U18178 (N_18178,N_17943,N_17596);
nor U18179 (N_18179,N_17975,N_17685);
nor U18180 (N_18180,N_17550,N_17641);
and U18181 (N_18181,N_17532,N_17663);
xnor U18182 (N_18182,N_17700,N_17932);
nor U18183 (N_18183,N_17876,N_17703);
xor U18184 (N_18184,N_17644,N_17632);
nand U18185 (N_18185,N_17578,N_17971);
or U18186 (N_18186,N_17731,N_17738);
or U18187 (N_18187,N_17806,N_17716);
or U18188 (N_18188,N_17697,N_17615);
nand U18189 (N_18189,N_17601,N_17925);
and U18190 (N_18190,N_17903,N_17709);
nor U18191 (N_18191,N_17872,N_17901);
and U18192 (N_18192,N_17630,N_17970);
and U18193 (N_18193,N_17734,N_17820);
xor U18194 (N_18194,N_17801,N_17812);
and U18195 (N_18195,N_17545,N_17799);
nor U18196 (N_18196,N_17927,N_17957);
nand U18197 (N_18197,N_17885,N_17688);
nand U18198 (N_18198,N_17989,N_17629);
and U18199 (N_18199,N_17610,N_17829);
nand U18200 (N_18200,N_17723,N_17984);
xor U18201 (N_18201,N_17869,N_17619);
xnor U18202 (N_18202,N_17667,N_17828);
and U18203 (N_18203,N_17564,N_17867);
and U18204 (N_18204,N_17525,N_17895);
and U18205 (N_18205,N_17669,N_17647);
nor U18206 (N_18206,N_17865,N_17816);
and U18207 (N_18207,N_17767,N_17600);
nand U18208 (N_18208,N_17673,N_17999);
or U18209 (N_18209,N_17548,N_17554);
nor U18210 (N_18210,N_17993,N_17717);
xor U18211 (N_18211,N_17768,N_17613);
xor U18212 (N_18212,N_17840,N_17506);
nand U18213 (N_18213,N_17785,N_17750);
nor U18214 (N_18214,N_17983,N_17933);
nand U18215 (N_18215,N_17888,N_17972);
nand U18216 (N_18216,N_17513,N_17842);
or U18217 (N_18217,N_17741,N_17534);
and U18218 (N_18218,N_17835,N_17706);
nor U18219 (N_18219,N_17637,N_17838);
or U18220 (N_18220,N_17643,N_17520);
and U18221 (N_18221,N_17648,N_17862);
or U18222 (N_18222,N_17789,N_17979);
nor U18223 (N_18223,N_17763,N_17718);
nand U18224 (N_18224,N_17832,N_17951);
and U18225 (N_18225,N_17661,N_17622);
nor U18226 (N_18226,N_17639,N_17570);
nor U18227 (N_18227,N_17618,N_17531);
nor U18228 (N_18228,N_17624,N_17772);
and U18229 (N_18229,N_17946,N_17656);
nor U18230 (N_18230,N_17902,N_17611);
nand U18231 (N_18231,N_17593,N_17651);
nor U18232 (N_18232,N_17590,N_17992);
nand U18233 (N_18233,N_17982,N_17945);
or U18234 (N_18234,N_17849,N_17794);
or U18235 (N_18235,N_17604,N_17539);
and U18236 (N_18236,N_17985,N_17908);
nand U18237 (N_18237,N_17671,N_17757);
nor U18238 (N_18238,N_17684,N_17952);
nand U18239 (N_18239,N_17934,N_17568);
nand U18240 (N_18240,N_17571,N_17696);
or U18241 (N_18241,N_17565,N_17808);
or U18242 (N_18242,N_17560,N_17530);
nor U18243 (N_18243,N_17963,N_17730);
and U18244 (N_18244,N_17955,N_17538);
nor U18245 (N_18245,N_17672,N_17617);
nand U18246 (N_18246,N_17834,N_17923);
nor U18247 (N_18247,N_17567,N_17636);
nor U18248 (N_18248,N_17563,N_17882);
or U18249 (N_18249,N_17890,N_17529);
or U18250 (N_18250,N_17562,N_17902);
or U18251 (N_18251,N_17918,N_17621);
nor U18252 (N_18252,N_17500,N_17571);
nor U18253 (N_18253,N_17799,N_17736);
and U18254 (N_18254,N_17867,N_17993);
and U18255 (N_18255,N_17697,N_17868);
nor U18256 (N_18256,N_17917,N_17718);
nor U18257 (N_18257,N_17762,N_17915);
and U18258 (N_18258,N_17943,N_17883);
and U18259 (N_18259,N_17941,N_17696);
xor U18260 (N_18260,N_17983,N_17919);
nor U18261 (N_18261,N_17567,N_17776);
and U18262 (N_18262,N_17671,N_17803);
nand U18263 (N_18263,N_17913,N_17692);
nand U18264 (N_18264,N_17646,N_17555);
xnor U18265 (N_18265,N_17603,N_17604);
or U18266 (N_18266,N_17977,N_17839);
nand U18267 (N_18267,N_17652,N_17782);
nor U18268 (N_18268,N_17721,N_17717);
or U18269 (N_18269,N_17911,N_17619);
or U18270 (N_18270,N_17987,N_17639);
and U18271 (N_18271,N_17742,N_17840);
nand U18272 (N_18272,N_17611,N_17883);
nor U18273 (N_18273,N_17952,N_17980);
or U18274 (N_18274,N_17687,N_17822);
or U18275 (N_18275,N_17835,N_17764);
xor U18276 (N_18276,N_17863,N_17949);
or U18277 (N_18277,N_17861,N_17985);
nand U18278 (N_18278,N_17996,N_17653);
nand U18279 (N_18279,N_17685,N_17568);
or U18280 (N_18280,N_17768,N_17807);
nand U18281 (N_18281,N_17673,N_17664);
xnor U18282 (N_18282,N_17756,N_17948);
nor U18283 (N_18283,N_17521,N_17872);
or U18284 (N_18284,N_17962,N_17683);
nor U18285 (N_18285,N_17785,N_17866);
nand U18286 (N_18286,N_17724,N_17739);
nor U18287 (N_18287,N_17543,N_17656);
nand U18288 (N_18288,N_17636,N_17776);
or U18289 (N_18289,N_17848,N_17766);
or U18290 (N_18290,N_17772,N_17982);
nand U18291 (N_18291,N_17920,N_17995);
nand U18292 (N_18292,N_17707,N_17509);
xnor U18293 (N_18293,N_17728,N_17644);
and U18294 (N_18294,N_17613,N_17843);
and U18295 (N_18295,N_17877,N_17845);
or U18296 (N_18296,N_17839,N_17993);
nand U18297 (N_18297,N_17741,N_17573);
nand U18298 (N_18298,N_17632,N_17564);
nor U18299 (N_18299,N_17705,N_17788);
nand U18300 (N_18300,N_17721,N_17842);
and U18301 (N_18301,N_17574,N_17833);
or U18302 (N_18302,N_17896,N_17747);
and U18303 (N_18303,N_17772,N_17524);
or U18304 (N_18304,N_17651,N_17523);
and U18305 (N_18305,N_17973,N_17980);
and U18306 (N_18306,N_17706,N_17522);
nor U18307 (N_18307,N_17540,N_17670);
xnor U18308 (N_18308,N_17726,N_17941);
nor U18309 (N_18309,N_17977,N_17783);
nor U18310 (N_18310,N_17764,N_17952);
and U18311 (N_18311,N_17897,N_17852);
nor U18312 (N_18312,N_17911,N_17962);
nand U18313 (N_18313,N_17841,N_17530);
nor U18314 (N_18314,N_17856,N_17514);
and U18315 (N_18315,N_17887,N_17704);
nor U18316 (N_18316,N_17672,N_17593);
nand U18317 (N_18317,N_17890,N_17630);
or U18318 (N_18318,N_17896,N_17577);
nand U18319 (N_18319,N_17905,N_17786);
or U18320 (N_18320,N_17741,N_17986);
or U18321 (N_18321,N_17662,N_17527);
or U18322 (N_18322,N_17587,N_17786);
nand U18323 (N_18323,N_17921,N_17553);
nor U18324 (N_18324,N_17506,N_17887);
nor U18325 (N_18325,N_17556,N_17842);
nor U18326 (N_18326,N_17834,N_17819);
nand U18327 (N_18327,N_17516,N_17940);
and U18328 (N_18328,N_17581,N_17688);
and U18329 (N_18329,N_17632,N_17680);
or U18330 (N_18330,N_17834,N_17584);
and U18331 (N_18331,N_17911,N_17991);
nand U18332 (N_18332,N_17906,N_17584);
nor U18333 (N_18333,N_17910,N_17916);
or U18334 (N_18334,N_17678,N_17646);
nand U18335 (N_18335,N_17968,N_17883);
nand U18336 (N_18336,N_17851,N_17534);
or U18337 (N_18337,N_17593,N_17862);
nor U18338 (N_18338,N_17896,N_17937);
xnor U18339 (N_18339,N_17805,N_17651);
nand U18340 (N_18340,N_17793,N_17912);
nor U18341 (N_18341,N_17596,N_17580);
or U18342 (N_18342,N_17985,N_17821);
nor U18343 (N_18343,N_17567,N_17708);
and U18344 (N_18344,N_17964,N_17890);
nand U18345 (N_18345,N_17538,N_17877);
nor U18346 (N_18346,N_17813,N_17849);
xnor U18347 (N_18347,N_17715,N_17974);
and U18348 (N_18348,N_17740,N_17935);
or U18349 (N_18349,N_17890,N_17916);
nor U18350 (N_18350,N_17954,N_17772);
or U18351 (N_18351,N_17731,N_17687);
and U18352 (N_18352,N_17566,N_17796);
or U18353 (N_18353,N_17866,N_17890);
and U18354 (N_18354,N_17621,N_17932);
nand U18355 (N_18355,N_17701,N_17849);
nor U18356 (N_18356,N_17551,N_17831);
and U18357 (N_18357,N_17931,N_17902);
and U18358 (N_18358,N_17803,N_17754);
or U18359 (N_18359,N_17853,N_17612);
and U18360 (N_18360,N_17616,N_17845);
and U18361 (N_18361,N_17717,N_17975);
nand U18362 (N_18362,N_17746,N_17531);
nand U18363 (N_18363,N_17818,N_17676);
and U18364 (N_18364,N_17691,N_17984);
nor U18365 (N_18365,N_17652,N_17767);
nand U18366 (N_18366,N_17993,N_17923);
xnor U18367 (N_18367,N_17664,N_17894);
or U18368 (N_18368,N_17992,N_17836);
nor U18369 (N_18369,N_17835,N_17581);
nor U18370 (N_18370,N_17992,N_17722);
or U18371 (N_18371,N_17593,N_17966);
nand U18372 (N_18372,N_17765,N_17825);
and U18373 (N_18373,N_17552,N_17922);
or U18374 (N_18374,N_17622,N_17730);
nor U18375 (N_18375,N_17707,N_17555);
or U18376 (N_18376,N_17693,N_17633);
or U18377 (N_18377,N_17573,N_17570);
nor U18378 (N_18378,N_17891,N_17819);
nand U18379 (N_18379,N_17784,N_17502);
and U18380 (N_18380,N_17571,N_17572);
nand U18381 (N_18381,N_17798,N_17771);
nor U18382 (N_18382,N_17878,N_17960);
or U18383 (N_18383,N_17931,N_17531);
nor U18384 (N_18384,N_17815,N_17573);
nand U18385 (N_18385,N_17846,N_17623);
nor U18386 (N_18386,N_17842,N_17580);
xor U18387 (N_18387,N_17805,N_17925);
nand U18388 (N_18388,N_17965,N_17779);
nand U18389 (N_18389,N_17717,N_17961);
and U18390 (N_18390,N_17968,N_17537);
nor U18391 (N_18391,N_17960,N_17595);
and U18392 (N_18392,N_17938,N_17991);
nand U18393 (N_18393,N_17774,N_17691);
xor U18394 (N_18394,N_17619,N_17757);
nor U18395 (N_18395,N_17602,N_17630);
nand U18396 (N_18396,N_17789,N_17961);
nor U18397 (N_18397,N_17991,N_17948);
nor U18398 (N_18398,N_17622,N_17974);
and U18399 (N_18399,N_17854,N_17805);
xnor U18400 (N_18400,N_17769,N_17568);
nor U18401 (N_18401,N_17646,N_17521);
nor U18402 (N_18402,N_17989,N_17557);
and U18403 (N_18403,N_17929,N_17999);
and U18404 (N_18404,N_17826,N_17641);
or U18405 (N_18405,N_17878,N_17552);
nor U18406 (N_18406,N_17566,N_17901);
and U18407 (N_18407,N_17571,N_17574);
and U18408 (N_18408,N_17528,N_17621);
or U18409 (N_18409,N_17884,N_17686);
nand U18410 (N_18410,N_17686,N_17711);
or U18411 (N_18411,N_17538,N_17861);
or U18412 (N_18412,N_17998,N_17777);
xor U18413 (N_18413,N_17704,N_17749);
nand U18414 (N_18414,N_17956,N_17913);
nand U18415 (N_18415,N_17805,N_17981);
and U18416 (N_18416,N_17881,N_17626);
nand U18417 (N_18417,N_17952,N_17645);
nor U18418 (N_18418,N_17572,N_17747);
nand U18419 (N_18419,N_17601,N_17818);
and U18420 (N_18420,N_17534,N_17818);
or U18421 (N_18421,N_17751,N_17901);
nor U18422 (N_18422,N_17974,N_17511);
nor U18423 (N_18423,N_17591,N_17704);
nand U18424 (N_18424,N_17593,N_17980);
or U18425 (N_18425,N_17599,N_17622);
and U18426 (N_18426,N_17649,N_17959);
and U18427 (N_18427,N_17831,N_17564);
nand U18428 (N_18428,N_17624,N_17840);
or U18429 (N_18429,N_17950,N_17805);
nor U18430 (N_18430,N_17766,N_17974);
or U18431 (N_18431,N_17668,N_17760);
nor U18432 (N_18432,N_17917,N_17929);
and U18433 (N_18433,N_17506,N_17760);
xnor U18434 (N_18434,N_17652,N_17754);
nor U18435 (N_18435,N_17844,N_17921);
nand U18436 (N_18436,N_17843,N_17676);
or U18437 (N_18437,N_17563,N_17847);
or U18438 (N_18438,N_17966,N_17764);
or U18439 (N_18439,N_17721,N_17747);
nand U18440 (N_18440,N_17517,N_17588);
nor U18441 (N_18441,N_17787,N_17769);
or U18442 (N_18442,N_17784,N_17807);
and U18443 (N_18443,N_17649,N_17609);
nand U18444 (N_18444,N_17930,N_17568);
nor U18445 (N_18445,N_17511,N_17993);
nand U18446 (N_18446,N_17758,N_17703);
or U18447 (N_18447,N_17814,N_17770);
nor U18448 (N_18448,N_17642,N_17816);
nor U18449 (N_18449,N_17833,N_17566);
nor U18450 (N_18450,N_17883,N_17516);
nor U18451 (N_18451,N_17816,N_17519);
xnor U18452 (N_18452,N_17648,N_17795);
nor U18453 (N_18453,N_17935,N_17529);
nand U18454 (N_18454,N_17707,N_17610);
xor U18455 (N_18455,N_17692,N_17995);
and U18456 (N_18456,N_17656,N_17515);
or U18457 (N_18457,N_17578,N_17540);
or U18458 (N_18458,N_17908,N_17837);
or U18459 (N_18459,N_17946,N_17753);
or U18460 (N_18460,N_17681,N_17614);
nor U18461 (N_18461,N_17597,N_17853);
xor U18462 (N_18462,N_17591,N_17612);
and U18463 (N_18463,N_17937,N_17872);
nor U18464 (N_18464,N_17959,N_17547);
nor U18465 (N_18465,N_17860,N_17693);
or U18466 (N_18466,N_17605,N_17786);
and U18467 (N_18467,N_17812,N_17961);
or U18468 (N_18468,N_17878,N_17510);
nor U18469 (N_18469,N_17559,N_17615);
nor U18470 (N_18470,N_17880,N_17984);
nor U18471 (N_18471,N_17997,N_17645);
nor U18472 (N_18472,N_17778,N_17801);
and U18473 (N_18473,N_17688,N_17848);
and U18474 (N_18474,N_17799,N_17800);
and U18475 (N_18475,N_17643,N_17814);
nor U18476 (N_18476,N_17776,N_17954);
nor U18477 (N_18477,N_17939,N_17590);
and U18478 (N_18478,N_17819,N_17805);
nor U18479 (N_18479,N_17691,N_17508);
nor U18480 (N_18480,N_17835,N_17838);
or U18481 (N_18481,N_17829,N_17934);
nand U18482 (N_18482,N_17907,N_17883);
or U18483 (N_18483,N_17703,N_17866);
nor U18484 (N_18484,N_17739,N_17610);
and U18485 (N_18485,N_17955,N_17519);
nand U18486 (N_18486,N_17715,N_17681);
nand U18487 (N_18487,N_17649,N_17960);
and U18488 (N_18488,N_17770,N_17754);
and U18489 (N_18489,N_17716,N_17614);
nand U18490 (N_18490,N_17555,N_17610);
nor U18491 (N_18491,N_17596,N_17956);
and U18492 (N_18492,N_17774,N_17616);
nor U18493 (N_18493,N_17706,N_17971);
nor U18494 (N_18494,N_17520,N_17702);
and U18495 (N_18495,N_17737,N_17883);
nor U18496 (N_18496,N_17561,N_17898);
or U18497 (N_18497,N_17860,N_17925);
nor U18498 (N_18498,N_17935,N_17799);
and U18499 (N_18499,N_17709,N_17586);
xnor U18500 (N_18500,N_18138,N_18449);
nand U18501 (N_18501,N_18110,N_18048);
nor U18502 (N_18502,N_18257,N_18098);
nand U18503 (N_18503,N_18192,N_18134);
xor U18504 (N_18504,N_18441,N_18456);
nor U18505 (N_18505,N_18323,N_18428);
and U18506 (N_18506,N_18238,N_18084);
nand U18507 (N_18507,N_18468,N_18370);
or U18508 (N_18508,N_18438,N_18211);
nor U18509 (N_18509,N_18044,N_18345);
xor U18510 (N_18510,N_18260,N_18436);
xnor U18511 (N_18511,N_18107,N_18418);
or U18512 (N_18512,N_18445,N_18161);
or U18513 (N_18513,N_18207,N_18312);
xnor U18514 (N_18514,N_18025,N_18489);
nand U18515 (N_18515,N_18473,N_18400);
or U18516 (N_18516,N_18195,N_18158);
and U18517 (N_18517,N_18146,N_18319);
xor U18518 (N_18518,N_18349,N_18163);
and U18519 (N_18519,N_18232,N_18014);
nand U18520 (N_18520,N_18381,N_18378);
or U18521 (N_18521,N_18470,N_18407);
nor U18522 (N_18522,N_18000,N_18113);
and U18523 (N_18523,N_18275,N_18149);
nor U18524 (N_18524,N_18205,N_18451);
nand U18525 (N_18525,N_18471,N_18300);
and U18526 (N_18526,N_18487,N_18332);
and U18527 (N_18527,N_18486,N_18437);
or U18528 (N_18528,N_18402,N_18208);
and U18529 (N_18529,N_18347,N_18039);
nand U18530 (N_18530,N_18484,N_18085);
or U18531 (N_18531,N_18005,N_18037);
xor U18532 (N_18532,N_18157,N_18492);
xor U18533 (N_18533,N_18322,N_18448);
or U18534 (N_18534,N_18364,N_18129);
xor U18535 (N_18535,N_18169,N_18118);
nor U18536 (N_18536,N_18054,N_18333);
and U18537 (N_18537,N_18384,N_18212);
nand U18538 (N_18538,N_18201,N_18204);
nand U18539 (N_18539,N_18066,N_18411);
nor U18540 (N_18540,N_18461,N_18019);
and U18541 (N_18541,N_18287,N_18472);
and U18542 (N_18542,N_18171,N_18308);
xor U18543 (N_18543,N_18071,N_18038);
nor U18544 (N_18544,N_18479,N_18123);
nand U18545 (N_18545,N_18168,N_18498);
xor U18546 (N_18546,N_18227,N_18064);
xor U18547 (N_18547,N_18453,N_18174);
nor U18548 (N_18548,N_18213,N_18467);
or U18549 (N_18549,N_18435,N_18070);
or U18550 (N_18550,N_18077,N_18193);
or U18551 (N_18551,N_18454,N_18065);
and U18552 (N_18552,N_18477,N_18111);
xnor U18553 (N_18553,N_18108,N_18268);
and U18554 (N_18554,N_18305,N_18124);
and U18555 (N_18555,N_18288,N_18112);
nand U18556 (N_18556,N_18426,N_18190);
and U18557 (N_18557,N_18075,N_18463);
nand U18558 (N_18558,N_18166,N_18221);
or U18559 (N_18559,N_18097,N_18156);
xnor U18560 (N_18560,N_18151,N_18313);
nor U18561 (N_18561,N_18068,N_18442);
nor U18562 (N_18562,N_18120,N_18177);
nand U18563 (N_18563,N_18363,N_18337);
and U18564 (N_18564,N_18405,N_18013);
and U18565 (N_18565,N_18234,N_18051);
or U18566 (N_18566,N_18175,N_18230);
nor U18567 (N_18567,N_18224,N_18457);
nor U18568 (N_18568,N_18385,N_18377);
or U18569 (N_18569,N_18248,N_18282);
nor U18570 (N_18570,N_18096,N_18395);
nand U18571 (N_18571,N_18277,N_18080);
or U18572 (N_18572,N_18247,N_18359);
and U18573 (N_18573,N_18041,N_18433);
nor U18574 (N_18574,N_18316,N_18246);
nand U18575 (N_18575,N_18458,N_18443);
nand U18576 (N_18576,N_18186,N_18189);
nor U18577 (N_18577,N_18339,N_18392);
or U18578 (N_18578,N_18265,N_18306);
xnor U18579 (N_18579,N_18088,N_18132);
nor U18580 (N_18580,N_18434,N_18202);
nor U18581 (N_18581,N_18105,N_18485);
and U18582 (N_18582,N_18002,N_18091);
nor U18583 (N_18583,N_18294,N_18376);
nand U18584 (N_18584,N_18496,N_18272);
nor U18585 (N_18585,N_18330,N_18021);
or U18586 (N_18586,N_18259,N_18444);
nand U18587 (N_18587,N_18226,N_18148);
nand U18588 (N_18588,N_18061,N_18301);
and U18589 (N_18589,N_18328,N_18320);
and U18590 (N_18590,N_18015,N_18131);
or U18591 (N_18591,N_18136,N_18035);
nand U18592 (N_18592,N_18455,N_18087);
and U18593 (N_18593,N_18340,N_18373);
or U18594 (N_18594,N_18414,N_18030);
and U18595 (N_18595,N_18165,N_18254);
or U18596 (N_18596,N_18170,N_18424);
nor U18597 (N_18597,N_18004,N_18310);
nand U18598 (N_18598,N_18043,N_18069);
or U18599 (N_18599,N_18490,N_18210);
and U18600 (N_18600,N_18459,N_18020);
nand U18601 (N_18601,N_18263,N_18278);
nor U18602 (N_18602,N_18033,N_18046);
or U18603 (N_18603,N_18432,N_18241);
and U18604 (N_18604,N_18140,N_18209);
and U18605 (N_18605,N_18419,N_18375);
and U18606 (N_18606,N_18430,N_18056);
or U18607 (N_18607,N_18235,N_18067);
nor U18608 (N_18608,N_18203,N_18142);
nand U18609 (N_18609,N_18012,N_18267);
nor U18610 (N_18610,N_18233,N_18253);
and U18611 (N_18611,N_18160,N_18427);
nor U18612 (N_18612,N_18052,N_18130);
and U18613 (N_18613,N_18144,N_18476);
nand U18614 (N_18614,N_18409,N_18079);
nand U18615 (N_18615,N_18104,N_18355);
and U18616 (N_18616,N_18040,N_18094);
and U18617 (N_18617,N_18351,N_18284);
nand U18618 (N_18618,N_18296,N_18317);
xnor U18619 (N_18619,N_18172,N_18314);
nor U18620 (N_18620,N_18245,N_18318);
nand U18621 (N_18621,N_18255,N_18388);
and U18622 (N_18622,N_18362,N_18249);
nor U18623 (N_18623,N_18464,N_18406);
nor U18624 (N_18624,N_18081,N_18421);
nor U18625 (N_18625,N_18483,N_18493);
and U18626 (N_18626,N_18011,N_18450);
or U18627 (N_18627,N_18133,N_18336);
nor U18628 (N_18628,N_18028,N_18236);
nor U18629 (N_18629,N_18354,N_18393);
nand U18630 (N_18630,N_18223,N_18394);
xor U18631 (N_18631,N_18237,N_18326);
nand U18632 (N_18632,N_18214,N_18127);
or U18633 (N_18633,N_18374,N_18194);
nor U18634 (N_18634,N_18341,N_18481);
xnor U18635 (N_18635,N_18198,N_18076);
and U18636 (N_18636,N_18285,N_18488);
nor U18637 (N_18637,N_18145,N_18217);
nand U18638 (N_18638,N_18178,N_18184);
and U18639 (N_18639,N_18474,N_18008);
nand U18640 (N_18640,N_18162,N_18290);
or U18641 (N_18641,N_18122,N_18420);
and U18642 (N_18642,N_18003,N_18431);
and U18643 (N_18643,N_18439,N_18007);
and U18644 (N_18644,N_18425,N_18137);
and U18645 (N_18645,N_18446,N_18159);
nand U18646 (N_18646,N_18386,N_18225);
nand U18647 (N_18647,N_18495,N_18229);
nand U18648 (N_18648,N_18219,N_18293);
or U18649 (N_18649,N_18042,N_18115);
xnor U18650 (N_18650,N_18244,N_18475);
or U18651 (N_18651,N_18185,N_18228);
xnor U18652 (N_18652,N_18415,N_18073);
or U18653 (N_18653,N_18422,N_18327);
nor U18654 (N_18654,N_18390,N_18022);
and U18655 (N_18655,N_18191,N_18139);
nor U18656 (N_18656,N_18478,N_18089);
or U18657 (N_18657,N_18009,N_18303);
xor U18658 (N_18658,N_18252,N_18371);
nand U18659 (N_18659,N_18251,N_18155);
and U18660 (N_18660,N_18126,N_18135);
and U18661 (N_18661,N_18304,N_18017);
and U18662 (N_18662,N_18215,N_18365);
and U18663 (N_18663,N_18216,N_18462);
nor U18664 (N_18664,N_18466,N_18083);
or U18665 (N_18665,N_18403,N_18297);
and U18666 (N_18666,N_18200,N_18045);
nor U18667 (N_18667,N_18413,N_18095);
or U18668 (N_18668,N_18482,N_18398);
or U18669 (N_18669,N_18289,N_18270);
and U18670 (N_18670,N_18173,N_18325);
nor U18671 (N_18671,N_18469,N_18024);
nand U18672 (N_18672,N_18429,N_18497);
and U18673 (N_18673,N_18334,N_18360);
and U18674 (N_18674,N_18206,N_18006);
nor U18675 (N_18675,N_18114,N_18342);
xor U18676 (N_18676,N_18276,N_18382);
xor U18677 (N_18677,N_18197,N_18343);
nor U18678 (N_18678,N_18179,N_18396);
or U18679 (N_18679,N_18016,N_18027);
and U18680 (N_18680,N_18283,N_18250);
nand U18681 (N_18681,N_18460,N_18292);
or U18682 (N_18682,N_18367,N_18366);
xor U18683 (N_18683,N_18356,N_18182);
nand U18684 (N_18684,N_18344,N_18417);
and U18685 (N_18685,N_18026,N_18147);
nor U18686 (N_18686,N_18031,N_18404);
nor U18687 (N_18687,N_18264,N_18032);
or U18688 (N_18688,N_18324,N_18286);
nor U18689 (N_18689,N_18412,N_18329);
xnor U18690 (N_18690,N_18291,N_18047);
nor U18691 (N_18691,N_18180,N_18188);
nor U18692 (N_18692,N_18102,N_18401);
and U18693 (N_18693,N_18167,N_18196);
xor U18694 (N_18694,N_18299,N_18408);
nor U18695 (N_18695,N_18266,N_18302);
nand U18696 (N_18696,N_18239,N_18380);
nor U18697 (N_18697,N_18348,N_18057);
or U18698 (N_18698,N_18036,N_18049);
nor U18699 (N_18699,N_18361,N_18358);
and U18700 (N_18700,N_18452,N_18387);
nor U18701 (N_18701,N_18335,N_18141);
nand U18702 (N_18702,N_18372,N_18256);
nor U18703 (N_18703,N_18109,N_18199);
or U18704 (N_18704,N_18357,N_18222);
nor U18705 (N_18705,N_18092,N_18295);
nor U18706 (N_18706,N_18331,N_18010);
or U18707 (N_18707,N_18074,N_18240);
nand U18708 (N_18708,N_18100,N_18261);
nor U18709 (N_18709,N_18298,N_18116);
nor U18710 (N_18710,N_18218,N_18279);
or U18711 (N_18711,N_18082,N_18050);
and U18712 (N_18712,N_18242,N_18018);
nor U18713 (N_18713,N_18311,N_18399);
or U18714 (N_18714,N_18423,N_18383);
and U18715 (N_18715,N_18280,N_18154);
nand U18716 (N_18716,N_18389,N_18125);
nand U18717 (N_18717,N_18090,N_18119);
or U18718 (N_18718,N_18063,N_18465);
nor U18719 (N_18719,N_18183,N_18499);
xnor U18720 (N_18720,N_18164,N_18128);
nand U18721 (N_18721,N_18315,N_18099);
or U18722 (N_18722,N_18101,N_18062);
and U18723 (N_18723,N_18143,N_18258);
or U18724 (N_18724,N_18023,N_18397);
or U18725 (N_18725,N_18034,N_18369);
nor U18726 (N_18726,N_18153,N_18309);
nor U18727 (N_18727,N_18281,N_18346);
and U18728 (N_18728,N_18072,N_18350);
nand U18729 (N_18729,N_18447,N_18053);
nor U18730 (N_18730,N_18121,N_18181);
nand U18731 (N_18731,N_18220,N_18078);
nand U18732 (N_18732,N_18103,N_18106);
xnor U18733 (N_18733,N_18001,N_18416);
nor U18734 (N_18734,N_18086,N_18269);
and U18735 (N_18735,N_18480,N_18440);
and U18736 (N_18736,N_18058,N_18262);
or U18737 (N_18737,N_18353,N_18410);
nor U18738 (N_18738,N_18152,N_18117);
and U18739 (N_18739,N_18176,N_18274);
xnor U18740 (N_18740,N_18338,N_18491);
nand U18741 (N_18741,N_18273,N_18271);
nor U18742 (N_18742,N_18060,N_18321);
nor U18743 (N_18743,N_18093,N_18352);
xnor U18744 (N_18744,N_18231,N_18391);
nand U18745 (N_18745,N_18494,N_18243);
nor U18746 (N_18746,N_18187,N_18150);
nand U18747 (N_18747,N_18029,N_18059);
or U18748 (N_18748,N_18379,N_18055);
and U18749 (N_18749,N_18368,N_18307);
nor U18750 (N_18750,N_18435,N_18259);
or U18751 (N_18751,N_18298,N_18205);
and U18752 (N_18752,N_18037,N_18130);
nand U18753 (N_18753,N_18476,N_18184);
and U18754 (N_18754,N_18294,N_18477);
and U18755 (N_18755,N_18372,N_18398);
and U18756 (N_18756,N_18289,N_18133);
or U18757 (N_18757,N_18067,N_18232);
nand U18758 (N_18758,N_18015,N_18428);
nor U18759 (N_18759,N_18358,N_18330);
xnor U18760 (N_18760,N_18329,N_18378);
nand U18761 (N_18761,N_18329,N_18073);
nand U18762 (N_18762,N_18135,N_18128);
xnor U18763 (N_18763,N_18304,N_18387);
and U18764 (N_18764,N_18326,N_18459);
xnor U18765 (N_18765,N_18203,N_18000);
xor U18766 (N_18766,N_18045,N_18419);
nand U18767 (N_18767,N_18317,N_18342);
nor U18768 (N_18768,N_18150,N_18239);
nor U18769 (N_18769,N_18497,N_18072);
nor U18770 (N_18770,N_18069,N_18328);
xnor U18771 (N_18771,N_18159,N_18137);
or U18772 (N_18772,N_18177,N_18270);
xor U18773 (N_18773,N_18389,N_18321);
nand U18774 (N_18774,N_18321,N_18209);
and U18775 (N_18775,N_18289,N_18397);
and U18776 (N_18776,N_18278,N_18038);
nor U18777 (N_18777,N_18336,N_18382);
nand U18778 (N_18778,N_18341,N_18059);
nor U18779 (N_18779,N_18456,N_18499);
nand U18780 (N_18780,N_18145,N_18311);
nand U18781 (N_18781,N_18082,N_18023);
and U18782 (N_18782,N_18179,N_18251);
nor U18783 (N_18783,N_18126,N_18366);
nor U18784 (N_18784,N_18499,N_18383);
nand U18785 (N_18785,N_18053,N_18343);
nor U18786 (N_18786,N_18470,N_18126);
or U18787 (N_18787,N_18351,N_18477);
xor U18788 (N_18788,N_18287,N_18048);
nor U18789 (N_18789,N_18408,N_18415);
nor U18790 (N_18790,N_18186,N_18150);
and U18791 (N_18791,N_18266,N_18455);
nor U18792 (N_18792,N_18162,N_18024);
nand U18793 (N_18793,N_18446,N_18197);
and U18794 (N_18794,N_18338,N_18327);
and U18795 (N_18795,N_18408,N_18460);
nor U18796 (N_18796,N_18079,N_18386);
and U18797 (N_18797,N_18282,N_18018);
xor U18798 (N_18798,N_18420,N_18341);
or U18799 (N_18799,N_18330,N_18281);
nand U18800 (N_18800,N_18151,N_18257);
xnor U18801 (N_18801,N_18358,N_18402);
nand U18802 (N_18802,N_18421,N_18404);
or U18803 (N_18803,N_18494,N_18009);
nor U18804 (N_18804,N_18153,N_18026);
and U18805 (N_18805,N_18483,N_18143);
and U18806 (N_18806,N_18492,N_18242);
nor U18807 (N_18807,N_18306,N_18159);
and U18808 (N_18808,N_18175,N_18336);
or U18809 (N_18809,N_18356,N_18457);
and U18810 (N_18810,N_18478,N_18180);
nor U18811 (N_18811,N_18360,N_18149);
nor U18812 (N_18812,N_18191,N_18265);
nand U18813 (N_18813,N_18139,N_18098);
or U18814 (N_18814,N_18421,N_18013);
nand U18815 (N_18815,N_18450,N_18309);
or U18816 (N_18816,N_18454,N_18211);
xor U18817 (N_18817,N_18310,N_18320);
and U18818 (N_18818,N_18138,N_18033);
and U18819 (N_18819,N_18337,N_18488);
or U18820 (N_18820,N_18073,N_18348);
nand U18821 (N_18821,N_18154,N_18011);
nand U18822 (N_18822,N_18204,N_18267);
or U18823 (N_18823,N_18002,N_18206);
nor U18824 (N_18824,N_18282,N_18016);
or U18825 (N_18825,N_18126,N_18039);
nand U18826 (N_18826,N_18095,N_18190);
nand U18827 (N_18827,N_18044,N_18385);
nor U18828 (N_18828,N_18442,N_18413);
or U18829 (N_18829,N_18104,N_18029);
and U18830 (N_18830,N_18148,N_18483);
and U18831 (N_18831,N_18108,N_18485);
and U18832 (N_18832,N_18013,N_18392);
nand U18833 (N_18833,N_18280,N_18283);
nor U18834 (N_18834,N_18086,N_18489);
or U18835 (N_18835,N_18212,N_18362);
xor U18836 (N_18836,N_18421,N_18157);
or U18837 (N_18837,N_18069,N_18166);
nor U18838 (N_18838,N_18380,N_18278);
and U18839 (N_18839,N_18453,N_18244);
nand U18840 (N_18840,N_18141,N_18253);
nor U18841 (N_18841,N_18380,N_18154);
xor U18842 (N_18842,N_18051,N_18069);
or U18843 (N_18843,N_18334,N_18486);
or U18844 (N_18844,N_18244,N_18396);
nand U18845 (N_18845,N_18468,N_18291);
nor U18846 (N_18846,N_18124,N_18199);
and U18847 (N_18847,N_18137,N_18028);
nor U18848 (N_18848,N_18213,N_18393);
nand U18849 (N_18849,N_18455,N_18145);
nor U18850 (N_18850,N_18346,N_18350);
xnor U18851 (N_18851,N_18071,N_18338);
or U18852 (N_18852,N_18090,N_18380);
xnor U18853 (N_18853,N_18104,N_18351);
and U18854 (N_18854,N_18130,N_18332);
and U18855 (N_18855,N_18173,N_18228);
nand U18856 (N_18856,N_18450,N_18238);
nor U18857 (N_18857,N_18269,N_18262);
nand U18858 (N_18858,N_18476,N_18056);
and U18859 (N_18859,N_18169,N_18051);
nand U18860 (N_18860,N_18286,N_18054);
and U18861 (N_18861,N_18322,N_18252);
nor U18862 (N_18862,N_18223,N_18464);
xor U18863 (N_18863,N_18240,N_18254);
nor U18864 (N_18864,N_18427,N_18102);
nor U18865 (N_18865,N_18402,N_18347);
or U18866 (N_18866,N_18329,N_18067);
nor U18867 (N_18867,N_18427,N_18305);
or U18868 (N_18868,N_18351,N_18415);
and U18869 (N_18869,N_18292,N_18220);
and U18870 (N_18870,N_18248,N_18144);
nor U18871 (N_18871,N_18168,N_18071);
nor U18872 (N_18872,N_18370,N_18355);
nand U18873 (N_18873,N_18078,N_18156);
nand U18874 (N_18874,N_18313,N_18055);
nor U18875 (N_18875,N_18231,N_18129);
or U18876 (N_18876,N_18227,N_18020);
and U18877 (N_18877,N_18304,N_18375);
nand U18878 (N_18878,N_18400,N_18186);
nand U18879 (N_18879,N_18255,N_18494);
nand U18880 (N_18880,N_18108,N_18049);
nand U18881 (N_18881,N_18065,N_18271);
or U18882 (N_18882,N_18185,N_18251);
xor U18883 (N_18883,N_18280,N_18458);
xnor U18884 (N_18884,N_18158,N_18080);
xor U18885 (N_18885,N_18429,N_18259);
nor U18886 (N_18886,N_18348,N_18120);
nand U18887 (N_18887,N_18059,N_18352);
nor U18888 (N_18888,N_18057,N_18012);
or U18889 (N_18889,N_18483,N_18262);
or U18890 (N_18890,N_18139,N_18094);
xnor U18891 (N_18891,N_18119,N_18009);
nand U18892 (N_18892,N_18358,N_18074);
nor U18893 (N_18893,N_18491,N_18379);
nor U18894 (N_18894,N_18354,N_18446);
and U18895 (N_18895,N_18295,N_18472);
nand U18896 (N_18896,N_18365,N_18307);
nand U18897 (N_18897,N_18404,N_18064);
or U18898 (N_18898,N_18494,N_18399);
xor U18899 (N_18899,N_18450,N_18024);
or U18900 (N_18900,N_18106,N_18135);
xnor U18901 (N_18901,N_18423,N_18030);
nand U18902 (N_18902,N_18067,N_18043);
nand U18903 (N_18903,N_18269,N_18255);
nor U18904 (N_18904,N_18159,N_18268);
or U18905 (N_18905,N_18441,N_18323);
and U18906 (N_18906,N_18233,N_18194);
nor U18907 (N_18907,N_18240,N_18416);
and U18908 (N_18908,N_18031,N_18419);
nand U18909 (N_18909,N_18232,N_18214);
nand U18910 (N_18910,N_18132,N_18345);
nor U18911 (N_18911,N_18390,N_18047);
and U18912 (N_18912,N_18296,N_18204);
or U18913 (N_18913,N_18028,N_18372);
or U18914 (N_18914,N_18018,N_18233);
nor U18915 (N_18915,N_18128,N_18461);
xor U18916 (N_18916,N_18417,N_18395);
and U18917 (N_18917,N_18261,N_18294);
nand U18918 (N_18918,N_18207,N_18344);
or U18919 (N_18919,N_18256,N_18453);
or U18920 (N_18920,N_18231,N_18277);
and U18921 (N_18921,N_18061,N_18202);
or U18922 (N_18922,N_18081,N_18071);
and U18923 (N_18923,N_18342,N_18119);
and U18924 (N_18924,N_18169,N_18376);
or U18925 (N_18925,N_18178,N_18221);
and U18926 (N_18926,N_18031,N_18117);
and U18927 (N_18927,N_18358,N_18065);
nand U18928 (N_18928,N_18229,N_18226);
nor U18929 (N_18929,N_18128,N_18217);
or U18930 (N_18930,N_18091,N_18429);
and U18931 (N_18931,N_18224,N_18407);
nand U18932 (N_18932,N_18295,N_18288);
nor U18933 (N_18933,N_18410,N_18036);
nand U18934 (N_18934,N_18255,N_18387);
nand U18935 (N_18935,N_18292,N_18285);
and U18936 (N_18936,N_18060,N_18346);
or U18937 (N_18937,N_18064,N_18224);
nor U18938 (N_18938,N_18072,N_18468);
xor U18939 (N_18939,N_18340,N_18220);
nor U18940 (N_18940,N_18424,N_18200);
nor U18941 (N_18941,N_18323,N_18158);
or U18942 (N_18942,N_18499,N_18344);
or U18943 (N_18943,N_18172,N_18164);
or U18944 (N_18944,N_18075,N_18440);
nand U18945 (N_18945,N_18161,N_18489);
nor U18946 (N_18946,N_18124,N_18033);
nor U18947 (N_18947,N_18143,N_18486);
nor U18948 (N_18948,N_18359,N_18182);
nor U18949 (N_18949,N_18153,N_18160);
nor U18950 (N_18950,N_18410,N_18417);
or U18951 (N_18951,N_18153,N_18401);
or U18952 (N_18952,N_18490,N_18306);
or U18953 (N_18953,N_18126,N_18004);
or U18954 (N_18954,N_18005,N_18413);
nand U18955 (N_18955,N_18461,N_18111);
or U18956 (N_18956,N_18335,N_18049);
or U18957 (N_18957,N_18492,N_18090);
xor U18958 (N_18958,N_18166,N_18019);
nand U18959 (N_18959,N_18279,N_18416);
nand U18960 (N_18960,N_18018,N_18452);
and U18961 (N_18961,N_18265,N_18037);
xor U18962 (N_18962,N_18020,N_18280);
and U18963 (N_18963,N_18454,N_18477);
xnor U18964 (N_18964,N_18183,N_18355);
and U18965 (N_18965,N_18404,N_18296);
nor U18966 (N_18966,N_18224,N_18031);
nor U18967 (N_18967,N_18200,N_18020);
nor U18968 (N_18968,N_18265,N_18307);
nor U18969 (N_18969,N_18199,N_18325);
nand U18970 (N_18970,N_18257,N_18072);
nand U18971 (N_18971,N_18168,N_18070);
nand U18972 (N_18972,N_18158,N_18398);
nand U18973 (N_18973,N_18155,N_18158);
nor U18974 (N_18974,N_18145,N_18281);
xor U18975 (N_18975,N_18378,N_18258);
or U18976 (N_18976,N_18095,N_18223);
and U18977 (N_18977,N_18361,N_18403);
and U18978 (N_18978,N_18119,N_18196);
or U18979 (N_18979,N_18074,N_18121);
and U18980 (N_18980,N_18036,N_18382);
or U18981 (N_18981,N_18376,N_18385);
and U18982 (N_18982,N_18371,N_18001);
nor U18983 (N_18983,N_18106,N_18410);
nor U18984 (N_18984,N_18057,N_18425);
and U18985 (N_18985,N_18222,N_18405);
or U18986 (N_18986,N_18202,N_18371);
nor U18987 (N_18987,N_18195,N_18016);
and U18988 (N_18988,N_18334,N_18344);
nor U18989 (N_18989,N_18245,N_18023);
and U18990 (N_18990,N_18125,N_18419);
or U18991 (N_18991,N_18483,N_18233);
and U18992 (N_18992,N_18499,N_18384);
xor U18993 (N_18993,N_18216,N_18294);
nor U18994 (N_18994,N_18390,N_18066);
or U18995 (N_18995,N_18354,N_18440);
nand U18996 (N_18996,N_18459,N_18464);
nand U18997 (N_18997,N_18474,N_18152);
xor U18998 (N_18998,N_18261,N_18000);
or U18999 (N_18999,N_18185,N_18372);
or U19000 (N_19000,N_18510,N_18728);
nand U19001 (N_19001,N_18910,N_18756);
nand U19002 (N_19002,N_18864,N_18852);
nand U19003 (N_19003,N_18558,N_18945);
and U19004 (N_19004,N_18940,N_18969);
and U19005 (N_19005,N_18554,N_18995);
or U19006 (N_19006,N_18622,N_18530);
nor U19007 (N_19007,N_18790,N_18529);
or U19008 (N_19008,N_18961,N_18538);
and U19009 (N_19009,N_18597,N_18572);
xnor U19010 (N_19010,N_18600,N_18641);
nand U19011 (N_19011,N_18994,N_18602);
nand U19012 (N_19012,N_18652,N_18761);
or U19013 (N_19013,N_18577,N_18640);
and U19014 (N_19014,N_18953,N_18542);
xor U19015 (N_19015,N_18585,N_18501);
nor U19016 (N_19016,N_18804,N_18786);
nand U19017 (N_19017,N_18776,N_18773);
xor U19018 (N_19018,N_18755,N_18942);
or U19019 (N_19019,N_18660,N_18527);
and U19020 (N_19020,N_18877,N_18788);
or U19021 (N_19021,N_18923,N_18734);
and U19022 (N_19022,N_18573,N_18733);
or U19023 (N_19023,N_18828,N_18789);
and U19024 (N_19024,N_18524,N_18943);
or U19025 (N_19025,N_18853,N_18717);
or U19026 (N_19026,N_18679,N_18875);
or U19027 (N_19027,N_18889,N_18837);
and U19028 (N_19028,N_18520,N_18534);
xnor U19029 (N_19029,N_18675,N_18583);
or U19030 (N_19030,N_18997,N_18691);
or U19031 (N_19031,N_18902,N_18627);
nand U19032 (N_19032,N_18601,N_18673);
nor U19033 (N_19033,N_18535,N_18898);
nand U19034 (N_19034,N_18962,N_18765);
xnor U19035 (N_19035,N_18590,N_18979);
and U19036 (N_19036,N_18854,N_18836);
nand U19037 (N_19037,N_18539,N_18571);
or U19038 (N_19038,N_18505,N_18745);
and U19039 (N_19039,N_18832,N_18705);
xor U19040 (N_19040,N_18649,N_18952);
and U19041 (N_19041,N_18643,N_18716);
nand U19042 (N_19042,N_18664,N_18680);
nand U19043 (N_19043,N_18906,N_18785);
nor U19044 (N_19044,N_18620,N_18744);
or U19045 (N_19045,N_18688,N_18835);
or U19046 (N_19046,N_18687,N_18516);
or U19047 (N_19047,N_18668,N_18706);
and U19048 (N_19048,N_18816,N_18781);
nand U19049 (N_19049,N_18580,N_18509);
and U19050 (N_19050,N_18960,N_18967);
and U19051 (N_19051,N_18644,N_18713);
and U19052 (N_19052,N_18915,N_18747);
xor U19053 (N_19053,N_18676,N_18711);
nor U19054 (N_19054,N_18857,N_18946);
xnor U19055 (N_19055,N_18657,N_18849);
or U19056 (N_19056,N_18861,N_18596);
or U19057 (N_19057,N_18515,N_18900);
and U19058 (N_19058,N_18896,N_18665);
or U19059 (N_19059,N_18645,N_18720);
nor U19060 (N_19060,N_18503,N_18586);
nand U19061 (N_19061,N_18842,N_18653);
and U19062 (N_19062,N_18506,N_18971);
and U19063 (N_19063,N_18701,N_18606);
nand U19064 (N_19064,N_18838,N_18860);
xnor U19065 (N_19065,N_18908,N_18958);
or U19066 (N_19066,N_18779,N_18780);
or U19067 (N_19067,N_18992,N_18693);
nor U19068 (N_19068,N_18768,N_18567);
xor U19069 (N_19069,N_18813,N_18922);
or U19070 (N_19070,N_18736,N_18569);
and U19071 (N_19071,N_18726,N_18553);
and U19072 (N_19072,N_18533,N_18632);
or U19073 (N_19073,N_18739,N_18662);
or U19074 (N_19074,N_18626,N_18592);
and U19075 (N_19075,N_18822,N_18646);
and U19076 (N_19076,N_18544,N_18579);
and U19077 (N_19077,N_18926,N_18973);
nor U19078 (N_19078,N_18760,N_18904);
xor U19079 (N_19079,N_18674,N_18683);
nand U19080 (N_19080,N_18689,N_18517);
and U19081 (N_19081,N_18708,N_18654);
nand U19082 (N_19082,N_18637,N_18612);
xor U19083 (N_19083,N_18872,N_18991);
and U19084 (N_19084,N_18619,N_18986);
xor U19085 (N_19085,N_18891,N_18762);
and U19086 (N_19086,N_18868,N_18532);
nor U19087 (N_19087,N_18801,N_18954);
or U19088 (N_19088,N_18631,N_18770);
nor U19089 (N_19089,N_18752,N_18564);
nor U19090 (N_19090,N_18984,N_18778);
nor U19091 (N_19091,N_18707,N_18678);
and U19092 (N_19092,N_18574,N_18695);
nand U19093 (N_19093,N_18883,N_18959);
nor U19094 (N_19094,N_18551,N_18557);
nor U19095 (N_19095,N_18727,N_18935);
and U19096 (N_19096,N_18661,N_18798);
nand U19097 (N_19097,N_18514,N_18880);
nand U19098 (N_19098,N_18607,N_18700);
and U19099 (N_19099,N_18947,N_18562);
xnor U19100 (N_19100,N_18859,N_18635);
nand U19101 (N_19101,N_18932,N_18570);
xnor U19102 (N_19102,N_18844,N_18621);
and U19103 (N_19103,N_18724,N_18797);
nor U19104 (N_19104,N_18565,N_18670);
or U19105 (N_19105,N_18783,N_18928);
nand U19106 (N_19106,N_18642,N_18924);
nor U19107 (N_19107,N_18598,N_18750);
nand U19108 (N_19108,N_18549,N_18833);
or U19109 (N_19109,N_18916,N_18671);
or U19110 (N_19110,N_18795,N_18893);
or U19111 (N_19111,N_18933,N_18806);
nand U19112 (N_19112,N_18787,N_18669);
or U19113 (N_19113,N_18681,N_18613);
nor U19114 (N_19114,N_18909,N_18913);
or U19115 (N_19115,N_18684,N_18759);
and U19116 (N_19116,N_18589,N_18983);
nand U19117 (N_19117,N_18903,N_18863);
and U19118 (N_19118,N_18876,N_18658);
nand U19119 (N_19119,N_18936,N_18865);
nor U19120 (N_19120,N_18823,N_18977);
nor U19121 (N_19121,N_18561,N_18771);
or U19122 (N_19122,N_18709,N_18805);
nor U19123 (N_19123,N_18886,N_18548);
or U19124 (N_19124,N_18576,N_18648);
xor U19125 (N_19125,N_18796,N_18829);
or U19126 (N_19126,N_18655,N_18630);
or U19127 (N_19127,N_18976,N_18899);
nand U19128 (N_19128,N_18792,N_18552);
nor U19129 (N_19129,N_18996,N_18782);
and U19130 (N_19130,N_18998,N_18625);
nor U19131 (N_19131,N_18841,N_18867);
nor U19132 (N_19132,N_18809,N_18966);
and U19133 (N_19133,N_18938,N_18748);
nand U19134 (N_19134,N_18767,N_18985);
nor U19135 (N_19135,N_18730,N_18604);
or U19136 (N_19136,N_18819,N_18757);
xor U19137 (N_19137,N_18599,N_18725);
nand U19138 (N_19138,N_18851,N_18988);
or U19139 (N_19139,N_18827,N_18907);
and U19140 (N_19140,N_18578,N_18871);
nand U19141 (N_19141,N_18970,N_18937);
nand U19142 (N_19142,N_18522,N_18581);
nand U19143 (N_19143,N_18702,N_18794);
and U19144 (N_19144,N_18667,N_18513);
nor U19145 (N_19145,N_18754,N_18616);
nor U19146 (N_19146,N_18696,N_18951);
nand U19147 (N_19147,N_18603,N_18541);
and U19148 (N_19148,N_18777,N_18888);
xor U19149 (N_19149,N_18981,N_18617);
and U19150 (N_19150,N_18814,N_18614);
or U19151 (N_19151,N_18856,N_18629);
nor U19152 (N_19152,N_18925,N_18672);
nor U19153 (N_19153,N_18870,N_18927);
nor U19154 (N_19154,N_18830,N_18944);
nand U19155 (N_19155,N_18500,N_18550);
or U19156 (N_19156,N_18566,N_18537);
xnor U19157 (N_19157,N_18609,N_18894);
nor U19158 (N_19158,N_18575,N_18885);
or U19159 (N_19159,N_18815,N_18628);
or U19160 (N_19160,N_18956,N_18807);
nand U19161 (N_19161,N_18507,N_18741);
or U19162 (N_19162,N_18595,N_18873);
and U19163 (N_19163,N_18525,N_18721);
xnor U19164 (N_19164,N_18545,N_18536);
xnor U19165 (N_19165,N_18897,N_18939);
nand U19166 (N_19166,N_18890,N_18519);
nand U19167 (N_19167,N_18699,N_18895);
nor U19168 (N_19168,N_18611,N_18593);
or U19169 (N_19169,N_18843,N_18698);
nand U19170 (N_19170,N_18948,N_18742);
xor U19171 (N_19171,N_18540,N_18824);
or U19172 (N_19172,N_18846,N_18735);
nor U19173 (N_19173,N_18518,N_18803);
xor U19174 (N_19174,N_18887,N_18784);
or U19175 (N_19175,N_18980,N_18704);
xnor U19176 (N_19176,N_18881,N_18839);
and U19177 (N_19177,N_18692,N_18582);
xnor U19178 (N_19178,N_18659,N_18821);
or U19179 (N_19179,N_18715,N_18764);
nand U19180 (N_19180,N_18543,N_18800);
xnor U19181 (N_19181,N_18845,N_18710);
and U19182 (N_19182,N_18957,N_18719);
or U19183 (N_19183,N_18663,N_18774);
nor U19184 (N_19184,N_18560,N_18531);
nand U19185 (N_19185,N_18950,N_18964);
and U19186 (N_19186,N_18753,N_18878);
xnor U19187 (N_19187,N_18694,N_18523);
xor U19188 (N_19188,N_18647,N_18905);
nand U19189 (N_19189,N_18690,N_18874);
xnor U19190 (N_19190,N_18931,N_18793);
nor U19191 (N_19191,N_18588,N_18610);
nor U19192 (N_19192,N_18989,N_18972);
and U19193 (N_19193,N_18639,N_18826);
or U19194 (N_19194,N_18656,N_18758);
nand U19195 (N_19195,N_18714,N_18901);
and U19196 (N_19196,N_18743,N_18556);
nor U19197 (N_19197,N_18978,N_18847);
nor U19198 (N_19198,N_18811,N_18919);
and U19199 (N_19199,N_18686,N_18563);
nand U19200 (N_19200,N_18502,N_18608);
nand U19201 (N_19201,N_18882,N_18825);
nand U19202 (N_19202,N_18740,N_18634);
or U19203 (N_19203,N_18769,N_18808);
nor U19204 (N_19204,N_18521,N_18812);
or U19205 (N_19205,N_18775,N_18850);
xnor U19206 (N_19206,N_18855,N_18555);
nor U19207 (N_19207,N_18965,N_18791);
nor U19208 (N_19208,N_18975,N_18831);
nor U19209 (N_19209,N_18638,N_18999);
nor U19210 (N_19210,N_18749,N_18930);
nand U19211 (N_19211,N_18974,N_18723);
or U19212 (N_19212,N_18869,N_18766);
and U19213 (N_19213,N_18718,N_18982);
nand U19214 (N_19214,N_18591,N_18993);
xnor U19215 (N_19215,N_18949,N_18605);
and U19216 (N_19216,N_18559,N_18862);
and U19217 (N_19217,N_18528,N_18990);
xor U19218 (N_19218,N_18729,N_18677);
nand U19219 (N_19219,N_18918,N_18615);
xor U19220 (N_19220,N_18968,N_18892);
nand U19221 (N_19221,N_18820,N_18772);
xnor U19222 (N_19222,N_18512,N_18685);
and U19223 (N_19223,N_18802,N_18840);
xnor U19224 (N_19224,N_18763,N_18848);
nand U19225 (N_19225,N_18568,N_18963);
nand U19226 (N_19226,N_18914,N_18712);
nand U19227 (N_19227,N_18682,N_18636);
nor U19228 (N_19228,N_18987,N_18934);
nor U19229 (N_19229,N_18955,N_18722);
xor U19230 (N_19230,N_18651,N_18504);
nand U19231 (N_19231,N_18941,N_18920);
or U19232 (N_19232,N_18697,N_18912);
and U19233 (N_19233,N_18703,N_18594);
or U19234 (N_19234,N_18618,N_18526);
nor U19235 (N_19235,N_18911,N_18751);
nand U19236 (N_19236,N_18587,N_18731);
nand U19237 (N_19237,N_18511,N_18921);
nand U19238 (N_19238,N_18624,N_18666);
nor U19239 (N_19239,N_18799,N_18547);
xnor U19240 (N_19240,N_18738,N_18508);
and U19241 (N_19241,N_18817,N_18546);
nand U19242 (N_19242,N_18879,N_18732);
nor U19243 (N_19243,N_18633,N_18884);
nor U19244 (N_19244,N_18834,N_18858);
nor U19245 (N_19245,N_18623,N_18866);
and U19246 (N_19246,N_18810,N_18917);
nand U19247 (N_19247,N_18746,N_18650);
nand U19248 (N_19248,N_18737,N_18929);
nor U19249 (N_19249,N_18584,N_18818);
nand U19250 (N_19250,N_18793,N_18779);
nand U19251 (N_19251,N_18831,N_18802);
nand U19252 (N_19252,N_18987,N_18767);
xor U19253 (N_19253,N_18723,N_18625);
and U19254 (N_19254,N_18982,N_18880);
or U19255 (N_19255,N_18639,N_18758);
and U19256 (N_19256,N_18920,N_18914);
and U19257 (N_19257,N_18528,N_18663);
or U19258 (N_19258,N_18639,N_18866);
and U19259 (N_19259,N_18675,N_18652);
and U19260 (N_19260,N_18657,N_18949);
and U19261 (N_19261,N_18801,N_18643);
nor U19262 (N_19262,N_18928,N_18632);
nor U19263 (N_19263,N_18678,N_18604);
nand U19264 (N_19264,N_18566,N_18784);
nand U19265 (N_19265,N_18848,N_18933);
nor U19266 (N_19266,N_18834,N_18559);
nand U19267 (N_19267,N_18508,N_18849);
or U19268 (N_19268,N_18775,N_18831);
or U19269 (N_19269,N_18689,N_18762);
and U19270 (N_19270,N_18537,N_18822);
and U19271 (N_19271,N_18689,N_18895);
nand U19272 (N_19272,N_18666,N_18644);
nand U19273 (N_19273,N_18590,N_18903);
or U19274 (N_19274,N_18597,N_18775);
and U19275 (N_19275,N_18924,N_18771);
and U19276 (N_19276,N_18781,N_18716);
or U19277 (N_19277,N_18816,N_18679);
and U19278 (N_19278,N_18900,N_18942);
nor U19279 (N_19279,N_18834,N_18577);
or U19280 (N_19280,N_18562,N_18823);
or U19281 (N_19281,N_18906,N_18909);
xnor U19282 (N_19282,N_18830,N_18904);
nor U19283 (N_19283,N_18534,N_18645);
nand U19284 (N_19284,N_18604,N_18676);
nand U19285 (N_19285,N_18675,N_18704);
or U19286 (N_19286,N_18991,N_18934);
or U19287 (N_19287,N_18785,N_18611);
nand U19288 (N_19288,N_18965,N_18684);
nand U19289 (N_19289,N_18800,N_18569);
nand U19290 (N_19290,N_18957,N_18949);
and U19291 (N_19291,N_18556,N_18887);
nand U19292 (N_19292,N_18978,N_18953);
xor U19293 (N_19293,N_18576,N_18909);
and U19294 (N_19294,N_18707,N_18973);
nand U19295 (N_19295,N_18565,N_18548);
nor U19296 (N_19296,N_18924,N_18811);
nand U19297 (N_19297,N_18939,N_18620);
nand U19298 (N_19298,N_18711,N_18949);
nand U19299 (N_19299,N_18789,N_18917);
and U19300 (N_19300,N_18606,N_18641);
and U19301 (N_19301,N_18533,N_18783);
or U19302 (N_19302,N_18525,N_18611);
nand U19303 (N_19303,N_18567,N_18967);
and U19304 (N_19304,N_18973,N_18505);
nand U19305 (N_19305,N_18514,N_18679);
nand U19306 (N_19306,N_18830,N_18834);
or U19307 (N_19307,N_18878,N_18880);
nand U19308 (N_19308,N_18927,N_18913);
nor U19309 (N_19309,N_18785,N_18932);
or U19310 (N_19310,N_18727,N_18902);
or U19311 (N_19311,N_18641,N_18902);
nand U19312 (N_19312,N_18753,N_18709);
or U19313 (N_19313,N_18866,N_18966);
nand U19314 (N_19314,N_18754,N_18570);
or U19315 (N_19315,N_18836,N_18901);
xnor U19316 (N_19316,N_18799,N_18843);
and U19317 (N_19317,N_18646,N_18524);
and U19318 (N_19318,N_18523,N_18517);
or U19319 (N_19319,N_18879,N_18612);
nor U19320 (N_19320,N_18947,N_18960);
or U19321 (N_19321,N_18710,N_18513);
and U19322 (N_19322,N_18553,N_18538);
and U19323 (N_19323,N_18634,N_18570);
and U19324 (N_19324,N_18604,N_18658);
nor U19325 (N_19325,N_18919,N_18693);
xnor U19326 (N_19326,N_18822,N_18512);
and U19327 (N_19327,N_18925,N_18928);
nand U19328 (N_19328,N_18668,N_18818);
xor U19329 (N_19329,N_18507,N_18814);
nand U19330 (N_19330,N_18698,N_18717);
nor U19331 (N_19331,N_18555,N_18975);
or U19332 (N_19332,N_18501,N_18697);
nand U19333 (N_19333,N_18602,N_18855);
nand U19334 (N_19334,N_18552,N_18838);
or U19335 (N_19335,N_18622,N_18871);
nand U19336 (N_19336,N_18983,N_18813);
xnor U19337 (N_19337,N_18718,N_18833);
nand U19338 (N_19338,N_18500,N_18852);
or U19339 (N_19339,N_18560,N_18895);
nor U19340 (N_19340,N_18701,N_18758);
and U19341 (N_19341,N_18804,N_18699);
nand U19342 (N_19342,N_18983,N_18649);
nand U19343 (N_19343,N_18966,N_18730);
or U19344 (N_19344,N_18804,N_18964);
nor U19345 (N_19345,N_18516,N_18593);
xor U19346 (N_19346,N_18750,N_18729);
xor U19347 (N_19347,N_18530,N_18900);
nand U19348 (N_19348,N_18528,N_18735);
and U19349 (N_19349,N_18711,N_18895);
nand U19350 (N_19350,N_18789,N_18742);
and U19351 (N_19351,N_18768,N_18873);
or U19352 (N_19352,N_18967,N_18623);
and U19353 (N_19353,N_18766,N_18963);
nand U19354 (N_19354,N_18585,N_18671);
nand U19355 (N_19355,N_18533,N_18547);
nor U19356 (N_19356,N_18893,N_18945);
or U19357 (N_19357,N_18945,N_18904);
and U19358 (N_19358,N_18803,N_18739);
or U19359 (N_19359,N_18860,N_18728);
and U19360 (N_19360,N_18687,N_18872);
or U19361 (N_19361,N_18746,N_18925);
and U19362 (N_19362,N_18643,N_18660);
or U19363 (N_19363,N_18932,N_18790);
and U19364 (N_19364,N_18654,N_18597);
nand U19365 (N_19365,N_18723,N_18508);
nand U19366 (N_19366,N_18584,N_18732);
nand U19367 (N_19367,N_18880,N_18702);
nor U19368 (N_19368,N_18853,N_18802);
and U19369 (N_19369,N_18829,N_18650);
nand U19370 (N_19370,N_18582,N_18524);
nand U19371 (N_19371,N_18756,N_18668);
xor U19372 (N_19372,N_18785,N_18602);
nand U19373 (N_19373,N_18559,N_18755);
nand U19374 (N_19374,N_18592,N_18873);
nor U19375 (N_19375,N_18964,N_18623);
nor U19376 (N_19376,N_18543,N_18577);
xor U19377 (N_19377,N_18779,N_18936);
xnor U19378 (N_19378,N_18571,N_18521);
nor U19379 (N_19379,N_18735,N_18801);
or U19380 (N_19380,N_18592,N_18931);
or U19381 (N_19381,N_18634,N_18785);
and U19382 (N_19382,N_18939,N_18596);
or U19383 (N_19383,N_18748,N_18816);
nand U19384 (N_19384,N_18847,N_18972);
nor U19385 (N_19385,N_18917,N_18706);
and U19386 (N_19386,N_18645,N_18864);
nor U19387 (N_19387,N_18537,N_18800);
or U19388 (N_19388,N_18871,N_18580);
or U19389 (N_19389,N_18536,N_18929);
or U19390 (N_19390,N_18796,N_18826);
and U19391 (N_19391,N_18661,N_18931);
nand U19392 (N_19392,N_18793,N_18726);
nand U19393 (N_19393,N_18909,N_18784);
nor U19394 (N_19394,N_18728,N_18994);
nor U19395 (N_19395,N_18988,N_18655);
nor U19396 (N_19396,N_18914,N_18874);
and U19397 (N_19397,N_18874,N_18981);
or U19398 (N_19398,N_18647,N_18897);
xnor U19399 (N_19399,N_18832,N_18637);
and U19400 (N_19400,N_18595,N_18830);
xor U19401 (N_19401,N_18920,N_18765);
and U19402 (N_19402,N_18652,N_18716);
nor U19403 (N_19403,N_18994,N_18627);
or U19404 (N_19404,N_18648,N_18881);
and U19405 (N_19405,N_18611,N_18822);
nand U19406 (N_19406,N_18901,N_18910);
and U19407 (N_19407,N_18636,N_18796);
or U19408 (N_19408,N_18748,N_18799);
and U19409 (N_19409,N_18846,N_18565);
nor U19410 (N_19410,N_18781,N_18664);
nand U19411 (N_19411,N_18670,N_18940);
nor U19412 (N_19412,N_18623,N_18676);
and U19413 (N_19413,N_18949,N_18701);
nor U19414 (N_19414,N_18513,N_18853);
or U19415 (N_19415,N_18777,N_18830);
xor U19416 (N_19416,N_18710,N_18824);
nand U19417 (N_19417,N_18915,N_18778);
or U19418 (N_19418,N_18608,N_18587);
or U19419 (N_19419,N_18934,N_18915);
nand U19420 (N_19420,N_18748,N_18523);
and U19421 (N_19421,N_18503,N_18572);
xor U19422 (N_19422,N_18674,N_18595);
or U19423 (N_19423,N_18593,N_18639);
nor U19424 (N_19424,N_18810,N_18888);
or U19425 (N_19425,N_18602,N_18880);
nand U19426 (N_19426,N_18840,N_18984);
nor U19427 (N_19427,N_18629,N_18553);
and U19428 (N_19428,N_18624,N_18650);
nand U19429 (N_19429,N_18618,N_18695);
nand U19430 (N_19430,N_18633,N_18766);
nand U19431 (N_19431,N_18544,N_18798);
nor U19432 (N_19432,N_18808,N_18556);
nand U19433 (N_19433,N_18538,N_18700);
and U19434 (N_19434,N_18665,N_18832);
or U19435 (N_19435,N_18822,N_18524);
nand U19436 (N_19436,N_18665,N_18638);
and U19437 (N_19437,N_18549,N_18877);
or U19438 (N_19438,N_18818,N_18761);
nor U19439 (N_19439,N_18936,N_18794);
nor U19440 (N_19440,N_18718,N_18687);
nand U19441 (N_19441,N_18618,N_18743);
nand U19442 (N_19442,N_18682,N_18685);
and U19443 (N_19443,N_18682,N_18677);
or U19444 (N_19444,N_18986,N_18991);
nand U19445 (N_19445,N_18623,N_18594);
or U19446 (N_19446,N_18601,N_18990);
nand U19447 (N_19447,N_18960,N_18989);
and U19448 (N_19448,N_18926,N_18641);
nand U19449 (N_19449,N_18525,N_18806);
or U19450 (N_19450,N_18717,N_18715);
and U19451 (N_19451,N_18791,N_18926);
nand U19452 (N_19452,N_18878,N_18923);
and U19453 (N_19453,N_18565,N_18920);
or U19454 (N_19454,N_18718,N_18658);
xor U19455 (N_19455,N_18966,N_18661);
or U19456 (N_19456,N_18986,N_18784);
and U19457 (N_19457,N_18974,N_18560);
and U19458 (N_19458,N_18780,N_18534);
xor U19459 (N_19459,N_18638,N_18690);
and U19460 (N_19460,N_18633,N_18692);
xnor U19461 (N_19461,N_18657,N_18923);
nor U19462 (N_19462,N_18763,N_18916);
and U19463 (N_19463,N_18964,N_18542);
nor U19464 (N_19464,N_18591,N_18770);
or U19465 (N_19465,N_18730,N_18926);
and U19466 (N_19466,N_18639,N_18892);
nor U19467 (N_19467,N_18573,N_18680);
or U19468 (N_19468,N_18571,N_18660);
nand U19469 (N_19469,N_18969,N_18646);
xnor U19470 (N_19470,N_18791,N_18960);
or U19471 (N_19471,N_18992,N_18819);
or U19472 (N_19472,N_18992,N_18967);
and U19473 (N_19473,N_18847,N_18530);
or U19474 (N_19474,N_18734,N_18630);
nand U19475 (N_19475,N_18653,N_18634);
xor U19476 (N_19476,N_18972,N_18589);
xor U19477 (N_19477,N_18772,N_18630);
nor U19478 (N_19478,N_18821,N_18695);
nor U19479 (N_19479,N_18652,N_18644);
or U19480 (N_19480,N_18603,N_18976);
or U19481 (N_19481,N_18984,N_18896);
and U19482 (N_19482,N_18570,N_18960);
nand U19483 (N_19483,N_18946,N_18982);
or U19484 (N_19484,N_18790,N_18994);
nor U19485 (N_19485,N_18701,N_18694);
nor U19486 (N_19486,N_18557,N_18795);
nand U19487 (N_19487,N_18753,N_18726);
xnor U19488 (N_19488,N_18892,N_18910);
and U19489 (N_19489,N_18962,N_18557);
nand U19490 (N_19490,N_18620,N_18717);
nor U19491 (N_19491,N_18781,N_18932);
or U19492 (N_19492,N_18771,N_18963);
xor U19493 (N_19493,N_18941,N_18560);
nand U19494 (N_19494,N_18788,N_18837);
nor U19495 (N_19495,N_18721,N_18841);
nor U19496 (N_19496,N_18779,N_18919);
nand U19497 (N_19497,N_18735,N_18794);
nand U19498 (N_19498,N_18782,N_18626);
xnor U19499 (N_19499,N_18992,N_18704);
or U19500 (N_19500,N_19452,N_19422);
nand U19501 (N_19501,N_19250,N_19117);
nand U19502 (N_19502,N_19197,N_19225);
nand U19503 (N_19503,N_19194,N_19484);
nor U19504 (N_19504,N_19086,N_19448);
nor U19505 (N_19505,N_19346,N_19491);
nor U19506 (N_19506,N_19060,N_19015);
and U19507 (N_19507,N_19005,N_19277);
nand U19508 (N_19508,N_19411,N_19386);
nor U19509 (N_19509,N_19393,N_19170);
or U19510 (N_19510,N_19327,N_19228);
nor U19511 (N_19511,N_19055,N_19283);
or U19512 (N_19512,N_19290,N_19066);
or U19513 (N_19513,N_19207,N_19017);
nor U19514 (N_19514,N_19367,N_19119);
nor U19515 (N_19515,N_19210,N_19082);
nand U19516 (N_19516,N_19404,N_19481);
xnor U19517 (N_19517,N_19300,N_19090);
nor U19518 (N_19518,N_19180,N_19103);
and U19519 (N_19519,N_19118,N_19128);
nor U19520 (N_19520,N_19043,N_19229);
and U19521 (N_19521,N_19172,N_19423);
nand U19522 (N_19522,N_19224,N_19319);
and U19523 (N_19523,N_19162,N_19465);
nor U19524 (N_19524,N_19062,N_19142);
nand U19525 (N_19525,N_19013,N_19303);
nand U19526 (N_19526,N_19173,N_19359);
nand U19527 (N_19527,N_19123,N_19392);
nand U19528 (N_19528,N_19397,N_19342);
or U19529 (N_19529,N_19489,N_19350);
nand U19530 (N_19530,N_19377,N_19253);
or U19531 (N_19531,N_19034,N_19219);
and U19532 (N_19532,N_19312,N_19395);
nand U19533 (N_19533,N_19265,N_19382);
and U19534 (N_19534,N_19094,N_19482);
nor U19535 (N_19535,N_19343,N_19193);
nor U19536 (N_19536,N_19054,N_19057);
nand U19537 (N_19537,N_19238,N_19234);
and U19538 (N_19538,N_19003,N_19487);
nand U19539 (N_19539,N_19376,N_19187);
or U19540 (N_19540,N_19361,N_19191);
and U19541 (N_19541,N_19420,N_19340);
nor U19542 (N_19542,N_19095,N_19209);
or U19543 (N_19543,N_19199,N_19112);
xor U19544 (N_19544,N_19063,N_19053);
or U19545 (N_19545,N_19202,N_19387);
nor U19546 (N_19546,N_19109,N_19488);
xor U19547 (N_19547,N_19278,N_19010);
or U19548 (N_19548,N_19485,N_19065);
nor U19549 (N_19549,N_19072,N_19284);
nor U19550 (N_19550,N_19499,N_19099);
nand U19551 (N_19551,N_19301,N_19334);
nor U19552 (N_19552,N_19433,N_19471);
and U19553 (N_19553,N_19074,N_19335);
or U19554 (N_19554,N_19154,N_19344);
nand U19555 (N_19555,N_19474,N_19051);
nand U19556 (N_19556,N_19365,N_19084);
nor U19557 (N_19557,N_19381,N_19133);
xor U19558 (N_19558,N_19476,N_19023);
nor U19559 (N_19559,N_19428,N_19092);
nand U19560 (N_19560,N_19431,N_19215);
and U19561 (N_19561,N_19497,N_19144);
and U19562 (N_19562,N_19231,N_19374);
nand U19563 (N_19563,N_19401,N_19155);
nand U19564 (N_19564,N_19473,N_19409);
or U19565 (N_19565,N_19035,N_19461);
and U19566 (N_19566,N_19220,N_19414);
nand U19567 (N_19567,N_19101,N_19379);
and U19568 (N_19568,N_19362,N_19449);
or U19569 (N_19569,N_19297,N_19490);
nand U19570 (N_19570,N_19130,N_19201);
and U19571 (N_19571,N_19432,N_19217);
and U19572 (N_19572,N_19388,N_19402);
xor U19573 (N_19573,N_19247,N_19195);
nand U19574 (N_19574,N_19111,N_19148);
or U19575 (N_19575,N_19316,N_19475);
nor U19576 (N_19576,N_19227,N_19114);
xor U19577 (N_19577,N_19178,N_19038);
and U19578 (N_19578,N_19174,N_19089);
or U19579 (N_19579,N_19218,N_19164);
and U19580 (N_19580,N_19002,N_19081);
or U19581 (N_19581,N_19368,N_19061);
nor U19582 (N_19582,N_19145,N_19143);
nor U19583 (N_19583,N_19263,N_19276);
and U19584 (N_19584,N_19059,N_19268);
and U19585 (N_19585,N_19458,N_19477);
and U19586 (N_19586,N_19168,N_19248);
nor U19587 (N_19587,N_19022,N_19236);
nand U19588 (N_19588,N_19456,N_19349);
nand U19589 (N_19589,N_19033,N_19427);
nand U19590 (N_19590,N_19241,N_19447);
or U19591 (N_19591,N_19364,N_19046);
nand U19592 (N_19592,N_19039,N_19157);
nand U19593 (N_19593,N_19026,N_19141);
and U19594 (N_19594,N_19203,N_19156);
nor U19595 (N_19595,N_19171,N_19439);
and U19596 (N_19596,N_19110,N_19345);
nand U19597 (N_19597,N_19080,N_19352);
or U19598 (N_19598,N_19434,N_19176);
nor U19599 (N_19599,N_19240,N_19208);
nand U19600 (N_19600,N_19494,N_19406);
nand U19601 (N_19601,N_19415,N_19307);
nand U19602 (N_19602,N_19037,N_19322);
or U19603 (N_19603,N_19299,N_19370);
xnor U19604 (N_19604,N_19047,N_19396);
xor U19605 (N_19605,N_19160,N_19314);
nor U19606 (N_19606,N_19271,N_19214);
xor U19607 (N_19607,N_19455,N_19151);
or U19608 (N_19608,N_19347,N_19189);
nand U19609 (N_19609,N_19252,N_19309);
nand U19610 (N_19610,N_19000,N_19177);
nand U19611 (N_19611,N_19009,N_19453);
nand U19612 (N_19612,N_19221,N_19163);
nand U19613 (N_19613,N_19104,N_19044);
nand U19614 (N_19614,N_19460,N_19242);
xor U19615 (N_19615,N_19019,N_19024);
and U19616 (N_19616,N_19320,N_19121);
and U19617 (N_19617,N_19410,N_19106);
and U19618 (N_19618,N_19318,N_19310);
and U19619 (N_19619,N_19093,N_19412);
nor U19620 (N_19620,N_19153,N_19262);
or U19621 (N_19621,N_19105,N_19042);
and U19622 (N_19622,N_19356,N_19496);
or U19623 (N_19623,N_19120,N_19472);
nor U19624 (N_19624,N_19389,N_19325);
and U19625 (N_19625,N_19182,N_19398);
nand U19626 (N_19626,N_19338,N_19069);
and U19627 (N_19627,N_19337,N_19244);
nand U19628 (N_19628,N_19048,N_19486);
or U19629 (N_19629,N_19399,N_19058);
nor U19630 (N_19630,N_19135,N_19279);
or U19631 (N_19631,N_19052,N_19152);
or U19632 (N_19632,N_19440,N_19073);
and U19633 (N_19633,N_19459,N_19137);
xor U19634 (N_19634,N_19246,N_19011);
and U19635 (N_19635,N_19351,N_19198);
nor U19636 (N_19636,N_19256,N_19190);
or U19637 (N_19637,N_19445,N_19070);
nor U19638 (N_19638,N_19281,N_19031);
nand U19639 (N_19639,N_19223,N_19298);
nand U19640 (N_19640,N_19371,N_19212);
nand U19641 (N_19641,N_19357,N_19493);
and U19642 (N_19642,N_19181,N_19492);
nor U19643 (N_19643,N_19289,N_19380);
and U19644 (N_19644,N_19341,N_19132);
and U19645 (N_19645,N_19226,N_19390);
and U19646 (N_19646,N_19408,N_19429);
xnor U19647 (N_19647,N_19235,N_19451);
or U19648 (N_19648,N_19188,N_19036);
and U19649 (N_19649,N_19165,N_19184);
nor U19650 (N_19650,N_19067,N_19331);
or U19651 (N_19651,N_19464,N_19435);
and U19652 (N_19652,N_19085,N_19071);
nor U19653 (N_19653,N_19161,N_19259);
nand U19654 (N_19654,N_19339,N_19498);
nand U19655 (N_19655,N_19267,N_19185);
nand U19656 (N_19656,N_19004,N_19463);
or U19657 (N_19657,N_19286,N_19016);
nor U19658 (N_19658,N_19025,N_19122);
nand U19659 (N_19659,N_19407,N_19315);
xor U19660 (N_19660,N_19134,N_19159);
nor U19661 (N_19661,N_19129,N_19358);
or U19662 (N_19662,N_19360,N_19293);
or U19663 (N_19663,N_19028,N_19332);
xor U19664 (N_19664,N_19313,N_19264);
and U19665 (N_19665,N_19329,N_19206);
and U19666 (N_19666,N_19027,N_19280);
and U19667 (N_19667,N_19311,N_19041);
nor U19668 (N_19668,N_19454,N_19091);
nand U19669 (N_19669,N_19323,N_19363);
nand U19670 (N_19670,N_19308,N_19317);
nand U19671 (N_19671,N_19251,N_19001);
or U19672 (N_19672,N_19083,N_19149);
or U19673 (N_19673,N_19302,N_19394);
nand U19674 (N_19674,N_19324,N_19419);
nor U19675 (N_19675,N_19478,N_19186);
or U19676 (N_19676,N_19258,N_19029);
nor U19677 (N_19677,N_19273,N_19436);
or U19678 (N_19678,N_19169,N_19125);
nand U19679 (N_19679,N_19403,N_19243);
and U19680 (N_19680,N_19049,N_19355);
nand U19681 (N_19681,N_19266,N_19348);
nor U19682 (N_19682,N_19115,N_19200);
and U19683 (N_19683,N_19075,N_19282);
and U19684 (N_19684,N_19469,N_19255);
xnor U19685 (N_19685,N_19336,N_19239);
nor U19686 (N_19686,N_19107,N_19372);
nor U19687 (N_19687,N_19450,N_19424);
nand U19688 (N_19688,N_19294,N_19088);
or U19689 (N_19689,N_19076,N_19183);
and U19690 (N_19690,N_19020,N_19369);
nor U19691 (N_19691,N_19045,N_19211);
or U19692 (N_19692,N_19012,N_19292);
and U19693 (N_19693,N_19230,N_19008);
nor U19694 (N_19694,N_19326,N_19426);
and U19695 (N_19695,N_19384,N_19295);
nor U19696 (N_19696,N_19079,N_19330);
nor U19697 (N_19697,N_19213,N_19416);
nor U19698 (N_19698,N_19442,N_19124);
and U19699 (N_19699,N_19175,N_19261);
and U19700 (N_19700,N_19275,N_19192);
nand U19701 (N_19701,N_19147,N_19158);
nand U19702 (N_19702,N_19040,N_19196);
and U19703 (N_19703,N_19288,N_19391);
and U19704 (N_19704,N_19333,N_19446);
nand U19705 (N_19705,N_19274,N_19050);
nor U19706 (N_19706,N_19366,N_19470);
nor U19707 (N_19707,N_19078,N_19405);
or U19708 (N_19708,N_19378,N_19462);
nand U19709 (N_19709,N_19006,N_19146);
nand U19710 (N_19710,N_19321,N_19131);
nor U19711 (N_19711,N_19296,N_19021);
xnor U19712 (N_19712,N_19437,N_19222);
or U19713 (N_19713,N_19413,N_19328);
and U19714 (N_19714,N_19139,N_19438);
and U19715 (N_19715,N_19400,N_19216);
or U19716 (N_19716,N_19291,N_19304);
and U19717 (N_19717,N_19441,N_19098);
nor U19718 (N_19718,N_19480,N_19064);
xnor U19719 (N_19719,N_19260,N_19254);
xnor U19720 (N_19720,N_19113,N_19425);
and U19721 (N_19721,N_19007,N_19421);
and U19722 (N_19722,N_19269,N_19237);
nand U19723 (N_19723,N_19272,N_19479);
or U19724 (N_19724,N_19375,N_19257);
and U19725 (N_19725,N_19443,N_19030);
nor U19726 (N_19726,N_19287,N_19285);
or U19727 (N_19727,N_19430,N_19127);
nand U19728 (N_19728,N_19097,N_19116);
nand U19729 (N_19729,N_19466,N_19373);
nor U19730 (N_19730,N_19150,N_19056);
nor U19731 (N_19731,N_19032,N_19245);
and U19732 (N_19732,N_19483,N_19204);
nand U19733 (N_19733,N_19249,N_19205);
or U19734 (N_19734,N_19495,N_19270);
xor U19735 (N_19735,N_19138,N_19306);
nor U19736 (N_19736,N_19468,N_19068);
xor U19737 (N_19737,N_19166,N_19100);
nor U19738 (N_19738,N_19385,N_19232);
nand U19739 (N_19739,N_19353,N_19305);
or U19740 (N_19740,N_19136,N_19417);
nor U19741 (N_19741,N_19467,N_19457);
nand U19742 (N_19742,N_19087,N_19444);
or U19743 (N_19743,N_19140,N_19018);
nand U19744 (N_19744,N_19096,N_19418);
nand U19745 (N_19745,N_19354,N_19126);
and U19746 (N_19746,N_19233,N_19167);
or U19747 (N_19747,N_19108,N_19383);
and U19748 (N_19748,N_19102,N_19179);
nand U19749 (N_19749,N_19077,N_19014);
or U19750 (N_19750,N_19290,N_19359);
and U19751 (N_19751,N_19240,N_19401);
or U19752 (N_19752,N_19120,N_19112);
and U19753 (N_19753,N_19213,N_19057);
nand U19754 (N_19754,N_19449,N_19125);
nor U19755 (N_19755,N_19241,N_19004);
xor U19756 (N_19756,N_19088,N_19077);
nor U19757 (N_19757,N_19139,N_19314);
or U19758 (N_19758,N_19051,N_19335);
nand U19759 (N_19759,N_19325,N_19318);
nand U19760 (N_19760,N_19155,N_19377);
nor U19761 (N_19761,N_19003,N_19285);
nand U19762 (N_19762,N_19265,N_19428);
xor U19763 (N_19763,N_19083,N_19324);
or U19764 (N_19764,N_19108,N_19430);
or U19765 (N_19765,N_19121,N_19482);
nor U19766 (N_19766,N_19148,N_19061);
nor U19767 (N_19767,N_19046,N_19447);
or U19768 (N_19768,N_19035,N_19244);
and U19769 (N_19769,N_19238,N_19350);
nand U19770 (N_19770,N_19134,N_19478);
nand U19771 (N_19771,N_19354,N_19268);
xor U19772 (N_19772,N_19175,N_19098);
and U19773 (N_19773,N_19346,N_19065);
nor U19774 (N_19774,N_19071,N_19347);
nand U19775 (N_19775,N_19235,N_19181);
nor U19776 (N_19776,N_19279,N_19342);
or U19777 (N_19777,N_19127,N_19182);
nand U19778 (N_19778,N_19498,N_19252);
nand U19779 (N_19779,N_19229,N_19062);
or U19780 (N_19780,N_19045,N_19373);
and U19781 (N_19781,N_19140,N_19152);
xor U19782 (N_19782,N_19009,N_19233);
nor U19783 (N_19783,N_19263,N_19494);
nand U19784 (N_19784,N_19028,N_19052);
and U19785 (N_19785,N_19447,N_19413);
nand U19786 (N_19786,N_19235,N_19494);
nor U19787 (N_19787,N_19366,N_19142);
xnor U19788 (N_19788,N_19075,N_19417);
or U19789 (N_19789,N_19005,N_19216);
or U19790 (N_19790,N_19288,N_19214);
nand U19791 (N_19791,N_19083,N_19294);
nor U19792 (N_19792,N_19366,N_19491);
nand U19793 (N_19793,N_19304,N_19444);
or U19794 (N_19794,N_19269,N_19160);
and U19795 (N_19795,N_19364,N_19297);
and U19796 (N_19796,N_19252,N_19408);
nor U19797 (N_19797,N_19296,N_19406);
nor U19798 (N_19798,N_19178,N_19377);
nand U19799 (N_19799,N_19425,N_19154);
and U19800 (N_19800,N_19318,N_19373);
xor U19801 (N_19801,N_19044,N_19258);
nand U19802 (N_19802,N_19454,N_19190);
and U19803 (N_19803,N_19088,N_19383);
nor U19804 (N_19804,N_19258,N_19071);
nor U19805 (N_19805,N_19360,N_19155);
nor U19806 (N_19806,N_19182,N_19259);
nor U19807 (N_19807,N_19041,N_19302);
nand U19808 (N_19808,N_19229,N_19169);
nor U19809 (N_19809,N_19089,N_19216);
nor U19810 (N_19810,N_19026,N_19151);
nand U19811 (N_19811,N_19339,N_19073);
xor U19812 (N_19812,N_19496,N_19067);
and U19813 (N_19813,N_19397,N_19259);
and U19814 (N_19814,N_19193,N_19483);
nand U19815 (N_19815,N_19133,N_19277);
nand U19816 (N_19816,N_19057,N_19296);
and U19817 (N_19817,N_19027,N_19278);
and U19818 (N_19818,N_19267,N_19440);
nor U19819 (N_19819,N_19406,N_19209);
nor U19820 (N_19820,N_19305,N_19230);
or U19821 (N_19821,N_19087,N_19314);
nand U19822 (N_19822,N_19367,N_19303);
and U19823 (N_19823,N_19242,N_19496);
and U19824 (N_19824,N_19466,N_19046);
nor U19825 (N_19825,N_19147,N_19133);
nand U19826 (N_19826,N_19262,N_19248);
and U19827 (N_19827,N_19384,N_19453);
nor U19828 (N_19828,N_19131,N_19163);
nor U19829 (N_19829,N_19095,N_19083);
nand U19830 (N_19830,N_19236,N_19230);
nand U19831 (N_19831,N_19435,N_19351);
nor U19832 (N_19832,N_19143,N_19204);
and U19833 (N_19833,N_19125,N_19319);
and U19834 (N_19834,N_19172,N_19119);
or U19835 (N_19835,N_19003,N_19021);
nor U19836 (N_19836,N_19342,N_19042);
nor U19837 (N_19837,N_19166,N_19281);
xnor U19838 (N_19838,N_19483,N_19421);
nor U19839 (N_19839,N_19330,N_19034);
nand U19840 (N_19840,N_19451,N_19319);
nand U19841 (N_19841,N_19231,N_19080);
nand U19842 (N_19842,N_19468,N_19465);
nand U19843 (N_19843,N_19067,N_19168);
and U19844 (N_19844,N_19454,N_19356);
or U19845 (N_19845,N_19350,N_19077);
nand U19846 (N_19846,N_19376,N_19226);
xnor U19847 (N_19847,N_19388,N_19300);
and U19848 (N_19848,N_19299,N_19077);
nor U19849 (N_19849,N_19190,N_19100);
and U19850 (N_19850,N_19107,N_19179);
and U19851 (N_19851,N_19027,N_19478);
or U19852 (N_19852,N_19092,N_19268);
nand U19853 (N_19853,N_19435,N_19295);
nor U19854 (N_19854,N_19310,N_19077);
and U19855 (N_19855,N_19033,N_19169);
or U19856 (N_19856,N_19493,N_19136);
and U19857 (N_19857,N_19078,N_19252);
nand U19858 (N_19858,N_19462,N_19013);
and U19859 (N_19859,N_19090,N_19356);
or U19860 (N_19860,N_19029,N_19031);
nand U19861 (N_19861,N_19238,N_19464);
nand U19862 (N_19862,N_19396,N_19456);
or U19863 (N_19863,N_19293,N_19421);
nor U19864 (N_19864,N_19075,N_19108);
nor U19865 (N_19865,N_19033,N_19126);
and U19866 (N_19866,N_19474,N_19285);
nor U19867 (N_19867,N_19097,N_19280);
and U19868 (N_19868,N_19245,N_19085);
nor U19869 (N_19869,N_19014,N_19092);
nand U19870 (N_19870,N_19474,N_19326);
and U19871 (N_19871,N_19473,N_19103);
xor U19872 (N_19872,N_19365,N_19190);
and U19873 (N_19873,N_19308,N_19272);
nor U19874 (N_19874,N_19194,N_19335);
nor U19875 (N_19875,N_19431,N_19017);
or U19876 (N_19876,N_19274,N_19350);
xnor U19877 (N_19877,N_19492,N_19344);
nor U19878 (N_19878,N_19149,N_19119);
nand U19879 (N_19879,N_19079,N_19296);
or U19880 (N_19880,N_19093,N_19008);
or U19881 (N_19881,N_19465,N_19029);
nor U19882 (N_19882,N_19036,N_19010);
or U19883 (N_19883,N_19193,N_19074);
nor U19884 (N_19884,N_19178,N_19085);
nor U19885 (N_19885,N_19002,N_19448);
or U19886 (N_19886,N_19156,N_19135);
nor U19887 (N_19887,N_19212,N_19341);
or U19888 (N_19888,N_19267,N_19143);
and U19889 (N_19889,N_19410,N_19335);
xor U19890 (N_19890,N_19143,N_19016);
or U19891 (N_19891,N_19034,N_19157);
nand U19892 (N_19892,N_19443,N_19201);
nand U19893 (N_19893,N_19002,N_19129);
nand U19894 (N_19894,N_19103,N_19122);
and U19895 (N_19895,N_19194,N_19097);
nand U19896 (N_19896,N_19311,N_19450);
nand U19897 (N_19897,N_19160,N_19258);
or U19898 (N_19898,N_19431,N_19188);
nand U19899 (N_19899,N_19279,N_19411);
nand U19900 (N_19900,N_19432,N_19440);
nand U19901 (N_19901,N_19457,N_19351);
xor U19902 (N_19902,N_19288,N_19079);
and U19903 (N_19903,N_19413,N_19025);
or U19904 (N_19904,N_19319,N_19169);
or U19905 (N_19905,N_19490,N_19423);
and U19906 (N_19906,N_19086,N_19349);
or U19907 (N_19907,N_19322,N_19064);
and U19908 (N_19908,N_19159,N_19215);
or U19909 (N_19909,N_19115,N_19169);
and U19910 (N_19910,N_19143,N_19223);
or U19911 (N_19911,N_19050,N_19380);
and U19912 (N_19912,N_19337,N_19051);
and U19913 (N_19913,N_19316,N_19057);
xnor U19914 (N_19914,N_19188,N_19455);
nand U19915 (N_19915,N_19482,N_19495);
and U19916 (N_19916,N_19168,N_19470);
and U19917 (N_19917,N_19066,N_19325);
nand U19918 (N_19918,N_19091,N_19002);
nand U19919 (N_19919,N_19122,N_19299);
xnor U19920 (N_19920,N_19158,N_19195);
nand U19921 (N_19921,N_19409,N_19317);
nand U19922 (N_19922,N_19357,N_19399);
nand U19923 (N_19923,N_19190,N_19370);
nand U19924 (N_19924,N_19222,N_19296);
nand U19925 (N_19925,N_19168,N_19162);
or U19926 (N_19926,N_19466,N_19375);
or U19927 (N_19927,N_19477,N_19342);
xnor U19928 (N_19928,N_19378,N_19275);
or U19929 (N_19929,N_19435,N_19349);
nor U19930 (N_19930,N_19407,N_19051);
nor U19931 (N_19931,N_19389,N_19398);
and U19932 (N_19932,N_19110,N_19358);
nor U19933 (N_19933,N_19283,N_19336);
and U19934 (N_19934,N_19280,N_19362);
and U19935 (N_19935,N_19178,N_19215);
and U19936 (N_19936,N_19399,N_19260);
nand U19937 (N_19937,N_19413,N_19271);
nor U19938 (N_19938,N_19456,N_19395);
nor U19939 (N_19939,N_19071,N_19150);
or U19940 (N_19940,N_19473,N_19480);
xnor U19941 (N_19941,N_19145,N_19044);
and U19942 (N_19942,N_19051,N_19323);
nor U19943 (N_19943,N_19456,N_19059);
and U19944 (N_19944,N_19168,N_19299);
nand U19945 (N_19945,N_19152,N_19098);
nor U19946 (N_19946,N_19384,N_19258);
nand U19947 (N_19947,N_19090,N_19152);
and U19948 (N_19948,N_19055,N_19015);
and U19949 (N_19949,N_19198,N_19126);
or U19950 (N_19950,N_19005,N_19332);
or U19951 (N_19951,N_19484,N_19128);
xor U19952 (N_19952,N_19181,N_19283);
nand U19953 (N_19953,N_19329,N_19080);
nor U19954 (N_19954,N_19482,N_19159);
and U19955 (N_19955,N_19488,N_19104);
nand U19956 (N_19956,N_19075,N_19232);
nand U19957 (N_19957,N_19489,N_19385);
nand U19958 (N_19958,N_19336,N_19267);
xnor U19959 (N_19959,N_19271,N_19029);
nand U19960 (N_19960,N_19461,N_19282);
nor U19961 (N_19961,N_19177,N_19327);
and U19962 (N_19962,N_19452,N_19328);
or U19963 (N_19963,N_19117,N_19273);
or U19964 (N_19964,N_19283,N_19377);
and U19965 (N_19965,N_19163,N_19029);
xnor U19966 (N_19966,N_19340,N_19375);
or U19967 (N_19967,N_19090,N_19331);
and U19968 (N_19968,N_19173,N_19054);
nand U19969 (N_19969,N_19246,N_19369);
xnor U19970 (N_19970,N_19294,N_19365);
nand U19971 (N_19971,N_19282,N_19038);
nand U19972 (N_19972,N_19328,N_19162);
nand U19973 (N_19973,N_19097,N_19453);
xor U19974 (N_19974,N_19490,N_19151);
nand U19975 (N_19975,N_19341,N_19251);
nor U19976 (N_19976,N_19410,N_19449);
or U19977 (N_19977,N_19122,N_19198);
nor U19978 (N_19978,N_19451,N_19453);
nand U19979 (N_19979,N_19081,N_19348);
nor U19980 (N_19980,N_19326,N_19013);
and U19981 (N_19981,N_19176,N_19466);
or U19982 (N_19982,N_19064,N_19182);
xor U19983 (N_19983,N_19338,N_19120);
and U19984 (N_19984,N_19304,N_19248);
nor U19985 (N_19985,N_19480,N_19108);
and U19986 (N_19986,N_19262,N_19238);
or U19987 (N_19987,N_19032,N_19186);
and U19988 (N_19988,N_19237,N_19206);
nand U19989 (N_19989,N_19103,N_19355);
and U19990 (N_19990,N_19045,N_19368);
xor U19991 (N_19991,N_19183,N_19084);
nand U19992 (N_19992,N_19361,N_19102);
and U19993 (N_19993,N_19191,N_19234);
nor U19994 (N_19994,N_19034,N_19254);
nor U19995 (N_19995,N_19252,N_19053);
nand U19996 (N_19996,N_19132,N_19326);
nand U19997 (N_19997,N_19386,N_19444);
nand U19998 (N_19998,N_19060,N_19107);
and U19999 (N_19999,N_19265,N_19466);
nor U20000 (N_20000,N_19833,N_19800);
or U20001 (N_20001,N_19652,N_19872);
and U20002 (N_20002,N_19842,N_19565);
nor U20003 (N_20003,N_19626,N_19932);
xor U20004 (N_20004,N_19628,N_19878);
xor U20005 (N_20005,N_19640,N_19887);
nor U20006 (N_20006,N_19982,N_19898);
nand U20007 (N_20007,N_19916,N_19763);
and U20008 (N_20008,N_19633,N_19503);
nor U20009 (N_20009,N_19750,N_19848);
nand U20010 (N_20010,N_19936,N_19637);
nor U20011 (N_20011,N_19873,N_19575);
or U20012 (N_20012,N_19632,N_19981);
nor U20013 (N_20013,N_19949,N_19972);
nor U20014 (N_20014,N_19723,N_19593);
and U20015 (N_20015,N_19894,N_19979);
nand U20016 (N_20016,N_19874,N_19529);
nand U20017 (N_20017,N_19561,N_19671);
or U20018 (N_20018,N_19557,N_19844);
nor U20019 (N_20019,N_19875,N_19850);
or U20020 (N_20020,N_19713,N_19762);
nor U20021 (N_20021,N_19854,N_19624);
xor U20022 (N_20022,N_19550,N_19920);
and U20023 (N_20023,N_19645,N_19797);
nor U20024 (N_20024,N_19798,N_19836);
xor U20025 (N_20025,N_19826,N_19794);
nor U20026 (N_20026,N_19885,N_19599);
or U20027 (N_20027,N_19735,N_19717);
nor U20028 (N_20028,N_19746,N_19992);
or U20029 (N_20029,N_19900,N_19741);
or U20030 (N_20030,N_19831,N_19657);
nor U20031 (N_20031,N_19896,N_19966);
and U20032 (N_20032,N_19748,N_19672);
nand U20033 (N_20033,N_19700,N_19879);
or U20034 (N_20034,N_19968,N_19930);
nor U20035 (N_20035,N_19917,N_19507);
and U20036 (N_20036,N_19870,N_19546);
or U20037 (N_20037,N_19967,N_19865);
nor U20038 (N_20038,N_19517,N_19654);
and U20039 (N_20039,N_19947,N_19569);
or U20040 (N_20040,N_19832,N_19564);
or U20041 (N_20041,N_19511,N_19845);
nand U20042 (N_20042,N_19918,N_19639);
nand U20043 (N_20043,N_19752,N_19704);
nor U20044 (N_20044,N_19744,N_19559);
nand U20045 (N_20045,N_19728,N_19786);
nor U20046 (N_20046,N_19883,N_19574);
or U20047 (N_20047,N_19812,N_19650);
nor U20048 (N_20048,N_19679,N_19606);
or U20049 (N_20049,N_19799,N_19998);
or U20050 (N_20050,N_19924,N_19609);
and U20051 (N_20051,N_19934,N_19975);
nor U20052 (N_20052,N_19818,N_19952);
nand U20053 (N_20053,N_19995,N_19644);
nor U20054 (N_20054,N_19675,N_19971);
xor U20055 (N_20055,N_19864,N_19931);
or U20056 (N_20056,N_19653,N_19997);
or U20057 (N_20057,N_19547,N_19510);
nand U20058 (N_20058,N_19567,N_19954);
xnor U20059 (N_20059,N_19810,N_19983);
nand U20060 (N_20060,N_19706,N_19527);
nor U20061 (N_20061,N_19835,N_19747);
nand U20062 (N_20062,N_19635,N_19803);
or U20063 (N_20063,N_19505,N_19858);
nor U20064 (N_20064,N_19587,N_19731);
nand U20065 (N_20065,N_19753,N_19525);
xor U20066 (N_20066,N_19610,N_19576);
or U20067 (N_20067,N_19780,N_19785);
nand U20068 (N_20068,N_19984,N_19862);
nor U20069 (N_20069,N_19642,N_19895);
nand U20070 (N_20070,N_19807,N_19683);
or U20071 (N_20071,N_19986,N_19751);
xnor U20072 (N_20072,N_19869,N_19777);
nor U20073 (N_20073,N_19951,N_19910);
and U20074 (N_20074,N_19915,N_19578);
nor U20075 (N_20075,N_19980,N_19860);
or U20076 (N_20076,N_19758,N_19961);
nor U20077 (N_20077,N_19891,N_19964);
xor U20078 (N_20078,N_19813,N_19715);
nor U20079 (N_20079,N_19816,N_19834);
xnor U20080 (N_20080,N_19526,N_19919);
nand U20081 (N_20081,N_19541,N_19694);
nor U20082 (N_20082,N_19782,N_19839);
nor U20083 (N_20083,N_19825,N_19781);
nand U20084 (N_20084,N_19540,N_19905);
nand U20085 (N_20085,N_19555,N_19655);
and U20086 (N_20086,N_19945,N_19608);
nand U20087 (N_20087,N_19532,N_19516);
nand U20088 (N_20088,N_19545,N_19703);
and U20089 (N_20089,N_19552,N_19745);
nand U20090 (N_20090,N_19853,N_19676);
or U20091 (N_20091,N_19535,N_19729);
nand U20092 (N_20092,N_19770,N_19793);
or U20093 (N_20093,N_19607,N_19948);
or U20094 (N_20094,N_19973,N_19674);
and U20095 (N_20095,N_19695,N_19809);
nor U20096 (N_20096,N_19987,N_19678);
xor U20097 (N_20097,N_19730,N_19859);
and U20098 (N_20098,N_19504,N_19840);
and U20099 (N_20099,N_19938,N_19590);
and U20100 (N_20100,N_19922,N_19823);
nand U20101 (N_20101,N_19696,N_19649);
nand U20102 (N_20102,N_19935,N_19778);
and U20103 (N_20103,N_19902,N_19710);
nor U20104 (N_20104,N_19620,N_19955);
or U20105 (N_20105,N_19892,N_19714);
and U20106 (N_20106,N_19913,N_19802);
nand U20107 (N_20107,N_19943,N_19662);
nand U20108 (N_20108,N_19976,N_19665);
nand U20109 (N_20109,N_19656,N_19712);
and U20110 (N_20110,N_19582,N_19542);
or U20111 (N_20111,N_19764,N_19739);
nand U20112 (N_20112,N_19629,N_19843);
xor U20113 (N_20113,N_19667,N_19549);
nand U20114 (N_20114,N_19658,N_19960);
nand U20115 (N_20115,N_19822,N_19589);
and U20116 (N_20116,N_19740,N_19824);
xnor U20117 (N_20117,N_19521,N_19876);
or U20118 (N_20118,N_19993,N_19784);
nor U20119 (N_20119,N_19937,N_19877);
nor U20120 (N_20120,N_19720,N_19779);
nand U20121 (N_20121,N_19602,N_19709);
and U20122 (N_20122,N_19622,N_19820);
xnor U20123 (N_20123,N_19737,N_19705);
nor U20124 (N_20124,N_19726,N_19698);
nor U20125 (N_20125,N_19756,N_19939);
xnor U20126 (N_20126,N_19890,N_19857);
xor U20127 (N_20127,N_19907,N_19551);
nand U20128 (N_20128,N_19994,N_19957);
and U20129 (N_20129,N_19631,N_19899);
nor U20130 (N_20130,N_19630,N_19769);
or U20131 (N_20131,N_19604,N_19861);
and U20132 (N_20132,N_19711,N_19806);
xor U20133 (N_20133,N_19623,N_19754);
or U20134 (N_20134,N_19680,N_19687);
nand U20135 (N_20135,N_19805,N_19908);
nand U20136 (N_20136,N_19722,N_19882);
nand U20137 (N_20137,N_19595,N_19940);
and U20138 (N_20138,N_19959,N_19884);
nand U20139 (N_20139,N_19988,N_19502);
nand U20140 (N_20140,N_19591,N_19742);
nor U20141 (N_20141,N_19929,N_19506);
or U20142 (N_20142,N_19594,N_19664);
nand U20143 (N_20143,N_19783,N_19603);
nor U20144 (N_20144,N_19830,N_19733);
or U20145 (N_20145,N_19787,N_19736);
and U20146 (N_20146,N_19886,N_19755);
nand U20147 (N_20147,N_19600,N_19725);
xnor U20148 (N_20148,N_19926,N_19682);
or U20149 (N_20149,N_19847,N_19871);
or U20150 (N_20150,N_19515,N_19509);
or U20151 (N_20151,N_19743,N_19612);
and U20152 (N_20152,N_19530,N_19881);
or U20153 (N_20153,N_19766,N_19566);
nor U20154 (N_20154,N_19625,N_19759);
xnor U20155 (N_20155,N_19601,N_19909);
and U20156 (N_20156,N_19911,N_19536);
nor U20157 (N_20157,N_19950,N_19841);
nor U20158 (N_20158,N_19903,N_19999);
nand U20159 (N_20159,N_19724,N_19906);
nand U20160 (N_20160,N_19627,N_19734);
nand U20161 (N_20161,N_19663,N_19942);
or U20162 (N_20162,N_19697,N_19985);
nand U20163 (N_20163,N_19651,N_19773);
nand U20164 (N_20164,N_19776,N_19838);
or U20165 (N_20165,N_19970,N_19563);
or U20166 (N_20166,N_19927,N_19866);
nor U20167 (N_20167,N_19855,N_19556);
nor U20168 (N_20168,N_19868,N_19914);
or U20169 (N_20169,N_19597,N_19904);
and U20170 (N_20170,N_19804,N_19670);
nand U20171 (N_20171,N_19923,N_19581);
and U20172 (N_20172,N_19889,N_19605);
or U20173 (N_20173,N_19958,N_19817);
nor U20174 (N_20174,N_19669,N_19821);
and U20175 (N_20175,N_19863,N_19661);
nor U20176 (N_20176,N_19962,N_19928);
nand U20177 (N_20177,N_19544,N_19616);
or U20178 (N_20178,N_19513,N_19638);
and U20179 (N_20179,N_19528,N_19636);
xnor U20180 (N_20180,N_19974,N_19522);
nand U20181 (N_20181,N_19646,N_19613);
xnor U20182 (N_20182,N_19659,N_19761);
nand U20183 (N_20183,N_19586,N_19719);
or U20184 (N_20184,N_19801,N_19888);
nor U20185 (N_20185,N_19691,N_19596);
and U20186 (N_20186,N_19965,N_19512);
or U20187 (N_20187,N_19953,N_19765);
nand U20188 (N_20188,N_19707,N_19775);
nor U20189 (N_20189,N_19757,N_19618);
nand U20190 (N_20190,N_19584,N_19690);
nor U20191 (N_20191,N_19615,N_19614);
and U20192 (N_20192,N_19538,N_19837);
or U20193 (N_20193,N_19815,N_19560);
or U20194 (N_20194,N_19641,N_19579);
nor U20195 (N_20195,N_19548,N_19956);
xor U20196 (N_20196,N_19772,N_19685);
or U20197 (N_20197,N_19553,N_19846);
or U20198 (N_20198,N_19668,N_19718);
and U20199 (N_20199,N_19933,N_19996);
nor U20200 (N_20200,N_19791,N_19851);
nor U20201 (N_20201,N_19537,N_19768);
or U20202 (N_20202,N_19583,N_19978);
xnor U20203 (N_20203,N_19539,N_19693);
and U20204 (N_20204,N_19508,N_19827);
and U20205 (N_20205,N_19666,N_19621);
and U20206 (N_20206,N_19598,N_19568);
and U20207 (N_20207,N_19963,N_19732);
nor U20208 (N_20208,N_19716,N_19558);
and U20209 (N_20209,N_19648,N_19788);
xnor U20210 (N_20210,N_19771,N_19514);
nand U20211 (N_20211,N_19727,N_19634);
and U20212 (N_20212,N_19533,N_19941);
nand U20213 (N_20213,N_19554,N_19789);
nand U20214 (N_20214,N_19760,N_19673);
and U20215 (N_20215,N_19585,N_19749);
xnor U20216 (N_20216,N_19702,N_19572);
nand U20217 (N_20217,N_19619,N_19795);
nand U20218 (N_20218,N_19944,N_19811);
nor U20219 (N_20219,N_19686,N_19808);
nor U20220 (N_20220,N_19880,N_19611);
and U20221 (N_20221,N_19699,N_19721);
or U20222 (N_20222,N_19819,N_19814);
nand U20223 (N_20223,N_19828,N_19534);
nor U20224 (N_20224,N_19774,N_19969);
and U20225 (N_20225,N_19708,N_19684);
and U20226 (N_20226,N_19588,N_19617);
and U20227 (N_20227,N_19796,N_19989);
nor U20228 (N_20228,N_19738,N_19893);
nand U20229 (N_20229,N_19571,N_19701);
nor U20230 (N_20230,N_19901,N_19991);
and U20231 (N_20231,N_19856,N_19562);
nand U20232 (N_20232,N_19523,N_19688);
nand U20233 (N_20233,N_19643,N_19501);
nand U20234 (N_20234,N_19647,N_19692);
and U20235 (N_20235,N_19580,N_19990);
or U20236 (N_20236,N_19925,N_19867);
xor U20237 (N_20237,N_19946,N_19660);
and U20238 (N_20238,N_19524,N_19573);
or U20239 (N_20239,N_19689,N_19790);
and U20240 (N_20240,N_19897,N_19829);
xor U20241 (N_20241,N_19500,N_19570);
and U20242 (N_20242,N_19912,N_19681);
nor U20243 (N_20243,N_19543,N_19921);
and U20244 (N_20244,N_19977,N_19520);
and U20245 (N_20245,N_19767,N_19519);
nor U20246 (N_20246,N_19792,N_19852);
and U20247 (N_20247,N_19849,N_19531);
nand U20248 (N_20248,N_19677,N_19577);
nand U20249 (N_20249,N_19518,N_19592);
xnor U20250 (N_20250,N_19987,N_19762);
or U20251 (N_20251,N_19733,N_19653);
nand U20252 (N_20252,N_19797,N_19848);
nand U20253 (N_20253,N_19747,N_19582);
nor U20254 (N_20254,N_19834,N_19688);
nand U20255 (N_20255,N_19568,N_19553);
and U20256 (N_20256,N_19801,N_19863);
or U20257 (N_20257,N_19651,N_19935);
or U20258 (N_20258,N_19955,N_19710);
or U20259 (N_20259,N_19742,N_19596);
nor U20260 (N_20260,N_19666,N_19795);
and U20261 (N_20261,N_19777,N_19668);
or U20262 (N_20262,N_19742,N_19799);
and U20263 (N_20263,N_19749,N_19741);
xor U20264 (N_20264,N_19931,N_19871);
nor U20265 (N_20265,N_19654,N_19513);
or U20266 (N_20266,N_19706,N_19994);
xnor U20267 (N_20267,N_19782,N_19845);
and U20268 (N_20268,N_19840,N_19887);
xnor U20269 (N_20269,N_19891,N_19967);
nand U20270 (N_20270,N_19540,N_19724);
nor U20271 (N_20271,N_19944,N_19983);
and U20272 (N_20272,N_19985,N_19991);
and U20273 (N_20273,N_19851,N_19895);
or U20274 (N_20274,N_19855,N_19896);
nand U20275 (N_20275,N_19555,N_19812);
nor U20276 (N_20276,N_19525,N_19851);
nor U20277 (N_20277,N_19585,N_19898);
or U20278 (N_20278,N_19512,N_19862);
nand U20279 (N_20279,N_19664,N_19578);
nor U20280 (N_20280,N_19736,N_19868);
nand U20281 (N_20281,N_19892,N_19736);
nor U20282 (N_20282,N_19834,N_19560);
or U20283 (N_20283,N_19800,N_19973);
and U20284 (N_20284,N_19573,N_19538);
nor U20285 (N_20285,N_19503,N_19711);
xor U20286 (N_20286,N_19621,N_19815);
nor U20287 (N_20287,N_19552,N_19548);
or U20288 (N_20288,N_19816,N_19652);
nand U20289 (N_20289,N_19735,N_19714);
nand U20290 (N_20290,N_19642,N_19915);
and U20291 (N_20291,N_19999,N_19888);
nand U20292 (N_20292,N_19569,N_19853);
and U20293 (N_20293,N_19643,N_19896);
and U20294 (N_20294,N_19653,N_19672);
xor U20295 (N_20295,N_19635,N_19688);
and U20296 (N_20296,N_19954,N_19631);
nor U20297 (N_20297,N_19619,N_19723);
nor U20298 (N_20298,N_19932,N_19678);
xnor U20299 (N_20299,N_19506,N_19886);
or U20300 (N_20300,N_19965,N_19999);
nor U20301 (N_20301,N_19577,N_19739);
xor U20302 (N_20302,N_19621,N_19910);
or U20303 (N_20303,N_19750,N_19585);
nor U20304 (N_20304,N_19681,N_19946);
nor U20305 (N_20305,N_19793,N_19577);
and U20306 (N_20306,N_19578,N_19903);
nand U20307 (N_20307,N_19710,N_19515);
or U20308 (N_20308,N_19601,N_19539);
xor U20309 (N_20309,N_19826,N_19522);
nor U20310 (N_20310,N_19848,N_19854);
xnor U20311 (N_20311,N_19582,N_19640);
nand U20312 (N_20312,N_19986,N_19891);
nor U20313 (N_20313,N_19837,N_19638);
or U20314 (N_20314,N_19590,N_19526);
nor U20315 (N_20315,N_19831,N_19762);
xor U20316 (N_20316,N_19811,N_19772);
xnor U20317 (N_20317,N_19815,N_19585);
nand U20318 (N_20318,N_19636,N_19576);
or U20319 (N_20319,N_19633,N_19995);
or U20320 (N_20320,N_19591,N_19670);
and U20321 (N_20321,N_19666,N_19956);
xor U20322 (N_20322,N_19758,N_19569);
and U20323 (N_20323,N_19537,N_19898);
nor U20324 (N_20324,N_19564,N_19961);
nand U20325 (N_20325,N_19652,N_19690);
xor U20326 (N_20326,N_19907,N_19660);
xor U20327 (N_20327,N_19910,N_19611);
nand U20328 (N_20328,N_19679,N_19716);
and U20329 (N_20329,N_19883,N_19918);
nand U20330 (N_20330,N_19943,N_19711);
xnor U20331 (N_20331,N_19634,N_19797);
and U20332 (N_20332,N_19906,N_19629);
and U20333 (N_20333,N_19891,N_19583);
and U20334 (N_20334,N_19537,N_19691);
nor U20335 (N_20335,N_19642,N_19947);
nand U20336 (N_20336,N_19938,N_19910);
and U20337 (N_20337,N_19928,N_19644);
nor U20338 (N_20338,N_19823,N_19802);
xor U20339 (N_20339,N_19610,N_19855);
xnor U20340 (N_20340,N_19886,N_19703);
or U20341 (N_20341,N_19947,N_19534);
nor U20342 (N_20342,N_19930,N_19948);
or U20343 (N_20343,N_19787,N_19968);
and U20344 (N_20344,N_19839,N_19930);
xnor U20345 (N_20345,N_19742,N_19597);
xnor U20346 (N_20346,N_19984,N_19504);
nand U20347 (N_20347,N_19745,N_19957);
or U20348 (N_20348,N_19623,N_19672);
nor U20349 (N_20349,N_19705,N_19974);
and U20350 (N_20350,N_19869,N_19624);
and U20351 (N_20351,N_19904,N_19522);
nor U20352 (N_20352,N_19856,N_19978);
or U20353 (N_20353,N_19669,N_19557);
and U20354 (N_20354,N_19922,N_19803);
or U20355 (N_20355,N_19514,N_19767);
or U20356 (N_20356,N_19830,N_19588);
nor U20357 (N_20357,N_19778,N_19627);
nor U20358 (N_20358,N_19883,N_19527);
and U20359 (N_20359,N_19822,N_19884);
and U20360 (N_20360,N_19705,N_19812);
and U20361 (N_20361,N_19649,N_19545);
and U20362 (N_20362,N_19652,N_19992);
xor U20363 (N_20363,N_19570,N_19651);
or U20364 (N_20364,N_19740,N_19879);
nand U20365 (N_20365,N_19593,N_19790);
nor U20366 (N_20366,N_19567,N_19505);
or U20367 (N_20367,N_19757,N_19729);
and U20368 (N_20368,N_19758,N_19860);
nand U20369 (N_20369,N_19741,N_19925);
nor U20370 (N_20370,N_19600,N_19976);
nand U20371 (N_20371,N_19945,N_19960);
or U20372 (N_20372,N_19751,N_19908);
or U20373 (N_20373,N_19772,N_19564);
nand U20374 (N_20374,N_19891,N_19714);
nand U20375 (N_20375,N_19972,N_19746);
nand U20376 (N_20376,N_19758,N_19506);
and U20377 (N_20377,N_19648,N_19553);
nor U20378 (N_20378,N_19681,N_19800);
and U20379 (N_20379,N_19957,N_19998);
nand U20380 (N_20380,N_19681,N_19635);
and U20381 (N_20381,N_19710,N_19605);
nand U20382 (N_20382,N_19533,N_19505);
or U20383 (N_20383,N_19574,N_19927);
and U20384 (N_20384,N_19660,N_19592);
or U20385 (N_20385,N_19774,N_19781);
nor U20386 (N_20386,N_19605,N_19846);
or U20387 (N_20387,N_19627,N_19798);
nor U20388 (N_20388,N_19738,N_19862);
nand U20389 (N_20389,N_19557,N_19956);
nor U20390 (N_20390,N_19928,N_19837);
nor U20391 (N_20391,N_19576,N_19633);
and U20392 (N_20392,N_19988,N_19630);
nor U20393 (N_20393,N_19627,N_19743);
and U20394 (N_20394,N_19670,N_19570);
and U20395 (N_20395,N_19688,N_19735);
xor U20396 (N_20396,N_19837,N_19789);
nor U20397 (N_20397,N_19582,N_19568);
and U20398 (N_20398,N_19596,N_19750);
nor U20399 (N_20399,N_19990,N_19828);
or U20400 (N_20400,N_19828,N_19930);
nand U20401 (N_20401,N_19568,N_19817);
nor U20402 (N_20402,N_19919,N_19914);
nand U20403 (N_20403,N_19569,N_19869);
nand U20404 (N_20404,N_19568,N_19722);
or U20405 (N_20405,N_19608,N_19879);
nor U20406 (N_20406,N_19842,N_19713);
and U20407 (N_20407,N_19506,N_19786);
nand U20408 (N_20408,N_19546,N_19858);
xnor U20409 (N_20409,N_19737,N_19849);
or U20410 (N_20410,N_19943,N_19736);
or U20411 (N_20411,N_19904,N_19943);
nor U20412 (N_20412,N_19704,N_19730);
or U20413 (N_20413,N_19659,N_19843);
nand U20414 (N_20414,N_19803,N_19633);
and U20415 (N_20415,N_19899,N_19689);
or U20416 (N_20416,N_19897,N_19996);
nand U20417 (N_20417,N_19771,N_19833);
nor U20418 (N_20418,N_19678,N_19772);
or U20419 (N_20419,N_19899,N_19779);
or U20420 (N_20420,N_19959,N_19955);
nand U20421 (N_20421,N_19644,N_19947);
nand U20422 (N_20422,N_19776,N_19581);
xor U20423 (N_20423,N_19582,N_19898);
nand U20424 (N_20424,N_19755,N_19941);
or U20425 (N_20425,N_19726,N_19559);
or U20426 (N_20426,N_19520,N_19727);
nor U20427 (N_20427,N_19970,N_19958);
nor U20428 (N_20428,N_19679,N_19741);
and U20429 (N_20429,N_19929,N_19773);
nand U20430 (N_20430,N_19709,N_19786);
or U20431 (N_20431,N_19802,N_19509);
nor U20432 (N_20432,N_19915,N_19950);
nand U20433 (N_20433,N_19657,N_19898);
and U20434 (N_20434,N_19909,N_19518);
nand U20435 (N_20435,N_19766,N_19896);
nor U20436 (N_20436,N_19600,N_19740);
and U20437 (N_20437,N_19986,N_19538);
xnor U20438 (N_20438,N_19583,N_19595);
xor U20439 (N_20439,N_19848,N_19818);
nand U20440 (N_20440,N_19666,N_19608);
and U20441 (N_20441,N_19806,N_19735);
or U20442 (N_20442,N_19880,N_19858);
and U20443 (N_20443,N_19958,N_19838);
and U20444 (N_20444,N_19965,N_19981);
and U20445 (N_20445,N_19640,N_19564);
nor U20446 (N_20446,N_19513,N_19689);
nor U20447 (N_20447,N_19978,N_19746);
nand U20448 (N_20448,N_19850,N_19543);
and U20449 (N_20449,N_19983,N_19698);
nand U20450 (N_20450,N_19934,N_19653);
and U20451 (N_20451,N_19631,N_19634);
xor U20452 (N_20452,N_19684,N_19846);
nand U20453 (N_20453,N_19831,N_19837);
nor U20454 (N_20454,N_19879,N_19818);
xor U20455 (N_20455,N_19893,N_19703);
and U20456 (N_20456,N_19772,N_19579);
and U20457 (N_20457,N_19768,N_19898);
nor U20458 (N_20458,N_19516,N_19830);
and U20459 (N_20459,N_19657,N_19560);
or U20460 (N_20460,N_19905,N_19799);
nor U20461 (N_20461,N_19999,N_19654);
nor U20462 (N_20462,N_19583,N_19640);
and U20463 (N_20463,N_19551,N_19582);
nand U20464 (N_20464,N_19639,N_19615);
or U20465 (N_20465,N_19686,N_19700);
nor U20466 (N_20466,N_19566,N_19599);
or U20467 (N_20467,N_19848,N_19627);
nor U20468 (N_20468,N_19527,N_19903);
or U20469 (N_20469,N_19594,N_19570);
xnor U20470 (N_20470,N_19761,N_19671);
nand U20471 (N_20471,N_19720,N_19691);
nor U20472 (N_20472,N_19806,N_19819);
nand U20473 (N_20473,N_19836,N_19735);
xor U20474 (N_20474,N_19993,N_19539);
xor U20475 (N_20475,N_19633,N_19771);
xnor U20476 (N_20476,N_19949,N_19631);
or U20477 (N_20477,N_19865,N_19782);
and U20478 (N_20478,N_19554,N_19944);
or U20479 (N_20479,N_19816,N_19782);
nor U20480 (N_20480,N_19754,N_19661);
xor U20481 (N_20481,N_19876,N_19943);
xnor U20482 (N_20482,N_19632,N_19594);
nor U20483 (N_20483,N_19729,N_19862);
nand U20484 (N_20484,N_19885,N_19668);
and U20485 (N_20485,N_19945,N_19631);
or U20486 (N_20486,N_19601,N_19662);
nor U20487 (N_20487,N_19642,N_19592);
nor U20488 (N_20488,N_19969,N_19763);
and U20489 (N_20489,N_19813,N_19944);
nor U20490 (N_20490,N_19947,N_19734);
or U20491 (N_20491,N_19739,N_19785);
or U20492 (N_20492,N_19681,N_19887);
xor U20493 (N_20493,N_19725,N_19959);
and U20494 (N_20494,N_19814,N_19601);
and U20495 (N_20495,N_19920,N_19609);
xnor U20496 (N_20496,N_19550,N_19940);
and U20497 (N_20497,N_19649,N_19668);
nor U20498 (N_20498,N_19938,N_19531);
nand U20499 (N_20499,N_19647,N_19948);
and U20500 (N_20500,N_20068,N_20004);
nand U20501 (N_20501,N_20234,N_20299);
nor U20502 (N_20502,N_20278,N_20070);
nor U20503 (N_20503,N_20294,N_20042);
or U20504 (N_20504,N_20178,N_20158);
nand U20505 (N_20505,N_20010,N_20033);
or U20506 (N_20506,N_20446,N_20157);
nand U20507 (N_20507,N_20451,N_20436);
and U20508 (N_20508,N_20409,N_20041);
xor U20509 (N_20509,N_20262,N_20413);
nor U20510 (N_20510,N_20470,N_20411);
nor U20511 (N_20511,N_20153,N_20443);
nand U20512 (N_20512,N_20031,N_20478);
and U20513 (N_20513,N_20013,N_20115);
and U20514 (N_20514,N_20452,N_20164);
nor U20515 (N_20515,N_20476,N_20160);
xnor U20516 (N_20516,N_20298,N_20114);
and U20517 (N_20517,N_20231,N_20295);
and U20518 (N_20518,N_20408,N_20496);
and U20519 (N_20519,N_20490,N_20005);
nand U20520 (N_20520,N_20019,N_20099);
nor U20521 (N_20521,N_20258,N_20350);
nand U20522 (N_20522,N_20483,N_20468);
nor U20523 (N_20523,N_20135,N_20291);
nand U20524 (N_20524,N_20080,N_20474);
or U20525 (N_20525,N_20089,N_20128);
or U20526 (N_20526,N_20312,N_20435);
xnor U20527 (N_20527,N_20123,N_20162);
nor U20528 (N_20528,N_20385,N_20392);
nand U20529 (N_20529,N_20370,N_20269);
nand U20530 (N_20530,N_20280,N_20419);
xor U20531 (N_20531,N_20210,N_20475);
nor U20532 (N_20532,N_20263,N_20473);
and U20533 (N_20533,N_20156,N_20069);
or U20534 (N_20534,N_20394,N_20060);
or U20535 (N_20535,N_20167,N_20283);
or U20536 (N_20536,N_20007,N_20108);
or U20537 (N_20537,N_20279,N_20437);
xnor U20538 (N_20538,N_20094,N_20445);
nor U20539 (N_20539,N_20239,N_20257);
xor U20540 (N_20540,N_20121,N_20377);
or U20541 (N_20541,N_20379,N_20093);
nor U20542 (N_20542,N_20259,N_20077);
and U20543 (N_20543,N_20332,N_20150);
nand U20544 (N_20544,N_20171,N_20120);
and U20545 (N_20545,N_20281,N_20139);
and U20546 (N_20546,N_20191,N_20096);
and U20547 (N_20547,N_20251,N_20368);
or U20548 (N_20548,N_20369,N_20462);
or U20549 (N_20549,N_20049,N_20039);
and U20550 (N_20550,N_20426,N_20354);
and U20551 (N_20551,N_20293,N_20497);
nor U20552 (N_20552,N_20040,N_20011);
nand U20553 (N_20553,N_20146,N_20220);
xor U20554 (N_20554,N_20087,N_20272);
nor U20555 (N_20555,N_20395,N_20481);
or U20556 (N_20556,N_20184,N_20378);
or U20557 (N_20557,N_20339,N_20166);
nor U20558 (N_20558,N_20083,N_20432);
or U20559 (N_20559,N_20499,N_20023);
or U20560 (N_20560,N_20480,N_20193);
xor U20561 (N_20561,N_20078,N_20017);
nor U20562 (N_20562,N_20075,N_20064);
nor U20563 (N_20563,N_20429,N_20202);
nor U20564 (N_20564,N_20037,N_20233);
nor U20565 (N_20565,N_20487,N_20073);
nand U20566 (N_20566,N_20381,N_20084);
nand U20567 (N_20567,N_20218,N_20058);
or U20568 (N_20568,N_20107,N_20209);
and U20569 (N_20569,N_20056,N_20386);
and U20570 (N_20570,N_20181,N_20104);
nor U20571 (N_20571,N_20255,N_20063);
and U20572 (N_20572,N_20091,N_20274);
nand U20573 (N_20573,N_20489,N_20131);
or U20574 (N_20574,N_20467,N_20149);
and U20575 (N_20575,N_20235,N_20397);
and U20576 (N_20576,N_20362,N_20217);
or U20577 (N_20577,N_20248,N_20453);
nor U20578 (N_20578,N_20138,N_20219);
or U20579 (N_20579,N_20196,N_20491);
nor U20580 (N_20580,N_20230,N_20036);
and U20581 (N_20581,N_20133,N_20169);
or U20582 (N_20582,N_20088,N_20173);
nor U20583 (N_20583,N_20389,N_20001);
nand U20584 (N_20584,N_20329,N_20079);
nor U20585 (N_20585,N_20222,N_20267);
xnor U20586 (N_20586,N_20243,N_20043);
nand U20587 (N_20587,N_20407,N_20441);
or U20588 (N_20588,N_20008,N_20309);
nand U20589 (N_20589,N_20223,N_20331);
nand U20590 (N_20590,N_20270,N_20140);
nand U20591 (N_20591,N_20029,N_20422);
or U20592 (N_20592,N_20152,N_20038);
nor U20593 (N_20593,N_20310,N_20323);
nor U20594 (N_20594,N_20137,N_20328);
nor U20595 (N_20595,N_20071,N_20449);
or U20596 (N_20596,N_20024,N_20292);
nand U20597 (N_20597,N_20410,N_20214);
nor U20598 (N_20598,N_20044,N_20003);
and U20599 (N_20599,N_20357,N_20469);
or U20600 (N_20600,N_20260,N_20117);
xor U20601 (N_20601,N_20053,N_20498);
or U20602 (N_20602,N_20431,N_20416);
nand U20603 (N_20603,N_20132,N_20225);
nor U20604 (N_20604,N_20351,N_20195);
or U20605 (N_20605,N_20006,N_20488);
or U20606 (N_20606,N_20460,N_20161);
nand U20607 (N_20607,N_20465,N_20192);
and U20608 (N_20608,N_20101,N_20126);
or U20609 (N_20609,N_20315,N_20175);
nor U20610 (N_20610,N_20335,N_20393);
or U20611 (N_20611,N_20401,N_20464);
nor U20612 (N_20612,N_20142,N_20244);
or U20613 (N_20613,N_20074,N_20485);
nor U20614 (N_20614,N_20095,N_20051);
and U20615 (N_20615,N_20026,N_20183);
nand U20616 (N_20616,N_20304,N_20418);
nor U20617 (N_20617,N_20317,N_20271);
nand U20618 (N_20618,N_20081,N_20284);
nand U20619 (N_20619,N_20247,N_20447);
nor U20620 (N_20620,N_20399,N_20287);
and U20621 (N_20621,N_20492,N_20198);
nor U20622 (N_20622,N_20384,N_20320);
nand U20623 (N_20623,N_20050,N_20415);
nor U20624 (N_20624,N_20207,N_20116);
and U20625 (N_20625,N_20296,N_20143);
and U20626 (N_20626,N_20105,N_20325);
or U20627 (N_20627,N_20085,N_20015);
nand U20628 (N_20628,N_20054,N_20176);
and U20629 (N_20629,N_20129,N_20454);
or U20630 (N_20630,N_20025,N_20308);
or U20631 (N_20631,N_20254,N_20240);
and U20632 (N_20632,N_20297,N_20012);
and U20633 (N_20633,N_20448,N_20398);
nor U20634 (N_20634,N_20282,N_20148);
xnor U20635 (N_20635,N_20159,N_20275);
nand U20636 (N_20636,N_20326,N_20302);
nor U20637 (N_20637,N_20179,N_20456);
xor U20638 (N_20638,N_20177,N_20364);
nor U20639 (N_20639,N_20215,N_20486);
or U20640 (N_20640,N_20110,N_20134);
xnor U20641 (N_20641,N_20165,N_20494);
or U20642 (N_20642,N_20034,N_20264);
xnor U20643 (N_20643,N_20414,N_20403);
or U20644 (N_20644,N_20327,N_20018);
or U20645 (N_20645,N_20402,N_20016);
nor U20646 (N_20646,N_20113,N_20337);
or U20647 (N_20647,N_20045,N_20186);
or U20648 (N_20648,N_20197,N_20185);
or U20649 (N_20649,N_20147,N_20348);
or U20650 (N_20650,N_20373,N_20000);
or U20651 (N_20651,N_20372,N_20118);
xor U20652 (N_20652,N_20366,N_20187);
nand U20653 (N_20653,N_20338,N_20450);
and U20654 (N_20654,N_20168,N_20365);
and U20655 (N_20655,N_20341,N_20122);
nand U20656 (N_20656,N_20375,N_20358);
nand U20657 (N_20657,N_20321,N_20300);
nor U20658 (N_20658,N_20330,N_20382);
or U20659 (N_20659,N_20433,N_20155);
and U20660 (N_20660,N_20180,N_20032);
and U20661 (N_20661,N_20289,N_20307);
nor U20662 (N_20662,N_20367,N_20493);
nand U20663 (N_20663,N_20380,N_20434);
or U20664 (N_20664,N_20374,N_20100);
nor U20665 (N_20665,N_20261,N_20249);
nand U20666 (N_20666,N_20438,N_20412);
xnor U20667 (N_20667,N_20022,N_20455);
nor U20668 (N_20668,N_20301,N_20216);
and U20669 (N_20669,N_20457,N_20333);
nor U20670 (N_20670,N_20232,N_20141);
nor U20671 (N_20671,N_20439,N_20027);
nor U20672 (N_20672,N_20082,N_20145);
or U20673 (N_20673,N_20065,N_20442);
nand U20674 (N_20674,N_20353,N_20406);
and U20675 (N_20675,N_20424,N_20086);
nand U20676 (N_20676,N_20371,N_20226);
nor U20677 (N_20677,N_20356,N_20035);
nand U20678 (N_20678,N_20421,N_20124);
nor U20679 (N_20679,N_20265,N_20242);
nand U20680 (N_20680,N_20224,N_20322);
nor U20681 (N_20681,N_20466,N_20163);
and U20682 (N_20682,N_20067,N_20172);
xor U20683 (N_20683,N_20072,N_20204);
or U20684 (N_20684,N_20256,N_20405);
nand U20685 (N_20685,N_20201,N_20319);
nand U20686 (N_20686,N_20046,N_20277);
nor U20687 (N_20687,N_20253,N_20286);
or U20688 (N_20688,N_20425,N_20387);
or U20689 (N_20689,N_20388,N_20237);
or U20690 (N_20690,N_20048,N_20349);
nor U20691 (N_20691,N_20288,N_20057);
or U20692 (N_20692,N_20252,N_20002);
nand U20693 (N_20693,N_20199,N_20190);
nand U20694 (N_20694,N_20154,N_20343);
or U20695 (N_20695,N_20276,N_20203);
and U20696 (N_20696,N_20189,N_20430);
nor U20697 (N_20697,N_20228,N_20363);
and U20698 (N_20698,N_20238,N_20174);
nor U20699 (N_20699,N_20344,N_20227);
or U20700 (N_20700,N_20427,N_20355);
or U20701 (N_20701,N_20484,N_20021);
nor U20702 (N_20702,N_20229,N_20090);
nor U20703 (N_20703,N_20334,N_20206);
and U20704 (N_20704,N_20318,N_20111);
or U20705 (N_20705,N_20340,N_20106);
nand U20706 (N_20706,N_20477,N_20458);
nor U20707 (N_20707,N_20324,N_20376);
nor U20708 (N_20708,N_20472,N_20311);
nand U20709 (N_20709,N_20245,N_20290);
nand U20710 (N_20710,N_20020,N_20200);
nor U20711 (N_20711,N_20052,N_20316);
nor U20712 (N_20712,N_20444,N_20306);
nor U20713 (N_20713,N_20188,N_20390);
nand U20714 (N_20714,N_20102,N_20047);
nor U20715 (N_20715,N_20213,N_20400);
nand U20716 (N_20716,N_20273,N_20030);
nand U20717 (N_20717,N_20471,N_20182);
nand U20718 (N_20718,N_20250,N_20420);
and U20719 (N_20719,N_20428,N_20144);
or U20720 (N_20720,N_20383,N_20440);
xor U20721 (N_20721,N_20266,N_20268);
and U20722 (N_20722,N_20482,N_20125);
nand U20723 (N_20723,N_20463,N_20352);
or U20724 (N_20724,N_20314,N_20055);
and U20725 (N_20725,N_20345,N_20479);
nor U20726 (N_20726,N_20130,N_20028);
nor U20727 (N_20727,N_20112,N_20396);
nand U20728 (N_20728,N_20059,N_20009);
nor U20729 (N_20729,N_20336,N_20313);
or U20730 (N_20730,N_20246,N_20423);
or U20731 (N_20731,N_20170,N_20062);
nand U20732 (N_20732,N_20359,N_20360);
nand U20733 (N_20733,N_20346,N_20212);
nor U20734 (N_20734,N_20361,N_20194);
or U20735 (N_20735,N_20461,N_20119);
and U20736 (N_20736,N_20205,N_20495);
or U20737 (N_20737,N_20061,N_20136);
or U20738 (N_20738,N_20347,N_20092);
and U20739 (N_20739,N_20066,N_20098);
nand U20740 (N_20740,N_20151,N_20391);
nor U20741 (N_20741,N_20076,N_20404);
and U20742 (N_20742,N_20417,N_20208);
nand U20743 (N_20743,N_20342,N_20014);
xor U20744 (N_20744,N_20285,N_20127);
xnor U20745 (N_20745,N_20097,N_20241);
and U20746 (N_20746,N_20305,N_20236);
and U20747 (N_20747,N_20459,N_20303);
nor U20748 (N_20748,N_20103,N_20109);
nand U20749 (N_20749,N_20211,N_20221);
nand U20750 (N_20750,N_20127,N_20434);
nand U20751 (N_20751,N_20352,N_20469);
and U20752 (N_20752,N_20161,N_20228);
nor U20753 (N_20753,N_20029,N_20129);
or U20754 (N_20754,N_20224,N_20004);
nor U20755 (N_20755,N_20063,N_20055);
nand U20756 (N_20756,N_20135,N_20029);
nor U20757 (N_20757,N_20482,N_20209);
nand U20758 (N_20758,N_20220,N_20324);
nand U20759 (N_20759,N_20444,N_20037);
nor U20760 (N_20760,N_20405,N_20080);
xnor U20761 (N_20761,N_20158,N_20133);
nand U20762 (N_20762,N_20051,N_20098);
nor U20763 (N_20763,N_20167,N_20002);
nor U20764 (N_20764,N_20034,N_20073);
or U20765 (N_20765,N_20069,N_20368);
nand U20766 (N_20766,N_20362,N_20304);
or U20767 (N_20767,N_20478,N_20264);
and U20768 (N_20768,N_20269,N_20497);
nor U20769 (N_20769,N_20180,N_20258);
nor U20770 (N_20770,N_20365,N_20101);
nand U20771 (N_20771,N_20161,N_20029);
or U20772 (N_20772,N_20207,N_20091);
nor U20773 (N_20773,N_20126,N_20473);
or U20774 (N_20774,N_20043,N_20078);
and U20775 (N_20775,N_20223,N_20275);
nor U20776 (N_20776,N_20168,N_20123);
xor U20777 (N_20777,N_20126,N_20035);
nor U20778 (N_20778,N_20119,N_20327);
nand U20779 (N_20779,N_20167,N_20470);
xnor U20780 (N_20780,N_20148,N_20061);
or U20781 (N_20781,N_20281,N_20389);
nand U20782 (N_20782,N_20113,N_20347);
xor U20783 (N_20783,N_20465,N_20492);
nand U20784 (N_20784,N_20466,N_20285);
or U20785 (N_20785,N_20173,N_20121);
or U20786 (N_20786,N_20060,N_20407);
or U20787 (N_20787,N_20181,N_20071);
nor U20788 (N_20788,N_20324,N_20031);
or U20789 (N_20789,N_20473,N_20491);
or U20790 (N_20790,N_20114,N_20285);
and U20791 (N_20791,N_20106,N_20353);
and U20792 (N_20792,N_20268,N_20447);
nand U20793 (N_20793,N_20393,N_20389);
nand U20794 (N_20794,N_20285,N_20005);
nor U20795 (N_20795,N_20020,N_20104);
or U20796 (N_20796,N_20428,N_20476);
nor U20797 (N_20797,N_20107,N_20246);
and U20798 (N_20798,N_20229,N_20375);
nand U20799 (N_20799,N_20429,N_20304);
nand U20800 (N_20800,N_20238,N_20434);
nor U20801 (N_20801,N_20472,N_20202);
and U20802 (N_20802,N_20116,N_20021);
nor U20803 (N_20803,N_20301,N_20237);
or U20804 (N_20804,N_20438,N_20115);
nor U20805 (N_20805,N_20079,N_20096);
or U20806 (N_20806,N_20382,N_20302);
xnor U20807 (N_20807,N_20111,N_20088);
or U20808 (N_20808,N_20301,N_20047);
and U20809 (N_20809,N_20362,N_20265);
nand U20810 (N_20810,N_20430,N_20381);
nand U20811 (N_20811,N_20010,N_20344);
and U20812 (N_20812,N_20248,N_20432);
or U20813 (N_20813,N_20234,N_20134);
or U20814 (N_20814,N_20350,N_20091);
nand U20815 (N_20815,N_20109,N_20040);
nand U20816 (N_20816,N_20312,N_20361);
and U20817 (N_20817,N_20136,N_20184);
nor U20818 (N_20818,N_20226,N_20197);
or U20819 (N_20819,N_20292,N_20079);
nand U20820 (N_20820,N_20293,N_20367);
and U20821 (N_20821,N_20297,N_20429);
nor U20822 (N_20822,N_20108,N_20453);
nand U20823 (N_20823,N_20250,N_20417);
and U20824 (N_20824,N_20010,N_20248);
or U20825 (N_20825,N_20134,N_20140);
nand U20826 (N_20826,N_20349,N_20375);
nand U20827 (N_20827,N_20352,N_20412);
or U20828 (N_20828,N_20361,N_20017);
or U20829 (N_20829,N_20473,N_20391);
nor U20830 (N_20830,N_20238,N_20457);
nand U20831 (N_20831,N_20219,N_20109);
or U20832 (N_20832,N_20066,N_20201);
nand U20833 (N_20833,N_20463,N_20360);
or U20834 (N_20834,N_20000,N_20346);
or U20835 (N_20835,N_20092,N_20275);
and U20836 (N_20836,N_20103,N_20041);
and U20837 (N_20837,N_20353,N_20297);
or U20838 (N_20838,N_20014,N_20144);
nand U20839 (N_20839,N_20089,N_20363);
nand U20840 (N_20840,N_20275,N_20326);
and U20841 (N_20841,N_20319,N_20197);
or U20842 (N_20842,N_20332,N_20002);
xnor U20843 (N_20843,N_20197,N_20348);
or U20844 (N_20844,N_20345,N_20415);
nor U20845 (N_20845,N_20387,N_20386);
nor U20846 (N_20846,N_20307,N_20019);
nand U20847 (N_20847,N_20348,N_20290);
nand U20848 (N_20848,N_20056,N_20127);
and U20849 (N_20849,N_20276,N_20383);
or U20850 (N_20850,N_20298,N_20382);
nand U20851 (N_20851,N_20222,N_20353);
or U20852 (N_20852,N_20376,N_20398);
xor U20853 (N_20853,N_20170,N_20266);
nor U20854 (N_20854,N_20487,N_20003);
and U20855 (N_20855,N_20200,N_20185);
nor U20856 (N_20856,N_20388,N_20299);
nor U20857 (N_20857,N_20152,N_20405);
nand U20858 (N_20858,N_20175,N_20417);
and U20859 (N_20859,N_20499,N_20411);
and U20860 (N_20860,N_20349,N_20311);
or U20861 (N_20861,N_20065,N_20179);
and U20862 (N_20862,N_20102,N_20442);
nor U20863 (N_20863,N_20349,N_20046);
or U20864 (N_20864,N_20218,N_20498);
and U20865 (N_20865,N_20118,N_20291);
nor U20866 (N_20866,N_20127,N_20218);
nand U20867 (N_20867,N_20332,N_20066);
nor U20868 (N_20868,N_20114,N_20439);
nor U20869 (N_20869,N_20265,N_20480);
nand U20870 (N_20870,N_20080,N_20277);
and U20871 (N_20871,N_20264,N_20337);
or U20872 (N_20872,N_20115,N_20126);
or U20873 (N_20873,N_20168,N_20083);
and U20874 (N_20874,N_20137,N_20397);
xnor U20875 (N_20875,N_20292,N_20035);
xnor U20876 (N_20876,N_20354,N_20263);
or U20877 (N_20877,N_20315,N_20424);
nand U20878 (N_20878,N_20051,N_20039);
and U20879 (N_20879,N_20045,N_20009);
and U20880 (N_20880,N_20102,N_20267);
and U20881 (N_20881,N_20369,N_20484);
nor U20882 (N_20882,N_20444,N_20419);
nand U20883 (N_20883,N_20101,N_20425);
and U20884 (N_20884,N_20467,N_20495);
nor U20885 (N_20885,N_20199,N_20340);
nor U20886 (N_20886,N_20018,N_20295);
nor U20887 (N_20887,N_20128,N_20391);
or U20888 (N_20888,N_20245,N_20239);
xor U20889 (N_20889,N_20440,N_20255);
or U20890 (N_20890,N_20130,N_20335);
nand U20891 (N_20891,N_20021,N_20423);
nand U20892 (N_20892,N_20499,N_20420);
nor U20893 (N_20893,N_20246,N_20093);
xor U20894 (N_20894,N_20353,N_20108);
and U20895 (N_20895,N_20283,N_20154);
nor U20896 (N_20896,N_20369,N_20360);
nor U20897 (N_20897,N_20070,N_20249);
and U20898 (N_20898,N_20299,N_20449);
or U20899 (N_20899,N_20036,N_20269);
or U20900 (N_20900,N_20308,N_20122);
nand U20901 (N_20901,N_20463,N_20387);
nor U20902 (N_20902,N_20041,N_20310);
and U20903 (N_20903,N_20213,N_20238);
or U20904 (N_20904,N_20000,N_20076);
or U20905 (N_20905,N_20288,N_20185);
nor U20906 (N_20906,N_20100,N_20044);
nand U20907 (N_20907,N_20292,N_20065);
xnor U20908 (N_20908,N_20143,N_20348);
or U20909 (N_20909,N_20228,N_20315);
nand U20910 (N_20910,N_20327,N_20081);
nand U20911 (N_20911,N_20297,N_20094);
nand U20912 (N_20912,N_20169,N_20318);
nand U20913 (N_20913,N_20187,N_20345);
nor U20914 (N_20914,N_20291,N_20275);
and U20915 (N_20915,N_20033,N_20131);
nor U20916 (N_20916,N_20118,N_20427);
nand U20917 (N_20917,N_20465,N_20098);
nor U20918 (N_20918,N_20318,N_20148);
nand U20919 (N_20919,N_20242,N_20084);
nor U20920 (N_20920,N_20140,N_20135);
nor U20921 (N_20921,N_20216,N_20374);
xnor U20922 (N_20922,N_20473,N_20274);
nand U20923 (N_20923,N_20131,N_20395);
nor U20924 (N_20924,N_20360,N_20310);
and U20925 (N_20925,N_20116,N_20432);
nor U20926 (N_20926,N_20027,N_20335);
nand U20927 (N_20927,N_20020,N_20423);
or U20928 (N_20928,N_20239,N_20128);
nand U20929 (N_20929,N_20120,N_20034);
nand U20930 (N_20930,N_20419,N_20071);
nor U20931 (N_20931,N_20152,N_20034);
nand U20932 (N_20932,N_20298,N_20008);
xor U20933 (N_20933,N_20453,N_20067);
nor U20934 (N_20934,N_20433,N_20432);
nand U20935 (N_20935,N_20442,N_20047);
xnor U20936 (N_20936,N_20451,N_20237);
nand U20937 (N_20937,N_20461,N_20185);
xnor U20938 (N_20938,N_20169,N_20099);
or U20939 (N_20939,N_20125,N_20403);
or U20940 (N_20940,N_20081,N_20306);
nand U20941 (N_20941,N_20024,N_20131);
and U20942 (N_20942,N_20458,N_20087);
or U20943 (N_20943,N_20305,N_20058);
and U20944 (N_20944,N_20102,N_20217);
or U20945 (N_20945,N_20334,N_20370);
or U20946 (N_20946,N_20444,N_20201);
or U20947 (N_20947,N_20309,N_20067);
nand U20948 (N_20948,N_20495,N_20310);
and U20949 (N_20949,N_20484,N_20497);
nand U20950 (N_20950,N_20120,N_20200);
and U20951 (N_20951,N_20310,N_20266);
nand U20952 (N_20952,N_20150,N_20090);
and U20953 (N_20953,N_20250,N_20383);
nand U20954 (N_20954,N_20032,N_20256);
nor U20955 (N_20955,N_20214,N_20173);
nor U20956 (N_20956,N_20473,N_20072);
and U20957 (N_20957,N_20370,N_20351);
or U20958 (N_20958,N_20297,N_20113);
nor U20959 (N_20959,N_20176,N_20154);
xor U20960 (N_20960,N_20078,N_20428);
nand U20961 (N_20961,N_20066,N_20047);
and U20962 (N_20962,N_20008,N_20455);
nor U20963 (N_20963,N_20317,N_20016);
nand U20964 (N_20964,N_20180,N_20300);
nor U20965 (N_20965,N_20058,N_20295);
and U20966 (N_20966,N_20185,N_20207);
nor U20967 (N_20967,N_20438,N_20177);
xnor U20968 (N_20968,N_20452,N_20091);
nor U20969 (N_20969,N_20111,N_20225);
nor U20970 (N_20970,N_20022,N_20353);
nand U20971 (N_20971,N_20319,N_20005);
or U20972 (N_20972,N_20320,N_20306);
nor U20973 (N_20973,N_20124,N_20258);
nor U20974 (N_20974,N_20051,N_20414);
or U20975 (N_20975,N_20365,N_20242);
nor U20976 (N_20976,N_20241,N_20348);
and U20977 (N_20977,N_20370,N_20080);
nor U20978 (N_20978,N_20260,N_20358);
and U20979 (N_20979,N_20038,N_20363);
or U20980 (N_20980,N_20164,N_20083);
or U20981 (N_20981,N_20381,N_20456);
or U20982 (N_20982,N_20478,N_20271);
and U20983 (N_20983,N_20225,N_20033);
or U20984 (N_20984,N_20315,N_20022);
xor U20985 (N_20985,N_20329,N_20196);
or U20986 (N_20986,N_20211,N_20169);
and U20987 (N_20987,N_20243,N_20471);
and U20988 (N_20988,N_20065,N_20268);
and U20989 (N_20989,N_20023,N_20472);
or U20990 (N_20990,N_20197,N_20201);
nand U20991 (N_20991,N_20128,N_20429);
nand U20992 (N_20992,N_20444,N_20018);
nand U20993 (N_20993,N_20087,N_20056);
nor U20994 (N_20994,N_20123,N_20350);
and U20995 (N_20995,N_20461,N_20358);
xor U20996 (N_20996,N_20167,N_20475);
and U20997 (N_20997,N_20183,N_20245);
and U20998 (N_20998,N_20144,N_20147);
nor U20999 (N_20999,N_20477,N_20487);
xor U21000 (N_21000,N_20921,N_20899);
nand U21001 (N_21001,N_20896,N_20573);
and U21002 (N_21002,N_20892,N_20676);
nand U21003 (N_21003,N_20660,N_20621);
nor U21004 (N_21004,N_20753,N_20993);
or U21005 (N_21005,N_20537,N_20666);
and U21006 (N_21006,N_20893,N_20647);
or U21007 (N_21007,N_20802,N_20694);
and U21008 (N_21008,N_20976,N_20517);
or U21009 (N_21009,N_20922,N_20655);
or U21010 (N_21010,N_20999,N_20989);
and U21011 (N_21011,N_20638,N_20630);
nor U21012 (N_21012,N_20816,N_20956);
nor U21013 (N_21013,N_20872,N_20757);
and U21014 (N_21014,N_20891,N_20553);
and U21015 (N_21015,N_20663,N_20978);
nor U21016 (N_21016,N_20811,N_20835);
and U21017 (N_21017,N_20618,N_20797);
nor U21018 (N_21018,N_20847,N_20657);
nor U21019 (N_21019,N_20939,N_20511);
nand U21020 (N_21020,N_20713,N_20724);
or U21021 (N_21021,N_20737,N_20840);
nor U21022 (N_21022,N_20503,N_20533);
nor U21023 (N_21023,N_20765,N_20581);
and U21024 (N_21024,N_20929,N_20813);
nand U21025 (N_21025,N_20826,N_20580);
nand U21026 (N_21026,N_20783,N_20843);
nand U21027 (N_21027,N_20874,N_20504);
and U21028 (N_21028,N_20550,N_20716);
nor U21029 (N_21029,N_20576,N_20602);
nor U21030 (N_21030,N_20667,N_20994);
nand U21031 (N_21031,N_20712,N_20572);
nand U21032 (N_21032,N_20617,N_20882);
and U21033 (N_21033,N_20910,N_20946);
and U21034 (N_21034,N_20933,N_20980);
nor U21035 (N_21035,N_20966,N_20991);
or U21036 (N_21036,N_20651,N_20865);
or U21037 (N_21037,N_20794,N_20658);
nand U21038 (N_21038,N_20743,N_20726);
xnor U21039 (N_21039,N_20941,N_20620);
or U21040 (N_21040,N_20687,N_20632);
nor U21041 (N_21041,N_20778,N_20914);
nand U21042 (N_21042,N_20556,N_20559);
and U21043 (N_21043,N_20858,N_20984);
nor U21044 (N_21044,N_20822,N_20803);
or U21045 (N_21045,N_20547,N_20680);
and U21046 (N_21046,N_20884,N_20661);
or U21047 (N_21047,N_20695,N_20943);
or U21048 (N_21048,N_20850,N_20997);
nor U21049 (N_21049,N_20628,N_20836);
nand U21050 (N_21050,N_20524,N_20672);
nor U21051 (N_21051,N_20586,N_20852);
nand U21052 (N_21052,N_20735,N_20972);
nor U21053 (N_21053,N_20948,N_20756);
nand U21054 (N_21054,N_20690,N_20988);
nand U21055 (N_21055,N_20679,N_20749);
and U21056 (N_21056,N_20876,N_20668);
nor U21057 (N_21057,N_20839,N_20605);
or U21058 (N_21058,N_20715,N_20886);
nand U21059 (N_21059,N_20842,N_20824);
nor U21060 (N_21060,N_20526,N_20619);
or U21061 (N_21061,N_20733,N_20534);
and U21062 (N_21062,N_20940,N_20745);
or U21063 (N_21063,N_20696,N_20755);
xnor U21064 (N_21064,N_20643,N_20830);
nor U21065 (N_21065,N_20564,N_20919);
nand U21066 (N_21066,N_20861,N_20913);
nand U21067 (N_21067,N_20810,N_20541);
and U21068 (N_21068,N_20648,N_20678);
xor U21069 (N_21069,N_20616,N_20649);
nand U21070 (N_21070,N_20624,N_20782);
and U21071 (N_21071,N_20578,N_20697);
nand U21072 (N_21072,N_20535,N_20877);
and U21073 (N_21073,N_20804,N_20799);
xor U21074 (N_21074,N_20562,N_20821);
or U21075 (N_21075,N_20645,N_20608);
nor U21076 (N_21076,N_20682,N_20543);
nand U21077 (N_21077,N_20570,N_20603);
or U21078 (N_21078,N_20700,N_20740);
and U21079 (N_21079,N_20805,N_20518);
xnor U21080 (N_21080,N_20729,N_20818);
xnor U21081 (N_21081,N_20554,N_20751);
or U21082 (N_21082,N_20525,N_20721);
and U21083 (N_21083,N_20633,N_20931);
nor U21084 (N_21084,N_20963,N_20831);
or U21085 (N_21085,N_20762,N_20641);
or U21086 (N_21086,N_20833,N_20942);
nand U21087 (N_21087,N_20841,N_20812);
nand U21088 (N_21088,N_20905,N_20703);
or U21089 (N_21089,N_20656,N_20760);
nand U21090 (N_21090,N_20631,N_20915);
nand U21091 (N_21091,N_20928,N_20873);
nor U21092 (N_21092,N_20869,N_20894);
nand U21093 (N_21093,N_20827,N_20702);
and U21094 (N_21094,N_20793,N_20857);
xor U21095 (N_21095,N_20654,N_20551);
nand U21096 (N_21096,N_20752,N_20860);
or U21097 (N_21097,N_20610,N_20856);
nand U21098 (N_21098,N_20814,N_20730);
nand U21099 (N_21099,N_20917,N_20685);
nor U21100 (N_21100,N_20834,N_20555);
nand U21101 (N_21101,N_20591,N_20722);
nand U21102 (N_21102,N_20775,N_20732);
and U21103 (N_21103,N_20817,N_20750);
nor U21104 (N_21104,N_20911,N_20614);
nor U21105 (N_21105,N_20625,N_20706);
nand U21106 (N_21106,N_20977,N_20952);
or U21107 (N_21107,N_20971,N_20998);
nor U21108 (N_21108,N_20781,N_20944);
nor U21109 (N_21109,N_20507,N_20934);
and U21110 (N_21110,N_20889,N_20653);
xor U21111 (N_21111,N_20888,N_20958);
xnor U21112 (N_21112,N_20851,N_20739);
or U21113 (N_21113,N_20809,N_20520);
nor U21114 (N_21114,N_20501,N_20642);
nand U21115 (N_21115,N_20711,N_20659);
or U21116 (N_21116,N_20574,N_20825);
and U21117 (N_21117,N_20776,N_20560);
or U21118 (N_21118,N_20594,N_20828);
nor U21119 (N_21119,N_20736,N_20837);
or U21120 (N_21120,N_20973,N_20592);
and U21121 (N_21121,N_20767,N_20612);
or U21122 (N_21122,N_20820,N_20965);
nor U21123 (N_21123,N_20954,N_20953);
nand U21124 (N_21124,N_20692,N_20968);
nor U21125 (N_21125,N_20981,N_20714);
xor U21126 (N_21126,N_20664,N_20925);
nand U21127 (N_21127,N_20741,N_20960);
and U21128 (N_21128,N_20890,N_20992);
nor U21129 (N_21129,N_20900,N_20883);
nand U21130 (N_21130,N_20975,N_20598);
nand U21131 (N_21131,N_20938,N_20774);
or U21132 (N_21132,N_20738,N_20587);
and U21133 (N_21133,N_20990,N_20565);
nand U21134 (N_21134,N_20916,N_20844);
nand U21135 (N_21135,N_20600,N_20561);
nor U21136 (N_21136,N_20719,N_20644);
nor U21137 (N_21137,N_20864,N_20540);
nor U21138 (N_21138,N_20969,N_20623);
nand U21139 (N_21139,N_20622,N_20806);
nand U21140 (N_21140,N_20516,N_20515);
and U21141 (N_21141,N_20684,N_20514);
nor U21142 (N_21142,N_20683,N_20611);
nor U21143 (N_21143,N_20780,N_20786);
nand U21144 (N_21144,N_20705,N_20800);
or U21145 (N_21145,N_20832,N_20704);
nor U21146 (N_21146,N_20639,N_20871);
xor U21147 (N_21147,N_20558,N_20571);
or U21148 (N_21148,N_20792,N_20635);
xor U21149 (N_21149,N_20523,N_20689);
nor U21150 (N_21150,N_20962,N_20878);
nor U21151 (N_21151,N_20652,N_20601);
nor U21152 (N_21152,N_20529,N_20568);
and U21153 (N_21153,N_20862,N_20609);
xnor U21154 (N_21154,N_20699,N_20983);
nor U21155 (N_21155,N_20848,N_20575);
or U21156 (N_21156,N_20508,N_20895);
xor U21157 (N_21157,N_20626,N_20771);
xor U21158 (N_21158,N_20538,N_20557);
nand U21159 (N_21159,N_20866,N_20909);
or U21160 (N_21160,N_20734,N_20770);
or U21161 (N_21161,N_20671,N_20717);
xor U21162 (N_21162,N_20691,N_20539);
or U21163 (N_21163,N_20789,N_20777);
nor U21164 (N_21164,N_20829,N_20881);
nand U21165 (N_21165,N_20807,N_20627);
nand U21166 (N_21166,N_20796,N_20903);
or U21167 (N_21167,N_20947,N_20901);
nor U21168 (N_21168,N_20823,N_20509);
nand U21169 (N_21169,N_20549,N_20763);
nand U21170 (N_21170,N_20588,N_20669);
or U21171 (N_21171,N_20701,N_20677);
nand U21172 (N_21172,N_20949,N_20566);
nand U21173 (N_21173,N_20838,N_20727);
nor U21174 (N_21174,N_20902,N_20589);
nand U21175 (N_21175,N_20926,N_20596);
or U21176 (N_21176,N_20819,N_20629);
or U21177 (N_21177,N_20674,N_20961);
nand U21178 (N_21178,N_20636,N_20924);
or U21179 (N_21179,N_20731,N_20552);
and U21180 (N_21180,N_20710,N_20747);
nor U21181 (N_21181,N_20808,N_20681);
or U21182 (N_21182,N_20646,N_20505);
or U21183 (N_21183,N_20885,N_20759);
and U21184 (N_21184,N_20613,N_20854);
and U21185 (N_21185,N_20599,N_20904);
or U21186 (N_21186,N_20791,N_20867);
and U21187 (N_21187,N_20521,N_20955);
nand U21188 (N_21188,N_20744,N_20887);
nor U21189 (N_21189,N_20606,N_20761);
nand U21190 (N_21190,N_20772,N_20615);
nand U21191 (N_21191,N_20723,N_20935);
and U21192 (N_21192,N_20546,N_20673);
and U21193 (N_21193,N_20502,N_20936);
or U21194 (N_21194,N_20579,N_20788);
nand U21195 (N_21195,N_20728,N_20879);
nand U21196 (N_21196,N_20569,N_20665);
or U21197 (N_21197,N_20506,N_20725);
or U21198 (N_21198,N_20979,N_20597);
and U21199 (N_21199,N_20920,N_20698);
nor U21200 (N_21200,N_20908,N_20531);
and U21201 (N_21201,N_20544,N_20951);
and U21202 (N_21202,N_20675,N_20906);
xor U21203 (N_21203,N_20964,N_20582);
or U21204 (N_21204,N_20742,N_20768);
and U21205 (N_21205,N_20764,N_20912);
nand U21206 (N_21206,N_20863,N_20959);
nand U21207 (N_21207,N_20593,N_20970);
nand U21208 (N_21208,N_20532,N_20512);
nor U21209 (N_21209,N_20693,N_20945);
nor U21210 (N_21210,N_20709,N_20640);
or U21211 (N_21211,N_20536,N_20996);
nor U21212 (N_21212,N_20985,N_20795);
and U21213 (N_21213,N_20986,N_20897);
or U21214 (N_21214,N_20748,N_20500);
or U21215 (N_21215,N_20987,N_20846);
and U21216 (N_21216,N_20798,N_20769);
or U21217 (N_21217,N_20662,N_20688);
nor U21218 (N_21218,N_20637,N_20585);
or U21219 (N_21219,N_20720,N_20787);
or U21220 (N_21220,N_20522,N_20583);
nand U21221 (N_21221,N_20670,N_20875);
and U21222 (N_21222,N_20974,N_20545);
and U21223 (N_21223,N_20584,N_20607);
or U21224 (N_21224,N_20950,N_20650);
and U21225 (N_21225,N_20849,N_20784);
or U21226 (N_21226,N_20758,N_20528);
or U21227 (N_21227,N_20927,N_20527);
and U21228 (N_21228,N_20779,N_20590);
and U21229 (N_21229,N_20982,N_20530);
nand U21230 (N_21230,N_20967,N_20930);
or U21231 (N_21231,N_20595,N_20932);
nand U21232 (N_21232,N_20577,N_20995);
or U21233 (N_21233,N_20542,N_20937);
nor U21234 (N_21234,N_20853,N_20790);
xor U21235 (N_21235,N_20957,N_20563);
xor U21236 (N_21236,N_20868,N_20855);
and U21237 (N_21237,N_20707,N_20548);
nand U21238 (N_21238,N_20567,N_20918);
and U21239 (N_21239,N_20870,N_20604);
nand U21240 (N_21240,N_20801,N_20510);
or U21241 (N_21241,N_20634,N_20513);
and U21242 (N_21242,N_20718,N_20766);
nor U21243 (N_21243,N_20708,N_20519);
nor U21244 (N_21244,N_20746,N_20898);
or U21245 (N_21245,N_20923,N_20773);
nand U21246 (N_21246,N_20845,N_20815);
nand U21247 (N_21247,N_20754,N_20880);
nand U21248 (N_21248,N_20859,N_20785);
nor U21249 (N_21249,N_20907,N_20686);
or U21250 (N_21250,N_20544,N_20626);
or U21251 (N_21251,N_20569,N_20912);
or U21252 (N_21252,N_20750,N_20689);
nor U21253 (N_21253,N_20869,N_20812);
or U21254 (N_21254,N_20771,N_20696);
xnor U21255 (N_21255,N_20593,N_20766);
or U21256 (N_21256,N_20855,N_20763);
nor U21257 (N_21257,N_20839,N_20867);
nor U21258 (N_21258,N_20902,N_20946);
xnor U21259 (N_21259,N_20970,N_20574);
and U21260 (N_21260,N_20820,N_20617);
and U21261 (N_21261,N_20841,N_20822);
and U21262 (N_21262,N_20710,N_20555);
or U21263 (N_21263,N_20537,N_20521);
and U21264 (N_21264,N_20891,N_20633);
nor U21265 (N_21265,N_20815,N_20705);
nand U21266 (N_21266,N_20504,N_20569);
or U21267 (N_21267,N_20529,N_20922);
nand U21268 (N_21268,N_20846,N_20954);
or U21269 (N_21269,N_20833,N_20762);
and U21270 (N_21270,N_20906,N_20640);
nand U21271 (N_21271,N_20509,N_20908);
or U21272 (N_21272,N_20966,N_20971);
nor U21273 (N_21273,N_20786,N_20708);
or U21274 (N_21274,N_20918,N_20895);
nand U21275 (N_21275,N_20975,N_20785);
and U21276 (N_21276,N_20584,N_20519);
and U21277 (N_21277,N_20829,N_20771);
or U21278 (N_21278,N_20797,N_20667);
or U21279 (N_21279,N_20565,N_20756);
or U21280 (N_21280,N_20749,N_20913);
and U21281 (N_21281,N_20721,N_20868);
nand U21282 (N_21282,N_20759,N_20862);
and U21283 (N_21283,N_20746,N_20967);
nand U21284 (N_21284,N_20938,N_20863);
nand U21285 (N_21285,N_20970,N_20797);
or U21286 (N_21286,N_20997,N_20718);
xnor U21287 (N_21287,N_20561,N_20980);
and U21288 (N_21288,N_20650,N_20686);
nor U21289 (N_21289,N_20937,N_20828);
xor U21290 (N_21290,N_20809,N_20723);
nor U21291 (N_21291,N_20626,N_20855);
or U21292 (N_21292,N_20607,N_20507);
nand U21293 (N_21293,N_20873,N_20816);
or U21294 (N_21294,N_20995,N_20890);
nor U21295 (N_21295,N_20534,N_20947);
nor U21296 (N_21296,N_20969,N_20748);
nand U21297 (N_21297,N_20641,N_20795);
or U21298 (N_21298,N_20596,N_20795);
or U21299 (N_21299,N_20669,N_20595);
or U21300 (N_21300,N_20764,N_20625);
nor U21301 (N_21301,N_20544,N_20973);
nor U21302 (N_21302,N_20728,N_20554);
nor U21303 (N_21303,N_20793,N_20790);
nor U21304 (N_21304,N_20964,N_20990);
and U21305 (N_21305,N_20592,N_20535);
nor U21306 (N_21306,N_20920,N_20606);
nor U21307 (N_21307,N_20890,N_20973);
or U21308 (N_21308,N_20976,N_20649);
nand U21309 (N_21309,N_20642,N_20808);
and U21310 (N_21310,N_20739,N_20843);
nor U21311 (N_21311,N_20598,N_20853);
and U21312 (N_21312,N_20763,N_20989);
nor U21313 (N_21313,N_20937,N_20509);
and U21314 (N_21314,N_20880,N_20833);
nand U21315 (N_21315,N_20921,N_20721);
nand U21316 (N_21316,N_20552,N_20758);
and U21317 (N_21317,N_20990,N_20908);
and U21318 (N_21318,N_20848,N_20574);
nand U21319 (N_21319,N_20858,N_20757);
nand U21320 (N_21320,N_20741,N_20860);
or U21321 (N_21321,N_20769,N_20725);
or U21322 (N_21322,N_20634,N_20859);
or U21323 (N_21323,N_20882,N_20865);
and U21324 (N_21324,N_20621,N_20737);
xor U21325 (N_21325,N_20820,N_20880);
nor U21326 (N_21326,N_20672,N_20879);
and U21327 (N_21327,N_20772,N_20764);
nor U21328 (N_21328,N_20910,N_20689);
or U21329 (N_21329,N_20772,N_20528);
nand U21330 (N_21330,N_20856,N_20731);
nor U21331 (N_21331,N_20918,N_20972);
or U21332 (N_21332,N_20672,N_20746);
and U21333 (N_21333,N_20566,N_20648);
nand U21334 (N_21334,N_20526,N_20799);
and U21335 (N_21335,N_20707,N_20986);
nand U21336 (N_21336,N_20812,N_20959);
nand U21337 (N_21337,N_20760,N_20715);
and U21338 (N_21338,N_20576,N_20744);
nor U21339 (N_21339,N_20826,N_20672);
nand U21340 (N_21340,N_20661,N_20918);
or U21341 (N_21341,N_20761,N_20982);
or U21342 (N_21342,N_20583,N_20542);
nand U21343 (N_21343,N_20800,N_20826);
xor U21344 (N_21344,N_20575,N_20769);
nor U21345 (N_21345,N_20995,N_20656);
nor U21346 (N_21346,N_20860,N_20799);
nand U21347 (N_21347,N_20783,N_20926);
nor U21348 (N_21348,N_20850,N_20979);
and U21349 (N_21349,N_20882,N_20607);
nor U21350 (N_21350,N_20575,N_20981);
or U21351 (N_21351,N_20787,N_20981);
or U21352 (N_21352,N_20973,N_20563);
and U21353 (N_21353,N_20705,N_20808);
nor U21354 (N_21354,N_20662,N_20577);
nand U21355 (N_21355,N_20591,N_20628);
xor U21356 (N_21356,N_20549,N_20702);
and U21357 (N_21357,N_20509,N_20898);
or U21358 (N_21358,N_20857,N_20708);
nor U21359 (N_21359,N_20679,N_20833);
nand U21360 (N_21360,N_20669,N_20871);
or U21361 (N_21361,N_20878,N_20676);
xor U21362 (N_21362,N_20625,N_20820);
nand U21363 (N_21363,N_20821,N_20620);
and U21364 (N_21364,N_20654,N_20594);
or U21365 (N_21365,N_20938,N_20531);
and U21366 (N_21366,N_20537,N_20556);
and U21367 (N_21367,N_20628,N_20814);
xnor U21368 (N_21368,N_20978,N_20654);
or U21369 (N_21369,N_20535,N_20583);
and U21370 (N_21370,N_20544,N_20821);
and U21371 (N_21371,N_20859,N_20579);
or U21372 (N_21372,N_20595,N_20518);
or U21373 (N_21373,N_20846,N_20861);
nand U21374 (N_21374,N_20651,N_20922);
nand U21375 (N_21375,N_20697,N_20910);
nor U21376 (N_21376,N_20667,N_20918);
xor U21377 (N_21377,N_20562,N_20972);
or U21378 (N_21378,N_20654,N_20655);
nor U21379 (N_21379,N_20838,N_20925);
nor U21380 (N_21380,N_20704,N_20975);
nand U21381 (N_21381,N_20989,N_20665);
or U21382 (N_21382,N_20810,N_20641);
nor U21383 (N_21383,N_20855,N_20740);
nor U21384 (N_21384,N_20605,N_20691);
or U21385 (N_21385,N_20990,N_20938);
nand U21386 (N_21386,N_20889,N_20865);
nor U21387 (N_21387,N_20515,N_20979);
and U21388 (N_21388,N_20730,N_20537);
nor U21389 (N_21389,N_20789,N_20687);
xor U21390 (N_21390,N_20964,N_20501);
nand U21391 (N_21391,N_20594,N_20821);
and U21392 (N_21392,N_20561,N_20929);
and U21393 (N_21393,N_20529,N_20729);
or U21394 (N_21394,N_20696,N_20808);
or U21395 (N_21395,N_20931,N_20834);
nand U21396 (N_21396,N_20844,N_20923);
nor U21397 (N_21397,N_20861,N_20838);
nand U21398 (N_21398,N_20785,N_20703);
nor U21399 (N_21399,N_20962,N_20697);
or U21400 (N_21400,N_20916,N_20541);
or U21401 (N_21401,N_20917,N_20985);
nand U21402 (N_21402,N_20709,N_20993);
nor U21403 (N_21403,N_20973,N_20998);
nand U21404 (N_21404,N_20811,N_20702);
nand U21405 (N_21405,N_20663,N_20899);
nand U21406 (N_21406,N_20881,N_20986);
xnor U21407 (N_21407,N_20714,N_20506);
nor U21408 (N_21408,N_20900,N_20773);
and U21409 (N_21409,N_20852,N_20985);
nand U21410 (N_21410,N_20803,N_20656);
nor U21411 (N_21411,N_20518,N_20513);
or U21412 (N_21412,N_20858,N_20705);
and U21413 (N_21413,N_20953,N_20522);
or U21414 (N_21414,N_20671,N_20555);
and U21415 (N_21415,N_20713,N_20526);
nand U21416 (N_21416,N_20855,N_20851);
or U21417 (N_21417,N_20685,N_20818);
and U21418 (N_21418,N_20918,N_20874);
or U21419 (N_21419,N_20898,N_20882);
and U21420 (N_21420,N_20679,N_20801);
or U21421 (N_21421,N_20684,N_20502);
and U21422 (N_21422,N_20639,N_20986);
or U21423 (N_21423,N_20668,N_20592);
nor U21424 (N_21424,N_20914,N_20538);
nor U21425 (N_21425,N_20933,N_20927);
nand U21426 (N_21426,N_20971,N_20852);
xor U21427 (N_21427,N_20885,N_20757);
or U21428 (N_21428,N_20529,N_20715);
nor U21429 (N_21429,N_20570,N_20557);
nor U21430 (N_21430,N_20656,N_20617);
nand U21431 (N_21431,N_20506,N_20710);
and U21432 (N_21432,N_20970,N_20954);
nand U21433 (N_21433,N_20850,N_20579);
or U21434 (N_21434,N_20827,N_20612);
and U21435 (N_21435,N_20622,N_20629);
nand U21436 (N_21436,N_20894,N_20792);
xor U21437 (N_21437,N_20816,N_20885);
or U21438 (N_21438,N_20767,N_20557);
xnor U21439 (N_21439,N_20506,N_20882);
and U21440 (N_21440,N_20687,N_20729);
xor U21441 (N_21441,N_20773,N_20777);
nand U21442 (N_21442,N_20909,N_20867);
and U21443 (N_21443,N_20808,N_20773);
nand U21444 (N_21444,N_20561,N_20933);
and U21445 (N_21445,N_20664,N_20780);
nand U21446 (N_21446,N_20526,N_20609);
and U21447 (N_21447,N_20755,N_20771);
nand U21448 (N_21448,N_20912,N_20793);
nor U21449 (N_21449,N_20795,N_20610);
nand U21450 (N_21450,N_20746,N_20801);
nand U21451 (N_21451,N_20832,N_20748);
nor U21452 (N_21452,N_20595,N_20624);
or U21453 (N_21453,N_20825,N_20779);
nor U21454 (N_21454,N_20532,N_20978);
or U21455 (N_21455,N_20755,N_20548);
or U21456 (N_21456,N_20918,N_20900);
nor U21457 (N_21457,N_20885,N_20964);
nor U21458 (N_21458,N_20814,N_20663);
xnor U21459 (N_21459,N_20849,N_20907);
nor U21460 (N_21460,N_20626,N_20779);
xor U21461 (N_21461,N_20791,N_20602);
and U21462 (N_21462,N_20836,N_20780);
or U21463 (N_21463,N_20770,N_20501);
nor U21464 (N_21464,N_20922,N_20864);
nor U21465 (N_21465,N_20980,N_20991);
or U21466 (N_21466,N_20665,N_20777);
nor U21467 (N_21467,N_20753,N_20909);
or U21468 (N_21468,N_20697,N_20846);
nor U21469 (N_21469,N_20922,N_20926);
and U21470 (N_21470,N_20865,N_20552);
nand U21471 (N_21471,N_20668,N_20675);
and U21472 (N_21472,N_20880,N_20705);
or U21473 (N_21473,N_20584,N_20518);
or U21474 (N_21474,N_20533,N_20944);
nand U21475 (N_21475,N_20642,N_20803);
and U21476 (N_21476,N_20661,N_20668);
nor U21477 (N_21477,N_20642,N_20591);
xnor U21478 (N_21478,N_20767,N_20803);
and U21479 (N_21479,N_20508,N_20796);
or U21480 (N_21480,N_20897,N_20674);
nand U21481 (N_21481,N_20858,N_20599);
and U21482 (N_21482,N_20904,N_20697);
nand U21483 (N_21483,N_20924,N_20716);
nor U21484 (N_21484,N_20730,N_20561);
and U21485 (N_21485,N_20872,N_20997);
nor U21486 (N_21486,N_20727,N_20667);
or U21487 (N_21487,N_20854,N_20756);
xor U21488 (N_21488,N_20751,N_20860);
and U21489 (N_21489,N_20768,N_20591);
xor U21490 (N_21490,N_20815,N_20556);
and U21491 (N_21491,N_20576,N_20618);
or U21492 (N_21492,N_20607,N_20621);
nand U21493 (N_21493,N_20874,N_20589);
or U21494 (N_21494,N_20652,N_20986);
nand U21495 (N_21495,N_20986,N_20728);
nor U21496 (N_21496,N_20566,N_20938);
and U21497 (N_21497,N_20845,N_20763);
xor U21498 (N_21498,N_20935,N_20912);
or U21499 (N_21499,N_20958,N_20803);
xnor U21500 (N_21500,N_21065,N_21276);
nand U21501 (N_21501,N_21334,N_21138);
nor U21502 (N_21502,N_21167,N_21035);
and U21503 (N_21503,N_21098,N_21487);
or U21504 (N_21504,N_21440,N_21243);
xnor U21505 (N_21505,N_21190,N_21110);
nor U21506 (N_21506,N_21090,N_21106);
or U21507 (N_21507,N_21315,N_21174);
nor U21508 (N_21508,N_21499,N_21385);
or U21509 (N_21509,N_21263,N_21235);
or U21510 (N_21510,N_21439,N_21317);
or U21511 (N_21511,N_21108,N_21053);
nand U21512 (N_21512,N_21456,N_21203);
and U21513 (N_21513,N_21102,N_21216);
and U21514 (N_21514,N_21311,N_21402);
or U21515 (N_21515,N_21394,N_21449);
nand U21516 (N_21516,N_21233,N_21044);
nand U21517 (N_21517,N_21472,N_21184);
and U21518 (N_21518,N_21146,N_21480);
or U21519 (N_21519,N_21457,N_21204);
and U21520 (N_21520,N_21361,N_21486);
xor U21521 (N_21521,N_21201,N_21023);
nor U21522 (N_21522,N_21401,N_21221);
and U21523 (N_21523,N_21058,N_21357);
nor U21524 (N_21524,N_21470,N_21337);
nand U21525 (N_21525,N_21194,N_21059);
nand U21526 (N_21526,N_21212,N_21448);
nand U21527 (N_21527,N_21326,N_21070);
and U21528 (N_21528,N_21378,N_21474);
nor U21529 (N_21529,N_21413,N_21368);
and U21530 (N_21530,N_21191,N_21262);
or U21531 (N_21531,N_21230,N_21034);
or U21532 (N_21532,N_21293,N_21393);
xnor U21533 (N_21533,N_21303,N_21002);
nor U21534 (N_21534,N_21005,N_21209);
and U21535 (N_21535,N_21389,N_21428);
and U21536 (N_21536,N_21080,N_21282);
or U21537 (N_21537,N_21195,N_21297);
or U21538 (N_21538,N_21224,N_21373);
or U21539 (N_21539,N_21313,N_21403);
or U21540 (N_21540,N_21485,N_21030);
nand U21541 (N_21541,N_21410,N_21051);
nor U21542 (N_21542,N_21495,N_21211);
and U21543 (N_21543,N_21148,N_21117);
xor U21544 (N_21544,N_21278,N_21291);
nor U21545 (N_21545,N_21241,N_21289);
nor U21546 (N_21546,N_21114,N_21140);
nand U21547 (N_21547,N_21196,N_21228);
xnor U21548 (N_21548,N_21013,N_21285);
and U21549 (N_21549,N_21476,N_21045);
and U21550 (N_21550,N_21478,N_21264);
or U21551 (N_21551,N_21255,N_21180);
and U21552 (N_21552,N_21037,N_21137);
nor U21553 (N_21553,N_21324,N_21046);
or U21554 (N_21554,N_21028,N_21238);
nor U21555 (N_21555,N_21181,N_21497);
nor U21556 (N_21556,N_21360,N_21185);
or U21557 (N_21557,N_21356,N_21436);
nand U21558 (N_21558,N_21288,N_21418);
nand U21559 (N_21559,N_21482,N_21222);
or U21560 (N_21560,N_21271,N_21392);
and U21561 (N_21561,N_21380,N_21049);
nand U21562 (N_21562,N_21060,N_21294);
nand U21563 (N_21563,N_21318,N_21284);
nand U21564 (N_21564,N_21341,N_21186);
or U21565 (N_21565,N_21157,N_21154);
nor U21566 (N_21566,N_21462,N_21340);
nand U21567 (N_21567,N_21141,N_21199);
or U21568 (N_21568,N_21375,N_21469);
xnor U21569 (N_21569,N_21111,N_21425);
and U21570 (N_21570,N_21121,N_21150);
nand U21571 (N_21571,N_21039,N_21004);
nor U21572 (N_21572,N_21197,N_21142);
nor U21573 (N_21573,N_21247,N_21447);
and U21574 (N_21574,N_21107,N_21084);
and U21575 (N_21575,N_21069,N_21163);
nand U21576 (N_21576,N_21144,N_21006);
and U21577 (N_21577,N_21493,N_21182);
and U21578 (N_21578,N_21043,N_21162);
or U21579 (N_21579,N_21423,N_21168);
and U21580 (N_21580,N_21352,N_21280);
nor U21581 (N_21581,N_21040,N_21434);
or U21582 (N_21582,N_21177,N_21089);
nor U21583 (N_21583,N_21379,N_21067);
xnor U21584 (N_21584,N_21173,N_21126);
or U21585 (N_21585,N_21187,N_21151);
nand U21586 (N_21586,N_21329,N_21075);
or U21587 (N_21587,N_21256,N_21036);
or U21588 (N_21588,N_21395,N_21412);
nand U21589 (N_21589,N_21330,N_21214);
or U21590 (N_21590,N_21419,N_21381);
xor U21591 (N_21591,N_21128,N_21279);
nor U21592 (N_21592,N_21015,N_21016);
nor U21593 (N_21593,N_21274,N_21268);
nand U21594 (N_21594,N_21261,N_21312);
or U21595 (N_21595,N_21104,N_21094);
and U21596 (N_21596,N_21057,N_21292);
or U21597 (N_21597,N_21275,N_21193);
nand U21598 (N_21598,N_21254,N_21359);
nand U21599 (N_21599,N_21076,N_21331);
nor U21600 (N_21600,N_21444,N_21236);
and U21601 (N_21601,N_21314,N_21160);
nand U21602 (N_21602,N_21112,N_21483);
nand U21603 (N_21603,N_21175,N_21012);
nand U21604 (N_21604,N_21073,N_21083);
nor U21605 (N_21605,N_21192,N_21454);
xor U21606 (N_21606,N_21158,N_21120);
or U21607 (N_21607,N_21129,N_21258);
or U21608 (N_21608,N_21382,N_21491);
nand U21609 (N_21609,N_21409,N_21091);
nand U21610 (N_21610,N_21429,N_21364);
or U21611 (N_21611,N_21398,N_21074);
or U21612 (N_21612,N_21430,N_21355);
xnor U21613 (N_21613,N_21072,N_21172);
xnor U21614 (N_21614,N_21253,N_21455);
xor U21615 (N_21615,N_21041,N_21363);
nor U21616 (N_21616,N_21450,N_21200);
nor U21617 (N_21617,N_21086,N_21215);
or U21618 (N_21618,N_21048,N_21475);
nand U21619 (N_21619,N_21229,N_21325);
nor U21620 (N_21620,N_21420,N_21219);
nor U21621 (N_21621,N_21047,N_21244);
nand U21622 (N_21622,N_21376,N_21459);
and U21623 (N_21623,N_21387,N_21479);
xor U21624 (N_21624,N_21103,N_21101);
or U21625 (N_21625,N_21490,N_21298);
nor U21626 (N_21626,N_21372,N_21404);
nand U21627 (N_21627,N_21464,N_21176);
and U21628 (N_21628,N_21097,N_21153);
nor U21629 (N_21629,N_21135,N_21115);
xnor U21630 (N_21630,N_21245,N_21122);
or U21631 (N_21631,N_21374,N_21159);
or U21632 (N_21632,N_21100,N_21477);
or U21633 (N_21633,N_21367,N_21328);
or U21634 (N_21634,N_21171,N_21198);
nand U21635 (N_21635,N_21446,N_21408);
or U21636 (N_21636,N_21061,N_21003);
nand U21637 (N_21637,N_21025,N_21345);
and U21638 (N_21638,N_21118,N_21347);
nand U21639 (N_21639,N_21309,N_21386);
nand U21640 (N_21640,N_21131,N_21068);
or U21641 (N_21641,N_21435,N_21250);
or U21642 (N_21642,N_21064,N_21437);
and U21643 (N_21643,N_21488,N_21252);
nor U21644 (N_21644,N_21000,N_21179);
nand U21645 (N_21645,N_21096,N_21400);
nand U21646 (N_21646,N_21283,N_21371);
nor U21647 (N_21647,N_21319,N_21422);
or U21648 (N_21648,N_21099,N_21332);
nor U21649 (N_21649,N_21390,N_21348);
nor U21650 (N_21650,N_21431,N_21169);
and U21651 (N_21651,N_21414,N_21277);
and U21652 (N_21652,N_21145,N_21052);
and U21653 (N_21653,N_21339,N_21259);
nand U21654 (N_21654,N_21316,N_21498);
nor U21655 (N_21655,N_21438,N_21147);
xor U21656 (N_21656,N_21270,N_21208);
and U21657 (N_21657,N_21333,N_21354);
nand U21658 (N_21658,N_21411,N_21489);
nand U21659 (N_21659,N_21161,N_21042);
nand U21660 (N_21660,N_21134,N_21239);
xnor U21661 (N_21661,N_21024,N_21467);
nor U21662 (N_21662,N_21082,N_21050);
nand U21663 (N_21663,N_21353,N_21077);
and U21664 (N_21664,N_21299,N_21442);
and U21665 (N_21665,N_21267,N_21205);
and U21666 (N_21666,N_21383,N_21266);
nor U21667 (N_21667,N_21071,N_21441);
or U21668 (N_21668,N_21471,N_21327);
xnor U21669 (N_21669,N_21170,N_21018);
or U21670 (N_21670,N_21246,N_21029);
nor U21671 (N_21671,N_21007,N_21105);
nand U21672 (N_21672,N_21249,N_21133);
or U21673 (N_21673,N_21451,N_21010);
xor U21674 (N_21674,N_21113,N_21321);
nand U21675 (N_21675,N_21066,N_21062);
or U21676 (N_21676,N_21468,N_21308);
and U21677 (N_21677,N_21139,N_21310);
and U21678 (N_21678,N_21484,N_21031);
and U21679 (N_21679,N_21188,N_21033);
or U21680 (N_21680,N_21492,N_21335);
and U21681 (N_21681,N_21286,N_21156);
or U21682 (N_21682,N_21362,N_21370);
or U21683 (N_21683,N_21295,N_21251);
or U21684 (N_21684,N_21009,N_21116);
and U21685 (N_21685,N_21225,N_21054);
nor U21686 (N_21686,N_21302,N_21384);
nor U21687 (N_21687,N_21088,N_21143);
and U21688 (N_21688,N_21453,N_21452);
and U21689 (N_21689,N_21183,N_21443);
or U21690 (N_21690,N_21269,N_21323);
nand U21691 (N_21691,N_21304,N_21217);
or U21692 (N_21692,N_21322,N_21405);
and U21693 (N_21693,N_21237,N_21032);
nand U21694 (N_21694,N_21306,N_21260);
nand U21695 (N_21695,N_21349,N_21272);
nor U21696 (N_21696,N_21206,N_21119);
nor U21697 (N_21697,N_21473,N_21377);
and U21698 (N_21698,N_21290,N_21223);
nor U21699 (N_21699,N_21008,N_21426);
or U21700 (N_21700,N_21095,N_21424);
nor U21701 (N_21701,N_21127,N_21458);
nand U21702 (N_21702,N_21369,N_21432);
nor U21703 (N_21703,N_21496,N_21078);
or U21704 (N_21704,N_21011,N_21242);
nand U21705 (N_21705,N_21001,N_21085);
nor U21706 (N_21706,N_21240,N_21027);
or U21707 (N_21707,N_21152,N_21218);
and U21708 (N_21708,N_21465,N_21130);
nor U21709 (N_21709,N_21336,N_21273);
or U21710 (N_21710,N_21366,N_21165);
nand U21711 (N_21711,N_21343,N_21155);
and U21712 (N_21712,N_21494,N_21307);
or U21713 (N_21713,N_21296,N_21227);
and U21714 (N_21714,N_21124,N_21358);
and U21715 (N_21715,N_21210,N_21460);
nand U21716 (N_21716,N_21092,N_21164);
or U21717 (N_21717,N_21399,N_21417);
nand U21718 (N_21718,N_21301,N_21081);
and U21719 (N_21719,N_21342,N_21463);
and U21720 (N_21720,N_21020,N_21351);
nor U21721 (N_21721,N_21406,N_21178);
or U21722 (N_21722,N_21466,N_21407);
xnor U21723 (N_21723,N_21166,N_21213);
nor U21724 (N_21724,N_21287,N_21391);
nand U21725 (N_21725,N_21014,N_21132);
and U21726 (N_21726,N_21189,N_21445);
nor U21727 (N_21727,N_21338,N_21346);
and U21728 (N_21728,N_21265,N_21149);
xor U21729 (N_21729,N_21427,N_21220);
and U21730 (N_21730,N_21021,N_21022);
nand U21731 (N_21731,N_21125,N_21231);
xor U21732 (N_21732,N_21397,N_21087);
or U21733 (N_21733,N_21461,N_21055);
xnor U21734 (N_21734,N_21232,N_21017);
nand U21735 (N_21735,N_21234,N_21056);
and U21736 (N_21736,N_21207,N_21109);
nand U21737 (N_21737,N_21257,N_21063);
or U21738 (N_21738,N_21093,N_21320);
xnor U21739 (N_21739,N_21433,N_21481);
nand U21740 (N_21740,N_21344,N_21305);
and U21741 (N_21741,N_21350,N_21226);
or U21742 (N_21742,N_21136,N_21038);
or U21743 (N_21743,N_21396,N_21416);
nor U21744 (N_21744,N_21415,N_21388);
and U21745 (N_21745,N_21281,N_21248);
nand U21746 (N_21746,N_21421,N_21300);
nor U21747 (N_21747,N_21026,N_21202);
nand U21748 (N_21748,N_21123,N_21365);
or U21749 (N_21749,N_21019,N_21079);
or U21750 (N_21750,N_21280,N_21125);
nand U21751 (N_21751,N_21138,N_21490);
or U21752 (N_21752,N_21098,N_21140);
nand U21753 (N_21753,N_21068,N_21117);
and U21754 (N_21754,N_21226,N_21242);
nand U21755 (N_21755,N_21363,N_21303);
or U21756 (N_21756,N_21000,N_21164);
xnor U21757 (N_21757,N_21260,N_21213);
and U21758 (N_21758,N_21008,N_21018);
nor U21759 (N_21759,N_21074,N_21176);
or U21760 (N_21760,N_21156,N_21219);
nor U21761 (N_21761,N_21262,N_21044);
and U21762 (N_21762,N_21327,N_21464);
nand U21763 (N_21763,N_21130,N_21297);
or U21764 (N_21764,N_21298,N_21115);
nand U21765 (N_21765,N_21315,N_21215);
nor U21766 (N_21766,N_21207,N_21400);
nand U21767 (N_21767,N_21481,N_21220);
nand U21768 (N_21768,N_21186,N_21352);
and U21769 (N_21769,N_21265,N_21014);
nand U21770 (N_21770,N_21170,N_21457);
nand U21771 (N_21771,N_21496,N_21256);
nor U21772 (N_21772,N_21082,N_21367);
nand U21773 (N_21773,N_21131,N_21290);
and U21774 (N_21774,N_21380,N_21406);
nor U21775 (N_21775,N_21021,N_21307);
nor U21776 (N_21776,N_21335,N_21188);
or U21777 (N_21777,N_21416,N_21368);
nor U21778 (N_21778,N_21460,N_21003);
xor U21779 (N_21779,N_21012,N_21379);
nor U21780 (N_21780,N_21033,N_21271);
or U21781 (N_21781,N_21475,N_21102);
and U21782 (N_21782,N_21002,N_21070);
and U21783 (N_21783,N_21425,N_21148);
nor U21784 (N_21784,N_21369,N_21181);
or U21785 (N_21785,N_21040,N_21394);
or U21786 (N_21786,N_21243,N_21482);
nand U21787 (N_21787,N_21111,N_21223);
nor U21788 (N_21788,N_21015,N_21498);
or U21789 (N_21789,N_21493,N_21041);
or U21790 (N_21790,N_21486,N_21027);
or U21791 (N_21791,N_21456,N_21144);
and U21792 (N_21792,N_21055,N_21323);
or U21793 (N_21793,N_21480,N_21286);
nor U21794 (N_21794,N_21352,N_21096);
nor U21795 (N_21795,N_21221,N_21277);
or U21796 (N_21796,N_21086,N_21484);
nand U21797 (N_21797,N_21035,N_21334);
xor U21798 (N_21798,N_21039,N_21126);
nor U21799 (N_21799,N_21172,N_21488);
nand U21800 (N_21800,N_21126,N_21340);
nor U21801 (N_21801,N_21020,N_21152);
nor U21802 (N_21802,N_21338,N_21248);
or U21803 (N_21803,N_21303,N_21335);
and U21804 (N_21804,N_21472,N_21251);
and U21805 (N_21805,N_21248,N_21372);
or U21806 (N_21806,N_21328,N_21081);
nor U21807 (N_21807,N_21324,N_21449);
nor U21808 (N_21808,N_21448,N_21173);
nand U21809 (N_21809,N_21128,N_21316);
nand U21810 (N_21810,N_21443,N_21164);
or U21811 (N_21811,N_21165,N_21078);
and U21812 (N_21812,N_21118,N_21015);
nand U21813 (N_21813,N_21179,N_21336);
and U21814 (N_21814,N_21185,N_21266);
and U21815 (N_21815,N_21069,N_21193);
or U21816 (N_21816,N_21408,N_21339);
nand U21817 (N_21817,N_21495,N_21454);
and U21818 (N_21818,N_21043,N_21020);
and U21819 (N_21819,N_21333,N_21308);
or U21820 (N_21820,N_21131,N_21393);
xnor U21821 (N_21821,N_21323,N_21261);
xnor U21822 (N_21822,N_21072,N_21232);
nor U21823 (N_21823,N_21036,N_21009);
and U21824 (N_21824,N_21072,N_21040);
nor U21825 (N_21825,N_21002,N_21356);
and U21826 (N_21826,N_21075,N_21040);
or U21827 (N_21827,N_21308,N_21442);
nand U21828 (N_21828,N_21244,N_21386);
or U21829 (N_21829,N_21350,N_21470);
or U21830 (N_21830,N_21135,N_21491);
or U21831 (N_21831,N_21444,N_21393);
nor U21832 (N_21832,N_21039,N_21119);
nor U21833 (N_21833,N_21011,N_21435);
or U21834 (N_21834,N_21418,N_21319);
nor U21835 (N_21835,N_21244,N_21352);
and U21836 (N_21836,N_21430,N_21178);
and U21837 (N_21837,N_21167,N_21106);
nand U21838 (N_21838,N_21450,N_21290);
nand U21839 (N_21839,N_21336,N_21491);
nand U21840 (N_21840,N_21024,N_21496);
and U21841 (N_21841,N_21264,N_21244);
nor U21842 (N_21842,N_21260,N_21386);
nand U21843 (N_21843,N_21282,N_21143);
nand U21844 (N_21844,N_21112,N_21393);
nor U21845 (N_21845,N_21201,N_21499);
xor U21846 (N_21846,N_21096,N_21265);
or U21847 (N_21847,N_21130,N_21099);
xnor U21848 (N_21848,N_21348,N_21420);
xor U21849 (N_21849,N_21000,N_21286);
and U21850 (N_21850,N_21400,N_21482);
and U21851 (N_21851,N_21242,N_21328);
or U21852 (N_21852,N_21163,N_21456);
nand U21853 (N_21853,N_21337,N_21267);
nor U21854 (N_21854,N_21274,N_21446);
or U21855 (N_21855,N_21151,N_21216);
or U21856 (N_21856,N_21470,N_21278);
nand U21857 (N_21857,N_21405,N_21482);
nor U21858 (N_21858,N_21101,N_21194);
xor U21859 (N_21859,N_21202,N_21446);
xor U21860 (N_21860,N_21386,N_21452);
and U21861 (N_21861,N_21301,N_21144);
or U21862 (N_21862,N_21332,N_21151);
nand U21863 (N_21863,N_21421,N_21403);
or U21864 (N_21864,N_21200,N_21269);
or U21865 (N_21865,N_21328,N_21378);
and U21866 (N_21866,N_21093,N_21475);
nand U21867 (N_21867,N_21403,N_21415);
nand U21868 (N_21868,N_21175,N_21490);
and U21869 (N_21869,N_21471,N_21261);
nor U21870 (N_21870,N_21010,N_21328);
and U21871 (N_21871,N_21332,N_21446);
or U21872 (N_21872,N_21210,N_21159);
or U21873 (N_21873,N_21448,N_21152);
or U21874 (N_21874,N_21266,N_21186);
and U21875 (N_21875,N_21136,N_21221);
xor U21876 (N_21876,N_21187,N_21052);
and U21877 (N_21877,N_21137,N_21009);
nor U21878 (N_21878,N_21308,N_21387);
or U21879 (N_21879,N_21135,N_21050);
or U21880 (N_21880,N_21287,N_21289);
nor U21881 (N_21881,N_21063,N_21248);
nand U21882 (N_21882,N_21187,N_21022);
nor U21883 (N_21883,N_21335,N_21349);
and U21884 (N_21884,N_21258,N_21213);
and U21885 (N_21885,N_21025,N_21128);
nand U21886 (N_21886,N_21403,N_21114);
xnor U21887 (N_21887,N_21085,N_21182);
and U21888 (N_21888,N_21039,N_21070);
or U21889 (N_21889,N_21355,N_21321);
and U21890 (N_21890,N_21365,N_21145);
nor U21891 (N_21891,N_21141,N_21119);
nand U21892 (N_21892,N_21161,N_21404);
nor U21893 (N_21893,N_21230,N_21288);
and U21894 (N_21894,N_21051,N_21172);
nand U21895 (N_21895,N_21430,N_21244);
nor U21896 (N_21896,N_21345,N_21293);
nand U21897 (N_21897,N_21343,N_21320);
xor U21898 (N_21898,N_21397,N_21417);
nand U21899 (N_21899,N_21462,N_21417);
nor U21900 (N_21900,N_21268,N_21156);
or U21901 (N_21901,N_21367,N_21343);
nand U21902 (N_21902,N_21114,N_21093);
nand U21903 (N_21903,N_21027,N_21406);
nor U21904 (N_21904,N_21287,N_21482);
nor U21905 (N_21905,N_21130,N_21471);
and U21906 (N_21906,N_21212,N_21131);
nand U21907 (N_21907,N_21020,N_21328);
nor U21908 (N_21908,N_21469,N_21452);
nor U21909 (N_21909,N_21442,N_21385);
or U21910 (N_21910,N_21345,N_21379);
nor U21911 (N_21911,N_21224,N_21393);
nand U21912 (N_21912,N_21307,N_21368);
nand U21913 (N_21913,N_21414,N_21243);
or U21914 (N_21914,N_21188,N_21283);
and U21915 (N_21915,N_21086,N_21204);
xnor U21916 (N_21916,N_21449,N_21145);
or U21917 (N_21917,N_21295,N_21468);
nand U21918 (N_21918,N_21012,N_21166);
nand U21919 (N_21919,N_21232,N_21324);
nor U21920 (N_21920,N_21028,N_21303);
and U21921 (N_21921,N_21102,N_21473);
nor U21922 (N_21922,N_21007,N_21328);
and U21923 (N_21923,N_21082,N_21323);
nor U21924 (N_21924,N_21449,N_21300);
or U21925 (N_21925,N_21462,N_21325);
nor U21926 (N_21926,N_21201,N_21068);
nand U21927 (N_21927,N_21475,N_21446);
and U21928 (N_21928,N_21055,N_21303);
and U21929 (N_21929,N_21321,N_21102);
nor U21930 (N_21930,N_21354,N_21007);
and U21931 (N_21931,N_21184,N_21150);
and U21932 (N_21932,N_21230,N_21389);
and U21933 (N_21933,N_21215,N_21353);
or U21934 (N_21934,N_21109,N_21485);
xor U21935 (N_21935,N_21405,N_21492);
xor U21936 (N_21936,N_21049,N_21416);
nor U21937 (N_21937,N_21088,N_21374);
and U21938 (N_21938,N_21327,N_21431);
nor U21939 (N_21939,N_21418,N_21459);
and U21940 (N_21940,N_21445,N_21293);
nand U21941 (N_21941,N_21215,N_21043);
xnor U21942 (N_21942,N_21065,N_21122);
and U21943 (N_21943,N_21152,N_21281);
or U21944 (N_21944,N_21214,N_21045);
and U21945 (N_21945,N_21278,N_21129);
and U21946 (N_21946,N_21124,N_21339);
nand U21947 (N_21947,N_21173,N_21223);
nor U21948 (N_21948,N_21352,N_21061);
or U21949 (N_21949,N_21255,N_21480);
nor U21950 (N_21950,N_21238,N_21420);
nor U21951 (N_21951,N_21430,N_21216);
nand U21952 (N_21952,N_21319,N_21062);
nand U21953 (N_21953,N_21317,N_21361);
nor U21954 (N_21954,N_21027,N_21003);
nor U21955 (N_21955,N_21324,N_21213);
xor U21956 (N_21956,N_21242,N_21498);
nor U21957 (N_21957,N_21034,N_21166);
xnor U21958 (N_21958,N_21429,N_21418);
or U21959 (N_21959,N_21008,N_21124);
and U21960 (N_21960,N_21196,N_21474);
nor U21961 (N_21961,N_21054,N_21193);
nor U21962 (N_21962,N_21136,N_21049);
nor U21963 (N_21963,N_21439,N_21437);
nand U21964 (N_21964,N_21155,N_21167);
and U21965 (N_21965,N_21181,N_21256);
and U21966 (N_21966,N_21412,N_21125);
or U21967 (N_21967,N_21161,N_21122);
and U21968 (N_21968,N_21038,N_21151);
xnor U21969 (N_21969,N_21019,N_21125);
or U21970 (N_21970,N_21155,N_21359);
or U21971 (N_21971,N_21445,N_21011);
xor U21972 (N_21972,N_21402,N_21490);
xnor U21973 (N_21973,N_21161,N_21088);
nor U21974 (N_21974,N_21042,N_21282);
or U21975 (N_21975,N_21141,N_21174);
nand U21976 (N_21976,N_21162,N_21369);
nand U21977 (N_21977,N_21266,N_21246);
nor U21978 (N_21978,N_21256,N_21120);
and U21979 (N_21979,N_21414,N_21216);
nor U21980 (N_21980,N_21183,N_21412);
and U21981 (N_21981,N_21313,N_21150);
nand U21982 (N_21982,N_21268,N_21172);
xor U21983 (N_21983,N_21204,N_21388);
and U21984 (N_21984,N_21266,N_21234);
and U21985 (N_21985,N_21317,N_21330);
or U21986 (N_21986,N_21018,N_21390);
nor U21987 (N_21987,N_21306,N_21104);
nor U21988 (N_21988,N_21098,N_21400);
nor U21989 (N_21989,N_21333,N_21352);
or U21990 (N_21990,N_21302,N_21075);
xor U21991 (N_21991,N_21288,N_21043);
or U21992 (N_21992,N_21276,N_21122);
or U21993 (N_21993,N_21201,N_21060);
or U21994 (N_21994,N_21453,N_21262);
nand U21995 (N_21995,N_21107,N_21095);
nand U21996 (N_21996,N_21119,N_21159);
or U21997 (N_21997,N_21278,N_21246);
and U21998 (N_21998,N_21074,N_21280);
and U21999 (N_21999,N_21405,N_21480);
and U22000 (N_22000,N_21949,N_21694);
or U22001 (N_22001,N_21827,N_21962);
xnor U22002 (N_22002,N_21762,N_21664);
and U22003 (N_22003,N_21638,N_21602);
and U22004 (N_22004,N_21929,N_21566);
and U22005 (N_22005,N_21980,N_21584);
nor U22006 (N_22006,N_21643,N_21511);
nor U22007 (N_22007,N_21658,N_21605);
nand U22008 (N_22008,N_21965,N_21868);
or U22009 (N_22009,N_21577,N_21579);
xor U22010 (N_22010,N_21955,N_21619);
nand U22011 (N_22011,N_21521,N_21812);
and U22012 (N_22012,N_21773,N_21911);
or U22013 (N_22013,N_21876,N_21716);
nor U22014 (N_22014,N_21870,N_21958);
nand U22015 (N_22015,N_21653,N_21981);
nand U22016 (N_22016,N_21938,N_21896);
or U22017 (N_22017,N_21997,N_21842);
xor U22018 (N_22018,N_21571,N_21907);
or U22019 (N_22019,N_21947,N_21708);
nor U22020 (N_22020,N_21613,N_21659);
or U22021 (N_22021,N_21975,N_21701);
and U22022 (N_22022,N_21909,N_21746);
nor U22023 (N_22023,N_21677,N_21927);
or U22024 (N_22024,N_21505,N_21525);
xnor U22025 (N_22025,N_21744,N_21633);
nand U22026 (N_22026,N_21632,N_21730);
nor U22027 (N_22027,N_21751,N_21721);
nor U22028 (N_22028,N_21514,N_21678);
xnor U22029 (N_22029,N_21673,N_21979);
nand U22030 (N_22030,N_21703,N_21946);
nand U22031 (N_22031,N_21686,N_21855);
nor U22032 (N_22032,N_21809,N_21583);
nor U22033 (N_22033,N_21957,N_21867);
nand U22034 (N_22034,N_21826,N_21887);
nand U22035 (N_22035,N_21657,N_21606);
nand U22036 (N_22036,N_21634,N_21555);
xor U22037 (N_22037,N_21596,N_21771);
or U22038 (N_22038,N_21609,N_21931);
or U22039 (N_22039,N_21908,N_21780);
and U22040 (N_22040,N_21551,N_21533);
nor U22041 (N_22041,N_21804,N_21950);
nor U22042 (N_22042,N_21704,N_21848);
and U22043 (N_22043,N_21801,N_21810);
nand U22044 (N_22044,N_21796,N_21996);
nand U22045 (N_22045,N_21737,N_21546);
and U22046 (N_22046,N_21523,N_21894);
or U22047 (N_22047,N_21817,N_21943);
nand U22048 (N_22048,N_21631,N_21942);
nor U22049 (N_22049,N_21699,N_21693);
nor U22050 (N_22050,N_21917,N_21770);
or U22051 (N_22051,N_21528,N_21578);
nand U22052 (N_22052,N_21742,N_21895);
nor U22053 (N_22053,N_21753,N_21562);
nor U22054 (N_22054,N_21984,N_21663);
or U22055 (N_22055,N_21961,N_21545);
or U22056 (N_22056,N_21798,N_21597);
nor U22057 (N_22057,N_21557,N_21871);
and U22058 (N_22058,N_21611,N_21889);
nor U22059 (N_22059,N_21846,N_21850);
nor U22060 (N_22060,N_21718,N_21507);
or U22061 (N_22061,N_21526,N_21539);
or U22062 (N_22062,N_21760,N_21681);
or U22063 (N_22063,N_21941,N_21574);
nand U22064 (N_22064,N_21900,N_21542);
and U22065 (N_22065,N_21860,N_21628);
xor U22066 (N_22066,N_21960,N_21757);
nor U22067 (N_22067,N_21768,N_21527);
and U22068 (N_22068,N_21513,N_21599);
nor U22069 (N_22069,N_21544,N_21992);
or U22070 (N_22070,N_21888,N_21549);
nor U22071 (N_22071,N_21696,N_21873);
or U22072 (N_22072,N_21591,N_21669);
or U22073 (N_22073,N_21783,N_21607);
and U22074 (N_22074,N_21590,N_21541);
or U22075 (N_22075,N_21772,N_21510);
and U22076 (N_22076,N_21923,N_21987);
nor U22077 (N_22077,N_21586,N_21790);
nand U22078 (N_22078,N_21913,N_21710);
or U22079 (N_22079,N_21926,N_21621);
nand U22080 (N_22080,N_21781,N_21624);
nand U22081 (N_22081,N_21794,N_21740);
nand U22082 (N_22082,N_21982,N_21680);
xor U22083 (N_22083,N_21518,N_21792);
or U22084 (N_22084,N_21836,N_21872);
or U22085 (N_22085,N_21723,N_21788);
nand U22086 (N_22086,N_21709,N_21558);
and U22087 (N_22087,N_21642,N_21845);
and U22088 (N_22088,N_21512,N_21959);
nand U22089 (N_22089,N_21930,N_21592);
and U22090 (N_22090,N_21805,N_21722);
nor U22091 (N_22091,N_21660,N_21815);
nor U22092 (N_22092,N_21822,N_21536);
and U22093 (N_22093,N_21806,N_21994);
nand U22094 (N_22094,N_21687,N_21635);
xnor U22095 (N_22095,N_21830,N_21530);
nand U22096 (N_22096,N_21884,N_21754);
or U22097 (N_22097,N_21844,N_21899);
or U22098 (N_22098,N_21503,N_21875);
nand U22099 (N_22099,N_21919,N_21682);
nand U22100 (N_22100,N_21799,N_21793);
nand U22101 (N_22101,N_21777,N_21779);
or U22102 (N_22102,N_21978,N_21874);
xor U22103 (N_22103,N_21552,N_21626);
and U22104 (N_22104,N_21862,N_21838);
or U22105 (N_22105,N_21849,N_21568);
and U22106 (N_22106,N_21890,N_21623);
nand U22107 (N_22107,N_21559,N_21985);
and U22108 (N_22108,N_21967,N_21863);
or U22109 (N_22109,N_21969,N_21733);
and U22110 (N_22110,N_21648,N_21707);
nor U22111 (N_22111,N_21936,N_21755);
nand U22112 (N_22112,N_21556,N_21553);
and U22113 (N_22113,N_21501,N_21977);
xor U22114 (N_22114,N_21999,N_21594);
and U22115 (N_22115,N_21688,N_21904);
or U22116 (N_22116,N_21925,N_21697);
xnor U22117 (N_22117,N_21647,N_21614);
nor U22118 (N_22118,N_21531,N_21778);
nor U22119 (N_22119,N_21901,N_21921);
and U22120 (N_22120,N_21561,N_21517);
nor U22121 (N_22121,N_21902,N_21854);
or U22122 (N_22122,N_21665,N_21750);
and U22123 (N_22123,N_21565,N_21878);
nand U22124 (N_22124,N_21720,N_21670);
nor U22125 (N_22125,N_21524,N_21719);
or U22126 (N_22126,N_21627,N_21729);
or U22127 (N_22127,N_21934,N_21581);
and U22128 (N_22128,N_21775,N_21617);
or U22129 (N_22129,N_21615,N_21550);
or U22130 (N_22130,N_21749,N_21535);
or U22131 (N_22131,N_21906,N_21666);
nand U22132 (N_22132,N_21933,N_21835);
and U22133 (N_22133,N_21713,N_21646);
nand U22134 (N_22134,N_21974,N_21612);
and U22135 (N_22135,N_21567,N_21784);
or U22136 (N_22136,N_21995,N_21944);
xor U22137 (N_22137,N_21679,N_21851);
or U22138 (N_22138,N_21522,N_21808);
nor U22139 (N_22139,N_21832,N_21534);
nand U22140 (N_22140,N_21725,N_21714);
or U22141 (N_22141,N_21645,N_21912);
and U22142 (N_22142,N_21575,N_21573);
xor U22143 (N_22143,N_21509,N_21973);
nor U22144 (N_22144,N_21758,N_21857);
or U22145 (N_22145,N_21728,N_21859);
nand U22146 (N_22146,N_21829,N_21502);
and U22147 (N_22147,N_21672,N_21706);
or U22148 (N_22148,N_21690,N_21731);
and U22149 (N_22149,N_21695,N_21765);
nand U22150 (N_22150,N_21864,N_21988);
and U22151 (N_22151,N_21971,N_21698);
and U22152 (N_22152,N_21986,N_21655);
xor U22153 (N_22153,N_21585,N_21877);
or U22154 (N_22154,N_21589,N_21785);
or U22155 (N_22155,N_21797,N_21764);
nor U22156 (N_22156,N_21903,N_21736);
nor U22157 (N_22157,N_21791,N_21756);
nand U22158 (N_22158,N_21519,N_21630);
nor U22159 (N_22159,N_21869,N_21735);
nand U22160 (N_22160,N_21662,N_21625);
nor U22161 (N_22161,N_21937,N_21563);
nor U22162 (N_22162,N_21789,N_21782);
or U22163 (N_22163,N_21689,N_21580);
or U22164 (N_22164,N_21920,N_21516);
or U22165 (N_22165,N_21861,N_21560);
or U22166 (N_22166,N_21548,N_21604);
or U22167 (N_22167,N_21824,N_21910);
or U22168 (N_22168,N_21508,N_21554);
nor U22169 (N_22169,N_21572,N_21892);
or U22170 (N_22170,N_21712,N_21833);
or U22171 (N_22171,N_21595,N_21841);
nor U22172 (N_22172,N_21963,N_21656);
xor U22173 (N_22173,N_21989,N_21667);
and U22174 (N_22174,N_21674,N_21547);
and U22175 (N_22175,N_21821,N_21993);
and U22176 (N_22176,N_21825,N_21811);
xnor U22177 (N_22177,N_21940,N_21671);
nor U22178 (N_22178,N_21651,N_21972);
or U22179 (N_22179,N_21598,N_21897);
nand U22180 (N_22180,N_21569,N_21748);
and U22181 (N_22181,N_21905,N_21898);
and U22182 (N_22182,N_21739,N_21676);
and U22183 (N_22183,N_21847,N_21866);
xor U22184 (N_22184,N_21640,N_21803);
xnor U22185 (N_22185,N_21620,N_21776);
nor U22186 (N_22186,N_21883,N_21795);
nand U22187 (N_22187,N_21787,N_21652);
and U22188 (N_22188,N_21691,N_21570);
or U22189 (N_22189,N_21865,N_21767);
nor U22190 (N_22190,N_21880,N_21564);
nand U22191 (N_22191,N_21763,N_21685);
or U22192 (N_22192,N_21727,N_21831);
xnor U22193 (N_22193,N_21818,N_21928);
xor U22194 (N_22194,N_21610,N_21891);
nor U22195 (N_22195,N_21816,N_21668);
nor U22196 (N_22196,N_21951,N_21636);
or U22197 (N_22197,N_21800,N_21692);
nor U22198 (N_22198,N_21600,N_21622);
xor U22199 (N_22199,N_21837,N_21774);
nand U22200 (N_22200,N_21576,N_21705);
and U22201 (N_22201,N_21601,N_21948);
and U22202 (N_22202,N_21840,N_21843);
xor U22203 (N_22203,N_21587,N_21715);
or U22204 (N_22204,N_21807,N_21644);
or U22205 (N_22205,N_21814,N_21922);
xor U22206 (N_22206,N_21820,N_21956);
nand U22207 (N_22207,N_21649,N_21603);
nor U22208 (N_22208,N_21700,N_21537);
nand U22209 (N_22209,N_21761,N_21769);
and U22210 (N_22210,N_21886,N_21734);
nor U22211 (N_22211,N_21743,N_21918);
and U22212 (N_22212,N_21914,N_21813);
and U22213 (N_22213,N_21856,N_21717);
and U22214 (N_22214,N_21879,N_21637);
or U22215 (N_22215,N_21654,N_21802);
nand U22216 (N_22216,N_21882,N_21702);
xnor U22217 (N_22217,N_21885,N_21954);
nand U22218 (N_22218,N_21532,N_21983);
nand U22219 (N_22219,N_21991,N_21766);
nand U22220 (N_22220,N_21819,N_21945);
or U22221 (N_22221,N_21745,N_21504);
or U22222 (N_22222,N_21747,N_21538);
nor U22223 (N_22223,N_21966,N_21506);
or U22224 (N_22224,N_21582,N_21608);
nor U22225 (N_22225,N_21529,N_21752);
nor U22226 (N_22226,N_21939,N_21970);
and U22227 (N_22227,N_21998,N_21675);
nor U22228 (N_22228,N_21520,N_21853);
and U22229 (N_22229,N_21732,N_21932);
xor U22230 (N_22230,N_21588,N_21500);
nor U22231 (N_22231,N_21839,N_21641);
and U22232 (N_22232,N_21711,N_21616);
and U22233 (N_22233,N_21759,N_21593);
nor U22234 (N_22234,N_21952,N_21786);
or U22235 (N_22235,N_21823,N_21684);
and U22236 (N_22236,N_21661,N_21726);
and U22237 (N_22237,N_21543,N_21953);
or U22238 (N_22238,N_21852,N_21515);
nand U22239 (N_22239,N_21935,N_21968);
and U22240 (N_22240,N_21650,N_21639);
nand U22241 (N_22241,N_21881,N_21618);
nand U22242 (N_22242,N_21540,N_21741);
and U22243 (N_22243,N_21964,N_21724);
or U22244 (N_22244,N_21834,N_21858);
and U22245 (N_22245,N_21990,N_21893);
nor U22246 (N_22246,N_21629,N_21828);
nor U22247 (N_22247,N_21738,N_21915);
and U22248 (N_22248,N_21976,N_21683);
and U22249 (N_22249,N_21924,N_21916);
nand U22250 (N_22250,N_21713,N_21641);
nor U22251 (N_22251,N_21789,N_21687);
nand U22252 (N_22252,N_21836,N_21784);
xor U22253 (N_22253,N_21780,N_21584);
and U22254 (N_22254,N_21818,N_21802);
or U22255 (N_22255,N_21585,N_21692);
nand U22256 (N_22256,N_21984,N_21763);
or U22257 (N_22257,N_21960,N_21598);
nor U22258 (N_22258,N_21594,N_21629);
nand U22259 (N_22259,N_21718,N_21880);
nor U22260 (N_22260,N_21542,N_21846);
nor U22261 (N_22261,N_21935,N_21830);
nor U22262 (N_22262,N_21653,N_21907);
or U22263 (N_22263,N_21517,N_21909);
nand U22264 (N_22264,N_21980,N_21721);
nor U22265 (N_22265,N_21989,N_21624);
and U22266 (N_22266,N_21787,N_21853);
or U22267 (N_22267,N_21863,N_21547);
nand U22268 (N_22268,N_21533,N_21929);
nor U22269 (N_22269,N_21629,N_21553);
nor U22270 (N_22270,N_21728,N_21751);
nor U22271 (N_22271,N_21537,N_21667);
nor U22272 (N_22272,N_21959,N_21678);
or U22273 (N_22273,N_21672,N_21726);
and U22274 (N_22274,N_21593,N_21943);
nor U22275 (N_22275,N_21787,N_21965);
or U22276 (N_22276,N_21975,N_21992);
or U22277 (N_22277,N_21847,N_21710);
nand U22278 (N_22278,N_21809,N_21591);
and U22279 (N_22279,N_21720,N_21534);
xor U22280 (N_22280,N_21716,N_21880);
or U22281 (N_22281,N_21718,N_21645);
or U22282 (N_22282,N_21748,N_21888);
and U22283 (N_22283,N_21718,N_21620);
or U22284 (N_22284,N_21959,N_21982);
nand U22285 (N_22285,N_21740,N_21593);
nor U22286 (N_22286,N_21674,N_21838);
nand U22287 (N_22287,N_21981,N_21679);
nor U22288 (N_22288,N_21799,N_21581);
or U22289 (N_22289,N_21544,N_21763);
xnor U22290 (N_22290,N_21811,N_21864);
nand U22291 (N_22291,N_21760,N_21959);
nand U22292 (N_22292,N_21563,N_21637);
nor U22293 (N_22293,N_21784,N_21712);
nand U22294 (N_22294,N_21505,N_21735);
nor U22295 (N_22295,N_21853,N_21623);
xor U22296 (N_22296,N_21768,N_21760);
xnor U22297 (N_22297,N_21953,N_21787);
or U22298 (N_22298,N_21942,N_21501);
nand U22299 (N_22299,N_21832,N_21793);
and U22300 (N_22300,N_21801,N_21578);
nand U22301 (N_22301,N_21738,N_21841);
and U22302 (N_22302,N_21774,N_21542);
nand U22303 (N_22303,N_21748,N_21759);
or U22304 (N_22304,N_21770,N_21994);
nor U22305 (N_22305,N_21606,N_21878);
xnor U22306 (N_22306,N_21956,N_21844);
and U22307 (N_22307,N_21568,N_21985);
xnor U22308 (N_22308,N_21524,N_21547);
xor U22309 (N_22309,N_21697,N_21578);
or U22310 (N_22310,N_21536,N_21720);
or U22311 (N_22311,N_21866,N_21680);
and U22312 (N_22312,N_21984,N_21564);
nor U22313 (N_22313,N_21948,N_21585);
and U22314 (N_22314,N_21873,N_21979);
xor U22315 (N_22315,N_21753,N_21844);
xor U22316 (N_22316,N_21835,N_21996);
or U22317 (N_22317,N_21631,N_21896);
or U22318 (N_22318,N_21612,N_21652);
and U22319 (N_22319,N_21969,N_21541);
and U22320 (N_22320,N_21766,N_21976);
nor U22321 (N_22321,N_21639,N_21837);
nand U22322 (N_22322,N_21534,N_21823);
and U22323 (N_22323,N_21677,N_21615);
and U22324 (N_22324,N_21698,N_21634);
nor U22325 (N_22325,N_21661,N_21978);
nor U22326 (N_22326,N_21521,N_21648);
nand U22327 (N_22327,N_21812,N_21971);
nand U22328 (N_22328,N_21516,N_21945);
and U22329 (N_22329,N_21704,N_21894);
nand U22330 (N_22330,N_21515,N_21568);
and U22331 (N_22331,N_21867,N_21966);
and U22332 (N_22332,N_21960,N_21640);
nor U22333 (N_22333,N_21861,N_21942);
nand U22334 (N_22334,N_21759,N_21803);
or U22335 (N_22335,N_21581,N_21715);
or U22336 (N_22336,N_21977,N_21706);
nor U22337 (N_22337,N_21994,N_21740);
nand U22338 (N_22338,N_21747,N_21769);
nand U22339 (N_22339,N_21930,N_21607);
nor U22340 (N_22340,N_21991,N_21566);
or U22341 (N_22341,N_21832,N_21648);
or U22342 (N_22342,N_21687,N_21805);
or U22343 (N_22343,N_21607,N_21633);
or U22344 (N_22344,N_21837,N_21985);
and U22345 (N_22345,N_21582,N_21661);
nand U22346 (N_22346,N_21648,N_21886);
nand U22347 (N_22347,N_21540,N_21718);
nor U22348 (N_22348,N_21504,N_21719);
and U22349 (N_22349,N_21651,N_21831);
nor U22350 (N_22350,N_21811,N_21856);
nor U22351 (N_22351,N_21670,N_21535);
and U22352 (N_22352,N_21748,N_21683);
or U22353 (N_22353,N_21730,N_21941);
or U22354 (N_22354,N_21914,N_21648);
nor U22355 (N_22355,N_21557,N_21977);
nand U22356 (N_22356,N_21627,N_21663);
nand U22357 (N_22357,N_21882,N_21648);
and U22358 (N_22358,N_21869,N_21797);
xor U22359 (N_22359,N_21617,N_21755);
or U22360 (N_22360,N_21921,N_21729);
xor U22361 (N_22361,N_21735,N_21651);
nand U22362 (N_22362,N_21615,N_21951);
xnor U22363 (N_22363,N_21706,N_21625);
or U22364 (N_22364,N_21504,N_21620);
nand U22365 (N_22365,N_21642,N_21953);
nand U22366 (N_22366,N_21902,N_21502);
and U22367 (N_22367,N_21595,N_21923);
nand U22368 (N_22368,N_21576,N_21821);
or U22369 (N_22369,N_21825,N_21778);
nor U22370 (N_22370,N_21644,N_21862);
or U22371 (N_22371,N_21979,N_21847);
or U22372 (N_22372,N_21737,N_21848);
nand U22373 (N_22373,N_21904,N_21796);
nand U22374 (N_22374,N_21930,N_21738);
nor U22375 (N_22375,N_21923,N_21796);
xnor U22376 (N_22376,N_21723,N_21917);
nand U22377 (N_22377,N_21814,N_21723);
or U22378 (N_22378,N_21650,N_21695);
nand U22379 (N_22379,N_21764,N_21812);
or U22380 (N_22380,N_21619,N_21948);
nand U22381 (N_22381,N_21883,N_21706);
xor U22382 (N_22382,N_21893,N_21641);
nand U22383 (N_22383,N_21879,N_21538);
nand U22384 (N_22384,N_21660,N_21829);
and U22385 (N_22385,N_21706,N_21522);
nand U22386 (N_22386,N_21712,N_21930);
or U22387 (N_22387,N_21502,N_21870);
nor U22388 (N_22388,N_21635,N_21717);
xor U22389 (N_22389,N_21943,N_21885);
or U22390 (N_22390,N_21821,N_21769);
or U22391 (N_22391,N_21625,N_21863);
or U22392 (N_22392,N_21846,N_21658);
nand U22393 (N_22393,N_21688,N_21925);
nor U22394 (N_22394,N_21736,N_21932);
nor U22395 (N_22395,N_21960,N_21993);
nand U22396 (N_22396,N_21866,N_21883);
nor U22397 (N_22397,N_21873,N_21585);
nor U22398 (N_22398,N_21853,N_21867);
xor U22399 (N_22399,N_21528,N_21592);
and U22400 (N_22400,N_21588,N_21751);
and U22401 (N_22401,N_21649,N_21870);
and U22402 (N_22402,N_21777,N_21927);
and U22403 (N_22403,N_21860,N_21776);
or U22404 (N_22404,N_21825,N_21933);
and U22405 (N_22405,N_21892,N_21584);
or U22406 (N_22406,N_21910,N_21947);
and U22407 (N_22407,N_21703,N_21515);
nor U22408 (N_22408,N_21996,N_21886);
or U22409 (N_22409,N_21834,N_21678);
or U22410 (N_22410,N_21589,N_21858);
and U22411 (N_22411,N_21872,N_21552);
nand U22412 (N_22412,N_21772,N_21643);
nor U22413 (N_22413,N_21613,N_21585);
nand U22414 (N_22414,N_21789,N_21929);
nand U22415 (N_22415,N_21966,N_21797);
or U22416 (N_22416,N_21669,N_21572);
and U22417 (N_22417,N_21681,N_21672);
or U22418 (N_22418,N_21848,N_21962);
nand U22419 (N_22419,N_21870,N_21683);
nor U22420 (N_22420,N_21631,N_21808);
or U22421 (N_22421,N_21525,N_21788);
and U22422 (N_22422,N_21521,N_21759);
and U22423 (N_22423,N_21778,N_21987);
nor U22424 (N_22424,N_21962,N_21511);
and U22425 (N_22425,N_21578,N_21658);
and U22426 (N_22426,N_21728,N_21733);
nand U22427 (N_22427,N_21667,N_21978);
nor U22428 (N_22428,N_21902,N_21651);
or U22429 (N_22429,N_21659,N_21527);
or U22430 (N_22430,N_21784,N_21597);
or U22431 (N_22431,N_21772,N_21644);
nand U22432 (N_22432,N_21810,N_21912);
nand U22433 (N_22433,N_21912,N_21930);
and U22434 (N_22434,N_21694,N_21858);
nand U22435 (N_22435,N_21609,N_21646);
nor U22436 (N_22436,N_21751,N_21605);
and U22437 (N_22437,N_21801,N_21910);
xnor U22438 (N_22438,N_21907,N_21783);
nand U22439 (N_22439,N_21647,N_21828);
and U22440 (N_22440,N_21855,N_21906);
or U22441 (N_22441,N_21726,N_21916);
and U22442 (N_22442,N_21892,N_21663);
or U22443 (N_22443,N_21737,N_21709);
or U22444 (N_22444,N_21734,N_21588);
or U22445 (N_22445,N_21753,N_21781);
and U22446 (N_22446,N_21883,N_21932);
or U22447 (N_22447,N_21976,N_21986);
nand U22448 (N_22448,N_21705,N_21661);
nand U22449 (N_22449,N_21669,N_21694);
nand U22450 (N_22450,N_21980,N_21914);
or U22451 (N_22451,N_21516,N_21581);
or U22452 (N_22452,N_21574,N_21938);
nand U22453 (N_22453,N_21779,N_21727);
nand U22454 (N_22454,N_21686,N_21556);
nand U22455 (N_22455,N_21947,N_21963);
xnor U22456 (N_22456,N_21951,N_21959);
nand U22457 (N_22457,N_21996,N_21519);
nand U22458 (N_22458,N_21790,N_21694);
nor U22459 (N_22459,N_21857,N_21966);
nand U22460 (N_22460,N_21505,N_21949);
or U22461 (N_22461,N_21563,N_21682);
and U22462 (N_22462,N_21574,N_21950);
xor U22463 (N_22463,N_21594,N_21945);
nor U22464 (N_22464,N_21565,N_21959);
and U22465 (N_22465,N_21655,N_21786);
and U22466 (N_22466,N_21813,N_21641);
xor U22467 (N_22467,N_21902,N_21774);
and U22468 (N_22468,N_21691,N_21983);
xnor U22469 (N_22469,N_21993,N_21636);
nor U22470 (N_22470,N_21500,N_21529);
nand U22471 (N_22471,N_21533,N_21740);
xnor U22472 (N_22472,N_21594,N_21534);
nand U22473 (N_22473,N_21578,N_21710);
nand U22474 (N_22474,N_21736,N_21609);
nor U22475 (N_22475,N_21764,N_21890);
or U22476 (N_22476,N_21682,N_21676);
nand U22477 (N_22477,N_21592,N_21726);
and U22478 (N_22478,N_21706,N_21984);
nand U22479 (N_22479,N_21946,N_21816);
nand U22480 (N_22480,N_21921,N_21544);
nand U22481 (N_22481,N_21769,N_21730);
and U22482 (N_22482,N_21889,N_21595);
nand U22483 (N_22483,N_21959,N_21767);
or U22484 (N_22484,N_21596,N_21556);
nand U22485 (N_22485,N_21664,N_21976);
xor U22486 (N_22486,N_21586,N_21948);
and U22487 (N_22487,N_21805,N_21858);
or U22488 (N_22488,N_21660,N_21582);
and U22489 (N_22489,N_21710,N_21560);
and U22490 (N_22490,N_21576,N_21557);
and U22491 (N_22491,N_21849,N_21914);
nor U22492 (N_22492,N_21803,N_21771);
and U22493 (N_22493,N_21962,N_21580);
nor U22494 (N_22494,N_21875,N_21770);
and U22495 (N_22495,N_21647,N_21978);
nand U22496 (N_22496,N_21562,N_21863);
xor U22497 (N_22497,N_21773,N_21728);
or U22498 (N_22498,N_21568,N_21824);
and U22499 (N_22499,N_21527,N_21939);
and U22500 (N_22500,N_22381,N_22401);
nor U22501 (N_22501,N_22222,N_22122);
and U22502 (N_22502,N_22166,N_22295);
and U22503 (N_22503,N_22125,N_22104);
xnor U22504 (N_22504,N_22250,N_22177);
or U22505 (N_22505,N_22073,N_22282);
and U22506 (N_22506,N_22397,N_22236);
and U22507 (N_22507,N_22372,N_22227);
and U22508 (N_22508,N_22064,N_22367);
nand U22509 (N_22509,N_22290,N_22441);
nor U22510 (N_22510,N_22330,N_22285);
nand U22511 (N_22511,N_22402,N_22395);
nand U22512 (N_22512,N_22337,N_22280);
nand U22513 (N_22513,N_22314,N_22034);
nor U22514 (N_22514,N_22208,N_22297);
nand U22515 (N_22515,N_22331,N_22488);
nand U22516 (N_22516,N_22086,N_22018);
nor U22517 (N_22517,N_22213,N_22007);
or U22518 (N_22518,N_22193,N_22374);
nor U22519 (N_22519,N_22003,N_22077);
nor U22520 (N_22520,N_22316,N_22145);
and U22521 (N_22521,N_22462,N_22202);
nand U22522 (N_22522,N_22065,N_22132);
or U22523 (N_22523,N_22383,N_22257);
nor U22524 (N_22524,N_22014,N_22309);
and U22525 (N_22525,N_22407,N_22161);
nand U22526 (N_22526,N_22475,N_22030);
and U22527 (N_22527,N_22165,N_22151);
and U22528 (N_22528,N_22042,N_22420);
nand U22529 (N_22529,N_22017,N_22090);
xnor U22530 (N_22530,N_22084,N_22204);
nand U22531 (N_22531,N_22072,N_22430);
or U22532 (N_22532,N_22069,N_22218);
or U22533 (N_22533,N_22300,N_22341);
or U22534 (N_22534,N_22413,N_22063);
nor U22535 (N_22535,N_22240,N_22472);
nor U22536 (N_22536,N_22192,N_22016);
nor U22537 (N_22537,N_22150,N_22378);
or U22538 (N_22538,N_22487,N_22276);
and U22539 (N_22539,N_22028,N_22264);
or U22540 (N_22540,N_22209,N_22414);
nor U22541 (N_22541,N_22451,N_22153);
and U22542 (N_22542,N_22343,N_22066);
nor U22543 (N_22543,N_22356,N_22113);
nand U22544 (N_22544,N_22274,N_22267);
nand U22545 (N_22545,N_22083,N_22326);
and U22546 (N_22546,N_22121,N_22091);
or U22547 (N_22547,N_22147,N_22307);
and U22548 (N_22548,N_22043,N_22315);
xnor U22549 (N_22549,N_22178,N_22245);
or U22550 (N_22550,N_22325,N_22220);
and U22551 (N_22551,N_22011,N_22020);
or U22552 (N_22552,N_22498,N_22163);
nand U22553 (N_22553,N_22100,N_22186);
or U22554 (N_22554,N_22001,N_22155);
nor U22555 (N_22555,N_22275,N_22459);
nor U22556 (N_22556,N_22425,N_22371);
or U22557 (N_22557,N_22226,N_22123);
nand U22558 (N_22558,N_22133,N_22393);
nand U22559 (N_22559,N_22434,N_22143);
xnor U22560 (N_22560,N_22468,N_22490);
and U22561 (N_22561,N_22474,N_22061);
nor U22562 (N_22562,N_22060,N_22197);
xor U22563 (N_22563,N_22156,N_22005);
xor U22564 (N_22564,N_22409,N_22461);
and U22565 (N_22565,N_22362,N_22056);
or U22566 (N_22566,N_22444,N_22266);
nor U22567 (N_22567,N_22366,N_22067);
or U22568 (N_22568,N_22438,N_22495);
nand U22569 (N_22569,N_22114,N_22046);
nand U22570 (N_22570,N_22242,N_22026);
and U22571 (N_22571,N_22312,N_22184);
and U22572 (N_22572,N_22134,N_22491);
nor U22573 (N_22573,N_22480,N_22399);
nor U22574 (N_22574,N_22433,N_22196);
and U22575 (N_22575,N_22247,N_22070);
nor U22576 (N_22576,N_22023,N_22322);
and U22577 (N_22577,N_22207,N_22336);
and U22578 (N_22578,N_22469,N_22308);
or U22579 (N_22579,N_22363,N_22442);
and U22580 (N_22580,N_22162,N_22353);
nor U22581 (N_22581,N_22416,N_22484);
nor U22582 (N_22582,N_22439,N_22109);
nand U22583 (N_22583,N_22176,N_22376);
and U22584 (N_22584,N_22085,N_22164);
and U22585 (N_22585,N_22251,N_22486);
and U22586 (N_22586,N_22033,N_22179);
nand U22587 (N_22587,N_22010,N_22059);
and U22588 (N_22588,N_22105,N_22327);
nor U22589 (N_22589,N_22172,N_22265);
and U22590 (N_22590,N_22306,N_22473);
nor U22591 (N_22591,N_22144,N_22201);
or U22592 (N_22592,N_22110,N_22294);
and U22593 (N_22593,N_22406,N_22435);
or U22594 (N_22594,N_22385,N_22195);
xnor U22595 (N_22595,N_22483,N_22169);
nand U22596 (N_22596,N_22149,N_22263);
nor U22597 (N_22597,N_22032,N_22157);
nand U22598 (N_22598,N_22270,N_22446);
nor U22599 (N_22599,N_22004,N_22291);
nor U22600 (N_22600,N_22349,N_22203);
nor U22601 (N_22601,N_22148,N_22478);
nor U22602 (N_22602,N_22025,N_22310);
and U22603 (N_22603,N_22106,N_22479);
nand U22604 (N_22604,N_22183,N_22449);
nor U22605 (N_22605,N_22055,N_22008);
and U22606 (N_22606,N_22443,N_22130);
and U22607 (N_22607,N_22191,N_22448);
and U22608 (N_22608,N_22051,N_22403);
or U22609 (N_22609,N_22277,N_22317);
and U22610 (N_22610,N_22037,N_22129);
nand U22611 (N_22611,N_22492,N_22233);
or U22612 (N_22612,N_22131,N_22002);
nand U22613 (N_22613,N_22256,N_22394);
nor U22614 (N_22614,N_22292,N_22380);
nand U22615 (N_22615,N_22424,N_22225);
or U22616 (N_22616,N_22296,N_22189);
xnor U22617 (N_22617,N_22111,N_22224);
xnor U22618 (N_22618,N_22058,N_22389);
or U22619 (N_22619,N_22467,N_22255);
nor U22620 (N_22620,N_22239,N_22452);
nand U22621 (N_22621,N_22365,N_22049);
or U22622 (N_22622,N_22436,N_22334);
xor U22623 (N_22623,N_22136,N_22035);
and U22624 (N_22624,N_22152,N_22135);
nor U22625 (N_22625,N_22278,N_22068);
xnor U22626 (N_22626,N_22421,N_22128);
or U22627 (N_22627,N_22426,N_22215);
and U22628 (N_22628,N_22158,N_22415);
and U22629 (N_22629,N_22238,N_22221);
and U22630 (N_22630,N_22427,N_22199);
or U22631 (N_22631,N_22379,N_22369);
or U22632 (N_22632,N_22454,N_22329);
nand U22633 (N_22633,N_22344,N_22006);
or U22634 (N_22634,N_22351,N_22279);
xor U22635 (N_22635,N_22481,N_22477);
nand U22636 (N_22636,N_22321,N_22429);
and U22637 (N_22637,N_22194,N_22261);
xor U22638 (N_22638,N_22140,N_22000);
and U22639 (N_22639,N_22460,N_22418);
nand U22640 (N_22640,N_22180,N_22071);
nor U22641 (N_22641,N_22107,N_22392);
or U22642 (N_22642,N_22160,N_22340);
or U22643 (N_22643,N_22181,N_22476);
nor U22644 (N_22644,N_22029,N_22092);
and U22645 (N_22645,N_22360,N_22246);
nor U22646 (N_22646,N_22405,N_22400);
nand U22647 (N_22647,N_22120,N_22087);
or U22648 (N_22648,N_22455,N_22062);
xor U22649 (N_22649,N_22410,N_22137);
or U22650 (N_22650,N_22283,N_22262);
or U22651 (N_22651,N_22496,N_22387);
or U22652 (N_22652,N_22214,N_22054);
nand U22653 (N_22653,N_22471,N_22258);
or U22654 (N_22654,N_22457,N_22345);
and U22655 (N_22655,N_22234,N_22388);
and U22656 (N_22656,N_22039,N_22335);
or U22657 (N_22657,N_22045,N_22252);
and U22658 (N_22658,N_22445,N_22338);
nand U22659 (N_22659,N_22319,N_22040);
or U22660 (N_22660,N_22463,N_22235);
and U22661 (N_22661,N_22038,N_22053);
nor U22662 (N_22662,N_22313,N_22089);
xnor U22663 (N_22663,N_22081,N_22364);
or U22664 (N_22664,N_22119,N_22223);
nand U22665 (N_22665,N_22361,N_22352);
nor U22666 (N_22666,N_22117,N_22108);
nor U22667 (N_22667,N_22219,N_22050);
and U22668 (N_22668,N_22103,N_22303);
nor U22669 (N_22669,N_22431,N_22447);
and U22670 (N_22670,N_22346,N_22302);
nor U22671 (N_22671,N_22244,N_22422);
nor U22672 (N_22672,N_22499,N_22182);
nor U22673 (N_22673,N_22021,N_22287);
nor U22674 (N_22674,N_22022,N_22357);
and U22675 (N_22675,N_22428,N_22370);
xnor U22676 (N_22676,N_22289,N_22146);
xor U22677 (N_22677,N_22013,N_22269);
xnor U22678 (N_22678,N_22171,N_22228);
and U22679 (N_22679,N_22355,N_22347);
nand U22680 (N_22680,N_22304,N_22118);
or U22681 (N_22681,N_22411,N_22206);
or U22682 (N_22682,N_22154,N_22368);
and U22683 (N_22683,N_22241,N_22332);
nand U22684 (N_22684,N_22350,N_22027);
and U22685 (N_22685,N_22324,N_22254);
and U22686 (N_22686,N_22281,N_22205);
nand U22687 (N_22687,N_22485,N_22139);
xnor U22688 (N_22688,N_22074,N_22138);
or U22689 (N_22689,N_22273,N_22339);
xnor U22690 (N_22690,N_22408,N_22286);
nand U22691 (N_22691,N_22078,N_22019);
xor U22692 (N_22692,N_22465,N_22124);
and U22693 (N_22693,N_22015,N_22079);
and U22694 (N_22694,N_22311,N_22057);
xnor U22695 (N_22695,N_22432,N_22450);
nand U22696 (N_22696,N_22482,N_22101);
and U22697 (N_22697,N_22440,N_22456);
and U22698 (N_22698,N_22096,N_22384);
nor U22699 (N_22699,N_22348,N_22359);
or U22700 (N_22700,N_22386,N_22052);
nand U22701 (N_22701,N_22116,N_22260);
nand U22702 (N_22702,N_22493,N_22047);
xnor U22703 (N_22703,N_22417,N_22185);
nor U22704 (N_22704,N_22230,N_22099);
nand U22705 (N_22705,N_22095,N_22396);
and U22706 (N_22706,N_22249,N_22142);
and U22707 (N_22707,N_22423,N_22377);
and U22708 (N_22708,N_22284,N_22453);
xnor U22709 (N_22709,N_22198,N_22097);
xor U22710 (N_22710,N_22323,N_22093);
nor U22711 (N_22711,N_22098,N_22259);
and U22712 (N_22712,N_22305,N_22088);
nand U22713 (N_22713,N_22012,N_22458);
nand U22714 (N_22714,N_22094,N_22318);
nand U22715 (N_22715,N_22187,N_22141);
nand U22716 (N_22716,N_22489,N_22112);
nor U22717 (N_22717,N_22390,N_22075);
nand U22718 (N_22718,N_22272,N_22080);
and U22719 (N_22719,N_22293,N_22174);
nor U22720 (N_22720,N_22404,N_22382);
and U22721 (N_22721,N_22298,N_22328);
and U22722 (N_22722,N_22212,N_22217);
nand U22723 (N_22723,N_22391,N_22115);
nor U22724 (N_22724,N_22188,N_22082);
and U22725 (N_22725,N_22048,N_22036);
nand U22726 (N_22726,N_22200,N_22271);
nor U22727 (N_22727,N_22253,N_22466);
nand U22728 (N_22728,N_22248,N_22301);
nand U22729 (N_22729,N_22358,N_22102);
and U22730 (N_22730,N_22237,N_22373);
nand U22731 (N_22731,N_22216,N_22211);
and U22732 (N_22732,N_22333,N_22243);
nand U22733 (N_22733,N_22076,N_22470);
nor U22734 (N_22734,N_22229,N_22170);
and U22735 (N_22735,N_22354,N_22127);
nor U22736 (N_22736,N_22210,N_22288);
or U22737 (N_22737,N_22041,N_22437);
or U22738 (N_22738,N_22342,N_22494);
or U22739 (N_22739,N_22299,N_22168);
or U22740 (N_22740,N_22024,N_22268);
xnor U22741 (N_22741,N_22190,N_22126);
nor U22742 (N_22742,N_22231,N_22173);
xnor U22743 (N_22743,N_22009,N_22497);
or U22744 (N_22744,N_22175,N_22320);
nor U22745 (N_22745,N_22044,N_22375);
nor U22746 (N_22746,N_22464,N_22232);
and U22747 (N_22747,N_22159,N_22412);
nand U22748 (N_22748,N_22419,N_22031);
or U22749 (N_22749,N_22167,N_22398);
and U22750 (N_22750,N_22493,N_22103);
nor U22751 (N_22751,N_22385,N_22450);
nor U22752 (N_22752,N_22268,N_22143);
or U22753 (N_22753,N_22066,N_22406);
or U22754 (N_22754,N_22125,N_22046);
and U22755 (N_22755,N_22392,N_22015);
or U22756 (N_22756,N_22357,N_22152);
or U22757 (N_22757,N_22136,N_22104);
nor U22758 (N_22758,N_22156,N_22006);
and U22759 (N_22759,N_22218,N_22458);
nand U22760 (N_22760,N_22274,N_22150);
and U22761 (N_22761,N_22447,N_22487);
or U22762 (N_22762,N_22020,N_22461);
nand U22763 (N_22763,N_22340,N_22052);
and U22764 (N_22764,N_22424,N_22264);
and U22765 (N_22765,N_22027,N_22340);
nor U22766 (N_22766,N_22487,N_22290);
or U22767 (N_22767,N_22269,N_22054);
nor U22768 (N_22768,N_22104,N_22094);
and U22769 (N_22769,N_22306,N_22364);
nor U22770 (N_22770,N_22306,N_22318);
and U22771 (N_22771,N_22161,N_22058);
or U22772 (N_22772,N_22077,N_22413);
nand U22773 (N_22773,N_22333,N_22456);
or U22774 (N_22774,N_22483,N_22438);
or U22775 (N_22775,N_22041,N_22130);
nor U22776 (N_22776,N_22298,N_22051);
or U22777 (N_22777,N_22057,N_22177);
and U22778 (N_22778,N_22168,N_22485);
nor U22779 (N_22779,N_22011,N_22153);
nor U22780 (N_22780,N_22484,N_22404);
nor U22781 (N_22781,N_22029,N_22467);
and U22782 (N_22782,N_22285,N_22007);
or U22783 (N_22783,N_22374,N_22107);
nor U22784 (N_22784,N_22391,N_22493);
nand U22785 (N_22785,N_22169,N_22448);
xor U22786 (N_22786,N_22305,N_22489);
nor U22787 (N_22787,N_22235,N_22076);
and U22788 (N_22788,N_22135,N_22249);
or U22789 (N_22789,N_22028,N_22119);
nand U22790 (N_22790,N_22426,N_22038);
nor U22791 (N_22791,N_22210,N_22253);
or U22792 (N_22792,N_22356,N_22292);
and U22793 (N_22793,N_22229,N_22495);
nand U22794 (N_22794,N_22215,N_22434);
nor U22795 (N_22795,N_22079,N_22230);
nand U22796 (N_22796,N_22460,N_22194);
nand U22797 (N_22797,N_22343,N_22127);
or U22798 (N_22798,N_22479,N_22164);
nand U22799 (N_22799,N_22255,N_22109);
xnor U22800 (N_22800,N_22256,N_22183);
and U22801 (N_22801,N_22307,N_22452);
nor U22802 (N_22802,N_22117,N_22247);
nand U22803 (N_22803,N_22253,N_22082);
nand U22804 (N_22804,N_22080,N_22312);
nand U22805 (N_22805,N_22372,N_22310);
and U22806 (N_22806,N_22061,N_22270);
and U22807 (N_22807,N_22458,N_22359);
nor U22808 (N_22808,N_22158,N_22458);
and U22809 (N_22809,N_22267,N_22130);
nor U22810 (N_22810,N_22152,N_22091);
nand U22811 (N_22811,N_22127,N_22276);
or U22812 (N_22812,N_22158,N_22497);
and U22813 (N_22813,N_22321,N_22096);
and U22814 (N_22814,N_22286,N_22482);
nor U22815 (N_22815,N_22308,N_22440);
nand U22816 (N_22816,N_22286,N_22029);
and U22817 (N_22817,N_22401,N_22326);
and U22818 (N_22818,N_22177,N_22407);
or U22819 (N_22819,N_22392,N_22420);
nand U22820 (N_22820,N_22063,N_22381);
and U22821 (N_22821,N_22189,N_22282);
nand U22822 (N_22822,N_22115,N_22049);
xor U22823 (N_22823,N_22226,N_22320);
or U22824 (N_22824,N_22275,N_22137);
or U22825 (N_22825,N_22450,N_22193);
and U22826 (N_22826,N_22287,N_22432);
xnor U22827 (N_22827,N_22358,N_22307);
nor U22828 (N_22828,N_22078,N_22416);
nand U22829 (N_22829,N_22497,N_22274);
nand U22830 (N_22830,N_22128,N_22355);
or U22831 (N_22831,N_22352,N_22363);
nor U22832 (N_22832,N_22447,N_22090);
or U22833 (N_22833,N_22343,N_22346);
nand U22834 (N_22834,N_22042,N_22055);
and U22835 (N_22835,N_22432,N_22212);
and U22836 (N_22836,N_22393,N_22159);
xnor U22837 (N_22837,N_22361,N_22320);
or U22838 (N_22838,N_22290,N_22142);
nand U22839 (N_22839,N_22375,N_22399);
or U22840 (N_22840,N_22374,N_22473);
or U22841 (N_22841,N_22232,N_22095);
and U22842 (N_22842,N_22490,N_22418);
or U22843 (N_22843,N_22081,N_22302);
nor U22844 (N_22844,N_22082,N_22340);
nor U22845 (N_22845,N_22238,N_22228);
nand U22846 (N_22846,N_22398,N_22228);
and U22847 (N_22847,N_22106,N_22032);
nor U22848 (N_22848,N_22045,N_22353);
nor U22849 (N_22849,N_22178,N_22100);
or U22850 (N_22850,N_22359,N_22202);
nor U22851 (N_22851,N_22429,N_22033);
and U22852 (N_22852,N_22150,N_22127);
or U22853 (N_22853,N_22302,N_22463);
nor U22854 (N_22854,N_22089,N_22069);
xnor U22855 (N_22855,N_22433,N_22466);
xnor U22856 (N_22856,N_22076,N_22383);
nand U22857 (N_22857,N_22381,N_22491);
nand U22858 (N_22858,N_22321,N_22022);
nor U22859 (N_22859,N_22452,N_22461);
or U22860 (N_22860,N_22420,N_22068);
nor U22861 (N_22861,N_22138,N_22176);
and U22862 (N_22862,N_22038,N_22493);
xnor U22863 (N_22863,N_22268,N_22456);
and U22864 (N_22864,N_22459,N_22046);
or U22865 (N_22865,N_22422,N_22152);
and U22866 (N_22866,N_22111,N_22231);
xor U22867 (N_22867,N_22309,N_22250);
and U22868 (N_22868,N_22282,N_22205);
nor U22869 (N_22869,N_22360,N_22218);
nand U22870 (N_22870,N_22243,N_22267);
nor U22871 (N_22871,N_22206,N_22467);
and U22872 (N_22872,N_22177,N_22319);
nor U22873 (N_22873,N_22335,N_22450);
nor U22874 (N_22874,N_22176,N_22039);
or U22875 (N_22875,N_22268,N_22329);
xor U22876 (N_22876,N_22385,N_22344);
nor U22877 (N_22877,N_22065,N_22370);
or U22878 (N_22878,N_22065,N_22071);
xor U22879 (N_22879,N_22271,N_22153);
and U22880 (N_22880,N_22220,N_22111);
or U22881 (N_22881,N_22323,N_22410);
nor U22882 (N_22882,N_22060,N_22079);
nor U22883 (N_22883,N_22426,N_22233);
nor U22884 (N_22884,N_22053,N_22454);
or U22885 (N_22885,N_22436,N_22375);
nor U22886 (N_22886,N_22239,N_22158);
nand U22887 (N_22887,N_22298,N_22074);
and U22888 (N_22888,N_22310,N_22291);
nand U22889 (N_22889,N_22122,N_22243);
xor U22890 (N_22890,N_22395,N_22085);
and U22891 (N_22891,N_22201,N_22276);
or U22892 (N_22892,N_22098,N_22391);
and U22893 (N_22893,N_22139,N_22310);
nor U22894 (N_22894,N_22409,N_22481);
xor U22895 (N_22895,N_22392,N_22057);
and U22896 (N_22896,N_22081,N_22418);
xor U22897 (N_22897,N_22303,N_22389);
xnor U22898 (N_22898,N_22354,N_22448);
nand U22899 (N_22899,N_22217,N_22413);
or U22900 (N_22900,N_22011,N_22456);
nor U22901 (N_22901,N_22367,N_22252);
or U22902 (N_22902,N_22468,N_22327);
or U22903 (N_22903,N_22077,N_22000);
or U22904 (N_22904,N_22300,N_22418);
nand U22905 (N_22905,N_22435,N_22173);
and U22906 (N_22906,N_22454,N_22216);
or U22907 (N_22907,N_22250,N_22350);
xnor U22908 (N_22908,N_22381,N_22333);
and U22909 (N_22909,N_22401,N_22201);
nand U22910 (N_22910,N_22138,N_22409);
and U22911 (N_22911,N_22238,N_22209);
nand U22912 (N_22912,N_22328,N_22285);
and U22913 (N_22913,N_22161,N_22279);
or U22914 (N_22914,N_22224,N_22378);
or U22915 (N_22915,N_22081,N_22389);
nand U22916 (N_22916,N_22299,N_22487);
nand U22917 (N_22917,N_22383,N_22191);
nand U22918 (N_22918,N_22453,N_22212);
and U22919 (N_22919,N_22196,N_22006);
or U22920 (N_22920,N_22365,N_22232);
nor U22921 (N_22921,N_22344,N_22407);
nor U22922 (N_22922,N_22287,N_22476);
nand U22923 (N_22923,N_22158,N_22475);
nor U22924 (N_22924,N_22204,N_22242);
or U22925 (N_22925,N_22036,N_22222);
and U22926 (N_22926,N_22036,N_22350);
or U22927 (N_22927,N_22217,N_22031);
and U22928 (N_22928,N_22398,N_22421);
xor U22929 (N_22929,N_22063,N_22139);
and U22930 (N_22930,N_22281,N_22321);
and U22931 (N_22931,N_22372,N_22004);
xor U22932 (N_22932,N_22198,N_22306);
or U22933 (N_22933,N_22131,N_22273);
nor U22934 (N_22934,N_22049,N_22339);
and U22935 (N_22935,N_22482,N_22425);
xnor U22936 (N_22936,N_22216,N_22452);
nor U22937 (N_22937,N_22069,N_22091);
and U22938 (N_22938,N_22008,N_22060);
nor U22939 (N_22939,N_22057,N_22488);
nor U22940 (N_22940,N_22087,N_22035);
nand U22941 (N_22941,N_22001,N_22429);
nand U22942 (N_22942,N_22049,N_22031);
nor U22943 (N_22943,N_22487,N_22008);
nand U22944 (N_22944,N_22226,N_22164);
nand U22945 (N_22945,N_22133,N_22001);
nor U22946 (N_22946,N_22103,N_22464);
xnor U22947 (N_22947,N_22273,N_22050);
nor U22948 (N_22948,N_22310,N_22087);
and U22949 (N_22949,N_22268,N_22390);
or U22950 (N_22950,N_22203,N_22441);
nor U22951 (N_22951,N_22446,N_22143);
or U22952 (N_22952,N_22137,N_22404);
nor U22953 (N_22953,N_22267,N_22385);
nor U22954 (N_22954,N_22387,N_22103);
nor U22955 (N_22955,N_22097,N_22072);
nor U22956 (N_22956,N_22218,N_22240);
nand U22957 (N_22957,N_22348,N_22251);
nor U22958 (N_22958,N_22226,N_22071);
xnor U22959 (N_22959,N_22459,N_22193);
or U22960 (N_22960,N_22323,N_22342);
xnor U22961 (N_22961,N_22237,N_22330);
nand U22962 (N_22962,N_22357,N_22085);
and U22963 (N_22963,N_22441,N_22494);
and U22964 (N_22964,N_22393,N_22373);
nor U22965 (N_22965,N_22269,N_22324);
nor U22966 (N_22966,N_22374,N_22314);
or U22967 (N_22967,N_22108,N_22243);
nor U22968 (N_22968,N_22493,N_22069);
nand U22969 (N_22969,N_22122,N_22286);
or U22970 (N_22970,N_22161,N_22280);
xnor U22971 (N_22971,N_22137,N_22053);
nand U22972 (N_22972,N_22229,N_22173);
nor U22973 (N_22973,N_22226,N_22201);
or U22974 (N_22974,N_22031,N_22317);
and U22975 (N_22975,N_22233,N_22429);
or U22976 (N_22976,N_22202,N_22076);
nor U22977 (N_22977,N_22440,N_22018);
or U22978 (N_22978,N_22322,N_22331);
nor U22979 (N_22979,N_22112,N_22266);
and U22980 (N_22980,N_22234,N_22274);
nand U22981 (N_22981,N_22453,N_22464);
nor U22982 (N_22982,N_22116,N_22107);
xnor U22983 (N_22983,N_22481,N_22469);
nand U22984 (N_22984,N_22214,N_22233);
or U22985 (N_22985,N_22097,N_22239);
nand U22986 (N_22986,N_22283,N_22251);
nand U22987 (N_22987,N_22383,N_22365);
nand U22988 (N_22988,N_22134,N_22051);
nand U22989 (N_22989,N_22492,N_22341);
or U22990 (N_22990,N_22456,N_22497);
and U22991 (N_22991,N_22194,N_22002);
and U22992 (N_22992,N_22096,N_22121);
nor U22993 (N_22993,N_22437,N_22072);
and U22994 (N_22994,N_22072,N_22393);
or U22995 (N_22995,N_22381,N_22010);
or U22996 (N_22996,N_22334,N_22323);
nor U22997 (N_22997,N_22004,N_22125);
and U22998 (N_22998,N_22268,N_22162);
xnor U22999 (N_22999,N_22389,N_22182);
or U23000 (N_23000,N_22902,N_22831);
or U23001 (N_23001,N_22683,N_22527);
xor U23002 (N_23002,N_22518,N_22936);
xor U23003 (N_23003,N_22553,N_22861);
nor U23004 (N_23004,N_22732,N_22719);
xnor U23005 (N_23005,N_22884,N_22841);
nor U23006 (N_23006,N_22923,N_22987);
and U23007 (N_23007,N_22524,N_22765);
nand U23008 (N_23008,N_22946,N_22977);
nor U23009 (N_23009,N_22857,N_22706);
nand U23010 (N_23010,N_22571,N_22692);
and U23011 (N_23011,N_22982,N_22508);
nand U23012 (N_23012,N_22979,N_22908);
xor U23013 (N_23013,N_22960,N_22651);
or U23014 (N_23014,N_22583,N_22696);
and U23015 (N_23015,N_22784,N_22818);
nor U23016 (N_23016,N_22921,N_22968);
nor U23017 (N_23017,N_22686,N_22890);
xor U23018 (N_23018,N_22638,N_22903);
nand U23019 (N_23019,N_22578,N_22992);
or U23020 (N_23020,N_22876,N_22544);
and U23021 (N_23021,N_22875,N_22601);
and U23022 (N_23022,N_22862,N_22560);
or U23023 (N_23023,N_22939,N_22617);
or U23024 (N_23024,N_22853,N_22926);
or U23025 (N_23025,N_22927,N_22859);
or U23026 (N_23026,N_22754,N_22776);
nand U23027 (N_23027,N_22827,N_22756);
nand U23028 (N_23028,N_22858,N_22600);
nand U23029 (N_23029,N_22625,N_22516);
and U23030 (N_23030,N_22856,N_22632);
nand U23031 (N_23031,N_22872,N_22805);
nor U23032 (N_23032,N_22990,N_22920);
and U23033 (N_23033,N_22773,N_22832);
xor U23034 (N_23034,N_22997,N_22514);
nand U23035 (N_23035,N_22536,N_22916);
or U23036 (N_23036,N_22891,N_22561);
and U23037 (N_23037,N_22947,N_22557);
or U23038 (N_23038,N_22948,N_22956);
nand U23039 (N_23039,N_22627,N_22656);
nand U23040 (N_23040,N_22628,N_22624);
nor U23041 (N_23041,N_22547,N_22563);
nand U23042 (N_23042,N_22526,N_22883);
nor U23043 (N_23043,N_22575,N_22576);
nor U23044 (N_23044,N_22952,N_22605);
nor U23045 (N_23045,N_22910,N_22593);
nand U23046 (N_23046,N_22584,N_22922);
nor U23047 (N_23047,N_22637,N_22500);
and U23048 (N_23048,N_22610,N_22866);
xor U23049 (N_23049,N_22852,N_22528);
nand U23050 (N_23050,N_22869,N_22878);
xor U23051 (N_23051,N_22835,N_22771);
or U23052 (N_23052,N_22865,N_22906);
or U23053 (N_23053,N_22677,N_22725);
and U23054 (N_23054,N_22871,N_22515);
or U23055 (N_23055,N_22636,N_22961);
or U23056 (N_23056,N_22967,N_22972);
nand U23057 (N_23057,N_22510,N_22542);
or U23058 (N_23058,N_22660,N_22667);
nand U23059 (N_23059,N_22572,N_22585);
nor U23060 (N_23060,N_22810,N_22602);
or U23061 (N_23061,N_22998,N_22840);
or U23062 (N_23062,N_22808,N_22888);
and U23063 (N_23063,N_22556,N_22604);
nand U23064 (N_23064,N_22727,N_22909);
nand U23065 (N_23065,N_22930,N_22792);
nor U23066 (N_23066,N_22887,N_22652);
and U23067 (N_23067,N_22940,N_22944);
nor U23068 (N_23068,N_22503,N_22897);
or U23069 (N_23069,N_22507,N_22789);
and U23070 (N_23070,N_22779,N_22894);
nand U23071 (N_23071,N_22864,N_22901);
nor U23072 (N_23072,N_22679,N_22963);
nor U23073 (N_23073,N_22893,N_22767);
or U23074 (N_23074,N_22882,N_22676);
and U23075 (N_23075,N_22971,N_22778);
nand U23076 (N_23076,N_22713,N_22693);
and U23077 (N_23077,N_22774,N_22760);
nand U23078 (N_23078,N_22834,N_22786);
or U23079 (N_23079,N_22520,N_22567);
nand U23080 (N_23080,N_22907,N_22672);
nor U23081 (N_23081,N_22519,N_22597);
nor U23082 (N_23082,N_22759,N_22665);
and U23083 (N_23083,N_22914,N_22750);
or U23084 (N_23084,N_22958,N_22829);
nand U23085 (N_23085,N_22819,N_22543);
and U23086 (N_23086,N_22534,N_22552);
nand U23087 (N_23087,N_22880,N_22645);
nand U23088 (N_23088,N_22658,N_22714);
or U23089 (N_23089,N_22621,N_22523);
nand U23090 (N_23090,N_22733,N_22650);
nand U23091 (N_23091,N_22648,N_22549);
nor U23092 (N_23092,N_22950,N_22622);
or U23093 (N_23093,N_22794,N_22795);
or U23094 (N_23094,N_22643,N_22877);
or U23095 (N_23095,N_22607,N_22501);
or U23096 (N_23096,N_22855,N_22994);
and U23097 (N_23097,N_22615,N_22881);
nand U23098 (N_23098,N_22517,N_22766);
or U23099 (N_23099,N_22634,N_22659);
and U23100 (N_23100,N_22845,N_22502);
xor U23101 (N_23101,N_22935,N_22775);
or U23102 (N_23102,N_22580,N_22989);
nand U23103 (N_23103,N_22635,N_22879);
and U23104 (N_23104,N_22976,N_22616);
xnor U23105 (N_23105,N_22886,N_22701);
and U23106 (N_23106,N_22816,N_22745);
nor U23107 (N_23107,N_22577,N_22629);
and U23108 (N_23108,N_22980,N_22904);
and U23109 (N_23109,N_22912,N_22991);
and U23110 (N_23110,N_22741,N_22685);
and U23111 (N_23111,N_22721,N_22757);
nor U23112 (N_23112,N_22964,N_22631);
nor U23113 (N_23113,N_22589,N_22983);
nor U23114 (N_23114,N_22731,N_22783);
nand U23115 (N_23115,N_22974,N_22854);
nor U23116 (N_23116,N_22565,N_22924);
xnor U23117 (N_23117,N_22895,N_22966);
nor U23118 (N_23118,N_22545,N_22870);
xnor U23119 (N_23119,N_22953,N_22995);
nand U23120 (N_23120,N_22868,N_22823);
or U23121 (N_23121,N_22642,N_22613);
and U23122 (N_23122,N_22905,N_22814);
nand U23123 (N_23123,N_22569,N_22847);
nand U23124 (N_23124,N_22700,N_22506);
nor U23125 (N_23125,N_22850,N_22566);
nor U23126 (N_23126,N_22669,N_22751);
xnor U23127 (N_23127,N_22668,N_22848);
nor U23128 (N_23128,N_22554,N_22531);
and U23129 (N_23129,N_22781,N_22743);
nor U23130 (N_23130,N_22680,N_22704);
nand U23131 (N_23131,N_22839,N_22873);
nor U23132 (N_23132,N_22815,N_22509);
nor U23133 (N_23133,N_22644,N_22999);
xnor U23134 (N_23134,N_22772,N_22782);
and U23135 (N_23135,N_22931,N_22712);
nand U23136 (N_23136,N_22603,N_22770);
and U23137 (N_23137,N_22801,N_22803);
nor U23138 (N_23138,N_22800,N_22970);
nor U23139 (N_23139,N_22532,N_22504);
or U23140 (N_23140,N_22595,N_22955);
or U23141 (N_23141,N_22694,N_22758);
nand U23142 (N_23142,N_22699,N_22984);
nor U23143 (N_23143,N_22978,N_22646);
nor U23144 (N_23144,N_22730,N_22568);
xnor U23145 (N_23145,N_22806,N_22729);
and U23146 (N_23146,N_22797,N_22740);
nand U23147 (N_23147,N_22540,N_22962);
xor U23148 (N_23148,N_22618,N_22537);
nor U23149 (N_23149,N_22551,N_22695);
or U23150 (N_23150,N_22647,N_22809);
nor U23151 (N_23151,N_22562,N_22820);
nand U23152 (N_23152,N_22763,N_22802);
or U23153 (N_23153,N_22737,N_22548);
nand U23154 (N_23154,N_22985,N_22720);
nor U23155 (N_23155,N_22860,N_22594);
or U23156 (N_23156,N_22599,N_22933);
and U23157 (N_23157,N_22851,N_22538);
nor U23158 (N_23158,N_22726,N_22619);
and U23159 (N_23159,N_22911,N_22555);
or U23160 (N_23160,N_22673,N_22591);
nand U23161 (N_23161,N_22777,N_22702);
nand U23162 (N_23162,N_22559,N_22722);
nor U23163 (N_23163,N_22917,N_22609);
and U23164 (N_23164,N_22521,N_22678);
nor U23165 (N_23165,N_22639,N_22812);
nand U23166 (N_23166,N_22535,N_22975);
and U23167 (N_23167,N_22804,N_22919);
nand U23168 (N_23168,N_22747,N_22993);
nand U23169 (N_23169,N_22570,N_22541);
nor U23170 (N_23170,N_22614,N_22937);
nand U23171 (N_23171,N_22611,N_22630);
or U23172 (N_23172,N_22697,N_22546);
nand U23173 (N_23173,N_22718,N_22558);
and U23174 (N_23174,N_22657,N_22959);
or U23175 (N_23175,N_22791,N_22842);
nor U23176 (N_23176,N_22550,N_22620);
xnor U23177 (N_23177,N_22705,N_22682);
nand U23178 (N_23178,N_22768,N_22899);
or U23179 (N_23179,N_22986,N_22711);
or U23180 (N_23180,N_22653,N_22954);
or U23181 (N_23181,N_22739,N_22799);
xor U23182 (N_23182,N_22674,N_22579);
xor U23183 (N_23183,N_22666,N_22932);
or U23184 (N_23184,N_22675,N_22530);
xor U23185 (N_23185,N_22654,N_22996);
and U23186 (N_23186,N_22564,N_22641);
xnor U23187 (N_23187,N_22670,N_22588);
nand U23188 (N_23188,N_22736,N_22762);
or U23189 (N_23189,N_22663,N_22981);
and U23190 (N_23190,N_22788,N_22826);
or U23191 (N_23191,N_22709,N_22780);
nor U23192 (N_23192,N_22690,N_22885);
or U23193 (N_23193,N_22691,N_22587);
nand U23194 (N_23194,N_22681,N_22836);
nor U23195 (N_23195,N_22539,N_22574);
nor U23196 (N_23196,N_22942,N_22825);
xor U23197 (N_23197,N_22837,N_22746);
or U23198 (N_23198,N_22761,N_22707);
nand U23199 (N_23199,N_22807,N_22626);
or U23200 (N_23200,N_22592,N_22703);
nand U23201 (N_23201,N_22671,N_22723);
or U23202 (N_23202,N_22817,N_22969);
xnor U23203 (N_23203,N_22661,N_22649);
or U23204 (N_23204,N_22846,N_22957);
nor U23205 (N_23205,N_22892,N_22742);
nand U23206 (N_23206,N_22748,N_22715);
nor U23207 (N_23207,N_22687,N_22724);
and U23208 (N_23208,N_22824,N_22934);
nor U23209 (N_23209,N_22590,N_22900);
and U23210 (N_23210,N_22623,N_22633);
nand U23211 (N_23211,N_22787,N_22813);
nor U23212 (N_23212,N_22811,N_22965);
and U23213 (N_23213,N_22929,N_22655);
nand U23214 (N_23214,N_22928,N_22698);
nand U23215 (N_23215,N_22752,N_22941);
xor U23216 (N_23216,N_22843,N_22988);
nand U23217 (N_23217,N_22581,N_22913);
nand U23218 (N_23218,N_22684,N_22790);
or U23219 (N_23219,N_22598,N_22525);
and U23220 (N_23220,N_22925,N_22949);
and U23221 (N_23221,N_22744,N_22533);
nor U23222 (N_23222,N_22938,N_22793);
or U23223 (N_23223,N_22664,N_22716);
and U23224 (N_23224,N_22688,N_22821);
nor U23225 (N_23225,N_22874,N_22662);
or U23226 (N_23226,N_22708,N_22945);
nor U23227 (N_23227,N_22728,N_22596);
xor U23228 (N_23228,N_22735,N_22973);
nand U23229 (N_23229,N_22951,N_22943);
nand U23230 (N_23230,N_22513,N_22918);
and U23231 (N_23231,N_22796,N_22867);
and U23232 (N_23232,N_22898,N_22512);
nand U23233 (N_23233,N_22511,N_22505);
nor U23234 (N_23234,N_22640,N_22764);
or U23235 (N_23235,N_22833,N_22798);
and U23236 (N_23236,N_22529,N_22889);
and U23237 (N_23237,N_22896,N_22753);
nor U23238 (N_23238,N_22915,N_22769);
nand U23239 (N_23239,N_22573,N_22734);
or U23240 (N_23240,N_22755,N_22822);
or U23241 (N_23241,N_22586,N_22710);
or U23242 (N_23242,N_22522,N_22863);
nor U23243 (N_23243,N_22717,N_22738);
xnor U23244 (N_23244,N_22689,N_22844);
xor U23245 (N_23245,N_22830,N_22582);
nand U23246 (N_23246,N_22749,N_22838);
or U23247 (N_23247,N_22608,N_22849);
nor U23248 (N_23248,N_22828,N_22785);
nor U23249 (N_23249,N_22606,N_22612);
nand U23250 (N_23250,N_22891,N_22893);
or U23251 (N_23251,N_22721,N_22695);
nor U23252 (N_23252,N_22576,N_22925);
nor U23253 (N_23253,N_22584,N_22820);
nor U23254 (N_23254,N_22649,N_22658);
or U23255 (N_23255,N_22704,N_22614);
or U23256 (N_23256,N_22740,N_22841);
or U23257 (N_23257,N_22563,N_22501);
or U23258 (N_23258,N_22808,N_22671);
nand U23259 (N_23259,N_22530,N_22846);
nor U23260 (N_23260,N_22866,N_22512);
and U23261 (N_23261,N_22940,N_22823);
and U23262 (N_23262,N_22714,N_22690);
nand U23263 (N_23263,N_22998,N_22987);
or U23264 (N_23264,N_22842,N_22599);
or U23265 (N_23265,N_22746,N_22502);
xnor U23266 (N_23266,N_22822,N_22628);
xnor U23267 (N_23267,N_22713,N_22799);
nor U23268 (N_23268,N_22642,N_22789);
nor U23269 (N_23269,N_22600,N_22706);
nor U23270 (N_23270,N_22635,N_22927);
or U23271 (N_23271,N_22947,N_22578);
and U23272 (N_23272,N_22869,N_22573);
nand U23273 (N_23273,N_22641,N_22573);
xor U23274 (N_23274,N_22610,N_22592);
and U23275 (N_23275,N_22692,N_22708);
and U23276 (N_23276,N_22717,N_22735);
nor U23277 (N_23277,N_22849,N_22931);
xnor U23278 (N_23278,N_22849,N_22541);
or U23279 (N_23279,N_22903,N_22720);
and U23280 (N_23280,N_22958,N_22844);
nand U23281 (N_23281,N_22716,N_22821);
xnor U23282 (N_23282,N_22656,N_22560);
nand U23283 (N_23283,N_22895,N_22646);
or U23284 (N_23284,N_22717,N_22992);
nand U23285 (N_23285,N_22799,N_22654);
nor U23286 (N_23286,N_22830,N_22838);
or U23287 (N_23287,N_22504,N_22729);
nor U23288 (N_23288,N_22692,N_22983);
and U23289 (N_23289,N_22515,N_22556);
or U23290 (N_23290,N_22594,N_22794);
nor U23291 (N_23291,N_22940,N_22899);
or U23292 (N_23292,N_22957,N_22525);
nor U23293 (N_23293,N_22571,N_22658);
nand U23294 (N_23294,N_22590,N_22501);
nor U23295 (N_23295,N_22534,N_22820);
and U23296 (N_23296,N_22994,N_22630);
or U23297 (N_23297,N_22505,N_22690);
nor U23298 (N_23298,N_22691,N_22544);
nand U23299 (N_23299,N_22964,N_22881);
xor U23300 (N_23300,N_22891,N_22731);
xor U23301 (N_23301,N_22684,N_22709);
nand U23302 (N_23302,N_22634,N_22503);
xor U23303 (N_23303,N_22724,N_22852);
and U23304 (N_23304,N_22548,N_22684);
nor U23305 (N_23305,N_22505,N_22734);
xnor U23306 (N_23306,N_22714,N_22754);
nor U23307 (N_23307,N_22515,N_22943);
nand U23308 (N_23308,N_22573,N_22914);
nor U23309 (N_23309,N_22977,N_22927);
or U23310 (N_23310,N_22673,N_22864);
nor U23311 (N_23311,N_22852,N_22960);
and U23312 (N_23312,N_22537,N_22990);
and U23313 (N_23313,N_22839,N_22713);
xnor U23314 (N_23314,N_22707,N_22615);
and U23315 (N_23315,N_22604,N_22500);
or U23316 (N_23316,N_22627,N_22698);
nor U23317 (N_23317,N_22601,N_22600);
xor U23318 (N_23318,N_22984,N_22530);
nor U23319 (N_23319,N_22536,N_22848);
or U23320 (N_23320,N_22786,N_22661);
nor U23321 (N_23321,N_22735,N_22913);
or U23322 (N_23322,N_22791,N_22709);
nand U23323 (N_23323,N_22998,N_22675);
nor U23324 (N_23324,N_22677,N_22817);
and U23325 (N_23325,N_22959,N_22849);
and U23326 (N_23326,N_22664,N_22673);
and U23327 (N_23327,N_22508,N_22952);
and U23328 (N_23328,N_22614,N_22583);
or U23329 (N_23329,N_22991,N_22977);
nor U23330 (N_23330,N_22909,N_22830);
xor U23331 (N_23331,N_22510,N_22821);
or U23332 (N_23332,N_22810,N_22980);
and U23333 (N_23333,N_22598,N_22607);
and U23334 (N_23334,N_22806,N_22984);
xor U23335 (N_23335,N_22960,N_22630);
and U23336 (N_23336,N_22937,N_22779);
or U23337 (N_23337,N_22706,N_22895);
and U23338 (N_23338,N_22709,N_22739);
nand U23339 (N_23339,N_22800,N_22807);
and U23340 (N_23340,N_22839,N_22690);
or U23341 (N_23341,N_22837,N_22510);
and U23342 (N_23342,N_22563,N_22711);
nand U23343 (N_23343,N_22917,N_22582);
or U23344 (N_23344,N_22835,N_22954);
or U23345 (N_23345,N_22896,N_22568);
nor U23346 (N_23346,N_22992,N_22562);
nand U23347 (N_23347,N_22627,N_22900);
and U23348 (N_23348,N_22547,N_22824);
or U23349 (N_23349,N_22749,N_22846);
and U23350 (N_23350,N_22747,N_22739);
xnor U23351 (N_23351,N_22741,N_22983);
and U23352 (N_23352,N_22938,N_22545);
xnor U23353 (N_23353,N_22849,N_22853);
or U23354 (N_23354,N_22798,N_22506);
xnor U23355 (N_23355,N_22757,N_22619);
or U23356 (N_23356,N_22729,N_22687);
xor U23357 (N_23357,N_22821,N_22864);
nand U23358 (N_23358,N_22520,N_22732);
xor U23359 (N_23359,N_22738,N_22805);
or U23360 (N_23360,N_22573,N_22782);
or U23361 (N_23361,N_22845,N_22909);
or U23362 (N_23362,N_22550,N_22626);
and U23363 (N_23363,N_22517,N_22852);
nand U23364 (N_23364,N_22978,N_22757);
nand U23365 (N_23365,N_22746,N_22960);
or U23366 (N_23366,N_22592,N_22511);
and U23367 (N_23367,N_22703,N_22781);
and U23368 (N_23368,N_22853,N_22977);
or U23369 (N_23369,N_22666,N_22700);
and U23370 (N_23370,N_22906,N_22607);
or U23371 (N_23371,N_22578,N_22554);
or U23372 (N_23372,N_22776,N_22640);
and U23373 (N_23373,N_22924,N_22610);
nand U23374 (N_23374,N_22907,N_22693);
nand U23375 (N_23375,N_22547,N_22837);
nor U23376 (N_23376,N_22906,N_22718);
nor U23377 (N_23377,N_22941,N_22827);
nand U23378 (N_23378,N_22621,N_22783);
nor U23379 (N_23379,N_22638,N_22648);
or U23380 (N_23380,N_22569,N_22778);
nand U23381 (N_23381,N_22795,N_22884);
xor U23382 (N_23382,N_22853,N_22685);
xnor U23383 (N_23383,N_22725,N_22622);
and U23384 (N_23384,N_22529,N_22605);
or U23385 (N_23385,N_22638,N_22883);
nor U23386 (N_23386,N_22705,N_22511);
nor U23387 (N_23387,N_22703,N_22706);
xnor U23388 (N_23388,N_22864,N_22623);
nor U23389 (N_23389,N_22635,N_22810);
xor U23390 (N_23390,N_22890,N_22567);
nand U23391 (N_23391,N_22925,N_22907);
xor U23392 (N_23392,N_22844,N_22858);
nand U23393 (N_23393,N_22869,N_22635);
nand U23394 (N_23394,N_22711,N_22543);
or U23395 (N_23395,N_22903,N_22640);
or U23396 (N_23396,N_22691,N_22743);
nand U23397 (N_23397,N_22826,N_22985);
and U23398 (N_23398,N_22797,N_22976);
nor U23399 (N_23399,N_22924,N_22928);
nand U23400 (N_23400,N_22754,N_22913);
nand U23401 (N_23401,N_22640,N_22675);
nand U23402 (N_23402,N_22597,N_22671);
or U23403 (N_23403,N_22929,N_22909);
and U23404 (N_23404,N_22899,N_22978);
nor U23405 (N_23405,N_22684,N_22504);
nor U23406 (N_23406,N_22612,N_22681);
nor U23407 (N_23407,N_22773,N_22821);
or U23408 (N_23408,N_22730,N_22539);
nor U23409 (N_23409,N_22998,N_22777);
and U23410 (N_23410,N_22825,N_22563);
nor U23411 (N_23411,N_22995,N_22842);
nand U23412 (N_23412,N_22559,N_22542);
nand U23413 (N_23413,N_22684,N_22848);
nor U23414 (N_23414,N_22851,N_22688);
xor U23415 (N_23415,N_22738,N_22842);
nor U23416 (N_23416,N_22629,N_22678);
or U23417 (N_23417,N_22616,N_22825);
xor U23418 (N_23418,N_22504,N_22549);
xnor U23419 (N_23419,N_22691,N_22857);
nor U23420 (N_23420,N_22907,N_22698);
nor U23421 (N_23421,N_22881,N_22834);
xor U23422 (N_23422,N_22533,N_22683);
nor U23423 (N_23423,N_22942,N_22743);
xor U23424 (N_23424,N_22998,N_22905);
nand U23425 (N_23425,N_22536,N_22907);
nor U23426 (N_23426,N_22719,N_22760);
or U23427 (N_23427,N_22870,N_22759);
xor U23428 (N_23428,N_22935,N_22789);
nor U23429 (N_23429,N_22997,N_22866);
and U23430 (N_23430,N_22775,N_22602);
or U23431 (N_23431,N_22974,N_22920);
nor U23432 (N_23432,N_22969,N_22624);
xor U23433 (N_23433,N_22911,N_22580);
or U23434 (N_23434,N_22602,N_22905);
nand U23435 (N_23435,N_22878,N_22689);
and U23436 (N_23436,N_22604,N_22953);
nor U23437 (N_23437,N_22874,N_22872);
and U23438 (N_23438,N_22736,N_22666);
or U23439 (N_23439,N_22512,N_22711);
nor U23440 (N_23440,N_22723,N_22945);
xor U23441 (N_23441,N_22988,N_22570);
and U23442 (N_23442,N_22940,N_22837);
nor U23443 (N_23443,N_22730,N_22995);
nand U23444 (N_23444,N_22639,N_22999);
and U23445 (N_23445,N_22808,N_22805);
nor U23446 (N_23446,N_22773,N_22914);
and U23447 (N_23447,N_22738,N_22729);
nand U23448 (N_23448,N_22720,N_22939);
nand U23449 (N_23449,N_22708,N_22621);
nand U23450 (N_23450,N_22988,N_22743);
and U23451 (N_23451,N_22859,N_22924);
nor U23452 (N_23452,N_22616,N_22687);
or U23453 (N_23453,N_22552,N_22956);
or U23454 (N_23454,N_22666,N_22676);
or U23455 (N_23455,N_22572,N_22724);
and U23456 (N_23456,N_22627,N_22598);
xor U23457 (N_23457,N_22628,N_22540);
or U23458 (N_23458,N_22983,N_22674);
nand U23459 (N_23459,N_22741,N_22818);
xor U23460 (N_23460,N_22871,N_22834);
and U23461 (N_23461,N_22609,N_22611);
or U23462 (N_23462,N_22771,N_22747);
nor U23463 (N_23463,N_22521,N_22655);
nand U23464 (N_23464,N_22726,N_22575);
nand U23465 (N_23465,N_22525,N_22828);
xor U23466 (N_23466,N_22513,N_22566);
xor U23467 (N_23467,N_22785,N_22617);
nor U23468 (N_23468,N_22786,N_22690);
xnor U23469 (N_23469,N_22930,N_22812);
nor U23470 (N_23470,N_22981,N_22723);
and U23471 (N_23471,N_22801,N_22710);
or U23472 (N_23472,N_22958,N_22526);
nor U23473 (N_23473,N_22619,N_22522);
nor U23474 (N_23474,N_22582,N_22800);
nor U23475 (N_23475,N_22705,N_22548);
nor U23476 (N_23476,N_22549,N_22743);
or U23477 (N_23477,N_22983,N_22646);
or U23478 (N_23478,N_22564,N_22646);
xor U23479 (N_23479,N_22792,N_22925);
and U23480 (N_23480,N_22673,N_22596);
nand U23481 (N_23481,N_22678,N_22941);
and U23482 (N_23482,N_22677,N_22607);
xor U23483 (N_23483,N_22782,N_22692);
nor U23484 (N_23484,N_22855,N_22953);
nand U23485 (N_23485,N_22605,N_22791);
or U23486 (N_23486,N_22615,N_22912);
nand U23487 (N_23487,N_22703,N_22894);
nor U23488 (N_23488,N_22893,N_22688);
nand U23489 (N_23489,N_22935,N_22633);
and U23490 (N_23490,N_22714,N_22783);
nor U23491 (N_23491,N_22830,N_22894);
or U23492 (N_23492,N_22585,N_22653);
or U23493 (N_23493,N_22738,N_22747);
and U23494 (N_23494,N_22922,N_22961);
nand U23495 (N_23495,N_22775,N_22870);
and U23496 (N_23496,N_22621,N_22908);
xnor U23497 (N_23497,N_22911,N_22998);
and U23498 (N_23498,N_22891,N_22645);
and U23499 (N_23499,N_22520,N_22914);
nand U23500 (N_23500,N_23204,N_23356);
xor U23501 (N_23501,N_23022,N_23064);
nand U23502 (N_23502,N_23327,N_23072);
nand U23503 (N_23503,N_23348,N_23266);
nor U23504 (N_23504,N_23218,N_23077);
nor U23505 (N_23505,N_23366,N_23316);
or U23506 (N_23506,N_23450,N_23180);
and U23507 (N_23507,N_23147,N_23340);
xnor U23508 (N_23508,N_23142,N_23200);
or U23509 (N_23509,N_23361,N_23258);
or U23510 (N_23510,N_23215,N_23250);
xor U23511 (N_23511,N_23487,N_23192);
and U23512 (N_23512,N_23078,N_23093);
and U23513 (N_23513,N_23449,N_23489);
nand U23514 (N_23514,N_23186,N_23482);
nand U23515 (N_23515,N_23293,N_23086);
xor U23516 (N_23516,N_23320,N_23211);
xor U23517 (N_23517,N_23338,N_23411);
nand U23518 (N_23518,N_23272,N_23029);
nand U23519 (N_23519,N_23013,N_23396);
nand U23520 (N_23520,N_23279,N_23058);
or U23521 (N_23521,N_23244,N_23498);
and U23522 (N_23522,N_23416,N_23301);
nand U23523 (N_23523,N_23299,N_23317);
or U23524 (N_23524,N_23453,N_23383);
xnor U23525 (N_23525,N_23443,N_23148);
and U23526 (N_23526,N_23295,N_23201);
nor U23527 (N_23527,N_23367,N_23420);
and U23528 (N_23528,N_23474,N_23097);
nand U23529 (N_23529,N_23100,N_23444);
or U23530 (N_23530,N_23079,N_23149);
xnor U23531 (N_23531,N_23214,N_23393);
nor U23532 (N_23532,N_23116,N_23398);
nor U23533 (N_23533,N_23263,N_23304);
nor U23534 (N_23534,N_23339,N_23095);
nor U23535 (N_23535,N_23016,N_23350);
nor U23536 (N_23536,N_23158,N_23036);
nand U23537 (N_23537,N_23395,N_23045);
nand U23538 (N_23538,N_23175,N_23108);
nor U23539 (N_23539,N_23207,N_23143);
nand U23540 (N_23540,N_23169,N_23236);
nand U23541 (N_23541,N_23289,N_23405);
or U23542 (N_23542,N_23471,N_23132);
xnor U23543 (N_23543,N_23242,N_23349);
xor U23544 (N_23544,N_23378,N_23027);
nand U23545 (N_23545,N_23082,N_23328);
nor U23546 (N_23546,N_23032,N_23018);
or U23547 (N_23547,N_23052,N_23206);
or U23548 (N_23548,N_23038,N_23425);
and U23549 (N_23549,N_23371,N_23085);
and U23550 (N_23550,N_23033,N_23160);
nor U23551 (N_23551,N_23240,N_23056);
nor U23552 (N_23552,N_23111,N_23238);
xor U23553 (N_23553,N_23434,N_23145);
or U23554 (N_23554,N_23172,N_23006);
xnor U23555 (N_23555,N_23456,N_23101);
and U23556 (N_23556,N_23277,N_23230);
and U23557 (N_23557,N_23460,N_23426);
xnor U23558 (N_23558,N_23020,N_23390);
xnor U23559 (N_23559,N_23008,N_23167);
and U23560 (N_23560,N_23099,N_23477);
or U23561 (N_23561,N_23457,N_23401);
and U23562 (N_23562,N_23462,N_23227);
nor U23563 (N_23563,N_23245,N_23294);
or U23564 (N_23564,N_23281,N_23499);
nand U23565 (N_23565,N_23166,N_23445);
xnor U23566 (N_23566,N_23494,N_23246);
or U23567 (N_23567,N_23259,N_23465);
and U23568 (N_23568,N_23387,N_23187);
nor U23569 (N_23569,N_23296,N_23406);
nand U23570 (N_23570,N_23189,N_23280);
nand U23571 (N_23571,N_23188,N_23312);
nand U23572 (N_23572,N_23203,N_23285);
nand U23573 (N_23573,N_23331,N_23105);
or U23574 (N_23574,N_23255,N_23384);
xor U23575 (N_23575,N_23380,N_23023);
nor U23576 (N_23576,N_23377,N_23291);
or U23577 (N_23577,N_23243,N_23408);
or U23578 (N_23578,N_23019,N_23297);
and U23579 (N_23579,N_23417,N_23357);
nand U23580 (N_23580,N_23268,N_23382);
and U23581 (N_23581,N_23113,N_23171);
xnor U23582 (N_23582,N_23184,N_23432);
nand U23583 (N_23583,N_23110,N_23446);
nor U23584 (N_23584,N_23427,N_23308);
nor U23585 (N_23585,N_23421,N_23212);
nand U23586 (N_23586,N_23333,N_23119);
nor U23587 (N_23587,N_23492,N_23091);
or U23588 (N_23588,N_23430,N_23412);
and U23589 (N_23589,N_23488,N_23083);
or U23590 (N_23590,N_23144,N_23220);
or U23591 (N_23591,N_23403,N_23060);
nor U23592 (N_23592,N_23496,N_23046);
nor U23593 (N_23593,N_23274,N_23223);
and U23594 (N_23594,N_23454,N_23003);
and U23595 (N_23595,N_23153,N_23248);
nor U23596 (N_23596,N_23141,N_23239);
and U23597 (N_23597,N_23005,N_23273);
xor U23598 (N_23598,N_23358,N_23418);
xor U23599 (N_23599,N_23183,N_23365);
nor U23600 (N_23600,N_23346,N_23400);
nand U23601 (N_23601,N_23126,N_23014);
or U23602 (N_23602,N_23190,N_23252);
nor U23603 (N_23603,N_23138,N_23044);
and U23604 (N_23604,N_23040,N_23355);
xnor U23605 (N_23605,N_23264,N_23440);
and U23606 (N_23606,N_23286,N_23422);
nor U23607 (N_23607,N_23102,N_23399);
nand U23608 (N_23608,N_23392,N_23485);
xnor U23609 (N_23609,N_23123,N_23219);
and U23610 (N_23610,N_23115,N_23322);
and U23611 (N_23611,N_23088,N_23224);
nand U23612 (N_23612,N_23424,N_23053);
nand U23613 (N_23613,N_23466,N_23484);
nor U23614 (N_23614,N_23007,N_23354);
nor U23615 (N_23615,N_23276,N_23069);
and U23616 (N_23616,N_23490,N_23155);
and U23617 (N_23617,N_23455,N_23042);
or U23618 (N_23618,N_23235,N_23409);
or U23619 (N_23619,N_23131,N_23084);
nand U23620 (N_23620,N_23257,N_23024);
nor U23621 (N_23621,N_23195,N_23210);
nand U23622 (N_23622,N_23130,N_23065);
xor U23623 (N_23623,N_23330,N_23323);
and U23624 (N_23624,N_23278,N_23269);
and U23625 (N_23625,N_23359,N_23347);
or U23626 (N_23626,N_23117,N_23306);
and U23627 (N_23627,N_23179,N_23163);
nor U23628 (N_23628,N_23198,N_23161);
nor U23629 (N_23629,N_23092,N_23114);
nand U23630 (N_23630,N_23232,N_23125);
and U23631 (N_23631,N_23067,N_23388);
nand U23632 (N_23632,N_23157,N_23178);
nor U23633 (N_23633,N_23237,N_23282);
or U23634 (N_23634,N_23270,N_23467);
nor U23635 (N_23635,N_23288,N_23152);
nand U23636 (N_23636,N_23074,N_23066);
xnor U23637 (N_23637,N_23000,N_23433);
nand U23638 (N_23638,N_23070,N_23298);
or U23639 (N_23639,N_23234,N_23021);
or U23640 (N_23640,N_23151,N_23028);
nand U23641 (N_23641,N_23461,N_23073);
xor U23642 (N_23642,N_23181,N_23463);
nand U23643 (N_23643,N_23050,N_23419);
xor U23644 (N_23644,N_23054,N_23231);
nor U23645 (N_23645,N_23493,N_23413);
and U23646 (N_23646,N_23229,N_23039);
or U23647 (N_23647,N_23197,N_23402);
or U23648 (N_23648,N_23080,N_23096);
nand U23649 (N_23649,N_23109,N_23368);
nor U23650 (N_23650,N_23314,N_23292);
or U23651 (N_23651,N_23217,N_23318);
nor U23652 (N_23652,N_23415,N_23254);
and U23653 (N_23653,N_23335,N_23055);
xnor U23654 (N_23654,N_23199,N_23407);
or U23655 (N_23655,N_23146,N_23370);
xor U23656 (N_23656,N_23122,N_23423);
and U23657 (N_23657,N_23373,N_23057);
xor U23658 (N_23658,N_23128,N_23213);
and U23659 (N_23659,N_23309,N_23043);
nor U23660 (N_23660,N_23351,N_23313);
xor U23661 (N_23661,N_23015,N_23385);
or U23662 (N_23662,N_23325,N_23154);
xnor U23663 (N_23663,N_23001,N_23394);
and U23664 (N_23664,N_23303,N_23098);
and U23665 (N_23665,N_23193,N_23174);
or U23666 (N_23666,N_23120,N_23075);
nor U23667 (N_23667,N_23369,N_23134);
nor U23668 (N_23668,N_23472,N_23094);
and U23669 (N_23669,N_23049,N_23451);
xnor U23670 (N_23670,N_23205,N_23360);
or U23671 (N_23671,N_23459,N_23479);
nand U23672 (N_23672,N_23265,N_23156);
nor U23673 (N_23673,N_23470,N_23256);
and U23674 (N_23674,N_23191,N_23300);
nand U23675 (N_23675,N_23087,N_23139);
nand U23676 (N_23676,N_23375,N_23324);
nor U23677 (N_23677,N_23150,N_23034);
nand U23678 (N_23678,N_23352,N_23004);
nor U23679 (N_23679,N_23475,N_23336);
nor U23680 (N_23680,N_23176,N_23321);
nor U23681 (N_23681,N_23374,N_23081);
or U23682 (N_23682,N_23051,N_23436);
nor U23683 (N_23683,N_23011,N_23241);
or U23684 (N_23684,N_23480,N_23302);
xor U23685 (N_23685,N_23253,N_23025);
nand U23686 (N_23686,N_23026,N_23112);
or U23687 (N_23687,N_23106,N_23090);
and U23688 (N_23688,N_23031,N_23226);
and U23689 (N_23689,N_23251,N_23124);
or U23690 (N_23690,N_23135,N_23047);
and U23691 (N_23691,N_23249,N_23159);
and U23692 (N_23692,N_23495,N_23089);
or U23693 (N_23693,N_23121,N_23464);
and U23694 (N_23694,N_23386,N_23364);
xor U23695 (N_23695,N_23486,N_23222);
nor U23696 (N_23696,N_23041,N_23397);
nor U23697 (N_23697,N_23068,N_23168);
or U23698 (N_23698,N_23376,N_23076);
or U23699 (N_23699,N_23469,N_23165);
and U23700 (N_23700,N_23202,N_23103);
xnor U23701 (N_23701,N_23315,N_23491);
and U23702 (N_23702,N_23337,N_23381);
nor U23703 (N_23703,N_23379,N_23476);
nand U23704 (N_23704,N_23129,N_23283);
nand U23705 (N_23705,N_23452,N_23136);
nor U23706 (N_23706,N_23438,N_23435);
nor U23707 (N_23707,N_23326,N_23290);
and U23708 (N_23708,N_23133,N_23061);
or U23709 (N_23709,N_23478,N_23118);
nor U23710 (N_23710,N_23391,N_23104);
or U23711 (N_23711,N_23329,N_23063);
nand U23712 (N_23712,N_23343,N_23448);
xnor U23713 (N_23713,N_23284,N_23010);
and U23714 (N_23714,N_23225,N_23196);
and U23715 (N_23715,N_23341,N_23262);
nor U23716 (N_23716,N_23404,N_23209);
and U23717 (N_23717,N_23247,N_23012);
nor U23718 (N_23718,N_23447,N_23271);
nand U23719 (N_23719,N_23307,N_23410);
or U23720 (N_23720,N_23185,N_23208);
or U23721 (N_23721,N_23137,N_23059);
or U23722 (N_23722,N_23228,N_23030);
nand U23723 (N_23723,N_23127,N_23305);
and U23724 (N_23724,N_23310,N_23334);
xnor U23725 (N_23725,N_23437,N_23353);
nor U23726 (N_23726,N_23458,N_23311);
nand U23727 (N_23727,N_23048,N_23431);
or U23728 (N_23728,N_23177,N_23332);
nor U23729 (N_23729,N_23267,N_23414);
nor U23730 (N_23730,N_23071,N_23344);
and U23731 (N_23731,N_23363,N_23233);
or U23732 (N_23732,N_23035,N_23441);
and U23733 (N_23733,N_23037,N_23372);
xnor U23734 (N_23734,N_23182,N_23389);
nor U23735 (N_23735,N_23342,N_23164);
nand U23736 (N_23736,N_23216,N_23173);
or U23737 (N_23737,N_23442,N_23428);
or U23738 (N_23738,N_23345,N_23162);
and U23739 (N_23739,N_23062,N_23260);
nor U23740 (N_23740,N_23275,N_23107);
and U23741 (N_23741,N_23439,N_23473);
nand U23742 (N_23742,N_23261,N_23009);
and U23743 (N_23743,N_23170,N_23221);
nand U23744 (N_23744,N_23468,N_23194);
and U23745 (N_23745,N_23362,N_23002);
nand U23746 (N_23746,N_23287,N_23429);
nand U23747 (N_23747,N_23319,N_23481);
or U23748 (N_23748,N_23497,N_23483);
and U23749 (N_23749,N_23140,N_23017);
and U23750 (N_23750,N_23482,N_23330);
nand U23751 (N_23751,N_23459,N_23209);
nor U23752 (N_23752,N_23432,N_23020);
nand U23753 (N_23753,N_23278,N_23258);
or U23754 (N_23754,N_23217,N_23187);
nor U23755 (N_23755,N_23260,N_23399);
or U23756 (N_23756,N_23462,N_23485);
or U23757 (N_23757,N_23218,N_23207);
and U23758 (N_23758,N_23406,N_23039);
nor U23759 (N_23759,N_23273,N_23431);
or U23760 (N_23760,N_23285,N_23268);
or U23761 (N_23761,N_23413,N_23059);
nand U23762 (N_23762,N_23326,N_23221);
xnor U23763 (N_23763,N_23045,N_23358);
and U23764 (N_23764,N_23403,N_23056);
nor U23765 (N_23765,N_23425,N_23017);
nor U23766 (N_23766,N_23059,N_23238);
nand U23767 (N_23767,N_23031,N_23437);
and U23768 (N_23768,N_23063,N_23260);
nand U23769 (N_23769,N_23289,N_23278);
or U23770 (N_23770,N_23253,N_23392);
xor U23771 (N_23771,N_23039,N_23058);
nand U23772 (N_23772,N_23262,N_23294);
or U23773 (N_23773,N_23191,N_23222);
and U23774 (N_23774,N_23413,N_23258);
nand U23775 (N_23775,N_23491,N_23192);
nand U23776 (N_23776,N_23086,N_23259);
or U23777 (N_23777,N_23011,N_23318);
and U23778 (N_23778,N_23371,N_23115);
and U23779 (N_23779,N_23200,N_23127);
or U23780 (N_23780,N_23097,N_23083);
xnor U23781 (N_23781,N_23193,N_23282);
nand U23782 (N_23782,N_23116,N_23455);
or U23783 (N_23783,N_23379,N_23138);
nor U23784 (N_23784,N_23316,N_23396);
nand U23785 (N_23785,N_23168,N_23296);
nand U23786 (N_23786,N_23320,N_23478);
and U23787 (N_23787,N_23305,N_23415);
nor U23788 (N_23788,N_23097,N_23260);
nand U23789 (N_23789,N_23311,N_23455);
or U23790 (N_23790,N_23335,N_23393);
and U23791 (N_23791,N_23461,N_23012);
nand U23792 (N_23792,N_23009,N_23401);
or U23793 (N_23793,N_23061,N_23157);
nor U23794 (N_23794,N_23234,N_23122);
nand U23795 (N_23795,N_23264,N_23176);
nor U23796 (N_23796,N_23411,N_23331);
or U23797 (N_23797,N_23015,N_23173);
or U23798 (N_23798,N_23064,N_23119);
and U23799 (N_23799,N_23194,N_23174);
nand U23800 (N_23800,N_23261,N_23148);
nand U23801 (N_23801,N_23459,N_23332);
nand U23802 (N_23802,N_23202,N_23143);
and U23803 (N_23803,N_23339,N_23160);
nor U23804 (N_23804,N_23094,N_23484);
nand U23805 (N_23805,N_23491,N_23280);
nand U23806 (N_23806,N_23042,N_23096);
and U23807 (N_23807,N_23023,N_23275);
nand U23808 (N_23808,N_23203,N_23221);
xnor U23809 (N_23809,N_23098,N_23187);
nand U23810 (N_23810,N_23426,N_23211);
or U23811 (N_23811,N_23066,N_23437);
xor U23812 (N_23812,N_23298,N_23039);
nand U23813 (N_23813,N_23452,N_23399);
xnor U23814 (N_23814,N_23394,N_23484);
nand U23815 (N_23815,N_23150,N_23494);
or U23816 (N_23816,N_23376,N_23158);
or U23817 (N_23817,N_23469,N_23286);
nor U23818 (N_23818,N_23317,N_23344);
and U23819 (N_23819,N_23065,N_23004);
or U23820 (N_23820,N_23402,N_23219);
or U23821 (N_23821,N_23206,N_23111);
nand U23822 (N_23822,N_23019,N_23040);
nand U23823 (N_23823,N_23456,N_23190);
and U23824 (N_23824,N_23372,N_23233);
or U23825 (N_23825,N_23073,N_23334);
nor U23826 (N_23826,N_23117,N_23140);
nand U23827 (N_23827,N_23393,N_23272);
nor U23828 (N_23828,N_23213,N_23246);
nor U23829 (N_23829,N_23416,N_23062);
nor U23830 (N_23830,N_23018,N_23195);
nand U23831 (N_23831,N_23202,N_23205);
nand U23832 (N_23832,N_23117,N_23137);
nor U23833 (N_23833,N_23167,N_23088);
nor U23834 (N_23834,N_23256,N_23499);
nand U23835 (N_23835,N_23262,N_23218);
xor U23836 (N_23836,N_23152,N_23230);
nand U23837 (N_23837,N_23142,N_23359);
nand U23838 (N_23838,N_23378,N_23236);
nand U23839 (N_23839,N_23437,N_23140);
nand U23840 (N_23840,N_23199,N_23323);
nand U23841 (N_23841,N_23424,N_23082);
nand U23842 (N_23842,N_23380,N_23388);
nand U23843 (N_23843,N_23195,N_23451);
or U23844 (N_23844,N_23167,N_23398);
and U23845 (N_23845,N_23020,N_23321);
xnor U23846 (N_23846,N_23165,N_23341);
nor U23847 (N_23847,N_23454,N_23402);
or U23848 (N_23848,N_23072,N_23044);
nand U23849 (N_23849,N_23250,N_23467);
nand U23850 (N_23850,N_23001,N_23383);
xor U23851 (N_23851,N_23271,N_23381);
xor U23852 (N_23852,N_23146,N_23317);
xor U23853 (N_23853,N_23294,N_23455);
nor U23854 (N_23854,N_23139,N_23472);
or U23855 (N_23855,N_23016,N_23308);
and U23856 (N_23856,N_23384,N_23241);
nand U23857 (N_23857,N_23080,N_23025);
and U23858 (N_23858,N_23200,N_23421);
and U23859 (N_23859,N_23429,N_23441);
or U23860 (N_23860,N_23133,N_23321);
and U23861 (N_23861,N_23109,N_23335);
nor U23862 (N_23862,N_23145,N_23247);
nor U23863 (N_23863,N_23000,N_23146);
or U23864 (N_23864,N_23465,N_23440);
and U23865 (N_23865,N_23376,N_23127);
or U23866 (N_23866,N_23199,N_23309);
xnor U23867 (N_23867,N_23491,N_23210);
nand U23868 (N_23868,N_23126,N_23159);
or U23869 (N_23869,N_23444,N_23014);
or U23870 (N_23870,N_23468,N_23199);
and U23871 (N_23871,N_23084,N_23386);
nor U23872 (N_23872,N_23481,N_23428);
nor U23873 (N_23873,N_23482,N_23169);
and U23874 (N_23874,N_23208,N_23216);
or U23875 (N_23875,N_23424,N_23250);
xor U23876 (N_23876,N_23080,N_23380);
nor U23877 (N_23877,N_23222,N_23446);
xor U23878 (N_23878,N_23415,N_23286);
xnor U23879 (N_23879,N_23224,N_23170);
or U23880 (N_23880,N_23450,N_23110);
nor U23881 (N_23881,N_23032,N_23384);
and U23882 (N_23882,N_23274,N_23389);
nand U23883 (N_23883,N_23041,N_23195);
nand U23884 (N_23884,N_23016,N_23428);
and U23885 (N_23885,N_23445,N_23237);
and U23886 (N_23886,N_23113,N_23108);
nand U23887 (N_23887,N_23104,N_23284);
nor U23888 (N_23888,N_23272,N_23090);
or U23889 (N_23889,N_23400,N_23032);
nor U23890 (N_23890,N_23293,N_23439);
xnor U23891 (N_23891,N_23100,N_23433);
and U23892 (N_23892,N_23312,N_23323);
nand U23893 (N_23893,N_23296,N_23393);
xnor U23894 (N_23894,N_23137,N_23315);
nand U23895 (N_23895,N_23487,N_23223);
nand U23896 (N_23896,N_23314,N_23113);
nor U23897 (N_23897,N_23211,N_23334);
and U23898 (N_23898,N_23138,N_23199);
xnor U23899 (N_23899,N_23398,N_23498);
or U23900 (N_23900,N_23150,N_23214);
nand U23901 (N_23901,N_23380,N_23387);
nor U23902 (N_23902,N_23126,N_23309);
nand U23903 (N_23903,N_23469,N_23157);
or U23904 (N_23904,N_23154,N_23390);
nor U23905 (N_23905,N_23376,N_23386);
nand U23906 (N_23906,N_23311,N_23051);
and U23907 (N_23907,N_23049,N_23294);
and U23908 (N_23908,N_23457,N_23293);
nand U23909 (N_23909,N_23125,N_23457);
or U23910 (N_23910,N_23401,N_23377);
or U23911 (N_23911,N_23361,N_23004);
or U23912 (N_23912,N_23411,N_23059);
nor U23913 (N_23913,N_23228,N_23044);
or U23914 (N_23914,N_23181,N_23067);
and U23915 (N_23915,N_23021,N_23345);
nand U23916 (N_23916,N_23172,N_23070);
and U23917 (N_23917,N_23301,N_23258);
or U23918 (N_23918,N_23148,N_23414);
nor U23919 (N_23919,N_23099,N_23446);
nand U23920 (N_23920,N_23360,N_23440);
nor U23921 (N_23921,N_23151,N_23327);
nand U23922 (N_23922,N_23140,N_23069);
and U23923 (N_23923,N_23223,N_23394);
nor U23924 (N_23924,N_23058,N_23311);
nand U23925 (N_23925,N_23453,N_23389);
or U23926 (N_23926,N_23266,N_23428);
and U23927 (N_23927,N_23176,N_23082);
or U23928 (N_23928,N_23414,N_23295);
and U23929 (N_23929,N_23057,N_23032);
nor U23930 (N_23930,N_23488,N_23421);
nor U23931 (N_23931,N_23090,N_23094);
xor U23932 (N_23932,N_23044,N_23220);
and U23933 (N_23933,N_23477,N_23486);
and U23934 (N_23934,N_23055,N_23359);
nand U23935 (N_23935,N_23377,N_23450);
nand U23936 (N_23936,N_23319,N_23075);
or U23937 (N_23937,N_23150,N_23186);
nand U23938 (N_23938,N_23209,N_23319);
nor U23939 (N_23939,N_23021,N_23463);
nand U23940 (N_23940,N_23434,N_23343);
and U23941 (N_23941,N_23351,N_23024);
or U23942 (N_23942,N_23013,N_23382);
and U23943 (N_23943,N_23477,N_23226);
nor U23944 (N_23944,N_23099,N_23494);
nand U23945 (N_23945,N_23015,N_23299);
nor U23946 (N_23946,N_23469,N_23444);
xnor U23947 (N_23947,N_23131,N_23074);
and U23948 (N_23948,N_23119,N_23372);
xnor U23949 (N_23949,N_23448,N_23222);
or U23950 (N_23950,N_23043,N_23201);
and U23951 (N_23951,N_23274,N_23147);
or U23952 (N_23952,N_23137,N_23201);
nor U23953 (N_23953,N_23159,N_23310);
nor U23954 (N_23954,N_23042,N_23118);
nand U23955 (N_23955,N_23329,N_23030);
xnor U23956 (N_23956,N_23007,N_23461);
nand U23957 (N_23957,N_23487,N_23441);
nor U23958 (N_23958,N_23182,N_23198);
nor U23959 (N_23959,N_23116,N_23088);
xor U23960 (N_23960,N_23266,N_23182);
nand U23961 (N_23961,N_23306,N_23259);
nand U23962 (N_23962,N_23322,N_23475);
nand U23963 (N_23963,N_23226,N_23032);
or U23964 (N_23964,N_23187,N_23340);
or U23965 (N_23965,N_23037,N_23296);
nand U23966 (N_23966,N_23242,N_23323);
nor U23967 (N_23967,N_23381,N_23164);
nor U23968 (N_23968,N_23420,N_23471);
and U23969 (N_23969,N_23116,N_23264);
or U23970 (N_23970,N_23386,N_23136);
xnor U23971 (N_23971,N_23330,N_23156);
nand U23972 (N_23972,N_23127,N_23106);
and U23973 (N_23973,N_23391,N_23191);
nand U23974 (N_23974,N_23162,N_23179);
xor U23975 (N_23975,N_23282,N_23311);
xor U23976 (N_23976,N_23337,N_23409);
and U23977 (N_23977,N_23365,N_23353);
nand U23978 (N_23978,N_23163,N_23308);
and U23979 (N_23979,N_23370,N_23352);
or U23980 (N_23980,N_23053,N_23428);
xor U23981 (N_23981,N_23422,N_23390);
and U23982 (N_23982,N_23479,N_23174);
nor U23983 (N_23983,N_23286,N_23169);
nand U23984 (N_23984,N_23416,N_23202);
or U23985 (N_23985,N_23164,N_23002);
and U23986 (N_23986,N_23201,N_23082);
or U23987 (N_23987,N_23214,N_23172);
and U23988 (N_23988,N_23246,N_23064);
or U23989 (N_23989,N_23266,N_23311);
xnor U23990 (N_23990,N_23074,N_23112);
nand U23991 (N_23991,N_23293,N_23461);
or U23992 (N_23992,N_23406,N_23260);
nor U23993 (N_23993,N_23498,N_23316);
nand U23994 (N_23994,N_23383,N_23075);
nand U23995 (N_23995,N_23017,N_23366);
and U23996 (N_23996,N_23111,N_23143);
and U23997 (N_23997,N_23444,N_23152);
or U23998 (N_23998,N_23166,N_23462);
nor U23999 (N_23999,N_23483,N_23419);
nor U24000 (N_24000,N_23794,N_23880);
and U24001 (N_24001,N_23565,N_23598);
or U24002 (N_24002,N_23904,N_23626);
or U24003 (N_24003,N_23676,N_23573);
and U24004 (N_24004,N_23640,N_23587);
nand U24005 (N_24005,N_23964,N_23684);
nand U24006 (N_24006,N_23705,N_23580);
xor U24007 (N_24007,N_23986,N_23527);
and U24008 (N_24008,N_23570,N_23538);
nor U24009 (N_24009,N_23581,N_23673);
nor U24010 (N_24010,N_23997,N_23928);
or U24011 (N_24011,N_23609,N_23825);
xor U24012 (N_24012,N_23808,N_23734);
nand U24013 (N_24013,N_23937,N_23903);
and U24014 (N_24014,N_23805,N_23911);
nor U24015 (N_24015,N_23681,N_23685);
and U24016 (N_24016,N_23731,N_23807);
xor U24017 (N_24017,N_23637,N_23860);
or U24018 (N_24018,N_23615,N_23641);
or U24019 (N_24019,N_23994,N_23711);
and U24020 (N_24020,N_23672,N_23765);
nand U24021 (N_24021,N_23848,N_23863);
nor U24022 (N_24022,N_23925,N_23520);
and U24023 (N_24023,N_23922,N_23920);
xor U24024 (N_24024,N_23783,N_23650);
and U24025 (N_24025,N_23844,N_23933);
nor U24026 (N_24026,N_23966,N_23504);
or U24027 (N_24027,N_23719,N_23832);
nor U24028 (N_24028,N_23514,N_23726);
and U24029 (N_24029,N_23768,N_23838);
nand U24030 (N_24030,N_23763,N_23916);
and U24031 (N_24031,N_23795,N_23568);
nand U24032 (N_24032,N_23655,N_23550);
nand U24033 (N_24033,N_23596,N_23965);
or U24034 (N_24034,N_23564,N_23842);
nor U24035 (N_24035,N_23739,N_23841);
nand U24036 (N_24036,N_23798,N_23625);
nor U24037 (N_24037,N_23762,N_23631);
xor U24038 (N_24038,N_23834,N_23542);
nand U24039 (N_24039,N_23978,N_23954);
nand U24040 (N_24040,N_23948,N_23628);
nand U24041 (N_24041,N_23981,N_23982);
nand U24042 (N_24042,N_23621,N_23942);
or U24043 (N_24043,N_23515,N_23712);
nand U24044 (N_24044,N_23718,N_23859);
nand U24045 (N_24045,N_23605,N_23559);
nand U24046 (N_24046,N_23836,N_23553);
nand U24047 (N_24047,N_23776,N_23599);
or U24048 (N_24048,N_23769,N_23635);
or U24049 (N_24049,N_23589,N_23699);
nand U24050 (N_24050,N_23503,N_23973);
nand U24051 (N_24051,N_23696,N_23691);
nor U24052 (N_24052,N_23968,N_23998);
nor U24053 (N_24053,N_23819,N_23634);
or U24054 (N_24054,N_23623,N_23584);
and U24055 (N_24055,N_23686,N_23567);
nand U24056 (N_24056,N_23680,N_23610);
nand U24057 (N_24057,N_23707,N_23622);
or U24058 (N_24058,N_23741,N_23619);
nand U24059 (N_24059,N_23850,N_23947);
xnor U24060 (N_24060,N_23992,N_23618);
nor U24061 (N_24061,N_23972,N_23921);
nand U24062 (N_24062,N_23732,N_23806);
and U24063 (N_24063,N_23714,N_23946);
nand U24064 (N_24064,N_23675,N_23989);
and U24065 (N_24065,N_23633,N_23751);
nor U24066 (N_24066,N_23821,N_23606);
nor U24067 (N_24067,N_23727,N_23613);
or U24068 (N_24068,N_23577,N_23535);
nor U24069 (N_24069,N_23582,N_23583);
nand U24070 (N_24070,N_23875,N_23758);
nor U24071 (N_24071,N_23887,N_23513);
and U24072 (N_24072,N_23638,N_23692);
xnor U24073 (N_24073,N_23840,N_23810);
or U24074 (N_24074,N_23594,N_23743);
and U24075 (N_24075,N_23730,N_23645);
and U24076 (N_24076,N_23669,N_23907);
xnor U24077 (N_24077,N_23649,N_23857);
xnor U24078 (N_24078,N_23725,N_23931);
and U24079 (N_24079,N_23752,N_23632);
nor U24080 (N_24080,N_23813,N_23918);
nand U24081 (N_24081,N_23979,N_23656);
xor U24082 (N_24082,N_23958,N_23865);
xnor U24083 (N_24083,N_23897,N_23658);
or U24084 (N_24084,N_23664,N_23800);
xnor U24085 (N_24085,N_23956,N_23824);
nand U24086 (N_24086,N_23845,N_23822);
xor U24087 (N_24087,N_23957,N_23679);
xor U24088 (N_24088,N_23502,N_23750);
and U24089 (N_24089,N_23646,N_23914);
and U24090 (N_24090,N_23539,N_23854);
or U24091 (N_24091,N_23869,N_23701);
or U24092 (N_24092,N_23930,N_23607);
or U24093 (N_24093,N_23940,N_23951);
or U24094 (N_24094,N_23505,N_23858);
and U24095 (N_24095,N_23747,N_23540);
and U24096 (N_24096,N_23851,N_23556);
and U24097 (N_24097,N_23816,N_23855);
or U24098 (N_24098,N_23700,N_23882);
and U24099 (N_24099,N_23704,N_23804);
or U24100 (N_24100,N_23737,N_23687);
or U24101 (N_24101,N_23585,N_23600);
or U24102 (N_24102,N_23608,N_23767);
and U24103 (N_24103,N_23815,N_23715);
and U24104 (N_24104,N_23661,N_23579);
nor U24105 (N_24105,N_23761,N_23666);
and U24106 (N_24106,N_23708,N_23549);
xnor U24107 (N_24107,N_23724,N_23936);
nor U24108 (N_24108,N_23566,N_23558);
or U24109 (N_24109,N_23934,N_23576);
nor U24110 (N_24110,N_23847,N_23562);
or U24111 (N_24111,N_23874,N_23908);
nand U24112 (N_24112,N_23820,N_23995);
nor U24113 (N_24113,N_23534,N_23512);
and U24114 (N_24114,N_23697,N_23766);
nand U24115 (N_24115,N_23643,N_23785);
or U24116 (N_24116,N_23745,N_23781);
and U24117 (N_24117,N_23915,N_23976);
nand U24118 (N_24118,N_23525,N_23817);
xor U24119 (N_24119,N_23663,N_23716);
and U24120 (N_24120,N_23575,N_23636);
and U24121 (N_24121,N_23709,N_23861);
nor U24122 (N_24122,N_23516,N_23560);
nand U24123 (N_24123,N_23843,N_23846);
and U24124 (N_24124,N_23668,N_23923);
and U24125 (N_24125,N_23885,N_23670);
nand U24126 (N_24126,N_23695,N_23953);
and U24127 (N_24127,N_23603,N_23864);
nand U24128 (N_24128,N_23900,N_23563);
nand U24129 (N_24129,N_23545,N_23917);
and U24130 (N_24130,N_23932,N_23710);
or U24131 (N_24131,N_23546,N_23879);
and U24132 (N_24132,N_23812,N_23993);
xor U24133 (N_24133,N_23678,N_23912);
nor U24134 (N_24134,N_23644,N_23571);
nor U24135 (N_24135,N_23604,N_23698);
nand U24136 (N_24136,N_23639,N_23617);
nor U24137 (N_24137,N_23884,N_23749);
nand U24138 (N_24138,N_23652,N_23620);
and U24139 (N_24139,N_23886,N_23780);
nand U24140 (N_24140,N_23990,N_23849);
and U24141 (N_24141,N_23764,N_23999);
nor U24142 (N_24142,N_23902,N_23839);
xor U24143 (N_24143,N_23983,N_23787);
or U24144 (N_24144,N_23757,N_23873);
and U24145 (N_24145,N_23996,N_23784);
nor U24146 (N_24146,N_23677,N_23592);
and U24147 (N_24147,N_23533,N_23630);
or U24148 (N_24148,N_23796,N_23557);
nand U24149 (N_24149,N_23510,N_23595);
nor U24150 (N_24150,N_23778,N_23755);
xnor U24151 (N_24151,N_23888,N_23597);
nor U24152 (N_24152,N_23554,N_23939);
and U24153 (N_24153,N_23541,N_23653);
nor U24154 (N_24154,N_23909,N_23627);
nor U24155 (N_24155,N_23890,N_23926);
nor U24156 (N_24156,N_23642,N_23960);
nand U24157 (N_24157,N_23789,N_23528);
xor U24158 (N_24158,N_23814,N_23975);
nor U24159 (N_24159,N_23959,N_23629);
and U24160 (N_24160,N_23831,N_23674);
xor U24161 (N_24161,N_23878,N_23742);
nor U24162 (N_24162,N_23586,N_23889);
or U24163 (N_24163,N_23665,N_23779);
and U24164 (N_24164,N_23703,N_23616);
xnor U24165 (N_24165,N_23905,N_23756);
nor U24166 (N_24166,N_23526,N_23590);
or U24167 (N_24167,N_23506,N_23835);
and U24168 (N_24168,N_23651,N_23729);
and U24169 (N_24169,N_23720,N_23984);
or U24170 (N_24170,N_23895,N_23818);
or U24171 (N_24171,N_23501,N_23561);
nand U24172 (N_24172,N_23523,N_23774);
nand U24173 (N_24173,N_23772,N_23593);
nand U24174 (N_24174,N_23662,N_23944);
nand U24175 (N_24175,N_23867,N_23702);
nor U24176 (N_24176,N_23531,N_23770);
nor U24177 (N_24177,N_23532,N_23728);
nor U24178 (N_24178,N_23508,N_23647);
xor U24179 (N_24179,N_23799,N_23688);
nand U24180 (N_24180,N_23740,N_23881);
and U24181 (N_24181,N_23574,N_23837);
xor U24182 (N_24182,N_23521,N_23736);
or U24183 (N_24183,N_23744,N_23927);
and U24184 (N_24184,N_23826,N_23547);
and U24185 (N_24185,N_23970,N_23517);
nand U24186 (N_24186,N_23987,N_23723);
or U24187 (N_24187,N_23775,N_23694);
nor U24188 (N_24188,N_23792,N_23777);
nand U24189 (N_24189,N_23913,N_23901);
and U24190 (N_24190,N_23530,N_23536);
and U24191 (N_24191,N_23782,N_23660);
or U24192 (N_24192,N_23833,N_23555);
nor U24193 (N_24193,N_23683,N_23853);
nand U24194 (N_24194,N_23519,N_23988);
nand U24195 (N_24195,N_23801,N_23738);
nand U24196 (N_24196,N_23793,N_23786);
nor U24197 (N_24197,N_23612,N_23943);
and U24198 (N_24198,N_23963,N_23689);
nor U24199 (N_24199,N_23823,N_23529);
nor U24200 (N_24200,N_23507,N_23548);
or U24201 (N_24201,N_23522,N_23569);
or U24202 (N_24202,N_23713,N_23962);
xor U24203 (N_24203,N_23754,N_23537);
xnor U24204 (N_24204,N_23511,N_23906);
and U24205 (N_24205,N_23827,N_23551);
nand U24206 (N_24206,N_23803,N_23892);
xnor U24207 (N_24207,N_23682,N_23667);
nor U24208 (N_24208,N_23924,N_23899);
nor U24209 (N_24209,N_23952,N_23955);
nor U24210 (N_24210,N_23601,N_23733);
nand U24211 (N_24211,N_23578,N_23870);
or U24212 (N_24212,N_23722,N_23748);
or U24213 (N_24213,N_23773,N_23898);
nand U24214 (N_24214,N_23830,N_23980);
nor U24215 (N_24215,N_23985,N_23721);
or U24216 (N_24216,N_23509,N_23828);
nor U24217 (N_24217,N_23929,N_23657);
nand U24218 (N_24218,N_23950,N_23788);
and U24219 (N_24219,N_23883,N_23614);
and U24220 (N_24220,N_23771,N_23910);
nand U24221 (N_24221,N_23690,N_23611);
or U24222 (N_24222,N_23524,N_23991);
nor U24223 (N_24223,N_23760,N_23971);
nand U24224 (N_24224,N_23791,N_23872);
or U24225 (N_24225,N_23938,N_23941);
and U24226 (N_24226,N_23809,N_23790);
or U24227 (N_24227,N_23717,N_23856);
nor U24228 (N_24228,N_23518,N_23735);
or U24229 (N_24229,N_23977,N_23659);
nand U24230 (N_24230,N_23797,N_23654);
nand U24231 (N_24231,N_23949,N_23693);
and U24232 (N_24232,N_23891,N_23602);
nor U24233 (N_24233,N_23871,N_23746);
nand U24234 (N_24234,N_23893,N_23935);
or U24235 (N_24235,N_23552,N_23974);
nand U24236 (N_24236,N_23591,N_23961);
or U24237 (N_24237,N_23945,N_23967);
or U24238 (N_24238,N_23919,N_23969);
and U24239 (N_24239,N_23862,N_23852);
or U24240 (N_24240,N_23544,N_23759);
or U24241 (N_24241,N_23894,N_23753);
and U24242 (N_24242,N_23706,N_23896);
nor U24243 (N_24243,N_23588,N_23802);
or U24244 (N_24244,N_23543,N_23866);
or U24245 (N_24245,N_23829,N_23572);
or U24246 (N_24246,N_23876,N_23671);
xor U24247 (N_24247,N_23811,N_23868);
or U24248 (N_24248,N_23500,N_23648);
and U24249 (N_24249,N_23624,N_23877);
nor U24250 (N_24250,N_23938,N_23804);
nand U24251 (N_24251,N_23644,N_23748);
and U24252 (N_24252,N_23701,N_23796);
or U24253 (N_24253,N_23757,N_23586);
and U24254 (N_24254,N_23707,N_23932);
nor U24255 (N_24255,N_23713,N_23756);
nor U24256 (N_24256,N_23633,N_23566);
or U24257 (N_24257,N_23810,N_23754);
nand U24258 (N_24258,N_23632,N_23534);
nand U24259 (N_24259,N_23774,N_23521);
and U24260 (N_24260,N_23768,N_23522);
xor U24261 (N_24261,N_23999,N_23656);
nor U24262 (N_24262,N_23734,N_23517);
and U24263 (N_24263,N_23576,N_23596);
nor U24264 (N_24264,N_23912,N_23763);
nor U24265 (N_24265,N_23612,N_23735);
xor U24266 (N_24266,N_23689,N_23955);
nand U24267 (N_24267,N_23605,N_23693);
nor U24268 (N_24268,N_23527,N_23802);
nand U24269 (N_24269,N_23619,N_23914);
nand U24270 (N_24270,N_23572,N_23612);
and U24271 (N_24271,N_23862,N_23984);
xor U24272 (N_24272,N_23671,N_23867);
xor U24273 (N_24273,N_23513,N_23510);
nor U24274 (N_24274,N_23536,N_23870);
or U24275 (N_24275,N_23855,N_23700);
xor U24276 (N_24276,N_23803,N_23836);
nor U24277 (N_24277,N_23943,N_23978);
nor U24278 (N_24278,N_23617,N_23921);
nand U24279 (N_24279,N_23970,N_23839);
or U24280 (N_24280,N_23777,N_23750);
and U24281 (N_24281,N_23935,N_23547);
nand U24282 (N_24282,N_23674,N_23814);
or U24283 (N_24283,N_23831,N_23590);
nand U24284 (N_24284,N_23894,N_23585);
or U24285 (N_24285,N_23682,N_23723);
nor U24286 (N_24286,N_23868,N_23623);
and U24287 (N_24287,N_23659,N_23995);
xnor U24288 (N_24288,N_23895,N_23658);
or U24289 (N_24289,N_23643,N_23683);
nand U24290 (N_24290,N_23928,N_23846);
or U24291 (N_24291,N_23865,N_23550);
nand U24292 (N_24292,N_23940,N_23771);
nor U24293 (N_24293,N_23515,N_23768);
xnor U24294 (N_24294,N_23975,N_23612);
and U24295 (N_24295,N_23978,N_23675);
xnor U24296 (N_24296,N_23683,N_23738);
and U24297 (N_24297,N_23631,N_23558);
and U24298 (N_24298,N_23518,N_23673);
nor U24299 (N_24299,N_23829,N_23730);
nand U24300 (N_24300,N_23560,N_23974);
xor U24301 (N_24301,N_23555,N_23516);
and U24302 (N_24302,N_23779,N_23815);
and U24303 (N_24303,N_23533,N_23779);
xnor U24304 (N_24304,N_23602,N_23996);
and U24305 (N_24305,N_23767,N_23867);
and U24306 (N_24306,N_23852,N_23521);
nor U24307 (N_24307,N_23829,N_23656);
nand U24308 (N_24308,N_23835,N_23843);
xnor U24309 (N_24309,N_23627,N_23931);
xnor U24310 (N_24310,N_23655,N_23854);
or U24311 (N_24311,N_23887,N_23651);
nand U24312 (N_24312,N_23944,N_23689);
nand U24313 (N_24313,N_23861,N_23983);
xnor U24314 (N_24314,N_23608,N_23515);
nand U24315 (N_24315,N_23575,N_23885);
nor U24316 (N_24316,N_23927,N_23844);
and U24317 (N_24317,N_23855,N_23697);
and U24318 (N_24318,N_23648,N_23680);
and U24319 (N_24319,N_23548,N_23534);
nor U24320 (N_24320,N_23709,N_23900);
nor U24321 (N_24321,N_23910,N_23621);
or U24322 (N_24322,N_23733,N_23609);
nor U24323 (N_24323,N_23739,N_23955);
or U24324 (N_24324,N_23707,N_23728);
nor U24325 (N_24325,N_23875,N_23935);
and U24326 (N_24326,N_23890,N_23791);
and U24327 (N_24327,N_23879,N_23810);
nand U24328 (N_24328,N_23606,N_23820);
xor U24329 (N_24329,N_23528,N_23689);
and U24330 (N_24330,N_23588,N_23884);
nor U24331 (N_24331,N_23771,N_23624);
nor U24332 (N_24332,N_23943,N_23780);
or U24333 (N_24333,N_23929,N_23964);
or U24334 (N_24334,N_23974,N_23525);
and U24335 (N_24335,N_23909,N_23969);
and U24336 (N_24336,N_23632,N_23889);
nand U24337 (N_24337,N_23850,N_23542);
or U24338 (N_24338,N_23808,N_23525);
or U24339 (N_24339,N_23800,N_23833);
nand U24340 (N_24340,N_23810,N_23707);
nand U24341 (N_24341,N_23616,N_23568);
nor U24342 (N_24342,N_23547,N_23813);
nor U24343 (N_24343,N_23711,N_23837);
and U24344 (N_24344,N_23615,N_23703);
nor U24345 (N_24345,N_23852,N_23754);
nand U24346 (N_24346,N_23973,N_23829);
and U24347 (N_24347,N_23888,N_23553);
and U24348 (N_24348,N_23870,N_23570);
and U24349 (N_24349,N_23648,N_23731);
or U24350 (N_24350,N_23711,N_23619);
and U24351 (N_24351,N_23862,N_23630);
xor U24352 (N_24352,N_23635,N_23560);
nor U24353 (N_24353,N_23925,N_23717);
xnor U24354 (N_24354,N_23761,N_23584);
or U24355 (N_24355,N_23704,N_23796);
nand U24356 (N_24356,N_23611,N_23810);
and U24357 (N_24357,N_23976,N_23974);
or U24358 (N_24358,N_23700,N_23811);
nand U24359 (N_24359,N_23767,N_23666);
nor U24360 (N_24360,N_23882,N_23765);
and U24361 (N_24361,N_23755,N_23826);
or U24362 (N_24362,N_23545,N_23763);
or U24363 (N_24363,N_23662,N_23846);
xor U24364 (N_24364,N_23856,N_23772);
or U24365 (N_24365,N_23903,N_23868);
or U24366 (N_24366,N_23825,N_23979);
and U24367 (N_24367,N_23676,N_23689);
or U24368 (N_24368,N_23934,N_23987);
or U24369 (N_24369,N_23579,N_23738);
nor U24370 (N_24370,N_23851,N_23889);
nor U24371 (N_24371,N_23632,N_23681);
or U24372 (N_24372,N_23902,N_23647);
and U24373 (N_24373,N_23696,N_23771);
nand U24374 (N_24374,N_23692,N_23596);
xor U24375 (N_24375,N_23618,N_23956);
nor U24376 (N_24376,N_23877,N_23505);
and U24377 (N_24377,N_23840,N_23622);
nor U24378 (N_24378,N_23665,N_23516);
or U24379 (N_24379,N_23686,N_23648);
nand U24380 (N_24380,N_23982,N_23524);
nor U24381 (N_24381,N_23591,N_23509);
nand U24382 (N_24382,N_23666,N_23902);
and U24383 (N_24383,N_23771,N_23659);
and U24384 (N_24384,N_23706,N_23839);
nor U24385 (N_24385,N_23730,N_23856);
or U24386 (N_24386,N_23913,N_23938);
and U24387 (N_24387,N_23821,N_23631);
or U24388 (N_24388,N_23956,N_23737);
nand U24389 (N_24389,N_23849,N_23763);
xnor U24390 (N_24390,N_23880,N_23537);
nand U24391 (N_24391,N_23875,N_23706);
xnor U24392 (N_24392,N_23836,N_23563);
or U24393 (N_24393,N_23912,N_23758);
or U24394 (N_24394,N_23813,N_23727);
or U24395 (N_24395,N_23562,N_23727);
nand U24396 (N_24396,N_23843,N_23916);
xor U24397 (N_24397,N_23908,N_23887);
and U24398 (N_24398,N_23623,N_23843);
nor U24399 (N_24399,N_23828,N_23841);
and U24400 (N_24400,N_23574,N_23874);
nor U24401 (N_24401,N_23540,N_23521);
xor U24402 (N_24402,N_23800,N_23895);
nor U24403 (N_24403,N_23812,N_23665);
or U24404 (N_24404,N_23594,N_23829);
and U24405 (N_24405,N_23550,N_23716);
and U24406 (N_24406,N_23526,N_23780);
nor U24407 (N_24407,N_23981,N_23716);
nor U24408 (N_24408,N_23986,N_23721);
or U24409 (N_24409,N_23993,N_23790);
nand U24410 (N_24410,N_23834,N_23796);
or U24411 (N_24411,N_23973,N_23997);
nand U24412 (N_24412,N_23841,N_23879);
nand U24413 (N_24413,N_23520,N_23658);
or U24414 (N_24414,N_23786,N_23816);
nor U24415 (N_24415,N_23618,N_23615);
nor U24416 (N_24416,N_23507,N_23990);
and U24417 (N_24417,N_23527,N_23841);
nand U24418 (N_24418,N_23833,N_23544);
nor U24419 (N_24419,N_23995,N_23900);
or U24420 (N_24420,N_23841,N_23516);
nand U24421 (N_24421,N_23534,N_23952);
nor U24422 (N_24422,N_23939,N_23688);
or U24423 (N_24423,N_23515,N_23756);
nor U24424 (N_24424,N_23601,N_23617);
or U24425 (N_24425,N_23606,N_23567);
and U24426 (N_24426,N_23597,N_23944);
or U24427 (N_24427,N_23880,N_23821);
xnor U24428 (N_24428,N_23825,N_23736);
or U24429 (N_24429,N_23939,N_23938);
and U24430 (N_24430,N_23676,N_23909);
nor U24431 (N_24431,N_23576,N_23594);
and U24432 (N_24432,N_23956,N_23615);
or U24433 (N_24433,N_23805,N_23973);
nor U24434 (N_24434,N_23839,N_23654);
xnor U24435 (N_24435,N_23797,N_23620);
or U24436 (N_24436,N_23588,N_23945);
and U24437 (N_24437,N_23820,N_23808);
or U24438 (N_24438,N_23998,N_23520);
and U24439 (N_24439,N_23903,N_23630);
nand U24440 (N_24440,N_23856,N_23807);
nand U24441 (N_24441,N_23542,N_23723);
nand U24442 (N_24442,N_23788,N_23585);
and U24443 (N_24443,N_23996,N_23829);
nand U24444 (N_24444,N_23594,N_23887);
nand U24445 (N_24445,N_23671,N_23652);
and U24446 (N_24446,N_23581,N_23920);
nor U24447 (N_24447,N_23810,N_23924);
nand U24448 (N_24448,N_23857,N_23896);
nand U24449 (N_24449,N_23994,N_23719);
nor U24450 (N_24450,N_23629,N_23815);
nand U24451 (N_24451,N_23715,N_23577);
or U24452 (N_24452,N_23643,N_23710);
nor U24453 (N_24453,N_23865,N_23944);
or U24454 (N_24454,N_23895,N_23856);
xnor U24455 (N_24455,N_23795,N_23818);
or U24456 (N_24456,N_23772,N_23701);
or U24457 (N_24457,N_23949,N_23695);
nand U24458 (N_24458,N_23645,N_23594);
and U24459 (N_24459,N_23733,N_23645);
or U24460 (N_24460,N_23616,N_23500);
and U24461 (N_24461,N_23535,N_23528);
xor U24462 (N_24462,N_23648,N_23936);
and U24463 (N_24463,N_23970,N_23716);
or U24464 (N_24464,N_23984,N_23500);
nand U24465 (N_24465,N_23695,N_23733);
and U24466 (N_24466,N_23908,N_23803);
or U24467 (N_24467,N_23674,N_23580);
nor U24468 (N_24468,N_23874,N_23982);
nand U24469 (N_24469,N_23918,N_23680);
and U24470 (N_24470,N_23634,N_23557);
and U24471 (N_24471,N_23862,N_23872);
nand U24472 (N_24472,N_23892,N_23752);
and U24473 (N_24473,N_23573,N_23579);
xor U24474 (N_24474,N_23739,N_23821);
nand U24475 (N_24475,N_23781,N_23914);
nand U24476 (N_24476,N_23835,N_23800);
nor U24477 (N_24477,N_23501,N_23970);
and U24478 (N_24478,N_23882,N_23670);
or U24479 (N_24479,N_23730,N_23790);
nor U24480 (N_24480,N_23887,N_23642);
xnor U24481 (N_24481,N_23571,N_23629);
xor U24482 (N_24482,N_23699,N_23790);
or U24483 (N_24483,N_23785,N_23705);
and U24484 (N_24484,N_23543,N_23798);
nor U24485 (N_24485,N_23701,N_23588);
nand U24486 (N_24486,N_23938,N_23547);
nand U24487 (N_24487,N_23682,N_23779);
and U24488 (N_24488,N_23826,N_23590);
xnor U24489 (N_24489,N_23506,N_23605);
nor U24490 (N_24490,N_23613,N_23979);
or U24491 (N_24491,N_23684,N_23976);
nand U24492 (N_24492,N_23947,N_23557);
and U24493 (N_24493,N_23610,N_23638);
nand U24494 (N_24494,N_23504,N_23726);
or U24495 (N_24495,N_23531,N_23537);
nor U24496 (N_24496,N_23589,N_23899);
and U24497 (N_24497,N_23511,N_23696);
xor U24498 (N_24498,N_23704,N_23904);
and U24499 (N_24499,N_23636,N_23689);
nand U24500 (N_24500,N_24116,N_24433);
nor U24501 (N_24501,N_24311,N_24127);
nand U24502 (N_24502,N_24218,N_24213);
and U24503 (N_24503,N_24372,N_24394);
or U24504 (N_24504,N_24148,N_24417);
and U24505 (N_24505,N_24019,N_24078);
or U24506 (N_24506,N_24304,N_24214);
and U24507 (N_24507,N_24217,N_24167);
and U24508 (N_24508,N_24442,N_24072);
nand U24509 (N_24509,N_24450,N_24077);
and U24510 (N_24510,N_24024,N_24239);
xor U24511 (N_24511,N_24081,N_24154);
nor U24512 (N_24512,N_24074,N_24174);
and U24513 (N_24513,N_24229,N_24306);
nand U24514 (N_24514,N_24481,N_24107);
nor U24515 (N_24515,N_24065,N_24408);
nor U24516 (N_24516,N_24048,N_24281);
nand U24517 (N_24517,N_24237,N_24123);
and U24518 (N_24518,N_24262,N_24470);
and U24519 (N_24519,N_24026,N_24429);
and U24520 (N_24520,N_24027,N_24216);
nand U24521 (N_24521,N_24042,N_24452);
xor U24522 (N_24522,N_24014,N_24058);
and U24523 (N_24523,N_24469,N_24140);
and U24524 (N_24524,N_24017,N_24185);
and U24525 (N_24525,N_24087,N_24161);
nand U24526 (N_24526,N_24318,N_24240);
nand U24527 (N_24527,N_24273,N_24303);
and U24528 (N_24528,N_24241,N_24360);
xnor U24529 (N_24529,N_24492,N_24326);
nand U24530 (N_24530,N_24238,N_24426);
and U24531 (N_24531,N_24449,N_24144);
and U24532 (N_24532,N_24244,N_24104);
and U24533 (N_24533,N_24235,N_24165);
xor U24534 (N_24534,N_24176,N_24317);
or U24535 (N_24535,N_24202,N_24029);
nand U24536 (N_24536,N_24220,N_24131);
or U24537 (N_24537,N_24499,N_24416);
nand U24538 (N_24538,N_24070,N_24211);
or U24539 (N_24539,N_24332,N_24483);
or U24540 (N_24540,N_24100,N_24310);
or U24541 (N_24541,N_24106,N_24249);
and U24542 (N_24542,N_24453,N_24378);
or U24543 (N_24543,N_24034,N_24390);
and U24544 (N_24544,N_24370,N_24191);
nand U24545 (N_24545,N_24298,N_24055);
nor U24546 (N_24546,N_24094,N_24091);
nor U24547 (N_24547,N_24059,N_24342);
or U24548 (N_24548,N_24462,N_24134);
xnor U24549 (N_24549,N_24115,N_24023);
or U24550 (N_24550,N_24009,N_24199);
nor U24551 (N_24551,N_24163,N_24487);
or U24552 (N_24552,N_24097,N_24195);
or U24553 (N_24553,N_24490,N_24219);
nor U24554 (N_24554,N_24261,N_24471);
and U24555 (N_24555,N_24286,N_24251);
nor U24556 (N_24556,N_24437,N_24007);
or U24557 (N_24557,N_24143,N_24410);
nor U24558 (N_24558,N_24109,N_24083);
and U24559 (N_24559,N_24121,N_24096);
nor U24560 (N_24560,N_24207,N_24400);
nand U24561 (N_24561,N_24412,N_24444);
nor U24562 (N_24562,N_24314,N_24321);
and U24563 (N_24563,N_24079,N_24435);
nor U24564 (N_24564,N_24371,N_24287);
xor U24565 (N_24565,N_24482,N_24343);
nand U24566 (N_24566,N_24114,N_24153);
nand U24567 (N_24567,N_24393,N_24118);
and U24568 (N_24568,N_24126,N_24198);
nor U24569 (N_24569,N_24020,N_24380);
or U24570 (N_24570,N_24376,N_24448);
and U24571 (N_24571,N_24132,N_24033);
nor U24572 (N_24572,N_24149,N_24264);
nand U24573 (N_24573,N_24129,N_24276);
nand U24574 (N_24574,N_24112,N_24162);
or U24575 (N_24575,N_24405,N_24139);
nor U24576 (N_24576,N_24395,N_24358);
nand U24577 (N_24577,N_24434,N_24322);
and U24578 (N_24578,N_24331,N_24349);
or U24579 (N_24579,N_24032,N_24312);
nor U24580 (N_24580,N_24184,N_24301);
nand U24581 (N_24581,N_24004,N_24436);
xnor U24582 (N_24582,N_24054,N_24397);
and U24583 (N_24583,N_24266,N_24497);
or U24584 (N_24584,N_24166,N_24117);
nand U24585 (N_24585,N_24383,N_24480);
or U24586 (N_24586,N_24049,N_24088);
nand U24587 (N_24587,N_24302,N_24151);
nand U24588 (N_24588,N_24459,N_24386);
and U24589 (N_24589,N_24284,N_24401);
and U24590 (N_24590,N_24455,N_24036);
or U24591 (N_24591,N_24082,N_24346);
or U24592 (N_24592,N_24008,N_24130);
or U24593 (N_24593,N_24186,N_24424);
nand U24594 (N_24594,N_24415,N_24341);
or U24595 (N_24595,N_24050,N_24037);
or U24596 (N_24596,N_24046,N_24413);
or U24597 (N_24597,N_24454,N_24090);
and U24598 (N_24598,N_24044,N_24085);
and U24599 (N_24599,N_24423,N_24254);
and U24600 (N_24600,N_24283,N_24291);
nand U24601 (N_24601,N_24045,N_24063);
nor U24602 (N_24602,N_24488,N_24293);
xnor U24603 (N_24603,N_24170,N_24022);
nor U24604 (N_24604,N_24141,N_24495);
xor U24605 (N_24605,N_24190,N_24086);
xor U24606 (N_24606,N_24041,N_24292);
and U24607 (N_24607,N_24060,N_24061);
or U24608 (N_24608,N_24025,N_24382);
and U24609 (N_24609,N_24498,N_24466);
and U24610 (N_24610,N_24280,N_24282);
and U24611 (N_24611,N_24122,N_24335);
and U24612 (N_24612,N_24226,N_24359);
nand U24613 (N_24613,N_24447,N_24461);
or U24614 (N_24614,N_24289,N_24067);
nor U24615 (N_24615,N_24399,N_24420);
xnor U24616 (N_24616,N_24253,N_24005);
nor U24617 (N_24617,N_24125,N_24236);
nand U24618 (N_24618,N_24002,N_24338);
or U24619 (N_24619,N_24098,N_24385);
xor U24620 (N_24620,N_24031,N_24150);
nor U24621 (N_24621,N_24197,N_24018);
nor U24622 (N_24622,N_24296,N_24245);
or U24623 (N_24623,N_24040,N_24035);
nand U24624 (N_24624,N_24446,N_24305);
or U24625 (N_24625,N_24362,N_24330);
nand U24626 (N_24626,N_24223,N_24493);
nor U24627 (N_24627,N_24428,N_24183);
or U24628 (N_24628,N_24006,N_24278);
or U24629 (N_24629,N_24193,N_24047);
and U24630 (N_24630,N_24248,N_24373);
nor U24631 (N_24631,N_24039,N_24189);
or U24632 (N_24632,N_24267,N_24344);
or U24633 (N_24633,N_24113,N_24486);
or U24634 (N_24634,N_24108,N_24368);
nor U24635 (N_24635,N_24396,N_24270);
or U24636 (N_24636,N_24379,N_24496);
and U24637 (N_24637,N_24173,N_24250);
or U24638 (N_24638,N_24354,N_24340);
and U24639 (N_24639,N_24076,N_24187);
and U24640 (N_24640,N_24111,N_24209);
nor U24641 (N_24641,N_24422,N_24208);
nand U24642 (N_24642,N_24308,N_24212);
and U24643 (N_24643,N_24353,N_24015);
and U24644 (N_24644,N_24155,N_24001);
or U24645 (N_24645,N_24464,N_24421);
nor U24646 (N_24646,N_24389,N_24328);
and U24647 (N_24647,N_24099,N_24438);
or U24648 (N_24648,N_24053,N_24327);
xnor U24649 (N_24649,N_24265,N_24407);
or U24650 (N_24650,N_24297,N_24419);
and U24651 (N_24651,N_24230,N_24105);
nor U24652 (N_24652,N_24095,N_24404);
nand U24653 (N_24653,N_24467,N_24227);
and U24654 (N_24654,N_24356,N_24384);
nor U24655 (N_24655,N_24485,N_24369);
nor U24656 (N_24656,N_24156,N_24247);
nand U24657 (N_24657,N_24246,N_24221);
or U24658 (N_24658,N_24120,N_24133);
and U24659 (N_24659,N_24479,N_24171);
xor U24660 (N_24660,N_24274,N_24336);
and U24661 (N_24661,N_24352,N_24158);
xnor U24662 (N_24662,N_24345,N_24391);
nor U24663 (N_24663,N_24175,N_24392);
nand U24664 (N_24664,N_24075,N_24196);
xor U24665 (N_24665,N_24159,N_24361);
or U24666 (N_24666,N_24204,N_24474);
or U24667 (N_24667,N_24409,N_24348);
and U24668 (N_24668,N_24146,N_24418);
nor U24669 (N_24669,N_24478,N_24071);
nand U24670 (N_24670,N_24411,N_24043);
and U24671 (N_24671,N_24398,N_24160);
nand U24672 (N_24672,N_24432,N_24279);
nand U24673 (N_24673,N_24092,N_24381);
nor U24674 (N_24674,N_24069,N_24333);
or U24675 (N_24675,N_24295,N_24124);
nor U24676 (N_24676,N_24316,N_24271);
and U24677 (N_24677,N_24307,N_24458);
nand U24678 (N_24678,N_24285,N_24259);
and U24679 (N_24679,N_24300,N_24313);
nand U24680 (N_24680,N_24030,N_24403);
nand U24681 (N_24681,N_24350,N_24288);
nor U24682 (N_24682,N_24255,N_24347);
and U24683 (N_24683,N_24365,N_24387);
xnor U24684 (N_24684,N_24089,N_24351);
or U24685 (N_24685,N_24210,N_24206);
xnor U24686 (N_24686,N_24013,N_24172);
nand U24687 (N_24687,N_24064,N_24073);
nand U24688 (N_24688,N_24177,N_24277);
nand U24689 (N_24689,N_24000,N_24275);
nor U24690 (N_24690,N_24080,N_24325);
nor U24691 (N_24691,N_24056,N_24137);
nand U24692 (N_24692,N_24425,N_24119);
or U24693 (N_24693,N_24334,N_24477);
or U24694 (N_24694,N_24068,N_24021);
and U24695 (N_24695,N_24366,N_24375);
nor U24696 (N_24696,N_24363,N_24203);
or U24697 (N_24697,N_24231,N_24324);
nor U24698 (N_24698,N_24299,N_24084);
and U24699 (N_24699,N_24252,N_24258);
and U24700 (N_24700,N_24355,N_24319);
and U24701 (N_24701,N_24272,N_24441);
and U24702 (N_24702,N_24168,N_24457);
or U24703 (N_24703,N_24456,N_24388);
nor U24704 (N_24704,N_24440,N_24491);
nand U24705 (N_24705,N_24257,N_24294);
and U24706 (N_24706,N_24135,N_24494);
nor U24707 (N_24707,N_24147,N_24337);
and U24708 (N_24708,N_24402,N_24468);
and U24709 (N_24709,N_24339,N_24263);
and U24710 (N_24710,N_24228,N_24445);
and U24711 (N_24711,N_24451,N_24243);
or U24712 (N_24712,N_24028,N_24038);
or U24713 (N_24713,N_24136,N_24169);
nor U24714 (N_24714,N_24101,N_24431);
and U24715 (N_24715,N_24182,N_24138);
or U24716 (N_24716,N_24443,N_24232);
nor U24717 (N_24717,N_24377,N_24233);
nor U24718 (N_24718,N_24011,N_24242);
nand U24719 (N_24719,N_24309,N_24142);
nor U24720 (N_24720,N_24215,N_24234);
nand U24721 (N_24721,N_24427,N_24357);
nand U24722 (N_24722,N_24051,N_24164);
nand U24723 (N_24723,N_24200,N_24016);
nor U24724 (N_24724,N_24364,N_24066);
xnor U24725 (N_24725,N_24329,N_24414);
xor U24726 (N_24726,N_24367,N_24489);
or U24727 (N_24727,N_24465,N_24260);
and U24728 (N_24728,N_24192,N_24102);
nand U24729 (N_24729,N_24003,N_24439);
and U24730 (N_24730,N_24062,N_24323);
nor U24731 (N_24731,N_24475,N_24460);
or U24732 (N_24732,N_24205,N_24110);
and U24733 (N_24733,N_24093,N_24181);
and U24734 (N_24734,N_24484,N_24472);
or U24735 (N_24735,N_24052,N_24157);
or U24736 (N_24736,N_24201,N_24406);
nand U24737 (N_24737,N_24269,N_24315);
or U24738 (N_24738,N_24476,N_24179);
or U24739 (N_24739,N_24222,N_24103);
nor U24740 (N_24740,N_24430,N_24320);
xnor U24741 (N_24741,N_24180,N_24152);
xor U24742 (N_24742,N_24145,N_24012);
nand U24743 (N_24743,N_24057,N_24010);
xnor U24744 (N_24744,N_24225,N_24268);
nor U24745 (N_24745,N_24188,N_24463);
nor U24746 (N_24746,N_24224,N_24194);
and U24747 (N_24747,N_24290,N_24473);
nor U24748 (N_24748,N_24128,N_24178);
nand U24749 (N_24749,N_24256,N_24374);
nor U24750 (N_24750,N_24133,N_24459);
and U24751 (N_24751,N_24237,N_24061);
nor U24752 (N_24752,N_24215,N_24258);
nor U24753 (N_24753,N_24466,N_24415);
xnor U24754 (N_24754,N_24421,N_24209);
and U24755 (N_24755,N_24446,N_24374);
nand U24756 (N_24756,N_24028,N_24425);
nand U24757 (N_24757,N_24005,N_24373);
nor U24758 (N_24758,N_24212,N_24271);
nor U24759 (N_24759,N_24024,N_24417);
or U24760 (N_24760,N_24480,N_24143);
and U24761 (N_24761,N_24254,N_24250);
nor U24762 (N_24762,N_24107,N_24415);
and U24763 (N_24763,N_24197,N_24066);
and U24764 (N_24764,N_24465,N_24056);
or U24765 (N_24765,N_24041,N_24220);
nor U24766 (N_24766,N_24290,N_24350);
and U24767 (N_24767,N_24492,N_24165);
nor U24768 (N_24768,N_24467,N_24184);
and U24769 (N_24769,N_24092,N_24116);
nand U24770 (N_24770,N_24217,N_24211);
nor U24771 (N_24771,N_24002,N_24029);
or U24772 (N_24772,N_24263,N_24112);
nand U24773 (N_24773,N_24326,N_24066);
and U24774 (N_24774,N_24464,N_24375);
xnor U24775 (N_24775,N_24053,N_24025);
nor U24776 (N_24776,N_24085,N_24315);
or U24777 (N_24777,N_24268,N_24474);
xor U24778 (N_24778,N_24132,N_24064);
or U24779 (N_24779,N_24062,N_24271);
or U24780 (N_24780,N_24089,N_24441);
xor U24781 (N_24781,N_24012,N_24051);
nand U24782 (N_24782,N_24283,N_24136);
nor U24783 (N_24783,N_24374,N_24323);
nor U24784 (N_24784,N_24473,N_24135);
and U24785 (N_24785,N_24215,N_24281);
and U24786 (N_24786,N_24324,N_24011);
and U24787 (N_24787,N_24331,N_24039);
nor U24788 (N_24788,N_24196,N_24087);
nand U24789 (N_24789,N_24165,N_24278);
nand U24790 (N_24790,N_24421,N_24006);
nor U24791 (N_24791,N_24087,N_24237);
nand U24792 (N_24792,N_24286,N_24194);
or U24793 (N_24793,N_24414,N_24313);
or U24794 (N_24794,N_24414,N_24444);
nand U24795 (N_24795,N_24097,N_24119);
xor U24796 (N_24796,N_24215,N_24336);
or U24797 (N_24797,N_24406,N_24266);
and U24798 (N_24798,N_24188,N_24166);
xnor U24799 (N_24799,N_24305,N_24047);
and U24800 (N_24800,N_24315,N_24176);
and U24801 (N_24801,N_24283,N_24056);
and U24802 (N_24802,N_24274,N_24162);
nor U24803 (N_24803,N_24426,N_24461);
nor U24804 (N_24804,N_24404,N_24069);
nand U24805 (N_24805,N_24409,N_24137);
nand U24806 (N_24806,N_24358,N_24136);
xnor U24807 (N_24807,N_24040,N_24309);
nand U24808 (N_24808,N_24174,N_24434);
and U24809 (N_24809,N_24315,N_24297);
or U24810 (N_24810,N_24401,N_24306);
nand U24811 (N_24811,N_24387,N_24431);
xor U24812 (N_24812,N_24364,N_24075);
nor U24813 (N_24813,N_24200,N_24191);
nand U24814 (N_24814,N_24407,N_24349);
or U24815 (N_24815,N_24053,N_24302);
nor U24816 (N_24816,N_24407,N_24454);
and U24817 (N_24817,N_24166,N_24208);
nor U24818 (N_24818,N_24470,N_24292);
or U24819 (N_24819,N_24129,N_24226);
nor U24820 (N_24820,N_24377,N_24312);
nand U24821 (N_24821,N_24389,N_24218);
nor U24822 (N_24822,N_24308,N_24277);
or U24823 (N_24823,N_24344,N_24265);
and U24824 (N_24824,N_24496,N_24054);
xnor U24825 (N_24825,N_24298,N_24147);
xnor U24826 (N_24826,N_24431,N_24003);
and U24827 (N_24827,N_24469,N_24274);
and U24828 (N_24828,N_24082,N_24313);
nor U24829 (N_24829,N_24455,N_24025);
and U24830 (N_24830,N_24385,N_24331);
nor U24831 (N_24831,N_24184,N_24432);
or U24832 (N_24832,N_24227,N_24311);
nor U24833 (N_24833,N_24317,N_24133);
nor U24834 (N_24834,N_24459,N_24337);
nand U24835 (N_24835,N_24397,N_24124);
or U24836 (N_24836,N_24077,N_24056);
or U24837 (N_24837,N_24426,N_24312);
nor U24838 (N_24838,N_24331,N_24121);
or U24839 (N_24839,N_24116,N_24094);
xor U24840 (N_24840,N_24238,N_24107);
or U24841 (N_24841,N_24273,N_24150);
or U24842 (N_24842,N_24428,N_24100);
or U24843 (N_24843,N_24123,N_24384);
or U24844 (N_24844,N_24132,N_24182);
and U24845 (N_24845,N_24242,N_24493);
nand U24846 (N_24846,N_24049,N_24073);
xor U24847 (N_24847,N_24359,N_24212);
or U24848 (N_24848,N_24401,N_24494);
nand U24849 (N_24849,N_24475,N_24352);
xor U24850 (N_24850,N_24366,N_24269);
xor U24851 (N_24851,N_24372,N_24236);
nand U24852 (N_24852,N_24499,N_24376);
or U24853 (N_24853,N_24420,N_24393);
nand U24854 (N_24854,N_24264,N_24367);
and U24855 (N_24855,N_24358,N_24226);
nand U24856 (N_24856,N_24411,N_24471);
and U24857 (N_24857,N_24199,N_24458);
nor U24858 (N_24858,N_24384,N_24378);
nand U24859 (N_24859,N_24357,N_24130);
nor U24860 (N_24860,N_24349,N_24133);
nand U24861 (N_24861,N_24478,N_24026);
and U24862 (N_24862,N_24297,N_24087);
nor U24863 (N_24863,N_24467,N_24038);
nand U24864 (N_24864,N_24198,N_24485);
nand U24865 (N_24865,N_24364,N_24344);
nand U24866 (N_24866,N_24057,N_24214);
nand U24867 (N_24867,N_24220,N_24331);
or U24868 (N_24868,N_24349,N_24084);
and U24869 (N_24869,N_24454,N_24354);
nor U24870 (N_24870,N_24039,N_24205);
or U24871 (N_24871,N_24328,N_24461);
xnor U24872 (N_24872,N_24390,N_24277);
nand U24873 (N_24873,N_24358,N_24213);
and U24874 (N_24874,N_24308,N_24184);
nor U24875 (N_24875,N_24381,N_24233);
nand U24876 (N_24876,N_24075,N_24473);
nand U24877 (N_24877,N_24280,N_24237);
nand U24878 (N_24878,N_24404,N_24378);
or U24879 (N_24879,N_24373,N_24240);
and U24880 (N_24880,N_24373,N_24356);
or U24881 (N_24881,N_24363,N_24443);
nand U24882 (N_24882,N_24155,N_24449);
nand U24883 (N_24883,N_24168,N_24076);
or U24884 (N_24884,N_24197,N_24360);
nand U24885 (N_24885,N_24388,N_24244);
and U24886 (N_24886,N_24155,N_24221);
nand U24887 (N_24887,N_24412,N_24351);
nand U24888 (N_24888,N_24381,N_24051);
and U24889 (N_24889,N_24034,N_24329);
nor U24890 (N_24890,N_24172,N_24322);
nor U24891 (N_24891,N_24363,N_24093);
and U24892 (N_24892,N_24471,N_24410);
nand U24893 (N_24893,N_24394,N_24118);
or U24894 (N_24894,N_24032,N_24197);
nand U24895 (N_24895,N_24314,N_24310);
and U24896 (N_24896,N_24039,N_24241);
xor U24897 (N_24897,N_24227,N_24364);
nand U24898 (N_24898,N_24234,N_24325);
nor U24899 (N_24899,N_24253,N_24415);
or U24900 (N_24900,N_24054,N_24099);
nand U24901 (N_24901,N_24426,N_24158);
nor U24902 (N_24902,N_24032,N_24210);
and U24903 (N_24903,N_24245,N_24286);
nor U24904 (N_24904,N_24477,N_24060);
xor U24905 (N_24905,N_24408,N_24210);
nor U24906 (N_24906,N_24399,N_24271);
nand U24907 (N_24907,N_24022,N_24189);
or U24908 (N_24908,N_24095,N_24258);
nand U24909 (N_24909,N_24062,N_24042);
or U24910 (N_24910,N_24385,N_24356);
or U24911 (N_24911,N_24148,N_24131);
nor U24912 (N_24912,N_24358,N_24069);
nand U24913 (N_24913,N_24235,N_24425);
or U24914 (N_24914,N_24317,N_24099);
nand U24915 (N_24915,N_24176,N_24422);
and U24916 (N_24916,N_24367,N_24108);
and U24917 (N_24917,N_24406,N_24207);
and U24918 (N_24918,N_24472,N_24048);
xnor U24919 (N_24919,N_24020,N_24495);
nor U24920 (N_24920,N_24174,N_24188);
or U24921 (N_24921,N_24236,N_24274);
and U24922 (N_24922,N_24394,N_24075);
or U24923 (N_24923,N_24034,N_24078);
or U24924 (N_24924,N_24278,N_24270);
or U24925 (N_24925,N_24130,N_24189);
nand U24926 (N_24926,N_24340,N_24228);
or U24927 (N_24927,N_24090,N_24276);
nand U24928 (N_24928,N_24203,N_24207);
nor U24929 (N_24929,N_24336,N_24312);
or U24930 (N_24930,N_24359,N_24335);
nor U24931 (N_24931,N_24238,N_24292);
xnor U24932 (N_24932,N_24134,N_24154);
nor U24933 (N_24933,N_24380,N_24094);
nor U24934 (N_24934,N_24265,N_24092);
or U24935 (N_24935,N_24044,N_24340);
xor U24936 (N_24936,N_24389,N_24124);
and U24937 (N_24937,N_24156,N_24258);
nand U24938 (N_24938,N_24300,N_24212);
and U24939 (N_24939,N_24144,N_24014);
or U24940 (N_24940,N_24052,N_24044);
xnor U24941 (N_24941,N_24277,N_24203);
xor U24942 (N_24942,N_24475,N_24367);
xnor U24943 (N_24943,N_24208,N_24152);
xor U24944 (N_24944,N_24220,N_24023);
nand U24945 (N_24945,N_24175,N_24195);
and U24946 (N_24946,N_24130,N_24207);
or U24947 (N_24947,N_24264,N_24423);
nor U24948 (N_24948,N_24256,N_24479);
or U24949 (N_24949,N_24011,N_24006);
nand U24950 (N_24950,N_24035,N_24140);
nand U24951 (N_24951,N_24049,N_24497);
and U24952 (N_24952,N_24466,N_24286);
or U24953 (N_24953,N_24157,N_24398);
nand U24954 (N_24954,N_24041,N_24425);
nand U24955 (N_24955,N_24121,N_24443);
nand U24956 (N_24956,N_24214,N_24493);
nand U24957 (N_24957,N_24216,N_24030);
xnor U24958 (N_24958,N_24385,N_24365);
nand U24959 (N_24959,N_24333,N_24127);
and U24960 (N_24960,N_24448,N_24330);
or U24961 (N_24961,N_24433,N_24022);
xnor U24962 (N_24962,N_24112,N_24486);
or U24963 (N_24963,N_24490,N_24408);
nor U24964 (N_24964,N_24426,N_24224);
xor U24965 (N_24965,N_24301,N_24228);
and U24966 (N_24966,N_24281,N_24339);
or U24967 (N_24967,N_24015,N_24297);
nor U24968 (N_24968,N_24280,N_24416);
or U24969 (N_24969,N_24240,N_24300);
nor U24970 (N_24970,N_24428,N_24095);
nand U24971 (N_24971,N_24094,N_24362);
or U24972 (N_24972,N_24432,N_24046);
nor U24973 (N_24973,N_24302,N_24378);
and U24974 (N_24974,N_24386,N_24251);
nand U24975 (N_24975,N_24125,N_24063);
and U24976 (N_24976,N_24446,N_24419);
nor U24977 (N_24977,N_24269,N_24426);
nand U24978 (N_24978,N_24432,N_24269);
xnor U24979 (N_24979,N_24108,N_24064);
or U24980 (N_24980,N_24404,N_24365);
or U24981 (N_24981,N_24247,N_24342);
or U24982 (N_24982,N_24364,N_24381);
nand U24983 (N_24983,N_24005,N_24068);
or U24984 (N_24984,N_24196,N_24326);
nor U24985 (N_24985,N_24197,N_24449);
nor U24986 (N_24986,N_24467,N_24453);
and U24987 (N_24987,N_24125,N_24225);
and U24988 (N_24988,N_24057,N_24213);
or U24989 (N_24989,N_24289,N_24415);
nand U24990 (N_24990,N_24245,N_24142);
nand U24991 (N_24991,N_24123,N_24161);
xnor U24992 (N_24992,N_24306,N_24347);
and U24993 (N_24993,N_24150,N_24303);
or U24994 (N_24994,N_24064,N_24139);
or U24995 (N_24995,N_24102,N_24091);
nand U24996 (N_24996,N_24456,N_24224);
or U24997 (N_24997,N_24217,N_24175);
nor U24998 (N_24998,N_24405,N_24059);
or U24999 (N_24999,N_24493,N_24098);
and UO_0 (O_0,N_24529,N_24913);
or UO_1 (O_1,N_24975,N_24520);
nand UO_2 (O_2,N_24857,N_24619);
nand UO_3 (O_3,N_24819,N_24550);
or UO_4 (O_4,N_24981,N_24729);
or UO_5 (O_5,N_24706,N_24671);
and UO_6 (O_6,N_24590,N_24504);
nor UO_7 (O_7,N_24828,N_24921);
or UO_8 (O_8,N_24612,N_24986);
and UO_9 (O_9,N_24652,N_24958);
nor UO_10 (O_10,N_24761,N_24528);
nor UO_11 (O_11,N_24995,N_24541);
xor UO_12 (O_12,N_24628,N_24740);
nand UO_13 (O_13,N_24714,N_24687);
nand UO_14 (O_14,N_24580,N_24607);
nand UO_15 (O_15,N_24843,N_24655);
and UO_16 (O_16,N_24577,N_24808);
or UO_17 (O_17,N_24930,N_24517);
nor UO_18 (O_18,N_24609,N_24928);
nand UO_19 (O_19,N_24833,N_24912);
or UO_20 (O_20,N_24683,N_24648);
nand UO_21 (O_21,N_24690,N_24601);
or UO_22 (O_22,N_24638,N_24964);
and UO_23 (O_23,N_24859,N_24746);
nand UO_24 (O_24,N_24689,N_24691);
or UO_25 (O_25,N_24610,N_24557);
and UO_26 (O_26,N_24634,N_24621);
or UO_27 (O_27,N_24873,N_24973);
nand UO_28 (O_28,N_24583,N_24954);
xor UO_29 (O_29,N_24855,N_24830);
and UO_30 (O_30,N_24844,N_24592);
nand UO_31 (O_31,N_24699,N_24821);
nand UO_32 (O_32,N_24936,N_24755);
xnor UO_33 (O_33,N_24796,N_24663);
nor UO_34 (O_34,N_24525,N_24717);
or UO_35 (O_35,N_24759,N_24965);
and UO_36 (O_36,N_24713,N_24503);
and UO_37 (O_37,N_24751,N_24733);
xnor UO_38 (O_38,N_24623,N_24994);
or UO_39 (O_39,N_24938,N_24910);
xnor UO_40 (O_40,N_24579,N_24667);
nor UO_41 (O_41,N_24640,N_24863);
nor UO_42 (O_42,N_24564,N_24510);
or UO_43 (O_43,N_24826,N_24664);
nand UO_44 (O_44,N_24716,N_24611);
nor UO_45 (O_45,N_24887,N_24603);
nor UO_46 (O_46,N_24811,N_24805);
and UO_47 (O_47,N_24825,N_24727);
or UO_48 (O_48,N_24862,N_24933);
nand UO_49 (O_49,N_24891,N_24702);
and UO_50 (O_50,N_24756,N_24556);
nor UO_51 (O_51,N_24822,N_24694);
nor UO_52 (O_52,N_24661,N_24858);
and UO_53 (O_53,N_24941,N_24851);
and UO_54 (O_54,N_24516,N_24861);
nor UO_55 (O_55,N_24688,N_24888);
nand UO_56 (O_56,N_24877,N_24831);
and UO_57 (O_57,N_24553,N_24974);
or UO_58 (O_58,N_24696,N_24884);
nor UO_59 (O_59,N_24939,N_24747);
or UO_60 (O_60,N_24565,N_24820);
or UO_61 (O_61,N_24934,N_24669);
or UO_62 (O_62,N_24952,N_24615);
nor UO_63 (O_63,N_24997,N_24660);
xnor UO_64 (O_64,N_24633,N_24723);
and UO_65 (O_65,N_24976,N_24818);
and UO_66 (O_66,N_24555,N_24650);
and UO_67 (O_67,N_24624,N_24540);
nor UO_68 (O_68,N_24585,N_24600);
and UO_69 (O_69,N_24507,N_24898);
or UO_70 (O_70,N_24876,N_24644);
nor UO_71 (O_71,N_24956,N_24736);
nor UO_72 (O_72,N_24878,N_24500);
nand UO_73 (O_73,N_24561,N_24763);
and UO_74 (O_74,N_24902,N_24719);
or UO_75 (O_75,N_24708,N_24942);
nor UO_76 (O_76,N_24718,N_24695);
nand UO_77 (O_77,N_24790,N_24591);
xor UO_78 (O_78,N_24904,N_24924);
and UO_79 (O_79,N_24743,N_24643);
and UO_80 (O_80,N_24674,N_24515);
nand UO_81 (O_81,N_24735,N_24935);
and UO_82 (O_82,N_24947,N_24840);
or UO_83 (O_83,N_24697,N_24800);
or UO_84 (O_84,N_24886,N_24931);
or UO_85 (O_85,N_24522,N_24552);
or UO_86 (O_86,N_24530,N_24745);
nor UO_87 (O_87,N_24606,N_24968);
nand UO_88 (O_88,N_24787,N_24707);
or UO_89 (O_89,N_24509,N_24998);
and UO_90 (O_90,N_24535,N_24532);
and UO_91 (O_91,N_24963,N_24685);
and UO_92 (O_92,N_24710,N_24527);
nor UO_93 (O_93,N_24883,N_24943);
nor UO_94 (O_94,N_24620,N_24693);
or UO_95 (O_95,N_24978,N_24874);
or UO_96 (O_96,N_24536,N_24996);
nand UO_97 (O_97,N_24666,N_24538);
xor UO_98 (O_98,N_24596,N_24872);
or UO_99 (O_99,N_24705,N_24834);
nor UO_100 (O_100,N_24715,N_24542);
nor UO_101 (O_101,N_24549,N_24584);
and UO_102 (O_102,N_24839,N_24841);
or UO_103 (O_103,N_24906,N_24518);
or UO_104 (O_104,N_24570,N_24670);
nand UO_105 (O_105,N_24682,N_24847);
nand UO_106 (O_106,N_24932,N_24959);
nand UO_107 (O_107,N_24742,N_24920);
nor UO_108 (O_108,N_24879,N_24792);
nor UO_109 (O_109,N_24618,N_24679);
nor UO_110 (O_110,N_24960,N_24778);
nor UO_111 (O_111,N_24780,N_24961);
xor UO_112 (O_112,N_24927,N_24793);
nand UO_113 (O_113,N_24649,N_24576);
nand UO_114 (O_114,N_24893,N_24869);
nor UO_115 (O_115,N_24642,N_24917);
nand UO_116 (O_116,N_24824,N_24575);
xor UO_117 (O_117,N_24750,N_24969);
and UO_118 (O_118,N_24867,N_24776);
nand UO_119 (O_119,N_24829,N_24845);
nand UO_120 (O_120,N_24734,N_24757);
or UO_121 (O_121,N_24572,N_24835);
xor UO_122 (O_122,N_24512,N_24786);
nand UO_123 (O_123,N_24881,N_24875);
nand UO_124 (O_124,N_24814,N_24676);
and UO_125 (O_125,N_24766,N_24657);
and UO_126 (O_126,N_24506,N_24760);
nor UO_127 (O_127,N_24738,N_24731);
nand UO_128 (O_128,N_24946,N_24653);
or UO_129 (O_129,N_24680,N_24508);
nor UO_130 (O_130,N_24905,N_24531);
and UO_131 (O_131,N_24885,N_24637);
and UO_132 (O_132,N_24636,N_24916);
and UO_133 (O_133,N_24514,N_24753);
and UO_134 (O_134,N_24901,N_24890);
and UO_135 (O_135,N_24578,N_24842);
nor UO_136 (O_136,N_24744,N_24758);
and UO_137 (O_137,N_24732,N_24537);
nand UO_138 (O_138,N_24672,N_24944);
nor UO_139 (O_139,N_24587,N_24654);
nor UO_140 (O_140,N_24999,N_24701);
nand UO_141 (O_141,N_24865,N_24922);
nand UO_142 (O_142,N_24992,N_24726);
nand UO_143 (O_143,N_24880,N_24779);
xnor UO_144 (O_144,N_24987,N_24772);
nand UO_145 (O_145,N_24809,N_24511);
or UO_146 (O_146,N_24558,N_24560);
or UO_147 (O_147,N_24810,N_24501);
and UO_148 (O_148,N_24647,N_24521);
nand UO_149 (O_149,N_24816,N_24967);
or UO_150 (O_150,N_24631,N_24769);
nand UO_151 (O_151,N_24854,N_24534);
and UO_152 (O_152,N_24907,N_24923);
nand UO_153 (O_153,N_24870,N_24721);
nor UO_154 (O_154,N_24681,N_24725);
or UO_155 (O_155,N_24949,N_24645);
xor UO_156 (O_156,N_24889,N_24673);
nor UO_157 (O_157,N_24817,N_24791);
xor UO_158 (O_158,N_24868,N_24684);
nor UO_159 (O_159,N_24768,N_24635);
and UO_160 (O_160,N_24526,N_24972);
and UO_161 (O_161,N_24709,N_24971);
nand UO_162 (O_162,N_24919,N_24505);
or UO_163 (O_163,N_24989,N_24546);
nand UO_164 (O_164,N_24703,N_24548);
or UO_165 (O_165,N_24784,N_24698);
nor UO_166 (O_166,N_24801,N_24523);
and UO_167 (O_167,N_24545,N_24748);
nand UO_168 (O_168,N_24581,N_24627);
or UO_169 (O_169,N_24752,N_24812);
and UO_170 (O_170,N_24539,N_24788);
and UO_171 (O_171,N_24914,N_24948);
nor UO_172 (O_172,N_24899,N_24985);
xor UO_173 (O_173,N_24739,N_24953);
or UO_174 (O_174,N_24728,N_24795);
and UO_175 (O_175,N_24594,N_24926);
nor UO_176 (O_176,N_24712,N_24856);
nor UO_177 (O_177,N_24908,N_24622);
nor UO_178 (O_178,N_24777,N_24864);
xor UO_179 (O_179,N_24799,N_24749);
or UO_180 (O_180,N_24559,N_24656);
nor UO_181 (O_181,N_24882,N_24533);
or UO_182 (O_182,N_24929,N_24765);
xnor UO_183 (O_183,N_24770,N_24602);
nor UO_184 (O_184,N_24806,N_24632);
nand UO_185 (O_185,N_24616,N_24614);
nand UO_186 (O_186,N_24982,N_24599);
or UO_187 (O_187,N_24807,N_24675);
or UO_188 (O_188,N_24962,N_24849);
or UO_189 (O_189,N_24945,N_24513);
nor UO_190 (O_190,N_24915,N_24774);
nand UO_191 (O_191,N_24569,N_24846);
or UO_192 (O_192,N_24771,N_24722);
xor UO_193 (O_193,N_24566,N_24641);
and UO_194 (O_194,N_24977,N_24866);
and UO_195 (O_195,N_24815,N_24617);
and UO_196 (O_196,N_24678,N_24692);
and UO_197 (O_197,N_24571,N_24502);
nor UO_198 (O_198,N_24911,N_24608);
nor UO_199 (O_199,N_24773,N_24895);
xnor UO_200 (O_200,N_24659,N_24589);
or UO_201 (O_201,N_24524,N_24794);
nand UO_202 (O_202,N_24988,N_24711);
and UO_203 (O_203,N_24551,N_24547);
nand UO_204 (O_204,N_24781,N_24955);
xor UO_205 (O_205,N_24903,N_24782);
and UO_206 (O_206,N_24900,N_24595);
or UO_207 (O_207,N_24813,N_24588);
or UO_208 (O_208,N_24918,N_24544);
nand UO_209 (O_209,N_24597,N_24574);
nor UO_210 (O_210,N_24860,N_24662);
nand UO_211 (O_211,N_24658,N_24951);
xnor UO_212 (O_212,N_24700,N_24767);
nand UO_213 (O_213,N_24827,N_24651);
or UO_214 (O_214,N_24730,N_24798);
nand UO_215 (O_215,N_24871,N_24892);
or UO_216 (O_216,N_24852,N_24737);
nand UO_217 (O_217,N_24785,N_24837);
nor UO_218 (O_218,N_24668,N_24665);
nor UO_219 (O_219,N_24626,N_24630);
or UO_220 (O_220,N_24563,N_24568);
and UO_221 (O_221,N_24677,N_24593);
nand UO_222 (O_222,N_24896,N_24991);
nor UO_223 (O_223,N_24629,N_24894);
or UO_224 (O_224,N_24848,N_24925);
nand UO_225 (O_225,N_24554,N_24970);
nand UO_226 (O_226,N_24613,N_24741);
nand UO_227 (O_227,N_24993,N_24686);
and UO_228 (O_228,N_24897,N_24720);
or UO_229 (O_229,N_24762,N_24604);
and UO_230 (O_230,N_24940,N_24598);
nand UO_231 (O_231,N_24823,N_24983);
and UO_232 (O_232,N_24966,N_24803);
and UO_233 (O_233,N_24586,N_24950);
nand UO_234 (O_234,N_24990,N_24573);
or UO_235 (O_235,N_24797,N_24783);
or UO_236 (O_236,N_24562,N_24836);
or UO_237 (O_237,N_24605,N_24567);
and UO_238 (O_238,N_24838,N_24789);
nand UO_239 (O_239,N_24957,N_24775);
xor UO_240 (O_240,N_24519,N_24804);
nand UO_241 (O_241,N_24764,N_24582);
xnor UO_242 (O_242,N_24724,N_24543);
nand UO_243 (O_243,N_24704,N_24984);
or UO_244 (O_244,N_24980,N_24853);
nand UO_245 (O_245,N_24802,N_24979);
or UO_246 (O_246,N_24639,N_24625);
nand UO_247 (O_247,N_24909,N_24937);
nor UO_248 (O_248,N_24832,N_24646);
xnor UO_249 (O_249,N_24754,N_24850);
nor UO_250 (O_250,N_24658,N_24664);
nor UO_251 (O_251,N_24663,N_24539);
nor UO_252 (O_252,N_24996,N_24947);
or UO_253 (O_253,N_24764,N_24822);
nor UO_254 (O_254,N_24569,N_24558);
nor UO_255 (O_255,N_24565,N_24704);
nor UO_256 (O_256,N_24879,N_24766);
and UO_257 (O_257,N_24797,N_24670);
and UO_258 (O_258,N_24774,N_24886);
and UO_259 (O_259,N_24881,N_24826);
and UO_260 (O_260,N_24860,N_24633);
and UO_261 (O_261,N_24845,N_24939);
xor UO_262 (O_262,N_24924,N_24820);
nand UO_263 (O_263,N_24760,N_24998);
nand UO_264 (O_264,N_24559,N_24573);
and UO_265 (O_265,N_24985,N_24864);
or UO_266 (O_266,N_24647,N_24703);
and UO_267 (O_267,N_24955,N_24817);
or UO_268 (O_268,N_24810,N_24591);
nor UO_269 (O_269,N_24586,N_24879);
xnor UO_270 (O_270,N_24835,N_24500);
nand UO_271 (O_271,N_24722,N_24953);
xnor UO_272 (O_272,N_24918,N_24624);
nand UO_273 (O_273,N_24843,N_24968);
nor UO_274 (O_274,N_24553,N_24793);
or UO_275 (O_275,N_24671,N_24987);
nand UO_276 (O_276,N_24998,N_24526);
and UO_277 (O_277,N_24557,N_24509);
or UO_278 (O_278,N_24703,N_24762);
xor UO_279 (O_279,N_24768,N_24805);
nor UO_280 (O_280,N_24549,N_24899);
nor UO_281 (O_281,N_24628,N_24946);
and UO_282 (O_282,N_24639,N_24844);
and UO_283 (O_283,N_24548,N_24633);
nand UO_284 (O_284,N_24860,N_24864);
or UO_285 (O_285,N_24684,N_24930);
or UO_286 (O_286,N_24629,N_24869);
nor UO_287 (O_287,N_24559,N_24754);
nand UO_288 (O_288,N_24676,N_24690);
xor UO_289 (O_289,N_24563,N_24570);
xnor UO_290 (O_290,N_24672,N_24939);
nand UO_291 (O_291,N_24994,N_24888);
xor UO_292 (O_292,N_24973,N_24908);
and UO_293 (O_293,N_24597,N_24656);
and UO_294 (O_294,N_24514,N_24805);
nor UO_295 (O_295,N_24825,N_24546);
and UO_296 (O_296,N_24991,N_24975);
nor UO_297 (O_297,N_24891,N_24779);
nor UO_298 (O_298,N_24736,N_24846);
nand UO_299 (O_299,N_24981,N_24568);
and UO_300 (O_300,N_24596,N_24732);
nand UO_301 (O_301,N_24845,N_24811);
or UO_302 (O_302,N_24971,N_24665);
nand UO_303 (O_303,N_24985,N_24788);
nor UO_304 (O_304,N_24848,N_24681);
or UO_305 (O_305,N_24946,N_24986);
nor UO_306 (O_306,N_24879,N_24953);
and UO_307 (O_307,N_24547,N_24990);
or UO_308 (O_308,N_24650,N_24815);
xor UO_309 (O_309,N_24919,N_24713);
nand UO_310 (O_310,N_24802,N_24864);
or UO_311 (O_311,N_24887,N_24811);
nand UO_312 (O_312,N_24754,N_24565);
and UO_313 (O_313,N_24792,N_24501);
nor UO_314 (O_314,N_24635,N_24652);
or UO_315 (O_315,N_24587,N_24719);
and UO_316 (O_316,N_24739,N_24631);
and UO_317 (O_317,N_24973,N_24805);
or UO_318 (O_318,N_24967,N_24852);
nand UO_319 (O_319,N_24800,N_24987);
nand UO_320 (O_320,N_24895,N_24763);
nor UO_321 (O_321,N_24575,N_24548);
or UO_322 (O_322,N_24688,N_24820);
or UO_323 (O_323,N_24803,N_24971);
or UO_324 (O_324,N_24959,N_24963);
and UO_325 (O_325,N_24980,N_24509);
or UO_326 (O_326,N_24892,N_24969);
or UO_327 (O_327,N_24735,N_24892);
nand UO_328 (O_328,N_24608,N_24891);
or UO_329 (O_329,N_24504,N_24822);
and UO_330 (O_330,N_24908,N_24676);
or UO_331 (O_331,N_24635,N_24984);
nand UO_332 (O_332,N_24978,N_24795);
xor UO_333 (O_333,N_24577,N_24836);
xor UO_334 (O_334,N_24616,N_24812);
and UO_335 (O_335,N_24969,N_24943);
nor UO_336 (O_336,N_24548,N_24963);
and UO_337 (O_337,N_24890,N_24889);
nand UO_338 (O_338,N_24571,N_24965);
nand UO_339 (O_339,N_24704,N_24727);
and UO_340 (O_340,N_24846,N_24803);
nor UO_341 (O_341,N_24567,N_24798);
or UO_342 (O_342,N_24747,N_24818);
and UO_343 (O_343,N_24574,N_24901);
nor UO_344 (O_344,N_24937,N_24822);
nor UO_345 (O_345,N_24634,N_24772);
and UO_346 (O_346,N_24865,N_24788);
or UO_347 (O_347,N_24838,N_24823);
and UO_348 (O_348,N_24735,N_24634);
and UO_349 (O_349,N_24895,N_24877);
nor UO_350 (O_350,N_24520,N_24753);
nand UO_351 (O_351,N_24761,N_24904);
or UO_352 (O_352,N_24911,N_24852);
nand UO_353 (O_353,N_24806,N_24574);
nand UO_354 (O_354,N_24911,N_24831);
nor UO_355 (O_355,N_24692,N_24936);
or UO_356 (O_356,N_24730,N_24603);
and UO_357 (O_357,N_24516,N_24766);
and UO_358 (O_358,N_24677,N_24653);
nor UO_359 (O_359,N_24718,N_24551);
and UO_360 (O_360,N_24720,N_24722);
and UO_361 (O_361,N_24644,N_24606);
nand UO_362 (O_362,N_24517,N_24788);
and UO_363 (O_363,N_24760,N_24755);
nand UO_364 (O_364,N_24814,N_24843);
nor UO_365 (O_365,N_24699,N_24515);
or UO_366 (O_366,N_24732,N_24769);
or UO_367 (O_367,N_24877,N_24793);
and UO_368 (O_368,N_24635,N_24606);
xor UO_369 (O_369,N_24953,N_24884);
nor UO_370 (O_370,N_24841,N_24909);
and UO_371 (O_371,N_24560,N_24605);
or UO_372 (O_372,N_24554,N_24889);
nor UO_373 (O_373,N_24774,N_24948);
and UO_374 (O_374,N_24578,N_24785);
nor UO_375 (O_375,N_24616,N_24569);
and UO_376 (O_376,N_24743,N_24831);
and UO_377 (O_377,N_24538,N_24577);
nor UO_378 (O_378,N_24756,N_24973);
or UO_379 (O_379,N_24664,N_24880);
nor UO_380 (O_380,N_24669,N_24721);
nor UO_381 (O_381,N_24592,N_24600);
nor UO_382 (O_382,N_24752,N_24917);
or UO_383 (O_383,N_24521,N_24903);
nand UO_384 (O_384,N_24749,N_24582);
nand UO_385 (O_385,N_24917,N_24904);
nand UO_386 (O_386,N_24793,N_24913);
or UO_387 (O_387,N_24621,N_24886);
nor UO_388 (O_388,N_24849,N_24884);
nand UO_389 (O_389,N_24798,N_24754);
nor UO_390 (O_390,N_24510,N_24783);
xnor UO_391 (O_391,N_24532,N_24765);
or UO_392 (O_392,N_24919,N_24544);
nor UO_393 (O_393,N_24546,N_24720);
or UO_394 (O_394,N_24573,N_24561);
or UO_395 (O_395,N_24626,N_24947);
nand UO_396 (O_396,N_24704,N_24944);
and UO_397 (O_397,N_24641,N_24556);
nor UO_398 (O_398,N_24916,N_24573);
or UO_399 (O_399,N_24782,N_24712);
or UO_400 (O_400,N_24603,N_24502);
or UO_401 (O_401,N_24839,N_24802);
or UO_402 (O_402,N_24554,N_24965);
nand UO_403 (O_403,N_24703,N_24680);
or UO_404 (O_404,N_24789,N_24602);
and UO_405 (O_405,N_24503,N_24769);
or UO_406 (O_406,N_24680,N_24794);
or UO_407 (O_407,N_24929,N_24607);
or UO_408 (O_408,N_24669,N_24584);
nor UO_409 (O_409,N_24819,N_24775);
nand UO_410 (O_410,N_24727,N_24521);
and UO_411 (O_411,N_24987,N_24938);
nand UO_412 (O_412,N_24959,N_24522);
xnor UO_413 (O_413,N_24886,N_24842);
or UO_414 (O_414,N_24513,N_24958);
nand UO_415 (O_415,N_24993,N_24810);
and UO_416 (O_416,N_24719,N_24718);
or UO_417 (O_417,N_24557,N_24818);
nor UO_418 (O_418,N_24797,N_24896);
and UO_419 (O_419,N_24515,N_24717);
or UO_420 (O_420,N_24837,N_24583);
nand UO_421 (O_421,N_24638,N_24652);
or UO_422 (O_422,N_24525,N_24932);
or UO_423 (O_423,N_24678,N_24572);
nor UO_424 (O_424,N_24730,N_24997);
or UO_425 (O_425,N_24535,N_24578);
nor UO_426 (O_426,N_24790,N_24922);
and UO_427 (O_427,N_24800,N_24594);
nor UO_428 (O_428,N_24691,N_24997);
nor UO_429 (O_429,N_24912,N_24735);
or UO_430 (O_430,N_24981,N_24842);
nor UO_431 (O_431,N_24909,N_24742);
or UO_432 (O_432,N_24830,N_24501);
or UO_433 (O_433,N_24501,N_24787);
nor UO_434 (O_434,N_24839,N_24709);
nor UO_435 (O_435,N_24571,N_24612);
nand UO_436 (O_436,N_24951,N_24547);
xnor UO_437 (O_437,N_24770,N_24977);
or UO_438 (O_438,N_24593,N_24619);
and UO_439 (O_439,N_24534,N_24640);
or UO_440 (O_440,N_24746,N_24786);
and UO_441 (O_441,N_24960,N_24648);
and UO_442 (O_442,N_24692,N_24512);
nand UO_443 (O_443,N_24588,N_24762);
nor UO_444 (O_444,N_24584,N_24949);
and UO_445 (O_445,N_24884,N_24893);
nand UO_446 (O_446,N_24971,N_24827);
nor UO_447 (O_447,N_24904,N_24659);
or UO_448 (O_448,N_24912,N_24986);
nand UO_449 (O_449,N_24910,N_24819);
nand UO_450 (O_450,N_24768,N_24621);
nand UO_451 (O_451,N_24811,N_24999);
or UO_452 (O_452,N_24707,N_24635);
and UO_453 (O_453,N_24827,N_24769);
nand UO_454 (O_454,N_24937,N_24747);
nor UO_455 (O_455,N_24560,N_24632);
xnor UO_456 (O_456,N_24650,N_24571);
nand UO_457 (O_457,N_24600,N_24502);
nor UO_458 (O_458,N_24668,N_24614);
nand UO_459 (O_459,N_24680,N_24588);
nor UO_460 (O_460,N_24509,N_24953);
nor UO_461 (O_461,N_24906,N_24968);
xnor UO_462 (O_462,N_24614,N_24758);
nor UO_463 (O_463,N_24827,N_24778);
or UO_464 (O_464,N_24727,N_24525);
nor UO_465 (O_465,N_24739,N_24768);
nor UO_466 (O_466,N_24626,N_24602);
nand UO_467 (O_467,N_24586,N_24906);
nor UO_468 (O_468,N_24701,N_24923);
or UO_469 (O_469,N_24610,N_24891);
and UO_470 (O_470,N_24679,N_24731);
nor UO_471 (O_471,N_24769,N_24544);
nand UO_472 (O_472,N_24792,N_24906);
and UO_473 (O_473,N_24905,N_24640);
nor UO_474 (O_474,N_24598,N_24822);
or UO_475 (O_475,N_24998,N_24589);
or UO_476 (O_476,N_24737,N_24877);
or UO_477 (O_477,N_24677,N_24940);
or UO_478 (O_478,N_24696,N_24855);
nor UO_479 (O_479,N_24689,N_24584);
or UO_480 (O_480,N_24882,N_24812);
nor UO_481 (O_481,N_24997,N_24524);
xnor UO_482 (O_482,N_24973,N_24605);
nor UO_483 (O_483,N_24911,N_24809);
xnor UO_484 (O_484,N_24817,N_24985);
nor UO_485 (O_485,N_24668,N_24779);
or UO_486 (O_486,N_24764,N_24991);
or UO_487 (O_487,N_24934,N_24514);
xnor UO_488 (O_488,N_24674,N_24605);
nor UO_489 (O_489,N_24988,N_24908);
nor UO_490 (O_490,N_24526,N_24931);
nor UO_491 (O_491,N_24848,N_24717);
nor UO_492 (O_492,N_24588,N_24881);
or UO_493 (O_493,N_24977,N_24845);
and UO_494 (O_494,N_24571,N_24854);
nand UO_495 (O_495,N_24755,N_24841);
and UO_496 (O_496,N_24778,N_24952);
nor UO_497 (O_497,N_24714,N_24598);
or UO_498 (O_498,N_24940,N_24524);
or UO_499 (O_499,N_24545,N_24994);
xor UO_500 (O_500,N_24688,N_24589);
nand UO_501 (O_501,N_24903,N_24749);
and UO_502 (O_502,N_24866,N_24958);
nor UO_503 (O_503,N_24572,N_24612);
and UO_504 (O_504,N_24913,N_24923);
xnor UO_505 (O_505,N_24962,N_24572);
and UO_506 (O_506,N_24679,N_24799);
nand UO_507 (O_507,N_24839,N_24693);
xnor UO_508 (O_508,N_24583,N_24824);
or UO_509 (O_509,N_24916,N_24801);
and UO_510 (O_510,N_24701,N_24941);
nor UO_511 (O_511,N_24773,N_24685);
or UO_512 (O_512,N_24695,N_24792);
and UO_513 (O_513,N_24595,N_24963);
or UO_514 (O_514,N_24959,N_24595);
nand UO_515 (O_515,N_24704,N_24961);
or UO_516 (O_516,N_24975,N_24983);
nor UO_517 (O_517,N_24657,N_24576);
or UO_518 (O_518,N_24835,N_24783);
and UO_519 (O_519,N_24851,N_24673);
or UO_520 (O_520,N_24612,N_24834);
nor UO_521 (O_521,N_24509,N_24798);
or UO_522 (O_522,N_24528,N_24534);
nand UO_523 (O_523,N_24519,N_24772);
or UO_524 (O_524,N_24947,N_24863);
and UO_525 (O_525,N_24506,N_24610);
nand UO_526 (O_526,N_24734,N_24911);
and UO_527 (O_527,N_24524,N_24775);
nor UO_528 (O_528,N_24544,N_24624);
or UO_529 (O_529,N_24799,N_24829);
nor UO_530 (O_530,N_24564,N_24742);
nand UO_531 (O_531,N_24704,N_24639);
nor UO_532 (O_532,N_24599,N_24797);
and UO_533 (O_533,N_24737,N_24661);
or UO_534 (O_534,N_24846,N_24741);
and UO_535 (O_535,N_24863,N_24738);
or UO_536 (O_536,N_24600,N_24936);
nor UO_537 (O_537,N_24705,N_24563);
nand UO_538 (O_538,N_24789,N_24615);
nor UO_539 (O_539,N_24644,N_24952);
nand UO_540 (O_540,N_24676,N_24853);
nand UO_541 (O_541,N_24596,N_24850);
nand UO_542 (O_542,N_24832,N_24688);
and UO_543 (O_543,N_24535,N_24584);
xnor UO_544 (O_544,N_24917,N_24950);
nor UO_545 (O_545,N_24519,N_24666);
and UO_546 (O_546,N_24604,N_24523);
or UO_547 (O_547,N_24996,N_24702);
and UO_548 (O_548,N_24698,N_24556);
nor UO_549 (O_549,N_24874,N_24635);
nor UO_550 (O_550,N_24717,N_24862);
nand UO_551 (O_551,N_24658,N_24803);
nor UO_552 (O_552,N_24783,N_24989);
nand UO_553 (O_553,N_24848,N_24804);
nand UO_554 (O_554,N_24620,N_24753);
and UO_555 (O_555,N_24680,N_24884);
nor UO_556 (O_556,N_24954,N_24825);
xnor UO_557 (O_557,N_24824,N_24570);
and UO_558 (O_558,N_24968,N_24567);
nand UO_559 (O_559,N_24895,N_24757);
or UO_560 (O_560,N_24854,N_24662);
nand UO_561 (O_561,N_24861,N_24680);
or UO_562 (O_562,N_24991,N_24905);
or UO_563 (O_563,N_24895,N_24732);
xnor UO_564 (O_564,N_24677,N_24781);
nand UO_565 (O_565,N_24980,N_24820);
nor UO_566 (O_566,N_24954,N_24864);
or UO_567 (O_567,N_24947,N_24724);
nand UO_568 (O_568,N_24598,N_24911);
and UO_569 (O_569,N_24632,N_24620);
nor UO_570 (O_570,N_24602,N_24520);
nand UO_571 (O_571,N_24921,N_24553);
nand UO_572 (O_572,N_24924,N_24915);
or UO_573 (O_573,N_24636,N_24594);
nor UO_574 (O_574,N_24654,N_24876);
or UO_575 (O_575,N_24959,N_24857);
nand UO_576 (O_576,N_24566,N_24931);
or UO_577 (O_577,N_24813,N_24752);
nand UO_578 (O_578,N_24536,N_24819);
and UO_579 (O_579,N_24696,N_24767);
and UO_580 (O_580,N_24919,N_24788);
nor UO_581 (O_581,N_24889,N_24762);
or UO_582 (O_582,N_24720,N_24998);
nor UO_583 (O_583,N_24917,N_24872);
nor UO_584 (O_584,N_24735,N_24515);
or UO_585 (O_585,N_24848,N_24744);
nor UO_586 (O_586,N_24781,N_24576);
and UO_587 (O_587,N_24501,N_24864);
nand UO_588 (O_588,N_24637,N_24513);
nor UO_589 (O_589,N_24811,N_24690);
nor UO_590 (O_590,N_24877,N_24516);
nor UO_591 (O_591,N_24641,N_24555);
nand UO_592 (O_592,N_24580,N_24598);
or UO_593 (O_593,N_24990,N_24988);
or UO_594 (O_594,N_24825,N_24890);
and UO_595 (O_595,N_24918,N_24851);
nand UO_596 (O_596,N_24843,N_24519);
or UO_597 (O_597,N_24567,N_24570);
nand UO_598 (O_598,N_24982,N_24853);
or UO_599 (O_599,N_24935,N_24778);
and UO_600 (O_600,N_24842,N_24977);
nand UO_601 (O_601,N_24783,N_24773);
nand UO_602 (O_602,N_24542,N_24580);
nand UO_603 (O_603,N_24938,N_24766);
xnor UO_604 (O_604,N_24926,N_24746);
nor UO_605 (O_605,N_24906,N_24780);
xnor UO_606 (O_606,N_24877,N_24927);
nor UO_607 (O_607,N_24932,N_24662);
or UO_608 (O_608,N_24702,N_24673);
and UO_609 (O_609,N_24959,N_24979);
nor UO_610 (O_610,N_24616,N_24860);
nand UO_611 (O_611,N_24977,N_24562);
nand UO_612 (O_612,N_24534,N_24716);
nand UO_613 (O_613,N_24634,N_24646);
or UO_614 (O_614,N_24583,N_24590);
and UO_615 (O_615,N_24622,N_24726);
nor UO_616 (O_616,N_24987,N_24698);
or UO_617 (O_617,N_24570,N_24913);
nand UO_618 (O_618,N_24680,N_24653);
and UO_619 (O_619,N_24886,N_24915);
nor UO_620 (O_620,N_24729,N_24674);
nand UO_621 (O_621,N_24677,N_24914);
or UO_622 (O_622,N_24575,N_24771);
nor UO_623 (O_623,N_24901,N_24647);
xor UO_624 (O_624,N_24835,N_24513);
or UO_625 (O_625,N_24870,N_24591);
or UO_626 (O_626,N_24909,N_24706);
or UO_627 (O_627,N_24663,N_24819);
nor UO_628 (O_628,N_24617,N_24982);
or UO_629 (O_629,N_24727,N_24717);
nor UO_630 (O_630,N_24856,N_24648);
and UO_631 (O_631,N_24733,N_24504);
nand UO_632 (O_632,N_24772,N_24754);
nor UO_633 (O_633,N_24742,N_24613);
or UO_634 (O_634,N_24707,N_24959);
or UO_635 (O_635,N_24852,N_24538);
and UO_636 (O_636,N_24925,N_24596);
and UO_637 (O_637,N_24881,N_24582);
nor UO_638 (O_638,N_24823,N_24709);
xnor UO_639 (O_639,N_24868,N_24864);
and UO_640 (O_640,N_24880,N_24862);
nand UO_641 (O_641,N_24824,N_24982);
nor UO_642 (O_642,N_24816,N_24916);
and UO_643 (O_643,N_24947,N_24953);
or UO_644 (O_644,N_24617,N_24814);
xor UO_645 (O_645,N_24820,N_24972);
and UO_646 (O_646,N_24841,N_24928);
nor UO_647 (O_647,N_24677,N_24865);
or UO_648 (O_648,N_24593,N_24777);
nor UO_649 (O_649,N_24783,N_24815);
nand UO_650 (O_650,N_24531,N_24692);
nor UO_651 (O_651,N_24550,N_24593);
and UO_652 (O_652,N_24724,N_24900);
nand UO_653 (O_653,N_24884,N_24617);
and UO_654 (O_654,N_24805,N_24538);
nor UO_655 (O_655,N_24741,N_24719);
and UO_656 (O_656,N_24629,N_24931);
nand UO_657 (O_657,N_24926,N_24975);
nand UO_658 (O_658,N_24898,N_24876);
or UO_659 (O_659,N_24772,N_24920);
xnor UO_660 (O_660,N_24838,N_24803);
nor UO_661 (O_661,N_24536,N_24672);
xor UO_662 (O_662,N_24999,N_24784);
nor UO_663 (O_663,N_24950,N_24954);
nor UO_664 (O_664,N_24728,N_24679);
and UO_665 (O_665,N_24862,N_24628);
or UO_666 (O_666,N_24583,N_24636);
nor UO_667 (O_667,N_24581,N_24736);
or UO_668 (O_668,N_24977,N_24654);
or UO_669 (O_669,N_24706,N_24786);
and UO_670 (O_670,N_24773,N_24908);
nor UO_671 (O_671,N_24860,N_24588);
nor UO_672 (O_672,N_24859,N_24626);
xor UO_673 (O_673,N_24880,N_24981);
nand UO_674 (O_674,N_24846,N_24609);
nand UO_675 (O_675,N_24786,N_24992);
xor UO_676 (O_676,N_24594,N_24745);
nor UO_677 (O_677,N_24608,N_24898);
and UO_678 (O_678,N_24945,N_24918);
nand UO_679 (O_679,N_24724,N_24961);
nand UO_680 (O_680,N_24689,N_24620);
and UO_681 (O_681,N_24605,N_24647);
nor UO_682 (O_682,N_24688,N_24627);
or UO_683 (O_683,N_24671,N_24928);
and UO_684 (O_684,N_24911,N_24581);
nand UO_685 (O_685,N_24828,N_24952);
or UO_686 (O_686,N_24973,N_24919);
nand UO_687 (O_687,N_24797,N_24820);
nor UO_688 (O_688,N_24843,N_24704);
nand UO_689 (O_689,N_24840,N_24622);
nand UO_690 (O_690,N_24567,N_24679);
or UO_691 (O_691,N_24640,N_24593);
and UO_692 (O_692,N_24815,N_24778);
and UO_693 (O_693,N_24985,N_24963);
nand UO_694 (O_694,N_24858,N_24689);
nand UO_695 (O_695,N_24648,N_24504);
nor UO_696 (O_696,N_24718,N_24777);
and UO_697 (O_697,N_24575,N_24560);
or UO_698 (O_698,N_24877,N_24523);
nor UO_699 (O_699,N_24871,N_24837);
nor UO_700 (O_700,N_24683,N_24965);
nor UO_701 (O_701,N_24643,N_24644);
xor UO_702 (O_702,N_24871,N_24547);
and UO_703 (O_703,N_24509,N_24872);
nor UO_704 (O_704,N_24619,N_24900);
and UO_705 (O_705,N_24904,N_24571);
nor UO_706 (O_706,N_24867,N_24648);
nor UO_707 (O_707,N_24889,N_24777);
nand UO_708 (O_708,N_24648,N_24825);
and UO_709 (O_709,N_24638,N_24533);
nor UO_710 (O_710,N_24729,N_24576);
xor UO_711 (O_711,N_24829,N_24744);
or UO_712 (O_712,N_24660,N_24913);
or UO_713 (O_713,N_24680,N_24545);
or UO_714 (O_714,N_24661,N_24727);
or UO_715 (O_715,N_24589,N_24986);
nand UO_716 (O_716,N_24523,N_24976);
nand UO_717 (O_717,N_24950,N_24988);
and UO_718 (O_718,N_24642,N_24747);
and UO_719 (O_719,N_24720,N_24733);
nand UO_720 (O_720,N_24631,N_24672);
or UO_721 (O_721,N_24609,N_24699);
nor UO_722 (O_722,N_24847,N_24858);
or UO_723 (O_723,N_24756,N_24734);
nor UO_724 (O_724,N_24764,N_24657);
or UO_725 (O_725,N_24890,N_24820);
nand UO_726 (O_726,N_24553,N_24509);
and UO_727 (O_727,N_24716,N_24583);
nand UO_728 (O_728,N_24603,N_24874);
or UO_729 (O_729,N_24584,N_24550);
and UO_730 (O_730,N_24812,N_24599);
xnor UO_731 (O_731,N_24585,N_24946);
or UO_732 (O_732,N_24633,N_24835);
and UO_733 (O_733,N_24872,N_24827);
or UO_734 (O_734,N_24896,N_24651);
and UO_735 (O_735,N_24616,N_24733);
or UO_736 (O_736,N_24586,N_24710);
and UO_737 (O_737,N_24504,N_24770);
or UO_738 (O_738,N_24913,N_24910);
nand UO_739 (O_739,N_24672,N_24533);
and UO_740 (O_740,N_24925,N_24560);
or UO_741 (O_741,N_24517,N_24612);
or UO_742 (O_742,N_24622,N_24819);
or UO_743 (O_743,N_24972,N_24678);
nand UO_744 (O_744,N_24810,N_24515);
or UO_745 (O_745,N_24837,N_24621);
nor UO_746 (O_746,N_24826,N_24740);
and UO_747 (O_747,N_24901,N_24820);
nor UO_748 (O_748,N_24823,N_24501);
and UO_749 (O_749,N_24520,N_24917);
xor UO_750 (O_750,N_24552,N_24844);
nand UO_751 (O_751,N_24525,N_24521);
nor UO_752 (O_752,N_24643,N_24989);
or UO_753 (O_753,N_24629,N_24746);
nand UO_754 (O_754,N_24719,N_24998);
and UO_755 (O_755,N_24523,N_24514);
nand UO_756 (O_756,N_24666,N_24887);
and UO_757 (O_757,N_24856,N_24716);
and UO_758 (O_758,N_24721,N_24928);
or UO_759 (O_759,N_24716,N_24921);
nand UO_760 (O_760,N_24747,N_24677);
or UO_761 (O_761,N_24880,N_24866);
nand UO_762 (O_762,N_24576,N_24974);
and UO_763 (O_763,N_24630,N_24789);
and UO_764 (O_764,N_24894,N_24931);
and UO_765 (O_765,N_24811,N_24806);
nand UO_766 (O_766,N_24693,N_24785);
and UO_767 (O_767,N_24995,N_24588);
nand UO_768 (O_768,N_24577,N_24775);
nand UO_769 (O_769,N_24937,N_24728);
or UO_770 (O_770,N_24734,N_24559);
and UO_771 (O_771,N_24925,N_24718);
or UO_772 (O_772,N_24868,N_24504);
and UO_773 (O_773,N_24737,N_24798);
nor UO_774 (O_774,N_24713,N_24686);
or UO_775 (O_775,N_24790,N_24821);
nor UO_776 (O_776,N_24656,N_24628);
nand UO_777 (O_777,N_24859,N_24723);
or UO_778 (O_778,N_24656,N_24633);
nor UO_779 (O_779,N_24703,N_24691);
xor UO_780 (O_780,N_24663,N_24652);
and UO_781 (O_781,N_24501,N_24646);
xnor UO_782 (O_782,N_24532,N_24924);
xnor UO_783 (O_783,N_24778,N_24692);
nor UO_784 (O_784,N_24949,N_24715);
and UO_785 (O_785,N_24686,N_24694);
nor UO_786 (O_786,N_24541,N_24691);
or UO_787 (O_787,N_24867,N_24964);
or UO_788 (O_788,N_24705,N_24968);
xnor UO_789 (O_789,N_24923,N_24722);
or UO_790 (O_790,N_24644,N_24771);
nand UO_791 (O_791,N_24569,N_24833);
or UO_792 (O_792,N_24876,N_24775);
or UO_793 (O_793,N_24523,N_24503);
and UO_794 (O_794,N_24820,N_24690);
or UO_795 (O_795,N_24693,N_24917);
and UO_796 (O_796,N_24760,N_24944);
and UO_797 (O_797,N_24672,N_24712);
xnor UO_798 (O_798,N_24811,N_24804);
and UO_799 (O_799,N_24808,N_24825);
nor UO_800 (O_800,N_24937,N_24842);
nor UO_801 (O_801,N_24808,N_24640);
nor UO_802 (O_802,N_24880,N_24985);
xor UO_803 (O_803,N_24933,N_24729);
nor UO_804 (O_804,N_24728,N_24710);
nor UO_805 (O_805,N_24696,N_24898);
nor UO_806 (O_806,N_24654,N_24844);
nor UO_807 (O_807,N_24821,N_24709);
nor UO_808 (O_808,N_24733,N_24772);
nor UO_809 (O_809,N_24694,N_24784);
and UO_810 (O_810,N_24645,N_24510);
nand UO_811 (O_811,N_24542,N_24790);
nand UO_812 (O_812,N_24584,N_24891);
xor UO_813 (O_813,N_24511,N_24573);
nand UO_814 (O_814,N_24591,N_24855);
and UO_815 (O_815,N_24835,N_24560);
and UO_816 (O_816,N_24963,N_24892);
or UO_817 (O_817,N_24594,N_24736);
and UO_818 (O_818,N_24940,N_24926);
or UO_819 (O_819,N_24737,N_24610);
nand UO_820 (O_820,N_24856,N_24972);
nand UO_821 (O_821,N_24927,N_24933);
and UO_822 (O_822,N_24593,N_24675);
nand UO_823 (O_823,N_24943,N_24993);
nor UO_824 (O_824,N_24752,N_24949);
and UO_825 (O_825,N_24829,N_24522);
nand UO_826 (O_826,N_24882,N_24632);
nand UO_827 (O_827,N_24969,N_24663);
nand UO_828 (O_828,N_24659,N_24856);
or UO_829 (O_829,N_24854,N_24543);
nor UO_830 (O_830,N_24649,N_24821);
or UO_831 (O_831,N_24567,N_24783);
nor UO_832 (O_832,N_24564,N_24844);
xnor UO_833 (O_833,N_24791,N_24577);
nor UO_834 (O_834,N_24817,N_24926);
nand UO_835 (O_835,N_24617,N_24599);
nor UO_836 (O_836,N_24599,N_24506);
nor UO_837 (O_837,N_24648,N_24912);
xor UO_838 (O_838,N_24643,N_24704);
nand UO_839 (O_839,N_24974,N_24902);
and UO_840 (O_840,N_24895,N_24665);
or UO_841 (O_841,N_24779,N_24533);
and UO_842 (O_842,N_24825,N_24854);
or UO_843 (O_843,N_24750,N_24978);
nand UO_844 (O_844,N_24912,N_24789);
or UO_845 (O_845,N_24560,N_24912);
nand UO_846 (O_846,N_24777,N_24605);
nor UO_847 (O_847,N_24564,N_24694);
nor UO_848 (O_848,N_24550,N_24580);
nor UO_849 (O_849,N_24902,N_24932);
nor UO_850 (O_850,N_24944,N_24973);
nand UO_851 (O_851,N_24765,N_24632);
xnor UO_852 (O_852,N_24640,N_24832);
or UO_853 (O_853,N_24900,N_24864);
nor UO_854 (O_854,N_24960,N_24881);
or UO_855 (O_855,N_24818,N_24514);
nor UO_856 (O_856,N_24529,N_24556);
nor UO_857 (O_857,N_24645,N_24539);
nor UO_858 (O_858,N_24816,N_24972);
or UO_859 (O_859,N_24736,N_24961);
and UO_860 (O_860,N_24508,N_24991);
and UO_861 (O_861,N_24529,N_24644);
xor UO_862 (O_862,N_24550,N_24716);
nand UO_863 (O_863,N_24863,N_24987);
nand UO_864 (O_864,N_24771,N_24911);
and UO_865 (O_865,N_24898,N_24716);
nor UO_866 (O_866,N_24732,N_24505);
nand UO_867 (O_867,N_24953,N_24984);
nand UO_868 (O_868,N_24798,N_24684);
nand UO_869 (O_869,N_24902,N_24827);
xor UO_870 (O_870,N_24732,N_24786);
nor UO_871 (O_871,N_24881,N_24596);
and UO_872 (O_872,N_24649,N_24653);
nor UO_873 (O_873,N_24713,N_24826);
or UO_874 (O_874,N_24569,N_24824);
nand UO_875 (O_875,N_24872,N_24691);
and UO_876 (O_876,N_24654,N_24532);
nand UO_877 (O_877,N_24951,N_24899);
nor UO_878 (O_878,N_24998,N_24809);
nand UO_879 (O_879,N_24727,N_24699);
and UO_880 (O_880,N_24945,N_24985);
nand UO_881 (O_881,N_24698,N_24840);
nor UO_882 (O_882,N_24715,N_24837);
nor UO_883 (O_883,N_24927,N_24558);
nand UO_884 (O_884,N_24853,N_24857);
and UO_885 (O_885,N_24597,N_24582);
xor UO_886 (O_886,N_24547,N_24623);
and UO_887 (O_887,N_24681,N_24912);
nand UO_888 (O_888,N_24929,N_24967);
or UO_889 (O_889,N_24580,N_24910);
and UO_890 (O_890,N_24987,N_24678);
or UO_891 (O_891,N_24509,N_24772);
xor UO_892 (O_892,N_24726,N_24566);
nand UO_893 (O_893,N_24852,N_24513);
nand UO_894 (O_894,N_24990,N_24828);
and UO_895 (O_895,N_24738,N_24856);
nor UO_896 (O_896,N_24997,N_24990);
and UO_897 (O_897,N_24639,N_24775);
xor UO_898 (O_898,N_24603,N_24959);
and UO_899 (O_899,N_24618,N_24881);
nor UO_900 (O_900,N_24811,N_24916);
xor UO_901 (O_901,N_24709,N_24941);
or UO_902 (O_902,N_24903,N_24586);
nand UO_903 (O_903,N_24934,N_24946);
nand UO_904 (O_904,N_24775,N_24534);
xor UO_905 (O_905,N_24787,N_24891);
nand UO_906 (O_906,N_24511,N_24659);
nor UO_907 (O_907,N_24707,N_24569);
or UO_908 (O_908,N_24856,N_24811);
nor UO_909 (O_909,N_24957,N_24607);
and UO_910 (O_910,N_24953,N_24614);
nor UO_911 (O_911,N_24501,N_24878);
nor UO_912 (O_912,N_24567,N_24976);
nand UO_913 (O_913,N_24580,N_24725);
or UO_914 (O_914,N_24922,N_24723);
and UO_915 (O_915,N_24575,N_24945);
and UO_916 (O_916,N_24500,N_24974);
or UO_917 (O_917,N_24700,N_24615);
nand UO_918 (O_918,N_24536,N_24537);
nand UO_919 (O_919,N_24864,N_24560);
nor UO_920 (O_920,N_24882,N_24740);
and UO_921 (O_921,N_24999,N_24996);
nor UO_922 (O_922,N_24568,N_24747);
and UO_923 (O_923,N_24713,N_24970);
or UO_924 (O_924,N_24831,N_24899);
nor UO_925 (O_925,N_24807,N_24975);
or UO_926 (O_926,N_24990,N_24608);
and UO_927 (O_927,N_24990,N_24901);
or UO_928 (O_928,N_24701,N_24594);
nor UO_929 (O_929,N_24682,N_24573);
nand UO_930 (O_930,N_24565,N_24966);
nor UO_931 (O_931,N_24944,N_24603);
nor UO_932 (O_932,N_24589,N_24989);
xor UO_933 (O_933,N_24919,N_24813);
nand UO_934 (O_934,N_24654,N_24636);
xor UO_935 (O_935,N_24987,N_24651);
and UO_936 (O_936,N_24553,N_24613);
nand UO_937 (O_937,N_24538,N_24691);
or UO_938 (O_938,N_24932,N_24586);
nor UO_939 (O_939,N_24740,N_24747);
or UO_940 (O_940,N_24981,N_24892);
nand UO_941 (O_941,N_24753,N_24750);
nor UO_942 (O_942,N_24692,N_24628);
nand UO_943 (O_943,N_24697,N_24960);
or UO_944 (O_944,N_24784,N_24642);
and UO_945 (O_945,N_24754,N_24682);
nor UO_946 (O_946,N_24621,N_24729);
or UO_947 (O_947,N_24696,N_24585);
nor UO_948 (O_948,N_24822,N_24884);
and UO_949 (O_949,N_24903,N_24701);
nand UO_950 (O_950,N_24906,N_24738);
or UO_951 (O_951,N_24945,N_24652);
or UO_952 (O_952,N_24953,N_24883);
or UO_953 (O_953,N_24785,N_24700);
nand UO_954 (O_954,N_24920,N_24623);
and UO_955 (O_955,N_24713,N_24638);
nor UO_956 (O_956,N_24566,N_24978);
nor UO_957 (O_957,N_24601,N_24679);
and UO_958 (O_958,N_24781,N_24656);
and UO_959 (O_959,N_24642,N_24745);
and UO_960 (O_960,N_24872,N_24661);
xor UO_961 (O_961,N_24576,N_24515);
nand UO_962 (O_962,N_24712,N_24555);
nand UO_963 (O_963,N_24774,N_24857);
nand UO_964 (O_964,N_24955,N_24959);
nor UO_965 (O_965,N_24563,N_24951);
nor UO_966 (O_966,N_24783,N_24881);
nand UO_967 (O_967,N_24845,N_24715);
nor UO_968 (O_968,N_24848,N_24630);
and UO_969 (O_969,N_24994,N_24927);
or UO_970 (O_970,N_24637,N_24897);
nor UO_971 (O_971,N_24738,N_24726);
xnor UO_972 (O_972,N_24687,N_24566);
nand UO_973 (O_973,N_24642,N_24875);
and UO_974 (O_974,N_24691,N_24590);
or UO_975 (O_975,N_24801,N_24834);
nor UO_976 (O_976,N_24788,N_24530);
and UO_977 (O_977,N_24842,N_24547);
and UO_978 (O_978,N_24512,N_24629);
nand UO_979 (O_979,N_24533,N_24712);
nor UO_980 (O_980,N_24892,N_24982);
nor UO_981 (O_981,N_24524,N_24569);
nor UO_982 (O_982,N_24570,N_24739);
and UO_983 (O_983,N_24604,N_24785);
nand UO_984 (O_984,N_24756,N_24708);
or UO_985 (O_985,N_24626,N_24555);
or UO_986 (O_986,N_24851,N_24850);
and UO_987 (O_987,N_24694,N_24671);
and UO_988 (O_988,N_24523,N_24538);
nor UO_989 (O_989,N_24961,N_24987);
and UO_990 (O_990,N_24651,N_24592);
and UO_991 (O_991,N_24817,N_24788);
or UO_992 (O_992,N_24640,N_24962);
or UO_993 (O_993,N_24625,N_24571);
and UO_994 (O_994,N_24562,N_24608);
xor UO_995 (O_995,N_24863,N_24513);
xnor UO_996 (O_996,N_24955,N_24793);
and UO_997 (O_997,N_24669,N_24873);
nand UO_998 (O_998,N_24815,N_24533);
or UO_999 (O_999,N_24887,N_24654);
nor UO_1000 (O_1000,N_24680,N_24901);
or UO_1001 (O_1001,N_24813,N_24709);
or UO_1002 (O_1002,N_24724,N_24654);
nand UO_1003 (O_1003,N_24816,N_24514);
nand UO_1004 (O_1004,N_24555,N_24873);
nand UO_1005 (O_1005,N_24650,N_24907);
nand UO_1006 (O_1006,N_24807,N_24513);
and UO_1007 (O_1007,N_24645,N_24561);
nor UO_1008 (O_1008,N_24908,N_24505);
and UO_1009 (O_1009,N_24874,N_24612);
nor UO_1010 (O_1010,N_24956,N_24749);
and UO_1011 (O_1011,N_24738,N_24589);
nor UO_1012 (O_1012,N_24745,N_24758);
nor UO_1013 (O_1013,N_24653,N_24798);
and UO_1014 (O_1014,N_24558,N_24843);
nand UO_1015 (O_1015,N_24955,N_24721);
nor UO_1016 (O_1016,N_24732,N_24787);
nor UO_1017 (O_1017,N_24825,N_24690);
and UO_1018 (O_1018,N_24924,N_24675);
or UO_1019 (O_1019,N_24771,N_24833);
nor UO_1020 (O_1020,N_24513,N_24631);
nand UO_1021 (O_1021,N_24813,N_24866);
or UO_1022 (O_1022,N_24730,N_24897);
nand UO_1023 (O_1023,N_24826,N_24948);
and UO_1024 (O_1024,N_24957,N_24703);
or UO_1025 (O_1025,N_24544,N_24592);
nor UO_1026 (O_1026,N_24831,N_24617);
or UO_1027 (O_1027,N_24617,N_24686);
nor UO_1028 (O_1028,N_24792,N_24929);
nor UO_1029 (O_1029,N_24863,N_24835);
nor UO_1030 (O_1030,N_24783,N_24907);
nor UO_1031 (O_1031,N_24508,N_24712);
and UO_1032 (O_1032,N_24910,N_24955);
nor UO_1033 (O_1033,N_24936,N_24797);
or UO_1034 (O_1034,N_24658,N_24994);
nand UO_1035 (O_1035,N_24528,N_24553);
and UO_1036 (O_1036,N_24989,N_24782);
nor UO_1037 (O_1037,N_24923,N_24995);
xor UO_1038 (O_1038,N_24527,N_24993);
nand UO_1039 (O_1039,N_24603,N_24846);
and UO_1040 (O_1040,N_24641,N_24638);
and UO_1041 (O_1041,N_24621,N_24996);
nand UO_1042 (O_1042,N_24970,N_24718);
nand UO_1043 (O_1043,N_24712,N_24703);
nor UO_1044 (O_1044,N_24511,N_24553);
nor UO_1045 (O_1045,N_24756,N_24819);
xor UO_1046 (O_1046,N_24735,N_24699);
and UO_1047 (O_1047,N_24851,N_24702);
nand UO_1048 (O_1048,N_24849,N_24556);
or UO_1049 (O_1049,N_24970,N_24980);
and UO_1050 (O_1050,N_24513,N_24878);
xnor UO_1051 (O_1051,N_24528,N_24748);
nand UO_1052 (O_1052,N_24627,N_24796);
xnor UO_1053 (O_1053,N_24714,N_24543);
nor UO_1054 (O_1054,N_24892,N_24739);
nor UO_1055 (O_1055,N_24665,N_24939);
or UO_1056 (O_1056,N_24595,N_24582);
or UO_1057 (O_1057,N_24973,N_24856);
nand UO_1058 (O_1058,N_24910,N_24951);
nor UO_1059 (O_1059,N_24803,N_24917);
nand UO_1060 (O_1060,N_24551,N_24945);
or UO_1061 (O_1061,N_24644,N_24603);
nand UO_1062 (O_1062,N_24857,N_24870);
or UO_1063 (O_1063,N_24713,N_24770);
nand UO_1064 (O_1064,N_24882,N_24808);
nand UO_1065 (O_1065,N_24655,N_24986);
nor UO_1066 (O_1066,N_24515,N_24611);
and UO_1067 (O_1067,N_24829,N_24603);
and UO_1068 (O_1068,N_24517,N_24500);
or UO_1069 (O_1069,N_24681,N_24607);
nand UO_1070 (O_1070,N_24599,N_24571);
or UO_1071 (O_1071,N_24549,N_24975);
or UO_1072 (O_1072,N_24879,N_24784);
and UO_1073 (O_1073,N_24744,N_24697);
and UO_1074 (O_1074,N_24905,N_24582);
and UO_1075 (O_1075,N_24819,N_24797);
xor UO_1076 (O_1076,N_24531,N_24527);
nand UO_1077 (O_1077,N_24756,N_24942);
nor UO_1078 (O_1078,N_24966,N_24544);
and UO_1079 (O_1079,N_24767,N_24745);
nor UO_1080 (O_1080,N_24830,N_24547);
or UO_1081 (O_1081,N_24679,N_24649);
and UO_1082 (O_1082,N_24743,N_24937);
and UO_1083 (O_1083,N_24679,N_24786);
nand UO_1084 (O_1084,N_24542,N_24620);
nor UO_1085 (O_1085,N_24536,N_24739);
or UO_1086 (O_1086,N_24928,N_24713);
and UO_1087 (O_1087,N_24502,N_24651);
or UO_1088 (O_1088,N_24694,N_24627);
or UO_1089 (O_1089,N_24799,N_24536);
nand UO_1090 (O_1090,N_24798,N_24942);
nand UO_1091 (O_1091,N_24960,N_24594);
or UO_1092 (O_1092,N_24776,N_24875);
and UO_1093 (O_1093,N_24743,N_24624);
and UO_1094 (O_1094,N_24692,N_24618);
nand UO_1095 (O_1095,N_24709,N_24531);
nand UO_1096 (O_1096,N_24730,N_24634);
nand UO_1097 (O_1097,N_24811,N_24702);
or UO_1098 (O_1098,N_24504,N_24686);
nand UO_1099 (O_1099,N_24852,N_24610);
and UO_1100 (O_1100,N_24527,N_24890);
nand UO_1101 (O_1101,N_24631,N_24921);
and UO_1102 (O_1102,N_24745,N_24892);
xnor UO_1103 (O_1103,N_24503,N_24589);
nor UO_1104 (O_1104,N_24858,N_24660);
nand UO_1105 (O_1105,N_24705,N_24722);
nand UO_1106 (O_1106,N_24528,N_24604);
nand UO_1107 (O_1107,N_24624,N_24559);
and UO_1108 (O_1108,N_24588,N_24698);
and UO_1109 (O_1109,N_24828,N_24873);
and UO_1110 (O_1110,N_24638,N_24911);
nand UO_1111 (O_1111,N_24761,N_24868);
nor UO_1112 (O_1112,N_24616,N_24798);
or UO_1113 (O_1113,N_24601,N_24672);
nand UO_1114 (O_1114,N_24917,N_24704);
nand UO_1115 (O_1115,N_24509,N_24928);
or UO_1116 (O_1116,N_24915,N_24648);
and UO_1117 (O_1117,N_24747,N_24589);
and UO_1118 (O_1118,N_24890,N_24828);
nand UO_1119 (O_1119,N_24962,N_24761);
and UO_1120 (O_1120,N_24694,N_24656);
nor UO_1121 (O_1121,N_24864,N_24694);
nand UO_1122 (O_1122,N_24688,N_24602);
xnor UO_1123 (O_1123,N_24676,N_24955);
and UO_1124 (O_1124,N_24722,N_24752);
and UO_1125 (O_1125,N_24851,N_24574);
and UO_1126 (O_1126,N_24597,N_24795);
or UO_1127 (O_1127,N_24682,N_24683);
or UO_1128 (O_1128,N_24794,N_24805);
xnor UO_1129 (O_1129,N_24837,N_24764);
or UO_1130 (O_1130,N_24567,N_24895);
nor UO_1131 (O_1131,N_24913,N_24528);
nor UO_1132 (O_1132,N_24580,N_24762);
nor UO_1133 (O_1133,N_24938,N_24689);
nand UO_1134 (O_1134,N_24637,N_24875);
xnor UO_1135 (O_1135,N_24968,N_24753);
nor UO_1136 (O_1136,N_24550,N_24507);
xnor UO_1137 (O_1137,N_24728,N_24843);
or UO_1138 (O_1138,N_24695,N_24958);
nor UO_1139 (O_1139,N_24634,N_24995);
nor UO_1140 (O_1140,N_24986,N_24835);
nand UO_1141 (O_1141,N_24603,N_24879);
and UO_1142 (O_1142,N_24639,N_24773);
xnor UO_1143 (O_1143,N_24654,N_24823);
or UO_1144 (O_1144,N_24578,N_24776);
xor UO_1145 (O_1145,N_24731,N_24663);
and UO_1146 (O_1146,N_24862,N_24639);
nand UO_1147 (O_1147,N_24958,N_24905);
or UO_1148 (O_1148,N_24743,N_24866);
or UO_1149 (O_1149,N_24872,N_24992);
nand UO_1150 (O_1150,N_24708,N_24811);
and UO_1151 (O_1151,N_24970,N_24621);
and UO_1152 (O_1152,N_24861,N_24815);
nand UO_1153 (O_1153,N_24821,N_24657);
nor UO_1154 (O_1154,N_24520,N_24601);
nor UO_1155 (O_1155,N_24688,N_24918);
and UO_1156 (O_1156,N_24602,N_24742);
nand UO_1157 (O_1157,N_24560,N_24792);
nand UO_1158 (O_1158,N_24747,N_24577);
or UO_1159 (O_1159,N_24675,N_24665);
and UO_1160 (O_1160,N_24854,N_24698);
nor UO_1161 (O_1161,N_24952,N_24622);
nand UO_1162 (O_1162,N_24870,N_24711);
or UO_1163 (O_1163,N_24578,N_24881);
xor UO_1164 (O_1164,N_24554,N_24744);
nand UO_1165 (O_1165,N_24888,N_24559);
nand UO_1166 (O_1166,N_24894,N_24646);
nand UO_1167 (O_1167,N_24779,N_24760);
nand UO_1168 (O_1168,N_24996,N_24615);
or UO_1169 (O_1169,N_24631,N_24819);
nand UO_1170 (O_1170,N_24504,N_24701);
or UO_1171 (O_1171,N_24937,N_24509);
nand UO_1172 (O_1172,N_24859,N_24818);
nor UO_1173 (O_1173,N_24982,N_24703);
nor UO_1174 (O_1174,N_24773,N_24504);
nor UO_1175 (O_1175,N_24644,N_24560);
and UO_1176 (O_1176,N_24758,N_24702);
xnor UO_1177 (O_1177,N_24661,N_24910);
nor UO_1178 (O_1178,N_24529,N_24899);
or UO_1179 (O_1179,N_24939,N_24777);
nand UO_1180 (O_1180,N_24823,N_24611);
xnor UO_1181 (O_1181,N_24507,N_24761);
or UO_1182 (O_1182,N_24971,N_24786);
and UO_1183 (O_1183,N_24804,N_24765);
and UO_1184 (O_1184,N_24536,N_24566);
nand UO_1185 (O_1185,N_24605,N_24628);
nand UO_1186 (O_1186,N_24797,N_24986);
nor UO_1187 (O_1187,N_24896,N_24613);
nand UO_1188 (O_1188,N_24887,N_24889);
nor UO_1189 (O_1189,N_24899,N_24922);
nand UO_1190 (O_1190,N_24649,N_24948);
or UO_1191 (O_1191,N_24841,N_24636);
nor UO_1192 (O_1192,N_24986,N_24963);
nand UO_1193 (O_1193,N_24791,N_24740);
nor UO_1194 (O_1194,N_24613,N_24526);
nor UO_1195 (O_1195,N_24806,N_24833);
and UO_1196 (O_1196,N_24645,N_24954);
nor UO_1197 (O_1197,N_24666,N_24534);
nand UO_1198 (O_1198,N_24546,N_24623);
xor UO_1199 (O_1199,N_24905,N_24821);
and UO_1200 (O_1200,N_24889,N_24690);
or UO_1201 (O_1201,N_24562,N_24814);
and UO_1202 (O_1202,N_24977,N_24925);
or UO_1203 (O_1203,N_24886,N_24531);
and UO_1204 (O_1204,N_24638,N_24511);
or UO_1205 (O_1205,N_24630,N_24795);
nand UO_1206 (O_1206,N_24681,N_24888);
nand UO_1207 (O_1207,N_24791,N_24646);
and UO_1208 (O_1208,N_24825,N_24904);
nor UO_1209 (O_1209,N_24686,N_24673);
nor UO_1210 (O_1210,N_24814,N_24574);
xor UO_1211 (O_1211,N_24751,N_24771);
nor UO_1212 (O_1212,N_24597,N_24821);
or UO_1213 (O_1213,N_24924,N_24954);
and UO_1214 (O_1214,N_24699,N_24689);
nor UO_1215 (O_1215,N_24666,N_24847);
or UO_1216 (O_1216,N_24930,N_24942);
or UO_1217 (O_1217,N_24904,N_24644);
or UO_1218 (O_1218,N_24720,N_24792);
nor UO_1219 (O_1219,N_24662,N_24990);
and UO_1220 (O_1220,N_24895,N_24764);
nand UO_1221 (O_1221,N_24801,N_24728);
nor UO_1222 (O_1222,N_24977,N_24516);
or UO_1223 (O_1223,N_24813,N_24695);
and UO_1224 (O_1224,N_24977,N_24605);
nor UO_1225 (O_1225,N_24516,N_24781);
or UO_1226 (O_1226,N_24588,N_24975);
nand UO_1227 (O_1227,N_24780,N_24584);
nor UO_1228 (O_1228,N_24917,N_24500);
and UO_1229 (O_1229,N_24752,N_24874);
xnor UO_1230 (O_1230,N_24801,N_24803);
and UO_1231 (O_1231,N_24578,N_24599);
nand UO_1232 (O_1232,N_24883,N_24850);
nor UO_1233 (O_1233,N_24820,N_24768);
or UO_1234 (O_1234,N_24583,N_24805);
nor UO_1235 (O_1235,N_24938,N_24515);
nor UO_1236 (O_1236,N_24811,N_24779);
nand UO_1237 (O_1237,N_24763,N_24510);
xor UO_1238 (O_1238,N_24993,N_24513);
nand UO_1239 (O_1239,N_24657,N_24814);
xnor UO_1240 (O_1240,N_24503,N_24728);
nand UO_1241 (O_1241,N_24743,N_24949);
and UO_1242 (O_1242,N_24845,N_24835);
and UO_1243 (O_1243,N_24655,N_24546);
or UO_1244 (O_1244,N_24737,N_24805);
or UO_1245 (O_1245,N_24961,N_24752);
or UO_1246 (O_1246,N_24904,N_24877);
nor UO_1247 (O_1247,N_24992,N_24863);
nor UO_1248 (O_1248,N_24608,N_24719);
nand UO_1249 (O_1249,N_24864,N_24679);
xor UO_1250 (O_1250,N_24880,N_24679);
nor UO_1251 (O_1251,N_24790,N_24660);
and UO_1252 (O_1252,N_24922,N_24956);
xnor UO_1253 (O_1253,N_24807,N_24797);
and UO_1254 (O_1254,N_24628,N_24951);
and UO_1255 (O_1255,N_24557,N_24819);
nand UO_1256 (O_1256,N_24549,N_24711);
nand UO_1257 (O_1257,N_24889,N_24519);
and UO_1258 (O_1258,N_24892,N_24936);
or UO_1259 (O_1259,N_24556,N_24937);
or UO_1260 (O_1260,N_24638,N_24719);
nor UO_1261 (O_1261,N_24675,N_24624);
or UO_1262 (O_1262,N_24651,N_24540);
nor UO_1263 (O_1263,N_24721,N_24930);
and UO_1264 (O_1264,N_24818,N_24517);
nor UO_1265 (O_1265,N_24631,N_24604);
nor UO_1266 (O_1266,N_24712,N_24784);
xor UO_1267 (O_1267,N_24617,N_24624);
xor UO_1268 (O_1268,N_24826,N_24973);
nor UO_1269 (O_1269,N_24726,N_24980);
nand UO_1270 (O_1270,N_24750,N_24721);
or UO_1271 (O_1271,N_24740,N_24859);
xnor UO_1272 (O_1272,N_24957,N_24822);
or UO_1273 (O_1273,N_24691,N_24881);
nand UO_1274 (O_1274,N_24818,N_24647);
or UO_1275 (O_1275,N_24946,N_24662);
or UO_1276 (O_1276,N_24672,N_24506);
or UO_1277 (O_1277,N_24887,N_24888);
nor UO_1278 (O_1278,N_24830,N_24777);
nor UO_1279 (O_1279,N_24968,N_24735);
nand UO_1280 (O_1280,N_24730,N_24633);
xor UO_1281 (O_1281,N_24609,N_24540);
or UO_1282 (O_1282,N_24660,N_24543);
and UO_1283 (O_1283,N_24762,N_24922);
and UO_1284 (O_1284,N_24720,N_24926);
nor UO_1285 (O_1285,N_24679,N_24769);
and UO_1286 (O_1286,N_24624,N_24696);
and UO_1287 (O_1287,N_24592,N_24607);
and UO_1288 (O_1288,N_24724,N_24926);
xor UO_1289 (O_1289,N_24614,N_24863);
nand UO_1290 (O_1290,N_24994,N_24525);
nor UO_1291 (O_1291,N_24744,N_24746);
xnor UO_1292 (O_1292,N_24995,N_24843);
and UO_1293 (O_1293,N_24802,N_24636);
or UO_1294 (O_1294,N_24697,N_24838);
or UO_1295 (O_1295,N_24758,N_24574);
and UO_1296 (O_1296,N_24618,N_24702);
nor UO_1297 (O_1297,N_24610,N_24886);
or UO_1298 (O_1298,N_24640,N_24502);
xor UO_1299 (O_1299,N_24996,N_24799);
nor UO_1300 (O_1300,N_24915,N_24738);
and UO_1301 (O_1301,N_24652,N_24772);
and UO_1302 (O_1302,N_24863,N_24696);
or UO_1303 (O_1303,N_24658,N_24527);
nand UO_1304 (O_1304,N_24882,N_24858);
xor UO_1305 (O_1305,N_24795,N_24863);
xor UO_1306 (O_1306,N_24987,N_24645);
and UO_1307 (O_1307,N_24800,N_24618);
nand UO_1308 (O_1308,N_24546,N_24612);
nand UO_1309 (O_1309,N_24737,N_24617);
nor UO_1310 (O_1310,N_24989,N_24808);
nor UO_1311 (O_1311,N_24860,N_24807);
nor UO_1312 (O_1312,N_24501,N_24650);
and UO_1313 (O_1313,N_24714,N_24641);
nand UO_1314 (O_1314,N_24850,N_24760);
nor UO_1315 (O_1315,N_24802,N_24885);
nor UO_1316 (O_1316,N_24854,N_24760);
and UO_1317 (O_1317,N_24883,N_24503);
or UO_1318 (O_1318,N_24755,N_24705);
or UO_1319 (O_1319,N_24587,N_24888);
nand UO_1320 (O_1320,N_24976,N_24948);
xnor UO_1321 (O_1321,N_24619,N_24925);
nand UO_1322 (O_1322,N_24973,N_24577);
nand UO_1323 (O_1323,N_24709,N_24599);
or UO_1324 (O_1324,N_24860,N_24717);
nor UO_1325 (O_1325,N_24546,N_24695);
xnor UO_1326 (O_1326,N_24661,N_24869);
and UO_1327 (O_1327,N_24950,N_24994);
or UO_1328 (O_1328,N_24614,N_24763);
nor UO_1329 (O_1329,N_24601,N_24801);
nor UO_1330 (O_1330,N_24876,N_24919);
or UO_1331 (O_1331,N_24940,N_24607);
nor UO_1332 (O_1332,N_24971,N_24648);
and UO_1333 (O_1333,N_24610,N_24863);
nor UO_1334 (O_1334,N_24871,N_24731);
and UO_1335 (O_1335,N_24533,N_24854);
xor UO_1336 (O_1336,N_24635,N_24743);
nor UO_1337 (O_1337,N_24903,N_24765);
and UO_1338 (O_1338,N_24894,N_24661);
xor UO_1339 (O_1339,N_24557,N_24622);
and UO_1340 (O_1340,N_24910,N_24861);
xnor UO_1341 (O_1341,N_24605,N_24725);
nand UO_1342 (O_1342,N_24901,N_24857);
or UO_1343 (O_1343,N_24918,N_24705);
xnor UO_1344 (O_1344,N_24772,N_24669);
or UO_1345 (O_1345,N_24779,N_24632);
nand UO_1346 (O_1346,N_24638,N_24501);
and UO_1347 (O_1347,N_24531,N_24569);
nand UO_1348 (O_1348,N_24985,N_24793);
and UO_1349 (O_1349,N_24852,N_24832);
and UO_1350 (O_1350,N_24648,N_24509);
xnor UO_1351 (O_1351,N_24738,N_24922);
nor UO_1352 (O_1352,N_24975,N_24768);
or UO_1353 (O_1353,N_24686,N_24606);
nand UO_1354 (O_1354,N_24834,N_24813);
and UO_1355 (O_1355,N_24994,N_24899);
nor UO_1356 (O_1356,N_24760,N_24673);
nand UO_1357 (O_1357,N_24757,N_24702);
and UO_1358 (O_1358,N_24531,N_24796);
nor UO_1359 (O_1359,N_24609,N_24636);
or UO_1360 (O_1360,N_24787,N_24797);
nand UO_1361 (O_1361,N_24683,N_24982);
and UO_1362 (O_1362,N_24714,N_24836);
nand UO_1363 (O_1363,N_24643,N_24920);
or UO_1364 (O_1364,N_24833,N_24620);
nand UO_1365 (O_1365,N_24878,N_24736);
or UO_1366 (O_1366,N_24829,N_24652);
and UO_1367 (O_1367,N_24700,N_24549);
and UO_1368 (O_1368,N_24908,N_24763);
nor UO_1369 (O_1369,N_24884,N_24634);
nand UO_1370 (O_1370,N_24521,N_24801);
or UO_1371 (O_1371,N_24609,N_24758);
nor UO_1372 (O_1372,N_24670,N_24863);
and UO_1373 (O_1373,N_24865,N_24609);
and UO_1374 (O_1374,N_24667,N_24566);
nor UO_1375 (O_1375,N_24742,N_24989);
and UO_1376 (O_1376,N_24546,N_24967);
nand UO_1377 (O_1377,N_24729,N_24613);
nand UO_1378 (O_1378,N_24593,N_24671);
and UO_1379 (O_1379,N_24558,N_24876);
nand UO_1380 (O_1380,N_24579,N_24715);
or UO_1381 (O_1381,N_24891,N_24590);
nand UO_1382 (O_1382,N_24807,N_24572);
xnor UO_1383 (O_1383,N_24500,N_24846);
nor UO_1384 (O_1384,N_24847,N_24572);
or UO_1385 (O_1385,N_24819,N_24755);
and UO_1386 (O_1386,N_24988,N_24644);
xor UO_1387 (O_1387,N_24521,N_24677);
or UO_1388 (O_1388,N_24678,N_24519);
or UO_1389 (O_1389,N_24701,N_24938);
nand UO_1390 (O_1390,N_24932,N_24999);
or UO_1391 (O_1391,N_24695,N_24746);
nor UO_1392 (O_1392,N_24656,N_24648);
and UO_1393 (O_1393,N_24698,N_24937);
nand UO_1394 (O_1394,N_24954,N_24674);
and UO_1395 (O_1395,N_24672,N_24675);
nor UO_1396 (O_1396,N_24578,N_24835);
nor UO_1397 (O_1397,N_24572,N_24830);
xnor UO_1398 (O_1398,N_24697,N_24741);
and UO_1399 (O_1399,N_24514,N_24970);
or UO_1400 (O_1400,N_24581,N_24770);
and UO_1401 (O_1401,N_24577,N_24684);
and UO_1402 (O_1402,N_24962,N_24908);
or UO_1403 (O_1403,N_24737,N_24866);
and UO_1404 (O_1404,N_24955,N_24799);
and UO_1405 (O_1405,N_24596,N_24897);
or UO_1406 (O_1406,N_24674,N_24829);
xnor UO_1407 (O_1407,N_24592,N_24582);
and UO_1408 (O_1408,N_24930,N_24979);
or UO_1409 (O_1409,N_24965,N_24944);
or UO_1410 (O_1410,N_24708,N_24591);
xnor UO_1411 (O_1411,N_24833,N_24615);
and UO_1412 (O_1412,N_24920,N_24861);
and UO_1413 (O_1413,N_24734,N_24577);
xnor UO_1414 (O_1414,N_24779,N_24534);
and UO_1415 (O_1415,N_24984,N_24626);
or UO_1416 (O_1416,N_24719,N_24515);
nand UO_1417 (O_1417,N_24637,N_24543);
or UO_1418 (O_1418,N_24528,N_24721);
or UO_1419 (O_1419,N_24736,N_24800);
xor UO_1420 (O_1420,N_24690,N_24523);
nand UO_1421 (O_1421,N_24997,N_24706);
or UO_1422 (O_1422,N_24976,N_24993);
nor UO_1423 (O_1423,N_24826,N_24547);
nand UO_1424 (O_1424,N_24716,N_24518);
nor UO_1425 (O_1425,N_24514,N_24841);
xor UO_1426 (O_1426,N_24636,N_24519);
nor UO_1427 (O_1427,N_24653,N_24973);
or UO_1428 (O_1428,N_24667,N_24867);
or UO_1429 (O_1429,N_24911,N_24777);
xor UO_1430 (O_1430,N_24962,N_24982);
and UO_1431 (O_1431,N_24710,N_24803);
and UO_1432 (O_1432,N_24614,N_24941);
or UO_1433 (O_1433,N_24730,N_24590);
xor UO_1434 (O_1434,N_24751,N_24937);
and UO_1435 (O_1435,N_24850,N_24785);
and UO_1436 (O_1436,N_24919,N_24943);
nand UO_1437 (O_1437,N_24646,N_24761);
and UO_1438 (O_1438,N_24990,N_24727);
xor UO_1439 (O_1439,N_24841,N_24977);
nand UO_1440 (O_1440,N_24808,N_24748);
xnor UO_1441 (O_1441,N_24654,N_24639);
nor UO_1442 (O_1442,N_24865,N_24720);
or UO_1443 (O_1443,N_24569,N_24952);
nand UO_1444 (O_1444,N_24987,N_24960);
nor UO_1445 (O_1445,N_24637,N_24764);
nand UO_1446 (O_1446,N_24576,N_24605);
nor UO_1447 (O_1447,N_24550,N_24861);
nand UO_1448 (O_1448,N_24588,N_24864);
nand UO_1449 (O_1449,N_24621,N_24504);
and UO_1450 (O_1450,N_24584,N_24661);
nand UO_1451 (O_1451,N_24678,N_24780);
nand UO_1452 (O_1452,N_24892,N_24901);
xnor UO_1453 (O_1453,N_24853,N_24986);
nor UO_1454 (O_1454,N_24586,N_24741);
or UO_1455 (O_1455,N_24595,N_24868);
nor UO_1456 (O_1456,N_24682,N_24757);
nand UO_1457 (O_1457,N_24641,N_24612);
or UO_1458 (O_1458,N_24939,N_24776);
or UO_1459 (O_1459,N_24966,N_24525);
nand UO_1460 (O_1460,N_24633,N_24753);
nand UO_1461 (O_1461,N_24734,N_24694);
nor UO_1462 (O_1462,N_24963,N_24566);
nor UO_1463 (O_1463,N_24760,N_24928);
or UO_1464 (O_1464,N_24515,N_24562);
nand UO_1465 (O_1465,N_24880,N_24678);
and UO_1466 (O_1466,N_24836,N_24798);
nor UO_1467 (O_1467,N_24536,N_24749);
and UO_1468 (O_1468,N_24661,N_24966);
and UO_1469 (O_1469,N_24824,N_24954);
and UO_1470 (O_1470,N_24574,N_24647);
or UO_1471 (O_1471,N_24676,N_24600);
nand UO_1472 (O_1472,N_24614,N_24716);
nor UO_1473 (O_1473,N_24896,N_24543);
nand UO_1474 (O_1474,N_24598,N_24664);
or UO_1475 (O_1475,N_24608,N_24789);
or UO_1476 (O_1476,N_24750,N_24615);
and UO_1477 (O_1477,N_24659,N_24809);
xor UO_1478 (O_1478,N_24867,N_24638);
or UO_1479 (O_1479,N_24999,N_24760);
xor UO_1480 (O_1480,N_24882,N_24657);
nand UO_1481 (O_1481,N_24621,N_24907);
or UO_1482 (O_1482,N_24980,N_24741);
nand UO_1483 (O_1483,N_24987,N_24586);
nand UO_1484 (O_1484,N_24872,N_24806);
nor UO_1485 (O_1485,N_24691,N_24843);
or UO_1486 (O_1486,N_24628,N_24631);
nand UO_1487 (O_1487,N_24542,N_24793);
nor UO_1488 (O_1488,N_24853,N_24770);
and UO_1489 (O_1489,N_24846,N_24942);
xor UO_1490 (O_1490,N_24994,N_24834);
and UO_1491 (O_1491,N_24650,N_24869);
and UO_1492 (O_1492,N_24718,N_24650);
and UO_1493 (O_1493,N_24748,N_24599);
or UO_1494 (O_1494,N_24824,N_24765);
xor UO_1495 (O_1495,N_24653,N_24638);
or UO_1496 (O_1496,N_24991,N_24724);
nand UO_1497 (O_1497,N_24771,N_24949);
nor UO_1498 (O_1498,N_24736,N_24850);
and UO_1499 (O_1499,N_24691,N_24746);
and UO_1500 (O_1500,N_24982,N_24816);
nand UO_1501 (O_1501,N_24935,N_24667);
and UO_1502 (O_1502,N_24532,N_24759);
nand UO_1503 (O_1503,N_24898,N_24749);
and UO_1504 (O_1504,N_24640,N_24596);
nor UO_1505 (O_1505,N_24831,N_24505);
and UO_1506 (O_1506,N_24588,N_24736);
xor UO_1507 (O_1507,N_24535,N_24888);
nor UO_1508 (O_1508,N_24785,N_24541);
or UO_1509 (O_1509,N_24991,N_24865);
nand UO_1510 (O_1510,N_24667,N_24978);
or UO_1511 (O_1511,N_24585,N_24567);
nor UO_1512 (O_1512,N_24591,N_24579);
xor UO_1513 (O_1513,N_24606,N_24945);
nor UO_1514 (O_1514,N_24523,N_24603);
nand UO_1515 (O_1515,N_24566,N_24915);
nand UO_1516 (O_1516,N_24865,N_24955);
or UO_1517 (O_1517,N_24910,N_24689);
xnor UO_1518 (O_1518,N_24685,N_24838);
nand UO_1519 (O_1519,N_24843,N_24553);
and UO_1520 (O_1520,N_24757,N_24735);
and UO_1521 (O_1521,N_24948,N_24995);
nor UO_1522 (O_1522,N_24584,N_24695);
nor UO_1523 (O_1523,N_24770,N_24925);
and UO_1524 (O_1524,N_24658,N_24600);
nor UO_1525 (O_1525,N_24820,N_24956);
or UO_1526 (O_1526,N_24585,N_24703);
or UO_1527 (O_1527,N_24754,N_24551);
xor UO_1528 (O_1528,N_24584,N_24617);
and UO_1529 (O_1529,N_24892,N_24579);
nand UO_1530 (O_1530,N_24695,N_24873);
nand UO_1531 (O_1531,N_24856,N_24861);
and UO_1532 (O_1532,N_24813,N_24920);
and UO_1533 (O_1533,N_24755,N_24551);
nand UO_1534 (O_1534,N_24902,N_24881);
nor UO_1535 (O_1535,N_24844,N_24524);
and UO_1536 (O_1536,N_24775,N_24820);
or UO_1537 (O_1537,N_24986,N_24957);
and UO_1538 (O_1538,N_24636,N_24669);
nor UO_1539 (O_1539,N_24551,N_24717);
nand UO_1540 (O_1540,N_24597,N_24848);
or UO_1541 (O_1541,N_24520,N_24877);
or UO_1542 (O_1542,N_24533,N_24762);
or UO_1543 (O_1543,N_24986,N_24553);
nor UO_1544 (O_1544,N_24716,N_24639);
or UO_1545 (O_1545,N_24899,N_24610);
or UO_1546 (O_1546,N_24923,N_24582);
xor UO_1547 (O_1547,N_24937,N_24744);
nand UO_1548 (O_1548,N_24841,N_24854);
nand UO_1549 (O_1549,N_24533,N_24748);
nand UO_1550 (O_1550,N_24877,N_24628);
and UO_1551 (O_1551,N_24581,N_24713);
xor UO_1552 (O_1552,N_24748,N_24537);
or UO_1553 (O_1553,N_24758,N_24909);
and UO_1554 (O_1554,N_24830,N_24967);
nand UO_1555 (O_1555,N_24885,N_24792);
or UO_1556 (O_1556,N_24718,N_24980);
nor UO_1557 (O_1557,N_24925,N_24615);
and UO_1558 (O_1558,N_24716,N_24983);
nand UO_1559 (O_1559,N_24582,N_24783);
or UO_1560 (O_1560,N_24996,N_24586);
or UO_1561 (O_1561,N_24678,N_24726);
and UO_1562 (O_1562,N_24787,N_24996);
and UO_1563 (O_1563,N_24911,N_24816);
and UO_1564 (O_1564,N_24908,N_24568);
and UO_1565 (O_1565,N_24721,N_24864);
nand UO_1566 (O_1566,N_24838,N_24899);
and UO_1567 (O_1567,N_24589,N_24897);
nor UO_1568 (O_1568,N_24758,N_24975);
or UO_1569 (O_1569,N_24845,N_24629);
nand UO_1570 (O_1570,N_24702,N_24937);
and UO_1571 (O_1571,N_24879,N_24686);
or UO_1572 (O_1572,N_24524,N_24994);
or UO_1573 (O_1573,N_24927,N_24546);
and UO_1574 (O_1574,N_24532,N_24693);
nor UO_1575 (O_1575,N_24747,N_24831);
and UO_1576 (O_1576,N_24738,N_24659);
and UO_1577 (O_1577,N_24723,N_24762);
nand UO_1578 (O_1578,N_24596,N_24968);
and UO_1579 (O_1579,N_24891,N_24576);
nand UO_1580 (O_1580,N_24938,N_24571);
or UO_1581 (O_1581,N_24818,N_24576);
nor UO_1582 (O_1582,N_24963,N_24845);
or UO_1583 (O_1583,N_24844,N_24722);
nand UO_1584 (O_1584,N_24531,N_24703);
nand UO_1585 (O_1585,N_24980,N_24830);
or UO_1586 (O_1586,N_24745,N_24612);
nand UO_1587 (O_1587,N_24854,N_24572);
and UO_1588 (O_1588,N_24544,N_24894);
nand UO_1589 (O_1589,N_24532,N_24773);
or UO_1590 (O_1590,N_24671,N_24771);
or UO_1591 (O_1591,N_24734,N_24533);
nand UO_1592 (O_1592,N_24638,N_24878);
nand UO_1593 (O_1593,N_24677,N_24924);
and UO_1594 (O_1594,N_24992,N_24683);
and UO_1595 (O_1595,N_24873,N_24975);
nor UO_1596 (O_1596,N_24826,N_24959);
or UO_1597 (O_1597,N_24776,N_24617);
nand UO_1598 (O_1598,N_24935,N_24671);
nand UO_1599 (O_1599,N_24759,N_24619);
and UO_1600 (O_1600,N_24600,N_24625);
nor UO_1601 (O_1601,N_24965,N_24967);
or UO_1602 (O_1602,N_24956,N_24904);
nand UO_1603 (O_1603,N_24546,N_24662);
nand UO_1604 (O_1604,N_24742,N_24815);
xnor UO_1605 (O_1605,N_24830,N_24981);
nand UO_1606 (O_1606,N_24747,N_24715);
nand UO_1607 (O_1607,N_24983,N_24708);
nand UO_1608 (O_1608,N_24918,N_24535);
and UO_1609 (O_1609,N_24542,N_24667);
nand UO_1610 (O_1610,N_24777,N_24633);
xnor UO_1611 (O_1611,N_24611,N_24551);
nand UO_1612 (O_1612,N_24969,N_24712);
xor UO_1613 (O_1613,N_24774,N_24734);
or UO_1614 (O_1614,N_24996,N_24899);
or UO_1615 (O_1615,N_24871,N_24736);
nor UO_1616 (O_1616,N_24563,N_24721);
nand UO_1617 (O_1617,N_24788,N_24857);
or UO_1618 (O_1618,N_24787,N_24970);
xnor UO_1619 (O_1619,N_24879,N_24920);
and UO_1620 (O_1620,N_24591,N_24804);
nor UO_1621 (O_1621,N_24686,N_24948);
or UO_1622 (O_1622,N_24667,N_24713);
and UO_1623 (O_1623,N_24995,N_24572);
or UO_1624 (O_1624,N_24702,N_24513);
or UO_1625 (O_1625,N_24777,N_24601);
or UO_1626 (O_1626,N_24618,N_24851);
and UO_1627 (O_1627,N_24511,N_24862);
and UO_1628 (O_1628,N_24630,N_24685);
or UO_1629 (O_1629,N_24913,N_24690);
nand UO_1630 (O_1630,N_24795,N_24547);
or UO_1631 (O_1631,N_24691,N_24752);
or UO_1632 (O_1632,N_24919,N_24552);
and UO_1633 (O_1633,N_24910,N_24932);
and UO_1634 (O_1634,N_24819,N_24837);
or UO_1635 (O_1635,N_24758,N_24831);
nor UO_1636 (O_1636,N_24572,N_24703);
or UO_1637 (O_1637,N_24712,N_24717);
and UO_1638 (O_1638,N_24612,N_24632);
nor UO_1639 (O_1639,N_24541,N_24858);
nor UO_1640 (O_1640,N_24589,N_24775);
or UO_1641 (O_1641,N_24541,N_24688);
nor UO_1642 (O_1642,N_24716,N_24646);
and UO_1643 (O_1643,N_24762,N_24737);
nor UO_1644 (O_1644,N_24967,N_24730);
and UO_1645 (O_1645,N_24877,N_24789);
nand UO_1646 (O_1646,N_24690,N_24524);
nand UO_1647 (O_1647,N_24587,N_24882);
and UO_1648 (O_1648,N_24771,N_24945);
nand UO_1649 (O_1649,N_24941,N_24660);
nand UO_1650 (O_1650,N_24861,N_24958);
nor UO_1651 (O_1651,N_24532,N_24819);
or UO_1652 (O_1652,N_24819,N_24556);
or UO_1653 (O_1653,N_24565,N_24941);
and UO_1654 (O_1654,N_24871,N_24585);
nor UO_1655 (O_1655,N_24764,N_24782);
nor UO_1656 (O_1656,N_24769,N_24554);
and UO_1657 (O_1657,N_24775,N_24809);
nor UO_1658 (O_1658,N_24607,N_24814);
nand UO_1659 (O_1659,N_24622,N_24994);
nand UO_1660 (O_1660,N_24998,N_24928);
nor UO_1661 (O_1661,N_24620,N_24917);
nor UO_1662 (O_1662,N_24985,N_24878);
and UO_1663 (O_1663,N_24978,N_24781);
xor UO_1664 (O_1664,N_24826,N_24751);
xnor UO_1665 (O_1665,N_24542,N_24735);
or UO_1666 (O_1666,N_24515,N_24554);
or UO_1667 (O_1667,N_24853,N_24586);
or UO_1668 (O_1668,N_24710,N_24998);
and UO_1669 (O_1669,N_24600,N_24716);
nor UO_1670 (O_1670,N_24904,N_24744);
or UO_1671 (O_1671,N_24940,N_24546);
and UO_1672 (O_1672,N_24687,N_24792);
or UO_1673 (O_1673,N_24552,N_24683);
xor UO_1674 (O_1674,N_24602,N_24999);
or UO_1675 (O_1675,N_24671,N_24998);
or UO_1676 (O_1676,N_24906,N_24531);
nor UO_1677 (O_1677,N_24648,N_24820);
nand UO_1678 (O_1678,N_24618,N_24823);
and UO_1679 (O_1679,N_24766,N_24576);
nand UO_1680 (O_1680,N_24569,N_24797);
nand UO_1681 (O_1681,N_24574,N_24505);
nand UO_1682 (O_1682,N_24644,N_24791);
xnor UO_1683 (O_1683,N_24739,N_24825);
xor UO_1684 (O_1684,N_24976,N_24741);
nor UO_1685 (O_1685,N_24908,N_24795);
nor UO_1686 (O_1686,N_24634,N_24973);
and UO_1687 (O_1687,N_24681,N_24975);
and UO_1688 (O_1688,N_24908,N_24766);
and UO_1689 (O_1689,N_24982,N_24671);
xor UO_1690 (O_1690,N_24697,N_24626);
nor UO_1691 (O_1691,N_24848,N_24688);
nand UO_1692 (O_1692,N_24754,N_24600);
nand UO_1693 (O_1693,N_24538,N_24600);
nand UO_1694 (O_1694,N_24693,N_24642);
nand UO_1695 (O_1695,N_24780,N_24827);
and UO_1696 (O_1696,N_24916,N_24871);
or UO_1697 (O_1697,N_24799,N_24818);
nand UO_1698 (O_1698,N_24539,N_24540);
nor UO_1699 (O_1699,N_24764,N_24564);
or UO_1700 (O_1700,N_24622,N_24967);
nand UO_1701 (O_1701,N_24911,N_24966);
or UO_1702 (O_1702,N_24858,N_24923);
and UO_1703 (O_1703,N_24719,N_24592);
nor UO_1704 (O_1704,N_24793,N_24678);
and UO_1705 (O_1705,N_24866,N_24984);
and UO_1706 (O_1706,N_24724,N_24835);
or UO_1707 (O_1707,N_24604,N_24853);
and UO_1708 (O_1708,N_24543,N_24893);
and UO_1709 (O_1709,N_24697,N_24603);
or UO_1710 (O_1710,N_24525,N_24536);
or UO_1711 (O_1711,N_24835,N_24725);
and UO_1712 (O_1712,N_24754,N_24596);
or UO_1713 (O_1713,N_24778,N_24824);
nand UO_1714 (O_1714,N_24573,N_24847);
or UO_1715 (O_1715,N_24815,N_24538);
or UO_1716 (O_1716,N_24764,N_24933);
and UO_1717 (O_1717,N_24850,N_24669);
nand UO_1718 (O_1718,N_24670,N_24855);
and UO_1719 (O_1719,N_24826,N_24872);
or UO_1720 (O_1720,N_24966,N_24716);
or UO_1721 (O_1721,N_24864,N_24595);
and UO_1722 (O_1722,N_24936,N_24592);
nor UO_1723 (O_1723,N_24954,N_24876);
xnor UO_1724 (O_1724,N_24646,N_24803);
nand UO_1725 (O_1725,N_24826,N_24500);
or UO_1726 (O_1726,N_24786,N_24723);
nand UO_1727 (O_1727,N_24891,N_24780);
nand UO_1728 (O_1728,N_24685,N_24641);
nand UO_1729 (O_1729,N_24522,N_24571);
nor UO_1730 (O_1730,N_24684,N_24665);
or UO_1731 (O_1731,N_24960,N_24923);
xor UO_1732 (O_1732,N_24618,N_24591);
and UO_1733 (O_1733,N_24518,N_24568);
or UO_1734 (O_1734,N_24616,N_24787);
nor UO_1735 (O_1735,N_24913,N_24749);
or UO_1736 (O_1736,N_24876,N_24844);
and UO_1737 (O_1737,N_24562,N_24894);
and UO_1738 (O_1738,N_24712,N_24777);
or UO_1739 (O_1739,N_24859,N_24927);
and UO_1740 (O_1740,N_24563,N_24871);
or UO_1741 (O_1741,N_24623,N_24732);
and UO_1742 (O_1742,N_24562,N_24950);
nand UO_1743 (O_1743,N_24747,N_24630);
or UO_1744 (O_1744,N_24619,N_24882);
and UO_1745 (O_1745,N_24947,N_24501);
nor UO_1746 (O_1746,N_24956,N_24989);
or UO_1747 (O_1747,N_24614,N_24675);
nor UO_1748 (O_1748,N_24792,N_24703);
xnor UO_1749 (O_1749,N_24600,N_24768);
or UO_1750 (O_1750,N_24525,N_24861);
xnor UO_1751 (O_1751,N_24777,N_24829);
or UO_1752 (O_1752,N_24531,N_24662);
nand UO_1753 (O_1753,N_24944,N_24846);
nand UO_1754 (O_1754,N_24692,N_24737);
or UO_1755 (O_1755,N_24580,N_24569);
nand UO_1756 (O_1756,N_24891,N_24535);
nor UO_1757 (O_1757,N_24834,N_24875);
nand UO_1758 (O_1758,N_24770,N_24540);
or UO_1759 (O_1759,N_24592,N_24835);
or UO_1760 (O_1760,N_24725,N_24772);
and UO_1761 (O_1761,N_24519,N_24606);
or UO_1762 (O_1762,N_24594,N_24599);
nor UO_1763 (O_1763,N_24587,N_24962);
xnor UO_1764 (O_1764,N_24722,N_24871);
nor UO_1765 (O_1765,N_24521,N_24989);
nor UO_1766 (O_1766,N_24779,N_24511);
and UO_1767 (O_1767,N_24941,N_24601);
and UO_1768 (O_1768,N_24536,N_24596);
and UO_1769 (O_1769,N_24889,N_24681);
nor UO_1770 (O_1770,N_24996,N_24596);
and UO_1771 (O_1771,N_24941,N_24847);
nand UO_1772 (O_1772,N_24897,N_24549);
nand UO_1773 (O_1773,N_24725,N_24990);
nor UO_1774 (O_1774,N_24931,N_24672);
nor UO_1775 (O_1775,N_24870,N_24682);
and UO_1776 (O_1776,N_24896,N_24682);
or UO_1777 (O_1777,N_24811,N_24901);
nor UO_1778 (O_1778,N_24622,N_24610);
nor UO_1779 (O_1779,N_24868,N_24654);
nor UO_1780 (O_1780,N_24680,N_24806);
nand UO_1781 (O_1781,N_24742,N_24944);
nor UO_1782 (O_1782,N_24578,N_24670);
or UO_1783 (O_1783,N_24826,N_24616);
nand UO_1784 (O_1784,N_24757,N_24837);
nor UO_1785 (O_1785,N_24894,N_24884);
xnor UO_1786 (O_1786,N_24613,N_24638);
nand UO_1787 (O_1787,N_24885,N_24810);
and UO_1788 (O_1788,N_24745,N_24553);
or UO_1789 (O_1789,N_24673,N_24620);
or UO_1790 (O_1790,N_24848,N_24588);
nand UO_1791 (O_1791,N_24780,N_24831);
and UO_1792 (O_1792,N_24889,N_24902);
nor UO_1793 (O_1793,N_24945,N_24570);
and UO_1794 (O_1794,N_24814,N_24521);
and UO_1795 (O_1795,N_24728,N_24686);
or UO_1796 (O_1796,N_24737,N_24952);
nor UO_1797 (O_1797,N_24951,N_24915);
xnor UO_1798 (O_1798,N_24871,N_24657);
and UO_1799 (O_1799,N_24762,N_24956);
and UO_1800 (O_1800,N_24910,N_24746);
xor UO_1801 (O_1801,N_24779,N_24733);
and UO_1802 (O_1802,N_24508,N_24621);
and UO_1803 (O_1803,N_24901,N_24876);
nand UO_1804 (O_1804,N_24753,N_24996);
or UO_1805 (O_1805,N_24825,N_24689);
nor UO_1806 (O_1806,N_24952,N_24582);
and UO_1807 (O_1807,N_24614,N_24600);
or UO_1808 (O_1808,N_24683,N_24740);
and UO_1809 (O_1809,N_24902,N_24679);
nor UO_1810 (O_1810,N_24862,N_24604);
and UO_1811 (O_1811,N_24541,N_24828);
and UO_1812 (O_1812,N_24822,N_24730);
nor UO_1813 (O_1813,N_24839,N_24652);
nand UO_1814 (O_1814,N_24849,N_24714);
nor UO_1815 (O_1815,N_24667,N_24583);
or UO_1816 (O_1816,N_24650,N_24971);
nand UO_1817 (O_1817,N_24724,N_24533);
or UO_1818 (O_1818,N_24772,N_24630);
nor UO_1819 (O_1819,N_24546,N_24977);
nor UO_1820 (O_1820,N_24779,N_24958);
or UO_1821 (O_1821,N_24908,N_24804);
and UO_1822 (O_1822,N_24926,N_24524);
nand UO_1823 (O_1823,N_24603,N_24943);
nor UO_1824 (O_1824,N_24550,N_24853);
nand UO_1825 (O_1825,N_24522,N_24729);
or UO_1826 (O_1826,N_24778,N_24688);
and UO_1827 (O_1827,N_24689,N_24747);
nor UO_1828 (O_1828,N_24907,N_24882);
and UO_1829 (O_1829,N_24896,N_24852);
and UO_1830 (O_1830,N_24642,N_24850);
or UO_1831 (O_1831,N_24821,N_24520);
nor UO_1832 (O_1832,N_24647,N_24620);
nand UO_1833 (O_1833,N_24523,N_24836);
and UO_1834 (O_1834,N_24688,N_24790);
nand UO_1835 (O_1835,N_24852,N_24743);
nor UO_1836 (O_1836,N_24854,N_24909);
nand UO_1837 (O_1837,N_24914,N_24656);
and UO_1838 (O_1838,N_24587,N_24958);
nand UO_1839 (O_1839,N_24785,N_24868);
and UO_1840 (O_1840,N_24662,N_24535);
nand UO_1841 (O_1841,N_24948,N_24742);
nand UO_1842 (O_1842,N_24780,N_24894);
or UO_1843 (O_1843,N_24639,N_24916);
and UO_1844 (O_1844,N_24510,N_24573);
or UO_1845 (O_1845,N_24616,N_24565);
or UO_1846 (O_1846,N_24545,N_24838);
or UO_1847 (O_1847,N_24923,N_24936);
and UO_1848 (O_1848,N_24906,N_24635);
nor UO_1849 (O_1849,N_24586,N_24765);
and UO_1850 (O_1850,N_24991,N_24597);
nor UO_1851 (O_1851,N_24602,N_24910);
or UO_1852 (O_1852,N_24539,N_24615);
nor UO_1853 (O_1853,N_24955,N_24577);
and UO_1854 (O_1854,N_24728,N_24582);
or UO_1855 (O_1855,N_24914,N_24691);
nor UO_1856 (O_1856,N_24949,N_24922);
xor UO_1857 (O_1857,N_24886,N_24773);
and UO_1858 (O_1858,N_24871,N_24602);
or UO_1859 (O_1859,N_24683,N_24809);
nor UO_1860 (O_1860,N_24521,N_24976);
nand UO_1861 (O_1861,N_24703,N_24692);
and UO_1862 (O_1862,N_24832,N_24514);
or UO_1863 (O_1863,N_24609,N_24628);
nand UO_1864 (O_1864,N_24547,N_24750);
nand UO_1865 (O_1865,N_24517,N_24617);
and UO_1866 (O_1866,N_24575,N_24993);
and UO_1867 (O_1867,N_24803,N_24555);
xor UO_1868 (O_1868,N_24990,N_24809);
nor UO_1869 (O_1869,N_24540,N_24982);
nand UO_1870 (O_1870,N_24743,N_24776);
and UO_1871 (O_1871,N_24824,N_24995);
xnor UO_1872 (O_1872,N_24876,N_24763);
nand UO_1873 (O_1873,N_24649,N_24751);
nand UO_1874 (O_1874,N_24741,N_24922);
and UO_1875 (O_1875,N_24786,N_24552);
nand UO_1876 (O_1876,N_24948,N_24851);
or UO_1877 (O_1877,N_24961,N_24815);
nand UO_1878 (O_1878,N_24784,N_24564);
or UO_1879 (O_1879,N_24902,N_24978);
nand UO_1880 (O_1880,N_24837,N_24926);
nand UO_1881 (O_1881,N_24667,N_24614);
and UO_1882 (O_1882,N_24740,N_24823);
nor UO_1883 (O_1883,N_24574,N_24793);
or UO_1884 (O_1884,N_24810,N_24578);
xor UO_1885 (O_1885,N_24658,N_24965);
or UO_1886 (O_1886,N_24596,N_24901);
and UO_1887 (O_1887,N_24798,N_24537);
nand UO_1888 (O_1888,N_24540,N_24561);
nor UO_1889 (O_1889,N_24852,N_24728);
or UO_1890 (O_1890,N_24526,N_24534);
nor UO_1891 (O_1891,N_24827,N_24979);
nor UO_1892 (O_1892,N_24733,N_24551);
or UO_1893 (O_1893,N_24995,N_24834);
nor UO_1894 (O_1894,N_24535,N_24898);
and UO_1895 (O_1895,N_24767,N_24928);
nor UO_1896 (O_1896,N_24631,N_24801);
nand UO_1897 (O_1897,N_24632,N_24611);
nand UO_1898 (O_1898,N_24907,N_24661);
and UO_1899 (O_1899,N_24997,N_24702);
or UO_1900 (O_1900,N_24555,N_24958);
and UO_1901 (O_1901,N_24653,N_24528);
nand UO_1902 (O_1902,N_24537,N_24994);
xor UO_1903 (O_1903,N_24584,N_24929);
and UO_1904 (O_1904,N_24513,N_24536);
and UO_1905 (O_1905,N_24789,N_24739);
nand UO_1906 (O_1906,N_24561,N_24990);
nor UO_1907 (O_1907,N_24860,N_24550);
or UO_1908 (O_1908,N_24929,N_24834);
and UO_1909 (O_1909,N_24910,N_24763);
nand UO_1910 (O_1910,N_24743,N_24864);
xnor UO_1911 (O_1911,N_24958,N_24898);
nor UO_1912 (O_1912,N_24935,N_24563);
or UO_1913 (O_1913,N_24999,N_24544);
or UO_1914 (O_1914,N_24911,N_24658);
and UO_1915 (O_1915,N_24999,N_24723);
xnor UO_1916 (O_1916,N_24646,N_24620);
xor UO_1917 (O_1917,N_24850,N_24657);
or UO_1918 (O_1918,N_24817,N_24546);
and UO_1919 (O_1919,N_24589,N_24787);
nor UO_1920 (O_1920,N_24862,N_24798);
or UO_1921 (O_1921,N_24800,N_24998);
or UO_1922 (O_1922,N_24597,N_24517);
xnor UO_1923 (O_1923,N_24597,N_24849);
and UO_1924 (O_1924,N_24968,N_24684);
and UO_1925 (O_1925,N_24540,N_24747);
nor UO_1926 (O_1926,N_24678,N_24925);
and UO_1927 (O_1927,N_24514,N_24636);
and UO_1928 (O_1928,N_24895,N_24742);
nor UO_1929 (O_1929,N_24638,N_24832);
nor UO_1930 (O_1930,N_24639,N_24769);
nor UO_1931 (O_1931,N_24522,N_24824);
or UO_1932 (O_1932,N_24705,N_24970);
or UO_1933 (O_1933,N_24508,N_24843);
nand UO_1934 (O_1934,N_24894,N_24696);
or UO_1935 (O_1935,N_24993,N_24603);
and UO_1936 (O_1936,N_24722,N_24674);
nand UO_1937 (O_1937,N_24544,N_24560);
nor UO_1938 (O_1938,N_24905,N_24586);
nor UO_1939 (O_1939,N_24649,N_24709);
xnor UO_1940 (O_1940,N_24633,N_24908);
and UO_1941 (O_1941,N_24717,N_24941);
or UO_1942 (O_1942,N_24507,N_24710);
or UO_1943 (O_1943,N_24921,N_24674);
xor UO_1944 (O_1944,N_24751,N_24709);
nand UO_1945 (O_1945,N_24888,N_24508);
nand UO_1946 (O_1946,N_24530,N_24682);
or UO_1947 (O_1947,N_24882,N_24654);
nor UO_1948 (O_1948,N_24624,N_24970);
or UO_1949 (O_1949,N_24658,N_24924);
xor UO_1950 (O_1950,N_24645,N_24554);
or UO_1951 (O_1951,N_24743,N_24716);
and UO_1952 (O_1952,N_24874,N_24672);
nand UO_1953 (O_1953,N_24690,N_24796);
xor UO_1954 (O_1954,N_24826,N_24633);
or UO_1955 (O_1955,N_24836,N_24928);
or UO_1956 (O_1956,N_24712,N_24864);
nand UO_1957 (O_1957,N_24956,N_24618);
nor UO_1958 (O_1958,N_24526,N_24561);
nor UO_1959 (O_1959,N_24707,N_24634);
nand UO_1960 (O_1960,N_24866,N_24766);
and UO_1961 (O_1961,N_24825,N_24692);
nand UO_1962 (O_1962,N_24535,N_24886);
xor UO_1963 (O_1963,N_24592,N_24861);
nand UO_1964 (O_1964,N_24890,N_24865);
and UO_1965 (O_1965,N_24704,N_24543);
or UO_1966 (O_1966,N_24766,N_24898);
xor UO_1967 (O_1967,N_24793,N_24633);
xnor UO_1968 (O_1968,N_24947,N_24971);
nor UO_1969 (O_1969,N_24875,N_24754);
or UO_1970 (O_1970,N_24726,N_24892);
or UO_1971 (O_1971,N_24633,N_24892);
and UO_1972 (O_1972,N_24925,N_24913);
xnor UO_1973 (O_1973,N_24995,N_24786);
and UO_1974 (O_1974,N_24965,N_24976);
nand UO_1975 (O_1975,N_24830,N_24822);
and UO_1976 (O_1976,N_24910,N_24981);
or UO_1977 (O_1977,N_24516,N_24622);
nand UO_1978 (O_1978,N_24596,N_24616);
and UO_1979 (O_1979,N_24619,N_24557);
nor UO_1980 (O_1980,N_24877,N_24655);
nor UO_1981 (O_1981,N_24760,N_24776);
and UO_1982 (O_1982,N_24785,N_24835);
nor UO_1983 (O_1983,N_24526,N_24553);
and UO_1984 (O_1984,N_24536,N_24693);
xor UO_1985 (O_1985,N_24707,N_24952);
nand UO_1986 (O_1986,N_24562,N_24649);
nand UO_1987 (O_1987,N_24677,N_24864);
xor UO_1988 (O_1988,N_24534,N_24877);
and UO_1989 (O_1989,N_24992,N_24704);
nor UO_1990 (O_1990,N_24999,N_24507);
nand UO_1991 (O_1991,N_24569,N_24684);
and UO_1992 (O_1992,N_24987,N_24555);
nand UO_1993 (O_1993,N_24616,N_24961);
nand UO_1994 (O_1994,N_24558,N_24567);
or UO_1995 (O_1995,N_24848,N_24820);
or UO_1996 (O_1996,N_24911,N_24960);
or UO_1997 (O_1997,N_24725,N_24838);
nand UO_1998 (O_1998,N_24506,N_24757);
xor UO_1999 (O_1999,N_24987,N_24688);
xnor UO_2000 (O_2000,N_24817,N_24589);
nand UO_2001 (O_2001,N_24837,N_24716);
and UO_2002 (O_2002,N_24728,N_24561);
nand UO_2003 (O_2003,N_24976,N_24863);
nand UO_2004 (O_2004,N_24827,N_24762);
or UO_2005 (O_2005,N_24532,N_24908);
nand UO_2006 (O_2006,N_24924,N_24746);
nor UO_2007 (O_2007,N_24901,N_24640);
nand UO_2008 (O_2008,N_24501,N_24756);
nor UO_2009 (O_2009,N_24704,N_24531);
xnor UO_2010 (O_2010,N_24907,N_24610);
or UO_2011 (O_2011,N_24691,N_24979);
nand UO_2012 (O_2012,N_24670,N_24827);
or UO_2013 (O_2013,N_24838,N_24904);
or UO_2014 (O_2014,N_24858,N_24591);
nand UO_2015 (O_2015,N_24790,N_24927);
nand UO_2016 (O_2016,N_24847,N_24668);
xor UO_2017 (O_2017,N_24540,N_24895);
and UO_2018 (O_2018,N_24920,N_24802);
nor UO_2019 (O_2019,N_24834,N_24768);
or UO_2020 (O_2020,N_24749,N_24781);
and UO_2021 (O_2021,N_24626,N_24669);
or UO_2022 (O_2022,N_24726,N_24514);
and UO_2023 (O_2023,N_24641,N_24963);
and UO_2024 (O_2024,N_24791,N_24978);
and UO_2025 (O_2025,N_24512,N_24844);
nand UO_2026 (O_2026,N_24644,N_24870);
nor UO_2027 (O_2027,N_24688,N_24653);
nand UO_2028 (O_2028,N_24625,N_24926);
nor UO_2029 (O_2029,N_24504,N_24850);
or UO_2030 (O_2030,N_24625,N_24834);
and UO_2031 (O_2031,N_24695,N_24558);
nor UO_2032 (O_2032,N_24900,N_24582);
nand UO_2033 (O_2033,N_24683,N_24954);
nand UO_2034 (O_2034,N_24748,N_24655);
or UO_2035 (O_2035,N_24768,N_24915);
and UO_2036 (O_2036,N_24854,N_24786);
nor UO_2037 (O_2037,N_24745,N_24701);
nor UO_2038 (O_2038,N_24641,N_24851);
and UO_2039 (O_2039,N_24585,N_24749);
nor UO_2040 (O_2040,N_24569,N_24586);
nand UO_2041 (O_2041,N_24744,N_24859);
and UO_2042 (O_2042,N_24666,N_24871);
nand UO_2043 (O_2043,N_24986,N_24972);
and UO_2044 (O_2044,N_24666,N_24612);
and UO_2045 (O_2045,N_24684,N_24762);
or UO_2046 (O_2046,N_24519,N_24960);
nor UO_2047 (O_2047,N_24899,N_24683);
or UO_2048 (O_2048,N_24702,N_24595);
nor UO_2049 (O_2049,N_24891,N_24783);
and UO_2050 (O_2050,N_24675,N_24774);
or UO_2051 (O_2051,N_24529,N_24802);
and UO_2052 (O_2052,N_24735,N_24712);
xor UO_2053 (O_2053,N_24706,N_24709);
nor UO_2054 (O_2054,N_24826,N_24871);
nand UO_2055 (O_2055,N_24501,N_24850);
and UO_2056 (O_2056,N_24508,N_24920);
and UO_2057 (O_2057,N_24646,N_24693);
and UO_2058 (O_2058,N_24878,N_24639);
or UO_2059 (O_2059,N_24558,N_24694);
or UO_2060 (O_2060,N_24570,N_24778);
or UO_2061 (O_2061,N_24820,N_24812);
nor UO_2062 (O_2062,N_24664,N_24702);
and UO_2063 (O_2063,N_24815,N_24730);
nor UO_2064 (O_2064,N_24974,N_24533);
or UO_2065 (O_2065,N_24636,N_24912);
and UO_2066 (O_2066,N_24760,N_24634);
nor UO_2067 (O_2067,N_24547,N_24525);
xnor UO_2068 (O_2068,N_24725,N_24985);
and UO_2069 (O_2069,N_24563,N_24881);
or UO_2070 (O_2070,N_24892,N_24979);
and UO_2071 (O_2071,N_24611,N_24582);
or UO_2072 (O_2072,N_24844,N_24617);
or UO_2073 (O_2073,N_24783,N_24827);
and UO_2074 (O_2074,N_24749,N_24780);
nor UO_2075 (O_2075,N_24759,N_24549);
and UO_2076 (O_2076,N_24733,N_24818);
nor UO_2077 (O_2077,N_24761,N_24790);
nor UO_2078 (O_2078,N_24707,N_24657);
nor UO_2079 (O_2079,N_24759,N_24612);
nor UO_2080 (O_2080,N_24552,N_24823);
nand UO_2081 (O_2081,N_24926,N_24506);
nand UO_2082 (O_2082,N_24882,N_24872);
nand UO_2083 (O_2083,N_24611,N_24554);
nor UO_2084 (O_2084,N_24522,N_24569);
or UO_2085 (O_2085,N_24578,N_24865);
or UO_2086 (O_2086,N_24844,N_24560);
xnor UO_2087 (O_2087,N_24911,N_24904);
nor UO_2088 (O_2088,N_24556,N_24904);
and UO_2089 (O_2089,N_24906,N_24560);
and UO_2090 (O_2090,N_24692,N_24677);
and UO_2091 (O_2091,N_24523,N_24512);
nor UO_2092 (O_2092,N_24562,N_24626);
and UO_2093 (O_2093,N_24902,N_24717);
nor UO_2094 (O_2094,N_24947,N_24831);
nor UO_2095 (O_2095,N_24691,N_24690);
and UO_2096 (O_2096,N_24656,N_24593);
nor UO_2097 (O_2097,N_24642,N_24551);
nor UO_2098 (O_2098,N_24565,N_24787);
nand UO_2099 (O_2099,N_24976,N_24983);
and UO_2100 (O_2100,N_24838,N_24738);
nor UO_2101 (O_2101,N_24875,N_24900);
nand UO_2102 (O_2102,N_24644,N_24515);
and UO_2103 (O_2103,N_24766,N_24697);
nand UO_2104 (O_2104,N_24742,N_24513);
or UO_2105 (O_2105,N_24568,N_24840);
or UO_2106 (O_2106,N_24719,N_24844);
nand UO_2107 (O_2107,N_24521,N_24580);
or UO_2108 (O_2108,N_24837,N_24725);
nand UO_2109 (O_2109,N_24610,N_24750);
and UO_2110 (O_2110,N_24648,N_24877);
or UO_2111 (O_2111,N_24637,N_24840);
nand UO_2112 (O_2112,N_24772,N_24701);
nand UO_2113 (O_2113,N_24669,N_24697);
and UO_2114 (O_2114,N_24722,N_24922);
nor UO_2115 (O_2115,N_24532,N_24965);
nand UO_2116 (O_2116,N_24816,N_24506);
or UO_2117 (O_2117,N_24714,N_24934);
nand UO_2118 (O_2118,N_24512,N_24703);
nand UO_2119 (O_2119,N_24725,N_24930);
or UO_2120 (O_2120,N_24546,N_24764);
and UO_2121 (O_2121,N_24614,N_24539);
or UO_2122 (O_2122,N_24976,N_24716);
nand UO_2123 (O_2123,N_24653,N_24641);
xor UO_2124 (O_2124,N_24781,N_24927);
and UO_2125 (O_2125,N_24693,N_24600);
and UO_2126 (O_2126,N_24709,N_24738);
nor UO_2127 (O_2127,N_24756,N_24706);
and UO_2128 (O_2128,N_24863,N_24882);
nand UO_2129 (O_2129,N_24997,N_24841);
nand UO_2130 (O_2130,N_24829,N_24682);
or UO_2131 (O_2131,N_24984,N_24753);
nand UO_2132 (O_2132,N_24701,N_24747);
nand UO_2133 (O_2133,N_24934,N_24732);
and UO_2134 (O_2134,N_24538,N_24831);
or UO_2135 (O_2135,N_24642,N_24613);
nor UO_2136 (O_2136,N_24508,N_24764);
nand UO_2137 (O_2137,N_24587,N_24675);
or UO_2138 (O_2138,N_24902,N_24658);
and UO_2139 (O_2139,N_24742,N_24594);
or UO_2140 (O_2140,N_24912,N_24639);
and UO_2141 (O_2141,N_24617,N_24855);
or UO_2142 (O_2142,N_24801,N_24751);
or UO_2143 (O_2143,N_24634,N_24750);
nand UO_2144 (O_2144,N_24806,N_24959);
nand UO_2145 (O_2145,N_24795,N_24946);
nand UO_2146 (O_2146,N_24556,N_24715);
or UO_2147 (O_2147,N_24591,N_24652);
nand UO_2148 (O_2148,N_24857,N_24677);
xnor UO_2149 (O_2149,N_24507,N_24851);
or UO_2150 (O_2150,N_24580,N_24696);
nand UO_2151 (O_2151,N_24757,N_24581);
nand UO_2152 (O_2152,N_24869,N_24862);
nand UO_2153 (O_2153,N_24787,N_24793);
or UO_2154 (O_2154,N_24549,N_24538);
nor UO_2155 (O_2155,N_24550,N_24936);
or UO_2156 (O_2156,N_24819,N_24742);
and UO_2157 (O_2157,N_24747,N_24702);
nor UO_2158 (O_2158,N_24582,N_24774);
or UO_2159 (O_2159,N_24728,N_24558);
nand UO_2160 (O_2160,N_24728,N_24742);
xor UO_2161 (O_2161,N_24904,N_24712);
and UO_2162 (O_2162,N_24793,N_24946);
and UO_2163 (O_2163,N_24552,N_24788);
and UO_2164 (O_2164,N_24747,N_24888);
nand UO_2165 (O_2165,N_24778,N_24853);
or UO_2166 (O_2166,N_24966,N_24539);
and UO_2167 (O_2167,N_24524,N_24907);
and UO_2168 (O_2168,N_24519,N_24609);
nor UO_2169 (O_2169,N_24752,N_24988);
and UO_2170 (O_2170,N_24768,N_24512);
nand UO_2171 (O_2171,N_24626,N_24809);
nand UO_2172 (O_2172,N_24979,N_24972);
and UO_2173 (O_2173,N_24852,N_24550);
xnor UO_2174 (O_2174,N_24515,N_24650);
nor UO_2175 (O_2175,N_24582,N_24660);
xnor UO_2176 (O_2176,N_24639,N_24913);
and UO_2177 (O_2177,N_24871,N_24974);
or UO_2178 (O_2178,N_24893,N_24604);
xnor UO_2179 (O_2179,N_24672,N_24948);
or UO_2180 (O_2180,N_24912,N_24617);
nand UO_2181 (O_2181,N_24935,N_24756);
nand UO_2182 (O_2182,N_24549,N_24661);
and UO_2183 (O_2183,N_24999,N_24741);
and UO_2184 (O_2184,N_24775,N_24730);
and UO_2185 (O_2185,N_24577,N_24576);
nor UO_2186 (O_2186,N_24543,N_24921);
nor UO_2187 (O_2187,N_24871,N_24942);
nand UO_2188 (O_2188,N_24564,N_24685);
xnor UO_2189 (O_2189,N_24735,N_24539);
nand UO_2190 (O_2190,N_24880,N_24837);
nand UO_2191 (O_2191,N_24900,N_24796);
or UO_2192 (O_2192,N_24564,N_24820);
nand UO_2193 (O_2193,N_24754,N_24605);
and UO_2194 (O_2194,N_24700,N_24927);
or UO_2195 (O_2195,N_24982,N_24634);
or UO_2196 (O_2196,N_24607,N_24586);
or UO_2197 (O_2197,N_24538,N_24578);
and UO_2198 (O_2198,N_24998,N_24846);
or UO_2199 (O_2199,N_24557,N_24901);
and UO_2200 (O_2200,N_24875,N_24947);
xnor UO_2201 (O_2201,N_24645,N_24972);
or UO_2202 (O_2202,N_24729,N_24831);
or UO_2203 (O_2203,N_24794,N_24975);
or UO_2204 (O_2204,N_24793,N_24936);
nand UO_2205 (O_2205,N_24857,N_24797);
nor UO_2206 (O_2206,N_24662,N_24831);
and UO_2207 (O_2207,N_24961,N_24574);
or UO_2208 (O_2208,N_24735,N_24857);
and UO_2209 (O_2209,N_24853,N_24723);
and UO_2210 (O_2210,N_24767,N_24755);
nand UO_2211 (O_2211,N_24915,N_24965);
or UO_2212 (O_2212,N_24957,N_24866);
nand UO_2213 (O_2213,N_24646,N_24872);
and UO_2214 (O_2214,N_24996,N_24628);
nand UO_2215 (O_2215,N_24849,N_24955);
and UO_2216 (O_2216,N_24830,N_24949);
nor UO_2217 (O_2217,N_24747,N_24984);
and UO_2218 (O_2218,N_24520,N_24772);
nand UO_2219 (O_2219,N_24964,N_24808);
xor UO_2220 (O_2220,N_24956,N_24863);
and UO_2221 (O_2221,N_24513,N_24758);
nor UO_2222 (O_2222,N_24891,N_24540);
or UO_2223 (O_2223,N_24812,N_24608);
nand UO_2224 (O_2224,N_24740,N_24975);
or UO_2225 (O_2225,N_24632,N_24927);
and UO_2226 (O_2226,N_24639,N_24804);
nand UO_2227 (O_2227,N_24745,N_24584);
and UO_2228 (O_2228,N_24873,N_24581);
or UO_2229 (O_2229,N_24662,N_24634);
nor UO_2230 (O_2230,N_24639,N_24810);
nor UO_2231 (O_2231,N_24521,N_24571);
and UO_2232 (O_2232,N_24628,N_24796);
and UO_2233 (O_2233,N_24607,N_24998);
nor UO_2234 (O_2234,N_24519,N_24523);
or UO_2235 (O_2235,N_24994,N_24586);
nand UO_2236 (O_2236,N_24799,N_24756);
or UO_2237 (O_2237,N_24682,N_24923);
and UO_2238 (O_2238,N_24834,N_24962);
and UO_2239 (O_2239,N_24728,N_24581);
nand UO_2240 (O_2240,N_24711,N_24784);
nand UO_2241 (O_2241,N_24839,N_24768);
nor UO_2242 (O_2242,N_24531,N_24503);
nand UO_2243 (O_2243,N_24687,N_24740);
nor UO_2244 (O_2244,N_24597,N_24883);
and UO_2245 (O_2245,N_24873,N_24590);
nand UO_2246 (O_2246,N_24620,N_24578);
and UO_2247 (O_2247,N_24529,N_24763);
and UO_2248 (O_2248,N_24673,N_24660);
or UO_2249 (O_2249,N_24677,N_24622);
or UO_2250 (O_2250,N_24576,N_24745);
and UO_2251 (O_2251,N_24916,N_24896);
nor UO_2252 (O_2252,N_24795,N_24537);
xor UO_2253 (O_2253,N_24728,N_24563);
and UO_2254 (O_2254,N_24968,N_24893);
nor UO_2255 (O_2255,N_24851,N_24726);
and UO_2256 (O_2256,N_24961,N_24861);
or UO_2257 (O_2257,N_24671,N_24838);
and UO_2258 (O_2258,N_24618,N_24631);
and UO_2259 (O_2259,N_24922,N_24564);
and UO_2260 (O_2260,N_24979,N_24917);
nand UO_2261 (O_2261,N_24510,N_24908);
nand UO_2262 (O_2262,N_24622,N_24709);
xor UO_2263 (O_2263,N_24790,N_24826);
or UO_2264 (O_2264,N_24661,N_24690);
nand UO_2265 (O_2265,N_24503,N_24850);
xnor UO_2266 (O_2266,N_24678,N_24643);
xor UO_2267 (O_2267,N_24956,N_24566);
and UO_2268 (O_2268,N_24958,N_24758);
nor UO_2269 (O_2269,N_24839,N_24571);
nor UO_2270 (O_2270,N_24969,N_24650);
and UO_2271 (O_2271,N_24997,N_24850);
or UO_2272 (O_2272,N_24895,N_24965);
nor UO_2273 (O_2273,N_24703,N_24723);
xor UO_2274 (O_2274,N_24705,N_24624);
or UO_2275 (O_2275,N_24603,N_24506);
and UO_2276 (O_2276,N_24885,N_24745);
nand UO_2277 (O_2277,N_24903,N_24918);
or UO_2278 (O_2278,N_24708,N_24563);
nand UO_2279 (O_2279,N_24794,N_24940);
nand UO_2280 (O_2280,N_24800,N_24944);
and UO_2281 (O_2281,N_24948,N_24980);
and UO_2282 (O_2282,N_24947,N_24786);
and UO_2283 (O_2283,N_24870,N_24593);
nor UO_2284 (O_2284,N_24744,N_24840);
and UO_2285 (O_2285,N_24604,N_24848);
nor UO_2286 (O_2286,N_24606,N_24619);
nor UO_2287 (O_2287,N_24509,N_24829);
nand UO_2288 (O_2288,N_24597,N_24857);
or UO_2289 (O_2289,N_24502,N_24607);
or UO_2290 (O_2290,N_24502,N_24937);
nand UO_2291 (O_2291,N_24844,N_24596);
nand UO_2292 (O_2292,N_24866,N_24504);
or UO_2293 (O_2293,N_24706,N_24585);
nor UO_2294 (O_2294,N_24639,N_24549);
and UO_2295 (O_2295,N_24511,N_24517);
and UO_2296 (O_2296,N_24664,N_24530);
and UO_2297 (O_2297,N_24780,N_24513);
nor UO_2298 (O_2298,N_24841,N_24920);
and UO_2299 (O_2299,N_24655,N_24894);
nor UO_2300 (O_2300,N_24503,N_24686);
nand UO_2301 (O_2301,N_24596,N_24670);
or UO_2302 (O_2302,N_24697,N_24953);
and UO_2303 (O_2303,N_24809,N_24767);
nand UO_2304 (O_2304,N_24743,N_24573);
nand UO_2305 (O_2305,N_24675,N_24959);
or UO_2306 (O_2306,N_24840,N_24741);
and UO_2307 (O_2307,N_24661,N_24753);
nor UO_2308 (O_2308,N_24872,N_24915);
nor UO_2309 (O_2309,N_24849,N_24516);
and UO_2310 (O_2310,N_24502,N_24504);
nor UO_2311 (O_2311,N_24945,N_24584);
and UO_2312 (O_2312,N_24846,N_24831);
and UO_2313 (O_2313,N_24800,N_24561);
nand UO_2314 (O_2314,N_24744,N_24666);
nand UO_2315 (O_2315,N_24724,N_24793);
or UO_2316 (O_2316,N_24934,N_24737);
and UO_2317 (O_2317,N_24653,N_24699);
nor UO_2318 (O_2318,N_24925,N_24633);
nor UO_2319 (O_2319,N_24671,N_24999);
nand UO_2320 (O_2320,N_24790,N_24555);
and UO_2321 (O_2321,N_24618,N_24734);
and UO_2322 (O_2322,N_24587,N_24707);
and UO_2323 (O_2323,N_24849,N_24664);
nor UO_2324 (O_2324,N_24962,N_24914);
and UO_2325 (O_2325,N_24635,N_24843);
and UO_2326 (O_2326,N_24906,N_24878);
nor UO_2327 (O_2327,N_24645,N_24543);
and UO_2328 (O_2328,N_24509,N_24737);
nor UO_2329 (O_2329,N_24742,N_24780);
nand UO_2330 (O_2330,N_24613,N_24906);
nor UO_2331 (O_2331,N_24807,N_24900);
nor UO_2332 (O_2332,N_24971,N_24559);
xnor UO_2333 (O_2333,N_24880,N_24668);
nor UO_2334 (O_2334,N_24920,N_24695);
or UO_2335 (O_2335,N_24749,N_24797);
nor UO_2336 (O_2336,N_24999,N_24552);
and UO_2337 (O_2337,N_24938,N_24861);
or UO_2338 (O_2338,N_24510,N_24999);
and UO_2339 (O_2339,N_24845,N_24996);
nor UO_2340 (O_2340,N_24704,N_24878);
and UO_2341 (O_2341,N_24667,N_24691);
nand UO_2342 (O_2342,N_24645,N_24720);
nor UO_2343 (O_2343,N_24733,N_24725);
nand UO_2344 (O_2344,N_24797,N_24852);
or UO_2345 (O_2345,N_24825,N_24799);
or UO_2346 (O_2346,N_24970,N_24616);
xnor UO_2347 (O_2347,N_24644,N_24967);
or UO_2348 (O_2348,N_24510,N_24797);
nor UO_2349 (O_2349,N_24556,N_24935);
or UO_2350 (O_2350,N_24836,N_24991);
nand UO_2351 (O_2351,N_24982,N_24895);
or UO_2352 (O_2352,N_24974,N_24616);
nand UO_2353 (O_2353,N_24559,N_24763);
nand UO_2354 (O_2354,N_24791,N_24539);
nor UO_2355 (O_2355,N_24776,N_24692);
or UO_2356 (O_2356,N_24864,N_24878);
and UO_2357 (O_2357,N_24889,N_24515);
nor UO_2358 (O_2358,N_24558,N_24646);
or UO_2359 (O_2359,N_24988,N_24883);
or UO_2360 (O_2360,N_24736,N_24612);
xor UO_2361 (O_2361,N_24726,N_24979);
xor UO_2362 (O_2362,N_24607,N_24939);
and UO_2363 (O_2363,N_24952,N_24511);
xnor UO_2364 (O_2364,N_24572,N_24666);
nor UO_2365 (O_2365,N_24711,N_24836);
and UO_2366 (O_2366,N_24916,N_24987);
or UO_2367 (O_2367,N_24606,N_24692);
nand UO_2368 (O_2368,N_24781,N_24757);
xnor UO_2369 (O_2369,N_24781,N_24887);
or UO_2370 (O_2370,N_24865,N_24766);
nand UO_2371 (O_2371,N_24572,N_24974);
nor UO_2372 (O_2372,N_24829,N_24505);
and UO_2373 (O_2373,N_24996,N_24507);
nor UO_2374 (O_2374,N_24858,N_24768);
and UO_2375 (O_2375,N_24836,N_24656);
xnor UO_2376 (O_2376,N_24939,N_24507);
or UO_2377 (O_2377,N_24571,N_24820);
or UO_2378 (O_2378,N_24869,N_24620);
and UO_2379 (O_2379,N_24851,N_24680);
or UO_2380 (O_2380,N_24822,N_24966);
or UO_2381 (O_2381,N_24612,N_24921);
and UO_2382 (O_2382,N_24737,N_24782);
and UO_2383 (O_2383,N_24757,N_24879);
nor UO_2384 (O_2384,N_24793,N_24908);
nand UO_2385 (O_2385,N_24562,N_24897);
xor UO_2386 (O_2386,N_24717,N_24583);
or UO_2387 (O_2387,N_24858,N_24934);
and UO_2388 (O_2388,N_24872,N_24921);
nor UO_2389 (O_2389,N_24771,N_24617);
or UO_2390 (O_2390,N_24651,N_24717);
nand UO_2391 (O_2391,N_24733,N_24917);
or UO_2392 (O_2392,N_24808,N_24815);
nand UO_2393 (O_2393,N_24936,N_24788);
or UO_2394 (O_2394,N_24833,N_24829);
nor UO_2395 (O_2395,N_24641,N_24520);
and UO_2396 (O_2396,N_24613,N_24707);
nor UO_2397 (O_2397,N_24623,N_24828);
nand UO_2398 (O_2398,N_24560,N_24714);
or UO_2399 (O_2399,N_24874,N_24743);
nand UO_2400 (O_2400,N_24967,N_24840);
nor UO_2401 (O_2401,N_24947,N_24617);
nand UO_2402 (O_2402,N_24561,N_24815);
and UO_2403 (O_2403,N_24641,N_24957);
and UO_2404 (O_2404,N_24881,N_24710);
and UO_2405 (O_2405,N_24919,N_24562);
and UO_2406 (O_2406,N_24894,N_24818);
nand UO_2407 (O_2407,N_24597,N_24895);
nor UO_2408 (O_2408,N_24881,N_24784);
nor UO_2409 (O_2409,N_24879,N_24841);
nand UO_2410 (O_2410,N_24935,N_24768);
and UO_2411 (O_2411,N_24657,N_24547);
or UO_2412 (O_2412,N_24891,N_24771);
nand UO_2413 (O_2413,N_24513,N_24818);
nand UO_2414 (O_2414,N_24580,N_24930);
nand UO_2415 (O_2415,N_24891,N_24620);
nand UO_2416 (O_2416,N_24870,N_24817);
nor UO_2417 (O_2417,N_24820,N_24560);
or UO_2418 (O_2418,N_24629,N_24825);
nand UO_2419 (O_2419,N_24935,N_24832);
or UO_2420 (O_2420,N_24607,N_24548);
nor UO_2421 (O_2421,N_24508,N_24808);
or UO_2422 (O_2422,N_24722,N_24507);
or UO_2423 (O_2423,N_24701,N_24525);
or UO_2424 (O_2424,N_24555,N_24729);
or UO_2425 (O_2425,N_24735,N_24893);
xor UO_2426 (O_2426,N_24590,N_24928);
or UO_2427 (O_2427,N_24887,N_24613);
nand UO_2428 (O_2428,N_24629,N_24995);
nor UO_2429 (O_2429,N_24777,N_24726);
nand UO_2430 (O_2430,N_24968,N_24587);
nor UO_2431 (O_2431,N_24566,N_24804);
or UO_2432 (O_2432,N_24739,N_24514);
nand UO_2433 (O_2433,N_24726,N_24606);
nor UO_2434 (O_2434,N_24815,N_24667);
nor UO_2435 (O_2435,N_24962,N_24546);
and UO_2436 (O_2436,N_24793,N_24853);
nand UO_2437 (O_2437,N_24926,N_24548);
nand UO_2438 (O_2438,N_24971,N_24664);
and UO_2439 (O_2439,N_24724,N_24958);
and UO_2440 (O_2440,N_24814,N_24826);
xnor UO_2441 (O_2441,N_24517,N_24996);
nor UO_2442 (O_2442,N_24801,N_24546);
nor UO_2443 (O_2443,N_24736,N_24915);
or UO_2444 (O_2444,N_24551,N_24881);
and UO_2445 (O_2445,N_24969,N_24730);
and UO_2446 (O_2446,N_24601,N_24687);
and UO_2447 (O_2447,N_24786,N_24844);
and UO_2448 (O_2448,N_24516,N_24540);
nor UO_2449 (O_2449,N_24501,N_24971);
nor UO_2450 (O_2450,N_24604,N_24792);
nand UO_2451 (O_2451,N_24596,N_24750);
nor UO_2452 (O_2452,N_24503,N_24817);
nor UO_2453 (O_2453,N_24628,N_24775);
and UO_2454 (O_2454,N_24600,N_24846);
nand UO_2455 (O_2455,N_24779,N_24964);
nand UO_2456 (O_2456,N_24647,N_24789);
or UO_2457 (O_2457,N_24605,N_24641);
nand UO_2458 (O_2458,N_24842,N_24808);
or UO_2459 (O_2459,N_24738,N_24607);
nor UO_2460 (O_2460,N_24637,N_24632);
nand UO_2461 (O_2461,N_24507,N_24528);
and UO_2462 (O_2462,N_24716,N_24896);
nor UO_2463 (O_2463,N_24533,N_24985);
and UO_2464 (O_2464,N_24836,N_24920);
or UO_2465 (O_2465,N_24964,N_24502);
or UO_2466 (O_2466,N_24578,N_24679);
or UO_2467 (O_2467,N_24848,N_24983);
or UO_2468 (O_2468,N_24829,N_24642);
nor UO_2469 (O_2469,N_24976,N_24865);
and UO_2470 (O_2470,N_24631,N_24612);
xor UO_2471 (O_2471,N_24503,N_24582);
nand UO_2472 (O_2472,N_24805,N_24580);
nor UO_2473 (O_2473,N_24855,N_24905);
or UO_2474 (O_2474,N_24973,N_24695);
nand UO_2475 (O_2475,N_24918,N_24876);
and UO_2476 (O_2476,N_24772,N_24899);
nor UO_2477 (O_2477,N_24532,N_24793);
or UO_2478 (O_2478,N_24981,N_24962);
nor UO_2479 (O_2479,N_24658,N_24869);
and UO_2480 (O_2480,N_24758,N_24979);
nor UO_2481 (O_2481,N_24767,N_24845);
or UO_2482 (O_2482,N_24555,N_24957);
nor UO_2483 (O_2483,N_24662,N_24588);
and UO_2484 (O_2484,N_24700,N_24635);
or UO_2485 (O_2485,N_24894,N_24905);
and UO_2486 (O_2486,N_24723,N_24910);
or UO_2487 (O_2487,N_24641,N_24587);
nor UO_2488 (O_2488,N_24611,N_24939);
xnor UO_2489 (O_2489,N_24741,N_24961);
nor UO_2490 (O_2490,N_24971,N_24698);
xor UO_2491 (O_2491,N_24500,N_24580);
nor UO_2492 (O_2492,N_24937,N_24624);
and UO_2493 (O_2493,N_24695,N_24872);
and UO_2494 (O_2494,N_24576,N_24712);
and UO_2495 (O_2495,N_24712,N_24729);
xor UO_2496 (O_2496,N_24562,N_24555);
xor UO_2497 (O_2497,N_24779,N_24931);
and UO_2498 (O_2498,N_24786,N_24954);
nor UO_2499 (O_2499,N_24888,N_24717);
or UO_2500 (O_2500,N_24646,N_24860);
and UO_2501 (O_2501,N_24553,N_24721);
nor UO_2502 (O_2502,N_24573,N_24760);
or UO_2503 (O_2503,N_24666,N_24605);
or UO_2504 (O_2504,N_24568,N_24987);
nor UO_2505 (O_2505,N_24973,N_24939);
nor UO_2506 (O_2506,N_24940,N_24827);
and UO_2507 (O_2507,N_24634,N_24508);
and UO_2508 (O_2508,N_24899,N_24563);
nand UO_2509 (O_2509,N_24887,N_24903);
nor UO_2510 (O_2510,N_24975,N_24715);
nand UO_2511 (O_2511,N_24568,N_24532);
nand UO_2512 (O_2512,N_24801,N_24813);
and UO_2513 (O_2513,N_24954,N_24515);
nand UO_2514 (O_2514,N_24846,N_24968);
or UO_2515 (O_2515,N_24895,N_24585);
and UO_2516 (O_2516,N_24981,N_24922);
xnor UO_2517 (O_2517,N_24576,N_24539);
nand UO_2518 (O_2518,N_24666,N_24753);
nand UO_2519 (O_2519,N_24994,N_24714);
nor UO_2520 (O_2520,N_24636,N_24680);
nand UO_2521 (O_2521,N_24707,N_24800);
nand UO_2522 (O_2522,N_24511,N_24984);
or UO_2523 (O_2523,N_24508,N_24857);
nor UO_2524 (O_2524,N_24701,N_24939);
nand UO_2525 (O_2525,N_24727,N_24664);
nand UO_2526 (O_2526,N_24537,N_24827);
or UO_2527 (O_2527,N_24708,N_24502);
nor UO_2528 (O_2528,N_24746,N_24785);
or UO_2529 (O_2529,N_24827,N_24910);
or UO_2530 (O_2530,N_24825,N_24529);
or UO_2531 (O_2531,N_24964,N_24915);
nor UO_2532 (O_2532,N_24583,N_24851);
or UO_2533 (O_2533,N_24974,N_24964);
or UO_2534 (O_2534,N_24746,N_24536);
nand UO_2535 (O_2535,N_24762,N_24645);
nand UO_2536 (O_2536,N_24520,N_24516);
nand UO_2537 (O_2537,N_24964,N_24538);
xor UO_2538 (O_2538,N_24712,N_24643);
and UO_2539 (O_2539,N_24909,N_24578);
nor UO_2540 (O_2540,N_24595,N_24972);
xor UO_2541 (O_2541,N_24522,N_24644);
nand UO_2542 (O_2542,N_24811,N_24593);
nand UO_2543 (O_2543,N_24848,N_24797);
or UO_2544 (O_2544,N_24507,N_24766);
nor UO_2545 (O_2545,N_24931,N_24579);
nor UO_2546 (O_2546,N_24681,N_24972);
nand UO_2547 (O_2547,N_24563,N_24934);
and UO_2548 (O_2548,N_24698,N_24910);
xor UO_2549 (O_2549,N_24808,N_24992);
or UO_2550 (O_2550,N_24871,N_24883);
nor UO_2551 (O_2551,N_24792,N_24974);
or UO_2552 (O_2552,N_24899,N_24809);
or UO_2553 (O_2553,N_24630,N_24875);
nand UO_2554 (O_2554,N_24951,N_24794);
and UO_2555 (O_2555,N_24996,N_24749);
nor UO_2556 (O_2556,N_24500,N_24955);
nand UO_2557 (O_2557,N_24595,N_24662);
or UO_2558 (O_2558,N_24664,N_24934);
or UO_2559 (O_2559,N_24601,N_24809);
xnor UO_2560 (O_2560,N_24921,N_24733);
or UO_2561 (O_2561,N_24893,N_24578);
and UO_2562 (O_2562,N_24805,N_24887);
or UO_2563 (O_2563,N_24810,N_24612);
nor UO_2564 (O_2564,N_24687,N_24560);
or UO_2565 (O_2565,N_24741,N_24744);
or UO_2566 (O_2566,N_24933,N_24990);
and UO_2567 (O_2567,N_24600,N_24666);
and UO_2568 (O_2568,N_24689,N_24706);
and UO_2569 (O_2569,N_24781,N_24755);
nor UO_2570 (O_2570,N_24970,N_24968);
and UO_2571 (O_2571,N_24564,N_24879);
and UO_2572 (O_2572,N_24678,N_24746);
nor UO_2573 (O_2573,N_24547,N_24534);
and UO_2574 (O_2574,N_24521,N_24623);
and UO_2575 (O_2575,N_24888,N_24942);
or UO_2576 (O_2576,N_24626,N_24573);
and UO_2577 (O_2577,N_24986,N_24623);
or UO_2578 (O_2578,N_24974,N_24535);
nand UO_2579 (O_2579,N_24785,N_24530);
and UO_2580 (O_2580,N_24921,N_24847);
or UO_2581 (O_2581,N_24939,N_24934);
xor UO_2582 (O_2582,N_24696,N_24788);
or UO_2583 (O_2583,N_24816,N_24966);
nor UO_2584 (O_2584,N_24713,N_24636);
nor UO_2585 (O_2585,N_24948,N_24866);
and UO_2586 (O_2586,N_24775,N_24647);
nor UO_2587 (O_2587,N_24723,N_24869);
nand UO_2588 (O_2588,N_24552,N_24527);
and UO_2589 (O_2589,N_24594,N_24572);
nor UO_2590 (O_2590,N_24964,N_24841);
and UO_2591 (O_2591,N_24823,N_24733);
xnor UO_2592 (O_2592,N_24726,N_24694);
or UO_2593 (O_2593,N_24677,N_24821);
nand UO_2594 (O_2594,N_24508,N_24707);
and UO_2595 (O_2595,N_24813,N_24812);
or UO_2596 (O_2596,N_24530,N_24540);
and UO_2597 (O_2597,N_24678,N_24774);
nand UO_2598 (O_2598,N_24857,N_24682);
and UO_2599 (O_2599,N_24820,N_24831);
and UO_2600 (O_2600,N_24799,N_24512);
nand UO_2601 (O_2601,N_24949,N_24542);
nor UO_2602 (O_2602,N_24860,N_24939);
or UO_2603 (O_2603,N_24697,N_24659);
xnor UO_2604 (O_2604,N_24880,N_24697);
or UO_2605 (O_2605,N_24738,N_24764);
or UO_2606 (O_2606,N_24636,N_24694);
or UO_2607 (O_2607,N_24671,N_24934);
nand UO_2608 (O_2608,N_24736,N_24849);
or UO_2609 (O_2609,N_24987,N_24774);
or UO_2610 (O_2610,N_24834,N_24904);
or UO_2611 (O_2611,N_24560,N_24621);
nand UO_2612 (O_2612,N_24581,N_24986);
and UO_2613 (O_2613,N_24981,N_24749);
and UO_2614 (O_2614,N_24975,N_24739);
xnor UO_2615 (O_2615,N_24817,N_24958);
or UO_2616 (O_2616,N_24581,N_24771);
and UO_2617 (O_2617,N_24901,N_24616);
and UO_2618 (O_2618,N_24568,N_24907);
and UO_2619 (O_2619,N_24887,N_24538);
or UO_2620 (O_2620,N_24598,N_24654);
xnor UO_2621 (O_2621,N_24639,N_24691);
nand UO_2622 (O_2622,N_24712,N_24649);
nand UO_2623 (O_2623,N_24774,N_24525);
and UO_2624 (O_2624,N_24616,N_24874);
and UO_2625 (O_2625,N_24811,N_24973);
nand UO_2626 (O_2626,N_24823,N_24808);
nor UO_2627 (O_2627,N_24531,N_24523);
or UO_2628 (O_2628,N_24805,N_24901);
or UO_2629 (O_2629,N_24807,N_24509);
and UO_2630 (O_2630,N_24547,N_24549);
and UO_2631 (O_2631,N_24897,N_24740);
nor UO_2632 (O_2632,N_24973,N_24831);
or UO_2633 (O_2633,N_24745,N_24830);
xnor UO_2634 (O_2634,N_24602,N_24987);
xor UO_2635 (O_2635,N_24875,N_24712);
nand UO_2636 (O_2636,N_24758,N_24517);
and UO_2637 (O_2637,N_24809,N_24792);
nand UO_2638 (O_2638,N_24707,N_24602);
or UO_2639 (O_2639,N_24535,N_24947);
xor UO_2640 (O_2640,N_24601,N_24947);
nor UO_2641 (O_2641,N_24712,N_24588);
or UO_2642 (O_2642,N_24781,N_24759);
or UO_2643 (O_2643,N_24998,N_24686);
and UO_2644 (O_2644,N_24618,N_24798);
nor UO_2645 (O_2645,N_24770,N_24501);
nor UO_2646 (O_2646,N_24836,N_24512);
nand UO_2647 (O_2647,N_24981,N_24570);
nor UO_2648 (O_2648,N_24762,N_24582);
or UO_2649 (O_2649,N_24930,N_24743);
nand UO_2650 (O_2650,N_24752,N_24614);
nand UO_2651 (O_2651,N_24766,N_24674);
nor UO_2652 (O_2652,N_24905,N_24641);
or UO_2653 (O_2653,N_24765,N_24966);
xor UO_2654 (O_2654,N_24664,N_24589);
and UO_2655 (O_2655,N_24832,N_24722);
nor UO_2656 (O_2656,N_24672,N_24517);
or UO_2657 (O_2657,N_24938,N_24674);
and UO_2658 (O_2658,N_24707,N_24583);
xor UO_2659 (O_2659,N_24926,N_24964);
or UO_2660 (O_2660,N_24533,N_24755);
or UO_2661 (O_2661,N_24733,N_24570);
or UO_2662 (O_2662,N_24875,N_24781);
and UO_2663 (O_2663,N_24662,N_24608);
nand UO_2664 (O_2664,N_24525,N_24772);
nand UO_2665 (O_2665,N_24579,N_24555);
nand UO_2666 (O_2666,N_24693,N_24938);
nor UO_2667 (O_2667,N_24611,N_24744);
nor UO_2668 (O_2668,N_24994,N_24867);
nand UO_2669 (O_2669,N_24815,N_24751);
and UO_2670 (O_2670,N_24765,N_24781);
nor UO_2671 (O_2671,N_24517,N_24504);
or UO_2672 (O_2672,N_24953,N_24562);
nand UO_2673 (O_2673,N_24757,N_24676);
nand UO_2674 (O_2674,N_24753,N_24956);
nor UO_2675 (O_2675,N_24689,N_24847);
nor UO_2676 (O_2676,N_24995,N_24501);
xnor UO_2677 (O_2677,N_24522,N_24855);
or UO_2678 (O_2678,N_24525,N_24663);
nor UO_2679 (O_2679,N_24779,N_24736);
or UO_2680 (O_2680,N_24904,N_24516);
or UO_2681 (O_2681,N_24819,N_24573);
and UO_2682 (O_2682,N_24964,N_24818);
nor UO_2683 (O_2683,N_24922,N_24714);
nand UO_2684 (O_2684,N_24969,N_24909);
or UO_2685 (O_2685,N_24594,N_24911);
nand UO_2686 (O_2686,N_24883,N_24801);
nor UO_2687 (O_2687,N_24854,N_24853);
xnor UO_2688 (O_2688,N_24947,N_24676);
or UO_2689 (O_2689,N_24544,N_24700);
nand UO_2690 (O_2690,N_24875,N_24611);
nand UO_2691 (O_2691,N_24815,N_24653);
nand UO_2692 (O_2692,N_24751,N_24580);
nand UO_2693 (O_2693,N_24957,N_24533);
and UO_2694 (O_2694,N_24729,N_24578);
and UO_2695 (O_2695,N_24653,N_24820);
nor UO_2696 (O_2696,N_24830,N_24753);
nor UO_2697 (O_2697,N_24696,N_24798);
nor UO_2698 (O_2698,N_24738,N_24940);
nor UO_2699 (O_2699,N_24919,N_24944);
and UO_2700 (O_2700,N_24702,N_24955);
nand UO_2701 (O_2701,N_24945,N_24680);
and UO_2702 (O_2702,N_24524,N_24543);
and UO_2703 (O_2703,N_24658,N_24620);
or UO_2704 (O_2704,N_24529,N_24933);
and UO_2705 (O_2705,N_24989,N_24951);
nand UO_2706 (O_2706,N_24927,N_24645);
nor UO_2707 (O_2707,N_24787,N_24613);
nand UO_2708 (O_2708,N_24860,N_24649);
and UO_2709 (O_2709,N_24752,N_24512);
xnor UO_2710 (O_2710,N_24688,N_24723);
nand UO_2711 (O_2711,N_24702,N_24945);
or UO_2712 (O_2712,N_24905,N_24707);
or UO_2713 (O_2713,N_24560,N_24704);
nor UO_2714 (O_2714,N_24678,N_24668);
or UO_2715 (O_2715,N_24663,N_24587);
xor UO_2716 (O_2716,N_24765,N_24574);
or UO_2717 (O_2717,N_24808,N_24831);
nand UO_2718 (O_2718,N_24555,N_24512);
or UO_2719 (O_2719,N_24986,N_24603);
and UO_2720 (O_2720,N_24671,N_24776);
and UO_2721 (O_2721,N_24689,N_24773);
and UO_2722 (O_2722,N_24895,N_24702);
xnor UO_2723 (O_2723,N_24869,N_24590);
nand UO_2724 (O_2724,N_24673,N_24752);
nor UO_2725 (O_2725,N_24927,N_24984);
nand UO_2726 (O_2726,N_24784,N_24830);
and UO_2727 (O_2727,N_24778,N_24639);
nor UO_2728 (O_2728,N_24755,N_24892);
nand UO_2729 (O_2729,N_24580,N_24730);
and UO_2730 (O_2730,N_24960,N_24993);
and UO_2731 (O_2731,N_24946,N_24788);
nor UO_2732 (O_2732,N_24926,N_24741);
and UO_2733 (O_2733,N_24739,N_24984);
or UO_2734 (O_2734,N_24816,N_24678);
nor UO_2735 (O_2735,N_24646,N_24909);
nand UO_2736 (O_2736,N_24879,N_24875);
nor UO_2737 (O_2737,N_24701,N_24584);
nor UO_2738 (O_2738,N_24620,N_24563);
or UO_2739 (O_2739,N_24961,N_24680);
nand UO_2740 (O_2740,N_24815,N_24755);
and UO_2741 (O_2741,N_24945,N_24533);
nand UO_2742 (O_2742,N_24874,N_24510);
or UO_2743 (O_2743,N_24812,N_24764);
nand UO_2744 (O_2744,N_24593,N_24696);
xnor UO_2745 (O_2745,N_24988,N_24704);
nand UO_2746 (O_2746,N_24909,N_24790);
xnor UO_2747 (O_2747,N_24680,N_24914);
and UO_2748 (O_2748,N_24970,N_24884);
and UO_2749 (O_2749,N_24841,N_24566);
or UO_2750 (O_2750,N_24788,N_24781);
and UO_2751 (O_2751,N_24696,N_24526);
or UO_2752 (O_2752,N_24637,N_24936);
and UO_2753 (O_2753,N_24527,N_24708);
nand UO_2754 (O_2754,N_24814,N_24721);
and UO_2755 (O_2755,N_24626,N_24616);
nor UO_2756 (O_2756,N_24995,N_24729);
or UO_2757 (O_2757,N_24691,N_24623);
and UO_2758 (O_2758,N_24945,N_24502);
nor UO_2759 (O_2759,N_24678,N_24991);
and UO_2760 (O_2760,N_24771,N_24780);
or UO_2761 (O_2761,N_24782,N_24723);
and UO_2762 (O_2762,N_24957,N_24772);
nor UO_2763 (O_2763,N_24529,N_24724);
nor UO_2764 (O_2764,N_24678,N_24979);
or UO_2765 (O_2765,N_24813,N_24825);
nand UO_2766 (O_2766,N_24513,N_24593);
nor UO_2767 (O_2767,N_24775,N_24917);
xor UO_2768 (O_2768,N_24588,N_24536);
and UO_2769 (O_2769,N_24729,N_24521);
or UO_2770 (O_2770,N_24716,N_24618);
nor UO_2771 (O_2771,N_24742,N_24540);
nand UO_2772 (O_2772,N_24520,N_24506);
and UO_2773 (O_2773,N_24656,N_24601);
or UO_2774 (O_2774,N_24992,N_24971);
nand UO_2775 (O_2775,N_24662,N_24672);
and UO_2776 (O_2776,N_24579,N_24824);
xor UO_2777 (O_2777,N_24704,N_24684);
nor UO_2778 (O_2778,N_24816,N_24502);
or UO_2779 (O_2779,N_24608,N_24561);
and UO_2780 (O_2780,N_24757,N_24528);
nor UO_2781 (O_2781,N_24552,N_24799);
and UO_2782 (O_2782,N_24769,N_24580);
nand UO_2783 (O_2783,N_24506,N_24907);
nand UO_2784 (O_2784,N_24546,N_24678);
and UO_2785 (O_2785,N_24957,N_24792);
nand UO_2786 (O_2786,N_24771,N_24758);
nor UO_2787 (O_2787,N_24821,N_24872);
and UO_2788 (O_2788,N_24550,N_24786);
or UO_2789 (O_2789,N_24679,N_24579);
or UO_2790 (O_2790,N_24619,N_24942);
and UO_2791 (O_2791,N_24904,N_24990);
or UO_2792 (O_2792,N_24901,N_24635);
and UO_2793 (O_2793,N_24516,N_24991);
or UO_2794 (O_2794,N_24908,N_24967);
nor UO_2795 (O_2795,N_24685,N_24843);
nor UO_2796 (O_2796,N_24706,N_24976);
xor UO_2797 (O_2797,N_24730,N_24927);
nand UO_2798 (O_2798,N_24895,N_24574);
and UO_2799 (O_2799,N_24812,N_24899);
xnor UO_2800 (O_2800,N_24923,N_24871);
nand UO_2801 (O_2801,N_24656,N_24521);
and UO_2802 (O_2802,N_24618,N_24554);
and UO_2803 (O_2803,N_24770,N_24761);
or UO_2804 (O_2804,N_24672,N_24966);
or UO_2805 (O_2805,N_24975,N_24774);
nand UO_2806 (O_2806,N_24567,N_24826);
or UO_2807 (O_2807,N_24585,N_24770);
and UO_2808 (O_2808,N_24962,N_24926);
or UO_2809 (O_2809,N_24692,N_24616);
xnor UO_2810 (O_2810,N_24684,N_24628);
nand UO_2811 (O_2811,N_24559,N_24711);
nor UO_2812 (O_2812,N_24732,N_24861);
nor UO_2813 (O_2813,N_24866,N_24817);
nand UO_2814 (O_2814,N_24829,N_24601);
nor UO_2815 (O_2815,N_24638,N_24588);
nand UO_2816 (O_2816,N_24681,N_24616);
and UO_2817 (O_2817,N_24758,N_24988);
xor UO_2818 (O_2818,N_24771,N_24509);
nor UO_2819 (O_2819,N_24635,N_24927);
and UO_2820 (O_2820,N_24708,N_24528);
or UO_2821 (O_2821,N_24679,N_24510);
or UO_2822 (O_2822,N_24869,N_24824);
nor UO_2823 (O_2823,N_24945,N_24644);
xnor UO_2824 (O_2824,N_24761,N_24576);
nand UO_2825 (O_2825,N_24921,N_24875);
xnor UO_2826 (O_2826,N_24699,N_24666);
nand UO_2827 (O_2827,N_24572,N_24682);
nand UO_2828 (O_2828,N_24956,N_24669);
xor UO_2829 (O_2829,N_24680,N_24917);
nand UO_2830 (O_2830,N_24767,N_24611);
and UO_2831 (O_2831,N_24805,N_24553);
and UO_2832 (O_2832,N_24996,N_24839);
or UO_2833 (O_2833,N_24540,N_24971);
or UO_2834 (O_2834,N_24868,N_24903);
or UO_2835 (O_2835,N_24758,N_24666);
nand UO_2836 (O_2836,N_24795,N_24958);
or UO_2837 (O_2837,N_24852,N_24694);
xor UO_2838 (O_2838,N_24619,N_24727);
nor UO_2839 (O_2839,N_24709,N_24897);
nand UO_2840 (O_2840,N_24768,N_24819);
and UO_2841 (O_2841,N_24927,N_24514);
nand UO_2842 (O_2842,N_24705,N_24622);
nor UO_2843 (O_2843,N_24599,N_24568);
nor UO_2844 (O_2844,N_24959,N_24597);
or UO_2845 (O_2845,N_24867,N_24602);
nand UO_2846 (O_2846,N_24976,N_24838);
nor UO_2847 (O_2847,N_24545,N_24991);
nor UO_2848 (O_2848,N_24926,N_24977);
nand UO_2849 (O_2849,N_24783,N_24838);
and UO_2850 (O_2850,N_24520,N_24939);
nor UO_2851 (O_2851,N_24626,N_24586);
nand UO_2852 (O_2852,N_24955,N_24845);
nand UO_2853 (O_2853,N_24946,N_24899);
or UO_2854 (O_2854,N_24820,N_24673);
nor UO_2855 (O_2855,N_24515,N_24988);
and UO_2856 (O_2856,N_24643,N_24884);
xnor UO_2857 (O_2857,N_24734,N_24984);
and UO_2858 (O_2858,N_24766,N_24995);
nand UO_2859 (O_2859,N_24876,N_24634);
nand UO_2860 (O_2860,N_24805,N_24832);
or UO_2861 (O_2861,N_24902,N_24954);
nor UO_2862 (O_2862,N_24905,N_24768);
nor UO_2863 (O_2863,N_24594,N_24813);
nand UO_2864 (O_2864,N_24518,N_24758);
nor UO_2865 (O_2865,N_24951,N_24520);
or UO_2866 (O_2866,N_24722,N_24963);
or UO_2867 (O_2867,N_24552,N_24587);
or UO_2868 (O_2868,N_24823,N_24775);
xnor UO_2869 (O_2869,N_24538,N_24677);
nand UO_2870 (O_2870,N_24893,N_24550);
xnor UO_2871 (O_2871,N_24856,N_24915);
nand UO_2872 (O_2872,N_24629,N_24535);
nor UO_2873 (O_2873,N_24500,N_24945);
nor UO_2874 (O_2874,N_24624,N_24765);
nand UO_2875 (O_2875,N_24986,N_24948);
and UO_2876 (O_2876,N_24989,N_24718);
nand UO_2877 (O_2877,N_24515,N_24558);
or UO_2878 (O_2878,N_24692,N_24838);
nand UO_2879 (O_2879,N_24556,N_24770);
or UO_2880 (O_2880,N_24596,N_24749);
and UO_2881 (O_2881,N_24877,N_24548);
nor UO_2882 (O_2882,N_24642,N_24565);
or UO_2883 (O_2883,N_24627,N_24600);
and UO_2884 (O_2884,N_24769,N_24663);
or UO_2885 (O_2885,N_24889,N_24787);
or UO_2886 (O_2886,N_24872,N_24565);
xor UO_2887 (O_2887,N_24751,N_24509);
xor UO_2888 (O_2888,N_24566,N_24736);
nand UO_2889 (O_2889,N_24777,N_24973);
or UO_2890 (O_2890,N_24884,N_24587);
and UO_2891 (O_2891,N_24691,N_24534);
or UO_2892 (O_2892,N_24758,N_24820);
xnor UO_2893 (O_2893,N_24820,N_24666);
nor UO_2894 (O_2894,N_24608,N_24705);
nor UO_2895 (O_2895,N_24693,N_24897);
and UO_2896 (O_2896,N_24528,N_24510);
nor UO_2897 (O_2897,N_24677,N_24506);
nor UO_2898 (O_2898,N_24946,N_24738);
or UO_2899 (O_2899,N_24769,N_24508);
nor UO_2900 (O_2900,N_24915,N_24531);
nor UO_2901 (O_2901,N_24526,N_24815);
xnor UO_2902 (O_2902,N_24583,N_24505);
nor UO_2903 (O_2903,N_24551,N_24564);
nor UO_2904 (O_2904,N_24893,N_24985);
nand UO_2905 (O_2905,N_24948,N_24718);
nand UO_2906 (O_2906,N_24975,N_24567);
and UO_2907 (O_2907,N_24888,N_24947);
or UO_2908 (O_2908,N_24541,N_24991);
nor UO_2909 (O_2909,N_24808,N_24515);
and UO_2910 (O_2910,N_24766,N_24804);
and UO_2911 (O_2911,N_24902,N_24845);
nand UO_2912 (O_2912,N_24521,N_24710);
and UO_2913 (O_2913,N_24952,N_24855);
nor UO_2914 (O_2914,N_24763,N_24878);
nand UO_2915 (O_2915,N_24531,N_24935);
or UO_2916 (O_2916,N_24902,N_24694);
nor UO_2917 (O_2917,N_24732,N_24735);
and UO_2918 (O_2918,N_24976,N_24780);
nand UO_2919 (O_2919,N_24762,N_24658);
xnor UO_2920 (O_2920,N_24642,N_24940);
or UO_2921 (O_2921,N_24549,N_24968);
nand UO_2922 (O_2922,N_24566,N_24898);
nand UO_2923 (O_2923,N_24670,N_24938);
and UO_2924 (O_2924,N_24866,N_24583);
nor UO_2925 (O_2925,N_24783,N_24982);
or UO_2926 (O_2926,N_24845,N_24557);
nand UO_2927 (O_2927,N_24801,N_24948);
and UO_2928 (O_2928,N_24622,N_24787);
nand UO_2929 (O_2929,N_24711,N_24959);
nor UO_2930 (O_2930,N_24930,N_24543);
or UO_2931 (O_2931,N_24907,N_24909);
xnor UO_2932 (O_2932,N_24567,N_24549);
xnor UO_2933 (O_2933,N_24876,N_24508);
xor UO_2934 (O_2934,N_24590,N_24565);
or UO_2935 (O_2935,N_24611,N_24511);
or UO_2936 (O_2936,N_24738,N_24602);
nor UO_2937 (O_2937,N_24529,N_24956);
nor UO_2938 (O_2938,N_24970,N_24931);
or UO_2939 (O_2939,N_24623,N_24905);
or UO_2940 (O_2940,N_24935,N_24793);
nand UO_2941 (O_2941,N_24839,N_24691);
or UO_2942 (O_2942,N_24560,N_24727);
and UO_2943 (O_2943,N_24966,N_24595);
xor UO_2944 (O_2944,N_24799,N_24929);
nor UO_2945 (O_2945,N_24565,N_24724);
xor UO_2946 (O_2946,N_24702,N_24638);
and UO_2947 (O_2947,N_24650,N_24672);
nand UO_2948 (O_2948,N_24864,N_24794);
and UO_2949 (O_2949,N_24685,N_24758);
or UO_2950 (O_2950,N_24603,N_24991);
and UO_2951 (O_2951,N_24860,N_24954);
nor UO_2952 (O_2952,N_24812,N_24623);
or UO_2953 (O_2953,N_24738,N_24827);
and UO_2954 (O_2954,N_24586,N_24938);
and UO_2955 (O_2955,N_24870,N_24813);
or UO_2956 (O_2956,N_24999,N_24611);
or UO_2957 (O_2957,N_24584,N_24598);
nor UO_2958 (O_2958,N_24878,N_24772);
or UO_2959 (O_2959,N_24587,N_24542);
nor UO_2960 (O_2960,N_24818,N_24565);
or UO_2961 (O_2961,N_24869,N_24513);
nor UO_2962 (O_2962,N_24851,N_24535);
nor UO_2963 (O_2963,N_24969,N_24772);
nand UO_2964 (O_2964,N_24819,N_24579);
or UO_2965 (O_2965,N_24819,N_24970);
xnor UO_2966 (O_2966,N_24865,N_24552);
nand UO_2967 (O_2967,N_24733,N_24918);
nand UO_2968 (O_2968,N_24654,N_24655);
and UO_2969 (O_2969,N_24987,N_24945);
nor UO_2970 (O_2970,N_24926,N_24740);
nor UO_2971 (O_2971,N_24510,N_24739);
nor UO_2972 (O_2972,N_24992,N_24749);
and UO_2973 (O_2973,N_24771,N_24566);
nor UO_2974 (O_2974,N_24744,N_24972);
or UO_2975 (O_2975,N_24826,N_24685);
or UO_2976 (O_2976,N_24757,N_24501);
nor UO_2977 (O_2977,N_24500,N_24818);
nor UO_2978 (O_2978,N_24893,N_24690);
xnor UO_2979 (O_2979,N_24694,N_24555);
or UO_2980 (O_2980,N_24770,N_24625);
nor UO_2981 (O_2981,N_24886,N_24851);
nand UO_2982 (O_2982,N_24552,N_24626);
nor UO_2983 (O_2983,N_24656,N_24826);
nor UO_2984 (O_2984,N_24795,N_24883);
or UO_2985 (O_2985,N_24626,N_24804);
nand UO_2986 (O_2986,N_24570,N_24693);
nor UO_2987 (O_2987,N_24861,N_24948);
nor UO_2988 (O_2988,N_24620,N_24790);
or UO_2989 (O_2989,N_24893,N_24995);
nor UO_2990 (O_2990,N_24611,N_24537);
and UO_2991 (O_2991,N_24986,N_24844);
nand UO_2992 (O_2992,N_24791,N_24632);
nor UO_2993 (O_2993,N_24852,N_24698);
or UO_2994 (O_2994,N_24573,N_24553);
nor UO_2995 (O_2995,N_24708,N_24695);
or UO_2996 (O_2996,N_24638,N_24521);
xor UO_2997 (O_2997,N_24796,N_24691);
nand UO_2998 (O_2998,N_24793,N_24956);
nand UO_2999 (O_2999,N_24968,N_24919);
endmodule