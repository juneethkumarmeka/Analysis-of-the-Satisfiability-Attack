module basic_500_3000_500_6_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_143,In_19);
nor U1 (N_1,In_237,In_108);
xor U2 (N_2,In_21,In_418);
and U3 (N_3,In_227,In_252);
nand U4 (N_4,In_469,In_359);
xor U5 (N_5,In_460,In_385);
nor U6 (N_6,In_56,In_485);
or U7 (N_7,In_4,In_24);
and U8 (N_8,In_194,In_284);
nor U9 (N_9,In_78,In_303);
and U10 (N_10,In_333,In_64);
xor U11 (N_11,In_435,In_294);
or U12 (N_12,In_457,In_126);
xnor U13 (N_13,In_90,In_258);
and U14 (N_14,In_100,In_117);
nor U15 (N_15,In_449,In_106);
or U16 (N_16,In_323,In_115);
xnor U17 (N_17,In_215,In_436);
and U18 (N_18,In_162,In_13);
nand U19 (N_19,In_369,In_132);
nor U20 (N_20,In_244,In_79);
or U21 (N_21,In_142,In_38);
and U22 (N_22,In_343,In_380);
nor U23 (N_23,In_297,In_494);
and U24 (N_24,In_482,In_468);
nor U25 (N_25,In_352,In_116);
xnor U26 (N_26,In_39,In_193);
nand U27 (N_27,In_170,In_372);
nor U28 (N_28,In_40,In_392);
nor U29 (N_29,In_61,In_319);
nand U30 (N_30,In_486,In_381);
nand U31 (N_31,In_20,In_83);
nand U32 (N_32,In_42,In_487);
and U33 (N_33,In_110,In_253);
or U34 (N_34,In_285,In_10);
or U35 (N_35,In_27,In_17);
and U36 (N_36,In_80,In_107);
or U37 (N_37,In_238,In_483);
nand U38 (N_38,In_348,In_339);
or U39 (N_39,In_277,In_85);
nand U40 (N_40,In_270,In_12);
nand U41 (N_41,In_321,In_497);
nand U42 (N_42,In_28,In_18);
or U43 (N_43,In_186,In_300);
or U44 (N_44,In_188,In_361);
nand U45 (N_45,In_37,In_423);
nand U46 (N_46,In_488,In_440);
nor U47 (N_47,In_311,In_416);
or U48 (N_48,In_394,In_0);
xnor U49 (N_49,In_474,In_57);
and U50 (N_50,In_223,In_140);
nand U51 (N_51,In_125,In_96);
nor U52 (N_52,In_130,In_426);
nand U53 (N_53,In_211,In_328);
or U54 (N_54,In_478,In_137);
xnor U55 (N_55,In_456,In_174);
xor U56 (N_56,In_357,In_172);
and U57 (N_57,In_371,In_113);
nor U58 (N_58,In_31,In_280);
nor U59 (N_59,In_322,In_324);
xor U60 (N_60,In_293,In_60);
xnor U61 (N_61,In_59,In_199);
or U62 (N_62,In_16,In_414);
xnor U63 (N_63,In_35,In_23);
nor U64 (N_64,In_93,In_5);
nor U65 (N_65,In_119,In_289);
nand U66 (N_66,In_171,In_152);
nand U67 (N_67,In_329,In_213);
or U68 (N_68,In_264,In_81);
nand U69 (N_69,In_232,In_43);
and U70 (N_70,In_221,In_434);
and U71 (N_71,In_287,In_376);
nand U72 (N_72,In_439,In_206);
nor U73 (N_73,In_209,In_356);
xnor U74 (N_74,In_459,In_66);
nor U75 (N_75,In_160,In_347);
xnor U76 (N_76,In_72,In_127);
nor U77 (N_77,In_58,In_427);
nor U78 (N_78,In_76,In_387);
nor U79 (N_79,In_46,In_175);
nand U80 (N_80,In_204,In_354);
or U81 (N_81,In_455,In_48);
and U82 (N_82,In_216,In_362);
xnor U83 (N_83,In_442,In_95);
nand U84 (N_84,In_370,In_453);
or U85 (N_85,In_476,In_30);
nor U86 (N_86,In_262,In_308);
and U87 (N_87,In_139,In_114);
nand U88 (N_88,In_377,In_67);
or U89 (N_89,In_71,In_399);
xnor U90 (N_90,In_393,In_86);
or U91 (N_91,In_181,In_379);
or U92 (N_92,In_250,In_34);
and U93 (N_93,In_411,In_458);
or U94 (N_94,In_136,In_92);
and U95 (N_95,In_446,In_334);
nand U96 (N_96,In_298,In_307);
nor U97 (N_97,In_197,In_6);
or U98 (N_98,In_150,In_169);
nor U99 (N_99,In_274,In_91);
and U100 (N_100,In_97,In_296);
xnor U101 (N_101,In_254,In_184);
or U102 (N_102,In_317,In_424);
or U103 (N_103,In_384,In_350);
or U104 (N_104,In_438,In_401);
xor U105 (N_105,In_290,In_326);
or U106 (N_106,In_178,In_164);
nor U107 (N_107,In_452,In_331);
and U108 (N_108,In_9,In_217);
xor U109 (N_109,In_220,In_383);
nand U110 (N_110,In_112,In_475);
nand U111 (N_111,In_261,In_69);
or U112 (N_112,In_367,In_2);
nor U113 (N_113,In_295,In_187);
nand U114 (N_114,In_498,In_11);
nand U115 (N_115,In_208,In_49);
nand U116 (N_116,In_242,In_149);
or U117 (N_117,In_433,In_443);
or U118 (N_118,In_395,In_88);
or U119 (N_119,In_465,In_25);
nand U120 (N_120,In_226,In_281);
nand U121 (N_121,In_473,In_183);
or U122 (N_122,In_398,In_70);
and U123 (N_123,In_121,In_282);
xor U124 (N_124,In_306,In_413);
or U125 (N_125,In_233,In_120);
or U126 (N_126,In_266,In_207);
or U127 (N_127,In_240,In_366);
nor U128 (N_128,In_153,In_405);
xor U129 (N_129,In_309,In_145);
nor U130 (N_130,In_421,In_415);
or U131 (N_131,In_1,In_180);
nand U132 (N_132,In_490,In_299);
and U133 (N_133,In_73,In_77);
nor U134 (N_134,In_163,In_463);
and U135 (N_135,In_340,In_15);
or U136 (N_136,In_26,In_431);
or U137 (N_137,In_271,In_391);
and U138 (N_138,In_396,In_353);
nor U139 (N_139,In_41,In_336);
nand U140 (N_140,In_315,In_467);
or U141 (N_141,In_466,In_246);
nand U142 (N_142,In_386,In_65);
nor U143 (N_143,In_103,In_190);
nor U144 (N_144,In_355,In_173);
nand U145 (N_145,In_241,In_330);
or U146 (N_146,In_243,In_68);
and U147 (N_147,In_291,In_288);
nand U148 (N_148,In_364,In_410);
or U149 (N_149,In_202,In_176);
nor U150 (N_150,In_346,In_144);
and U151 (N_151,In_256,In_55);
nand U152 (N_152,In_400,In_337);
nand U153 (N_153,In_146,In_419);
and U154 (N_154,In_236,In_159);
and U155 (N_155,In_138,In_420);
nand U156 (N_156,In_259,In_109);
and U157 (N_157,In_363,In_52);
or U158 (N_158,In_229,In_345);
nand U159 (N_159,In_47,In_304);
and U160 (N_160,In_429,In_445);
nand U161 (N_161,In_218,In_477);
nand U162 (N_162,In_8,In_156);
xnor U163 (N_163,In_255,In_320);
and U164 (N_164,In_374,In_462);
nor U165 (N_165,In_332,In_74);
nand U166 (N_166,In_491,In_407);
and U167 (N_167,In_368,In_135);
nor U168 (N_168,In_484,In_260);
and U169 (N_169,In_245,In_404);
xor U170 (N_170,In_129,In_200);
xnor U171 (N_171,In_118,In_235);
nor U172 (N_172,In_192,In_402);
xor U173 (N_173,In_33,In_87);
and U174 (N_174,In_316,In_406);
and U175 (N_175,In_189,In_177);
xor U176 (N_176,In_104,In_257);
nand U177 (N_177,In_151,In_45);
or U178 (N_178,In_157,In_335);
nor U179 (N_179,In_122,In_373);
or U180 (N_180,In_481,In_276);
or U181 (N_181,In_239,In_283);
or U182 (N_182,In_408,In_447);
xor U183 (N_183,In_249,In_210);
nor U184 (N_184,In_279,In_480);
xor U185 (N_185,In_32,In_417);
or U186 (N_186,In_205,In_148);
or U187 (N_187,In_472,In_349);
or U188 (N_188,In_212,In_185);
nand U189 (N_189,In_313,In_50);
or U190 (N_190,In_286,In_451);
nor U191 (N_191,In_430,In_147);
xnor U192 (N_192,In_251,In_231);
nor U193 (N_193,In_432,In_195);
or U194 (N_194,In_29,In_166);
and U195 (N_195,In_36,In_168);
xnor U196 (N_196,In_44,In_305);
and U197 (N_197,In_247,In_214);
and U198 (N_198,In_448,In_75);
and U199 (N_199,In_464,In_388);
nand U200 (N_200,In_167,In_248);
and U201 (N_201,In_428,In_128);
nand U202 (N_202,In_89,In_123);
nor U203 (N_203,In_437,In_365);
or U204 (N_204,In_131,In_318);
or U205 (N_205,In_94,In_224);
and U206 (N_206,In_302,In_63);
nor U207 (N_207,In_219,In_155);
or U208 (N_208,In_22,In_182);
nor U209 (N_209,In_111,In_158);
and U210 (N_210,In_338,In_310);
nor U211 (N_211,In_351,In_272);
nor U212 (N_212,In_495,In_360);
or U213 (N_213,In_124,In_325);
xnor U214 (N_214,In_191,In_496);
nand U215 (N_215,In_461,In_7);
and U216 (N_216,In_450,In_493);
xor U217 (N_217,In_470,In_422);
nor U218 (N_218,In_269,In_82);
and U219 (N_219,In_389,In_196);
or U220 (N_220,In_425,In_341);
nand U221 (N_221,In_382,In_327);
or U222 (N_222,In_312,In_273);
xor U223 (N_223,In_105,In_134);
nand U224 (N_224,In_141,In_265);
and U225 (N_225,In_489,In_198);
nor U226 (N_226,In_292,In_278);
nor U227 (N_227,In_161,In_479);
and U228 (N_228,In_412,In_441);
nor U229 (N_229,In_444,In_301);
and U230 (N_230,In_344,In_222);
and U231 (N_231,In_101,In_201);
nand U232 (N_232,In_234,In_133);
nand U233 (N_233,In_267,In_99);
and U234 (N_234,In_53,In_228);
and U235 (N_235,In_342,In_14);
and U236 (N_236,In_390,In_225);
nand U237 (N_237,In_378,In_471);
nand U238 (N_238,In_165,In_230);
or U239 (N_239,In_102,In_179);
or U240 (N_240,In_62,In_84);
nand U241 (N_241,In_154,In_54);
and U242 (N_242,In_492,In_314);
nor U243 (N_243,In_499,In_454);
nand U244 (N_244,In_409,In_397);
and U245 (N_245,In_275,In_375);
nor U246 (N_246,In_268,In_403);
and U247 (N_247,In_263,In_51);
and U248 (N_248,In_3,In_203);
xnor U249 (N_249,In_98,In_358);
nand U250 (N_250,In_120,In_462);
nor U251 (N_251,In_205,In_51);
nand U252 (N_252,In_276,In_126);
or U253 (N_253,In_215,In_342);
and U254 (N_254,In_457,In_441);
xor U255 (N_255,In_357,In_14);
xnor U256 (N_256,In_469,In_319);
xor U257 (N_257,In_63,In_325);
or U258 (N_258,In_210,In_365);
nor U259 (N_259,In_67,In_484);
or U260 (N_260,In_173,In_47);
and U261 (N_261,In_308,In_399);
or U262 (N_262,In_202,In_487);
and U263 (N_263,In_369,In_349);
or U264 (N_264,In_434,In_224);
nor U265 (N_265,In_316,In_128);
and U266 (N_266,In_168,In_465);
and U267 (N_267,In_358,In_355);
xnor U268 (N_268,In_459,In_411);
nor U269 (N_269,In_298,In_252);
nand U270 (N_270,In_356,In_11);
or U271 (N_271,In_499,In_117);
and U272 (N_272,In_398,In_98);
nand U273 (N_273,In_243,In_433);
xor U274 (N_274,In_36,In_397);
and U275 (N_275,In_191,In_255);
nor U276 (N_276,In_115,In_403);
or U277 (N_277,In_419,In_52);
and U278 (N_278,In_368,In_228);
nand U279 (N_279,In_348,In_245);
or U280 (N_280,In_288,In_137);
nor U281 (N_281,In_142,In_292);
and U282 (N_282,In_108,In_114);
xnor U283 (N_283,In_187,In_107);
or U284 (N_284,In_320,In_275);
and U285 (N_285,In_405,In_370);
or U286 (N_286,In_211,In_317);
and U287 (N_287,In_165,In_149);
or U288 (N_288,In_452,In_203);
nand U289 (N_289,In_312,In_230);
or U290 (N_290,In_304,In_475);
or U291 (N_291,In_443,In_414);
or U292 (N_292,In_359,In_195);
nand U293 (N_293,In_272,In_459);
nand U294 (N_294,In_200,In_183);
and U295 (N_295,In_417,In_13);
or U296 (N_296,In_94,In_306);
nand U297 (N_297,In_178,In_296);
nand U298 (N_298,In_419,In_108);
nand U299 (N_299,In_164,In_127);
and U300 (N_300,In_433,In_377);
and U301 (N_301,In_363,In_206);
nand U302 (N_302,In_83,In_58);
xnor U303 (N_303,In_370,In_0);
and U304 (N_304,In_299,In_42);
and U305 (N_305,In_107,In_250);
nand U306 (N_306,In_255,In_55);
or U307 (N_307,In_431,In_149);
and U308 (N_308,In_404,In_199);
nor U309 (N_309,In_104,In_334);
or U310 (N_310,In_345,In_383);
and U311 (N_311,In_144,In_175);
or U312 (N_312,In_472,In_133);
nand U313 (N_313,In_476,In_237);
nand U314 (N_314,In_9,In_393);
and U315 (N_315,In_413,In_246);
nand U316 (N_316,In_312,In_432);
nor U317 (N_317,In_212,In_395);
and U318 (N_318,In_318,In_435);
nand U319 (N_319,In_69,In_337);
nor U320 (N_320,In_270,In_451);
or U321 (N_321,In_239,In_213);
nor U322 (N_322,In_323,In_25);
nand U323 (N_323,In_408,In_236);
or U324 (N_324,In_49,In_201);
xor U325 (N_325,In_64,In_27);
xnor U326 (N_326,In_51,In_232);
and U327 (N_327,In_421,In_144);
and U328 (N_328,In_242,In_384);
nand U329 (N_329,In_439,In_428);
or U330 (N_330,In_266,In_245);
nand U331 (N_331,In_148,In_274);
nor U332 (N_332,In_1,In_405);
nand U333 (N_333,In_390,In_214);
nand U334 (N_334,In_51,In_13);
or U335 (N_335,In_21,In_433);
nor U336 (N_336,In_23,In_282);
and U337 (N_337,In_151,In_464);
nand U338 (N_338,In_404,In_243);
and U339 (N_339,In_44,In_156);
or U340 (N_340,In_98,In_36);
xnor U341 (N_341,In_454,In_226);
or U342 (N_342,In_203,In_463);
nand U343 (N_343,In_478,In_452);
nor U344 (N_344,In_336,In_377);
or U345 (N_345,In_46,In_181);
nand U346 (N_346,In_115,In_334);
and U347 (N_347,In_312,In_83);
nor U348 (N_348,In_147,In_95);
and U349 (N_349,In_499,In_290);
and U350 (N_350,In_371,In_161);
or U351 (N_351,In_178,In_285);
xnor U352 (N_352,In_440,In_198);
and U353 (N_353,In_14,In_429);
nor U354 (N_354,In_76,In_417);
nand U355 (N_355,In_420,In_96);
nor U356 (N_356,In_307,In_322);
nand U357 (N_357,In_207,In_427);
or U358 (N_358,In_414,In_173);
nor U359 (N_359,In_432,In_302);
nor U360 (N_360,In_472,In_237);
nor U361 (N_361,In_263,In_52);
and U362 (N_362,In_220,In_130);
and U363 (N_363,In_36,In_307);
or U364 (N_364,In_483,In_473);
nor U365 (N_365,In_196,In_486);
nor U366 (N_366,In_205,In_152);
or U367 (N_367,In_103,In_109);
and U368 (N_368,In_433,In_352);
or U369 (N_369,In_280,In_64);
and U370 (N_370,In_234,In_94);
nand U371 (N_371,In_225,In_53);
nor U372 (N_372,In_44,In_98);
nor U373 (N_373,In_266,In_331);
nand U374 (N_374,In_268,In_111);
and U375 (N_375,In_193,In_14);
xor U376 (N_376,In_352,In_330);
nand U377 (N_377,In_64,In_256);
xor U378 (N_378,In_190,In_352);
and U379 (N_379,In_123,In_20);
nor U380 (N_380,In_132,In_162);
nor U381 (N_381,In_107,In_363);
or U382 (N_382,In_467,In_483);
xor U383 (N_383,In_355,In_210);
xor U384 (N_384,In_424,In_151);
xor U385 (N_385,In_77,In_299);
and U386 (N_386,In_84,In_440);
nand U387 (N_387,In_329,In_292);
nor U388 (N_388,In_214,In_127);
nor U389 (N_389,In_202,In_405);
or U390 (N_390,In_297,In_163);
or U391 (N_391,In_461,In_211);
or U392 (N_392,In_386,In_499);
nor U393 (N_393,In_468,In_473);
nand U394 (N_394,In_130,In_454);
or U395 (N_395,In_41,In_297);
nand U396 (N_396,In_28,In_104);
and U397 (N_397,In_459,In_258);
xor U398 (N_398,In_387,In_80);
or U399 (N_399,In_211,In_339);
xnor U400 (N_400,In_3,In_129);
nand U401 (N_401,In_39,In_27);
nor U402 (N_402,In_357,In_18);
nor U403 (N_403,In_278,In_478);
xor U404 (N_404,In_409,In_236);
or U405 (N_405,In_455,In_87);
or U406 (N_406,In_242,In_50);
xor U407 (N_407,In_94,In_296);
and U408 (N_408,In_478,In_252);
or U409 (N_409,In_365,In_92);
or U410 (N_410,In_327,In_491);
xor U411 (N_411,In_374,In_484);
or U412 (N_412,In_453,In_14);
and U413 (N_413,In_452,In_244);
or U414 (N_414,In_8,In_110);
xnor U415 (N_415,In_82,In_30);
and U416 (N_416,In_457,In_181);
or U417 (N_417,In_347,In_442);
nand U418 (N_418,In_355,In_300);
or U419 (N_419,In_88,In_402);
nor U420 (N_420,In_30,In_356);
or U421 (N_421,In_177,In_51);
xor U422 (N_422,In_196,In_189);
nand U423 (N_423,In_120,In_138);
and U424 (N_424,In_234,In_177);
and U425 (N_425,In_476,In_363);
nand U426 (N_426,In_67,In_483);
and U427 (N_427,In_183,In_38);
nor U428 (N_428,In_402,In_105);
nand U429 (N_429,In_477,In_356);
nor U430 (N_430,In_402,In_15);
nand U431 (N_431,In_487,In_196);
nor U432 (N_432,In_277,In_263);
xor U433 (N_433,In_321,In_114);
and U434 (N_434,In_116,In_254);
or U435 (N_435,In_36,In_214);
nor U436 (N_436,In_206,In_292);
and U437 (N_437,In_258,In_273);
xnor U438 (N_438,In_277,In_39);
nor U439 (N_439,In_52,In_197);
nand U440 (N_440,In_87,In_308);
or U441 (N_441,In_359,In_494);
nand U442 (N_442,In_387,In_180);
or U443 (N_443,In_402,In_147);
nor U444 (N_444,In_3,In_467);
or U445 (N_445,In_137,In_381);
or U446 (N_446,In_194,In_437);
or U447 (N_447,In_216,In_291);
nor U448 (N_448,In_226,In_65);
or U449 (N_449,In_112,In_458);
or U450 (N_450,In_369,In_144);
or U451 (N_451,In_90,In_216);
nand U452 (N_452,In_303,In_311);
or U453 (N_453,In_141,In_317);
xor U454 (N_454,In_183,In_215);
or U455 (N_455,In_452,In_260);
nand U456 (N_456,In_269,In_136);
nor U457 (N_457,In_361,In_303);
and U458 (N_458,In_121,In_90);
nand U459 (N_459,In_148,In_228);
and U460 (N_460,In_471,In_115);
nor U461 (N_461,In_205,In_428);
nand U462 (N_462,In_302,In_452);
nand U463 (N_463,In_69,In_107);
and U464 (N_464,In_38,In_284);
or U465 (N_465,In_58,In_136);
and U466 (N_466,In_486,In_67);
or U467 (N_467,In_437,In_49);
nor U468 (N_468,In_348,In_224);
or U469 (N_469,In_258,In_366);
and U470 (N_470,In_219,In_343);
or U471 (N_471,In_99,In_466);
or U472 (N_472,In_95,In_166);
nand U473 (N_473,In_423,In_251);
xor U474 (N_474,In_383,In_278);
or U475 (N_475,In_429,In_36);
or U476 (N_476,In_46,In_398);
nand U477 (N_477,In_476,In_172);
nor U478 (N_478,In_144,In_138);
nor U479 (N_479,In_271,In_132);
nand U480 (N_480,In_415,In_57);
nand U481 (N_481,In_98,In_8);
or U482 (N_482,In_59,In_234);
nor U483 (N_483,In_130,In_15);
and U484 (N_484,In_343,In_103);
or U485 (N_485,In_204,In_105);
nand U486 (N_486,In_266,In_268);
xor U487 (N_487,In_220,In_239);
nor U488 (N_488,In_348,In_109);
xnor U489 (N_489,In_261,In_216);
nor U490 (N_490,In_397,In_148);
nand U491 (N_491,In_467,In_499);
and U492 (N_492,In_188,In_161);
nand U493 (N_493,In_183,In_106);
nand U494 (N_494,In_178,In_350);
nor U495 (N_495,In_69,In_120);
or U496 (N_496,In_31,In_222);
nand U497 (N_497,In_178,In_122);
or U498 (N_498,In_64,In_474);
nor U499 (N_499,In_400,In_471);
and U500 (N_500,N_97,N_147);
xor U501 (N_501,N_398,N_123);
nand U502 (N_502,N_391,N_446);
or U503 (N_503,N_247,N_171);
nand U504 (N_504,N_331,N_357);
or U505 (N_505,N_22,N_176);
nand U506 (N_506,N_134,N_328);
and U507 (N_507,N_33,N_237);
nand U508 (N_508,N_89,N_369);
or U509 (N_509,N_58,N_196);
nand U510 (N_510,N_379,N_81);
or U511 (N_511,N_35,N_359);
xor U512 (N_512,N_309,N_169);
and U513 (N_513,N_343,N_71);
and U514 (N_514,N_349,N_469);
xnor U515 (N_515,N_430,N_300);
or U516 (N_516,N_73,N_318);
nand U517 (N_517,N_383,N_117);
xnor U518 (N_518,N_222,N_76);
nand U519 (N_519,N_385,N_184);
xnor U520 (N_520,N_185,N_473);
or U521 (N_521,N_387,N_397);
nor U522 (N_522,N_307,N_198);
nand U523 (N_523,N_396,N_354);
nor U524 (N_524,N_101,N_288);
nand U525 (N_525,N_182,N_201);
and U526 (N_526,N_461,N_295);
and U527 (N_527,N_294,N_94);
nand U528 (N_528,N_130,N_297);
nand U529 (N_529,N_28,N_374);
or U530 (N_530,N_50,N_141);
xnor U531 (N_531,N_395,N_137);
and U532 (N_532,N_335,N_488);
or U533 (N_533,N_353,N_450);
and U534 (N_534,N_301,N_104);
nand U535 (N_535,N_421,N_191);
nand U536 (N_536,N_166,N_437);
xnor U537 (N_537,N_41,N_484);
nand U538 (N_538,N_20,N_471);
and U539 (N_539,N_240,N_106);
nand U540 (N_540,N_313,N_490);
nor U541 (N_541,N_13,N_116);
nand U542 (N_542,N_0,N_333);
nor U543 (N_543,N_95,N_175);
or U544 (N_544,N_87,N_299);
nand U545 (N_545,N_355,N_377);
nand U546 (N_546,N_161,N_75);
xor U547 (N_547,N_142,N_212);
nand U548 (N_548,N_495,N_216);
nand U549 (N_549,N_316,N_485);
nor U550 (N_550,N_466,N_146);
nor U551 (N_551,N_246,N_2);
nand U552 (N_552,N_483,N_168);
and U553 (N_553,N_193,N_36);
xor U554 (N_554,N_467,N_152);
and U555 (N_555,N_48,N_443);
or U556 (N_556,N_39,N_157);
and U557 (N_557,N_497,N_428);
and U558 (N_558,N_454,N_350);
and U559 (N_559,N_144,N_177);
xor U560 (N_560,N_487,N_429);
nor U561 (N_561,N_17,N_389);
or U562 (N_562,N_348,N_90);
nand U563 (N_563,N_289,N_218);
nand U564 (N_564,N_179,N_435);
and U565 (N_565,N_274,N_40);
nor U566 (N_566,N_455,N_470);
nor U567 (N_567,N_432,N_125);
and U568 (N_568,N_227,N_7);
and U569 (N_569,N_108,N_463);
or U570 (N_570,N_21,N_111);
nor U571 (N_571,N_115,N_336);
and U572 (N_572,N_149,N_439);
nor U573 (N_573,N_415,N_252);
or U574 (N_574,N_105,N_59);
and U575 (N_575,N_329,N_405);
xor U576 (N_576,N_154,N_230);
nand U577 (N_577,N_314,N_189);
or U578 (N_578,N_213,N_478);
nand U579 (N_579,N_255,N_18);
nor U580 (N_580,N_244,N_165);
xor U581 (N_581,N_481,N_458);
or U582 (N_582,N_56,N_468);
nand U583 (N_583,N_31,N_225);
nor U584 (N_584,N_129,N_302);
and U585 (N_585,N_228,N_209);
or U586 (N_586,N_140,N_127);
or U587 (N_587,N_204,N_224);
and U588 (N_588,N_410,N_453);
nand U589 (N_589,N_205,N_464);
and U590 (N_590,N_107,N_30);
nand U591 (N_591,N_390,N_86);
and U592 (N_592,N_100,N_342);
nand U593 (N_593,N_386,N_339);
and U594 (N_594,N_474,N_11);
and U595 (N_595,N_411,N_164);
nand U596 (N_596,N_317,N_338);
or U597 (N_597,N_170,N_284);
nand U598 (N_598,N_372,N_298);
and U599 (N_599,N_358,N_235);
nor U600 (N_600,N_138,N_351);
nand U601 (N_601,N_283,N_188);
or U602 (N_602,N_214,N_53);
and U603 (N_603,N_187,N_434);
nor U604 (N_604,N_160,N_279);
xor U605 (N_605,N_438,N_256);
nor U606 (N_606,N_424,N_131);
nor U607 (N_607,N_99,N_126);
nor U608 (N_608,N_345,N_67);
nor U609 (N_609,N_47,N_186);
or U610 (N_610,N_239,N_273);
or U611 (N_611,N_211,N_475);
and U612 (N_612,N_311,N_57);
nand U613 (N_613,N_49,N_286);
or U614 (N_614,N_150,N_456);
nor U615 (N_615,N_234,N_148);
or U616 (N_616,N_489,N_32);
nor U617 (N_617,N_124,N_1);
nand U618 (N_618,N_414,N_406);
nor U619 (N_619,N_19,N_327);
or U620 (N_620,N_326,N_136);
and U621 (N_621,N_44,N_375);
nand U622 (N_622,N_324,N_420);
and U623 (N_623,N_180,N_442);
nand U624 (N_624,N_77,N_217);
or U625 (N_625,N_321,N_363);
or U626 (N_626,N_445,N_278);
nand U627 (N_627,N_323,N_308);
nor U628 (N_628,N_55,N_163);
nor U629 (N_629,N_480,N_479);
nor U630 (N_630,N_332,N_482);
nand U631 (N_631,N_400,N_269);
xnor U632 (N_632,N_210,N_14);
or U633 (N_633,N_296,N_291);
and U634 (N_634,N_96,N_3);
nor U635 (N_635,N_8,N_145);
or U636 (N_636,N_61,N_268);
nand U637 (N_637,N_356,N_413);
or U638 (N_638,N_208,N_371);
or U639 (N_639,N_259,N_407);
or U640 (N_640,N_26,N_194);
and U641 (N_641,N_380,N_9);
or U642 (N_642,N_465,N_121);
or U643 (N_643,N_72,N_404);
and U644 (N_644,N_93,N_496);
nor U645 (N_645,N_419,N_120);
or U646 (N_646,N_427,N_280);
nand U647 (N_647,N_325,N_452);
and U648 (N_648,N_320,N_236);
xnor U649 (N_649,N_203,N_63);
or U650 (N_650,N_366,N_394);
and U651 (N_651,N_277,N_6);
and U652 (N_652,N_114,N_346);
nand U653 (N_653,N_472,N_223);
or U654 (N_654,N_80,N_418);
nand U655 (N_655,N_221,N_376);
or U656 (N_656,N_233,N_98);
and U657 (N_657,N_493,N_181);
nand U658 (N_658,N_449,N_271);
nor U659 (N_659,N_368,N_436);
xnor U660 (N_660,N_392,N_287);
nor U661 (N_661,N_84,N_103);
or U662 (N_662,N_231,N_51);
or U663 (N_663,N_499,N_29);
nor U664 (N_664,N_282,N_315);
nand U665 (N_665,N_162,N_250);
nand U666 (N_666,N_352,N_293);
and U667 (N_667,N_242,N_85);
nand U668 (N_668,N_38,N_66);
or U669 (N_669,N_401,N_42);
or U670 (N_670,N_447,N_118);
or U671 (N_671,N_88,N_74);
nor U672 (N_672,N_462,N_334);
nand U673 (N_673,N_365,N_251);
nor U674 (N_674,N_370,N_498);
or U675 (N_675,N_276,N_69);
and U676 (N_676,N_10,N_70);
nor U677 (N_677,N_4,N_128);
or U678 (N_678,N_440,N_24);
and U679 (N_679,N_330,N_64);
and U680 (N_680,N_245,N_344);
xnor U681 (N_681,N_494,N_215);
or U682 (N_682,N_79,N_423);
and U683 (N_683,N_382,N_285);
or U684 (N_684,N_158,N_119);
xor U685 (N_685,N_143,N_229);
or U686 (N_686,N_249,N_78);
nor U687 (N_687,N_190,N_448);
nor U688 (N_688,N_27,N_425);
xnor U689 (N_689,N_486,N_457);
and U690 (N_690,N_207,N_172);
nor U691 (N_691,N_159,N_337);
nor U692 (N_692,N_82,N_347);
and U693 (N_693,N_409,N_304);
xnor U694 (N_694,N_270,N_167);
nor U695 (N_695,N_422,N_192);
xor U696 (N_696,N_281,N_206);
xnor U697 (N_697,N_477,N_305);
nor U698 (N_698,N_312,N_403);
xor U699 (N_699,N_367,N_340);
nor U700 (N_700,N_267,N_292);
xor U701 (N_701,N_220,N_361);
nand U702 (N_702,N_156,N_364);
or U703 (N_703,N_393,N_360);
or U704 (N_704,N_202,N_5);
nor U705 (N_705,N_253,N_112);
nor U706 (N_706,N_65,N_83);
or U707 (N_707,N_92,N_153);
nand U708 (N_708,N_381,N_476);
nand U709 (N_709,N_254,N_441);
nor U710 (N_710,N_341,N_257);
nor U711 (N_711,N_417,N_109);
nor U712 (N_712,N_460,N_43);
or U713 (N_713,N_110,N_37);
and U714 (N_714,N_306,N_408);
nand U715 (N_715,N_46,N_23);
and U716 (N_716,N_373,N_15);
or U717 (N_717,N_226,N_290);
or U718 (N_718,N_54,N_34);
nor U719 (N_719,N_200,N_272);
nor U720 (N_720,N_261,N_155);
and U721 (N_721,N_174,N_362);
nor U722 (N_722,N_491,N_262);
or U723 (N_723,N_402,N_433);
and U724 (N_724,N_60,N_52);
nand U725 (N_725,N_263,N_195);
nor U726 (N_726,N_303,N_62);
nor U727 (N_727,N_135,N_258);
nor U728 (N_728,N_16,N_412);
nand U729 (N_729,N_431,N_232);
or U730 (N_730,N_12,N_173);
nor U731 (N_731,N_444,N_219);
and U732 (N_732,N_265,N_388);
or U733 (N_733,N_151,N_113);
or U734 (N_734,N_264,N_45);
nor U735 (N_735,N_139,N_91);
nand U736 (N_736,N_199,N_275);
and U737 (N_737,N_260,N_122);
and U738 (N_738,N_451,N_197);
and U739 (N_739,N_178,N_266);
and U740 (N_740,N_378,N_102);
and U741 (N_741,N_68,N_241);
nand U742 (N_742,N_426,N_399);
nor U743 (N_743,N_248,N_310);
nand U744 (N_744,N_416,N_322);
nand U745 (N_745,N_243,N_183);
nand U746 (N_746,N_133,N_492);
and U747 (N_747,N_319,N_459);
nand U748 (N_748,N_25,N_132);
xor U749 (N_749,N_238,N_384);
nor U750 (N_750,N_443,N_361);
or U751 (N_751,N_79,N_466);
xor U752 (N_752,N_169,N_36);
or U753 (N_753,N_178,N_147);
and U754 (N_754,N_372,N_386);
or U755 (N_755,N_210,N_420);
nor U756 (N_756,N_455,N_163);
nand U757 (N_757,N_435,N_373);
or U758 (N_758,N_359,N_198);
and U759 (N_759,N_212,N_410);
or U760 (N_760,N_3,N_425);
or U761 (N_761,N_482,N_68);
nand U762 (N_762,N_484,N_409);
and U763 (N_763,N_115,N_99);
nor U764 (N_764,N_381,N_269);
and U765 (N_765,N_193,N_19);
or U766 (N_766,N_78,N_362);
and U767 (N_767,N_221,N_38);
nand U768 (N_768,N_225,N_426);
nor U769 (N_769,N_398,N_230);
and U770 (N_770,N_10,N_448);
and U771 (N_771,N_121,N_404);
nor U772 (N_772,N_311,N_213);
nand U773 (N_773,N_428,N_423);
and U774 (N_774,N_396,N_494);
nor U775 (N_775,N_313,N_119);
or U776 (N_776,N_155,N_497);
xor U777 (N_777,N_73,N_165);
nor U778 (N_778,N_209,N_130);
or U779 (N_779,N_446,N_463);
nor U780 (N_780,N_258,N_15);
nor U781 (N_781,N_315,N_460);
nand U782 (N_782,N_62,N_402);
nor U783 (N_783,N_19,N_185);
or U784 (N_784,N_279,N_71);
xnor U785 (N_785,N_367,N_482);
and U786 (N_786,N_456,N_312);
or U787 (N_787,N_96,N_72);
or U788 (N_788,N_365,N_488);
nand U789 (N_789,N_169,N_33);
and U790 (N_790,N_450,N_43);
or U791 (N_791,N_28,N_82);
nor U792 (N_792,N_438,N_356);
and U793 (N_793,N_242,N_110);
nand U794 (N_794,N_271,N_410);
or U795 (N_795,N_290,N_491);
nor U796 (N_796,N_10,N_8);
nor U797 (N_797,N_126,N_54);
nor U798 (N_798,N_127,N_490);
or U799 (N_799,N_280,N_67);
nand U800 (N_800,N_232,N_200);
nor U801 (N_801,N_478,N_462);
and U802 (N_802,N_295,N_233);
nor U803 (N_803,N_237,N_289);
nor U804 (N_804,N_488,N_172);
or U805 (N_805,N_181,N_192);
and U806 (N_806,N_124,N_221);
and U807 (N_807,N_376,N_322);
and U808 (N_808,N_438,N_14);
xnor U809 (N_809,N_163,N_230);
xnor U810 (N_810,N_239,N_338);
nor U811 (N_811,N_110,N_405);
and U812 (N_812,N_131,N_343);
xor U813 (N_813,N_389,N_8);
nand U814 (N_814,N_327,N_493);
or U815 (N_815,N_393,N_417);
or U816 (N_816,N_294,N_481);
or U817 (N_817,N_131,N_297);
nand U818 (N_818,N_467,N_282);
and U819 (N_819,N_207,N_311);
or U820 (N_820,N_201,N_277);
and U821 (N_821,N_5,N_210);
or U822 (N_822,N_187,N_296);
or U823 (N_823,N_179,N_174);
or U824 (N_824,N_447,N_232);
nor U825 (N_825,N_315,N_290);
or U826 (N_826,N_157,N_410);
and U827 (N_827,N_243,N_484);
nand U828 (N_828,N_154,N_16);
or U829 (N_829,N_86,N_427);
nand U830 (N_830,N_335,N_132);
nor U831 (N_831,N_496,N_40);
or U832 (N_832,N_395,N_153);
nor U833 (N_833,N_213,N_398);
and U834 (N_834,N_233,N_34);
nor U835 (N_835,N_248,N_87);
nor U836 (N_836,N_241,N_145);
nand U837 (N_837,N_344,N_187);
and U838 (N_838,N_186,N_323);
and U839 (N_839,N_353,N_72);
or U840 (N_840,N_422,N_132);
or U841 (N_841,N_177,N_59);
nor U842 (N_842,N_184,N_228);
nand U843 (N_843,N_412,N_153);
xor U844 (N_844,N_216,N_148);
xor U845 (N_845,N_35,N_363);
or U846 (N_846,N_155,N_202);
or U847 (N_847,N_137,N_440);
nor U848 (N_848,N_472,N_149);
or U849 (N_849,N_81,N_270);
nor U850 (N_850,N_277,N_223);
and U851 (N_851,N_318,N_7);
or U852 (N_852,N_97,N_298);
nand U853 (N_853,N_47,N_196);
nand U854 (N_854,N_119,N_118);
nand U855 (N_855,N_275,N_155);
xnor U856 (N_856,N_342,N_212);
nor U857 (N_857,N_166,N_347);
and U858 (N_858,N_440,N_47);
nand U859 (N_859,N_50,N_297);
and U860 (N_860,N_186,N_483);
xnor U861 (N_861,N_113,N_328);
and U862 (N_862,N_47,N_178);
or U863 (N_863,N_164,N_466);
nor U864 (N_864,N_187,N_51);
or U865 (N_865,N_155,N_258);
nand U866 (N_866,N_485,N_321);
or U867 (N_867,N_333,N_32);
xnor U868 (N_868,N_384,N_273);
and U869 (N_869,N_189,N_329);
nor U870 (N_870,N_310,N_23);
nand U871 (N_871,N_195,N_168);
xnor U872 (N_872,N_359,N_370);
or U873 (N_873,N_52,N_277);
xor U874 (N_874,N_124,N_490);
nand U875 (N_875,N_134,N_416);
nor U876 (N_876,N_404,N_421);
nor U877 (N_877,N_141,N_184);
or U878 (N_878,N_335,N_251);
nor U879 (N_879,N_435,N_193);
nor U880 (N_880,N_383,N_257);
nor U881 (N_881,N_466,N_103);
xor U882 (N_882,N_127,N_366);
nand U883 (N_883,N_190,N_307);
nand U884 (N_884,N_159,N_281);
xor U885 (N_885,N_371,N_362);
or U886 (N_886,N_392,N_185);
nand U887 (N_887,N_47,N_161);
and U888 (N_888,N_441,N_329);
or U889 (N_889,N_201,N_281);
or U890 (N_890,N_101,N_34);
nand U891 (N_891,N_123,N_452);
and U892 (N_892,N_419,N_33);
nand U893 (N_893,N_15,N_306);
and U894 (N_894,N_213,N_82);
or U895 (N_895,N_493,N_413);
nand U896 (N_896,N_449,N_25);
nor U897 (N_897,N_29,N_108);
and U898 (N_898,N_11,N_57);
and U899 (N_899,N_132,N_274);
xnor U900 (N_900,N_67,N_367);
and U901 (N_901,N_128,N_37);
nand U902 (N_902,N_149,N_246);
and U903 (N_903,N_373,N_168);
xor U904 (N_904,N_264,N_468);
and U905 (N_905,N_117,N_455);
nor U906 (N_906,N_117,N_67);
or U907 (N_907,N_448,N_200);
or U908 (N_908,N_45,N_346);
or U909 (N_909,N_480,N_48);
xor U910 (N_910,N_36,N_105);
nand U911 (N_911,N_128,N_221);
and U912 (N_912,N_247,N_372);
and U913 (N_913,N_294,N_446);
nor U914 (N_914,N_461,N_305);
and U915 (N_915,N_93,N_448);
and U916 (N_916,N_158,N_317);
nand U917 (N_917,N_315,N_263);
xor U918 (N_918,N_459,N_478);
and U919 (N_919,N_175,N_257);
nor U920 (N_920,N_465,N_74);
and U921 (N_921,N_79,N_340);
or U922 (N_922,N_493,N_306);
or U923 (N_923,N_89,N_114);
and U924 (N_924,N_408,N_6);
and U925 (N_925,N_191,N_363);
nor U926 (N_926,N_307,N_220);
nor U927 (N_927,N_383,N_390);
nor U928 (N_928,N_347,N_120);
and U929 (N_929,N_362,N_124);
or U930 (N_930,N_54,N_380);
and U931 (N_931,N_446,N_64);
nand U932 (N_932,N_265,N_387);
and U933 (N_933,N_322,N_154);
nor U934 (N_934,N_370,N_65);
and U935 (N_935,N_253,N_269);
or U936 (N_936,N_425,N_481);
and U937 (N_937,N_68,N_332);
and U938 (N_938,N_357,N_88);
or U939 (N_939,N_94,N_374);
or U940 (N_940,N_264,N_60);
nand U941 (N_941,N_59,N_398);
or U942 (N_942,N_226,N_452);
or U943 (N_943,N_15,N_251);
or U944 (N_944,N_473,N_455);
or U945 (N_945,N_196,N_249);
nor U946 (N_946,N_98,N_278);
xnor U947 (N_947,N_432,N_422);
or U948 (N_948,N_383,N_234);
nand U949 (N_949,N_439,N_400);
xnor U950 (N_950,N_460,N_368);
nor U951 (N_951,N_26,N_481);
nand U952 (N_952,N_499,N_449);
or U953 (N_953,N_195,N_268);
and U954 (N_954,N_78,N_311);
xor U955 (N_955,N_408,N_175);
and U956 (N_956,N_5,N_128);
or U957 (N_957,N_494,N_452);
nand U958 (N_958,N_397,N_479);
nand U959 (N_959,N_176,N_411);
or U960 (N_960,N_146,N_299);
nand U961 (N_961,N_336,N_76);
or U962 (N_962,N_416,N_75);
or U963 (N_963,N_492,N_195);
and U964 (N_964,N_113,N_428);
nand U965 (N_965,N_114,N_440);
and U966 (N_966,N_412,N_342);
nor U967 (N_967,N_366,N_162);
and U968 (N_968,N_321,N_21);
nand U969 (N_969,N_370,N_410);
and U970 (N_970,N_9,N_466);
nand U971 (N_971,N_41,N_328);
and U972 (N_972,N_80,N_315);
and U973 (N_973,N_462,N_244);
xnor U974 (N_974,N_24,N_241);
and U975 (N_975,N_81,N_34);
or U976 (N_976,N_100,N_482);
and U977 (N_977,N_276,N_152);
or U978 (N_978,N_379,N_57);
or U979 (N_979,N_114,N_123);
nand U980 (N_980,N_434,N_225);
nand U981 (N_981,N_438,N_8);
or U982 (N_982,N_169,N_435);
nand U983 (N_983,N_9,N_146);
or U984 (N_984,N_246,N_159);
or U985 (N_985,N_477,N_473);
and U986 (N_986,N_455,N_191);
nor U987 (N_987,N_346,N_28);
or U988 (N_988,N_310,N_358);
nand U989 (N_989,N_230,N_336);
and U990 (N_990,N_76,N_166);
or U991 (N_991,N_53,N_307);
and U992 (N_992,N_483,N_326);
and U993 (N_993,N_74,N_193);
and U994 (N_994,N_354,N_436);
and U995 (N_995,N_191,N_402);
or U996 (N_996,N_305,N_489);
nor U997 (N_997,N_27,N_93);
xor U998 (N_998,N_173,N_160);
nand U999 (N_999,N_247,N_195);
and U1000 (N_1000,N_877,N_679);
nor U1001 (N_1001,N_927,N_507);
nand U1002 (N_1002,N_599,N_727);
and U1003 (N_1003,N_936,N_934);
nand U1004 (N_1004,N_772,N_520);
nand U1005 (N_1005,N_832,N_904);
and U1006 (N_1006,N_884,N_974);
xor U1007 (N_1007,N_728,N_981);
nor U1008 (N_1008,N_920,N_880);
or U1009 (N_1009,N_970,N_821);
nor U1010 (N_1010,N_574,N_778);
or U1011 (N_1011,N_533,N_606);
or U1012 (N_1012,N_871,N_590);
nor U1013 (N_1013,N_749,N_817);
nand U1014 (N_1014,N_966,N_989);
nand U1015 (N_1015,N_508,N_563);
nand U1016 (N_1016,N_947,N_743);
nor U1017 (N_1017,N_940,N_837);
or U1018 (N_1018,N_584,N_500);
or U1019 (N_1019,N_765,N_995);
nor U1020 (N_1020,N_654,N_651);
nand U1021 (N_1021,N_839,N_828);
or U1022 (N_1022,N_650,N_935);
nor U1023 (N_1023,N_648,N_805);
or U1024 (N_1024,N_907,N_949);
nand U1025 (N_1025,N_838,N_754);
and U1026 (N_1026,N_763,N_781);
nand U1027 (N_1027,N_597,N_776);
nor U1028 (N_1028,N_703,N_626);
and U1029 (N_1029,N_802,N_850);
nor U1030 (N_1030,N_867,N_916);
nor U1031 (N_1031,N_609,N_566);
nor U1032 (N_1032,N_761,N_784);
and U1033 (N_1033,N_572,N_782);
nand U1034 (N_1034,N_511,N_512);
nand U1035 (N_1035,N_742,N_843);
nand U1036 (N_1036,N_738,N_660);
or U1037 (N_1037,N_799,N_893);
xor U1038 (N_1038,N_918,N_993);
and U1039 (N_1039,N_774,N_810);
xor U1040 (N_1040,N_720,N_676);
or U1041 (N_1041,N_960,N_543);
or U1042 (N_1042,N_580,N_865);
and U1043 (N_1043,N_717,N_962);
nand U1044 (N_1044,N_823,N_898);
nand U1045 (N_1045,N_620,N_542);
nand U1046 (N_1046,N_640,N_712);
nor U1047 (N_1047,N_662,N_631);
nand U1048 (N_1048,N_564,N_524);
nor U1049 (N_1049,N_596,N_589);
nand U1050 (N_1050,N_702,N_967);
xor U1051 (N_1051,N_538,N_900);
and U1052 (N_1052,N_509,N_675);
xor U1053 (N_1053,N_922,N_856);
nor U1054 (N_1054,N_642,N_892);
nor U1055 (N_1055,N_943,N_889);
and U1056 (N_1056,N_753,N_536);
nor U1057 (N_1057,N_766,N_602);
or U1058 (N_1058,N_629,N_909);
nor U1059 (N_1059,N_628,N_658);
or U1060 (N_1060,N_671,N_687);
nand U1061 (N_1061,N_822,N_777);
and U1062 (N_1062,N_638,N_605);
and U1063 (N_1063,N_591,N_630);
or U1064 (N_1064,N_780,N_689);
and U1065 (N_1065,N_722,N_968);
nor U1066 (N_1066,N_706,N_724);
and U1067 (N_1067,N_827,N_721);
or U1068 (N_1068,N_692,N_562);
nor U1069 (N_1069,N_731,N_540);
and U1070 (N_1070,N_645,N_636);
or U1071 (N_1071,N_700,N_503);
nand U1072 (N_1072,N_846,N_882);
and U1073 (N_1073,N_764,N_812);
and U1074 (N_1074,N_614,N_710);
xor U1075 (N_1075,N_545,N_565);
and U1076 (N_1076,N_891,N_773);
or U1077 (N_1077,N_999,N_725);
nand U1078 (N_1078,N_752,N_746);
and U1079 (N_1079,N_635,N_548);
nand U1080 (N_1080,N_957,N_965);
xor U1081 (N_1081,N_866,N_627);
or U1082 (N_1082,N_872,N_969);
nor U1083 (N_1083,N_750,N_946);
and U1084 (N_1084,N_901,N_973);
nor U1085 (N_1085,N_905,N_992);
and U1086 (N_1086,N_868,N_666);
and U1087 (N_1087,N_632,N_885);
nand U1088 (N_1088,N_567,N_514);
and U1089 (N_1089,N_659,N_528);
and U1090 (N_1090,N_502,N_734);
nand U1091 (N_1091,N_762,N_751);
nor U1092 (N_1092,N_959,N_921);
and U1093 (N_1093,N_532,N_544);
nor U1094 (N_1094,N_852,N_816);
or U1095 (N_1095,N_860,N_622);
or U1096 (N_1096,N_719,N_624);
nand U1097 (N_1097,N_917,N_890);
nand U1098 (N_1098,N_757,N_771);
or U1099 (N_1099,N_558,N_896);
xor U1100 (N_1100,N_549,N_906);
nand U1101 (N_1101,N_996,N_691);
and U1102 (N_1102,N_678,N_581);
nor U1103 (N_1103,N_699,N_911);
and U1104 (N_1104,N_519,N_570);
nor U1105 (N_1105,N_547,N_997);
or U1106 (N_1106,N_736,N_592);
or U1107 (N_1107,N_539,N_815);
or U1108 (N_1108,N_732,N_663);
or U1109 (N_1109,N_579,N_932);
nor U1110 (N_1110,N_561,N_941);
nor U1111 (N_1111,N_861,N_914);
nor U1112 (N_1112,N_933,N_991);
and U1113 (N_1113,N_980,N_677);
nor U1114 (N_1114,N_615,N_505);
and U1115 (N_1115,N_972,N_859);
nor U1116 (N_1116,N_963,N_745);
and U1117 (N_1117,N_554,N_575);
xnor U1118 (N_1118,N_937,N_798);
or U1119 (N_1119,N_858,N_876);
nand U1120 (N_1120,N_600,N_644);
or U1121 (N_1121,N_652,N_744);
and U1122 (N_1122,N_740,N_693);
nand U1123 (N_1123,N_931,N_864);
and U1124 (N_1124,N_739,N_623);
and U1125 (N_1125,N_595,N_790);
and U1126 (N_1126,N_718,N_797);
and U1127 (N_1127,N_954,N_577);
and U1128 (N_1128,N_713,N_783);
and U1129 (N_1129,N_583,N_748);
and U1130 (N_1130,N_848,N_908);
nor U1131 (N_1131,N_930,N_964);
and U1132 (N_1132,N_515,N_836);
xnor U1133 (N_1133,N_696,N_851);
and U1134 (N_1134,N_842,N_807);
and U1135 (N_1135,N_813,N_681);
and U1136 (N_1136,N_715,N_986);
and U1137 (N_1137,N_804,N_688);
or U1138 (N_1138,N_534,N_811);
or U1139 (N_1139,N_793,N_814);
nand U1140 (N_1140,N_611,N_985);
nand U1141 (N_1141,N_801,N_573);
and U1142 (N_1142,N_690,N_958);
nor U1143 (N_1143,N_525,N_704);
nor U1144 (N_1144,N_618,N_879);
and U1145 (N_1145,N_672,N_741);
and U1146 (N_1146,N_521,N_910);
xnor U1147 (N_1147,N_998,N_786);
xnor U1148 (N_1148,N_919,N_598);
nand U1149 (N_1149,N_616,N_944);
nand U1150 (N_1150,N_705,N_818);
nor U1151 (N_1151,N_779,N_735);
or U1152 (N_1152,N_853,N_594);
or U1153 (N_1153,N_729,N_560);
nand U1154 (N_1154,N_601,N_657);
nand U1155 (N_1155,N_621,N_894);
and U1156 (N_1156,N_950,N_593);
xor U1157 (N_1157,N_878,N_669);
and U1158 (N_1158,N_559,N_956);
or U1159 (N_1159,N_707,N_613);
xor U1160 (N_1160,N_951,N_803);
or U1161 (N_1161,N_926,N_808);
nand U1162 (N_1162,N_637,N_646);
and U1163 (N_1163,N_768,N_649);
nand U1164 (N_1164,N_923,N_902);
or U1165 (N_1165,N_586,N_869);
and U1166 (N_1166,N_546,N_874);
nor U1167 (N_1167,N_979,N_854);
or U1168 (N_1168,N_971,N_684);
nor U1169 (N_1169,N_955,N_711);
nor U1170 (N_1170,N_826,N_915);
and U1171 (N_1171,N_552,N_680);
and U1172 (N_1172,N_903,N_953);
nor U1173 (N_1173,N_990,N_819);
and U1174 (N_1174,N_588,N_845);
or U1175 (N_1175,N_568,N_501);
or U1176 (N_1176,N_526,N_571);
xnor U1177 (N_1177,N_862,N_840);
nand U1178 (N_1178,N_978,N_531);
nand U1179 (N_1179,N_697,N_504);
nor U1180 (N_1180,N_683,N_523);
nor U1181 (N_1181,N_849,N_556);
nand U1182 (N_1182,N_714,N_643);
nor U1183 (N_1183,N_983,N_608);
or U1184 (N_1184,N_756,N_555);
nor U1185 (N_1185,N_834,N_899);
nand U1186 (N_1186,N_755,N_551);
nor U1187 (N_1187,N_825,N_716);
nand U1188 (N_1188,N_833,N_939);
and U1189 (N_1189,N_886,N_775);
and U1190 (N_1190,N_855,N_913);
nor U1191 (N_1191,N_708,N_875);
or U1192 (N_1192,N_661,N_800);
and U1193 (N_1193,N_888,N_522);
and U1194 (N_1194,N_550,N_948);
nor U1195 (N_1195,N_945,N_767);
or U1196 (N_1196,N_831,N_988);
nand U1197 (N_1197,N_794,N_977);
and U1198 (N_1198,N_639,N_517);
nand U1199 (N_1199,N_510,N_607);
nand U1200 (N_1200,N_667,N_938);
nor U1201 (N_1201,N_942,N_895);
and U1202 (N_1202,N_537,N_673);
or U1203 (N_1203,N_747,N_625);
or U1204 (N_1204,N_952,N_634);
and U1205 (N_1205,N_527,N_653);
nor U1206 (N_1206,N_610,N_604);
or U1207 (N_1207,N_694,N_857);
nand U1208 (N_1208,N_881,N_835);
and U1209 (N_1209,N_976,N_789);
or U1210 (N_1210,N_760,N_737);
and U1211 (N_1211,N_820,N_994);
and U1212 (N_1212,N_925,N_987);
nand U1213 (N_1213,N_770,N_529);
nand U1214 (N_1214,N_809,N_824);
nor U1215 (N_1215,N_733,N_576);
nor U1216 (N_1216,N_578,N_655);
and U1217 (N_1217,N_829,N_723);
nand U1218 (N_1218,N_730,N_769);
and U1219 (N_1219,N_695,N_633);
nand U1220 (N_1220,N_674,N_535);
nand U1221 (N_1221,N_665,N_518);
nand U1222 (N_1222,N_569,N_641);
xor U1223 (N_1223,N_830,N_787);
or U1224 (N_1224,N_796,N_582);
nand U1225 (N_1225,N_668,N_603);
xor U1226 (N_1226,N_788,N_897);
nor U1227 (N_1227,N_506,N_785);
nand U1228 (N_1228,N_585,N_928);
nand U1229 (N_1229,N_612,N_759);
nand U1230 (N_1230,N_686,N_726);
xnor U1231 (N_1231,N_806,N_887);
or U1232 (N_1232,N_587,N_791);
nor U1233 (N_1233,N_883,N_841);
xor U1234 (N_1234,N_541,N_984);
and U1235 (N_1235,N_758,N_844);
nand U1236 (N_1236,N_873,N_557);
nor U1237 (N_1237,N_617,N_513);
nand U1238 (N_1238,N_929,N_619);
nor U1239 (N_1239,N_792,N_847);
nand U1240 (N_1240,N_647,N_912);
xor U1241 (N_1241,N_982,N_795);
nand U1242 (N_1242,N_924,N_670);
and U1243 (N_1243,N_863,N_975);
xor U1244 (N_1244,N_870,N_701);
nor U1245 (N_1245,N_709,N_698);
nor U1246 (N_1246,N_553,N_656);
nand U1247 (N_1247,N_664,N_682);
or U1248 (N_1248,N_530,N_961);
and U1249 (N_1249,N_516,N_685);
nand U1250 (N_1250,N_645,N_930);
nand U1251 (N_1251,N_903,N_982);
nand U1252 (N_1252,N_891,N_606);
and U1253 (N_1253,N_610,N_807);
or U1254 (N_1254,N_825,N_687);
and U1255 (N_1255,N_971,N_654);
nand U1256 (N_1256,N_636,N_565);
and U1257 (N_1257,N_969,N_987);
nand U1258 (N_1258,N_540,N_723);
nand U1259 (N_1259,N_516,N_597);
nand U1260 (N_1260,N_575,N_685);
xor U1261 (N_1261,N_530,N_709);
xor U1262 (N_1262,N_933,N_595);
and U1263 (N_1263,N_754,N_749);
nand U1264 (N_1264,N_731,N_884);
and U1265 (N_1265,N_945,N_787);
xnor U1266 (N_1266,N_550,N_963);
and U1267 (N_1267,N_621,N_519);
nand U1268 (N_1268,N_552,N_933);
nor U1269 (N_1269,N_807,N_627);
nand U1270 (N_1270,N_813,N_610);
and U1271 (N_1271,N_775,N_808);
and U1272 (N_1272,N_731,N_801);
xnor U1273 (N_1273,N_550,N_568);
nand U1274 (N_1274,N_843,N_998);
nor U1275 (N_1275,N_593,N_926);
or U1276 (N_1276,N_739,N_610);
and U1277 (N_1277,N_851,N_975);
nor U1278 (N_1278,N_851,N_770);
nand U1279 (N_1279,N_828,N_883);
nand U1280 (N_1280,N_611,N_777);
xnor U1281 (N_1281,N_621,N_616);
or U1282 (N_1282,N_699,N_632);
nand U1283 (N_1283,N_661,N_509);
or U1284 (N_1284,N_726,N_594);
nand U1285 (N_1285,N_942,N_640);
or U1286 (N_1286,N_845,N_780);
nor U1287 (N_1287,N_529,N_938);
or U1288 (N_1288,N_658,N_579);
nand U1289 (N_1289,N_643,N_634);
nand U1290 (N_1290,N_929,N_930);
and U1291 (N_1291,N_780,N_677);
nand U1292 (N_1292,N_579,N_869);
and U1293 (N_1293,N_572,N_692);
or U1294 (N_1294,N_695,N_872);
nor U1295 (N_1295,N_686,N_846);
nand U1296 (N_1296,N_771,N_837);
nor U1297 (N_1297,N_999,N_534);
or U1298 (N_1298,N_761,N_956);
and U1299 (N_1299,N_719,N_503);
nand U1300 (N_1300,N_782,N_784);
or U1301 (N_1301,N_695,N_723);
nand U1302 (N_1302,N_927,N_833);
nand U1303 (N_1303,N_941,N_864);
or U1304 (N_1304,N_729,N_922);
nand U1305 (N_1305,N_838,N_940);
or U1306 (N_1306,N_621,N_506);
or U1307 (N_1307,N_858,N_905);
nor U1308 (N_1308,N_936,N_560);
or U1309 (N_1309,N_609,N_712);
nor U1310 (N_1310,N_918,N_666);
nand U1311 (N_1311,N_764,N_855);
nand U1312 (N_1312,N_910,N_951);
and U1313 (N_1313,N_545,N_933);
or U1314 (N_1314,N_751,N_641);
nor U1315 (N_1315,N_564,N_502);
and U1316 (N_1316,N_957,N_884);
or U1317 (N_1317,N_900,N_703);
nor U1318 (N_1318,N_517,N_539);
nand U1319 (N_1319,N_991,N_727);
and U1320 (N_1320,N_989,N_619);
and U1321 (N_1321,N_747,N_965);
xor U1322 (N_1322,N_897,N_595);
and U1323 (N_1323,N_921,N_955);
or U1324 (N_1324,N_686,N_963);
nor U1325 (N_1325,N_634,N_549);
or U1326 (N_1326,N_844,N_900);
and U1327 (N_1327,N_720,N_812);
and U1328 (N_1328,N_621,N_861);
or U1329 (N_1329,N_609,N_528);
nor U1330 (N_1330,N_907,N_993);
nand U1331 (N_1331,N_932,N_948);
and U1332 (N_1332,N_817,N_768);
nand U1333 (N_1333,N_996,N_582);
or U1334 (N_1334,N_602,N_876);
and U1335 (N_1335,N_987,N_606);
and U1336 (N_1336,N_785,N_875);
or U1337 (N_1337,N_559,N_766);
nor U1338 (N_1338,N_933,N_588);
nor U1339 (N_1339,N_617,N_960);
nor U1340 (N_1340,N_972,N_935);
or U1341 (N_1341,N_614,N_868);
and U1342 (N_1342,N_690,N_618);
or U1343 (N_1343,N_666,N_665);
nand U1344 (N_1344,N_804,N_865);
nor U1345 (N_1345,N_558,N_646);
nand U1346 (N_1346,N_953,N_651);
nand U1347 (N_1347,N_847,N_882);
nand U1348 (N_1348,N_947,N_642);
or U1349 (N_1349,N_913,N_628);
or U1350 (N_1350,N_679,N_631);
nor U1351 (N_1351,N_894,N_619);
nand U1352 (N_1352,N_706,N_730);
or U1353 (N_1353,N_531,N_900);
nor U1354 (N_1354,N_864,N_719);
and U1355 (N_1355,N_627,N_500);
or U1356 (N_1356,N_794,N_938);
or U1357 (N_1357,N_811,N_710);
or U1358 (N_1358,N_750,N_569);
xor U1359 (N_1359,N_683,N_657);
nand U1360 (N_1360,N_791,N_665);
and U1361 (N_1361,N_633,N_959);
nor U1362 (N_1362,N_798,N_563);
nor U1363 (N_1363,N_526,N_653);
and U1364 (N_1364,N_954,N_710);
nor U1365 (N_1365,N_993,N_825);
nand U1366 (N_1366,N_998,N_763);
nand U1367 (N_1367,N_575,N_611);
nand U1368 (N_1368,N_575,N_602);
or U1369 (N_1369,N_637,N_666);
or U1370 (N_1370,N_780,N_886);
nor U1371 (N_1371,N_591,N_578);
nor U1372 (N_1372,N_554,N_959);
and U1373 (N_1373,N_670,N_559);
or U1374 (N_1374,N_653,N_545);
nor U1375 (N_1375,N_689,N_610);
xnor U1376 (N_1376,N_884,N_682);
nand U1377 (N_1377,N_711,N_774);
or U1378 (N_1378,N_886,N_623);
nor U1379 (N_1379,N_621,N_577);
nand U1380 (N_1380,N_864,N_717);
or U1381 (N_1381,N_582,N_816);
nor U1382 (N_1382,N_519,N_810);
xnor U1383 (N_1383,N_949,N_791);
nor U1384 (N_1384,N_929,N_516);
nand U1385 (N_1385,N_601,N_861);
nor U1386 (N_1386,N_547,N_830);
nor U1387 (N_1387,N_824,N_784);
nand U1388 (N_1388,N_748,N_700);
nor U1389 (N_1389,N_580,N_601);
or U1390 (N_1390,N_636,N_691);
nand U1391 (N_1391,N_758,N_649);
or U1392 (N_1392,N_627,N_677);
and U1393 (N_1393,N_616,N_608);
nand U1394 (N_1394,N_513,N_764);
or U1395 (N_1395,N_646,N_843);
nor U1396 (N_1396,N_791,N_749);
nor U1397 (N_1397,N_693,N_679);
or U1398 (N_1398,N_864,N_824);
nor U1399 (N_1399,N_919,N_909);
and U1400 (N_1400,N_564,N_606);
or U1401 (N_1401,N_768,N_564);
xnor U1402 (N_1402,N_928,N_533);
or U1403 (N_1403,N_724,N_776);
nor U1404 (N_1404,N_778,N_641);
or U1405 (N_1405,N_567,N_854);
or U1406 (N_1406,N_840,N_835);
nand U1407 (N_1407,N_642,N_666);
nor U1408 (N_1408,N_515,N_707);
nor U1409 (N_1409,N_639,N_610);
nor U1410 (N_1410,N_586,N_713);
nand U1411 (N_1411,N_554,N_791);
and U1412 (N_1412,N_675,N_680);
nor U1413 (N_1413,N_788,N_826);
or U1414 (N_1414,N_788,N_813);
nand U1415 (N_1415,N_841,N_801);
and U1416 (N_1416,N_987,N_746);
nand U1417 (N_1417,N_686,N_955);
nor U1418 (N_1418,N_705,N_512);
or U1419 (N_1419,N_708,N_929);
xor U1420 (N_1420,N_963,N_988);
nor U1421 (N_1421,N_786,N_513);
nor U1422 (N_1422,N_797,N_921);
xnor U1423 (N_1423,N_611,N_683);
xor U1424 (N_1424,N_635,N_514);
xor U1425 (N_1425,N_977,N_943);
nor U1426 (N_1426,N_666,N_872);
nor U1427 (N_1427,N_658,N_983);
and U1428 (N_1428,N_638,N_624);
nand U1429 (N_1429,N_891,N_677);
nor U1430 (N_1430,N_744,N_562);
and U1431 (N_1431,N_616,N_689);
or U1432 (N_1432,N_870,N_647);
and U1433 (N_1433,N_699,N_639);
or U1434 (N_1434,N_932,N_711);
nand U1435 (N_1435,N_502,N_730);
and U1436 (N_1436,N_576,N_505);
nor U1437 (N_1437,N_937,N_569);
nand U1438 (N_1438,N_838,N_761);
and U1439 (N_1439,N_827,N_708);
nand U1440 (N_1440,N_676,N_939);
nand U1441 (N_1441,N_905,N_739);
xor U1442 (N_1442,N_594,N_788);
xnor U1443 (N_1443,N_915,N_657);
nor U1444 (N_1444,N_715,N_724);
and U1445 (N_1445,N_925,N_555);
and U1446 (N_1446,N_609,N_726);
nand U1447 (N_1447,N_589,N_996);
nand U1448 (N_1448,N_725,N_524);
and U1449 (N_1449,N_506,N_728);
nand U1450 (N_1450,N_567,N_776);
nor U1451 (N_1451,N_766,N_953);
nand U1452 (N_1452,N_683,N_688);
and U1453 (N_1453,N_948,N_639);
xnor U1454 (N_1454,N_962,N_983);
and U1455 (N_1455,N_863,N_890);
or U1456 (N_1456,N_771,N_549);
xnor U1457 (N_1457,N_729,N_972);
xnor U1458 (N_1458,N_755,N_629);
nand U1459 (N_1459,N_850,N_654);
or U1460 (N_1460,N_740,N_618);
nor U1461 (N_1461,N_892,N_566);
or U1462 (N_1462,N_849,N_723);
or U1463 (N_1463,N_860,N_789);
xor U1464 (N_1464,N_713,N_757);
nand U1465 (N_1465,N_953,N_865);
nand U1466 (N_1466,N_854,N_841);
or U1467 (N_1467,N_981,N_580);
and U1468 (N_1468,N_830,N_822);
nand U1469 (N_1469,N_985,N_856);
nand U1470 (N_1470,N_842,N_829);
xnor U1471 (N_1471,N_602,N_790);
and U1472 (N_1472,N_528,N_893);
and U1473 (N_1473,N_933,N_994);
nor U1474 (N_1474,N_791,N_612);
nor U1475 (N_1475,N_604,N_817);
xnor U1476 (N_1476,N_849,N_620);
and U1477 (N_1477,N_607,N_637);
and U1478 (N_1478,N_870,N_822);
nor U1479 (N_1479,N_568,N_796);
nor U1480 (N_1480,N_784,N_516);
nor U1481 (N_1481,N_755,N_520);
or U1482 (N_1482,N_924,N_890);
nand U1483 (N_1483,N_846,N_849);
or U1484 (N_1484,N_543,N_752);
nor U1485 (N_1485,N_544,N_994);
xor U1486 (N_1486,N_842,N_515);
nand U1487 (N_1487,N_504,N_644);
and U1488 (N_1488,N_662,N_879);
nor U1489 (N_1489,N_670,N_593);
nand U1490 (N_1490,N_564,N_504);
nor U1491 (N_1491,N_742,N_649);
nor U1492 (N_1492,N_976,N_518);
or U1493 (N_1493,N_553,N_506);
nor U1494 (N_1494,N_575,N_771);
nor U1495 (N_1495,N_761,N_803);
nand U1496 (N_1496,N_646,N_984);
nor U1497 (N_1497,N_905,N_598);
nand U1498 (N_1498,N_865,N_792);
nor U1499 (N_1499,N_740,N_593);
nand U1500 (N_1500,N_1404,N_1017);
and U1501 (N_1501,N_1417,N_1368);
nor U1502 (N_1502,N_1282,N_1449);
and U1503 (N_1503,N_1107,N_1366);
nor U1504 (N_1504,N_1038,N_1408);
and U1505 (N_1505,N_1188,N_1491);
nand U1506 (N_1506,N_1314,N_1388);
nand U1507 (N_1507,N_1042,N_1421);
and U1508 (N_1508,N_1485,N_1353);
and U1509 (N_1509,N_1114,N_1145);
xnor U1510 (N_1510,N_1395,N_1091);
nor U1511 (N_1511,N_1046,N_1078);
and U1512 (N_1512,N_1482,N_1202);
and U1513 (N_1513,N_1250,N_1195);
nand U1514 (N_1514,N_1229,N_1105);
xnor U1515 (N_1515,N_1182,N_1120);
xnor U1516 (N_1516,N_1310,N_1129);
or U1517 (N_1517,N_1080,N_1071);
nand U1518 (N_1518,N_1049,N_1255);
nor U1519 (N_1519,N_1471,N_1010);
nand U1520 (N_1520,N_1242,N_1397);
or U1521 (N_1521,N_1062,N_1407);
and U1522 (N_1522,N_1389,N_1492);
nor U1523 (N_1523,N_1064,N_1293);
xor U1524 (N_1524,N_1086,N_1462);
xnor U1525 (N_1525,N_1138,N_1193);
and U1526 (N_1526,N_1127,N_1169);
or U1527 (N_1527,N_1094,N_1158);
nand U1528 (N_1528,N_1377,N_1439);
nor U1529 (N_1529,N_1416,N_1263);
nor U1530 (N_1530,N_1192,N_1300);
nand U1531 (N_1531,N_1348,N_1331);
nand U1532 (N_1532,N_1019,N_1164);
or U1533 (N_1533,N_1066,N_1065);
xnor U1534 (N_1534,N_1330,N_1000);
and U1535 (N_1535,N_1179,N_1464);
or U1536 (N_1536,N_1296,N_1484);
nand U1537 (N_1537,N_1026,N_1034);
or U1538 (N_1538,N_1171,N_1432);
or U1539 (N_1539,N_1170,N_1266);
xnor U1540 (N_1540,N_1394,N_1362);
and U1541 (N_1541,N_1496,N_1039);
or U1542 (N_1542,N_1008,N_1381);
or U1543 (N_1543,N_1470,N_1097);
or U1544 (N_1544,N_1092,N_1116);
or U1545 (N_1545,N_1458,N_1288);
and U1546 (N_1546,N_1048,N_1396);
nand U1547 (N_1547,N_1441,N_1117);
nor U1548 (N_1548,N_1316,N_1084);
and U1549 (N_1549,N_1390,N_1385);
nor U1550 (N_1550,N_1118,N_1443);
xor U1551 (N_1551,N_1328,N_1299);
nor U1552 (N_1552,N_1350,N_1361);
nand U1553 (N_1553,N_1246,N_1448);
nor U1554 (N_1554,N_1486,N_1455);
or U1555 (N_1555,N_1355,N_1196);
and U1556 (N_1556,N_1096,N_1338);
nand U1557 (N_1557,N_1302,N_1332);
and U1558 (N_1558,N_1254,N_1445);
and U1559 (N_1559,N_1208,N_1378);
xnor U1560 (N_1560,N_1317,N_1498);
nor U1561 (N_1561,N_1480,N_1004);
nand U1562 (N_1562,N_1075,N_1274);
nand U1563 (N_1563,N_1037,N_1359);
and U1564 (N_1564,N_1043,N_1015);
nand U1565 (N_1565,N_1121,N_1234);
and U1566 (N_1566,N_1029,N_1238);
xor U1567 (N_1567,N_1052,N_1200);
nor U1568 (N_1568,N_1349,N_1167);
and U1569 (N_1569,N_1313,N_1028);
nand U1570 (N_1570,N_1468,N_1183);
and U1571 (N_1571,N_1420,N_1499);
nand U1572 (N_1572,N_1303,N_1356);
nand U1573 (N_1573,N_1024,N_1122);
and U1574 (N_1574,N_1239,N_1237);
xnor U1575 (N_1575,N_1184,N_1190);
or U1576 (N_1576,N_1232,N_1228);
nand U1577 (N_1577,N_1260,N_1321);
nor U1578 (N_1578,N_1156,N_1241);
nand U1579 (N_1579,N_1067,N_1281);
nand U1580 (N_1580,N_1447,N_1344);
and U1581 (N_1581,N_1068,N_1273);
nor U1582 (N_1582,N_1459,N_1128);
or U1583 (N_1583,N_1176,N_1002);
nand U1584 (N_1584,N_1110,N_1093);
or U1585 (N_1585,N_1370,N_1055);
nor U1586 (N_1586,N_1283,N_1469);
nor U1587 (N_1587,N_1044,N_1473);
and U1588 (N_1588,N_1279,N_1376);
nor U1589 (N_1589,N_1380,N_1419);
nand U1590 (N_1590,N_1379,N_1392);
or U1591 (N_1591,N_1347,N_1318);
or U1592 (N_1592,N_1460,N_1206);
and U1593 (N_1593,N_1157,N_1222);
or U1594 (N_1594,N_1166,N_1187);
nand U1595 (N_1595,N_1141,N_1324);
xnor U1596 (N_1596,N_1357,N_1178);
nand U1597 (N_1597,N_1087,N_1375);
nor U1598 (N_1598,N_1415,N_1005);
or U1599 (N_1599,N_1257,N_1382);
and U1600 (N_1600,N_1494,N_1259);
nand U1601 (N_1601,N_1467,N_1453);
and U1602 (N_1602,N_1147,N_1016);
nor U1603 (N_1603,N_1069,N_1213);
nor U1604 (N_1604,N_1082,N_1045);
and U1605 (N_1605,N_1223,N_1033);
and U1606 (N_1606,N_1051,N_1360);
or U1607 (N_1607,N_1411,N_1267);
or U1608 (N_1608,N_1103,N_1403);
or U1609 (N_1609,N_1053,N_1315);
or U1610 (N_1610,N_1244,N_1233);
nand U1611 (N_1611,N_1327,N_1493);
or U1612 (N_1612,N_1099,N_1150);
or U1613 (N_1613,N_1275,N_1134);
nand U1614 (N_1614,N_1210,N_1346);
and U1615 (N_1615,N_1027,N_1189);
nand U1616 (N_1616,N_1077,N_1427);
and U1617 (N_1617,N_1256,N_1426);
nand U1618 (N_1618,N_1262,N_1140);
nand U1619 (N_1619,N_1339,N_1104);
or U1620 (N_1620,N_1204,N_1144);
nor U1621 (N_1621,N_1336,N_1290);
or U1622 (N_1622,N_1240,N_1216);
xnor U1623 (N_1623,N_1139,N_1136);
or U1624 (N_1624,N_1444,N_1124);
xnor U1625 (N_1625,N_1334,N_1243);
and U1626 (N_1626,N_1225,N_1456);
nand U1627 (N_1627,N_1264,N_1333);
nor U1628 (N_1628,N_1374,N_1436);
or U1629 (N_1629,N_1474,N_1036);
or U1630 (N_1630,N_1387,N_1070);
and U1631 (N_1631,N_1047,N_1035);
and U1632 (N_1632,N_1154,N_1265);
nand U1633 (N_1633,N_1020,N_1161);
nand U1634 (N_1634,N_1384,N_1115);
xor U1635 (N_1635,N_1340,N_1323);
nand U1636 (N_1636,N_1088,N_1442);
nand U1637 (N_1637,N_1057,N_1422);
or U1638 (N_1638,N_1247,N_1292);
or U1639 (N_1639,N_1297,N_1220);
or U1640 (N_1640,N_1197,N_1011);
or U1641 (N_1641,N_1177,N_1412);
and U1642 (N_1642,N_1450,N_1325);
xor U1643 (N_1643,N_1351,N_1320);
and U1644 (N_1644,N_1425,N_1059);
nand U1645 (N_1645,N_1009,N_1423);
nand U1646 (N_1646,N_1430,N_1497);
nor U1647 (N_1647,N_1090,N_1476);
and U1648 (N_1648,N_1413,N_1245);
xnor U1649 (N_1649,N_1372,N_1060);
nor U1650 (N_1650,N_1341,N_1101);
nand U1651 (N_1651,N_1304,N_1072);
xnor U1652 (N_1652,N_1465,N_1386);
and U1653 (N_1653,N_1106,N_1214);
xor U1654 (N_1654,N_1174,N_1143);
or U1655 (N_1655,N_1477,N_1130);
nand U1656 (N_1656,N_1226,N_1481);
xnor U1657 (N_1657,N_1451,N_1074);
or U1658 (N_1658,N_1058,N_1218);
and U1659 (N_1659,N_1311,N_1146);
nor U1660 (N_1660,N_1235,N_1018);
nand U1661 (N_1661,N_1402,N_1014);
xnor U1662 (N_1662,N_1123,N_1006);
nor U1663 (N_1663,N_1001,N_1335);
or U1664 (N_1664,N_1148,N_1230);
or U1665 (N_1665,N_1312,N_1209);
nor U1666 (N_1666,N_1367,N_1406);
or U1667 (N_1667,N_1050,N_1268);
and U1668 (N_1668,N_1440,N_1405);
xnor U1669 (N_1669,N_1424,N_1270);
nand U1670 (N_1670,N_1112,N_1085);
and U1671 (N_1671,N_1261,N_1199);
xnor U1672 (N_1672,N_1137,N_1463);
nand U1673 (N_1673,N_1201,N_1021);
nand U1674 (N_1674,N_1227,N_1398);
or U1675 (N_1675,N_1152,N_1061);
or U1676 (N_1676,N_1369,N_1194);
nor U1677 (N_1677,N_1181,N_1249);
and U1678 (N_1678,N_1013,N_1354);
nand U1679 (N_1679,N_1475,N_1373);
nand U1680 (N_1680,N_1025,N_1163);
nand U1681 (N_1681,N_1291,N_1253);
or U1682 (N_1682,N_1248,N_1159);
xnor U1683 (N_1683,N_1278,N_1012);
xor U1684 (N_1684,N_1102,N_1433);
or U1685 (N_1685,N_1098,N_1337);
nor U1686 (N_1686,N_1400,N_1032);
nor U1687 (N_1687,N_1149,N_1211);
nor U1688 (N_1688,N_1217,N_1329);
nor U1689 (N_1689,N_1003,N_1095);
xnor U1690 (N_1690,N_1393,N_1488);
or U1691 (N_1691,N_1364,N_1111);
or U1692 (N_1692,N_1457,N_1073);
or U1693 (N_1693,N_1186,N_1126);
and U1694 (N_1694,N_1132,N_1414);
xor U1695 (N_1695,N_1461,N_1089);
nor U1696 (N_1696,N_1221,N_1401);
and U1697 (N_1697,N_1125,N_1345);
and U1698 (N_1698,N_1307,N_1434);
and U1699 (N_1699,N_1435,N_1454);
nand U1700 (N_1700,N_1295,N_1446);
and U1701 (N_1701,N_1437,N_1487);
nor U1702 (N_1702,N_1391,N_1277);
xor U1703 (N_1703,N_1284,N_1083);
nand U1704 (N_1704,N_1185,N_1478);
nand U1705 (N_1705,N_1041,N_1180);
or U1706 (N_1706,N_1276,N_1215);
nor U1707 (N_1707,N_1322,N_1151);
nor U1708 (N_1708,N_1198,N_1483);
and U1709 (N_1709,N_1258,N_1286);
nor U1710 (N_1710,N_1289,N_1172);
nand U1711 (N_1711,N_1131,N_1119);
nand U1712 (N_1712,N_1162,N_1142);
nand U1713 (N_1713,N_1438,N_1301);
nand U1714 (N_1714,N_1294,N_1219);
or U1715 (N_1715,N_1030,N_1113);
or U1716 (N_1716,N_1452,N_1371);
and U1717 (N_1717,N_1495,N_1022);
nand U1718 (N_1718,N_1272,N_1409);
and U1719 (N_1719,N_1358,N_1054);
nor U1720 (N_1720,N_1431,N_1287);
and U1721 (N_1721,N_1363,N_1175);
nand U1722 (N_1722,N_1207,N_1383);
xnor U1723 (N_1723,N_1203,N_1133);
xor U1724 (N_1724,N_1271,N_1490);
nor U1725 (N_1725,N_1489,N_1165);
nor U1726 (N_1726,N_1399,N_1472);
nor U1727 (N_1727,N_1056,N_1040);
nor U1728 (N_1728,N_1479,N_1173);
xnor U1729 (N_1729,N_1343,N_1280);
or U1730 (N_1730,N_1410,N_1305);
nor U1731 (N_1731,N_1079,N_1269);
and U1732 (N_1732,N_1160,N_1063);
or U1733 (N_1733,N_1251,N_1236);
nor U1734 (N_1734,N_1428,N_1135);
or U1735 (N_1735,N_1252,N_1309);
and U1736 (N_1736,N_1298,N_1224);
nand U1737 (N_1737,N_1076,N_1231);
and U1738 (N_1738,N_1205,N_1308);
nand U1739 (N_1739,N_1212,N_1108);
or U1740 (N_1740,N_1326,N_1081);
nand U1741 (N_1741,N_1153,N_1352);
and U1742 (N_1742,N_1155,N_1342);
nand U1743 (N_1743,N_1100,N_1285);
and U1744 (N_1744,N_1466,N_1007);
or U1745 (N_1745,N_1306,N_1365);
xnor U1746 (N_1746,N_1319,N_1191);
or U1747 (N_1747,N_1168,N_1418);
and U1748 (N_1748,N_1109,N_1429);
xor U1749 (N_1749,N_1031,N_1023);
xor U1750 (N_1750,N_1322,N_1055);
nand U1751 (N_1751,N_1162,N_1417);
nor U1752 (N_1752,N_1034,N_1161);
nand U1753 (N_1753,N_1362,N_1285);
or U1754 (N_1754,N_1467,N_1142);
and U1755 (N_1755,N_1097,N_1384);
xnor U1756 (N_1756,N_1280,N_1089);
or U1757 (N_1757,N_1101,N_1289);
nor U1758 (N_1758,N_1311,N_1144);
or U1759 (N_1759,N_1107,N_1471);
or U1760 (N_1760,N_1110,N_1042);
nand U1761 (N_1761,N_1348,N_1086);
or U1762 (N_1762,N_1299,N_1260);
nor U1763 (N_1763,N_1015,N_1494);
or U1764 (N_1764,N_1489,N_1189);
nor U1765 (N_1765,N_1053,N_1389);
or U1766 (N_1766,N_1320,N_1137);
or U1767 (N_1767,N_1083,N_1262);
or U1768 (N_1768,N_1471,N_1198);
nand U1769 (N_1769,N_1325,N_1338);
and U1770 (N_1770,N_1069,N_1241);
and U1771 (N_1771,N_1082,N_1312);
nor U1772 (N_1772,N_1096,N_1016);
and U1773 (N_1773,N_1309,N_1105);
nand U1774 (N_1774,N_1113,N_1480);
or U1775 (N_1775,N_1009,N_1344);
nand U1776 (N_1776,N_1018,N_1254);
xnor U1777 (N_1777,N_1453,N_1318);
or U1778 (N_1778,N_1049,N_1330);
nor U1779 (N_1779,N_1439,N_1387);
nor U1780 (N_1780,N_1029,N_1188);
xnor U1781 (N_1781,N_1056,N_1226);
and U1782 (N_1782,N_1265,N_1033);
nor U1783 (N_1783,N_1260,N_1002);
nor U1784 (N_1784,N_1474,N_1407);
and U1785 (N_1785,N_1424,N_1227);
and U1786 (N_1786,N_1385,N_1141);
or U1787 (N_1787,N_1034,N_1486);
and U1788 (N_1788,N_1278,N_1109);
nor U1789 (N_1789,N_1198,N_1005);
or U1790 (N_1790,N_1339,N_1473);
or U1791 (N_1791,N_1177,N_1319);
and U1792 (N_1792,N_1144,N_1073);
nor U1793 (N_1793,N_1278,N_1329);
or U1794 (N_1794,N_1219,N_1103);
nand U1795 (N_1795,N_1209,N_1414);
or U1796 (N_1796,N_1434,N_1405);
or U1797 (N_1797,N_1042,N_1408);
nand U1798 (N_1798,N_1309,N_1321);
and U1799 (N_1799,N_1453,N_1332);
nand U1800 (N_1800,N_1203,N_1329);
and U1801 (N_1801,N_1175,N_1426);
or U1802 (N_1802,N_1276,N_1233);
and U1803 (N_1803,N_1019,N_1313);
xor U1804 (N_1804,N_1131,N_1296);
nor U1805 (N_1805,N_1056,N_1152);
nand U1806 (N_1806,N_1106,N_1255);
nand U1807 (N_1807,N_1135,N_1083);
xnor U1808 (N_1808,N_1116,N_1122);
nor U1809 (N_1809,N_1308,N_1285);
nor U1810 (N_1810,N_1154,N_1001);
nor U1811 (N_1811,N_1047,N_1416);
and U1812 (N_1812,N_1063,N_1022);
xor U1813 (N_1813,N_1326,N_1177);
or U1814 (N_1814,N_1051,N_1171);
and U1815 (N_1815,N_1363,N_1118);
and U1816 (N_1816,N_1326,N_1377);
or U1817 (N_1817,N_1210,N_1291);
and U1818 (N_1818,N_1440,N_1028);
or U1819 (N_1819,N_1103,N_1430);
nor U1820 (N_1820,N_1119,N_1413);
and U1821 (N_1821,N_1444,N_1337);
nor U1822 (N_1822,N_1395,N_1171);
nor U1823 (N_1823,N_1442,N_1140);
nor U1824 (N_1824,N_1483,N_1068);
xnor U1825 (N_1825,N_1348,N_1007);
or U1826 (N_1826,N_1250,N_1415);
nand U1827 (N_1827,N_1209,N_1416);
xor U1828 (N_1828,N_1305,N_1252);
and U1829 (N_1829,N_1044,N_1209);
or U1830 (N_1830,N_1028,N_1356);
and U1831 (N_1831,N_1343,N_1071);
and U1832 (N_1832,N_1371,N_1312);
nand U1833 (N_1833,N_1189,N_1429);
nor U1834 (N_1834,N_1243,N_1031);
or U1835 (N_1835,N_1031,N_1294);
or U1836 (N_1836,N_1341,N_1195);
nand U1837 (N_1837,N_1274,N_1011);
and U1838 (N_1838,N_1278,N_1083);
nand U1839 (N_1839,N_1026,N_1055);
nand U1840 (N_1840,N_1046,N_1122);
nor U1841 (N_1841,N_1029,N_1288);
and U1842 (N_1842,N_1128,N_1360);
nand U1843 (N_1843,N_1333,N_1404);
and U1844 (N_1844,N_1160,N_1198);
xnor U1845 (N_1845,N_1202,N_1322);
and U1846 (N_1846,N_1051,N_1207);
and U1847 (N_1847,N_1483,N_1046);
and U1848 (N_1848,N_1381,N_1370);
nor U1849 (N_1849,N_1175,N_1275);
nor U1850 (N_1850,N_1460,N_1345);
nor U1851 (N_1851,N_1496,N_1319);
xnor U1852 (N_1852,N_1399,N_1103);
nor U1853 (N_1853,N_1234,N_1466);
xnor U1854 (N_1854,N_1340,N_1334);
or U1855 (N_1855,N_1187,N_1005);
and U1856 (N_1856,N_1316,N_1083);
and U1857 (N_1857,N_1310,N_1146);
and U1858 (N_1858,N_1377,N_1425);
or U1859 (N_1859,N_1388,N_1453);
xnor U1860 (N_1860,N_1215,N_1413);
nor U1861 (N_1861,N_1255,N_1493);
and U1862 (N_1862,N_1371,N_1290);
nand U1863 (N_1863,N_1242,N_1358);
or U1864 (N_1864,N_1133,N_1427);
nor U1865 (N_1865,N_1176,N_1450);
or U1866 (N_1866,N_1392,N_1414);
and U1867 (N_1867,N_1165,N_1111);
and U1868 (N_1868,N_1476,N_1093);
nor U1869 (N_1869,N_1209,N_1212);
and U1870 (N_1870,N_1314,N_1309);
and U1871 (N_1871,N_1107,N_1179);
nand U1872 (N_1872,N_1388,N_1139);
or U1873 (N_1873,N_1195,N_1268);
and U1874 (N_1874,N_1442,N_1487);
nand U1875 (N_1875,N_1129,N_1388);
and U1876 (N_1876,N_1026,N_1235);
and U1877 (N_1877,N_1382,N_1351);
nor U1878 (N_1878,N_1052,N_1076);
and U1879 (N_1879,N_1406,N_1322);
nor U1880 (N_1880,N_1225,N_1126);
nand U1881 (N_1881,N_1425,N_1283);
or U1882 (N_1882,N_1250,N_1316);
or U1883 (N_1883,N_1409,N_1379);
and U1884 (N_1884,N_1192,N_1433);
and U1885 (N_1885,N_1149,N_1476);
or U1886 (N_1886,N_1381,N_1417);
xor U1887 (N_1887,N_1003,N_1404);
and U1888 (N_1888,N_1173,N_1319);
nor U1889 (N_1889,N_1363,N_1135);
nand U1890 (N_1890,N_1319,N_1379);
or U1891 (N_1891,N_1303,N_1113);
or U1892 (N_1892,N_1174,N_1087);
nand U1893 (N_1893,N_1445,N_1159);
and U1894 (N_1894,N_1175,N_1095);
and U1895 (N_1895,N_1488,N_1249);
nor U1896 (N_1896,N_1055,N_1223);
xor U1897 (N_1897,N_1262,N_1183);
or U1898 (N_1898,N_1028,N_1099);
or U1899 (N_1899,N_1308,N_1317);
xor U1900 (N_1900,N_1030,N_1495);
and U1901 (N_1901,N_1256,N_1393);
or U1902 (N_1902,N_1482,N_1445);
and U1903 (N_1903,N_1163,N_1201);
and U1904 (N_1904,N_1020,N_1134);
nor U1905 (N_1905,N_1120,N_1079);
nor U1906 (N_1906,N_1189,N_1252);
or U1907 (N_1907,N_1330,N_1044);
and U1908 (N_1908,N_1269,N_1292);
xor U1909 (N_1909,N_1249,N_1025);
and U1910 (N_1910,N_1316,N_1498);
and U1911 (N_1911,N_1187,N_1240);
nor U1912 (N_1912,N_1057,N_1232);
nand U1913 (N_1913,N_1167,N_1102);
xor U1914 (N_1914,N_1220,N_1027);
and U1915 (N_1915,N_1469,N_1480);
or U1916 (N_1916,N_1015,N_1206);
and U1917 (N_1917,N_1329,N_1361);
and U1918 (N_1918,N_1365,N_1256);
xor U1919 (N_1919,N_1204,N_1232);
or U1920 (N_1920,N_1343,N_1329);
nor U1921 (N_1921,N_1100,N_1430);
or U1922 (N_1922,N_1349,N_1240);
nor U1923 (N_1923,N_1041,N_1066);
and U1924 (N_1924,N_1395,N_1033);
nand U1925 (N_1925,N_1221,N_1304);
and U1926 (N_1926,N_1008,N_1014);
nand U1927 (N_1927,N_1353,N_1468);
nor U1928 (N_1928,N_1038,N_1037);
nand U1929 (N_1929,N_1161,N_1446);
nand U1930 (N_1930,N_1214,N_1114);
nand U1931 (N_1931,N_1093,N_1375);
nand U1932 (N_1932,N_1461,N_1292);
or U1933 (N_1933,N_1377,N_1271);
or U1934 (N_1934,N_1304,N_1440);
nand U1935 (N_1935,N_1313,N_1201);
nand U1936 (N_1936,N_1241,N_1493);
nor U1937 (N_1937,N_1142,N_1381);
or U1938 (N_1938,N_1171,N_1496);
nand U1939 (N_1939,N_1293,N_1005);
or U1940 (N_1940,N_1227,N_1328);
xnor U1941 (N_1941,N_1107,N_1375);
nand U1942 (N_1942,N_1383,N_1444);
nand U1943 (N_1943,N_1061,N_1307);
nor U1944 (N_1944,N_1315,N_1415);
and U1945 (N_1945,N_1031,N_1432);
or U1946 (N_1946,N_1240,N_1360);
and U1947 (N_1947,N_1142,N_1240);
or U1948 (N_1948,N_1080,N_1471);
nor U1949 (N_1949,N_1260,N_1369);
nand U1950 (N_1950,N_1365,N_1467);
nor U1951 (N_1951,N_1320,N_1142);
or U1952 (N_1952,N_1497,N_1124);
nor U1953 (N_1953,N_1033,N_1419);
nand U1954 (N_1954,N_1480,N_1256);
and U1955 (N_1955,N_1278,N_1310);
nor U1956 (N_1956,N_1013,N_1422);
or U1957 (N_1957,N_1132,N_1492);
nor U1958 (N_1958,N_1201,N_1329);
or U1959 (N_1959,N_1453,N_1010);
nand U1960 (N_1960,N_1429,N_1168);
or U1961 (N_1961,N_1297,N_1062);
nand U1962 (N_1962,N_1260,N_1150);
nor U1963 (N_1963,N_1267,N_1129);
nor U1964 (N_1964,N_1115,N_1054);
and U1965 (N_1965,N_1351,N_1263);
nor U1966 (N_1966,N_1474,N_1041);
nor U1967 (N_1967,N_1087,N_1177);
nor U1968 (N_1968,N_1014,N_1193);
nand U1969 (N_1969,N_1087,N_1225);
nor U1970 (N_1970,N_1232,N_1323);
nor U1971 (N_1971,N_1119,N_1463);
or U1972 (N_1972,N_1397,N_1069);
and U1973 (N_1973,N_1058,N_1435);
and U1974 (N_1974,N_1197,N_1203);
xnor U1975 (N_1975,N_1263,N_1366);
xnor U1976 (N_1976,N_1105,N_1074);
and U1977 (N_1977,N_1389,N_1403);
nand U1978 (N_1978,N_1035,N_1444);
nor U1979 (N_1979,N_1112,N_1194);
nand U1980 (N_1980,N_1020,N_1056);
nor U1981 (N_1981,N_1031,N_1262);
or U1982 (N_1982,N_1003,N_1014);
and U1983 (N_1983,N_1362,N_1380);
nand U1984 (N_1984,N_1177,N_1068);
and U1985 (N_1985,N_1192,N_1491);
nand U1986 (N_1986,N_1251,N_1360);
and U1987 (N_1987,N_1094,N_1364);
nor U1988 (N_1988,N_1303,N_1042);
nand U1989 (N_1989,N_1104,N_1386);
xor U1990 (N_1990,N_1175,N_1044);
and U1991 (N_1991,N_1350,N_1456);
xor U1992 (N_1992,N_1027,N_1314);
and U1993 (N_1993,N_1425,N_1149);
nor U1994 (N_1994,N_1148,N_1323);
nand U1995 (N_1995,N_1083,N_1173);
and U1996 (N_1996,N_1484,N_1261);
nor U1997 (N_1997,N_1197,N_1024);
or U1998 (N_1998,N_1334,N_1324);
nand U1999 (N_1999,N_1365,N_1318);
nand U2000 (N_2000,N_1985,N_1884);
xnor U2001 (N_2001,N_1777,N_1801);
xor U2002 (N_2002,N_1935,N_1946);
and U2003 (N_2003,N_1846,N_1864);
nand U2004 (N_2004,N_1664,N_1829);
xor U2005 (N_2005,N_1578,N_1926);
nor U2006 (N_2006,N_1780,N_1530);
or U2007 (N_2007,N_1959,N_1599);
nand U2008 (N_2008,N_1845,N_1942);
nand U2009 (N_2009,N_1533,N_1671);
xor U2010 (N_2010,N_1859,N_1726);
and U2011 (N_2011,N_1774,N_1873);
xor U2012 (N_2012,N_1830,N_1644);
and U2013 (N_2013,N_1963,N_1584);
or U2014 (N_2014,N_1746,N_1535);
nand U2015 (N_2015,N_1580,N_1814);
nand U2016 (N_2016,N_1922,N_1849);
nor U2017 (N_2017,N_1760,N_1765);
or U2018 (N_2018,N_1515,N_1994);
and U2019 (N_2019,N_1811,N_1508);
xor U2020 (N_2020,N_1800,N_1835);
nor U2021 (N_2021,N_1501,N_1652);
nand U2022 (N_2022,N_1653,N_1502);
and U2023 (N_2023,N_1895,N_1917);
nor U2024 (N_2024,N_1853,N_1976);
and U2025 (N_2025,N_1860,N_1759);
and U2026 (N_2026,N_1719,N_1862);
and U2027 (N_2027,N_1991,N_1907);
nand U2028 (N_2028,N_1758,N_1891);
xor U2029 (N_2029,N_1747,N_1617);
and U2030 (N_2030,N_1544,N_1868);
or U2031 (N_2031,N_1978,N_1951);
and U2032 (N_2032,N_1673,N_1661);
nand U2033 (N_2033,N_1950,N_1945);
or U2034 (N_2034,N_1659,N_1754);
or U2035 (N_2035,N_1875,N_1893);
nand U2036 (N_2036,N_1904,N_1972);
xor U2037 (N_2037,N_1813,N_1771);
and U2038 (N_2038,N_1697,N_1700);
nand U2039 (N_2039,N_1648,N_1822);
nand U2040 (N_2040,N_1762,N_1626);
nand U2041 (N_2041,N_1756,N_1637);
nor U2042 (N_2042,N_1952,N_1748);
nand U2043 (N_2043,N_1795,N_1657);
or U2044 (N_2044,N_1979,N_1753);
or U2045 (N_2045,N_1755,N_1647);
nor U2046 (N_2046,N_1931,N_1715);
nand U2047 (N_2047,N_1910,N_1990);
nand U2048 (N_2048,N_1505,N_1730);
nor U2049 (N_2049,N_1890,N_1871);
nand U2050 (N_2050,N_1838,N_1908);
or U2051 (N_2051,N_1670,N_1779);
or U2052 (N_2052,N_1510,N_1769);
and U2053 (N_2053,N_1820,N_1679);
and U2054 (N_2054,N_1596,N_1770);
nor U2055 (N_2055,N_1782,N_1609);
and U2056 (N_2056,N_1621,N_1879);
nand U2057 (N_2057,N_1579,N_1555);
nor U2058 (N_2058,N_1526,N_1943);
nand U2059 (N_2059,N_1553,N_1713);
or U2060 (N_2060,N_1752,N_1523);
nand U2061 (N_2061,N_1764,N_1568);
nand U2062 (N_2062,N_1655,N_1678);
nor U2063 (N_2063,N_1767,N_1642);
or U2064 (N_2064,N_1902,N_1792);
xor U2065 (N_2065,N_1744,N_1799);
xnor U2066 (N_2066,N_1798,N_1882);
nand U2067 (N_2067,N_1723,N_1545);
and U2068 (N_2068,N_1724,N_1582);
nand U2069 (N_2069,N_1714,N_1870);
or U2070 (N_2070,N_1881,N_1690);
nand U2071 (N_2071,N_1939,N_1852);
nor U2072 (N_2072,N_1923,N_1831);
nand U2073 (N_2073,N_1768,N_1572);
nor U2074 (N_2074,N_1815,N_1836);
nor U2075 (N_2075,N_1825,N_1929);
or U2076 (N_2076,N_1589,N_1731);
or U2077 (N_2077,N_1969,N_1808);
or U2078 (N_2078,N_1785,N_1522);
nand U2079 (N_2079,N_1818,N_1934);
and U2080 (N_2080,N_1745,N_1970);
or U2081 (N_2081,N_1741,N_1751);
nand U2082 (N_2082,N_1672,N_1602);
or U2083 (N_2083,N_1840,N_1682);
and U2084 (N_2084,N_1761,N_1608);
nand U2085 (N_2085,N_1577,N_1607);
and U2086 (N_2086,N_1680,N_1689);
and U2087 (N_2087,N_1720,N_1900);
nand U2088 (N_2088,N_1911,N_1973);
nand U2089 (N_2089,N_1532,N_1790);
or U2090 (N_2090,N_1841,N_1666);
nor U2091 (N_2091,N_1695,N_1827);
xor U2092 (N_2092,N_1927,N_1658);
or U2093 (N_2093,N_1773,N_1603);
xor U2094 (N_2094,N_1967,N_1901);
and U2095 (N_2095,N_1867,N_1512);
and U2096 (N_2096,N_1699,N_1639);
nor U2097 (N_2097,N_1591,N_1737);
nor U2098 (N_2098,N_1735,N_1948);
and U2099 (N_2099,N_1665,N_1620);
or U2100 (N_2100,N_1826,N_1614);
nor U2101 (N_2101,N_1615,N_1616);
or U2102 (N_2102,N_1783,N_1855);
or U2103 (N_2103,N_1576,N_1804);
nand U2104 (N_2104,N_1581,N_1966);
or U2105 (N_2105,N_1992,N_1705);
nor U2106 (N_2106,N_1877,N_1691);
and U2107 (N_2107,N_1736,N_1763);
or U2108 (N_2108,N_1794,N_1633);
or U2109 (N_2109,N_1850,N_1560);
and U2110 (N_2110,N_1725,N_1776);
nor U2111 (N_2111,N_1681,N_1539);
and U2112 (N_2112,N_1880,N_1778);
or U2113 (N_2113,N_1663,N_1806);
nand U2114 (N_2114,N_1612,N_1885);
nand U2115 (N_2115,N_1909,N_1983);
nor U2116 (N_2116,N_1551,N_1878);
nor U2117 (N_2117,N_1817,N_1722);
nor U2118 (N_2118,N_1604,N_1623);
and U2119 (N_2119,N_1631,N_1993);
nor U2120 (N_2120,N_1977,N_1894);
or U2121 (N_2121,N_1613,N_1660);
and U2122 (N_2122,N_1872,N_1667);
xnor U2123 (N_2123,N_1635,N_1574);
nand U2124 (N_2124,N_1843,N_1823);
and U2125 (N_2125,N_1955,N_1688);
or U2126 (N_2126,N_1793,N_1645);
nand U2127 (N_2127,N_1554,N_1636);
and U2128 (N_2128,N_1619,N_1940);
nor U2129 (N_2129,N_1598,N_1938);
and U2130 (N_2130,N_1742,N_1587);
and U2131 (N_2131,N_1564,N_1932);
nand U2132 (N_2132,N_1865,N_1651);
or U2133 (N_2133,N_1721,N_1692);
nor U2134 (N_2134,N_1789,N_1874);
nand U2135 (N_2135,N_1915,N_1707);
or U2136 (N_2136,N_1772,N_1944);
and U2137 (N_2137,N_1540,N_1937);
nor U2138 (N_2138,N_1941,N_1858);
and U2139 (N_2139,N_1677,N_1650);
xnor U2140 (N_2140,N_1567,N_1669);
nand U2141 (N_2141,N_1590,N_1962);
or U2142 (N_2142,N_1674,N_1654);
or U2143 (N_2143,N_1834,N_1866);
xnor U2144 (N_2144,N_1916,N_1987);
or U2145 (N_2145,N_1861,N_1750);
and U2146 (N_2146,N_1525,N_1628);
nand U2147 (N_2147,N_1733,N_1982);
and U2148 (N_2148,N_1989,N_1953);
nor U2149 (N_2149,N_1583,N_1848);
or U2150 (N_2150,N_1729,N_1738);
nand U2151 (N_2151,N_1988,N_1912);
nor U2152 (N_2152,N_1588,N_1784);
nand U2153 (N_2153,N_1629,N_1562);
nor U2154 (N_2154,N_1698,N_1534);
and U2155 (N_2155,N_1928,N_1566);
or U2156 (N_2156,N_1824,N_1837);
nand U2157 (N_2157,N_1610,N_1775);
nand U2158 (N_2158,N_1503,N_1593);
nand U2159 (N_2159,N_1625,N_1570);
xnor U2160 (N_2160,N_1640,N_1821);
nor U2161 (N_2161,N_1518,N_1743);
or U2162 (N_2162,N_1734,N_1529);
and U2163 (N_2163,N_1749,N_1857);
nand U2164 (N_2164,N_1624,N_1936);
nor U2165 (N_2165,N_1847,N_1693);
or U2166 (N_2166,N_1513,N_1556);
nand U2167 (N_2167,N_1844,N_1531);
and U2168 (N_2168,N_1924,N_1524);
nor U2169 (N_2169,N_1543,N_1981);
nor U2170 (N_2170,N_1728,N_1630);
xor U2171 (N_2171,N_1507,N_1896);
and U2172 (N_2172,N_1797,N_1727);
and U2173 (N_2173,N_1717,N_1905);
nor U2174 (N_2174,N_1632,N_1833);
nor U2175 (N_2175,N_1984,N_1996);
nor U2176 (N_2176,N_1965,N_1899);
nand U2177 (N_2177,N_1914,N_1999);
or U2178 (N_2178,N_1892,N_1686);
nor U2179 (N_2179,N_1887,N_1611);
and U2180 (N_2180,N_1883,N_1732);
nor U2181 (N_2181,N_1803,N_1668);
nor U2182 (N_2182,N_1514,N_1696);
and U2183 (N_2183,N_1930,N_1649);
or U2184 (N_2184,N_1561,N_1646);
and U2185 (N_2185,N_1920,N_1956);
nand U2186 (N_2186,N_1605,N_1863);
and U2187 (N_2187,N_1684,N_1839);
and U2188 (N_2188,N_1563,N_1791);
nand U2189 (N_2189,N_1516,N_1933);
nand U2190 (N_2190,N_1842,N_1676);
and U2191 (N_2191,N_1569,N_1675);
and U2192 (N_2192,N_1627,N_1519);
nand U2193 (N_2193,N_1706,N_1997);
xnor U2194 (N_2194,N_1802,N_1704);
nand U2195 (N_2195,N_1711,N_1573);
and U2196 (N_2196,N_1964,N_1968);
nor U2197 (N_2197,N_1541,N_1788);
nor U2198 (N_2198,N_1549,N_1716);
nand U2199 (N_2199,N_1876,N_1906);
xor U2200 (N_2200,N_1954,N_1638);
and U2201 (N_2201,N_1919,N_1851);
nor U2202 (N_2202,N_1537,N_1509);
nor U2203 (N_2203,N_1662,N_1781);
and U2204 (N_2204,N_1856,N_1961);
and U2205 (N_2205,N_1558,N_1897);
and U2206 (N_2206,N_1527,N_1592);
xnor U2207 (N_2207,N_1957,N_1595);
or U2208 (N_2208,N_1712,N_1918);
nor U2209 (N_2209,N_1656,N_1601);
and U2210 (N_2210,N_1618,N_1889);
xor U2211 (N_2211,N_1766,N_1812);
nand U2212 (N_2212,N_1528,N_1807);
nand U2213 (N_2213,N_1739,N_1709);
and U2214 (N_2214,N_1974,N_1980);
or U2215 (N_2215,N_1913,N_1557);
and U2216 (N_2216,N_1542,N_1520);
and U2217 (N_2217,N_1995,N_1548);
nor U2218 (N_2218,N_1643,N_1809);
nor U2219 (N_2219,N_1854,N_1546);
xnor U2220 (N_2220,N_1685,N_1622);
and U2221 (N_2221,N_1694,N_1786);
nand U2222 (N_2222,N_1921,N_1559);
nor U2223 (N_2223,N_1586,N_1998);
nand U2224 (N_2224,N_1757,N_1975);
or U2225 (N_2225,N_1634,N_1703);
xnor U2226 (N_2226,N_1506,N_1600);
or U2227 (N_2227,N_1949,N_1550);
nor U2228 (N_2228,N_1816,N_1585);
and U2229 (N_2229,N_1538,N_1504);
and U2230 (N_2230,N_1869,N_1710);
or U2231 (N_2231,N_1832,N_1960);
nand U2232 (N_2232,N_1925,N_1971);
or U2233 (N_2233,N_1571,N_1606);
or U2234 (N_2234,N_1597,N_1958);
nor U2235 (N_2235,N_1701,N_1500);
or U2236 (N_2236,N_1986,N_1718);
xor U2237 (N_2237,N_1947,N_1565);
nor U2238 (N_2238,N_1787,N_1511);
and U2239 (N_2239,N_1702,N_1687);
or U2240 (N_2240,N_1536,N_1886);
nor U2241 (N_2241,N_1805,N_1594);
xnor U2242 (N_2242,N_1575,N_1903);
nand U2243 (N_2243,N_1641,N_1521);
and U2244 (N_2244,N_1683,N_1828);
or U2245 (N_2245,N_1517,N_1810);
nand U2246 (N_2246,N_1740,N_1552);
nand U2247 (N_2247,N_1547,N_1898);
xnor U2248 (N_2248,N_1819,N_1708);
nor U2249 (N_2249,N_1888,N_1796);
nor U2250 (N_2250,N_1684,N_1535);
and U2251 (N_2251,N_1658,N_1887);
nand U2252 (N_2252,N_1688,N_1857);
nand U2253 (N_2253,N_1846,N_1878);
and U2254 (N_2254,N_1744,N_1990);
and U2255 (N_2255,N_1943,N_1750);
or U2256 (N_2256,N_1808,N_1840);
or U2257 (N_2257,N_1957,N_1995);
and U2258 (N_2258,N_1528,N_1808);
or U2259 (N_2259,N_1720,N_1951);
or U2260 (N_2260,N_1915,N_1763);
and U2261 (N_2261,N_1945,N_1894);
nand U2262 (N_2262,N_1721,N_1775);
nor U2263 (N_2263,N_1665,N_1617);
and U2264 (N_2264,N_1914,N_1819);
or U2265 (N_2265,N_1608,N_1556);
or U2266 (N_2266,N_1831,N_1868);
and U2267 (N_2267,N_1835,N_1518);
or U2268 (N_2268,N_1604,N_1708);
and U2269 (N_2269,N_1574,N_1787);
and U2270 (N_2270,N_1938,N_1701);
nor U2271 (N_2271,N_1685,N_1681);
nor U2272 (N_2272,N_1690,N_1860);
nor U2273 (N_2273,N_1785,N_1932);
nor U2274 (N_2274,N_1722,N_1705);
nand U2275 (N_2275,N_1973,N_1765);
nand U2276 (N_2276,N_1903,N_1555);
and U2277 (N_2277,N_1761,N_1697);
and U2278 (N_2278,N_1738,N_1836);
or U2279 (N_2279,N_1778,N_1886);
nor U2280 (N_2280,N_1945,N_1804);
and U2281 (N_2281,N_1782,N_1766);
and U2282 (N_2282,N_1618,N_1653);
and U2283 (N_2283,N_1996,N_1549);
nor U2284 (N_2284,N_1678,N_1834);
or U2285 (N_2285,N_1609,N_1640);
nand U2286 (N_2286,N_1577,N_1784);
or U2287 (N_2287,N_1797,N_1569);
xor U2288 (N_2288,N_1975,N_1685);
nand U2289 (N_2289,N_1700,N_1706);
and U2290 (N_2290,N_1640,N_1858);
or U2291 (N_2291,N_1531,N_1972);
and U2292 (N_2292,N_1703,N_1901);
nand U2293 (N_2293,N_1584,N_1790);
nor U2294 (N_2294,N_1875,N_1723);
and U2295 (N_2295,N_1767,N_1835);
xor U2296 (N_2296,N_1882,N_1932);
and U2297 (N_2297,N_1861,N_1981);
nor U2298 (N_2298,N_1540,N_1862);
nor U2299 (N_2299,N_1972,N_1815);
xor U2300 (N_2300,N_1971,N_1630);
or U2301 (N_2301,N_1932,N_1747);
and U2302 (N_2302,N_1889,N_1898);
nor U2303 (N_2303,N_1773,N_1556);
nand U2304 (N_2304,N_1929,N_1587);
nand U2305 (N_2305,N_1979,N_1645);
and U2306 (N_2306,N_1719,N_1829);
and U2307 (N_2307,N_1533,N_1527);
nor U2308 (N_2308,N_1593,N_1920);
nor U2309 (N_2309,N_1513,N_1791);
nor U2310 (N_2310,N_1908,N_1527);
and U2311 (N_2311,N_1519,N_1561);
and U2312 (N_2312,N_1520,N_1719);
nor U2313 (N_2313,N_1522,N_1896);
nand U2314 (N_2314,N_1724,N_1820);
or U2315 (N_2315,N_1739,N_1877);
or U2316 (N_2316,N_1739,N_1929);
xnor U2317 (N_2317,N_1819,N_1666);
or U2318 (N_2318,N_1674,N_1588);
and U2319 (N_2319,N_1834,N_1619);
nor U2320 (N_2320,N_1980,N_1710);
nor U2321 (N_2321,N_1875,N_1583);
nand U2322 (N_2322,N_1968,N_1930);
and U2323 (N_2323,N_1927,N_1793);
nor U2324 (N_2324,N_1744,N_1574);
nor U2325 (N_2325,N_1989,N_1849);
and U2326 (N_2326,N_1689,N_1926);
or U2327 (N_2327,N_1659,N_1826);
or U2328 (N_2328,N_1649,N_1894);
nor U2329 (N_2329,N_1712,N_1708);
or U2330 (N_2330,N_1735,N_1802);
nand U2331 (N_2331,N_1816,N_1690);
nand U2332 (N_2332,N_1676,N_1678);
nand U2333 (N_2333,N_1917,N_1809);
xor U2334 (N_2334,N_1770,N_1572);
and U2335 (N_2335,N_1545,N_1663);
xnor U2336 (N_2336,N_1975,N_1977);
or U2337 (N_2337,N_1642,N_1918);
and U2338 (N_2338,N_1530,N_1948);
nand U2339 (N_2339,N_1887,N_1710);
or U2340 (N_2340,N_1971,N_1618);
nand U2341 (N_2341,N_1545,N_1909);
nor U2342 (N_2342,N_1748,N_1793);
nor U2343 (N_2343,N_1946,N_1819);
xnor U2344 (N_2344,N_1912,N_1903);
and U2345 (N_2345,N_1943,N_1710);
nand U2346 (N_2346,N_1802,N_1958);
and U2347 (N_2347,N_1832,N_1805);
nor U2348 (N_2348,N_1925,N_1862);
nor U2349 (N_2349,N_1739,N_1803);
or U2350 (N_2350,N_1782,N_1971);
and U2351 (N_2351,N_1509,N_1620);
nand U2352 (N_2352,N_1541,N_1621);
nand U2353 (N_2353,N_1671,N_1897);
nor U2354 (N_2354,N_1887,N_1908);
or U2355 (N_2355,N_1851,N_1951);
xor U2356 (N_2356,N_1805,N_1847);
nand U2357 (N_2357,N_1519,N_1860);
or U2358 (N_2358,N_1540,N_1585);
nor U2359 (N_2359,N_1778,N_1740);
and U2360 (N_2360,N_1798,N_1797);
and U2361 (N_2361,N_1629,N_1805);
nand U2362 (N_2362,N_1806,N_1639);
or U2363 (N_2363,N_1611,N_1988);
nand U2364 (N_2364,N_1866,N_1572);
xor U2365 (N_2365,N_1637,N_1821);
xnor U2366 (N_2366,N_1711,N_1802);
nor U2367 (N_2367,N_1589,N_1734);
nor U2368 (N_2368,N_1891,N_1632);
xnor U2369 (N_2369,N_1666,N_1739);
nand U2370 (N_2370,N_1688,N_1596);
nor U2371 (N_2371,N_1964,N_1845);
or U2372 (N_2372,N_1883,N_1801);
nor U2373 (N_2373,N_1949,N_1888);
nand U2374 (N_2374,N_1780,N_1556);
nor U2375 (N_2375,N_1835,N_1841);
and U2376 (N_2376,N_1958,N_1937);
and U2377 (N_2377,N_1601,N_1598);
or U2378 (N_2378,N_1892,N_1607);
nor U2379 (N_2379,N_1565,N_1712);
nand U2380 (N_2380,N_1524,N_1802);
xnor U2381 (N_2381,N_1795,N_1868);
or U2382 (N_2382,N_1504,N_1889);
nor U2383 (N_2383,N_1862,N_1647);
nand U2384 (N_2384,N_1966,N_1708);
and U2385 (N_2385,N_1717,N_1842);
nor U2386 (N_2386,N_1992,N_1502);
nor U2387 (N_2387,N_1845,N_1841);
nor U2388 (N_2388,N_1680,N_1724);
nand U2389 (N_2389,N_1857,N_1661);
and U2390 (N_2390,N_1628,N_1880);
and U2391 (N_2391,N_1523,N_1759);
or U2392 (N_2392,N_1837,N_1828);
and U2393 (N_2393,N_1698,N_1862);
and U2394 (N_2394,N_1866,N_1841);
nand U2395 (N_2395,N_1812,N_1784);
nand U2396 (N_2396,N_1918,N_1942);
and U2397 (N_2397,N_1994,N_1975);
nand U2398 (N_2398,N_1723,N_1993);
nand U2399 (N_2399,N_1595,N_1762);
and U2400 (N_2400,N_1821,N_1927);
nor U2401 (N_2401,N_1785,N_1511);
nor U2402 (N_2402,N_1590,N_1919);
and U2403 (N_2403,N_1925,N_1874);
nand U2404 (N_2404,N_1754,N_1631);
and U2405 (N_2405,N_1653,N_1738);
and U2406 (N_2406,N_1554,N_1912);
and U2407 (N_2407,N_1697,N_1691);
nor U2408 (N_2408,N_1610,N_1718);
nor U2409 (N_2409,N_1535,N_1993);
nand U2410 (N_2410,N_1755,N_1526);
or U2411 (N_2411,N_1696,N_1650);
nor U2412 (N_2412,N_1558,N_1938);
xnor U2413 (N_2413,N_1979,N_1688);
nand U2414 (N_2414,N_1574,N_1995);
nand U2415 (N_2415,N_1557,N_1894);
or U2416 (N_2416,N_1586,N_1740);
or U2417 (N_2417,N_1706,N_1604);
nor U2418 (N_2418,N_1853,N_1673);
and U2419 (N_2419,N_1572,N_1638);
and U2420 (N_2420,N_1741,N_1558);
nand U2421 (N_2421,N_1585,N_1677);
and U2422 (N_2422,N_1550,N_1895);
nand U2423 (N_2423,N_1730,N_1998);
and U2424 (N_2424,N_1638,N_1562);
nand U2425 (N_2425,N_1727,N_1693);
and U2426 (N_2426,N_1715,N_1517);
xnor U2427 (N_2427,N_1659,N_1544);
nand U2428 (N_2428,N_1676,N_1541);
nand U2429 (N_2429,N_1962,N_1785);
nand U2430 (N_2430,N_1742,N_1915);
nand U2431 (N_2431,N_1502,N_1945);
nand U2432 (N_2432,N_1652,N_1894);
or U2433 (N_2433,N_1720,N_1744);
nand U2434 (N_2434,N_1799,N_1552);
or U2435 (N_2435,N_1606,N_1759);
nor U2436 (N_2436,N_1623,N_1944);
nor U2437 (N_2437,N_1760,N_1660);
nor U2438 (N_2438,N_1908,N_1935);
and U2439 (N_2439,N_1738,N_1688);
and U2440 (N_2440,N_1824,N_1635);
or U2441 (N_2441,N_1878,N_1983);
nand U2442 (N_2442,N_1905,N_1588);
nand U2443 (N_2443,N_1622,N_1876);
and U2444 (N_2444,N_1803,N_1595);
nor U2445 (N_2445,N_1593,N_1993);
and U2446 (N_2446,N_1765,N_1784);
xor U2447 (N_2447,N_1612,N_1536);
nand U2448 (N_2448,N_1969,N_1764);
or U2449 (N_2449,N_1753,N_1964);
xor U2450 (N_2450,N_1773,N_1959);
or U2451 (N_2451,N_1826,N_1688);
xor U2452 (N_2452,N_1658,N_1621);
or U2453 (N_2453,N_1944,N_1840);
or U2454 (N_2454,N_1854,N_1992);
nor U2455 (N_2455,N_1779,N_1821);
nand U2456 (N_2456,N_1830,N_1520);
or U2457 (N_2457,N_1888,N_1704);
or U2458 (N_2458,N_1891,N_1538);
and U2459 (N_2459,N_1792,N_1536);
or U2460 (N_2460,N_1837,N_1759);
or U2461 (N_2461,N_1523,N_1644);
or U2462 (N_2462,N_1650,N_1501);
nand U2463 (N_2463,N_1627,N_1668);
nand U2464 (N_2464,N_1980,N_1571);
nor U2465 (N_2465,N_1566,N_1851);
and U2466 (N_2466,N_1972,N_1835);
nand U2467 (N_2467,N_1809,N_1739);
and U2468 (N_2468,N_1669,N_1863);
or U2469 (N_2469,N_1935,N_1771);
xnor U2470 (N_2470,N_1828,N_1972);
nand U2471 (N_2471,N_1686,N_1640);
and U2472 (N_2472,N_1919,N_1571);
and U2473 (N_2473,N_1627,N_1666);
and U2474 (N_2474,N_1923,N_1898);
xnor U2475 (N_2475,N_1597,N_1753);
nand U2476 (N_2476,N_1874,N_1632);
xnor U2477 (N_2477,N_1860,N_1526);
nor U2478 (N_2478,N_1823,N_1927);
nor U2479 (N_2479,N_1755,N_1731);
or U2480 (N_2480,N_1641,N_1529);
nand U2481 (N_2481,N_1718,N_1638);
nand U2482 (N_2482,N_1961,N_1798);
nand U2483 (N_2483,N_1559,N_1962);
or U2484 (N_2484,N_1643,N_1508);
nand U2485 (N_2485,N_1630,N_1584);
nand U2486 (N_2486,N_1767,N_1994);
nand U2487 (N_2487,N_1941,N_1677);
nor U2488 (N_2488,N_1566,N_1710);
nor U2489 (N_2489,N_1999,N_1635);
or U2490 (N_2490,N_1799,N_1752);
and U2491 (N_2491,N_1895,N_1748);
and U2492 (N_2492,N_1658,N_1811);
nand U2493 (N_2493,N_1844,N_1982);
and U2494 (N_2494,N_1888,N_1565);
nand U2495 (N_2495,N_1948,N_1890);
xnor U2496 (N_2496,N_1949,N_1865);
or U2497 (N_2497,N_1990,N_1624);
and U2498 (N_2498,N_1568,N_1713);
or U2499 (N_2499,N_1872,N_1946);
and U2500 (N_2500,N_2049,N_2297);
nor U2501 (N_2501,N_2265,N_2310);
and U2502 (N_2502,N_2097,N_2336);
nor U2503 (N_2503,N_2398,N_2025);
nor U2504 (N_2504,N_2114,N_2161);
and U2505 (N_2505,N_2158,N_2242);
and U2506 (N_2506,N_2477,N_2475);
nor U2507 (N_2507,N_2276,N_2246);
nand U2508 (N_2508,N_2466,N_2442);
nor U2509 (N_2509,N_2355,N_2459);
nor U2510 (N_2510,N_2261,N_2122);
nor U2511 (N_2511,N_2068,N_2282);
and U2512 (N_2512,N_2417,N_2176);
and U2513 (N_2513,N_2094,N_2160);
nor U2514 (N_2514,N_2346,N_2362);
nand U2515 (N_2515,N_2418,N_2035);
and U2516 (N_2516,N_2038,N_2012);
nor U2517 (N_2517,N_2199,N_2054);
or U2518 (N_2518,N_2013,N_2472);
nor U2519 (N_2519,N_2034,N_2145);
or U2520 (N_2520,N_2020,N_2167);
or U2521 (N_2521,N_2454,N_2345);
nor U2522 (N_2522,N_2298,N_2203);
or U2523 (N_2523,N_2439,N_2016);
or U2524 (N_2524,N_2092,N_2209);
or U2525 (N_2525,N_2048,N_2385);
and U2526 (N_2526,N_2070,N_2351);
or U2527 (N_2527,N_2347,N_2078);
and U2528 (N_2528,N_2372,N_2189);
nor U2529 (N_2529,N_2350,N_2273);
or U2530 (N_2530,N_2124,N_2118);
nand U2531 (N_2531,N_2131,N_2208);
xnor U2532 (N_2532,N_2060,N_2028);
nor U2533 (N_2533,N_2381,N_2178);
xnor U2534 (N_2534,N_2322,N_2149);
nand U2535 (N_2535,N_2264,N_2043);
or U2536 (N_2536,N_2415,N_2295);
and U2537 (N_2537,N_2134,N_2349);
xnor U2538 (N_2538,N_2227,N_2460);
nand U2539 (N_2539,N_2109,N_2206);
nand U2540 (N_2540,N_2168,N_2403);
and U2541 (N_2541,N_2247,N_2443);
nand U2542 (N_2542,N_2011,N_2154);
nor U2543 (N_2543,N_2366,N_2485);
or U2544 (N_2544,N_2027,N_2329);
nand U2545 (N_2545,N_2113,N_2159);
and U2546 (N_2546,N_2179,N_2087);
xnor U2547 (N_2547,N_2422,N_2104);
and U2548 (N_2548,N_2486,N_2008);
or U2549 (N_2549,N_2093,N_2238);
xor U2550 (N_2550,N_2000,N_2338);
nand U2551 (N_2551,N_2467,N_2047);
or U2552 (N_2552,N_2280,N_2374);
or U2553 (N_2553,N_2434,N_2389);
and U2554 (N_2554,N_2191,N_2436);
or U2555 (N_2555,N_2481,N_2074);
or U2556 (N_2556,N_2296,N_2402);
nand U2557 (N_2557,N_2042,N_2305);
or U2558 (N_2558,N_2435,N_2218);
and U2559 (N_2559,N_2153,N_2059);
nor U2560 (N_2560,N_2450,N_2330);
or U2561 (N_2561,N_2077,N_2235);
xnor U2562 (N_2562,N_2195,N_2036);
nand U2563 (N_2563,N_2480,N_2021);
nand U2564 (N_2564,N_2210,N_2185);
xnor U2565 (N_2565,N_2215,N_2063);
nor U2566 (N_2566,N_2431,N_2323);
nand U2567 (N_2567,N_2426,N_2052);
nor U2568 (N_2568,N_2483,N_2111);
nor U2569 (N_2569,N_2250,N_2232);
or U2570 (N_2570,N_2157,N_2237);
or U2571 (N_2571,N_2339,N_2465);
xnor U2572 (N_2572,N_2233,N_2286);
nand U2573 (N_2573,N_2207,N_2437);
and U2574 (N_2574,N_2184,N_2311);
nand U2575 (N_2575,N_2123,N_2230);
and U2576 (N_2576,N_2337,N_2190);
xnor U2577 (N_2577,N_2066,N_2173);
or U2578 (N_2578,N_2395,N_2102);
nand U2579 (N_2579,N_2119,N_2086);
nand U2580 (N_2580,N_2169,N_2107);
and U2581 (N_2581,N_2257,N_2138);
or U2582 (N_2582,N_2262,N_2427);
or U2583 (N_2583,N_2129,N_2005);
nand U2584 (N_2584,N_2175,N_2499);
nand U2585 (N_2585,N_2320,N_2010);
xor U2586 (N_2586,N_2388,N_2284);
or U2587 (N_2587,N_2044,N_2018);
nand U2588 (N_2588,N_2002,N_2384);
or U2589 (N_2589,N_2105,N_2463);
nor U2590 (N_2590,N_2363,N_2127);
nand U2591 (N_2591,N_2164,N_2268);
nand U2592 (N_2592,N_2429,N_2380);
nand U2593 (N_2593,N_2015,N_2353);
nor U2594 (N_2594,N_2003,N_2306);
nand U2595 (N_2595,N_2260,N_2067);
xnor U2596 (N_2596,N_2419,N_2019);
or U2597 (N_2597,N_2244,N_2072);
nor U2598 (N_2598,N_2030,N_2468);
and U2599 (N_2599,N_2430,N_2132);
and U2600 (N_2600,N_2332,N_2056);
or U2601 (N_2601,N_2302,N_2331);
or U2602 (N_2602,N_2196,N_2461);
nor U2603 (N_2603,N_2075,N_2083);
nand U2604 (N_2604,N_2391,N_2292);
and U2605 (N_2605,N_2299,N_2407);
xor U2606 (N_2606,N_2228,N_2361);
nor U2607 (N_2607,N_2263,N_2394);
nor U2608 (N_2608,N_2281,N_2474);
and U2609 (N_2609,N_2112,N_2289);
or U2610 (N_2610,N_2492,N_2200);
and U2611 (N_2611,N_2014,N_2476);
nand U2612 (N_2612,N_2141,N_2152);
nor U2613 (N_2613,N_2006,N_2342);
xnor U2614 (N_2614,N_2321,N_2441);
and U2615 (N_2615,N_2307,N_2193);
xor U2616 (N_2616,N_2071,N_2090);
and U2617 (N_2617,N_2423,N_2009);
or U2618 (N_2618,N_2236,N_2377);
and U2619 (N_2619,N_2098,N_2358);
and U2620 (N_2620,N_2221,N_2414);
and U2621 (N_2621,N_2166,N_2309);
nand U2622 (N_2622,N_2393,N_2082);
nor U2623 (N_2623,N_2103,N_2490);
xnor U2624 (N_2624,N_2137,N_2354);
xor U2625 (N_2625,N_2272,N_2359);
nor U2626 (N_2626,N_2404,N_2458);
and U2627 (N_2627,N_2065,N_2294);
nor U2628 (N_2628,N_2115,N_2327);
nand U2629 (N_2629,N_2340,N_2088);
or U2630 (N_2630,N_2438,N_2308);
nor U2631 (N_2631,N_2073,N_2051);
nand U2632 (N_2632,N_2448,N_2416);
xnor U2633 (N_2633,N_2379,N_2022);
or U2634 (N_2634,N_2186,N_2165);
nand U2635 (N_2635,N_2192,N_2187);
or U2636 (N_2636,N_2333,N_2026);
and U2637 (N_2637,N_2128,N_2266);
and U2638 (N_2638,N_2279,N_2446);
nand U2639 (N_2639,N_2285,N_2133);
nand U2640 (N_2640,N_2183,N_2151);
nor U2641 (N_2641,N_2357,N_2143);
nor U2642 (N_2642,N_2312,N_2081);
and U2643 (N_2643,N_2445,N_2375);
or U2644 (N_2644,N_2100,N_2277);
nor U2645 (N_2645,N_2456,N_2024);
or U2646 (N_2646,N_2300,N_2204);
and U2647 (N_2647,N_2494,N_2314);
and U2648 (N_2648,N_2291,N_2064);
nand U2649 (N_2649,N_2062,N_2479);
and U2650 (N_2650,N_2121,N_2313);
nand U2651 (N_2651,N_2211,N_2253);
or U2652 (N_2652,N_2224,N_2231);
nand U2653 (N_2653,N_2290,N_2489);
xnor U2654 (N_2654,N_2392,N_2045);
nor U2655 (N_2655,N_2162,N_2023);
or U2656 (N_2656,N_2373,N_2213);
xor U2657 (N_2657,N_2382,N_2447);
and U2658 (N_2658,N_2130,N_2155);
nand U2659 (N_2659,N_2258,N_2343);
nor U2660 (N_2660,N_2135,N_2239);
nor U2661 (N_2661,N_2455,N_2079);
nor U2662 (N_2662,N_2163,N_2469);
nand U2663 (N_2663,N_2144,N_2270);
nand U2664 (N_2664,N_2405,N_2096);
nand U2665 (N_2665,N_2400,N_2453);
nand U2666 (N_2666,N_2255,N_2488);
or U2667 (N_2667,N_2288,N_2069);
and U2668 (N_2668,N_2223,N_2214);
nor U2669 (N_2669,N_2198,N_2376);
or U2670 (N_2670,N_2371,N_2278);
and U2671 (N_2671,N_2116,N_2449);
and U2672 (N_2672,N_2039,N_2055);
nor U2673 (N_2673,N_2267,N_2147);
nor U2674 (N_2674,N_2348,N_2222);
xor U2675 (N_2675,N_2146,N_2220);
nor U2676 (N_2676,N_2029,N_2383);
xor U2677 (N_2677,N_2140,N_2058);
or U2678 (N_2678,N_2360,N_2365);
or U2679 (N_2679,N_2399,N_2080);
nor U2680 (N_2680,N_2462,N_2007);
nand U2681 (N_2681,N_2356,N_2219);
nand U2682 (N_2682,N_2188,N_2254);
xor U2683 (N_2683,N_2212,N_2170);
nor U2684 (N_2684,N_2205,N_2274);
nor U2685 (N_2685,N_2108,N_2241);
and U2686 (N_2686,N_2471,N_2110);
nand U2687 (N_2687,N_2197,N_2420);
nand U2688 (N_2688,N_2032,N_2271);
xnor U2689 (N_2689,N_2061,N_2495);
nand U2690 (N_2690,N_2352,N_2317);
and U2691 (N_2691,N_2370,N_2440);
nor U2692 (N_2692,N_2177,N_2301);
nand U2693 (N_2693,N_2136,N_2125);
xnor U2694 (N_2694,N_2180,N_2148);
nor U2695 (N_2695,N_2318,N_2303);
and U2696 (N_2696,N_2287,N_2139);
nand U2697 (N_2697,N_2491,N_2316);
and U2698 (N_2698,N_2275,N_2057);
nor U2699 (N_2699,N_2085,N_2259);
or U2700 (N_2700,N_2334,N_2243);
or U2701 (N_2701,N_2464,N_2150);
xnor U2702 (N_2702,N_2397,N_2451);
nor U2703 (N_2703,N_2106,N_2408);
or U2704 (N_2704,N_2304,N_2493);
or U2705 (N_2705,N_2248,N_2390);
nor U2706 (N_2706,N_2194,N_2487);
xnor U2707 (N_2707,N_2229,N_2174);
or U2708 (N_2708,N_2252,N_2324);
nand U2709 (N_2709,N_2410,N_2344);
nand U2710 (N_2710,N_2378,N_2367);
and U2711 (N_2711,N_2182,N_2269);
or U2712 (N_2712,N_2084,N_2293);
and U2713 (N_2713,N_2473,N_2181);
and U2714 (N_2714,N_2099,N_2484);
and U2715 (N_2715,N_2031,N_2033);
or U2716 (N_2716,N_2040,N_2171);
or U2717 (N_2717,N_2216,N_2457);
or U2718 (N_2718,N_2328,N_2341);
nand U2719 (N_2719,N_2283,N_2050);
nand U2720 (N_2720,N_2425,N_2041);
nor U2721 (N_2721,N_2406,N_2249);
xnor U2722 (N_2722,N_2217,N_2496);
and U2723 (N_2723,N_2401,N_2319);
nor U2724 (N_2724,N_2368,N_2315);
nand U2725 (N_2725,N_2498,N_2095);
or U2726 (N_2726,N_2424,N_2202);
and U2727 (N_2727,N_2364,N_2396);
or U2728 (N_2728,N_2245,N_2076);
or U2729 (N_2729,N_2142,N_2433);
or U2730 (N_2730,N_2412,N_2101);
nor U2731 (N_2731,N_2156,N_2326);
and U2732 (N_2732,N_2226,N_2428);
and U2733 (N_2733,N_2234,N_2117);
or U2734 (N_2734,N_2470,N_2120);
xor U2735 (N_2735,N_2201,N_2172);
nor U2736 (N_2736,N_2325,N_2037);
nand U2737 (N_2737,N_2409,N_2478);
or U2738 (N_2738,N_2251,N_2126);
and U2739 (N_2739,N_2225,N_2482);
xnor U2740 (N_2740,N_2386,N_2387);
nor U2741 (N_2741,N_2432,N_2497);
nor U2742 (N_2742,N_2444,N_2335);
nand U2743 (N_2743,N_2240,N_2046);
and U2744 (N_2744,N_2369,N_2089);
and U2745 (N_2745,N_2411,N_2421);
nor U2746 (N_2746,N_2413,N_2053);
or U2747 (N_2747,N_2452,N_2091);
and U2748 (N_2748,N_2001,N_2017);
nor U2749 (N_2749,N_2004,N_2256);
nand U2750 (N_2750,N_2376,N_2092);
nor U2751 (N_2751,N_2186,N_2161);
nand U2752 (N_2752,N_2491,N_2088);
nand U2753 (N_2753,N_2201,N_2336);
or U2754 (N_2754,N_2233,N_2393);
nor U2755 (N_2755,N_2070,N_2092);
and U2756 (N_2756,N_2067,N_2143);
xor U2757 (N_2757,N_2156,N_2292);
and U2758 (N_2758,N_2295,N_2416);
nor U2759 (N_2759,N_2087,N_2473);
and U2760 (N_2760,N_2084,N_2473);
xnor U2761 (N_2761,N_2344,N_2435);
nand U2762 (N_2762,N_2103,N_2162);
nand U2763 (N_2763,N_2368,N_2040);
nor U2764 (N_2764,N_2224,N_2456);
nand U2765 (N_2765,N_2222,N_2232);
or U2766 (N_2766,N_2021,N_2485);
nor U2767 (N_2767,N_2247,N_2462);
nand U2768 (N_2768,N_2253,N_2155);
xor U2769 (N_2769,N_2203,N_2077);
nor U2770 (N_2770,N_2002,N_2134);
or U2771 (N_2771,N_2202,N_2436);
and U2772 (N_2772,N_2277,N_2328);
nand U2773 (N_2773,N_2058,N_2351);
or U2774 (N_2774,N_2454,N_2315);
nand U2775 (N_2775,N_2115,N_2061);
and U2776 (N_2776,N_2225,N_2235);
nor U2777 (N_2777,N_2059,N_2125);
and U2778 (N_2778,N_2321,N_2073);
and U2779 (N_2779,N_2442,N_2018);
or U2780 (N_2780,N_2251,N_2233);
xor U2781 (N_2781,N_2435,N_2467);
or U2782 (N_2782,N_2399,N_2009);
nor U2783 (N_2783,N_2469,N_2175);
and U2784 (N_2784,N_2390,N_2121);
xor U2785 (N_2785,N_2150,N_2151);
or U2786 (N_2786,N_2320,N_2404);
or U2787 (N_2787,N_2347,N_2334);
xnor U2788 (N_2788,N_2002,N_2396);
nand U2789 (N_2789,N_2318,N_2328);
nand U2790 (N_2790,N_2365,N_2078);
nand U2791 (N_2791,N_2453,N_2362);
xor U2792 (N_2792,N_2417,N_2415);
nand U2793 (N_2793,N_2030,N_2154);
and U2794 (N_2794,N_2341,N_2333);
nand U2795 (N_2795,N_2217,N_2495);
and U2796 (N_2796,N_2261,N_2016);
and U2797 (N_2797,N_2473,N_2171);
nand U2798 (N_2798,N_2409,N_2101);
or U2799 (N_2799,N_2186,N_2318);
nand U2800 (N_2800,N_2350,N_2192);
and U2801 (N_2801,N_2255,N_2073);
nor U2802 (N_2802,N_2015,N_2270);
and U2803 (N_2803,N_2111,N_2394);
and U2804 (N_2804,N_2100,N_2214);
or U2805 (N_2805,N_2232,N_2463);
xnor U2806 (N_2806,N_2327,N_2361);
nand U2807 (N_2807,N_2216,N_2294);
or U2808 (N_2808,N_2171,N_2131);
and U2809 (N_2809,N_2129,N_2066);
and U2810 (N_2810,N_2476,N_2140);
nor U2811 (N_2811,N_2408,N_2261);
and U2812 (N_2812,N_2212,N_2008);
nand U2813 (N_2813,N_2308,N_2456);
nand U2814 (N_2814,N_2167,N_2378);
or U2815 (N_2815,N_2263,N_2383);
nor U2816 (N_2816,N_2343,N_2337);
nor U2817 (N_2817,N_2130,N_2008);
nand U2818 (N_2818,N_2110,N_2464);
or U2819 (N_2819,N_2023,N_2435);
or U2820 (N_2820,N_2416,N_2215);
nand U2821 (N_2821,N_2143,N_2480);
or U2822 (N_2822,N_2466,N_2216);
and U2823 (N_2823,N_2490,N_2136);
or U2824 (N_2824,N_2006,N_2001);
nand U2825 (N_2825,N_2036,N_2429);
nor U2826 (N_2826,N_2023,N_2455);
nor U2827 (N_2827,N_2369,N_2090);
nand U2828 (N_2828,N_2356,N_2411);
nand U2829 (N_2829,N_2150,N_2199);
nand U2830 (N_2830,N_2189,N_2040);
nor U2831 (N_2831,N_2449,N_2119);
and U2832 (N_2832,N_2346,N_2306);
and U2833 (N_2833,N_2116,N_2092);
or U2834 (N_2834,N_2368,N_2046);
and U2835 (N_2835,N_2473,N_2132);
nand U2836 (N_2836,N_2046,N_2346);
or U2837 (N_2837,N_2284,N_2293);
nor U2838 (N_2838,N_2008,N_2348);
and U2839 (N_2839,N_2030,N_2219);
or U2840 (N_2840,N_2073,N_2333);
or U2841 (N_2841,N_2466,N_2317);
or U2842 (N_2842,N_2055,N_2010);
or U2843 (N_2843,N_2059,N_2451);
nand U2844 (N_2844,N_2428,N_2373);
nor U2845 (N_2845,N_2214,N_2135);
nor U2846 (N_2846,N_2266,N_2084);
and U2847 (N_2847,N_2427,N_2353);
and U2848 (N_2848,N_2088,N_2338);
nor U2849 (N_2849,N_2046,N_2369);
and U2850 (N_2850,N_2138,N_2468);
nand U2851 (N_2851,N_2053,N_2131);
nand U2852 (N_2852,N_2153,N_2259);
or U2853 (N_2853,N_2170,N_2032);
or U2854 (N_2854,N_2340,N_2063);
xor U2855 (N_2855,N_2319,N_2298);
or U2856 (N_2856,N_2411,N_2458);
and U2857 (N_2857,N_2004,N_2063);
nand U2858 (N_2858,N_2324,N_2109);
xnor U2859 (N_2859,N_2177,N_2383);
or U2860 (N_2860,N_2359,N_2035);
or U2861 (N_2861,N_2460,N_2051);
nor U2862 (N_2862,N_2087,N_2105);
xor U2863 (N_2863,N_2279,N_2351);
xor U2864 (N_2864,N_2047,N_2020);
and U2865 (N_2865,N_2032,N_2435);
and U2866 (N_2866,N_2248,N_2198);
or U2867 (N_2867,N_2190,N_2022);
and U2868 (N_2868,N_2138,N_2156);
and U2869 (N_2869,N_2009,N_2225);
or U2870 (N_2870,N_2449,N_2222);
nor U2871 (N_2871,N_2267,N_2392);
or U2872 (N_2872,N_2187,N_2020);
nand U2873 (N_2873,N_2105,N_2452);
nand U2874 (N_2874,N_2387,N_2162);
nor U2875 (N_2875,N_2319,N_2481);
nand U2876 (N_2876,N_2079,N_2118);
nor U2877 (N_2877,N_2102,N_2036);
xor U2878 (N_2878,N_2409,N_2395);
nor U2879 (N_2879,N_2386,N_2399);
and U2880 (N_2880,N_2208,N_2082);
nand U2881 (N_2881,N_2016,N_2087);
nor U2882 (N_2882,N_2304,N_2392);
or U2883 (N_2883,N_2372,N_2323);
or U2884 (N_2884,N_2161,N_2271);
nor U2885 (N_2885,N_2365,N_2490);
or U2886 (N_2886,N_2304,N_2183);
nor U2887 (N_2887,N_2392,N_2294);
and U2888 (N_2888,N_2153,N_2299);
and U2889 (N_2889,N_2125,N_2169);
nor U2890 (N_2890,N_2208,N_2229);
nor U2891 (N_2891,N_2036,N_2237);
nor U2892 (N_2892,N_2261,N_2120);
nand U2893 (N_2893,N_2124,N_2458);
or U2894 (N_2894,N_2329,N_2449);
nor U2895 (N_2895,N_2161,N_2192);
xnor U2896 (N_2896,N_2450,N_2155);
xnor U2897 (N_2897,N_2309,N_2374);
or U2898 (N_2898,N_2085,N_2010);
nor U2899 (N_2899,N_2299,N_2056);
or U2900 (N_2900,N_2259,N_2167);
or U2901 (N_2901,N_2045,N_2086);
nand U2902 (N_2902,N_2441,N_2301);
or U2903 (N_2903,N_2309,N_2088);
xnor U2904 (N_2904,N_2061,N_2174);
nor U2905 (N_2905,N_2324,N_2364);
nand U2906 (N_2906,N_2422,N_2094);
nor U2907 (N_2907,N_2052,N_2078);
or U2908 (N_2908,N_2369,N_2138);
or U2909 (N_2909,N_2441,N_2414);
nor U2910 (N_2910,N_2009,N_2400);
nand U2911 (N_2911,N_2266,N_2161);
nand U2912 (N_2912,N_2312,N_2196);
nand U2913 (N_2913,N_2347,N_2468);
xnor U2914 (N_2914,N_2113,N_2457);
xor U2915 (N_2915,N_2420,N_2236);
and U2916 (N_2916,N_2077,N_2451);
and U2917 (N_2917,N_2046,N_2357);
xor U2918 (N_2918,N_2056,N_2245);
and U2919 (N_2919,N_2409,N_2177);
nand U2920 (N_2920,N_2135,N_2354);
nand U2921 (N_2921,N_2263,N_2228);
or U2922 (N_2922,N_2137,N_2440);
xor U2923 (N_2923,N_2025,N_2203);
nor U2924 (N_2924,N_2053,N_2324);
and U2925 (N_2925,N_2383,N_2123);
or U2926 (N_2926,N_2049,N_2237);
nor U2927 (N_2927,N_2451,N_2415);
nor U2928 (N_2928,N_2491,N_2186);
xnor U2929 (N_2929,N_2011,N_2290);
nand U2930 (N_2930,N_2211,N_2081);
nor U2931 (N_2931,N_2314,N_2273);
nor U2932 (N_2932,N_2434,N_2183);
nand U2933 (N_2933,N_2346,N_2451);
and U2934 (N_2934,N_2125,N_2131);
or U2935 (N_2935,N_2126,N_2116);
nand U2936 (N_2936,N_2363,N_2195);
and U2937 (N_2937,N_2110,N_2458);
nor U2938 (N_2938,N_2266,N_2345);
or U2939 (N_2939,N_2022,N_2402);
or U2940 (N_2940,N_2218,N_2397);
nand U2941 (N_2941,N_2006,N_2004);
and U2942 (N_2942,N_2365,N_2052);
nand U2943 (N_2943,N_2373,N_2425);
nand U2944 (N_2944,N_2309,N_2297);
and U2945 (N_2945,N_2133,N_2418);
xnor U2946 (N_2946,N_2234,N_2353);
and U2947 (N_2947,N_2408,N_2195);
nand U2948 (N_2948,N_2275,N_2395);
or U2949 (N_2949,N_2027,N_2237);
and U2950 (N_2950,N_2197,N_2018);
nor U2951 (N_2951,N_2023,N_2244);
and U2952 (N_2952,N_2487,N_2116);
nor U2953 (N_2953,N_2301,N_2135);
nor U2954 (N_2954,N_2171,N_2187);
or U2955 (N_2955,N_2392,N_2434);
xor U2956 (N_2956,N_2271,N_2445);
and U2957 (N_2957,N_2418,N_2027);
nor U2958 (N_2958,N_2019,N_2080);
nand U2959 (N_2959,N_2182,N_2235);
nor U2960 (N_2960,N_2341,N_2080);
or U2961 (N_2961,N_2002,N_2415);
or U2962 (N_2962,N_2416,N_2457);
or U2963 (N_2963,N_2370,N_2034);
xor U2964 (N_2964,N_2087,N_2052);
nor U2965 (N_2965,N_2094,N_2389);
or U2966 (N_2966,N_2497,N_2017);
and U2967 (N_2967,N_2054,N_2097);
or U2968 (N_2968,N_2307,N_2088);
xor U2969 (N_2969,N_2405,N_2087);
and U2970 (N_2970,N_2164,N_2263);
nand U2971 (N_2971,N_2317,N_2338);
nor U2972 (N_2972,N_2215,N_2456);
nor U2973 (N_2973,N_2224,N_2299);
nor U2974 (N_2974,N_2256,N_2361);
nand U2975 (N_2975,N_2417,N_2308);
and U2976 (N_2976,N_2359,N_2050);
or U2977 (N_2977,N_2064,N_2247);
and U2978 (N_2978,N_2472,N_2047);
and U2979 (N_2979,N_2008,N_2264);
nor U2980 (N_2980,N_2490,N_2125);
and U2981 (N_2981,N_2044,N_2190);
nand U2982 (N_2982,N_2028,N_2252);
nand U2983 (N_2983,N_2217,N_2292);
nor U2984 (N_2984,N_2400,N_2389);
and U2985 (N_2985,N_2327,N_2276);
xnor U2986 (N_2986,N_2175,N_2350);
nand U2987 (N_2987,N_2296,N_2154);
nand U2988 (N_2988,N_2348,N_2368);
and U2989 (N_2989,N_2243,N_2372);
and U2990 (N_2990,N_2439,N_2442);
xnor U2991 (N_2991,N_2049,N_2287);
xor U2992 (N_2992,N_2329,N_2070);
and U2993 (N_2993,N_2327,N_2062);
nor U2994 (N_2994,N_2311,N_2056);
nand U2995 (N_2995,N_2074,N_2039);
nand U2996 (N_2996,N_2366,N_2071);
nor U2997 (N_2997,N_2282,N_2345);
nand U2998 (N_2998,N_2009,N_2499);
nor U2999 (N_2999,N_2004,N_2139);
or UO_0 (O_0,N_2526,N_2673);
or UO_1 (O_1,N_2508,N_2986);
nor UO_2 (O_2,N_2612,N_2515);
or UO_3 (O_3,N_2662,N_2513);
or UO_4 (O_4,N_2649,N_2582);
or UO_5 (O_5,N_2829,N_2545);
xor UO_6 (O_6,N_2932,N_2831);
nor UO_7 (O_7,N_2512,N_2753);
xnor UO_8 (O_8,N_2683,N_2953);
and UO_9 (O_9,N_2656,N_2905);
and UO_10 (O_10,N_2856,N_2989);
nor UO_11 (O_11,N_2786,N_2821);
nor UO_12 (O_12,N_2762,N_2985);
or UO_13 (O_13,N_2535,N_2590);
or UO_14 (O_14,N_2594,N_2852);
and UO_15 (O_15,N_2653,N_2850);
xnor UO_16 (O_16,N_2972,N_2922);
and UO_17 (O_17,N_2849,N_2933);
and UO_18 (O_18,N_2685,N_2613);
nor UO_19 (O_19,N_2518,N_2614);
or UO_20 (O_20,N_2659,N_2519);
nor UO_21 (O_21,N_2992,N_2584);
nand UO_22 (O_22,N_2628,N_2763);
and UO_23 (O_23,N_2892,N_2714);
nor UO_24 (O_24,N_2709,N_2550);
or UO_25 (O_25,N_2864,N_2899);
nand UO_26 (O_26,N_2689,N_2845);
nand UO_27 (O_27,N_2925,N_2681);
or UO_28 (O_28,N_2926,N_2570);
and UO_29 (O_29,N_2901,N_2765);
and UO_30 (O_30,N_2643,N_2872);
or UO_31 (O_31,N_2720,N_2959);
and UO_32 (O_32,N_2573,N_2732);
nand UO_33 (O_33,N_2760,N_2835);
xnor UO_34 (O_34,N_2622,N_2780);
or UO_35 (O_35,N_2994,N_2517);
and UO_36 (O_36,N_2587,N_2878);
nand UO_37 (O_37,N_2657,N_2525);
or UO_38 (O_38,N_2826,N_2772);
or UO_39 (O_39,N_2722,N_2546);
nand UO_40 (O_40,N_2956,N_2748);
nor UO_41 (O_41,N_2975,N_2798);
or UO_42 (O_42,N_2589,N_2710);
or UO_43 (O_43,N_2946,N_2877);
nand UO_44 (O_44,N_2883,N_2941);
xnor UO_45 (O_45,N_2961,N_2898);
or UO_46 (O_46,N_2869,N_2815);
or UO_47 (O_47,N_2991,N_2900);
xor UO_48 (O_48,N_2810,N_2547);
nor UO_49 (O_49,N_2910,N_2749);
nor UO_50 (O_50,N_2718,N_2970);
nor UO_51 (O_51,N_2644,N_2897);
and UO_52 (O_52,N_2706,N_2504);
nand UO_53 (O_53,N_2781,N_2995);
nor UO_54 (O_54,N_2527,N_2880);
nand UO_55 (O_55,N_2971,N_2670);
nand UO_56 (O_56,N_2853,N_2549);
xnor UO_57 (O_57,N_2832,N_2741);
or UO_58 (O_58,N_2819,N_2603);
or UO_59 (O_59,N_2500,N_2928);
or UO_60 (O_60,N_2875,N_2640);
nor UO_61 (O_61,N_2945,N_2949);
and UO_62 (O_62,N_2574,N_2564);
nand UO_63 (O_63,N_2632,N_2509);
or UO_64 (O_64,N_2827,N_2935);
nand UO_65 (O_65,N_2936,N_2805);
nand UO_66 (O_66,N_2777,N_2522);
nor UO_67 (O_67,N_2750,N_2598);
and UO_68 (O_68,N_2544,N_2555);
and UO_69 (O_69,N_2881,N_2999);
nand UO_70 (O_70,N_2811,N_2967);
nand UO_71 (O_71,N_2822,N_2693);
nand UO_72 (O_72,N_2551,N_2755);
nand UO_73 (O_73,N_2723,N_2968);
nor UO_74 (O_74,N_2704,N_2793);
nand UO_75 (O_75,N_2839,N_2571);
or UO_76 (O_76,N_2752,N_2966);
nor UO_77 (O_77,N_2863,N_2751);
nand UO_78 (O_78,N_2982,N_2888);
xnor UO_79 (O_79,N_2857,N_2828);
nor UO_80 (O_80,N_2539,N_2784);
nand UO_81 (O_81,N_2562,N_2913);
nand UO_82 (O_82,N_2833,N_2609);
and UO_83 (O_83,N_2937,N_2838);
or UO_84 (O_84,N_2648,N_2756);
or UO_85 (O_85,N_2542,N_2813);
nor UO_86 (O_86,N_2785,N_2843);
nor UO_87 (O_87,N_2687,N_2896);
and UO_88 (O_88,N_2927,N_2615);
or UO_89 (O_89,N_2906,N_2511);
nor UO_90 (O_90,N_2879,N_2911);
or UO_91 (O_91,N_2783,N_2507);
nor UO_92 (O_92,N_2668,N_2619);
nor UO_93 (O_93,N_2791,N_2921);
xnor UO_94 (O_94,N_2778,N_2909);
and UO_95 (O_95,N_2894,N_2620);
nor UO_96 (O_96,N_2684,N_2672);
nand UO_97 (O_97,N_2637,N_2682);
and UO_98 (O_98,N_2737,N_2680);
or UO_99 (O_99,N_2596,N_2981);
and UO_100 (O_100,N_2770,N_2830);
nand UO_101 (O_101,N_2954,N_2804);
or UO_102 (O_102,N_2788,N_2583);
or UO_103 (O_103,N_2931,N_2803);
or UO_104 (O_104,N_2908,N_2721);
xnor UO_105 (O_105,N_2758,N_2903);
nand UO_106 (O_106,N_2579,N_2987);
nand UO_107 (O_107,N_2824,N_2635);
and UO_108 (O_108,N_2563,N_2790);
or UO_109 (O_109,N_2825,N_2608);
nand UO_110 (O_110,N_2731,N_2980);
nand UO_111 (O_111,N_2739,N_2536);
or UO_112 (O_112,N_2501,N_2963);
or UO_113 (O_113,N_2585,N_2516);
or UO_114 (O_114,N_2624,N_2934);
or UO_115 (O_115,N_2727,N_2862);
xor UO_116 (O_116,N_2923,N_2520);
nand UO_117 (O_117,N_2743,N_2617);
or UO_118 (O_118,N_2602,N_2746);
and UO_119 (O_119,N_2887,N_2707);
or UO_120 (O_120,N_2865,N_2634);
or UO_121 (O_121,N_2600,N_2918);
nor UO_122 (O_122,N_2974,N_2797);
or UO_123 (O_123,N_2965,N_2642);
nor UO_124 (O_124,N_2920,N_2776);
nor UO_125 (O_125,N_2745,N_2715);
xnor UO_126 (O_126,N_2559,N_2904);
nand UO_127 (O_127,N_2868,N_2983);
and UO_128 (O_128,N_2919,N_2766);
and UO_129 (O_129,N_2876,N_2728);
nor UO_130 (O_130,N_2537,N_2917);
nor UO_131 (O_131,N_2789,N_2979);
nand UO_132 (O_132,N_2686,N_2502);
or UO_133 (O_133,N_2695,N_2747);
nand UO_134 (O_134,N_2625,N_2725);
nor UO_135 (O_135,N_2565,N_2719);
nand UO_136 (O_136,N_2667,N_2675);
or UO_137 (O_137,N_2969,N_2611);
and UO_138 (O_138,N_2769,N_2817);
nand UO_139 (O_139,N_2976,N_2802);
nand UO_140 (O_140,N_2978,N_2627);
nand UO_141 (O_141,N_2767,N_2698);
or UO_142 (O_142,N_2738,N_2740);
nor UO_143 (O_143,N_2834,N_2993);
and UO_144 (O_144,N_2629,N_2990);
nand UO_145 (O_145,N_2604,N_2572);
nand UO_146 (O_146,N_2599,N_2799);
and UO_147 (O_147,N_2794,N_2807);
nand UO_148 (O_148,N_2616,N_2757);
nor UO_149 (O_149,N_2534,N_2957);
nor UO_150 (O_150,N_2854,N_2962);
and UO_151 (O_151,N_2702,N_2703);
nand UO_152 (O_152,N_2669,N_2960);
nor UO_153 (O_153,N_2568,N_2840);
and UO_154 (O_154,N_2688,N_2601);
and UO_155 (O_155,N_2855,N_2950);
nand UO_156 (O_156,N_2581,N_2801);
nor UO_157 (O_157,N_2633,N_2606);
nand UO_158 (O_158,N_2610,N_2891);
nand UO_159 (O_159,N_2697,N_2650);
nand UO_160 (O_160,N_2779,N_2692);
nand UO_161 (O_161,N_2848,N_2889);
nor UO_162 (O_162,N_2605,N_2543);
xor UO_163 (O_163,N_2859,N_2973);
nor UO_164 (O_164,N_2506,N_2586);
nor UO_165 (O_165,N_2618,N_2711);
or UO_166 (O_166,N_2996,N_2890);
nand UO_167 (O_167,N_2955,N_2576);
or UO_168 (O_168,N_2561,N_2665);
and UO_169 (O_169,N_2787,N_2958);
nand UO_170 (O_170,N_2663,N_2735);
nor UO_171 (O_171,N_2503,N_2597);
and UO_172 (O_172,N_2567,N_2858);
and UO_173 (O_173,N_2588,N_2851);
or UO_174 (O_174,N_2691,N_2699);
nand UO_175 (O_175,N_2924,N_2800);
or UO_176 (O_176,N_2676,N_2532);
xnor UO_177 (O_177,N_2912,N_2929);
nor UO_178 (O_178,N_2837,N_2951);
or UO_179 (O_179,N_2523,N_2893);
nand UO_180 (O_180,N_2948,N_2874);
nand UO_181 (O_181,N_2771,N_2623);
nor UO_182 (O_182,N_2882,N_2631);
or UO_183 (O_183,N_2754,N_2884);
and UO_184 (O_184,N_2595,N_2538);
nand UO_185 (O_185,N_2809,N_2942);
and UO_186 (O_186,N_2846,N_2541);
and UO_187 (O_187,N_2867,N_2655);
nor UO_188 (O_188,N_2907,N_2510);
nor UO_189 (O_189,N_2836,N_2694);
or UO_190 (O_190,N_2774,N_2964);
xor UO_191 (O_191,N_2870,N_2666);
nand UO_192 (O_192,N_2998,N_2895);
or UO_193 (O_193,N_2560,N_2700);
xnor UO_194 (O_194,N_2873,N_2806);
nor UO_195 (O_195,N_2690,N_2742);
nand UO_196 (O_196,N_2915,N_2708);
nand UO_197 (O_197,N_2592,N_2651);
and UO_198 (O_198,N_2871,N_2768);
and UO_199 (O_199,N_2569,N_2736);
and UO_200 (O_200,N_2729,N_2658);
nand UO_201 (O_201,N_2553,N_2591);
and UO_202 (O_202,N_2943,N_2820);
xnor UO_203 (O_203,N_2795,N_2626);
and UO_204 (O_204,N_2930,N_2885);
nor UO_205 (O_205,N_2952,N_2944);
nand UO_206 (O_206,N_2947,N_2664);
nand UO_207 (O_207,N_2733,N_2808);
and UO_208 (O_208,N_2938,N_2679);
or UO_209 (O_209,N_2764,N_2621);
or UO_210 (O_210,N_2671,N_2902);
nor UO_211 (O_211,N_2726,N_2782);
nand UO_212 (O_212,N_2548,N_2652);
xor UO_213 (O_213,N_2540,N_2775);
and UO_214 (O_214,N_2812,N_2713);
and UO_215 (O_215,N_2984,N_2524);
nor UO_216 (O_216,N_2531,N_2639);
xnor UO_217 (O_217,N_2557,N_2734);
and UO_218 (O_218,N_2844,N_2660);
xor UO_219 (O_219,N_2696,N_2552);
or UO_220 (O_220,N_2886,N_2940);
nor UO_221 (O_221,N_2578,N_2717);
and UO_222 (O_222,N_2505,N_2654);
nor UO_223 (O_223,N_2533,N_2712);
nor UO_224 (O_224,N_2554,N_2530);
nand UO_225 (O_225,N_2792,N_2641);
or UO_226 (O_226,N_2914,N_2773);
nand UO_227 (O_227,N_2916,N_2638);
nand UO_228 (O_228,N_2796,N_2842);
nand UO_229 (O_229,N_2577,N_2705);
xnor UO_230 (O_230,N_2939,N_2730);
nor UO_231 (O_231,N_2645,N_2716);
nand UO_232 (O_232,N_2761,N_2636);
xor UO_233 (O_233,N_2661,N_2529);
xnor UO_234 (O_234,N_2674,N_2575);
and UO_235 (O_235,N_2566,N_2866);
xor UO_236 (O_236,N_2630,N_2823);
xor UO_237 (O_237,N_2847,N_2997);
nand UO_238 (O_238,N_2814,N_2818);
nor UO_239 (O_239,N_2860,N_2607);
nand UO_240 (O_240,N_2724,N_2580);
or UO_241 (O_241,N_2593,N_2744);
nor UO_242 (O_242,N_2677,N_2816);
or UO_243 (O_243,N_2514,N_2558);
nand UO_244 (O_244,N_2759,N_2528);
or UO_245 (O_245,N_2977,N_2988);
nand UO_246 (O_246,N_2841,N_2521);
xor UO_247 (O_247,N_2647,N_2646);
or UO_248 (O_248,N_2678,N_2861);
or UO_249 (O_249,N_2556,N_2701);
nand UO_250 (O_250,N_2610,N_2511);
nand UO_251 (O_251,N_2528,N_2511);
nor UO_252 (O_252,N_2750,N_2636);
and UO_253 (O_253,N_2976,N_2957);
nor UO_254 (O_254,N_2891,N_2911);
nor UO_255 (O_255,N_2764,N_2624);
and UO_256 (O_256,N_2681,N_2505);
nand UO_257 (O_257,N_2942,N_2930);
or UO_258 (O_258,N_2949,N_2606);
nor UO_259 (O_259,N_2596,N_2755);
nand UO_260 (O_260,N_2985,N_2818);
or UO_261 (O_261,N_2779,N_2709);
xor UO_262 (O_262,N_2667,N_2947);
and UO_263 (O_263,N_2788,N_2557);
nor UO_264 (O_264,N_2545,N_2849);
or UO_265 (O_265,N_2884,N_2671);
nor UO_266 (O_266,N_2729,N_2524);
and UO_267 (O_267,N_2854,N_2500);
nand UO_268 (O_268,N_2601,N_2876);
nor UO_269 (O_269,N_2872,N_2740);
or UO_270 (O_270,N_2780,N_2755);
nand UO_271 (O_271,N_2831,N_2649);
and UO_272 (O_272,N_2910,N_2538);
and UO_273 (O_273,N_2869,N_2739);
nor UO_274 (O_274,N_2542,N_2652);
nand UO_275 (O_275,N_2997,N_2844);
nor UO_276 (O_276,N_2502,N_2716);
nor UO_277 (O_277,N_2710,N_2533);
or UO_278 (O_278,N_2930,N_2812);
nor UO_279 (O_279,N_2584,N_2510);
nor UO_280 (O_280,N_2671,N_2966);
nor UO_281 (O_281,N_2896,N_2742);
nand UO_282 (O_282,N_2670,N_2587);
nor UO_283 (O_283,N_2796,N_2826);
nand UO_284 (O_284,N_2530,N_2865);
and UO_285 (O_285,N_2754,N_2578);
nand UO_286 (O_286,N_2793,N_2650);
and UO_287 (O_287,N_2504,N_2777);
nand UO_288 (O_288,N_2615,N_2503);
and UO_289 (O_289,N_2795,N_2972);
nor UO_290 (O_290,N_2919,N_2999);
nor UO_291 (O_291,N_2692,N_2897);
nor UO_292 (O_292,N_2627,N_2678);
and UO_293 (O_293,N_2737,N_2801);
and UO_294 (O_294,N_2728,N_2935);
xor UO_295 (O_295,N_2733,N_2876);
nor UO_296 (O_296,N_2807,N_2983);
nand UO_297 (O_297,N_2777,N_2658);
or UO_298 (O_298,N_2786,N_2802);
and UO_299 (O_299,N_2617,N_2803);
xor UO_300 (O_300,N_2988,N_2876);
nand UO_301 (O_301,N_2721,N_2796);
nand UO_302 (O_302,N_2794,N_2957);
and UO_303 (O_303,N_2613,N_2973);
nor UO_304 (O_304,N_2832,N_2564);
or UO_305 (O_305,N_2835,N_2671);
nand UO_306 (O_306,N_2862,N_2582);
xor UO_307 (O_307,N_2644,N_2795);
and UO_308 (O_308,N_2855,N_2649);
and UO_309 (O_309,N_2774,N_2944);
and UO_310 (O_310,N_2628,N_2589);
or UO_311 (O_311,N_2719,N_2917);
or UO_312 (O_312,N_2850,N_2888);
nand UO_313 (O_313,N_2794,N_2970);
nand UO_314 (O_314,N_2783,N_2564);
xor UO_315 (O_315,N_2892,N_2975);
and UO_316 (O_316,N_2916,N_2644);
nor UO_317 (O_317,N_2973,N_2756);
and UO_318 (O_318,N_2962,N_2630);
and UO_319 (O_319,N_2618,N_2735);
nor UO_320 (O_320,N_2891,N_2558);
nor UO_321 (O_321,N_2592,N_2572);
nor UO_322 (O_322,N_2797,N_2549);
or UO_323 (O_323,N_2570,N_2634);
and UO_324 (O_324,N_2996,N_2885);
nor UO_325 (O_325,N_2946,N_2977);
nor UO_326 (O_326,N_2646,N_2684);
and UO_327 (O_327,N_2937,N_2519);
or UO_328 (O_328,N_2635,N_2650);
or UO_329 (O_329,N_2540,N_2666);
or UO_330 (O_330,N_2921,N_2799);
nor UO_331 (O_331,N_2622,N_2857);
nor UO_332 (O_332,N_2861,N_2661);
or UO_333 (O_333,N_2689,N_2559);
nand UO_334 (O_334,N_2602,N_2950);
and UO_335 (O_335,N_2642,N_2629);
nand UO_336 (O_336,N_2696,N_2712);
nand UO_337 (O_337,N_2915,N_2888);
nand UO_338 (O_338,N_2583,N_2530);
nand UO_339 (O_339,N_2795,N_2549);
or UO_340 (O_340,N_2853,N_2723);
nand UO_341 (O_341,N_2934,N_2594);
xnor UO_342 (O_342,N_2925,N_2764);
and UO_343 (O_343,N_2892,N_2998);
and UO_344 (O_344,N_2809,N_2574);
nand UO_345 (O_345,N_2900,N_2515);
and UO_346 (O_346,N_2777,N_2966);
or UO_347 (O_347,N_2617,N_2579);
nor UO_348 (O_348,N_2842,N_2783);
nor UO_349 (O_349,N_2685,N_2853);
or UO_350 (O_350,N_2990,N_2979);
xor UO_351 (O_351,N_2788,N_2732);
nand UO_352 (O_352,N_2682,N_2904);
nor UO_353 (O_353,N_2752,N_2880);
nand UO_354 (O_354,N_2691,N_2767);
xor UO_355 (O_355,N_2864,N_2941);
nand UO_356 (O_356,N_2644,N_2692);
or UO_357 (O_357,N_2507,N_2822);
nor UO_358 (O_358,N_2522,N_2832);
nand UO_359 (O_359,N_2819,N_2977);
or UO_360 (O_360,N_2581,N_2714);
nor UO_361 (O_361,N_2873,N_2733);
nand UO_362 (O_362,N_2776,N_2834);
or UO_363 (O_363,N_2628,N_2700);
nor UO_364 (O_364,N_2874,N_2598);
and UO_365 (O_365,N_2823,N_2613);
xor UO_366 (O_366,N_2539,N_2710);
or UO_367 (O_367,N_2989,N_2950);
nand UO_368 (O_368,N_2838,N_2680);
or UO_369 (O_369,N_2513,N_2755);
or UO_370 (O_370,N_2894,N_2743);
nand UO_371 (O_371,N_2712,N_2711);
nand UO_372 (O_372,N_2661,N_2714);
and UO_373 (O_373,N_2752,N_2794);
nor UO_374 (O_374,N_2657,N_2580);
xor UO_375 (O_375,N_2630,N_2606);
or UO_376 (O_376,N_2783,N_2824);
or UO_377 (O_377,N_2531,N_2723);
and UO_378 (O_378,N_2629,N_2624);
and UO_379 (O_379,N_2965,N_2808);
or UO_380 (O_380,N_2516,N_2695);
or UO_381 (O_381,N_2725,N_2700);
nor UO_382 (O_382,N_2662,N_2553);
and UO_383 (O_383,N_2895,N_2595);
or UO_384 (O_384,N_2707,N_2540);
nand UO_385 (O_385,N_2813,N_2957);
xor UO_386 (O_386,N_2930,N_2515);
or UO_387 (O_387,N_2524,N_2505);
and UO_388 (O_388,N_2653,N_2828);
xnor UO_389 (O_389,N_2976,N_2789);
nand UO_390 (O_390,N_2774,N_2928);
nor UO_391 (O_391,N_2981,N_2985);
nor UO_392 (O_392,N_2552,N_2834);
nand UO_393 (O_393,N_2787,N_2967);
xnor UO_394 (O_394,N_2516,N_2932);
nand UO_395 (O_395,N_2682,N_2511);
nand UO_396 (O_396,N_2525,N_2771);
and UO_397 (O_397,N_2965,N_2683);
nand UO_398 (O_398,N_2772,N_2830);
or UO_399 (O_399,N_2867,N_2568);
nand UO_400 (O_400,N_2641,N_2663);
and UO_401 (O_401,N_2586,N_2727);
or UO_402 (O_402,N_2946,N_2862);
nand UO_403 (O_403,N_2717,N_2896);
nor UO_404 (O_404,N_2950,N_2780);
or UO_405 (O_405,N_2920,N_2902);
and UO_406 (O_406,N_2920,N_2879);
nand UO_407 (O_407,N_2924,N_2710);
and UO_408 (O_408,N_2891,N_2861);
nor UO_409 (O_409,N_2527,N_2687);
and UO_410 (O_410,N_2760,N_2836);
nor UO_411 (O_411,N_2772,N_2885);
or UO_412 (O_412,N_2696,N_2791);
and UO_413 (O_413,N_2936,N_2953);
nand UO_414 (O_414,N_2916,N_2890);
and UO_415 (O_415,N_2943,N_2958);
and UO_416 (O_416,N_2777,N_2543);
nand UO_417 (O_417,N_2951,N_2587);
nor UO_418 (O_418,N_2618,N_2667);
nand UO_419 (O_419,N_2806,N_2547);
or UO_420 (O_420,N_2752,N_2643);
nor UO_421 (O_421,N_2824,N_2893);
or UO_422 (O_422,N_2693,N_2679);
nor UO_423 (O_423,N_2556,N_2650);
or UO_424 (O_424,N_2574,N_2956);
nor UO_425 (O_425,N_2965,N_2543);
and UO_426 (O_426,N_2782,N_2507);
and UO_427 (O_427,N_2806,N_2697);
nor UO_428 (O_428,N_2599,N_2801);
nor UO_429 (O_429,N_2610,N_2508);
nand UO_430 (O_430,N_2839,N_2776);
nand UO_431 (O_431,N_2899,N_2815);
nand UO_432 (O_432,N_2938,N_2681);
nand UO_433 (O_433,N_2602,N_2774);
and UO_434 (O_434,N_2577,N_2930);
nand UO_435 (O_435,N_2797,N_2708);
nand UO_436 (O_436,N_2756,N_2932);
xnor UO_437 (O_437,N_2966,N_2774);
nor UO_438 (O_438,N_2973,N_2622);
nand UO_439 (O_439,N_2899,N_2992);
or UO_440 (O_440,N_2742,N_2658);
or UO_441 (O_441,N_2977,N_2901);
and UO_442 (O_442,N_2826,N_2730);
and UO_443 (O_443,N_2777,N_2598);
and UO_444 (O_444,N_2776,N_2644);
or UO_445 (O_445,N_2876,N_2873);
nor UO_446 (O_446,N_2759,N_2722);
nor UO_447 (O_447,N_2805,N_2884);
or UO_448 (O_448,N_2863,N_2694);
nor UO_449 (O_449,N_2950,N_2841);
or UO_450 (O_450,N_2651,N_2952);
and UO_451 (O_451,N_2762,N_2608);
nor UO_452 (O_452,N_2592,N_2537);
nand UO_453 (O_453,N_2513,N_2748);
nand UO_454 (O_454,N_2873,N_2839);
and UO_455 (O_455,N_2601,N_2672);
and UO_456 (O_456,N_2740,N_2976);
or UO_457 (O_457,N_2717,N_2835);
nor UO_458 (O_458,N_2892,N_2699);
or UO_459 (O_459,N_2530,N_2682);
or UO_460 (O_460,N_2711,N_2944);
or UO_461 (O_461,N_2638,N_2704);
xor UO_462 (O_462,N_2720,N_2529);
or UO_463 (O_463,N_2915,N_2599);
nand UO_464 (O_464,N_2541,N_2947);
and UO_465 (O_465,N_2580,N_2569);
nand UO_466 (O_466,N_2797,N_2618);
xnor UO_467 (O_467,N_2836,N_2565);
nand UO_468 (O_468,N_2775,N_2649);
or UO_469 (O_469,N_2766,N_2770);
nand UO_470 (O_470,N_2614,N_2757);
nand UO_471 (O_471,N_2989,N_2613);
and UO_472 (O_472,N_2625,N_2992);
nor UO_473 (O_473,N_2949,N_2615);
and UO_474 (O_474,N_2861,N_2583);
or UO_475 (O_475,N_2710,N_2978);
and UO_476 (O_476,N_2900,N_2721);
or UO_477 (O_477,N_2605,N_2601);
nor UO_478 (O_478,N_2862,N_2803);
and UO_479 (O_479,N_2637,N_2791);
nor UO_480 (O_480,N_2738,N_2945);
and UO_481 (O_481,N_2605,N_2945);
nor UO_482 (O_482,N_2711,N_2511);
and UO_483 (O_483,N_2813,N_2839);
nor UO_484 (O_484,N_2735,N_2613);
nor UO_485 (O_485,N_2504,N_2918);
or UO_486 (O_486,N_2734,N_2890);
or UO_487 (O_487,N_2505,N_2619);
nor UO_488 (O_488,N_2752,N_2757);
nand UO_489 (O_489,N_2640,N_2849);
nand UO_490 (O_490,N_2664,N_2574);
xnor UO_491 (O_491,N_2780,N_2783);
or UO_492 (O_492,N_2898,N_2691);
and UO_493 (O_493,N_2794,N_2871);
xor UO_494 (O_494,N_2611,N_2868);
and UO_495 (O_495,N_2694,N_2794);
or UO_496 (O_496,N_2995,N_2645);
nand UO_497 (O_497,N_2517,N_2814);
nand UO_498 (O_498,N_2825,N_2619);
nor UO_499 (O_499,N_2752,N_2888);
endmodule