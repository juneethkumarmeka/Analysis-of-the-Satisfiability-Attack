module basic_1000_10000_1500_4_levels_2xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_646,In_695);
nand U1 (N_1,In_318,In_937);
or U2 (N_2,In_362,In_792);
or U3 (N_3,In_209,In_854);
nand U4 (N_4,In_418,In_847);
nand U5 (N_5,In_867,In_578);
and U6 (N_6,In_402,In_324);
xnor U7 (N_7,In_316,In_896);
and U8 (N_8,In_672,In_832);
nor U9 (N_9,In_950,In_165);
or U10 (N_10,In_149,In_132);
nand U11 (N_11,In_167,In_448);
or U12 (N_12,In_178,In_888);
or U13 (N_13,In_617,In_211);
nand U14 (N_14,In_295,In_258);
nor U15 (N_15,In_637,In_986);
nand U16 (N_16,In_887,In_882);
nand U17 (N_17,In_341,In_837);
or U18 (N_18,In_797,In_838);
and U19 (N_19,In_640,In_535);
and U20 (N_20,In_962,In_726);
nor U21 (N_21,In_493,In_667);
and U22 (N_22,In_115,In_243);
or U23 (N_23,In_782,In_984);
nand U24 (N_24,In_154,In_928);
and U25 (N_25,In_199,In_465);
nand U26 (N_26,In_90,In_459);
nand U27 (N_27,In_260,In_565);
or U28 (N_28,In_456,In_284);
or U29 (N_29,In_57,In_377);
nand U30 (N_30,In_993,In_959);
nor U31 (N_31,In_319,In_985);
and U32 (N_32,In_357,In_277);
nor U33 (N_33,In_879,In_643);
and U34 (N_34,In_813,In_666);
or U35 (N_35,In_8,In_970);
nand U36 (N_36,In_487,In_796);
xor U37 (N_37,In_486,In_768);
nor U38 (N_38,In_698,In_711);
and U39 (N_39,In_831,In_185);
nor U40 (N_40,In_676,In_148);
nand U41 (N_41,In_670,In_688);
and U42 (N_42,In_50,In_771);
and U43 (N_43,In_411,In_5);
nor U44 (N_44,In_395,In_923);
nor U45 (N_45,In_592,In_337);
or U46 (N_46,In_735,In_495);
nand U47 (N_47,In_684,In_146);
nand U48 (N_48,In_292,In_889);
xnor U49 (N_49,In_127,In_938);
nand U50 (N_50,In_464,In_124);
or U51 (N_51,In_326,In_363);
nand U52 (N_52,In_836,In_811);
and U53 (N_53,In_91,In_692);
and U54 (N_54,In_399,In_681);
or U55 (N_55,In_259,In_225);
nand U56 (N_56,In_375,In_351);
and U57 (N_57,In_182,In_651);
nor U58 (N_58,In_415,In_496);
or U59 (N_59,In_957,In_77);
nand U60 (N_60,In_435,In_931);
and U61 (N_61,In_95,In_783);
or U62 (N_62,In_886,In_151);
or U63 (N_63,In_475,In_97);
and U64 (N_64,In_300,In_170);
or U65 (N_65,In_786,In_273);
nor U66 (N_66,In_791,In_562);
nand U67 (N_67,In_851,In_787);
nor U68 (N_68,In_530,In_668);
nor U69 (N_69,In_54,In_370);
nor U70 (N_70,In_102,In_850);
nand U71 (N_71,In_502,In_274);
nor U72 (N_72,In_999,In_972);
nor U73 (N_73,In_463,In_618);
and U74 (N_74,In_433,In_848);
and U75 (N_75,In_400,In_874);
nand U76 (N_76,In_864,In_113);
and U77 (N_77,In_757,In_344);
xnor U78 (N_78,In_653,In_358);
nand U79 (N_79,In_752,In_569);
and U80 (N_80,In_65,In_620);
or U81 (N_81,In_247,In_120);
nor U82 (N_82,In_539,In_43);
or U83 (N_83,In_145,In_511);
and U84 (N_84,In_858,In_648);
and U85 (N_85,In_437,In_571);
or U86 (N_86,In_169,In_673);
nand U87 (N_87,In_980,In_829);
nand U88 (N_88,In_86,In_443);
nor U89 (N_89,In_275,In_122);
nor U90 (N_90,In_389,In_899);
or U91 (N_91,In_594,In_195);
or U92 (N_92,In_62,In_770);
or U93 (N_93,In_164,In_656);
nor U94 (N_94,In_215,In_631);
and U95 (N_95,In_731,In_743);
nor U96 (N_96,In_559,In_407);
and U97 (N_97,In_379,In_71);
or U98 (N_98,In_368,In_333);
or U99 (N_99,In_373,In_348);
and U100 (N_100,In_955,In_480);
or U101 (N_101,In_349,In_966);
nand U102 (N_102,In_208,In_834);
nor U103 (N_103,In_466,In_645);
or U104 (N_104,In_366,In_983);
or U105 (N_105,In_23,In_343);
xnor U106 (N_106,In_194,In_59);
nor U107 (N_107,In_642,In_206);
and U108 (N_108,In_558,In_416);
or U109 (N_109,In_100,In_925);
nand U110 (N_110,In_892,In_222);
nor U111 (N_111,In_807,In_736);
nor U112 (N_112,In_941,In_184);
nor U113 (N_113,In_755,In_545);
nand U114 (N_114,In_626,In_34);
nand U115 (N_115,In_803,In_320);
nor U116 (N_116,In_678,In_25);
or U117 (N_117,In_898,In_556);
nor U118 (N_118,In_682,In_239);
or U119 (N_119,In_136,In_897);
nor U120 (N_120,In_18,In_360);
nor U121 (N_121,In_614,In_88);
nand U122 (N_122,In_629,In_778);
or U123 (N_123,In_111,In_805);
nor U124 (N_124,In_779,In_537);
nand U125 (N_125,In_514,In_451);
nand U126 (N_126,In_309,In_623);
nor U127 (N_127,In_622,In_598);
nand U128 (N_128,In_975,In_152);
nor U129 (N_129,In_762,In_795);
and U130 (N_130,In_595,In_74);
nand U131 (N_131,In_80,In_760);
or U132 (N_132,In_608,In_953);
and U133 (N_133,In_905,In_104);
and U134 (N_134,In_526,In_754);
or U135 (N_135,In_491,In_586);
nor U136 (N_136,In_554,In_20);
xnor U137 (N_137,In_956,In_665);
nor U138 (N_138,In_340,In_103);
nor U139 (N_139,In_262,In_912);
nand U140 (N_140,In_193,In_265);
or U141 (N_141,In_188,In_15);
nor U142 (N_142,In_890,In_790);
nand U143 (N_143,In_301,In_60);
and U144 (N_144,In_424,In_374);
and U145 (N_145,In_677,In_991);
and U146 (N_146,In_744,In_290);
and U147 (N_147,In_429,In_609);
or U148 (N_148,In_179,In_244);
and U149 (N_149,In_878,In_106);
nand U150 (N_150,In_426,In_588);
or U151 (N_151,In_24,In_322);
and U152 (N_152,In_764,In_428);
nand U153 (N_153,In_973,In_998);
nand U154 (N_154,In_599,In_442);
nor U155 (N_155,In_506,In_914);
xor U156 (N_156,In_974,In_432);
nor U157 (N_157,In_427,In_128);
and U158 (N_158,In_885,In_249);
and U159 (N_159,In_745,In_781);
nor U160 (N_160,In_553,In_489);
and U161 (N_161,In_187,In_647);
and U162 (N_162,In_474,In_392);
nor U163 (N_163,In_235,In_661);
xor U164 (N_164,In_460,In_384);
nor U165 (N_165,In_982,In_849);
nor U166 (N_166,In_141,In_978);
or U167 (N_167,In_388,In_621);
nor U168 (N_168,In_328,In_131);
and U169 (N_169,In_257,In_561);
nand U170 (N_170,In_439,In_968);
or U171 (N_171,In_61,In_627);
nor U172 (N_172,In_21,In_523);
nand U173 (N_173,In_823,In_250);
nand U174 (N_174,In_761,In_458);
nand U175 (N_175,In_995,In_660);
or U176 (N_176,In_963,In_822);
and U177 (N_177,In_630,In_910);
xnor U178 (N_178,In_632,In_172);
nand U179 (N_179,In_160,In_875);
nand U180 (N_180,In_338,In_902);
or U181 (N_181,In_72,In_943);
nand U182 (N_182,In_446,In_810);
nor U183 (N_183,In_236,In_305);
nor U184 (N_184,In_671,In_650);
or U185 (N_185,In_721,In_53);
or U186 (N_186,In_767,In_430);
nor U187 (N_187,In_306,In_347);
nand U188 (N_188,In_585,In_94);
nor U189 (N_189,In_518,In_470);
nand U190 (N_190,In_177,In_840);
nor U191 (N_191,In_738,In_68);
and U192 (N_192,In_253,In_212);
nor U193 (N_193,In_230,In_143);
and U194 (N_194,In_855,In_175);
nor U195 (N_195,In_278,In_254);
and U196 (N_196,In_500,In_323);
or U197 (N_197,In_525,In_335);
or U198 (N_198,In_334,In_583);
nor U199 (N_199,In_830,In_775);
nor U200 (N_200,In_64,In_107);
nor U201 (N_201,In_935,In_683);
nand U202 (N_202,In_266,In_376);
nand U203 (N_203,In_505,In_288);
or U204 (N_204,In_602,In_971);
nand U205 (N_205,In_593,In_483);
nand U206 (N_206,In_891,In_529);
nand U207 (N_207,In_719,In_503);
or U208 (N_208,In_380,In_741);
nand U209 (N_209,In_546,In_150);
nor U210 (N_210,In_951,In_210);
xor U211 (N_211,In_156,In_297);
and U212 (N_212,In_990,In_996);
and U213 (N_213,In_99,In_261);
or U214 (N_214,In_272,In_397);
or U215 (N_215,In_203,In_12);
nand U216 (N_216,In_733,In_659);
or U217 (N_217,In_478,In_16);
or U218 (N_218,In_447,In_157);
nand U219 (N_219,In_2,In_139);
nor U220 (N_220,In_844,In_516);
nand U221 (N_221,In_66,In_445);
and U222 (N_222,In_624,In_354);
and U223 (N_223,In_385,In_96);
nor U224 (N_224,In_317,In_939);
nand U225 (N_225,In_461,In_469);
nor U226 (N_226,In_521,In_276);
or U227 (N_227,In_784,In_863);
and U228 (N_228,In_965,In_490);
or U229 (N_229,In_229,In_785);
nand U230 (N_230,In_454,In_730);
nor U231 (N_231,In_11,In_158);
nor U232 (N_232,In_381,In_204);
and U233 (N_233,In_36,In_270);
nor U234 (N_234,In_180,In_920);
xnor U235 (N_235,In_872,In_765);
and U236 (N_236,In_406,In_28);
and U237 (N_237,In_135,In_927);
nor U238 (N_238,In_192,In_37);
and U239 (N_239,In_828,In_710);
or U240 (N_240,In_126,In_815);
or U241 (N_241,In_308,In_409);
or U242 (N_242,In_967,In_241);
and U243 (N_243,In_960,In_142);
nor U244 (N_244,In_232,In_843);
and U245 (N_245,In_138,In_689);
and U246 (N_246,In_93,In_255);
nand U247 (N_247,In_728,In_331);
nand U248 (N_248,In_285,In_75);
nor U249 (N_249,In_748,In_568);
nor U250 (N_250,In_436,In_371);
nand U251 (N_251,In_940,In_410);
nand U252 (N_252,In_657,In_528);
and U253 (N_253,In_52,In_664);
and U254 (N_254,In_549,In_234);
nand U255 (N_255,In_669,In_176);
nand U256 (N_256,In_48,In_520);
nor U257 (N_257,In_922,In_981);
and U258 (N_258,In_9,In_13);
or U259 (N_259,In_788,In_361);
nand U260 (N_260,In_299,In_751);
or U261 (N_261,In_870,In_641);
or U262 (N_262,In_507,In_425);
or U263 (N_263,In_693,In_31);
xor U264 (N_264,In_625,In_223);
or U265 (N_265,In_233,In_33);
nand U266 (N_266,In_694,In_871);
and U267 (N_267,In_680,In_396);
and U268 (N_268,In_155,In_27);
nor U269 (N_269,In_312,In_687);
nand U270 (N_270,In_574,In_263);
nor U271 (N_271,In_359,In_110);
or U272 (N_272,In_540,In_703);
and U273 (N_273,In_67,In_383);
nor U274 (N_274,In_824,In_367);
nand U275 (N_275,In_945,In_708);
nand U276 (N_276,In_596,In_378);
or U277 (N_277,In_41,In_699);
or U278 (N_278,In_42,In_504);
and U279 (N_279,In_917,In_512);
and U280 (N_280,In_524,In_189);
or U281 (N_281,In_311,In_325);
or U282 (N_282,In_780,In_551);
and U283 (N_283,In_296,In_531);
and U284 (N_284,In_382,In_936);
nor U285 (N_285,In_964,In_423);
and U286 (N_286,In_774,In_701);
nor U287 (N_287,In_286,In_32);
nand U288 (N_288,In_987,In_513);
or U289 (N_289,In_582,In_841);
or U290 (N_290,In_471,In_499);
and U291 (N_291,In_462,In_481);
nor U292 (N_292,In_268,In_716);
nor U293 (N_293,In_579,In_712);
nand U294 (N_294,In_809,In_605);
nand U295 (N_295,In_720,In_509);
nor U296 (N_296,In_597,In_707);
nand U297 (N_297,In_314,In_183);
nand U298 (N_298,In_421,In_747);
or U299 (N_299,In_759,In_134);
nand U300 (N_300,In_394,In_477);
and U301 (N_301,In_70,In_422);
and U302 (N_302,In_919,In_538);
nor U303 (N_303,In_994,In_918);
nand U304 (N_304,In_536,In_746);
and U305 (N_305,In_825,In_600);
nand U306 (N_306,In_619,In_22);
and U307 (N_307,In_412,In_214);
or U308 (N_308,In_452,In_527);
and U309 (N_309,In_772,In_1);
and U310 (N_310,In_457,In_85);
nor U311 (N_311,In_654,In_369);
or U312 (N_312,In_789,In_390);
nand U313 (N_313,In_4,In_205);
or U314 (N_314,In_353,In_532);
nand U315 (N_315,In_638,In_915);
and U316 (N_316,In_827,In_900);
and U317 (N_317,In_181,In_812);
nor U318 (N_318,In_894,In_329);
nand U319 (N_319,In_954,In_227);
or U320 (N_320,In_794,In_391);
nor U321 (N_321,In_611,In_476);
nor U322 (N_322,In_769,In_417);
nand U323 (N_323,In_799,In_674);
nor U324 (N_324,In_560,In_472);
nand U325 (N_325,In_419,In_880);
xor U326 (N_326,In_649,In_269);
nand U327 (N_327,In_218,In_753);
nor U328 (N_328,In_921,In_550);
and U329 (N_329,In_715,In_35);
xnor U330 (N_330,In_542,In_281);
and U331 (N_331,In_804,In_818);
nor U332 (N_332,In_663,In_352);
or U333 (N_333,In_144,In_814);
or U334 (N_334,In_979,In_201);
nand U335 (N_335,In_750,In_833);
nor U336 (N_336,In_387,In_977);
nor U337 (N_337,In_413,In_846);
nor U338 (N_338,In_207,In_658);
and U339 (N_339,In_817,In_685);
nor U340 (N_340,In_81,In_130);
or U341 (N_341,In_434,In_55);
or U342 (N_342,In_821,In_116);
nor U343 (N_343,In_566,In_372);
nor U344 (N_344,In_853,In_264);
or U345 (N_345,In_294,In_246);
nor U346 (N_346,In_332,In_226);
or U347 (N_347,In_958,In_793);
and U348 (N_348,In_946,In_522);
nor U349 (N_349,In_237,In_570);
or U350 (N_350,In_961,In_901);
nor U351 (N_351,In_635,In_0);
or U352 (N_352,In_404,In_479);
or U353 (N_353,In_129,In_533);
nand U354 (N_354,In_628,In_238);
or U355 (N_355,In_14,In_808);
nand U356 (N_356,In_168,In_904);
or U357 (N_357,In_162,In_510);
and U358 (N_358,In_845,In_916);
nor U359 (N_359,In_860,In_137);
nand U360 (N_360,In_112,In_679);
nand U361 (N_361,In_929,In_355);
nor U362 (N_362,In_603,In_842);
and U363 (N_363,In_153,In_908);
or U364 (N_364,In_909,In_947);
or U365 (N_365,In_310,In_856);
nor U366 (N_366,In_515,In_161);
or U367 (N_367,In_932,In_87);
or U368 (N_368,In_644,In_44);
or U369 (N_369,In_220,In_826);
nor U370 (N_370,In_729,In_756);
and U371 (N_371,In_557,In_484);
xor U372 (N_372,In_576,In_776);
nand U373 (N_373,In_485,In_873);
and U374 (N_374,In_655,In_49);
nand U375 (N_375,In_58,In_287);
or U376 (N_376,In_98,In_604);
or U377 (N_377,In_587,In_488);
and U378 (N_378,In_766,In_444);
nor U379 (N_379,In_39,In_607);
nand U380 (N_380,In_173,In_267);
and U381 (N_381,In_125,In_198);
or U382 (N_382,In_690,In_877);
nand U383 (N_383,In_302,In_816);
or U384 (N_384,In_572,In_298);
and U385 (N_385,In_83,In_934);
or U386 (N_386,In_467,In_200);
nor U387 (N_387,In_453,In_590);
nand U388 (N_388,In_256,In_398);
and U389 (N_389,In_926,In_386);
nor U390 (N_390,In_580,In_541);
or U391 (N_391,In_911,In_327);
nor U392 (N_392,In_19,In_700);
and U393 (N_393,In_903,In_802);
nand U394 (N_394,In_722,In_517);
or U395 (N_395,In_691,In_497);
nand U396 (N_396,In_989,In_171);
or U397 (N_397,In_202,In_108);
and U398 (N_398,In_997,In_543);
and U399 (N_399,In_547,In_866);
nand U400 (N_400,In_252,In_835);
and U401 (N_401,In_73,In_7);
or U402 (N_402,In_573,In_865);
or U403 (N_403,In_702,In_468);
nand U404 (N_404,In_612,In_304);
and U405 (N_405,In_219,In_868);
or U406 (N_406,In_742,In_705);
or U407 (N_407,In_723,In_952);
nor U408 (N_408,In_405,In_408);
or U409 (N_409,In_248,In_633);
nor U410 (N_410,In_924,In_763);
and U411 (N_411,In_589,In_801);
or U412 (N_412,In_534,In_662);
and U413 (N_413,In_186,In_696);
and U414 (N_414,In_555,In_508);
nor U415 (N_415,In_438,In_675);
or U416 (N_416,In_321,In_76);
nor U417 (N_417,In_40,In_345);
and U418 (N_418,In_289,In_51);
and U419 (N_419,In_140,In_652);
or U420 (N_420,In_29,In_820);
xor U421 (N_421,In_197,In_26);
nor U422 (N_422,In_401,In_293);
nor U423 (N_423,In_913,In_330);
and U424 (N_424,In_17,In_519);
nand U425 (N_425,In_431,In_3);
nor U426 (N_426,In_615,In_852);
or U427 (N_427,In_283,In_717);
and U428 (N_428,In_706,In_307);
xnor U429 (N_429,In_591,In_216);
and U430 (N_430,In_450,In_231);
or U431 (N_431,In_869,In_101);
nand U432 (N_432,In_105,In_893);
or U433 (N_433,In_365,In_739);
nand U434 (N_434,In_117,In_713);
or U435 (N_435,In_906,In_191);
or U436 (N_436,In_806,In_933);
or U437 (N_437,In_414,In_686);
or U438 (N_438,In_190,In_271);
and U439 (N_439,In_174,In_240);
or U440 (N_440,In_46,In_196);
nor U441 (N_441,In_291,In_969);
and U442 (N_442,In_133,In_876);
or U443 (N_443,In_494,In_455);
and U444 (N_444,In_988,In_714);
or U445 (N_445,In_734,In_84);
or U446 (N_446,In_709,In_303);
or U447 (N_447,In_861,In_224);
nand U448 (N_448,In_548,In_704);
or U449 (N_449,In_242,In_119);
or U450 (N_450,In_501,In_732);
and U451 (N_451,In_773,In_563);
nor U452 (N_452,In_393,In_616);
and U453 (N_453,In_159,In_949);
nor U454 (N_454,In_123,In_948);
nor U455 (N_455,In_737,In_581);
or U456 (N_456,In_819,In_839);
and U457 (N_457,In_279,In_564);
or U458 (N_458,In_498,In_881);
or U459 (N_459,In_10,In_567);
nand U460 (N_460,In_163,In_610);
nor U461 (N_461,In_47,In_639);
nand U462 (N_462,In_92,In_976);
or U463 (N_463,In_492,In_749);
nor U464 (N_464,In_883,In_441);
or U465 (N_465,In_109,In_575);
nand U466 (N_466,In_56,In_482);
nand U467 (N_467,In_944,In_473);
nand U468 (N_468,In_89,In_217);
and U469 (N_469,In_859,In_166);
or U470 (N_470,In_30,In_552);
nand U471 (N_471,In_634,In_758);
and U472 (N_472,In_356,In_992);
or U473 (N_473,In_544,In_346);
nand U474 (N_474,In_577,In_601);
and U475 (N_475,In_800,In_895);
or U476 (N_476,In_336,In_740);
nand U477 (N_477,In_907,In_147);
xor U478 (N_478,In_727,In_38);
nor U479 (N_479,In_350,In_342);
nand U480 (N_480,In_724,In_725);
or U481 (N_481,In_280,In_6);
nand U482 (N_482,In_584,In_213);
and U483 (N_483,In_697,In_339);
or U484 (N_484,In_121,In_942);
nor U485 (N_485,In_63,In_613);
or U486 (N_486,In_245,In_78);
nor U487 (N_487,In_440,In_606);
nor U488 (N_488,In_420,In_69);
or U489 (N_489,In_228,In_118);
nand U490 (N_490,In_282,In_313);
or U491 (N_491,In_636,In_221);
and U492 (N_492,In_930,In_449);
nand U493 (N_493,In_82,In_364);
or U494 (N_494,In_798,In_718);
or U495 (N_495,In_403,In_315);
nor U496 (N_496,In_114,In_79);
nand U497 (N_497,In_251,In_862);
and U498 (N_498,In_777,In_884);
or U499 (N_499,In_45,In_857);
nor U500 (N_500,In_685,In_159);
nand U501 (N_501,In_584,In_709);
xnor U502 (N_502,In_533,In_669);
or U503 (N_503,In_217,In_495);
nor U504 (N_504,In_308,In_260);
and U505 (N_505,In_216,In_902);
nand U506 (N_506,In_126,In_716);
and U507 (N_507,In_888,In_833);
and U508 (N_508,In_481,In_415);
or U509 (N_509,In_57,In_401);
and U510 (N_510,In_961,In_271);
and U511 (N_511,In_214,In_362);
and U512 (N_512,In_206,In_851);
or U513 (N_513,In_865,In_477);
nor U514 (N_514,In_627,In_120);
xnor U515 (N_515,In_662,In_657);
and U516 (N_516,In_715,In_410);
and U517 (N_517,In_723,In_549);
or U518 (N_518,In_431,In_184);
or U519 (N_519,In_637,In_104);
or U520 (N_520,In_30,In_484);
nand U521 (N_521,In_877,In_83);
nand U522 (N_522,In_35,In_942);
and U523 (N_523,In_266,In_6);
nand U524 (N_524,In_727,In_849);
and U525 (N_525,In_93,In_283);
nor U526 (N_526,In_638,In_213);
nor U527 (N_527,In_621,In_504);
nor U528 (N_528,In_264,In_266);
or U529 (N_529,In_576,In_466);
nor U530 (N_530,In_4,In_114);
and U531 (N_531,In_728,In_777);
and U532 (N_532,In_784,In_662);
nand U533 (N_533,In_472,In_89);
nand U534 (N_534,In_325,In_466);
or U535 (N_535,In_183,In_385);
nand U536 (N_536,In_508,In_424);
xor U537 (N_537,In_25,In_348);
nand U538 (N_538,In_894,In_824);
nand U539 (N_539,In_826,In_723);
nor U540 (N_540,In_433,In_487);
nor U541 (N_541,In_217,In_127);
and U542 (N_542,In_898,In_128);
nand U543 (N_543,In_242,In_54);
nor U544 (N_544,In_728,In_134);
nand U545 (N_545,In_870,In_192);
or U546 (N_546,In_521,In_149);
nor U547 (N_547,In_152,In_154);
nor U548 (N_548,In_747,In_797);
nand U549 (N_549,In_403,In_96);
or U550 (N_550,In_708,In_975);
or U551 (N_551,In_883,In_206);
nor U552 (N_552,In_692,In_389);
nand U553 (N_553,In_811,In_565);
nand U554 (N_554,In_70,In_864);
and U555 (N_555,In_460,In_532);
nor U556 (N_556,In_371,In_46);
nand U557 (N_557,In_501,In_622);
or U558 (N_558,In_912,In_439);
nor U559 (N_559,In_502,In_665);
and U560 (N_560,In_710,In_321);
nand U561 (N_561,In_670,In_859);
and U562 (N_562,In_386,In_73);
xor U563 (N_563,In_767,In_807);
nand U564 (N_564,In_534,In_256);
and U565 (N_565,In_59,In_485);
and U566 (N_566,In_150,In_862);
nor U567 (N_567,In_485,In_393);
nand U568 (N_568,In_117,In_396);
or U569 (N_569,In_240,In_499);
nand U570 (N_570,In_466,In_548);
or U571 (N_571,In_587,In_977);
nand U572 (N_572,In_418,In_338);
and U573 (N_573,In_323,In_719);
or U574 (N_574,In_799,In_964);
or U575 (N_575,In_459,In_986);
and U576 (N_576,In_96,In_985);
or U577 (N_577,In_776,In_507);
nor U578 (N_578,In_462,In_663);
nor U579 (N_579,In_474,In_377);
nand U580 (N_580,In_920,In_980);
nor U581 (N_581,In_421,In_128);
and U582 (N_582,In_978,In_54);
nand U583 (N_583,In_535,In_469);
nor U584 (N_584,In_878,In_771);
or U585 (N_585,In_144,In_89);
or U586 (N_586,In_508,In_453);
nand U587 (N_587,In_957,In_193);
and U588 (N_588,In_871,In_480);
or U589 (N_589,In_570,In_288);
or U590 (N_590,In_191,In_500);
nand U591 (N_591,In_648,In_148);
xor U592 (N_592,In_709,In_477);
nor U593 (N_593,In_571,In_471);
and U594 (N_594,In_87,In_103);
xor U595 (N_595,In_471,In_768);
or U596 (N_596,In_194,In_141);
or U597 (N_597,In_696,In_385);
nor U598 (N_598,In_614,In_744);
and U599 (N_599,In_208,In_911);
or U600 (N_600,In_641,In_386);
xnor U601 (N_601,In_87,In_115);
nor U602 (N_602,In_393,In_443);
nand U603 (N_603,In_930,In_98);
nor U604 (N_604,In_458,In_772);
nor U605 (N_605,In_946,In_400);
nor U606 (N_606,In_414,In_802);
or U607 (N_607,In_340,In_307);
and U608 (N_608,In_777,In_817);
nand U609 (N_609,In_492,In_875);
or U610 (N_610,In_93,In_56);
nand U611 (N_611,In_660,In_834);
xnor U612 (N_612,In_329,In_808);
nand U613 (N_613,In_736,In_841);
nor U614 (N_614,In_902,In_316);
or U615 (N_615,In_511,In_551);
nand U616 (N_616,In_896,In_49);
and U617 (N_617,In_162,In_196);
or U618 (N_618,In_489,In_526);
and U619 (N_619,In_886,In_173);
and U620 (N_620,In_849,In_827);
nand U621 (N_621,In_265,In_156);
and U622 (N_622,In_219,In_651);
nor U623 (N_623,In_492,In_9);
or U624 (N_624,In_314,In_145);
or U625 (N_625,In_187,In_293);
nand U626 (N_626,In_282,In_491);
nor U627 (N_627,In_948,In_497);
and U628 (N_628,In_45,In_637);
nor U629 (N_629,In_356,In_660);
or U630 (N_630,In_674,In_145);
or U631 (N_631,In_194,In_757);
nand U632 (N_632,In_39,In_913);
nor U633 (N_633,In_195,In_985);
and U634 (N_634,In_148,In_663);
and U635 (N_635,In_580,In_121);
and U636 (N_636,In_193,In_628);
nand U637 (N_637,In_777,In_638);
or U638 (N_638,In_337,In_759);
or U639 (N_639,In_75,In_982);
or U640 (N_640,In_201,In_80);
nor U641 (N_641,In_704,In_151);
or U642 (N_642,In_422,In_684);
nand U643 (N_643,In_197,In_500);
nand U644 (N_644,In_317,In_15);
or U645 (N_645,In_271,In_237);
and U646 (N_646,In_163,In_118);
or U647 (N_647,In_463,In_222);
or U648 (N_648,In_113,In_213);
and U649 (N_649,In_2,In_827);
and U650 (N_650,In_104,In_837);
nand U651 (N_651,In_771,In_579);
and U652 (N_652,In_579,In_542);
nand U653 (N_653,In_314,In_229);
or U654 (N_654,In_253,In_313);
nand U655 (N_655,In_133,In_491);
and U656 (N_656,In_667,In_699);
nor U657 (N_657,In_356,In_586);
nand U658 (N_658,In_77,In_622);
and U659 (N_659,In_893,In_14);
and U660 (N_660,In_207,In_790);
or U661 (N_661,In_381,In_574);
nand U662 (N_662,In_712,In_289);
and U663 (N_663,In_590,In_374);
nand U664 (N_664,In_131,In_752);
and U665 (N_665,In_322,In_11);
or U666 (N_666,In_580,In_349);
nand U667 (N_667,In_849,In_170);
xor U668 (N_668,In_40,In_606);
and U669 (N_669,In_408,In_189);
nand U670 (N_670,In_983,In_346);
nand U671 (N_671,In_312,In_72);
xnor U672 (N_672,In_673,In_496);
or U673 (N_673,In_106,In_11);
and U674 (N_674,In_969,In_836);
and U675 (N_675,In_930,In_851);
and U676 (N_676,In_884,In_652);
nor U677 (N_677,In_737,In_638);
nor U678 (N_678,In_142,In_874);
nand U679 (N_679,In_743,In_857);
nand U680 (N_680,In_594,In_659);
nor U681 (N_681,In_961,In_763);
and U682 (N_682,In_372,In_788);
nor U683 (N_683,In_981,In_174);
nand U684 (N_684,In_419,In_249);
nor U685 (N_685,In_183,In_611);
and U686 (N_686,In_15,In_372);
nand U687 (N_687,In_440,In_268);
and U688 (N_688,In_496,In_151);
or U689 (N_689,In_861,In_438);
nor U690 (N_690,In_462,In_129);
nor U691 (N_691,In_878,In_429);
and U692 (N_692,In_807,In_823);
or U693 (N_693,In_639,In_618);
nand U694 (N_694,In_496,In_359);
and U695 (N_695,In_706,In_377);
nor U696 (N_696,In_134,In_309);
nand U697 (N_697,In_111,In_414);
and U698 (N_698,In_247,In_93);
nand U699 (N_699,In_314,In_816);
and U700 (N_700,In_275,In_676);
nand U701 (N_701,In_570,In_400);
nand U702 (N_702,In_670,In_388);
nand U703 (N_703,In_768,In_377);
xor U704 (N_704,In_301,In_847);
or U705 (N_705,In_127,In_744);
and U706 (N_706,In_171,In_820);
nor U707 (N_707,In_219,In_685);
nor U708 (N_708,In_101,In_176);
nor U709 (N_709,In_559,In_973);
nand U710 (N_710,In_193,In_400);
or U711 (N_711,In_768,In_429);
nor U712 (N_712,In_505,In_694);
nor U713 (N_713,In_694,In_740);
and U714 (N_714,In_699,In_654);
or U715 (N_715,In_892,In_201);
xor U716 (N_716,In_492,In_975);
nand U717 (N_717,In_186,In_8);
and U718 (N_718,In_855,In_545);
or U719 (N_719,In_366,In_931);
xnor U720 (N_720,In_2,In_876);
nand U721 (N_721,In_581,In_103);
xnor U722 (N_722,In_677,In_225);
or U723 (N_723,In_564,In_504);
and U724 (N_724,In_916,In_214);
and U725 (N_725,In_121,In_550);
nand U726 (N_726,In_431,In_252);
and U727 (N_727,In_503,In_870);
or U728 (N_728,In_856,In_784);
and U729 (N_729,In_83,In_582);
and U730 (N_730,In_159,In_908);
and U731 (N_731,In_387,In_239);
nor U732 (N_732,In_580,In_156);
nor U733 (N_733,In_125,In_940);
nand U734 (N_734,In_619,In_450);
nor U735 (N_735,In_518,In_725);
or U736 (N_736,In_140,In_19);
nand U737 (N_737,In_533,In_132);
xnor U738 (N_738,In_863,In_426);
or U739 (N_739,In_254,In_337);
or U740 (N_740,In_519,In_82);
nor U741 (N_741,In_318,In_445);
nor U742 (N_742,In_659,In_869);
nand U743 (N_743,In_290,In_823);
nor U744 (N_744,In_315,In_948);
or U745 (N_745,In_928,In_865);
or U746 (N_746,In_74,In_197);
nor U747 (N_747,In_11,In_749);
nor U748 (N_748,In_252,In_9);
and U749 (N_749,In_142,In_763);
nand U750 (N_750,In_942,In_228);
or U751 (N_751,In_676,In_909);
nor U752 (N_752,In_929,In_184);
and U753 (N_753,In_318,In_670);
and U754 (N_754,In_145,In_822);
nor U755 (N_755,In_467,In_544);
or U756 (N_756,In_770,In_275);
nand U757 (N_757,In_707,In_411);
or U758 (N_758,In_931,In_304);
nand U759 (N_759,In_642,In_680);
and U760 (N_760,In_286,In_804);
xnor U761 (N_761,In_611,In_138);
and U762 (N_762,In_697,In_56);
and U763 (N_763,In_568,In_195);
and U764 (N_764,In_431,In_36);
xor U765 (N_765,In_373,In_498);
and U766 (N_766,In_969,In_87);
nand U767 (N_767,In_447,In_724);
and U768 (N_768,In_431,In_982);
or U769 (N_769,In_194,In_604);
nor U770 (N_770,In_118,In_504);
and U771 (N_771,In_850,In_482);
nand U772 (N_772,In_827,In_969);
nor U773 (N_773,In_382,In_562);
nor U774 (N_774,In_798,In_348);
and U775 (N_775,In_605,In_185);
and U776 (N_776,In_500,In_318);
and U777 (N_777,In_709,In_243);
nor U778 (N_778,In_681,In_444);
and U779 (N_779,In_553,In_905);
nor U780 (N_780,In_858,In_734);
nor U781 (N_781,In_63,In_947);
nand U782 (N_782,In_621,In_15);
nand U783 (N_783,In_454,In_994);
nor U784 (N_784,In_643,In_780);
and U785 (N_785,In_893,In_697);
nand U786 (N_786,In_210,In_108);
nand U787 (N_787,In_676,In_101);
or U788 (N_788,In_302,In_17);
or U789 (N_789,In_795,In_251);
and U790 (N_790,In_237,In_803);
nand U791 (N_791,In_699,In_706);
nor U792 (N_792,In_170,In_532);
or U793 (N_793,In_35,In_681);
or U794 (N_794,In_507,In_738);
or U795 (N_795,In_353,In_196);
nand U796 (N_796,In_48,In_915);
nor U797 (N_797,In_683,In_38);
and U798 (N_798,In_154,In_692);
or U799 (N_799,In_272,In_927);
and U800 (N_800,In_257,In_368);
nand U801 (N_801,In_455,In_564);
and U802 (N_802,In_78,In_434);
nor U803 (N_803,In_220,In_266);
nand U804 (N_804,In_449,In_574);
or U805 (N_805,In_332,In_431);
or U806 (N_806,In_186,In_146);
nor U807 (N_807,In_629,In_30);
nand U808 (N_808,In_0,In_893);
nand U809 (N_809,In_926,In_337);
or U810 (N_810,In_832,In_29);
or U811 (N_811,In_895,In_197);
and U812 (N_812,In_399,In_72);
and U813 (N_813,In_760,In_594);
nor U814 (N_814,In_148,In_435);
and U815 (N_815,In_619,In_869);
and U816 (N_816,In_596,In_271);
nand U817 (N_817,In_88,In_179);
nand U818 (N_818,In_966,In_500);
or U819 (N_819,In_526,In_930);
and U820 (N_820,In_918,In_303);
and U821 (N_821,In_75,In_77);
nor U822 (N_822,In_531,In_146);
nand U823 (N_823,In_23,In_243);
or U824 (N_824,In_401,In_650);
nor U825 (N_825,In_577,In_301);
nand U826 (N_826,In_198,In_975);
xnor U827 (N_827,In_158,In_816);
and U828 (N_828,In_603,In_158);
and U829 (N_829,In_244,In_486);
nor U830 (N_830,In_933,In_224);
and U831 (N_831,In_923,In_646);
nand U832 (N_832,In_953,In_246);
nor U833 (N_833,In_450,In_222);
nor U834 (N_834,In_953,In_390);
and U835 (N_835,In_901,In_516);
nor U836 (N_836,In_28,In_978);
and U837 (N_837,In_193,In_25);
or U838 (N_838,In_885,In_999);
or U839 (N_839,In_660,In_665);
and U840 (N_840,In_735,In_776);
or U841 (N_841,In_798,In_674);
or U842 (N_842,In_306,In_96);
or U843 (N_843,In_222,In_187);
nor U844 (N_844,In_247,In_980);
and U845 (N_845,In_390,In_846);
and U846 (N_846,In_586,In_253);
or U847 (N_847,In_104,In_15);
or U848 (N_848,In_241,In_345);
nand U849 (N_849,In_874,In_950);
or U850 (N_850,In_455,In_764);
xor U851 (N_851,In_197,In_706);
nand U852 (N_852,In_582,In_643);
nor U853 (N_853,In_741,In_884);
or U854 (N_854,In_189,In_388);
or U855 (N_855,In_627,In_37);
and U856 (N_856,In_798,In_925);
nor U857 (N_857,In_508,In_185);
nand U858 (N_858,In_873,In_311);
or U859 (N_859,In_342,In_92);
and U860 (N_860,In_813,In_929);
nor U861 (N_861,In_478,In_266);
nand U862 (N_862,In_128,In_585);
nor U863 (N_863,In_209,In_351);
nand U864 (N_864,In_288,In_742);
and U865 (N_865,In_722,In_800);
or U866 (N_866,In_761,In_396);
nor U867 (N_867,In_52,In_60);
or U868 (N_868,In_163,In_10);
and U869 (N_869,In_187,In_995);
nor U870 (N_870,In_149,In_584);
and U871 (N_871,In_77,In_522);
or U872 (N_872,In_636,In_275);
nand U873 (N_873,In_792,In_849);
and U874 (N_874,In_685,In_99);
nor U875 (N_875,In_82,In_319);
or U876 (N_876,In_992,In_437);
or U877 (N_877,In_515,In_859);
and U878 (N_878,In_558,In_621);
and U879 (N_879,In_933,In_265);
and U880 (N_880,In_327,In_368);
and U881 (N_881,In_540,In_556);
xnor U882 (N_882,In_856,In_261);
nor U883 (N_883,In_825,In_115);
nor U884 (N_884,In_342,In_585);
and U885 (N_885,In_825,In_64);
nor U886 (N_886,In_776,In_6);
nor U887 (N_887,In_550,In_125);
and U888 (N_888,In_868,In_392);
nor U889 (N_889,In_977,In_568);
xor U890 (N_890,In_614,In_232);
or U891 (N_891,In_552,In_474);
xnor U892 (N_892,In_698,In_848);
or U893 (N_893,In_996,In_196);
or U894 (N_894,In_354,In_864);
nor U895 (N_895,In_248,In_433);
nor U896 (N_896,In_491,In_433);
and U897 (N_897,In_210,In_417);
or U898 (N_898,In_267,In_781);
nor U899 (N_899,In_933,In_519);
or U900 (N_900,In_135,In_741);
and U901 (N_901,In_368,In_791);
nand U902 (N_902,In_739,In_492);
nor U903 (N_903,In_208,In_989);
nor U904 (N_904,In_55,In_893);
nand U905 (N_905,In_610,In_673);
nand U906 (N_906,In_898,In_910);
nand U907 (N_907,In_295,In_949);
or U908 (N_908,In_285,In_8);
and U909 (N_909,In_779,In_443);
nor U910 (N_910,In_264,In_649);
or U911 (N_911,In_307,In_581);
or U912 (N_912,In_886,In_410);
nor U913 (N_913,In_629,In_973);
or U914 (N_914,In_965,In_73);
nor U915 (N_915,In_734,In_320);
nor U916 (N_916,In_829,In_748);
nor U917 (N_917,In_928,In_851);
and U918 (N_918,In_563,In_180);
nor U919 (N_919,In_333,In_779);
and U920 (N_920,In_278,In_738);
and U921 (N_921,In_725,In_680);
and U922 (N_922,In_7,In_823);
and U923 (N_923,In_483,In_826);
and U924 (N_924,In_922,In_885);
nor U925 (N_925,In_759,In_327);
and U926 (N_926,In_476,In_631);
nor U927 (N_927,In_825,In_255);
nor U928 (N_928,In_457,In_453);
and U929 (N_929,In_79,In_279);
nand U930 (N_930,In_944,In_799);
and U931 (N_931,In_188,In_325);
or U932 (N_932,In_429,In_695);
nand U933 (N_933,In_72,In_15);
or U934 (N_934,In_859,In_324);
nand U935 (N_935,In_529,In_451);
or U936 (N_936,In_796,In_987);
nand U937 (N_937,In_550,In_839);
nand U938 (N_938,In_243,In_927);
nor U939 (N_939,In_159,In_168);
or U940 (N_940,In_364,In_552);
nand U941 (N_941,In_696,In_953);
nor U942 (N_942,In_600,In_982);
and U943 (N_943,In_622,In_318);
and U944 (N_944,In_869,In_794);
and U945 (N_945,In_234,In_236);
nand U946 (N_946,In_686,In_868);
nor U947 (N_947,In_844,In_203);
nor U948 (N_948,In_949,In_88);
nand U949 (N_949,In_523,In_291);
xor U950 (N_950,In_314,In_905);
or U951 (N_951,In_497,In_728);
xor U952 (N_952,In_79,In_643);
nand U953 (N_953,In_876,In_228);
nor U954 (N_954,In_216,In_299);
nor U955 (N_955,In_873,In_937);
nand U956 (N_956,In_566,In_933);
or U957 (N_957,In_604,In_591);
and U958 (N_958,In_742,In_802);
nor U959 (N_959,In_941,In_300);
nand U960 (N_960,In_27,In_322);
and U961 (N_961,In_392,In_631);
nor U962 (N_962,In_521,In_180);
and U963 (N_963,In_600,In_506);
or U964 (N_964,In_920,In_949);
nand U965 (N_965,In_758,In_646);
and U966 (N_966,In_20,In_992);
or U967 (N_967,In_381,In_387);
nor U968 (N_968,In_742,In_956);
nand U969 (N_969,In_38,In_339);
nand U970 (N_970,In_66,In_862);
nor U971 (N_971,In_291,In_102);
and U972 (N_972,In_432,In_3);
nor U973 (N_973,In_3,In_369);
nand U974 (N_974,In_473,In_59);
nand U975 (N_975,In_644,In_556);
nand U976 (N_976,In_184,In_315);
and U977 (N_977,In_376,In_876);
nand U978 (N_978,In_713,In_3);
and U979 (N_979,In_302,In_728);
and U980 (N_980,In_356,In_143);
nand U981 (N_981,In_629,In_386);
nand U982 (N_982,In_597,In_873);
nand U983 (N_983,In_396,In_356);
or U984 (N_984,In_122,In_227);
nand U985 (N_985,In_727,In_554);
nand U986 (N_986,In_165,In_513);
nand U987 (N_987,In_763,In_749);
and U988 (N_988,In_560,In_62);
nand U989 (N_989,In_914,In_245);
and U990 (N_990,In_844,In_721);
nor U991 (N_991,In_592,In_773);
and U992 (N_992,In_779,In_272);
nor U993 (N_993,In_590,In_670);
and U994 (N_994,In_933,In_601);
nand U995 (N_995,In_183,In_136);
or U996 (N_996,In_351,In_658);
nor U997 (N_997,In_207,In_544);
or U998 (N_998,In_74,In_356);
nor U999 (N_999,In_696,In_141);
nor U1000 (N_1000,In_434,In_129);
and U1001 (N_1001,In_844,In_103);
or U1002 (N_1002,In_671,In_165);
nand U1003 (N_1003,In_284,In_770);
xnor U1004 (N_1004,In_84,In_470);
or U1005 (N_1005,In_69,In_455);
or U1006 (N_1006,In_194,In_23);
and U1007 (N_1007,In_168,In_348);
or U1008 (N_1008,In_946,In_969);
and U1009 (N_1009,In_995,In_396);
nor U1010 (N_1010,In_402,In_383);
nand U1011 (N_1011,In_594,In_821);
and U1012 (N_1012,In_295,In_588);
and U1013 (N_1013,In_209,In_374);
nand U1014 (N_1014,In_520,In_591);
and U1015 (N_1015,In_626,In_976);
and U1016 (N_1016,In_905,In_592);
and U1017 (N_1017,In_511,In_683);
and U1018 (N_1018,In_233,In_696);
nor U1019 (N_1019,In_97,In_318);
nand U1020 (N_1020,In_410,In_131);
nand U1021 (N_1021,In_344,In_68);
and U1022 (N_1022,In_49,In_774);
and U1023 (N_1023,In_616,In_185);
nor U1024 (N_1024,In_604,In_257);
nand U1025 (N_1025,In_302,In_95);
nand U1026 (N_1026,In_356,In_253);
nor U1027 (N_1027,In_308,In_720);
and U1028 (N_1028,In_974,In_235);
nor U1029 (N_1029,In_414,In_328);
nand U1030 (N_1030,In_30,In_622);
nor U1031 (N_1031,In_552,In_855);
and U1032 (N_1032,In_863,In_524);
nor U1033 (N_1033,In_49,In_193);
or U1034 (N_1034,In_998,In_610);
nor U1035 (N_1035,In_953,In_276);
or U1036 (N_1036,In_516,In_817);
or U1037 (N_1037,In_93,In_130);
or U1038 (N_1038,In_973,In_3);
xor U1039 (N_1039,In_577,In_290);
nor U1040 (N_1040,In_700,In_663);
or U1041 (N_1041,In_510,In_447);
nor U1042 (N_1042,In_974,In_966);
nand U1043 (N_1043,In_708,In_866);
or U1044 (N_1044,In_879,In_608);
nand U1045 (N_1045,In_375,In_338);
or U1046 (N_1046,In_217,In_267);
and U1047 (N_1047,In_432,In_412);
or U1048 (N_1048,In_507,In_861);
nor U1049 (N_1049,In_283,In_353);
nand U1050 (N_1050,In_756,In_484);
nand U1051 (N_1051,In_118,In_984);
nor U1052 (N_1052,In_175,In_836);
nor U1053 (N_1053,In_8,In_866);
and U1054 (N_1054,In_483,In_217);
nand U1055 (N_1055,In_589,In_539);
nand U1056 (N_1056,In_54,In_461);
or U1057 (N_1057,In_294,In_515);
and U1058 (N_1058,In_162,In_182);
nor U1059 (N_1059,In_45,In_714);
nor U1060 (N_1060,In_69,In_328);
or U1061 (N_1061,In_985,In_60);
or U1062 (N_1062,In_728,In_117);
nor U1063 (N_1063,In_888,In_697);
nor U1064 (N_1064,In_608,In_571);
or U1065 (N_1065,In_373,In_864);
xor U1066 (N_1066,In_158,In_705);
and U1067 (N_1067,In_495,In_210);
and U1068 (N_1068,In_728,In_739);
and U1069 (N_1069,In_800,In_644);
nand U1070 (N_1070,In_176,In_882);
and U1071 (N_1071,In_944,In_361);
and U1072 (N_1072,In_615,In_241);
and U1073 (N_1073,In_492,In_994);
nand U1074 (N_1074,In_174,In_654);
nand U1075 (N_1075,In_358,In_228);
nor U1076 (N_1076,In_340,In_678);
nand U1077 (N_1077,In_27,In_619);
or U1078 (N_1078,In_292,In_920);
and U1079 (N_1079,In_324,In_257);
nor U1080 (N_1080,In_553,In_689);
nor U1081 (N_1081,In_806,In_567);
and U1082 (N_1082,In_2,In_966);
nand U1083 (N_1083,In_893,In_460);
nor U1084 (N_1084,In_136,In_593);
nor U1085 (N_1085,In_807,In_515);
and U1086 (N_1086,In_972,In_466);
nor U1087 (N_1087,In_134,In_929);
or U1088 (N_1088,In_527,In_593);
nor U1089 (N_1089,In_799,In_54);
nand U1090 (N_1090,In_3,In_7);
nand U1091 (N_1091,In_136,In_148);
and U1092 (N_1092,In_283,In_79);
nand U1093 (N_1093,In_37,In_9);
or U1094 (N_1094,In_830,In_569);
and U1095 (N_1095,In_416,In_24);
nor U1096 (N_1096,In_663,In_952);
nand U1097 (N_1097,In_983,In_731);
and U1098 (N_1098,In_836,In_484);
nor U1099 (N_1099,In_45,In_613);
nor U1100 (N_1100,In_7,In_407);
or U1101 (N_1101,In_54,In_427);
nor U1102 (N_1102,In_192,In_895);
and U1103 (N_1103,In_7,In_139);
nand U1104 (N_1104,In_457,In_976);
and U1105 (N_1105,In_507,In_505);
nor U1106 (N_1106,In_755,In_566);
nor U1107 (N_1107,In_404,In_548);
and U1108 (N_1108,In_480,In_156);
and U1109 (N_1109,In_930,In_814);
or U1110 (N_1110,In_65,In_442);
and U1111 (N_1111,In_385,In_147);
and U1112 (N_1112,In_928,In_657);
and U1113 (N_1113,In_418,In_78);
nor U1114 (N_1114,In_606,In_107);
nand U1115 (N_1115,In_601,In_672);
and U1116 (N_1116,In_299,In_708);
and U1117 (N_1117,In_907,In_478);
nand U1118 (N_1118,In_360,In_423);
and U1119 (N_1119,In_290,In_583);
or U1120 (N_1120,In_968,In_211);
and U1121 (N_1121,In_597,In_451);
nor U1122 (N_1122,In_948,In_397);
and U1123 (N_1123,In_926,In_583);
nand U1124 (N_1124,In_694,In_955);
or U1125 (N_1125,In_22,In_855);
or U1126 (N_1126,In_103,In_624);
nand U1127 (N_1127,In_161,In_162);
nand U1128 (N_1128,In_853,In_132);
and U1129 (N_1129,In_343,In_219);
nand U1130 (N_1130,In_650,In_261);
and U1131 (N_1131,In_64,In_520);
nor U1132 (N_1132,In_765,In_991);
and U1133 (N_1133,In_449,In_839);
or U1134 (N_1134,In_703,In_152);
nor U1135 (N_1135,In_891,In_637);
nand U1136 (N_1136,In_470,In_568);
or U1137 (N_1137,In_351,In_825);
or U1138 (N_1138,In_6,In_470);
or U1139 (N_1139,In_613,In_337);
nand U1140 (N_1140,In_964,In_102);
and U1141 (N_1141,In_328,In_849);
nand U1142 (N_1142,In_230,In_577);
and U1143 (N_1143,In_834,In_289);
or U1144 (N_1144,In_684,In_56);
and U1145 (N_1145,In_740,In_175);
and U1146 (N_1146,In_579,In_791);
or U1147 (N_1147,In_534,In_35);
xnor U1148 (N_1148,In_32,In_724);
nor U1149 (N_1149,In_265,In_204);
nand U1150 (N_1150,In_99,In_762);
nand U1151 (N_1151,In_634,In_836);
or U1152 (N_1152,In_263,In_229);
or U1153 (N_1153,In_855,In_20);
nand U1154 (N_1154,In_113,In_187);
nand U1155 (N_1155,In_284,In_300);
nor U1156 (N_1156,In_911,In_562);
nand U1157 (N_1157,In_567,In_633);
nand U1158 (N_1158,In_124,In_86);
nand U1159 (N_1159,In_530,In_162);
or U1160 (N_1160,In_552,In_854);
and U1161 (N_1161,In_451,In_70);
nor U1162 (N_1162,In_642,In_275);
or U1163 (N_1163,In_718,In_511);
xnor U1164 (N_1164,In_206,In_204);
nor U1165 (N_1165,In_369,In_928);
nor U1166 (N_1166,In_50,In_613);
or U1167 (N_1167,In_805,In_253);
and U1168 (N_1168,In_471,In_708);
nand U1169 (N_1169,In_402,In_391);
or U1170 (N_1170,In_10,In_501);
and U1171 (N_1171,In_973,In_602);
nor U1172 (N_1172,In_252,In_490);
nor U1173 (N_1173,In_790,In_113);
nor U1174 (N_1174,In_576,In_316);
nor U1175 (N_1175,In_602,In_441);
nand U1176 (N_1176,In_766,In_74);
or U1177 (N_1177,In_774,In_784);
nor U1178 (N_1178,In_884,In_556);
or U1179 (N_1179,In_253,In_530);
and U1180 (N_1180,In_721,In_13);
nand U1181 (N_1181,In_964,In_907);
nand U1182 (N_1182,In_10,In_760);
and U1183 (N_1183,In_255,In_22);
and U1184 (N_1184,In_481,In_733);
and U1185 (N_1185,In_249,In_616);
nand U1186 (N_1186,In_767,In_96);
nand U1187 (N_1187,In_879,In_916);
or U1188 (N_1188,In_22,In_183);
nand U1189 (N_1189,In_146,In_956);
or U1190 (N_1190,In_137,In_488);
nor U1191 (N_1191,In_579,In_790);
or U1192 (N_1192,In_446,In_794);
and U1193 (N_1193,In_651,In_89);
or U1194 (N_1194,In_968,In_0);
xor U1195 (N_1195,In_789,In_861);
and U1196 (N_1196,In_54,In_613);
or U1197 (N_1197,In_497,In_754);
nor U1198 (N_1198,In_73,In_907);
and U1199 (N_1199,In_935,In_179);
and U1200 (N_1200,In_268,In_75);
nor U1201 (N_1201,In_714,In_657);
xor U1202 (N_1202,In_967,In_502);
nor U1203 (N_1203,In_173,In_284);
and U1204 (N_1204,In_932,In_996);
nor U1205 (N_1205,In_276,In_172);
or U1206 (N_1206,In_994,In_501);
nand U1207 (N_1207,In_907,In_91);
and U1208 (N_1208,In_417,In_934);
and U1209 (N_1209,In_662,In_991);
and U1210 (N_1210,In_321,In_469);
or U1211 (N_1211,In_194,In_94);
and U1212 (N_1212,In_182,In_290);
or U1213 (N_1213,In_302,In_115);
or U1214 (N_1214,In_385,In_930);
nor U1215 (N_1215,In_769,In_572);
nand U1216 (N_1216,In_645,In_77);
nor U1217 (N_1217,In_672,In_813);
nor U1218 (N_1218,In_975,In_120);
or U1219 (N_1219,In_851,In_751);
and U1220 (N_1220,In_893,In_254);
or U1221 (N_1221,In_229,In_351);
and U1222 (N_1222,In_67,In_834);
and U1223 (N_1223,In_193,In_279);
nor U1224 (N_1224,In_184,In_592);
xnor U1225 (N_1225,In_795,In_997);
or U1226 (N_1226,In_543,In_643);
and U1227 (N_1227,In_646,In_431);
or U1228 (N_1228,In_498,In_212);
xnor U1229 (N_1229,In_303,In_346);
and U1230 (N_1230,In_862,In_79);
nor U1231 (N_1231,In_988,In_259);
nor U1232 (N_1232,In_440,In_206);
nand U1233 (N_1233,In_233,In_789);
nor U1234 (N_1234,In_519,In_212);
nor U1235 (N_1235,In_498,In_0);
or U1236 (N_1236,In_413,In_473);
nand U1237 (N_1237,In_49,In_918);
nor U1238 (N_1238,In_661,In_607);
xnor U1239 (N_1239,In_640,In_328);
or U1240 (N_1240,In_128,In_775);
and U1241 (N_1241,In_409,In_808);
nor U1242 (N_1242,In_915,In_82);
nor U1243 (N_1243,In_864,In_997);
or U1244 (N_1244,In_458,In_396);
nand U1245 (N_1245,In_686,In_845);
or U1246 (N_1246,In_728,In_146);
nand U1247 (N_1247,In_996,In_404);
and U1248 (N_1248,In_532,In_673);
nand U1249 (N_1249,In_279,In_204);
and U1250 (N_1250,In_237,In_840);
and U1251 (N_1251,In_160,In_290);
nand U1252 (N_1252,In_331,In_509);
nand U1253 (N_1253,In_357,In_959);
and U1254 (N_1254,In_871,In_544);
or U1255 (N_1255,In_34,In_673);
nand U1256 (N_1256,In_63,In_782);
nand U1257 (N_1257,In_607,In_103);
and U1258 (N_1258,In_301,In_981);
or U1259 (N_1259,In_326,In_717);
nor U1260 (N_1260,In_510,In_275);
nand U1261 (N_1261,In_48,In_198);
or U1262 (N_1262,In_252,In_753);
and U1263 (N_1263,In_498,In_325);
and U1264 (N_1264,In_15,In_52);
nor U1265 (N_1265,In_916,In_100);
nor U1266 (N_1266,In_56,In_76);
or U1267 (N_1267,In_41,In_609);
and U1268 (N_1268,In_642,In_756);
or U1269 (N_1269,In_318,In_644);
and U1270 (N_1270,In_568,In_112);
nor U1271 (N_1271,In_300,In_351);
or U1272 (N_1272,In_932,In_885);
or U1273 (N_1273,In_58,In_955);
or U1274 (N_1274,In_369,In_530);
nand U1275 (N_1275,In_452,In_250);
xor U1276 (N_1276,In_549,In_374);
nor U1277 (N_1277,In_533,In_548);
nand U1278 (N_1278,In_373,In_875);
nor U1279 (N_1279,In_194,In_576);
nand U1280 (N_1280,In_848,In_181);
nand U1281 (N_1281,In_950,In_122);
nand U1282 (N_1282,In_815,In_685);
and U1283 (N_1283,In_916,In_510);
or U1284 (N_1284,In_654,In_921);
nand U1285 (N_1285,In_912,In_234);
nand U1286 (N_1286,In_335,In_904);
nor U1287 (N_1287,In_106,In_426);
xnor U1288 (N_1288,In_792,In_395);
nand U1289 (N_1289,In_108,In_396);
nand U1290 (N_1290,In_543,In_783);
nand U1291 (N_1291,In_687,In_292);
or U1292 (N_1292,In_406,In_909);
nand U1293 (N_1293,In_167,In_765);
nand U1294 (N_1294,In_999,In_524);
and U1295 (N_1295,In_379,In_59);
and U1296 (N_1296,In_499,In_905);
xor U1297 (N_1297,In_138,In_628);
nand U1298 (N_1298,In_598,In_788);
and U1299 (N_1299,In_553,In_699);
and U1300 (N_1300,In_231,In_814);
nor U1301 (N_1301,In_136,In_998);
and U1302 (N_1302,In_167,In_961);
nand U1303 (N_1303,In_86,In_10);
nand U1304 (N_1304,In_890,In_947);
xnor U1305 (N_1305,In_654,In_720);
nand U1306 (N_1306,In_337,In_19);
and U1307 (N_1307,In_581,In_670);
and U1308 (N_1308,In_586,In_477);
xnor U1309 (N_1309,In_296,In_455);
or U1310 (N_1310,In_40,In_376);
and U1311 (N_1311,In_720,In_524);
nor U1312 (N_1312,In_885,In_84);
and U1313 (N_1313,In_322,In_203);
and U1314 (N_1314,In_825,In_168);
and U1315 (N_1315,In_725,In_242);
and U1316 (N_1316,In_497,In_778);
nor U1317 (N_1317,In_836,In_998);
nor U1318 (N_1318,In_573,In_490);
and U1319 (N_1319,In_969,In_900);
and U1320 (N_1320,In_10,In_602);
nor U1321 (N_1321,In_553,In_627);
nand U1322 (N_1322,In_438,In_954);
nand U1323 (N_1323,In_159,In_406);
and U1324 (N_1324,In_535,In_210);
nand U1325 (N_1325,In_746,In_621);
nor U1326 (N_1326,In_406,In_847);
nand U1327 (N_1327,In_11,In_844);
nor U1328 (N_1328,In_382,In_69);
nor U1329 (N_1329,In_718,In_370);
and U1330 (N_1330,In_881,In_606);
nand U1331 (N_1331,In_432,In_126);
and U1332 (N_1332,In_818,In_154);
nor U1333 (N_1333,In_98,In_579);
nor U1334 (N_1334,In_322,In_184);
nand U1335 (N_1335,In_49,In_517);
and U1336 (N_1336,In_475,In_284);
nand U1337 (N_1337,In_583,In_810);
or U1338 (N_1338,In_962,In_899);
nand U1339 (N_1339,In_300,In_108);
and U1340 (N_1340,In_411,In_573);
nand U1341 (N_1341,In_723,In_367);
nand U1342 (N_1342,In_594,In_250);
or U1343 (N_1343,In_923,In_53);
and U1344 (N_1344,In_254,In_342);
and U1345 (N_1345,In_440,In_71);
nor U1346 (N_1346,In_579,In_142);
xnor U1347 (N_1347,In_911,In_13);
nor U1348 (N_1348,In_478,In_294);
nor U1349 (N_1349,In_532,In_616);
nand U1350 (N_1350,In_503,In_996);
and U1351 (N_1351,In_530,In_875);
and U1352 (N_1352,In_443,In_23);
nor U1353 (N_1353,In_150,In_829);
and U1354 (N_1354,In_681,In_772);
or U1355 (N_1355,In_148,In_138);
nand U1356 (N_1356,In_471,In_703);
nand U1357 (N_1357,In_770,In_931);
or U1358 (N_1358,In_73,In_285);
and U1359 (N_1359,In_995,In_826);
and U1360 (N_1360,In_560,In_366);
or U1361 (N_1361,In_545,In_535);
or U1362 (N_1362,In_711,In_212);
and U1363 (N_1363,In_517,In_558);
or U1364 (N_1364,In_594,In_174);
xnor U1365 (N_1365,In_499,In_49);
and U1366 (N_1366,In_996,In_263);
or U1367 (N_1367,In_594,In_534);
nor U1368 (N_1368,In_382,In_752);
nand U1369 (N_1369,In_899,In_969);
or U1370 (N_1370,In_267,In_423);
and U1371 (N_1371,In_998,In_373);
nor U1372 (N_1372,In_663,In_345);
xnor U1373 (N_1373,In_702,In_200);
nand U1374 (N_1374,In_775,In_774);
or U1375 (N_1375,In_226,In_747);
nor U1376 (N_1376,In_43,In_643);
nor U1377 (N_1377,In_227,In_543);
nand U1378 (N_1378,In_22,In_296);
and U1379 (N_1379,In_635,In_196);
and U1380 (N_1380,In_229,In_956);
or U1381 (N_1381,In_748,In_252);
or U1382 (N_1382,In_537,In_27);
nand U1383 (N_1383,In_875,In_610);
nor U1384 (N_1384,In_622,In_573);
nor U1385 (N_1385,In_588,In_306);
or U1386 (N_1386,In_352,In_32);
nand U1387 (N_1387,In_609,In_735);
nor U1388 (N_1388,In_222,In_93);
xnor U1389 (N_1389,In_338,In_0);
and U1390 (N_1390,In_899,In_273);
and U1391 (N_1391,In_670,In_901);
nor U1392 (N_1392,In_676,In_919);
or U1393 (N_1393,In_934,In_433);
and U1394 (N_1394,In_908,In_867);
and U1395 (N_1395,In_38,In_312);
or U1396 (N_1396,In_987,In_708);
or U1397 (N_1397,In_161,In_720);
nor U1398 (N_1398,In_622,In_937);
or U1399 (N_1399,In_750,In_668);
or U1400 (N_1400,In_509,In_79);
or U1401 (N_1401,In_589,In_720);
nand U1402 (N_1402,In_434,In_307);
or U1403 (N_1403,In_339,In_646);
xnor U1404 (N_1404,In_227,In_392);
nand U1405 (N_1405,In_642,In_82);
nor U1406 (N_1406,In_939,In_791);
or U1407 (N_1407,In_314,In_714);
nor U1408 (N_1408,In_476,In_878);
nor U1409 (N_1409,In_719,In_46);
xnor U1410 (N_1410,In_65,In_652);
nor U1411 (N_1411,In_700,In_739);
or U1412 (N_1412,In_810,In_726);
nand U1413 (N_1413,In_67,In_423);
and U1414 (N_1414,In_541,In_579);
xor U1415 (N_1415,In_875,In_494);
nor U1416 (N_1416,In_990,In_385);
or U1417 (N_1417,In_575,In_796);
or U1418 (N_1418,In_135,In_804);
nor U1419 (N_1419,In_305,In_711);
and U1420 (N_1420,In_685,In_974);
nand U1421 (N_1421,In_674,In_660);
and U1422 (N_1422,In_362,In_331);
xor U1423 (N_1423,In_262,In_950);
or U1424 (N_1424,In_518,In_900);
or U1425 (N_1425,In_366,In_852);
or U1426 (N_1426,In_192,In_601);
nand U1427 (N_1427,In_390,In_74);
and U1428 (N_1428,In_652,In_517);
nand U1429 (N_1429,In_81,In_471);
or U1430 (N_1430,In_330,In_400);
and U1431 (N_1431,In_173,In_783);
nand U1432 (N_1432,In_163,In_625);
or U1433 (N_1433,In_972,In_562);
or U1434 (N_1434,In_339,In_66);
nand U1435 (N_1435,In_898,In_509);
and U1436 (N_1436,In_401,In_38);
or U1437 (N_1437,In_981,In_373);
and U1438 (N_1438,In_105,In_743);
nor U1439 (N_1439,In_940,In_368);
or U1440 (N_1440,In_730,In_831);
or U1441 (N_1441,In_221,In_537);
and U1442 (N_1442,In_656,In_127);
nor U1443 (N_1443,In_224,In_846);
xor U1444 (N_1444,In_202,In_933);
and U1445 (N_1445,In_116,In_569);
or U1446 (N_1446,In_860,In_747);
xor U1447 (N_1447,In_627,In_649);
and U1448 (N_1448,In_7,In_629);
nand U1449 (N_1449,In_606,In_93);
and U1450 (N_1450,In_565,In_227);
and U1451 (N_1451,In_749,In_365);
nand U1452 (N_1452,In_835,In_10);
and U1453 (N_1453,In_855,In_648);
or U1454 (N_1454,In_649,In_915);
or U1455 (N_1455,In_778,In_480);
or U1456 (N_1456,In_795,In_432);
or U1457 (N_1457,In_779,In_771);
and U1458 (N_1458,In_117,In_444);
and U1459 (N_1459,In_973,In_68);
and U1460 (N_1460,In_690,In_116);
nand U1461 (N_1461,In_991,In_795);
nor U1462 (N_1462,In_915,In_861);
xnor U1463 (N_1463,In_978,In_90);
and U1464 (N_1464,In_693,In_455);
or U1465 (N_1465,In_656,In_384);
or U1466 (N_1466,In_741,In_604);
nand U1467 (N_1467,In_680,In_369);
nor U1468 (N_1468,In_595,In_317);
xnor U1469 (N_1469,In_789,In_801);
and U1470 (N_1470,In_670,In_240);
nor U1471 (N_1471,In_231,In_193);
nor U1472 (N_1472,In_497,In_987);
and U1473 (N_1473,In_978,In_690);
nor U1474 (N_1474,In_14,In_475);
or U1475 (N_1475,In_495,In_106);
nor U1476 (N_1476,In_498,In_610);
or U1477 (N_1477,In_51,In_121);
nand U1478 (N_1478,In_761,In_262);
nand U1479 (N_1479,In_231,In_993);
nor U1480 (N_1480,In_117,In_399);
nand U1481 (N_1481,In_16,In_800);
nand U1482 (N_1482,In_773,In_844);
nand U1483 (N_1483,In_113,In_393);
nand U1484 (N_1484,In_202,In_373);
or U1485 (N_1485,In_73,In_797);
or U1486 (N_1486,In_758,In_345);
nor U1487 (N_1487,In_917,In_395);
nand U1488 (N_1488,In_184,In_379);
and U1489 (N_1489,In_613,In_118);
or U1490 (N_1490,In_634,In_536);
nand U1491 (N_1491,In_130,In_576);
or U1492 (N_1492,In_344,In_256);
nand U1493 (N_1493,In_882,In_330);
or U1494 (N_1494,In_833,In_547);
nand U1495 (N_1495,In_476,In_41);
nand U1496 (N_1496,In_470,In_582);
xor U1497 (N_1497,In_54,In_33);
nor U1498 (N_1498,In_305,In_600);
or U1499 (N_1499,In_460,In_387);
or U1500 (N_1500,In_406,In_718);
or U1501 (N_1501,In_792,In_101);
and U1502 (N_1502,In_323,In_187);
and U1503 (N_1503,In_146,In_211);
nand U1504 (N_1504,In_708,In_462);
nand U1505 (N_1505,In_818,In_379);
nor U1506 (N_1506,In_749,In_816);
nor U1507 (N_1507,In_135,In_70);
nor U1508 (N_1508,In_713,In_151);
xnor U1509 (N_1509,In_37,In_411);
nand U1510 (N_1510,In_131,In_914);
and U1511 (N_1511,In_160,In_32);
nor U1512 (N_1512,In_512,In_464);
nor U1513 (N_1513,In_361,In_398);
nand U1514 (N_1514,In_969,In_173);
or U1515 (N_1515,In_239,In_289);
nor U1516 (N_1516,In_346,In_858);
and U1517 (N_1517,In_68,In_717);
nand U1518 (N_1518,In_87,In_480);
and U1519 (N_1519,In_764,In_32);
nand U1520 (N_1520,In_340,In_352);
nand U1521 (N_1521,In_971,In_498);
or U1522 (N_1522,In_355,In_10);
and U1523 (N_1523,In_44,In_155);
or U1524 (N_1524,In_447,In_754);
and U1525 (N_1525,In_479,In_199);
and U1526 (N_1526,In_805,In_897);
nand U1527 (N_1527,In_710,In_820);
and U1528 (N_1528,In_941,In_545);
and U1529 (N_1529,In_208,In_288);
or U1530 (N_1530,In_860,In_887);
and U1531 (N_1531,In_801,In_350);
nor U1532 (N_1532,In_683,In_765);
and U1533 (N_1533,In_711,In_640);
nand U1534 (N_1534,In_844,In_626);
nor U1535 (N_1535,In_752,In_288);
nand U1536 (N_1536,In_977,In_243);
and U1537 (N_1537,In_57,In_324);
and U1538 (N_1538,In_789,In_505);
or U1539 (N_1539,In_226,In_390);
or U1540 (N_1540,In_357,In_168);
or U1541 (N_1541,In_225,In_503);
or U1542 (N_1542,In_86,In_320);
and U1543 (N_1543,In_474,In_844);
nor U1544 (N_1544,In_233,In_218);
nand U1545 (N_1545,In_983,In_699);
and U1546 (N_1546,In_66,In_893);
and U1547 (N_1547,In_724,In_371);
nand U1548 (N_1548,In_383,In_795);
nand U1549 (N_1549,In_880,In_432);
or U1550 (N_1550,In_263,In_886);
and U1551 (N_1551,In_394,In_531);
nor U1552 (N_1552,In_175,In_636);
nor U1553 (N_1553,In_202,In_309);
nor U1554 (N_1554,In_88,In_922);
and U1555 (N_1555,In_613,In_946);
nand U1556 (N_1556,In_549,In_841);
and U1557 (N_1557,In_862,In_307);
or U1558 (N_1558,In_663,In_327);
or U1559 (N_1559,In_360,In_197);
and U1560 (N_1560,In_17,In_522);
nand U1561 (N_1561,In_176,In_879);
nor U1562 (N_1562,In_484,In_916);
and U1563 (N_1563,In_500,In_465);
nor U1564 (N_1564,In_547,In_317);
nor U1565 (N_1565,In_95,In_292);
or U1566 (N_1566,In_96,In_418);
and U1567 (N_1567,In_417,In_955);
nor U1568 (N_1568,In_522,In_248);
or U1569 (N_1569,In_271,In_531);
or U1570 (N_1570,In_508,In_601);
nand U1571 (N_1571,In_321,In_919);
or U1572 (N_1572,In_553,In_380);
and U1573 (N_1573,In_195,In_114);
nor U1574 (N_1574,In_601,In_710);
or U1575 (N_1575,In_696,In_985);
xnor U1576 (N_1576,In_57,In_367);
and U1577 (N_1577,In_925,In_520);
nand U1578 (N_1578,In_135,In_0);
nand U1579 (N_1579,In_519,In_353);
nand U1580 (N_1580,In_656,In_573);
and U1581 (N_1581,In_499,In_562);
or U1582 (N_1582,In_503,In_962);
and U1583 (N_1583,In_941,In_268);
or U1584 (N_1584,In_670,In_232);
nand U1585 (N_1585,In_507,In_657);
nand U1586 (N_1586,In_879,In_967);
and U1587 (N_1587,In_43,In_296);
or U1588 (N_1588,In_942,In_896);
nor U1589 (N_1589,In_346,In_420);
and U1590 (N_1590,In_521,In_93);
and U1591 (N_1591,In_79,In_599);
nor U1592 (N_1592,In_52,In_923);
or U1593 (N_1593,In_807,In_898);
nor U1594 (N_1594,In_256,In_288);
and U1595 (N_1595,In_407,In_296);
or U1596 (N_1596,In_907,In_739);
nor U1597 (N_1597,In_59,In_864);
nor U1598 (N_1598,In_789,In_917);
nand U1599 (N_1599,In_871,In_941);
and U1600 (N_1600,In_978,In_18);
or U1601 (N_1601,In_456,In_512);
nand U1602 (N_1602,In_45,In_725);
or U1603 (N_1603,In_3,In_691);
and U1604 (N_1604,In_382,In_563);
xnor U1605 (N_1605,In_189,In_413);
xnor U1606 (N_1606,In_324,In_721);
nand U1607 (N_1607,In_336,In_717);
nand U1608 (N_1608,In_506,In_441);
nand U1609 (N_1609,In_435,In_486);
nor U1610 (N_1610,In_754,In_863);
nor U1611 (N_1611,In_968,In_20);
or U1612 (N_1612,In_874,In_414);
nand U1613 (N_1613,In_42,In_231);
or U1614 (N_1614,In_981,In_733);
nand U1615 (N_1615,In_876,In_907);
and U1616 (N_1616,In_216,In_247);
or U1617 (N_1617,In_993,In_825);
xor U1618 (N_1618,In_63,In_558);
or U1619 (N_1619,In_879,In_752);
nand U1620 (N_1620,In_105,In_967);
or U1621 (N_1621,In_828,In_614);
nand U1622 (N_1622,In_905,In_114);
or U1623 (N_1623,In_924,In_100);
and U1624 (N_1624,In_963,In_356);
and U1625 (N_1625,In_821,In_521);
nand U1626 (N_1626,In_208,In_502);
nand U1627 (N_1627,In_903,In_293);
nand U1628 (N_1628,In_191,In_343);
or U1629 (N_1629,In_569,In_219);
nor U1630 (N_1630,In_71,In_368);
and U1631 (N_1631,In_387,In_631);
and U1632 (N_1632,In_724,In_425);
nand U1633 (N_1633,In_681,In_371);
or U1634 (N_1634,In_617,In_598);
and U1635 (N_1635,In_909,In_135);
nand U1636 (N_1636,In_531,In_721);
or U1637 (N_1637,In_896,In_203);
and U1638 (N_1638,In_272,In_208);
xnor U1639 (N_1639,In_324,In_31);
nand U1640 (N_1640,In_355,In_584);
nand U1641 (N_1641,In_595,In_571);
nand U1642 (N_1642,In_520,In_442);
or U1643 (N_1643,In_844,In_665);
and U1644 (N_1644,In_768,In_430);
nor U1645 (N_1645,In_10,In_954);
nand U1646 (N_1646,In_480,In_748);
nand U1647 (N_1647,In_824,In_684);
or U1648 (N_1648,In_823,In_670);
or U1649 (N_1649,In_280,In_519);
nor U1650 (N_1650,In_902,In_853);
nand U1651 (N_1651,In_975,In_908);
or U1652 (N_1652,In_111,In_62);
nand U1653 (N_1653,In_845,In_273);
nor U1654 (N_1654,In_728,In_79);
or U1655 (N_1655,In_220,In_801);
and U1656 (N_1656,In_156,In_607);
nand U1657 (N_1657,In_953,In_772);
or U1658 (N_1658,In_870,In_372);
and U1659 (N_1659,In_870,In_685);
and U1660 (N_1660,In_999,In_80);
nand U1661 (N_1661,In_181,In_817);
and U1662 (N_1662,In_322,In_71);
nor U1663 (N_1663,In_313,In_397);
or U1664 (N_1664,In_878,In_581);
and U1665 (N_1665,In_537,In_455);
nand U1666 (N_1666,In_848,In_272);
or U1667 (N_1667,In_882,In_311);
nor U1668 (N_1668,In_44,In_218);
nand U1669 (N_1669,In_109,In_515);
and U1670 (N_1670,In_94,In_733);
or U1671 (N_1671,In_556,In_215);
nand U1672 (N_1672,In_701,In_855);
nor U1673 (N_1673,In_873,In_498);
nand U1674 (N_1674,In_449,In_676);
or U1675 (N_1675,In_118,In_54);
or U1676 (N_1676,In_611,In_173);
nand U1677 (N_1677,In_217,In_210);
nor U1678 (N_1678,In_656,In_789);
and U1679 (N_1679,In_562,In_5);
nand U1680 (N_1680,In_482,In_113);
nor U1681 (N_1681,In_702,In_836);
nand U1682 (N_1682,In_687,In_830);
or U1683 (N_1683,In_145,In_828);
or U1684 (N_1684,In_121,In_951);
nand U1685 (N_1685,In_864,In_99);
nand U1686 (N_1686,In_939,In_772);
nor U1687 (N_1687,In_733,In_577);
nand U1688 (N_1688,In_668,In_394);
and U1689 (N_1689,In_706,In_962);
and U1690 (N_1690,In_6,In_921);
nand U1691 (N_1691,In_344,In_466);
nand U1692 (N_1692,In_859,In_780);
and U1693 (N_1693,In_189,In_252);
nor U1694 (N_1694,In_540,In_806);
nor U1695 (N_1695,In_631,In_86);
or U1696 (N_1696,In_80,In_167);
nor U1697 (N_1697,In_277,In_706);
nand U1698 (N_1698,In_214,In_444);
nor U1699 (N_1699,In_966,In_835);
or U1700 (N_1700,In_154,In_535);
or U1701 (N_1701,In_394,In_93);
xnor U1702 (N_1702,In_52,In_720);
or U1703 (N_1703,In_882,In_990);
and U1704 (N_1704,In_325,In_840);
nand U1705 (N_1705,In_541,In_442);
or U1706 (N_1706,In_451,In_235);
or U1707 (N_1707,In_522,In_75);
or U1708 (N_1708,In_778,In_224);
nor U1709 (N_1709,In_824,In_968);
nor U1710 (N_1710,In_872,In_391);
and U1711 (N_1711,In_986,In_676);
nand U1712 (N_1712,In_911,In_678);
and U1713 (N_1713,In_478,In_438);
nor U1714 (N_1714,In_349,In_589);
or U1715 (N_1715,In_915,In_711);
nor U1716 (N_1716,In_508,In_212);
or U1717 (N_1717,In_61,In_648);
nand U1718 (N_1718,In_543,In_912);
nand U1719 (N_1719,In_328,In_413);
nor U1720 (N_1720,In_220,In_362);
nor U1721 (N_1721,In_80,In_869);
nand U1722 (N_1722,In_361,In_849);
nor U1723 (N_1723,In_372,In_847);
and U1724 (N_1724,In_319,In_474);
or U1725 (N_1725,In_816,In_533);
or U1726 (N_1726,In_446,In_205);
or U1727 (N_1727,In_423,In_648);
and U1728 (N_1728,In_857,In_625);
and U1729 (N_1729,In_259,In_594);
and U1730 (N_1730,In_804,In_730);
nor U1731 (N_1731,In_587,In_755);
or U1732 (N_1732,In_681,In_565);
nand U1733 (N_1733,In_717,In_676);
nand U1734 (N_1734,In_456,In_159);
or U1735 (N_1735,In_937,In_28);
nor U1736 (N_1736,In_664,In_802);
or U1737 (N_1737,In_465,In_367);
and U1738 (N_1738,In_566,In_42);
or U1739 (N_1739,In_769,In_713);
or U1740 (N_1740,In_332,In_845);
or U1741 (N_1741,In_625,In_59);
and U1742 (N_1742,In_107,In_180);
xor U1743 (N_1743,In_392,In_38);
nor U1744 (N_1744,In_594,In_673);
nand U1745 (N_1745,In_924,In_29);
and U1746 (N_1746,In_706,In_766);
nand U1747 (N_1747,In_42,In_485);
or U1748 (N_1748,In_559,In_486);
and U1749 (N_1749,In_378,In_162);
nand U1750 (N_1750,In_602,In_67);
and U1751 (N_1751,In_947,In_570);
and U1752 (N_1752,In_137,In_698);
or U1753 (N_1753,In_260,In_643);
nand U1754 (N_1754,In_56,In_679);
or U1755 (N_1755,In_916,In_672);
nand U1756 (N_1756,In_540,In_10);
nor U1757 (N_1757,In_175,In_349);
and U1758 (N_1758,In_824,In_884);
nand U1759 (N_1759,In_109,In_248);
nor U1760 (N_1760,In_407,In_886);
and U1761 (N_1761,In_34,In_253);
nand U1762 (N_1762,In_956,In_543);
or U1763 (N_1763,In_859,In_49);
nand U1764 (N_1764,In_313,In_909);
nor U1765 (N_1765,In_954,In_719);
nor U1766 (N_1766,In_580,In_672);
nand U1767 (N_1767,In_471,In_915);
or U1768 (N_1768,In_470,In_893);
or U1769 (N_1769,In_101,In_139);
or U1770 (N_1770,In_832,In_87);
and U1771 (N_1771,In_527,In_218);
and U1772 (N_1772,In_657,In_587);
nand U1773 (N_1773,In_132,In_767);
or U1774 (N_1774,In_77,In_354);
nand U1775 (N_1775,In_75,In_744);
and U1776 (N_1776,In_928,In_821);
nor U1777 (N_1777,In_72,In_948);
and U1778 (N_1778,In_441,In_589);
or U1779 (N_1779,In_996,In_884);
nand U1780 (N_1780,In_191,In_7);
nor U1781 (N_1781,In_635,In_433);
nand U1782 (N_1782,In_96,In_22);
or U1783 (N_1783,In_742,In_662);
or U1784 (N_1784,In_599,In_514);
nor U1785 (N_1785,In_737,In_829);
and U1786 (N_1786,In_704,In_973);
nor U1787 (N_1787,In_764,In_919);
nand U1788 (N_1788,In_134,In_955);
and U1789 (N_1789,In_721,In_553);
and U1790 (N_1790,In_936,In_642);
and U1791 (N_1791,In_295,In_571);
and U1792 (N_1792,In_144,In_786);
and U1793 (N_1793,In_796,In_968);
or U1794 (N_1794,In_43,In_81);
or U1795 (N_1795,In_777,In_439);
nor U1796 (N_1796,In_136,In_594);
or U1797 (N_1797,In_130,In_733);
or U1798 (N_1798,In_266,In_342);
and U1799 (N_1799,In_702,In_675);
nor U1800 (N_1800,In_898,In_727);
or U1801 (N_1801,In_224,In_123);
and U1802 (N_1802,In_54,In_795);
nand U1803 (N_1803,In_808,In_18);
nand U1804 (N_1804,In_916,In_503);
nor U1805 (N_1805,In_590,In_331);
nor U1806 (N_1806,In_256,In_948);
nor U1807 (N_1807,In_941,In_496);
and U1808 (N_1808,In_200,In_767);
and U1809 (N_1809,In_721,In_774);
nand U1810 (N_1810,In_928,In_395);
nor U1811 (N_1811,In_742,In_810);
nor U1812 (N_1812,In_415,In_927);
nor U1813 (N_1813,In_86,In_488);
and U1814 (N_1814,In_392,In_418);
and U1815 (N_1815,In_532,In_775);
or U1816 (N_1816,In_471,In_786);
nand U1817 (N_1817,In_830,In_18);
or U1818 (N_1818,In_113,In_462);
or U1819 (N_1819,In_619,In_252);
and U1820 (N_1820,In_210,In_515);
or U1821 (N_1821,In_605,In_132);
or U1822 (N_1822,In_867,In_304);
or U1823 (N_1823,In_745,In_112);
or U1824 (N_1824,In_446,In_221);
nand U1825 (N_1825,In_18,In_866);
xnor U1826 (N_1826,In_80,In_248);
and U1827 (N_1827,In_635,In_537);
and U1828 (N_1828,In_47,In_48);
nor U1829 (N_1829,In_476,In_77);
nand U1830 (N_1830,In_904,In_7);
nand U1831 (N_1831,In_13,In_95);
or U1832 (N_1832,In_202,In_507);
and U1833 (N_1833,In_773,In_207);
or U1834 (N_1834,In_459,In_196);
nand U1835 (N_1835,In_187,In_79);
or U1836 (N_1836,In_815,In_410);
or U1837 (N_1837,In_354,In_936);
nand U1838 (N_1838,In_222,In_363);
and U1839 (N_1839,In_787,In_96);
and U1840 (N_1840,In_770,In_392);
nand U1841 (N_1841,In_24,In_868);
nor U1842 (N_1842,In_932,In_448);
nor U1843 (N_1843,In_947,In_29);
and U1844 (N_1844,In_605,In_139);
or U1845 (N_1845,In_955,In_740);
nand U1846 (N_1846,In_831,In_494);
and U1847 (N_1847,In_946,In_688);
or U1848 (N_1848,In_905,In_595);
nand U1849 (N_1849,In_373,In_760);
and U1850 (N_1850,In_78,In_747);
and U1851 (N_1851,In_447,In_548);
nor U1852 (N_1852,In_342,In_802);
nand U1853 (N_1853,In_415,In_380);
nor U1854 (N_1854,In_673,In_171);
or U1855 (N_1855,In_615,In_505);
or U1856 (N_1856,In_728,In_64);
nor U1857 (N_1857,In_912,In_368);
and U1858 (N_1858,In_45,In_380);
nand U1859 (N_1859,In_920,In_715);
nand U1860 (N_1860,In_630,In_109);
nor U1861 (N_1861,In_842,In_662);
nor U1862 (N_1862,In_964,In_681);
nor U1863 (N_1863,In_883,In_318);
nor U1864 (N_1864,In_995,In_417);
or U1865 (N_1865,In_972,In_654);
nor U1866 (N_1866,In_709,In_266);
or U1867 (N_1867,In_751,In_82);
or U1868 (N_1868,In_512,In_557);
and U1869 (N_1869,In_492,In_68);
and U1870 (N_1870,In_450,In_983);
nor U1871 (N_1871,In_694,In_682);
nand U1872 (N_1872,In_817,In_869);
and U1873 (N_1873,In_238,In_818);
xor U1874 (N_1874,In_568,In_577);
or U1875 (N_1875,In_826,In_670);
and U1876 (N_1876,In_559,In_899);
and U1877 (N_1877,In_957,In_247);
nand U1878 (N_1878,In_735,In_143);
nor U1879 (N_1879,In_37,In_593);
nand U1880 (N_1880,In_586,In_427);
or U1881 (N_1881,In_448,In_473);
or U1882 (N_1882,In_790,In_857);
or U1883 (N_1883,In_177,In_885);
and U1884 (N_1884,In_930,In_807);
and U1885 (N_1885,In_584,In_239);
and U1886 (N_1886,In_411,In_825);
or U1887 (N_1887,In_529,In_406);
nand U1888 (N_1888,In_561,In_68);
or U1889 (N_1889,In_729,In_68);
or U1890 (N_1890,In_263,In_241);
nand U1891 (N_1891,In_344,In_970);
nand U1892 (N_1892,In_885,In_534);
nand U1893 (N_1893,In_668,In_851);
or U1894 (N_1894,In_296,In_304);
and U1895 (N_1895,In_544,In_616);
and U1896 (N_1896,In_323,In_126);
nor U1897 (N_1897,In_186,In_29);
nor U1898 (N_1898,In_980,In_697);
and U1899 (N_1899,In_926,In_629);
or U1900 (N_1900,In_746,In_375);
and U1901 (N_1901,In_565,In_948);
nand U1902 (N_1902,In_130,In_456);
nor U1903 (N_1903,In_170,In_552);
nand U1904 (N_1904,In_13,In_316);
or U1905 (N_1905,In_345,In_752);
nor U1906 (N_1906,In_528,In_224);
nand U1907 (N_1907,In_66,In_698);
nor U1908 (N_1908,In_707,In_624);
or U1909 (N_1909,In_314,In_653);
or U1910 (N_1910,In_628,In_554);
and U1911 (N_1911,In_540,In_360);
xnor U1912 (N_1912,In_518,In_430);
nand U1913 (N_1913,In_126,In_105);
and U1914 (N_1914,In_219,In_861);
and U1915 (N_1915,In_741,In_39);
or U1916 (N_1916,In_437,In_14);
or U1917 (N_1917,In_493,In_644);
nand U1918 (N_1918,In_877,In_616);
nor U1919 (N_1919,In_100,In_678);
nor U1920 (N_1920,In_130,In_39);
nand U1921 (N_1921,In_497,In_709);
and U1922 (N_1922,In_474,In_364);
or U1923 (N_1923,In_619,In_416);
nor U1924 (N_1924,In_924,In_571);
nand U1925 (N_1925,In_813,In_616);
and U1926 (N_1926,In_717,In_404);
nand U1927 (N_1927,In_16,In_763);
nand U1928 (N_1928,In_505,In_64);
or U1929 (N_1929,In_790,In_509);
or U1930 (N_1930,In_953,In_510);
xnor U1931 (N_1931,In_834,In_179);
and U1932 (N_1932,In_685,In_437);
nand U1933 (N_1933,In_341,In_172);
or U1934 (N_1934,In_147,In_239);
and U1935 (N_1935,In_573,In_645);
nor U1936 (N_1936,In_954,In_654);
nand U1937 (N_1937,In_396,In_444);
or U1938 (N_1938,In_191,In_565);
nor U1939 (N_1939,In_911,In_436);
and U1940 (N_1940,In_876,In_312);
nor U1941 (N_1941,In_206,In_310);
or U1942 (N_1942,In_878,In_4);
and U1943 (N_1943,In_504,In_858);
nor U1944 (N_1944,In_897,In_675);
nor U1945 (N_1945,In_593,In_409);
nand U1946 (N_1946,In_380,In_54);
or U1947 (N_1947,In_858,In_494);
nand U1948 (N_1948,In_658,In_180);
and U1949 (N_1949,In_101,In_862);
or U1950 (N_1950,In_245,In_695);
and U1951 (N_1951,In_744,In_7);
nor U1952 (N_1952,In_855,In_96);
or U1953 (N_1953,In_222,In_599);
or U1954 (N_1954,In_659,In_12);
nand U1955 (N_1955,In_320,In_689);
xnor U1956 (N_1956,In_43,In_345);
xor U1957 (N_1957,In_996,In_388);
nand U1958 (N_1958,In_54,In_675);
and U1959 (N_1959,In_477,In_504);
or U1960 (N_1960,In_972,In_314);
and U1961 (N_1961,In_234,In_370);
nor U1962 (N_1962,In_879,In_932);
nand U1963 (N_1963,In_248,In_216);
nor U1964 (N_1964,In_41,In_720);
and U1965 (N_1965,In_633,In_653);
nor U1966 (N_1966,In_273,In_208);
or U1967 (N_1967,In_684,In_958);
nor U1968 (N_1968,In_815,In_25);
or U1969 (N_1969,In_308,In_772);
nor U1970 (N_1970,In_821,In_101);
nand U1971 (N_1971,In_445,In_254);
and U1972 (N_1972,In_658,In_379);
and U1973 (N_1973,In_205,In_768);
or U1974 (N_1974,In_977,In_619);
and U1975 (N_1975,In_514,In_823);
nand U1976 (N_1976,In_868,In_411);
or U1977 (N_1977,In_976,In_818);
nor U1978 (N_1978,In_308,In_793);
nor U1979 (N_1979,In_167,In_685);
nor U1980 (N_1980,In_901,In_677);
nand U1981 (N_1981,In_877,In_608);
nor U1982 (N_1982,In_909,In_176);
nand U1983 (N_1983,In_171,In_925);
or U1984 (N_1984,In_42,In_576);
nand U1985 (N_1985,In_273,In_132);
nand U1986 (N_1986,In_47,In_670);
nor U1987 (N_1987,In_144,In_988);
nand U1988 (N_1988,In_137,In_621);
nand U1989 (N_1989,In_296,In_634);
and U1990 (N_1990,In_936,In_856);
nor U1991 (N_1991,In_341,In_967);
nor U1992 (N_1992,In_230,In_864);
nor U1993 (N_1993,In_81,In_214);
and U1994 (N_1994,In_253,In_20);
nor U1995 (N_1995,In_402,In_102);
or U1996 (N_1996,In_103,In_794);
or U1997 (N_1997,In_249,In_170);
nor U1998 (N_1998,In_706,In_826);
and U1999 (N_1999,In_563,In_482);
or U2000 (N_2000,In_484,In_466);
xnor U2001 (N_2001,In_729,In_67);
nor U2002 (N_2002,In_987,In_941);
and U2003 (N_2003,In_193,In_576);
or U2004 (N_2004,In_717,In_260);
nand U2005 (N_2005,In_855,In_116);
nor U2006 (N_2006,In_725,In_346);
xnor U2007 (N_2007,In_336,In_948);
nand U2008 (N_2008,In_771,In_319);
nand U2009 (N_2009,In_200,In_711);
and U2010 (N_2010,In_12,In_290);
and U2011 (N_2011,In_535,In_692);
or U2012 (N_2012,In_633,In_472);
or U2013 (N_2013,In_707,In_571);
nand U2014 (N_2014,In_745,In_780);
or U2015 (N_2015,In_84,In_227);
nor U2016 (N_2016,In_215,In_757);
nor U2017 (N_2017,In_106,In_89);
nor U2018 (N_2018,In_542,In_822);
or U2019 (N_2019,In_85,In_337);
nand U2020 (N_2020,In_571,In_366);
nor U2021 (N_2021,In_761,In_783);
nand U2022 (N_2022,In_265,In_470);
or U2023 (N_2023,In_646,In_174);
nor U2024 (N_2024,In_19,In_677);
and U2025 (N_2025,In_588,In_864);
nand U2026 (N_2026,In_721,In_479);
nor U2027 (N_2027,In_935,In_975);
or U2028 (N_2028,In_428,In_982);
nor U2029 (N_2029,In_989,In_315);
nor U2030 (N_2030,In_595,In_12);
nand U2031 (N_2031,In_593,In_10);
xnor U2032 (N_2032,In_330,In_968);
and U2033 (N_2033,In_685,In_500);
or U2034 (N_2034,In_483,In_622);
nand U2035 (N_2035,In_167,In_860);
or U2036 (N_2036,In_677,In_403);
or U2037 (N_2037,In_918,In_556);
nand U2038 (N_2038,In_820,In_725);
and U2039 (N_2039,In_414,In_124);
or U2040 (N_2040,In_849,In_450);
nand U2041 (N_2041,In_651,In_355);
nand U2042 (N_2042,In_31,In_201);
xor U2043 (N_2043,In_79,In_733);
nand U2044 (N_2044,In_189,In_320);
and U2045 (N_2045,In_616,In_273);
and U2046 (N_2046,In_411,In_528);
and U2047 (N_2047,In_91,In_437);
nand U2048 (N_2048,In_505,In_748);
or U2049 (N_2049,In_202,In_257);
nand U2050 (N_2050,In_758,In_133);
nor U2051 (N_2051,In_230,In_43);
and U2052 (N_2052,In_675,In_427);
or U2053 (N_2053,In_380,In_296);
nand U2054 (N_2054,In_309,In_225);
nor U2055 (N_2055,In_394,In_719);
nand U2056 (N_2056,In_146,In_248);
xnor U2057 (N_2057,In_672,In_178);
or U2058 (N_2058,In_72,In_20);
or U2059 (N_2059,In_206,In_446);
nand U2060 (N_2060,In_655,In_462);
and U2061 (N_2061,In_44,In_564);
nand U2062 (N_2062,In_150,In_416);
nand U2063 (N_2063,In_818,In_109);
nor U2064 (N_2064,In_100,In_169);
and U2065 (N_2065,In_772,In_500);
xor U2066 (N_2066,In_832,In_753);
nor U2067 (N_2067,In_958,In_613);
xnor U2068 (N_2068,In_85,In_994);
nor U2069 (N_2069,In_804,In_888);
and U2070 (N_2070,In_73,In_925);
and U2071 (N_2071,In_777,In_877);
nand U2072 (N_2072,In_968,In_938);
xnor U2073 (N_2073,In_872,In_922);
and U2074 (N_2074,In_758,In_680);
nand U2075 (N_2075,In_375,In_943);
or U2076 (N_2076,In_39,In_988);
nor U2077 (N_2077,In_76,In_191);
and U2078 (N_2078,In_509,In_432);
nor U2079 (N_2079,In_994,In_886);
nor U2080 (N_2080,In_620,In_212);
or U2081 (N_2081,In_519,In_39);
and U2082 (N_2082,In_952,In_62);
and U2083 (N_2083,In_558,In_133);
nor U2084 (N_2084,In_844,In_238);
and U2085 (N_2085,In_460,In_378);
and U2086 (N_2086,In_516,In_703);
nor U2087 (N_2087,In_36,In_434);
nor U2088 (N_2088,In_73,In_589);
or U2089 (N_2089,In_200,In_596);
and U2090 (N_2090,In_893,In_790);
nand U2091 (N_2091,In_603,In_504);
nor U2092 (N_2092,In_87,In_738);
and U2093 (N_2093,In_328,In_909);
or U2094 (N_2094,In_742,In_611);
nand U2095 (N_2095,In_714,In_328);
or U2096 (N_2096,In_86,In_962);
xor U2097 (N_2097,In_811,In_723);
and U2098 (N_2098,In_352,In_772);
or U2099 (N_2099,In_414,In_497);
or U2100 (N_2100,In_619,In_317);
nor U2101 (N_2101,In_17,In_136);
nand U2102 (N_2102,In_723,In_509);
nor U2103 (N_2103,In_910,In_269);
or U2104 (N_2104,In_940,In_199);
or U2105 (N_2105,In_361,In_306);
and U2106 (N_2106,In_10,In_406);
or U2107 (N_2107,In_799,In_512);
and U2108 (N_2108,In_954,In_528);
or U2109 (N_2109,In_951,In_823);
nand U2110 (N_2110,In_334,In_773);
or U2111 (N_2111,In_474,In_533);
nand U2112 (N_2112,In_368,In_235);
nor U2113 (N_2113,In_957,In_746);
nand U2114 (N_2114,In_209,In_682);
or U2115 (N_2115,In_975,In_705);
nand U2116 (N_2116,In_14,In_392);
and U2117 (N_2117,In_822,In_196);
and U2118 (N_2118,In_423,In_323);
or U2119 (N_2119,In_312,In_361);
and U2120 (N_2120,In_929,In_377);
and U2121 (N_2121,In_461,In_804);
or U2122 (N_2122,In_10,In_122);
and U2123 (N_2123,In_206,In_575);
and U2124 (N_2124,In_70,In_677);
nor U2125 (N_2125,In_673,In_270);
or U2126 (N_2126,In_112,In_78);
or U2127 (N_2127,In_964,In_848);
or U2128 (N_2128,In_316,In_470);
and U2129 (N_2129,In_194,In_187);
and U2130 (N_2130,In_398,In_704);
or U2131 (N_2131,In_146,In_29);
nand U2132 (N_2132,In_902,In_719);
and U2133 (N_2133,In_203,In_658);
xnor U2134 (N_2134,In_231,In_944);
nand U2135 (N_2135,In_235,In_422);
nand U2136 (N_2136,In_178,In_274);
or U2137 (N_2137,In_930,In_791);
or U2138 (N_2138,In_426,In_153);
or U2139 (N_2139,In_976,In_183);
nand U2140 (N_2140,In_481,In_189);
or U2141 (N_2141,In_288,In_150);
nand U2142 (N_2142,In_938,In_432);
nand U2143 (N_2143,In_981,In_640);
nor U2144 (N_2144,In_896,In_80);
nand U2145 (N_2145,In_777,In_375);
nor U2146 (N_2146,In_343,In_476);
nand U2147 (N_2147,In_796,In_326);
or U2148 (N_2148,In_28,In_446);
nor U2149 (N_2149,In_264,In_764);
and U2150 (N_2150,In_903,In_180);
nand U2151 (N_2151,In_576,In_222);
nand U2152 (N_2152,In_829,In_778);
nor U2153 (N_2153,In_973,In_618);
and U2154 (N_2154,In_302,In_396);
nor U2155 (N_2155,In_44,In_21);
or U2156 (N_2156,In_872,In_185);
or U2157 (N_2157,In_628,In_426);
nor U2158 (N_2158,In_317,In_365);
or U2159 (N_2159,In_603,In_734);
nand U2160 (N_2160,In_860,In_218);
or U2161 (N_2161,In_605,In_421);
xnor U2162 (N_2162,In_64,In_93);
nor U2163 (N_2163,In_522,In_19);
nor U2164 (N_2164,In_15,In_594);
nand U2165 (N_2165,In_203,In_115);
or U2166 (N_2166,In_405,In_334);
or U2167 (N_2167,In_984,In_951);
nor U2168 (N_2168,In_143,In_578);
or U2169 (N_2169,In_295,In_831);
nor U2170 (N_2170,In_702,In_117);
nand U2171 (N_2171,In_849,In_330);
and U2172 (N_2172,In_530,In_191);
nor U2173 (N_2173,In_217,In_338);
and U2174 (N_2174,In_783,In_262);
nand U2175 (N_2175,In_665,In_995);
nor U2176 (N_2176,In_830,In_236);
or U2177 (N_2177,In_861,In_989);
nor U2178 (N_2178,In_218,In_917);
or U2179 (N_2179,In_943,In_743);
and U2180 (N_2180,In_559,In_768);
nand U2181 (N_2181,In_355,In_874);
nand U2182 (N_2182,In_75,In_225);
nor U2183 (N_2183,In_47,In_733);
nand U2184 (N_2184,In_254,In_730);
or U2185 (N_2185,In_321,In_595);
and U2186 (N_2186,In_777,In_857);
nand U2187 (N_2187,In_752,In_601);
and U2188 (N_2188,In_294,In_712);
nand U2189 (N_2189,In_747,In_523);
nor U2190 (N_2190,In_227,In_79);
nand U2191 (N_2191,In_957,In_26);
nand U2192 (N_2192,In_162,In_881);
nand U2193 (N_2193,In_823,In_172);
or U2194 (N_2194,In_956,In_50);
nor U2195 (N_2195,In_411,In_490);
nor U2196 (N_2196,In_817,In_735);
or U2197 (N_2197,In_200,In_665);
and U2198 (N_2198,In_836,In_72);
nor U2199 (N_2199,In_8,In_99);
nand U2200 (N_2200,In_504,In_403);
and U2201 (N_2201,In_169,In_730);
and U2202 (N_2202,In_730,In_869);
nand U2203 (N_2203,In_314,In_414);
or U2204 (N_2204,In_945,In_736);
nor U2205 (N_2205,In_730,In_541);
and U2206 (N_2206,In_711,In_107);
nor U2207 (N_2207,In_388,In_607);
nor U2208 (N_2208,In_386,In_200);
or U2209 (N_2209,In_24,In_313);
nor U2210 (N_2210,In_410,In_973);
nand U2211 (N_2211,In_79,In_786);
nand U2212 (N_2212,In_133,In_210);
and U2213 (N_2213,In_721,In_486);
nand U2214 (N_2214,In_248,In_102);
and U2215 (N_2215,In_182,In_465);
or U2216 (N_2216,In_557,In_768);
nand U2217 (N_2217,In_536,In_693);
nand U2218 (N_2218,In_52,In_179);
nand U2219 (N_2219,In_659,In_138);
and U2220 (N_2220,In_289,In_576);
nor U2221 (N_2221,In_853,In_46);
or U2222 (N_2222,In_956,In_946);
or U2223 (N_2223,In_279,In_407);
nor U2224 (N_2224,In_329,In_856);
and U2225 (N_2225,In_10,In_564);
nand U2226 (N_2226,In_50,In_990);
or U2227 (N_2227,In_402,In_709);
or U2228 (N_2228,In_156,In_371);
and U2229 (N_2229,In_272,In_33);
and U2230 (N_2230,In_681,In_106);
nand U2231 (N_2231,In_366,In_208);
and U2232 (N_2232,In_813,In_499);
and U2233 (N_2233,In_71,In_803);
nor U2234 (N_2234,In_702,In_154);
and U2235 (N_2235,In_503,In_409);
nand U2236 (N_2236,In_395,In_485);
nand U2237 (N_2237,In_361,In_57);
nor U2238 (N_2238,In_66,In_1);
nor U2239 (N_2239,In_548,In_485);
nor U2240 (N_2240,In_372,In_809);
nor U2241 (N_2241,In_145,In_768);
xnor U2242 (N_2242,In_222,In_266);
nand U2243 (N_2243,In_613,In_228);
or U2244 (N_2244,In_455,In_700);
nand U2245 (N_2245,In_780,In_685);
or U2246 (N_2246,In_263,In_689);
and U2247 (N_2247,In_544,In_693);
or U2248 (N_2248,In_803,In_419);
nand U2249 (N_2249,In_16,In_406);
xor U2250 (N_2250,In_143,In_857);
nand U2251 (N_2251,In_582,In_884);
and U2252 (N_2252,In_117,In_556);
nand U2253 (N_2253,In_550,In_89);
nand U2254 (N_2254,In_453,In_238);
and U2255 (N_2255,In_172,In_321);
and U2256 (N_2256,In_885,In_322);
or U2257 (N_2257,In_292,In_151);
or U2258 (N_2258,In_990,In_677);
or U2259 (N_2259,In_670,In_549);
and U2260 (N_2260,In_838,In_564);
xor U2261 (N_2261,In_111,In_462);
nor U2262 (N_2262,In_903,In_907);
and U2263 (N_2263,In_267,In_304);
or U2264 (N_2264,In_651,In_896);
or U2265 (N_2265,In_638,In_475);
or U2266 (N_2266,In_348,In_493);
nor U2267 (N_2267,In_247,In_626);
and U2268 (N_2268,In_945,In_438);
and U2269 (N_2269,In_654,In_451);
or U2270 (N_2270,In_993,In_736);
or U2271 (N_2271,In_436,In_702);
and U2272 (N_2272,In_752,In_850);
nor U2273 (N_2273,In_960,In_483);
nand U2274 (N_2274,In_747,In_907);
and U2275 (N_2275,In_730,In_578);
or U2276 (N_2276,In_99,In_250);
or U2277 (N_2277,In_964,In_758);
or U2278 (N_2278,In_550,In_108);
and U2279 (N_2279,In_992,In_311);
and U2280 (N_2280,In_713,In_627);
and U2281 (N_2281,In_311,In_875);
or U2282 (N_2282,In_768,In_122);
nor U2283 (N_2283,In_180,In_310);
and U2284 (N_2284,In_197,In_17);
or U2285 (N_2285,In_951,In_859);
nor U2286 (N_2286,In_991,In_541);
or U2287 (N_2287,In_652,In_384);
and U2288 (N_2288,In_294,In_391);
and U2289 (N_2289,In_279,In_825);
nand U2290 (N_2290,In_884,In_9);
or U2291 (N_2291,In_536,In_61);
and U2292 (N_2292,In_20,In_39);
and U2293 (N_2293,In_760,In_269);
nand U2294 (N_2294,In_569,In_583);
nand U2295 (N_2295,In_739,In_760);
nor U2296 (N_2296,In_343,In_236);
nor U2297 (N_2297,In_687,In_850);
nand U2298 (N_2298,In_294,In_795);
nor U2299 (N_2299,In_210,In_58);
or U2300 (N_2300,In_787,In_144);
and U2301 (N_2301,In_59,In_345);
nor U2302 (N_2302,In_494,In_892);
or U2303 (N_2303,In_354,In_102);
and U2304 (N_2304,In_985,In_473);
and U2305 (N_2305,In_786,In_815);
and U2306 (N_2306,In_560,In_13);
nand U2307 (N_2307,In_261,In_251);
or U2308 (N_2308,In_71,In_573);
and U2309 (N_2309,In_870,In_669);
and U2310 (N_2310,In_985,In_203);
and U2311 (N_2311,In_649,In_670);
nor U2312 (N_2312,In_24,In_54);
xnor U2313 (N_2313,In_88,In_632);
nand U2314 (N_2314,In_756,In_630);
nand U2315 (N_2315,In_442,In_948);
nor U2316 (N_2316,In_900,In_629);
nor U2317 (N_2317,In_488,In_39);
or U2318 (N_2318,In_502,In_595);
nor U2319 (N_2319,In_574,In_871);
or U2320 (N_2320,In_782,In_645);
nand U2321 (N_2321,In_389,In_915);
and U2322 (N_2322,In_597,In_878);
and U2323 (N_2323,In_892,In_876);
and U2324 (N_2324,In_861,In_975);
or U2325 (N_2325,In_217,In_733);
and U2326 (N_2326,In_994,In_152);
or U2327 (N_2327,In_307,In_164);
nor U2328 (N_2328,In_961,In_190);
and U2329 (N_2329,In_319,In_994);
nand U2330 (N_2330,In_237,In_474);
and U2331 (N_2331,In_133,In_392);
or U2332 (N_2332,In_397,In_704);
and U2333 (N_2333,In_358,In_522);
nor U2334 (N_2334,In_331,In_468);
and U2335 (N_2335,In_730,In_479);
nand U2336 (N_2336,In_881,In_971);
nand U2337 (N_2337,In_713,In_577);
nor U2338 (N_2338,In_233,In_15);
and U2339 (N_2339,In_560,In_666);
or U2340 (N_2340,In_463,In_951);
nand U2341 (N_2341,In_81,In_517);
and U2342 (N_2342,In_184,In_688);
or U2343 (N_2343,In_410,In_904);
or U2344 (N_2344,In_716,In_89);
and U2345 (N_2345,In_475,In_87);
or U2346 (N_2346,In_965,In_153);
nor U2347 (N_2347,In_57,In_403);
nand U2348 (N_2348,In_367,In_47);
nand U2349 (N_2349,In_742,In_145);
nor U2350 (N_2350,In_773,In_502);
nor U2351 (N_2351,In_781,In_737);
nor U2352 (N_2352,In_933,In_45);
and U2353 (N_2353,In_65,In_655);
nand U2354 (N_2354,In_100,In_974);
and U2355 (N_2355,In_501,In_753);
nand U2356 (N_2356,In_258,In_578);
nand U2357 (N_2357,In_479,In_71);
or U2358 (N_2358,In_950,In_1);
nor U2359 (N_2359,In_424,In_423);
nor U2360 (N_2360,In_707,In_719);
nor U2361 (N_2361,In_33,In_933);
and U2362 (N_2362,In_517,In_541);
nand U2363 (N_2363,In_11,In_360);
and U2364 (N_2364,In_855,In_983);
and U2365 (N_2365,In_877,In_785);
nor U2366 (N_2366,In_408,In_199);
nor U2367 (N_2367,In_583,In_937);
nor U2368 (N_2368,In_323,In_476);
nor U2369 (N_2369,In_537,In_260);
and U2370 (N_2370,In_708,In_275);
and U2371 (N_2371,In_818,In_57);
xnor U2372 (N_2372,In_894,In_13);
nor U2373 (N_2373,In_668,In_845);
and U2374 (N_2374,In_721,In_912);
nor U2375 (N_2375,In_585,In_313);
nor U2376 (N_2376,In_725,In_652);
nand U2377 (N_2377,In_270,In_296);
nand U2378 (N_2378,In_351,In_32);
and U2379 (N_2379,In_967,In_124);
nand U2380 (N_2380,In_915,In_326);
nor U2381 (N_2381,In_528,In_24);
nand U2382 (N_2382,In_169,In_181);
nor U2383 (N_2383,In_133,In_987);
nor U2384 (N_2384,In_244,In_959);
or U2385 (N_2385,In_95,In_111);
nor U2386 (N_2386,In_331,In_891);
nor U2387 (N_2387,In_637,In_529);
nor U2388 (N_2388,In_358,In_436);
and U2389 (N_2389,In_750,In_857);
nand U2390 (N_2390,In_498,In_479);
nand U2391 (N_2391,In_801,In_150);
nand U2392 (N_2392,In_137,In_614);
and U2393 (N_2393,In_383,In_980);
or U2394 (N_2394,In_767,In_947);
or U2395 (N_2395,In_589,In_160);
nand U2396 (N_2396,In_624,In_520);
and U2397 (N_2397,In_387,In_658);
nor U2398 (N_2398,In_293,In_796);
nor U2399 (N_2399,In_541,In_250);
or U2400 (N_2400,In_508,In_415);
or U2401 (N_2401,In_618,In_272);
nand U2402 (N_2402,In_642,In_594);
and U2403 (N_2403,In_875,In_647);
nor U2404 (N_2404,In_218,In_295);
or U2405 (N_2405,In_785,In_407);
nand U2406 (N_2406,In_15,In_678);
and U2407 (N_2407,In_245,In_861);
nor U2408 (N_2408,In_902,In_899);
nor U2409 (N_2409,In_505,In_556);
and U2410 (N_2410,In_985,In_852);
and U2411 (N_2411,In_617,In_86);
and U2412 (N_2412,In_977,In_606);
xor U2413 (N_2413,In_33,In_208);
nor U2414 (N_2414,In_299,In_858);
and U2415 (N_2415,In_959,In_575);
nand U2416 (N_2416,In_412,In_853);
nand U2417 (N_2417,In_935,In_714);
and U2418 (N_2418,In_903,In_708);
and U2419 (N_2419,In_121,In_651);
and U2420 (N_2420,In_610,In_511);
nand U2421 (N_2421,In_544,In_359);
or U2422 (N_2422,In_948,In_982);
or U2423 (N_2423,In_300,In_569);
or U2424 (N_2424,In_97,In_420);
and U2425 (N_2425,In_836,In_165);
or U2426 (N_2426,In_225,In_346);
or U2427 (N_2427,In_276,In_689);
nand U2428 (N_2428,In_472,In_524);
nor U2429 (N_2429,In_216,In_910);
nor U2430 (N_2430,In_861,In_880);
nor U2431 (N_2431,In_372,In_517);
nand U2432 (N_2432,In_598,In_478);
or U2433 (N_2433,In_521,In_90);
nand U2434 (N_2434,In_699,In_432);
and U2435 (N_2435,In_445,In_325);
and U2436 (N_2436,In_90,In_998);
or U2437 (N_2437,In_504,In_375);
nor U2438 (N_2438,In_466,In_150);
nand U2439 (N_2439,In_690,In_507);
nor U2440 (N_2440,In_923,In_776);
xor U2441 (N_2441,In_593,In_819);
nand U2442 (N_2442,In_490,In_330);
and U2443 (N_2443,In_395,In_114);
nor U2444 (N_2444,In_39,In_661);
and U2445 (N_2445,In_304,In_504);
nand U2446 (N_2446,In_243,In_4);
nand U2447 (N_2447,In_821,In_190);
or U2448 (N_2448,In_970,In_893);
or U2449 (N_2449,In_170,In_307);
or U2450 (N_2450,In_796,In_283);
nand U2451 (N_2451,In_165,In_83);
or U2452 (N_2452,In_329,In_698);
or U2453 (N_2453,In_166,In_402);
and U2454 (N_2454,In_98,In_903);
and U2455 (N_2455,In_135,In_115);
nor U2456 (N_2456,In_680,In_138);
nand U2457 (N_2457,In_422,In_353);
nor U2458 (N_2458,In_157,In_437);
and U2459 (N_2459,In_490,In_227);
and U2460 (N_2460,In_592,In_651);
nand U2461 (N_2461,In_5,In_9);
nor U2462 (N_2462,In_188,In_427);
and U2463 (N_2463,In_652,In_948);
nand U2464 (N_2464,In_258,In_150);
and U2465 (N_2465,In_104,In_409);
nor U2466 (N_2466,In_903,In_393);
nand U2467 (N_2467,In_142,In_191);
or U2468 (N_2468,In_571,In_213);
or U2469 (N_2469,In_291,In_521);
nor U2470 (N_2470,In_411,In_200);
and U2471 (N_2471,In_603,In_587);
and U2472 (N_2472,In_130,In_502);
nor U2473 (N_2473,In_539,In_362);
and U2474 (N_2474,In_319,In_795);
and U2475 (N_2475,In_327,In_7);
nor U2476 (N_2476,In_774,In_128);
and U2477 (N_2477,In_123,In_931);
nand U2478 (N_2478,In_65,In_864);
or U2479 (N_2479,In_248,In_888);
nand U2480 (N_2480,In_103,In_710);
nand U2481 (N_2481,In_262,In_245);
or U2482 (N_2482,In_61,In_624);
xor U2483 (N_2483,In_590,In_163);
and U2484 (N_2484,In_983,In_609);
nor U2485 (N_2485,In_227,In_508);
nor U2486 (N_2486,In_711,In_112);
or U2487 (N_2487,In_159,In_151);
and U2488 (N_2488,In_79,In_559);
nand U2489 (N_2489,In_366,In_818);
nor U2490 (N_2490,In_964,In_879);
and U2491 (N_2491,In_780,In_154);
nor U2492 (N_2492,In_580,In_730);
nand U2493 (N_2493,In_231,In_831);
nor U2494 (N_2494,In_478,In_312);
nand U2495 (N_2495,In_377,In_15);
nand U2496 (N_2496,In_657,In_98);
and U2497 (N_2497,In_228,In_81);
and U2498 (N_2498,In_245,In_24);
or U2499 (N_2499,In_233,In_152);
or U2500 (N_2500,N_458,N_1892);
nand U2501 (N_2501,N_2292,N_1020);
nor U2502 (N_2502,N_1001,N_2381);
or U2503 (N_2503,N_1548,N_325);
nor U2504 (N_2504,N_1799,N_1201);
or U2505 (N_2505,N_2445,N_1278);
nand U2506 (N_2506,N_1304,N_2173);
nand U2507 (N_2507,N_1835,N_454);
or U2508 (N_2508,N_38,N_2464);
and U2509 (N_2509,N_736,N_1557);
or U2510 (N_2510,N_149,N_1767);
or U2511 (N_2511,N_1568,N_1874);
nor U2512 (N_2512,N_2247,N_2108);
or U2513 (N_2513,N_250,N_1083);
or U2514 (N_2514,N_1421,N_1919);
and U2515 (N_2515,N_2291,N_771);
nand U2516 (N_2516,N_2006,N_1039);
and U2517 (N_2517,N_1402,N_1348);
nor U2518 (N_2518,N_1978,N_2094);
nand U2519 (N_2519,N_2142,N_116);
nor U2520 (N_2520,N_714,N_2446);
or U2521 (N_2521,N_2125,N_2440);
and U2522 (N_2522,N_31,N_1409);
nor U2523 (N_2523,N_472,N_777);
nand U2524 (N_2524,N_1647,N_977);
nor U2525 (N_2525,N_1173,N_1111);
nor U2526 (N_2526,N_17,N_1938);
nor U2527 (N_2527,N_547,N_1556);
nand U2528 (N_2528,N_1109,N_194);
nand U2529 (N_2529,N_1240,N_578);
and U2530 (N_2530,N_2060,N_326);
and U2531 (N_2531,N_536,N_610);
nand U2532 (N_2532,N_2074,N_1853);
nand U2533 (N_2533,N_1117,N_752);
nor U2534 (N_2534,N_2226,N_385);
nor U2535 (N_2535,N_783,N_373);
and U2536 (N_2536,N_798,N_950);
nor U2537 (N_2537,N_2050,N_350);
or U2538 (N_2538,N_2063,N_543);
nor U2539 (N_2539,N_1762,N_1666);
nor U2540 (N_2540,N_986,N_2251);
nand U2541 (N_2541,N_556,N_2218);
and U2542 (N_2542,N_1145,N_1144);
nor U2543 (N_2543,N_344,N_1552);
nand U2544 (N_2544,N_1852,N_2105);
and U2545 (N_2545,N_1953,N_683);
or U2546 (N_2546,N_2237,N_2376);
or U2547 (N_2547,N_2229,N_2433);
nor U2548 (N_2548,N_1102,N_744);
nand U2549 (N_2549,N_1178,N_708);
or U2550 (N_2550,N_530,N_1975);
and U2551 (N_2551,N_1417,N_1336);
nor U2552 (N_2552,N_2203,N_2438);
or U2553 (N_2553,N_1549,N_1808);
or U2554 (N_2554,N_1828,N_1299);
nor U2555 (N_2555,N_2136,N_1207);
or U2556 (N_2556,N_1352,N_706);
xor U2557 (N_2557,N_844,N_416);
or U2558 (N_2558,N_979,N_2283);
nand U2559 (N_2559,N_1035,N_258);
or U2560 (N_2560,N_1256,N_658);
nand U2561 (N_2561,N_606,N_1472);
or U2562 (N_2562,N_2472,N_1063);
nor U2563 (N_2563,N_473,N_247);
xor U2564 (N_2564,N_1644,N_2047);
and U2565 (N_2565,N_352,N_424);
nor U2566 (N_2566,N_949,N_2099);
and U2567 (N_2567,N_308,N_813);
xnor U2568 (N_2568,N_1079,N_967);
and U2569 (N_2569,N_877,N_1106);
nor U2570 (N_2570,N_1213,N_1915);
or U2571 (N_2571,N_668,N_689);
nor U2572 (N_2572,N_1135,N_985);
nand U2573 (N_2573,N_329,N_457);
nor U2574 (N_2574,N_1362,N_1765);
nor U2575 (N_2575,N_1452,N_1846);
or U2576 (N_2576,N_1252,N_1338);
and U2577 (N_2577,N_220,N_947);
nand U2578 (N_2578,N_1040,N_829);
nor U2579 (N_2579,N_1608,N_1047);
nor U2580 (N_2580,N_16,N_1021);
nand U2581 (N_2581,N_188,N_167);
or U2582 (N_2582,N_522,N_943);
nand U2583 (N_2583,N_427,N_1528);
nand U2584 (N_2584,N_927,N_317);
nor U2585 (N_2585,N_1725,N_918);
or U2586 (N_2586,N_93,N_2430);
and U2587 (N_2587,N_1501,N_1006);
nor U2588 (N_2588,N_973,N_501);
or U2589 (N_2589,N_1776,N_2068);
or U2590 (N_2590,N_430,N_770);
and U2591 (N_2591,N_1378,N_371);
or U2592 (N_2592,N_1507,N_896);
nor U2593 (N_2593,N_814,N_591);
nand U2594 (N_2594,N_1536,N_931);
or U2595 (N_2595,N_1890,N_564);
or U2596 (N_2596,N_1343,N_795);
nor U2597 (N_2597,N_1208,N_2289);
nor U2598 (N_2598,N_348,N_2332);
nand U2599 (N_2599,N_1830,N_1763);
and U2600 (N_2600,N_1984,N_551);
and U2601 (N_2601,N_1255,N_2185);
nand U2602 (N_2602,N_2081,N_2129);
and U2603 (N_2603,N_1330,N_1425);
or U2604 (N_2604,N_255,N_1972);
nor U2605 (N_2605,N_872,N_225);
or U2606 (N_2606,N_651,N_954);
nor U2607 (N_2607,N_2205,N_2184);
nor U2608 (N_2608,N_41,N_2124);
and U2609 (N_2609,N_769,N_1420);
nor U2610 (N_2610,N_1573,N_890);
nand U2611 (N_2611,N_2034,N_1467);
nand U2612 (N_2612,N_202,N_634);
and U2613 (N_2613,N_479,N_1658);
or U2614 (N_2614,N_1239,N_2336);
and U2615 (N_2615,N_552,N_842);
nand U2616 (N_2616,N_2313,N_1926);
nor U2617 (N_2617,N_2286,N_1395);
and U2618 (N_2618,N_1317,N_2007);
nand U2619 (N_2619,N_171,N_2409);
or U2620 (N_2620,N_1462,N_1685);
and U2621 (N_2621,N_1679,N_2232);
nor U2622 (N_2622,N_2491,N_414);
and U2623 (N_2623,N_1199,N_1586);
nand U2624 (N_2624,N_1993,N_1577);
and U2625 (N_2625,N_987,N_874);
and U2626 (N_2626,N_153,N_1719);
nand U2627 (N_2627,N_42,N_1598);
or U2628 (N_2628,N_2273,N_135);
or U2629 (N_2629,N_1313,N_1324);
nand U2630 (N_2630,N_1061,N_1641);
and U2631 (N_2631,N_924,N_2059);
and U2632 (N_2632,N_2150,N_1443);
nand U2633 (N_2633,N_711,N_2486);
and U2634 (N_2634,N_345,N_2194);
xor U2635 (N_2635,N_735,N_1792);
and U2636 (N_2636,N_2039,N_299);
and U2637 (N_2637,N_1314,N_1119);
and U2638 (N_2638,N_83,N_1414);
or U2639 (N_2639,N_1800,N_399);
or U2640 (N_2640,N_2485,N_2394);
nor U2641 (N_2641,N_1718,N_252);
nand U2642 (N_2642,N_1560,N_2419);
nand U2643 (N_2643,N_1244,N_2387);
and U2644 (N_2644,N_2272,N_542);
nand U2645 (N_2645,N_2462,N_1990);
nor U2646 (N_2646,N_2493,N_411);
or U2647 (N_2647,N_984,N_1454);
and U2648 (N_2648,N_2127,N_1387);
nor U2649 (N_2649,N_1151,N_2104);
or U2650 (N_2650,N_1939,N_616);
and U2651 (N_2651,N_1910,N_846);
nor U2652 (N_2652,N_2244,N_2155);
or U2653 (N_2653,N_1758,N_2449);
and U2654 (N_2654,N_1356,N_1216);
nand U2655 (N_2655,N_466,N_205);
nor U2656 (N_2656,N_1126,N_2294);
xor U2657 (N_2657,N_2069,N_923);
nand U2658 (N_2658,N_1347,N_2174);
nor U2659 (N_2659,N_781,N_2078);
or U2660 (N_2660,N_751,N_277);
or U2661 (N_2661,N_792,N_1519);
nor U2662 (N_2662,N_817,N_1947);
or U2663 (N_2663,N_1113,N_7);
or U2664 (N_2664,N_2023,N_1535);
xnor U2665 (N_2665,N_242,N_1029);
and U2666 (N_2666,N_174,N_2466);
or U2667 (N_2667,N_510,N_187);
or U2668 (N_2668,N_1675,N_1388);
or U2669 (N_2669,N_1322,N_2117);
and U2670 (N_2670,N_1152,N_1226);
and U2671 (N_2671,N_851,N_1477);
nand U2672 (N_2672,N_2231,N_160);
or U2673 (N_2673,N_239,N_2391);
or U2674 (N_2674,N_617,N_1385);
nand U2675 (N_2675,N_1863,N_2181);
nor U2676 (N_2676,N_132,N_2100);
nand U2677 (N_2677,N_138,N_235);
nor U2678 (N_2678,N_1961,N_1249);
and U2679 (N_2679,N_2178,N_2320);
nor U2680 (N_2680,N_1637,N_1115);
and U2681 (N_2681,N_67,N_396);
and U2682 (N_2682,N_811,N_1968);
nor U2683 (N_2683,N_2022,N_2013);
nand U2684 (N_2684,N_869,N_797);
nand U2685 (N_2685,N_2368,N_2358);
or U2686 (N_2686,N_793,N_2159);
xor U2687 (N_2687,N_1609,N_1293);
and U2688 (N_2688,N_1617,N_1078);
and U2689 (N_2689,N_441,N_1907);
nand U2690 (N_2690,N_749,N_1790);
nand U2691 (N_2691,N_1855,N_1948);
and U2692 (N_2692,N_133,N_213);
nand U2693 (N_2693,N_2441,N_2329);
and U2694 (N_2694,N_2204,N_624);
nand U2695 (N_2695,N_1985,N_1341);
and U2696 (N_2696,N_1309,N_840);
and U2697 (N_2697,N_2379,N_1936);
or U2698 (N_2698,N_1405,N_854);
nor U2699 (N_2699,N_1950,N_2221);
or U2700 (N_2700,N_1665,N_337);
and U2701 (N_2701,N_1381,N_621);
and U2702 (N_2702,N_1994,N_1429);
nor U2703 (N_2703,N_1529,N_2041);
nand U2704 (N_2704,N_2024,N_568);
nor U2705 (N_2705,N_692,N_1946);
or U2706 (N_2706,N_1735,N_1991);
or U2707 (N_2707,N_9,N_59);
nor U2708 (N_2708,N_2361,N_876);
or U2709 (N_2709,N_1143,N_268);
nor U2710 (N_2710,N_521,N_524);
or U2711 (N_2711,N_1349,N_1060);
or U2712 (N_2712,N_1784,N_1533);
or U2713 (N_2713,N_1812,N_594);
and U2714 (N_2714,N_131,N_1311);
or U2715 (N_2715,N_1704,N_2439);
nor U2716 (N_2716,N_387,N_1455);
nor U2717 (N_2717,N_110,N_2064);
or U2718 (N_2718,N_477,N_1399);
nand U2719 (N_2719,N_1866,N_1242);
and U2720 (N_2720,N_143,N_2260);
nand U2721 (N_2721,N_32,N_1840);
or U2722 (N_2722,N_538,N_700);
or U2723 (N_2723,N_701,N_628);
nand U2724 (N_2724,N_1905,N_2224);
nand U2725 (N_2725,N_1380,N_483);
and U2726 (N_2726,N_857,N_703);
nor U2727 (N_2727,N_2375,N_511);
and U2728 (N_2728,N_2249,N_1510);
and U2729 (N_2729,N_2325,N_1218);
nand U2730 (N_2730,N_1614,N_750);
nand U2731 (N_2731,N_847,N_1632);
nand U2732 (N_2732,N_1464,N_1486);
nand U2733 (N_2733,N_2279,N_117);
nand U2734 (N_2734,N_264,N_1008);
and U2735 (N_2735,N_1913,N_2384);
nor U2736 (N_2736,N_1657,N_733);
nor U2737 (N_2737,N_2367,N_1674);
nand U2738 (N_2738,N_2036,N_2119);
or U2739 (N_2739,N_1241,N_570);
or U2740 (N_2740,N_801,N_359);
or U2741 (N_2741,N_1284,N_1764);
nor U2742 (N_2742,N_917,N_1629);
nor U2743 (N_2743,N_2451,N_356);
or U2744 (N_2744,N_388,N_1332);
nor U2745 (N_2745,N_1634,N_163);
and U2746 (N_2746,N_741,N_429);
or U2747 (N_2747,N_2479,N_77);
nor U2748 (N_2748,N_2167,N_439);
and U2749 (N_2749,N_1396,N_1316);
and U2750 (N_2750,N_1271,N_2072);
nor U2751 (N_2751,N_1407,N_2355);
or U2752 (N_2752,N_773,N_837);
or U2753 (N_2753,N_378,N_1945);
nand U2754 (N_2754,N_335,N_2457);
nor U2755 (N_2755,N_1653,N_1358);
nor U2756 (N_2756,N_1748,N_1831);
and U2757 (N_2757,N_1128,N_1859);
nand U2758 (N_2758,N_2305,N_963);
and U2759 (N_2759,N_2045,N_833);
nand U2760 (N_2760,N_922,N_118);
or U2761 (N_2761,N_1091,N_231);
nor U2762 (N_2762,N_978,N_261);
nand U2763 (N_2763,N_169,N_630);
nand U2764 (N_2764,N_1937,N_2046);
nor U2765 (N_2765,N_2234,N_107);
or U2766 (N_2766,N_637,N_464);
nor U2767 (N_2767,N_2453,N_573);
nor U2768 (N_2768,N_1605,N_1285);
nand U2769 (N_2769,N_721,N_2400);
or U2770 (N_2770,N_1518,N_760);
nand U2771 (N_2771,N_64,N_690);
and U2772 (N_2772,N_1400,N_2000);
or U2773 (N_2773,N_2153,N_1900);
and U2774 (N_2774,N_787,N_1565);
and U2775 (N_2775,N_2357,N_2135);
nand U2776 (N_2776,N_830,N_1066);
nand U2777 (N_2777,N_15,N_81);
or U2778 (N_2778,N_697,N_2437);
nand U2779 (N_2779,N_2423,N_1814);
nor U2780 (N_2780,N_391,N_1401);
nor U2781 (N_2781,N_285,N_73);
or U2782 (N_2782,N_1896,N_318);
and U2783 (N_2783,N_320,N_957);
or U2784 (N_2784,N_1346,N_1248);
or U2785 (N_2785,N_407,N_413);
nand U2786 (N_2786,N_1458,N_2349);
xor U2787 (N_2787,N_1524,N_2442);
nand U2788 (N_2788,N_1424,N_1023);
and U2789 (N_2789,N_2406,N_2053);
nand U2790 (N_2790,N_1716,N_1333);
nand U2791 (N_2791,N_180,N_1099);
nor U2792 (N_2792,N_1430,N_1832);
and U2793 (N_2793,N_301,N_298);
and U2794 (N_2794,N_1011,N_204);
nand U2795 (N_2795,N_1394,N_535);
and U2796 (N_2796,N_2311,N_51);
nand U2797 (N_2797,N_1841,N_2404);
or U2798 (N_2798,N_2192,N_362);
nor U2799 (N_2799,N_336,N_1893);
nand U2800 (N_2800,N_450,N_418);
or U2801 (N_2801,N_1253,N_1624);
or U2802 (N_2802,N_2296,N_1941);
nand U2803 (N_2803,N_2304,N_981);
and U2804 (N_2804,N_2315,N_1772);
or U2805 (N_2805,N_2395,N_283);
and U2806 (N_2806,N_340,N_1924);
or U2807 (N_2807,N_1933,N_2350);
nand U2808 (N_2808,N_2342,N_2293);
nand U2809 (N_2809,N_1729,N_461);
or U2810 (N_2810,N_1575,N_372);
nand U2811 (N_2811,N_2147,N_2471);
xor U2812 (N_2812,N_587,N_1042);
nor U2813 (N_2813,N_297,N_1157);
or U2814 (N_2814,N_1465,N_660);
and U2815 (N_2815,N_1137,N_1664);
nand U2816 (N_2816,N_804,N_2463);
and U2817 (N_2817,N_2424,N_363);
or U2818 (N_2818,N_1131,N_1171);
and U2819 (N_2819,N_859,N_295);
or U2820 (N_2820,N_87,N_2415);
xnor U2821 (N_2821,N_181,N_1705);
or U2822 (N_2822,N_748,N_504);
nand U2823 (N_2823,N_1925,N_1268);
or U2824 (N_2824,N_157,N_1476);
or U2825 (N_2825,N_2301,N_904);
nand U2826 (N_2826,N_1667,N_2353);
and U2827 (N_2827,N_1471,N_1555);
nand U2828 (N_2828,N_2323,N_1325);
nor U2829 (N_2829,N_1331,N_357);
nand U2830 (N_2830,N_2360,N_2393);
and U2831 (N_2831,N_236,N_1646);
or U2832 (N_2832,N_1631,N_2211);
or U2833 (N_2833,N_410,N_2475);
nand U2834 (N_2834,N_1908,N_2284);
nor U2835 (N_2835,N_680,N_370);
nor U2836 (N_2836,N_2188,N_1597);
nor U2837 (N_2837,N_1326,N_932);
and U2838 (N_2838,N_810,N_2145);
or U2839 (N_2839,N_1934,N_702);
and U2840 (N_2840,N_2163,N_1923);
nand U2841 (N_2841,N_65,N_1775);
nor U2842 (N_2842,N_892,N_1522);
or U2843 (N_2843,N_1418,N_284);
nor U2844 (N_2844,N_199,N_550);
xor U2845 (N_2845,N_2001,N_866);
nor U2846 (N_2846,N_653,N_1504);
nor U2847 (N_2847,N_129,N_2429);
nand U2848 (N_2848,N_589,N_2008);
and U2849 (N_2849,N_155,N_397);
or U2850 (N_2850,N_1583,N_1283);
nand U2851 (N_2851,N_442,N_1403);
and U2852 (N_2852,N_2262,N_1123);
nor U2853 (N_2853,N_124,N_2465);
nor U2854 (N_2854,N_2175,N_49);
and U2855 (N_2855,N_2425,N_695);
and U2856 (N_2856,N_1426,N_1703);
nor U2857 (N_2857,N_2253,N_1964);
or U2858 (N_2858,N_90,N_838);
nand U2859 (N_2859,N_1659,N_240);
nor U2860 (N_2860,N_1466,N_47);
and U2861 (N_2861,N_2456,N_1164);
and U2862 (N_2862,N_1599,N_759);
and U2863 (N_2863,N_1191,N_2373);
or U2864 (N_2864,N_691,N_909);
and U2865 (N_2865,N_2374,N_1876);
nor U2866 (N_2866,N_22,N_1543);
xnor U2867 (N_2867,N_1076,N_2151);
and U2868 (N_2868,N_1980,N_1138);
and U2869 (N_2869,N_926,N_2132);
nand U2870 (N_2870,N_2228,N_279);
and U2871 (N_2871,N_2003,N_2265);
nand U2872 (N_2872,N_878,N_92);
and U2873 (N_2873,N_2019,N_2206);
or U2874 (N_2874,N_894,N_1177);
and U2875 (N_2875,N_2454,N_1158);
nor U2876 (N_2876,N_1186,N_1788);
nand U2877 (N_2877,N_1232,N_426);
nor U2878 (N_2878,N_1613,N_1340);
xnor U2879 (N_2879,N_1377,N_2280);
and U2880 (N_2880,N_588,N_209);
nor U2881 (N_2881,N_982,N_103);
nand U2882 (N_2882,N_1247,N_470);
and U2883 (N_2883,N_1379,N_423);
and U2884 (N_2884,N_48,N_1072);
nand U2885 (N_2885,N_1959,N_1234);
or U2886 (N_2886,N_273,N_1848);
and U2887 (N_2887,N_217,N_1492);
or U2888 (N_2888,N_1965,N_212);
and U2889 (N_2889,N_2410,N_1306);
nor U2890 (N_2890,N_1392,N_2141);
nor U2891 (N_2891,N_2048,N_1404);
and U2892 (N_2892,N_2295,N_835);
nor U2893 (N_2893,N_78,N_1438);
or U2894 (N_2894,N_498,N_2263);
nor U2895 (N_2895,N_1431,N_1798);
or U2896 (N_2896,N_1497,N_351);
nor U2897 (N_2897,N_971,N_1988);
nor U2898 (N_2898,N_34,N_1711);
or U2899 (N_2899,N_2213,N_2207);
nand U2900 (N_2900,N_1744,N_696);
and U2901 (N_2901,N_99,N_1879);
or U2902 (N_2902,N_1585,N_1049);
or U2903 (N_2903,N_1981,N_780);
xor U2904 (N_2904,N_1521,N_1806);
nor U2905 (N_2905,N_481,N_2354);
and U2906 (N_2906,N_2436,N_1470);
nand U2907 (N_2907,N_1491,N_2252);
or U2908 (N_2908,N_929,N_2364);
and U2909 (N_2909,N_1563,N_148);
xor U2910 (N_2910,N_1633,N_1889);
and U2911 (N_2911,N_1734,N_227);
or U2912 (N_2912,N_165,N_1289);
nand U2913 (N_2913,N_743,N_1364);
or U2914 (N_2914,N_1645,N_2321);
and U2915 (N_2915,N_2474,N_559);
or U2916 (N_2916,N_767,N_33);
nor U2917 (N_2917,N_1733,N_1095);
or U2918 (N_2918,N_2026,N_1805);
nand U2919 (N_2919,N_2487,N_919);
or U2920 (N_2920,N_1165,N_253);
or U2921 (N_2921,N_600,N_302);
and U2922 (N_2922,N_1662,N_1016);
and U2923 (N_2923,N_74,N_224);
nor U2924 (N_2924,N_1822,N_1087);
or U2925 (N_2925,N_1742,N_1129);
nand U2926 (N_2926,N_1139,N_910);
nand U2927 (N_2927,N_2341,N_647);
or U2928 (N_2928,N_1150,N_1355);
nand U2929 (N_2929,N_1259,N_282);
or U2930 (N_2930,N_1554,N_666);
and U2931 (N_2931,N_1147,N_1391);
or U2932 (N_2932,N_1816,N_1625);
nand U2933 (N_2933,N_1279,N_393);
nor U2934 (N_2934,N_126,N_826);
or U2935 (N_2935,N_1044,N_1930);
xnor U2936 (N_2936,N_1081,N_900);
and U2937 (N_2937,N_2222,N_2326);
nand U2938 (N_2938,N_1018,N_434);
or U2939 (N_2939,N_1786,N_2484);
nand U2940 (N_2940,N_1678,N_2062);
nand U2941 (N_2941,N_360,N_1434);
and U2942 (N_2942,N_1727,N_289);
and U2943 (N_2943,N_2219,N_88);
xor U2944 (N_2944,N_1071,N_377);
or U2945 (N_2945,N_1690,N_2271);
or U2946 (N_2946,N_2044,N_1161);
nor U2947 (N_2947,N_1844,N_2306);
and U2948 (N_2948,N_1251,N_2372);
and U2949 (N_2949,N_1415,N_1702);
nor U2950 (N_2950,N_349,N_1101);
nand U2951 (N_2951,N_1484,N_1683);
nor U2952 (N_2952,N_1260,N_365);
and U2953 (N_2953,N_1789,N_1615);
or U2954 (N_2954,N_774,N_561);
nor U2955 (N_2955,N_1749,N_2233);
and U2956 (N_2956,N_2385,N_2071);
and U2957 (N_2957,N_305,N_2040);
or U2958 (N_2958,N_2298,N_512);
nor U2959 (N_2959,N_2243,N_718);
nand U2960 (N_2960,N_796,N_822);
nor U2961 (N_2961,N_1211,N_1570);
nand U2962 (N_2962,N_2176,N_885);
nor U2963 (N_2963,N_2343,N_2431);
xor U2964 (N_2964,N_2149,N_1944);
nand U2965 (N_2965,N_531,N_1196);
nor U2966 (N_2966,N_1530,N_1303);
or U2967 (N_2967,N_1747,N_593);
and U2968 (N_2968,N_141,N_554);
nand U2969 (N_2969,N_1759,N_1982);
or U2970 (N_2970,N_316,N_4);
xor U2971 (N_2971,N_715,N_1618);
nor U2972 (N_2972,N_2066,N_8);
nand U2973 (N_2973,N_2093,N_852);
or U2974 (N_2974,N_2427,N_281);
nand U2975 (N_2975,N_1098,N_952);
or U2976 (N_2976,N_489,N_2356);
and U2977 (N_2977,N_1757,N_1694);
xnor U2978 (N_2978,N_1114,N_2112);
or U2979 (N_2979,N_1538,N_25);
nor U2980 (N_2980,N_361,N_791);
or U2981 (N_2981,N_128,N_462);
nor U2982 (N_2982,N_908,N_1928);
nand U2983 (N_2983,N_193,N_2086);
or U2984 (N_2984,N_1136,N_1801);
nor U2985 (N_2985,N_933,N_1033);
and U2986 (N_2986,N_1979,N_836);
nor U2987 (N_2987,N_386,N_1263);
nand U2988 (N_2988,N_1811,N_884);
or U2989 (N_2989,N_82,N_1302);
nand U2990 (N_2990,N_1621,N_10);
nor U2991 (N_2991,N_207,N_580);
and U2992 (N_2992,N_762,N_1180);
nor U2993 (N_2993,N_571,N_907);
nor U2994 (N_2994,N_2158,N_913);
nor U2995 (N_2995,N_2146,N_2309);
nor U2996 (N_2996,N_819,N_1093);
or U2997 (N_2997,N_1670,N_1483);
nand U2998 (N_2998,N_596,N_215);
or U2999 (N_2999,N_1881,N_786);
and U3000 (N_3000,N_2370,N_998);
and U3001 (N_3001,N_259,N_2106);
nand U3002 (N_3002,N_768,N_1235);
and U3003 (N_3003,N_2399,N_146);
and U3004 (N_3004,N_860,N_2397);
and U3005 (N_3005,N_1185,N_256);
nand U3006 (N_3006,N_784,N_1771);
nand U3007 (N_3007,N_68,N_27);
or U3008 (N_3008,N_323,N_379);
nor U3009 (N_3009,N_1579,N_1870);
or U3010 (N_3010,N_1294,N_1869);
nand U3011 (N_3011,N_421,N_1059);
nor U3012 (N_3012,N_1473,N_137);
nand U3013 (N_3013,N_1967,N_970);
or U3014 (N_3014,N_1793,N_641);
nor U3015 (N_3015,N_684,N_2435);
nand U3016 (N_3016,N_1198,N_662);
or U3017 (N_3017,N_485,N_725);
nand U3018 (N_3018,N_1661,N_1300);
nor U3019 (N_3019,N_1397,N_2168);
nor U3020 (N_3020,N_803,N_1693);
or U3021 (N_3021,N_1444,N_368);
or U3022 (N_3022,N_848,N_287);
or U3023 (N_3023,N_1227,N_2411);
nor U3024 (N_3024,N_106,N_1656);
nor U3025 (N_3025,N_1110,N_1532);
nor U3026 (N_3026,N_2010,N_1969);
nand U3027 (N_3027,N_1709,N_2092);
and U3028 (N_3028,N_91,N_1456);
or U3029 (N_3029,N_76,N_23);
nor U3030 (N_3030,N_1236,N_1103);
nand U3031 (N_3031,N_1836,N_1373);
or U3032 (N_3032,N_881,N_1361);
or U3033 (N_3033,N_1527,N_1499);
nand U3034 (N_3034,N_1043,N_1531);
and U3035 (N_3035,N_2362,N_127);
or U3036 (N_3036,N_2310,N_392);
nor U3037 (N_3037,N_557,N_353);
and U3038 (N_3038,N_2164,N_790);
nand U3039 (N_3039,N_1159,N_1080);
xnor U3040 (N_3040,N_2096,N_1514);
or U3041 (N_3041,N_2130,N_112);
nor U3042 (N_3042,N_509,N_2230);
or U3043 (N_3043,N_1419,N_983);
and U3044 (N_3044,N_677,N_558);
or U3045 (N_3045,N_2426,N_159);
nor U3046 (N_3046,N_2190,N_2365);
nor U3047 (N_3047,N_2377,N_2084);
nand U3048 (N_3048,N_471,N_1731);
nor U3049 (N_3049,N_1069,N_487);
or U3050 (N_3050,N_1824,N_710);
nor U3051 (N_3051,N_546,N_670);
nand U3052 (N_3052,N_2494,N_2087);
nor U3053 (N_3053,N_1359,N_1275);
nor U3054 (N_3054,N_1374,N_1372);
and U3055 (N_3055,N_1055,N_1062);
or U3056 (N_3056,N_1500,N_585);
or U3057 (N_3057,N_2021,N_1515);
and U3058 (N_3058,N_951,N_889);
nor U3059 (N_3059,N_1867,N_300);
or U3060 (N_3060,N_72,N_334);
nand U3061 (N_3061,N_310,N_682);
nor U3062 (N_3062,N_6,N_720);
or U3063 (N_3063,N_1031,N_906);
and U3064 (N_3064,N_376,N_1745);
nor U3065 (N_3065,N_520,N_1795);
and U3066 (N_3066,N_856,N_1017);
nand U3067 (N_3067,N_1276,N_1320);
and U3068 (N_3068,N_2037,N_290);
and U3069 (N_3069,N_1116,N_2258);
nand U3070 (N_3070,N_30,N_94);
nor U3071 (N_3071,N_1920,N_1286);
nor U3072 (N_3072,N_681,N_1668);
nand U3073 (N_3073,N_799,N_208);
or U3074 (N_3074,N_408,N_147);
and U3075 (N_3075,N_945,N_404);
nor U3076 (N_3076,N_1408,N_2182);
nand U3077 (N_3077,N_1104,N_1188);
nand U3078 (N_3078,N_1457,N_727);
nand U3079 (N_3079,N_496,N_491);
nor U3080 (N_3080,N_196,N_5);
nand U3081 (N_3081,N_505,N_219);
nand U3082 (N_3082,N_494,N_440);
nor U3083 (N_3083,N_1172,N_747);
and U3084 (N_3084,N_577,N_1834);
or U3085 (N_3085,N_1474,N_1539);
or U3086 (N_3086,N_2090,N_976);
or U3087 (N_3087,N_1935,N_1682);
nor U3088 (N_3088,N_2285,N_2223);
and U3089 (N_3089,N_2344,N_1176);
or U3090 (N_3090,N_1045,N_1435);
nor U3091 (N_3091,N_1440,N_657);
nor U3092 (N_3092,N_2469,N_108);
nand U3093 (N_3093,N_503,N_649);
nand U3094 (N_3094,N_597,N_2448);
nor U3095 (N_3095,N_667,N_1883);
or U3096 (N_3096,N_687,N_1288);
nor U3097 (N_3097,N_1509,N_2483);
nor U3098 (N_3098,N_507,N_1264);
nor U3099 (N_3099,N_1073,N_1534);
nand U3100 (N_3100,N_806,N_100);
or U3101 (N_3101,N_1272,N_518);
and U3102 (N_3102,N_1818,N_802);
or U3103 (N_3103,N_1551,N_2248);
nor U3104 (N_3104,N_2398,N_603);
nand U3105 (N_3105,N_338,N_1865);
and U3106 (N_3106,N_1616,N_1121);
and U3107 (N_3107,N_314,N_1155);
nor U3108 (N_3108,N_161,N_1699);
nor U3109 (N_3109,N_152,N_2359);
or U3110 (N_3110,N_1567,N_381);
nand U3111 (N_3111,N_2134,N_366);
or U3112 (N_3112,N_2352,N_2076);
and U3113 (N_3113,N_216,N_409);
and U3114 (N_3114,N_1700,N_1602);
and U3115 (N_3115,N_1442,N_85);
or U3116 (N_3116,N_1423,N_1885);
nor U3117 (N_3117,N_130,N_868);
and U3118 (N_3118,N_182,N_1212);
and U3119 (N_3119,N_2459,N_257);
or U3120 (N_3120,N_1014,N_1371);
or U3121 (N_3121,N_1205,N_1025);
or U3122 (N_3122,N_1823,N_643);
and U3123 (N_3123,N_928,N_2216);
or U3124 (N_3124,N_549,N_341);
and U3125 (N_3125,N_645,N_2482);
or U3126 (N_3126,N_265,N_1581);
nor U3127 (N_3127,N_1872,N_2177);
and U3128 (N_3128,N_172,N_2281);
nor U3129 (N_3129,N_1219,N_262);
nor U3130 (N_3130,N_867,N_605);
nand U3131 (N_3131,N_1269,N_993);
nor U3132 (N_3132,N_1672,N_332);
xor U3133 (N_3133,N_1221,N_2070);
nor U3134 (N_3134,N_2144,N_232);
or U3135 (N_3135,N_686,N_1292);
nand U3136 (N_3136,N_75,N_460);
or U3137 (N_3137,N_1197,N_459);
nor U3138 (N_3138,N_1013,N_2111);
or U3139 (N_3139,N_2257,N_586);
nor U3140 (N_3140,N_1493,N_14);
and U3141 (N_3141,N_1987,N_2363);
or U3142 (N_3142,N_2267,N_2489);
nor U3143 (N_3143,N_567,N_673);
nand U3144 (N_3144,N_1574,N_2470);
and U3145 (N_3145,N_2241,N_125);
nand U3146 (N_3146,N_1012,N_584);
nor U3147 (N_3147,N_375,N_26);
and U3148 (N_3148,N_693,N_2300);
nand U3149 (N_3149,N_291,N_1446);
and U3150 (N_3150,N_794,N_2477);
nor U3151 (N_3151,N_1607,N_1760);
and U3152 (N_3152,N_1383,N_961);
nand U3153 (N_3153,N_1932,N_1469);
or U3154 (N_3154,N_1622,N_1706);
nand U3155 (N_3155,N_1175,N_2402);
nand U3156 (N_3156,N_1971,N_178);
nor U3157 (N_3157,N_2274,N_1334);
nand U3158 (N_3158,N_1148,N_2210);
nor U3159 (N_3159,N_2165,N_330);
and U3160 (N_3160,N_2196,N_97);
nor U3161 (N_3161,N_939,N_1342);
nor U3162 (N_3162,N_1721,N_2481);
nor U3163 (N_3163,N_625,N_1791);
nand U3164 (N_3164,N_1254,N_1297);
nand U3165 (N_3165,N_1257,N_2334);
nor U3166 (N_3166,N_2290,N_966);
nand U3167 (N_3167,N_955,N_475);
or U3168 (N_3168,N_2498,N_1630);
or U3169 (N_3169,N_1643,N_2256);
and U3170 (N_3170,N_861,N_2392);
and U3171 (N_3171,N_815,N_779);
nand U3172 (N_3172,N_1281,N_1973);
or U3173 (N_3173,N_936,N_1717);
or U3174 (N_3174,N_1540,N_537);
and U3175 (N_3175,N_2242,N_824);
or U3176 (N_3176,N_234,N_821);
or U3177 (N_3177,N_1740,N_1190);
and U3178 (N_3178,N_223,N_1635);
or U3179 (N_3179,N_883,N_36);
or U3180 (N_3180,N_2478,N_1280);
or U3181 (N_3181,N_709,N_1751);
or U3182 (N_3182,N_825,N_1902);
and U3183 (N_3183,N_595,N_24);
or U3184 (N_3184,N_1817,N_863);
and U3185 (N_3185,N_456,N_631);
and U3186 (N_3186,N_398,N_354);
and U3187 (N_3187,N_1162,N_1669);
or U3188 (N_3188,N_2270,N_105);
xor U3189 (N_3189,N_2468,N_1541);
nand U3190 (N_3190,N_1130,N_1140);
nand U3191 (N_3191,N_1912,N_69);
and U3192 (N_3192,N_1441,N_1692);
nor U3193 (N_3193,N_1754,N_2307);
nand U3194 (N_3194,N_2009,N_946);
and U3195 (N_3195,N_2250,N_1027);
nor U3196 (N_3196,N_2148,N_761);
nor U3197 (N_3197,N_895,N_832);
or U3198 (N_3198,N_1345,N_1189);
or U3199 (N_3199,N_1648,N_903);
nand U3200 (N_3200,N_953,N_355);
xor U3201 (N_3201,N_468,N_996);
nor U3202 (N_3202,N_539,N_2299);
or U3203 (N_3203,N_1558,N_1127);
or U3204 (N_3204,N_1450,N_1886);
and U3205 (N_3205,N_2382,N_1638);
or U3206 (N_3206,N_11,N_280);
nor U3207 (N_3207,N_183,N_1956);
nor U3208 (N_3208,N_436,N_1619);
and U3209 (N_3209,N_2015,N_2166);
or U3210 (N_3210,N_1034,N_2156);
nor U3211 (N_3211,N_331,N_1783);
nor U3212 (N_3212,N_1898,N_98);
or U3213 (N_3213,N_2098,N_739);
and U3214 (N_3214,N_579,N_493);
nor U3215 (N_3215,N_2049,N_2369);
nor U3216 (N_3216,N_1231,N_1942);
or U3217 (N_3217,N_705,N_1921);
and U3218 (N_3218,N_694,N_719);
or U3219 (N_3219,N_1009,N_944);
and U3220 (N_3220,N_1488,N_622);
nor U3221 (N_3221,N_1479,N_1873);
nor U3222 (N_3222,N_663,N_1998);
and U3223 (N_3223,N_1960,N_1032);
and U3224 (N_3224,N_197,N_140);
nand U3225 (N_3225,N_425,N_1246);
nand U3226 (N_3226,N_619,N_80);
nand U3227 (N_3227,N_251,N_2083);
or U3228 (N_3228,N_2312,N_2030);
nand U3229 (N_3229,N_1517,N_514);
or U3230 (N_3230,N_123,N_1878);
and U3231 (N_3231,N_2169,N_2057);
xnor U3232 (N_3232,N_688,N_1958);
nor U3233 (N_3233,N_1951,N_2288);
nor U3234 (N_3234,N_1927,N_2079);
nand U3235 (N_3235,N_1671,N_1782);
nand U3236 (N_3236,N_1726,N_1398);
and U3237 (N_3237,N_2085,N_1997);
and U3238 (N_3238,N_1000,N_772);
or U3239 (N_3239,N_1589,N_1200);
or U3240 (N_3240,N_1884,N_2499);
or U3241 (N_3241,N_206,N_2444);
nor U3242 (N_3242,N_1714,N_1652);
nand U3243 (N_3243,N_2137,N_1995);
or U3244 (N_3244,N_1545,N_296);
and U3245 (N_3245,N_1677,N_611);
and U3246 (N_3246,N_1369,N_1202);
and U3247 (N_3247,N_2314,N_164);
and U3248 (N_3248,N_346,N_1124);
nand U3249 (N_3249,N_195,N_2443);
and U3250 (N_3250,N_2434,N_2017);
nor U3251 (N_3251,N_254,N_839);
or U3252 (N_3252,N_415,N_560);
nor U3253 (N_3253,N_1753,N_1451);
and U3254 (N_3254,N_1833,N_1761);
and U3255 (N_3255,N_428,N_1074);
nor U3256 (N_3256,N_405,N_754);
and U3257 (N_3257,N_534,N_467);
and U3258 (N_3258,N_1389,N_1267);
nand U3259 (N_3259,N_1696,N_785);
and U3260 (N_3260,N_1701,N_306);
xor U3261 (N_3261,N_1918,N_2236);
or U3262 (N_3262,N_738,N_455);
nand U3263 (N_3263,N_948,N_2208);
nor U3264 (N_3264,N_1708,N_1899);
or U3265 (N_3265,N_2191,N_2183);
or U3266 (N_3266,N_1118,N_1882);
nor U3267 (N_3267,N_1999,N_655);
nor U3268 (N_3268,N_1092,N_704);
nand U3269 (N_3269,N_1511,N_1943);
and U3270 (N_3270,N_1897,N_1738);
nor U3271 (N_3271,N_1917,N_114);
nor U3272 (N_3272,N_1636,N_2209);
nor U3273 (N_3273,N_656,N_1712);
nand U3274 (N_3274,N_519,N_446);
or U3275 (N_3275,N_674,N_2220);
nor U3276 (N_3276,N_2217,N_2179);
nor U3277 (N_3277,N_1827,N_1564);
nand U3278 (N_3278,N_2193,N_1591);
or U3279 (N_3279,N_991,N_2421);
or U3280 (N_3280,N_672,N_57);
and U3281 (N_3281,N_2455,N_1604);
or U3282 (N_3282,N_1513,N_2139);
and U3283 (N_3283,N_865,N_136);
or U3284 (N_3284,N_1482,N_576);
nand U3285 (N_3285,N_1723,N_1680);
and U3286 (N_3286,N_728,N_115);
xnor U3287 (N_3287,N_887,N_453);
and U3288 (N_3288,N_2412,N_1977);
and U3289 (N_3289,N_1516,N_1911);
nor U3290 (N_3290,N_1030,N_1051);
nand U3291 (N_3291,N_1097,N_2238);
and U3292 (N_3292,N_834,N_1495);
nor U3293 (N_3293,N_499,N_1295);
or U3294 (N_3294,N_2322,N_1743);
nand U3295 (N_3295,N_1026,N_1594);
nor U3296 (N_3296,N_2261,N_304);
and U3297 (N_3297,N_713,N_104);
nand U3298 (N_3298,N_1238,N_12);
or U3299 (N_3299,N_2199,N_2275);
nand U3300 (N_3300,N_2133,N_1803);
nand U3301 (N_3301,N_1262,N_1837);
nor U3302 (N_3302,N_2016,N_1861);
nor U3303 (N_3303,N_1590,N_1277);
and U3304 (N_3304,N_189,N_1024);
or U3305 (N_3305,N_2029,N_1321);
or U3306 (N_3306,N_488,N_2186);
and U3307 (N_3307,N_1453,N_1357);
and U3308 (N_3308,N_2212,N_1307);
or U3309 (N_3309,N_1720,N_1350);
nor U3310 (N_3310,N_402,N_1940);
nor U3311 (N_3311,N_553,N_1593);
or U3312 (N_3312,N_1512,N_465);
nor U3313 (N_3313,N_342,N_925);
nand U3314 (N_3314,N_19,N_1481);
and U3315 (N_3315,N_2380,N_111);
or U3316 (N_3316,N_1732,N_731);
nand U3317 (N_3317,N_2113,N_1949);
or U3318 (N_3318,N_1245,N_2065);
nor U3319 (N_3319,N_2172,N_969);
nand U3320 (N_3320,N_664,N_893);
nand U3321 (N_3321,N_1170,N_1406);
nor U3322 (N_3322,N_176,N_2197);
nand U3323 (N_3323,N_565,N_941);
and U3324 (N_3324,N_1433,N_1639);
or U3325 (N_3325,N_109,N_607);
nand U3326 (N_3326,N_756,N_319);
nand U3327 (N_3327,N_2043,N_1606);
nand U3328 (N_3328,N_2089,N_1337);
nor U3329 (N_3329,N_260,N_158);
nand U3330 (N_3330,N_2131,N_1084);
or U3331 (N_3331,N_101,N_716);
nor U3332 (N_3332,N_2126,N_732);
nor U3333 (N_3333,N_1502,N_1587);
and U3334 (N_3334,N_1146,N_1210);
and U3335 (N_3335,N_1163,N_1755);
nand U3336 (N_3336,N_2418,N_1412);
nand U3337 (N_3337,N_2051,N_1088);
and U3338 (N_3338,N_2157,N_1328);
and U3339 (N_3339,N_490,N_1181);
nor U3340 (N_3340,N_54,N_608);
nand U3341 (N_3341,N_121,N_134);
or U3342 (N_3342,N_745,N_1375);
nand U3343 (N_3343,N_1774,N_1880);
and U3344 (N_3344,N_1888,N_2259);
nor U3345 (N_3345,N_71,N_1750);
nand U3346 (N_3346,N_1825,N_1769);
nand U3347 (N_3347,N_66,N_122);
nand U3348 (N_3348,N_827,N_1766);
nor U3349 (N_3349,N_55,N_1627);
nand U3350 (N_3350,N_627,N_1461);
or U3351 (N_3351,N_853,N_1955);
and U3352 (N_3352,N_1360,N_1057);
nor U3353 (N_3353,N_1864,N_1983);
nor U3354 (N_3354,N_2345,N_1485);
or U3355 (N_3355,N_1906,N_2195);
nand U3356 (N_3356,N_1224,N_1037);
or U3357 (N_3357,N_2480,N_333);
and U3358 (N_3358,N_1167,N_312);
nand U3359 (N_3359,N_1542,N_934);
nand U3360 (N_3360,N_420,N_891);
and U3361 (N_3361,N_1220,N_214);
and U3362 (N_3362,N_276,N_2123);
nand U3363 (N_3363,N_639,N_990);
and U3364 (N_3364,N_914,N_1777);
nor U3365 (N_3365,N_1547,N_1689);
or U3366 (N_3366,N_184,N_230);
nor U3367 (N_3367,N_1050,N_2154);
nand U3368 (N_3368,N_526,N_2114);
and U3369 (N_3369,N_1642,N_2056);
or U3370 (N_3370,N_2091,N_1108);
or U3371 (N_3371,N_912,N_228);
nand U3372 (N_3372,N_2407,N_1459);
nor U3373 (N_3373,N_347,N_389);
nor U3374 (N_3374,N_95,N_322);
or U3375 (N_3375,N_800,N_862);
xnor U3376 (N_3376,N_566,N_582);
nand U3377 (N_3377,N_2389,N_1077);
or U3378 (N_3378,N_898,N_500);
and U3379 (N_3379,N_513,N_1193);
nor U3380 (N_3380,N_992,N_2028);
nand U3381 (N_3381,N_1739,N_1182);
or U3382 (N_3382,N_1468,N_1858);
and U3383 (N_3383,N_807,N_1310);
nor U3384 (N_3384,N_1237,N_1494);
nand U3385 (N_3385,N_238,N_364);
nor U3386 (N_3386,N_2383,N_445);
nand U3387 (N_3387,N_937,N_1217);
nor U3388 (N_3388,N_210,N_2335);
or U3389 (N_3389,N_2330,N_2);
nor U3390 (N_3390,N_1174,N_2189);
and U3391 (N_3391,N_1105,N_435);
or U3392 (N_3392,N_1781,N_911);
nand U3393 (N_3393,N_831,N_168);
and U3394 (N_3394,N_1676,N_2428);
or U3395 (N_3395,N_2058,N_198);
and U3396 (N_3396,N_968,N_486);
or U3397 (N_3397,N_2340,N_1230);
and U3398 (N_3398,N_432,N_640);
and U3399 (N_3399,N_2496,N_633);
nor U3400 (N_3400,N_845,N_1085);
or U3401 (N_3401,N_1002,N_2413);
or U3402 (N_3402,N_374,N_1386);
nor U3403 (N_3403,N_763,N_56);
xor U3404 (N_3404,N_2246,N_618);
nor U3405 (N_3405,N_523,N_263);
or U3406 (N_3406,N_286,N_1868);
nor U3407 (N_3407,N_2011,N_1036);
or U3408 (N_3408,N_525,N_1184);
nor U3409 (N_3409,N_1525,N_722);
nand U3410 (N_3410,N_2004,N_1003);
nor U3411 (N_3411,N_1339,N_2031);
and U3412 (N_3412,N_598,N_449);
nand U3413 (N_3413,N_1436,N_2005);
nor U3414 (N_3414,N_717,N_1301);
nor U3415 (N_3415,N_1298,N_2115);
and U3416 (N_3416,N_229,N_13);
and U3417 (N_3417,N_18,N_1603);
nand U3418 (N_3418,N_1007,N_723);
nor U3419 (N_3419,N_1487,N_484);
nor U3420 (N_3420,N_162,N_166);
nand U3421 (N_3421,N_1323,N_1204);
and U3422 (N_3422,N_79,N_1655);
nand U3423 (N_3423,N_89,N_1142);
nor U3424 (N_3424,N_1366,N_2171);
nand U3425 (N_3425,N_339,N_1390);
nor U3426 (N_3426,N_2339,N_1);
nand U3427 (N_3427,N_2198,N_1695);
nand U3428 (N_3428,N_1064,N_1505);
and U3429 (N_3429,N_311,N_650);
and U3430 (N_3430,N_173,N_2240);
or U3431 (N_3431,N_2308,N_1651);
and U3432 (N_3432,N_1610,N_113);
nand U3433 (N_3433,N_1503,N_62);
nand U3434 (N_3434,N_1222,N_1422);
or U3435 (N_3435,N_2495,N_463);
nor U3436 (N_3436,N_186,N_1909);
xnor U3437 (N_3437,N_1821,N_1931);
nand U3438 (N_3438,N_145,N_294);
nand U3439 (N_3439,N_1132,N_1427);
nand U3440 (N_3440,N_1986,N_1315);
nor U3441 (N_3441,N_1856,N_60);
and U3442 (N_3442,N_84,N_191);
nor U3443 (N_3443,N_899,N_139);
nand U3444 (N_3444,N_1056,N_243);
or U3445 (N_3445,N_438,N_1626);
nor U3446 (N_3446,N_636,N_2324);
nand U3447 (N_3447,N_823,N_1707);
or U3448 (N_3448,N_1376,N_1233);
or U3449 (N_3449,N_1370,N_412);
and U3450 (N_3450,N_1741,N_1229);
and U3451 (N_3451,N_604,N_994);
and U3452 (N_3452,N_2458,N_2348);
xor U3453 (N_3453,N_1225,N_1537);
nand U3454 (N_3454,N_1363,N_2420);
and U3455 (N_3455,N_1660,N_448);
or U3456 (N_3456,N_2401,N_1141);
and U3457 (N_3457,N_1875,N_2225);
nor U3458 (N_3458,N_2082,N_515);
or U3459 (N_3459,N_1901,N_614);
and U3460 (N_3460,N_2287,N_185);
and U3461 (N_3461,N_1089,N_659);
or U3462 (N_3462,N_20,N_2318);
and U3463 (N_3463,N_921,N_1203);
or U3464 (N_3464,N_175,N_1523);
and U3465 (N_3465,N_144,N_2067);
or U3466 (N_3466,N_1952,N_1650);
or U3467 (N_3467,N_778,N_313);
nand U3468 (N_3468,N_901,N_1736);
and U3469 (N_3469,N_888,N_679);
or U3470 (N_3470,N_2390,N_975);
nand U3471 (N_3471,N_35,N_1929);
and U3472 (N_3472,N_1319,N_707);
nor U3473 (N_3473,N_635,N_757);
or U3474 (N_3474,N_1058,N_1722);
or U3475 (N_3475,N_43,N_1877);
and U3476 (N_3476,N_1963,N_1654);
nand U3477 (N_3477,N_1445,N_1710);
or U3478 (N_3478,N_2214,N_1691);
and U3479 (N_3479,N_270,N_1195);
and U3480 (N_3480,N_665,N_940);
nand U3481 (N_3481,N_1090,N_40);
or U3482 (N_3482,N_699,N_2027);
nand U3483 (N_3483,N_1209,N_1447);
nor U3484 (N_3484,N_962,N_1582);
or U3485 (N_3485,N_2388,N_1329);
or U3486 (N_3486,N_1544,N_1891);
nand U3487 (N_3487,N_2095,N_1839);
and U3488 (N_3488,N_2276,N_1628);
or U3489 (N_3489,N_1820,N_1166);
or U3490 (N_3490,N_1794,N_808);
and U3491 (N_3491,N_2025,N_1439);
nor U3492 (N_3492,N_2054,N_233);
and U3493 (N_3493,N_1010,N_775);
nand U3494 (N_3494,N_63,N_1214);
nand U3495 (N_3495,N_482,N_935);
xor U3496 (N_3496,N_742,N_1845);
nand U3497 (N_3497,N_1681,N_1838);
xnor U3498 (N_3498,N_1353,N_698);
nor U3499 (N_3499,N_1187,N_2118);
or U3500 (N_3500,N_1075,N_1914);
or U3501 (N_3501,N_905,N_612);
nand U3502 (N_3502,N_2327,N_1094);
nor U3503 (N_3503,N_1862,N_2180);
or U3504 (N_3504,N_2014,N_480);
or U3505 (N_3505,N_671,N_383);
or U3506 (N_3506,N_956,N_1305);
nor U3507 (N_3507,N_669,N_39);
or U3508 (N_3508,N_1601,N_293);
nor U3509 (N_3509,N_1966,N_2032);
and U3510 (N_3510,N_599,N_1640);
nand U3511 (N_3511,N_278,N_843);
or U3512 (N_3512,N_871,N_1623);
or U3513 (N_3513,N_2331,N_545);
nor U3514 (N_3514,N_1287,N_1819);
nor U3515 (N_3515,N_2033,N_850);
xor U3516 (N_3516,N_2102,N_855);
nand U3517 (N_3517,N_965,N_2116);
or U3518 (N_3518,N_828,N_602);
nand U3519 (N_3519,N_1992,N_452);
nor U3520 (N_3520,N_2497,N_1976);
nor U3521 (N_3521,N_1318,N_1120);
and U3522 (N_3522,N_849,N_1291);
and U3523 (N_3523,N_678,N_1611);
or U3524 (N_3524,N_1854,N_367);
and U3525 (N_3525,N_1382,N_583);
and U3526 (N_3526,N_1282,N_1107);
or U3527 (N_3527,N_2386,N_1600);
and U3528 (N_3528,N_1086,N_2254);
nand U3529 (N_3529,N_384,N_46);
nand U3530 (N_3530,N_2378,N_1096);
nor U3531 (N_3531,N_0,N_274);
or U3532 (N_3532,N_1004,N_1005);
or U3533 (N_3533,N_2120,N_1895);
or U3534 (N_3534,N_237,N_2473);
nor U3535 (N_3535,N_2110,N_897);
or U3536 (N_3536,N_200,N_431);
nor U3537 (N_3537,N_2042,N_151);
nor U3538 (N_3538,N_529,N_1261);
nor U3539 (N_3539,N_2351,N_380);
nor U3540 (N_3540,N_2461,N_818);
nor U3541 (N_3541,N_527,N_203);
or U3542 (N_3542,N_2187,N_2052);
or U3543 (N_3543,N_2396,N_395);
nor U3544 (N_3544,N_403,N_451);
and U3545 (N_3545,N_211,N_1112);
nor U3546 (N_3546,N_2138,N_1989);
and U3547 (N_3547,N_2235,N_581);
nor U3548 (N_3548,N_249,N_190);
nand U3549 (N_3549,N_882,N_1779);
or U3550 (N_3550,N_2101,N_809);
nor U3551 (N_3551,N_1687,N_177);
or U3552 (N_3552,N_2264,N_915);
nand U3553 (N_3553,N_2245,N_1153);
nand U3554 (N_3554,N_2075,N_2317);
or U3555 (N_3555,N_601,N_1698);
nand U3556 (N_3556,N_623,N_1368);
nor U3557 (N_3557,N_730,N_632);
nand U3558 (N_3558,N_1697,N_615);
or U3559 (N_3559,N_1724,N_1572);
or U3560 (N_3560,N_1688,N_2316);
and U3561 (N_3561,N_1773,N_1206);
and U3562 (N_3562,N_1562,N_1367);
nand U3563 (N_3563,N_86,N_886);
or U3564 (N_3564,N_995,N_1730);
and U3565 (N_3565,N_1428,N_1052);
nand U3566 (N_3566,N_734,N_563);
nor U3567 (N_3567,N_1028,N_1728);
and U3568 (N_3568,N_532,N_1046);
or U3569 (N_3569,N_2414,N_572);
nand U3570 (N_3570,N_764,N_1569);
nand U3571 (N_3571,N_2038,N_1215);
nor U3572 (N_3572,N_2269,N_2417);
and U3573 (N_3573,N_1796,N_1715);
or U3574 (N_3574,N_652,N_2161);
nand U3575 (N_3575,N_1571,N_2302);
or U3576 (N_3576,N_1850,N_502);
and U3577 (N_3577,N_1228,N_1270);
or U3578 (N_3578,N_2035,N_1578);
nor U3579 (N_3579,N_2268,N_120);
and U3580 (N_3580,N_1673,N_1553);
and U3581 (N_3581,N_2152,N_2346);
or U3582 (N_3582,N_495,N_1133);
nand U3583 (N_3583,N_1448,N_1559);
and U3584 (N_3584,N_343,N_1156);
nand U3585 (N_3585,N_150,N_492);
or U3586 (N_3586,N_1068,N_841);
nand U3587 (N_3587,N_1048,N_1169);
or U3588 (N_3588,N_1576,N_1922);
nor U3589 (N_3589,N_740,N_1335);
and U3590 (N_3590,N_328,N_805);
and U3591 (N_3591,N_1179,N_2337);
nand U3592 (N_3592,N_1756,N_575);
nand U3593 (N_3593,N_476,N_613);
and U3594 (N_3594,N_1273,N_2490);
or U3595 (N_3595,N_1019,N_642);
or U3596 (N_3596,N_156,N_1065);
nor U3597 (N_3597,N_222,N_358);
and U3598 (N_3598,N_2200,N_244);
nor U3599 (N_3599,N_1550,N_2170);
or U3600 (N_3600,N_1384,N_2447);
nor U3601 (N_3601,N_648,N_638);
or U3602 (N_3602,N_321,N_21);
or U3603 (N_3603,N_2277,N_2371);
or U3604 (N_3604,N_1768,N_1460);
or U3605 (N_3605,N_2020,N_1770);
and U3606 (N_3606,N_2460,N_1125);
and U3607 (N_3607,N_400,N_959);
or U3608 (N_3608,N_447,N_201);
nand U3609 (N_3609,N_474,N_1847);
nor U3610 (N_3610,N_2297,N_292);
nor U3611 (N_3611,N_989,N_1787);
or U3612 (N_3612,N_469,N_1149);
nor U3613 (N_3613,N_2452,N_1737);
xor U3614 (N_3614,N_1916,N_307);
or U3615 (N_3615,N_541,N_1894);
nor U3616 (N_3616,N_776,N_2255);
xor U3617 (N_3617,N_1663,N_1480);
or U3618 (N_3618,N_729,N_1746);
or U3619 (N_3619,N_288,N_1810);
nor U3620 (N_3620,N_626,N_2002);
or U3621 (N_3621,N_1308,N_1957);
nor U3622 (N_3622,N_1752,N_1413);
xor U3623 (N_3623,N_309,N_1463);
nor U3624 (N_3624,N_1804,N_29);
or U3625 (N_3625,N_654,N_517);
nand U3626 (N_3626,N_960,N_1807);
or U3627 (N_3627,N_2077,N_1312);
or U3628 (N_3628,N_218,N_1684);
nor U3629 (N_3629,N_1154,N_1996);
nand U3630 (N_3630,N_685,N_765);
nor U3631 (N_3631,N_2266,N_2319);
nand U3632 (N_3632,N_2416,N_562);
and U3633 (N_3633,N_170,N_2128);
and U3634 (N_3634,N_1410,N_2109);
nand U3635 (N_3635,N_2405,N_269);
nor U3636 (N_3636,N_433,N_629);
or U3637 (N_3637,N_609,N_873);
nand U3638 (N_3638,N_812,N_1584);
nand U3639 (N_3639,N_1478,N_96);
nor U3640 (N_3640,N_726,N_782);
nor U3641 (N_3641,N_1416,N_1327);
nor U3642 (N_3642,N_2303,N_2467);
and U3643 (N_3643,N_1904,N_241);
and U3644 (N_3644,N_1566,N_2097);
nor U3645 (N_3645,N_324,N_437);
and U3646 (N_3646,N_401,N_997);
and U3647 (N_3647,N_3,N_1506);
or U3648 (N_3648,N_422,N_753);
nand U3649 (N_3649,N_548,N_142);
nor U3650 (N_3650,N_271,N_1038);
and U3651 (N_3651,N_1612,N_1802);
or U3652 (N_3652,N_506,N_988);
and U3653 (N_3653,N_2012,N_1194);
nor U3654 (N_3654,N_2239,N_1067);
or U3655 (N_3655,N_2162,N_2122);
or U3656 (N_3656,N_119,N_2432);
nand U3657 (N_3657,N_1411,N_1054);
and U3658 (N_3658,N_1489,N_1649);
and U3659 (N_3659,N_1829,N_1871);
nand U3660 (N_3660,N_58,N_1785);
or U3661 (N_3661,N_755,N_2282);
or U3662 (N_3662,N_50,N_1595);
or U3663 (N_3663,N_1849,N_2328);
nand U3664 (N_3664,N_61,N_1100);
nor U3665 (N_3665,N_676,N_999);
nand U3666 (N_3666,N_1134,N_1592);
xnor U3667 (N_3667,N_528,N_1265);
or U3668 (N_3668,N_1351,N_788);
and U3669 (N_3669,N_1580,N_820);
and U3670 (N_3670,N_644,N_2422);
nand U3671 (N_3671,N_443,N_2215);
and U3672 (N_3672,N_1860,N_1970);
nor U3673 (N_3673,N_2201,N_102);
and U3674 (N_3674,N_1449,N_419);
xor U3675 (N_3675,N_406,N_1250);
or U3676 (N_3676,N_1851,N_1354);
nand U3677 (N_3677,N_1432,N_246);
nand U3678 (N_3678,N_2107,N_758);
nand U3679 (N_3679,N_2061,N_1490);
and U3680 (N_3680,N_1070,N_1160);
nand U3681 (N_3681,N_1508,N_1496);
nor U3682 (N_3682,N_1843,N_870);
nand U3683 (N_3683,N_864,N_980);
nand U3684 (N_3684,N_1365,N_816);
nand U3685 (N_3685,N_2088,N_2492);
and U3686 (N_3686,N_497,N_1561);
nor U3687 (N_3687,N_920,N_746);
and U3688 (N_3688,N_1826,N_2488);
nor U3689 (N_3689,N_592,N_1266);
or U3690 (N_3690,N_916,N_2143);
nand U3691 (N_3691,N_266,N_444);
or U3692 (N_3692,N_1815,N_766);
or U3693 (N_3693,N_964,N_1546);
and U3694 (N_3694,N_1393,N_327);
and U3695 (N_3695,N_1290,N_2476);
and U3696 (N_3696,N_2338,N_275);
nor U3697 (N_3697,N_44,N_569);
or U3698 (N_3698,N_478,N_533);
and U3699 (N_3699,N_52,N_1974);
and U3700 (N_3700,N_382,N_1526);
nor U3701 (N_3701,N_789,N_902);
or U3702 (N_3702,N_369,N_620);
or U3703 (N_3703,N_646,N_2073);
and U3704 (N_3704,N_1903,N_2366);
nor U3705 (N_3705,N_1168,N_1713);
or U3706 (N_3706,N_248,N_226);
nand U3707 (N_3707,N_661,N_1437);
nor U3708 (N_3708,N_2408,N_1041);
and U3709 (N_3709,N_45,N_1015);
and U3710 (N_3710,N_192,N_1296);
nor U3711 (N_3711,N_28,N_2450);
nor U3712 (N_3712,N_1842,N_2160);
and U3713 (N_3713,N_958,N_574);
nand U3714 (N_3714,N_1498,N_2202);
nand U3715 (N_3715,N_555,N_1022);
nor U3716 (N_3716,N_267,N_938);
and U3717 (N_3717,N_37,N_315);
nand U3718 (N_3718,N_1274,N_2403);
nor U3719 (N_3719,N_245,N_544);
nand U3720 (N_3720,N_1243,N_508);
nand U3721 (N_3721,N_2347,N_540);
and U3722 (N_3722,N_1887,N_1475);
nand U3723 (N_3723,N_1223,N_303);
and U3724 (N_3724,N_1962,N_2103);
nand U3725 (N_3725,N_1258,N_1192);
nor U3726 (N_3726,N_2278,N_972);
and U3727 (N_3727,N_394,N_272);
nor U3728 (N_3728,N_1053,N_675);
nor U3729 (N_3729,N_2018,N_1813);
or U3730 (N_3730,N_390,N_942);
nand U3731 (N_3731,N_1183,N_1778);
or U3732 (N_3732,N_1596,N_858);
or U3733 (N_3733,N_1620,N_154);
nor U3734 (N_3734,N_2080,N_880);
nand U3735 (N_3735,N_2140,N_516);
nand U3736 (N_3736,N_1122,N_417);
nand U3737 (N_3737,N_590,N_70);
nand U3738 (N_3738,N_53,N_1686);
or U3739 (N_3739,N_1954,N_221);
and U3740 (N_3740,N_1857,N_2121);
or U3741 (N_3741,N_1588,N_179);
nand U3742 (N_3742,N_2227,N_737);
nor U3743 (N_3743,N_724,N_2055);
nand U3744 (N_3744,N_1082,N_1797);
and U3745 (N_3745,N_875,N_2333);
or U3746 (N_3746,N_879,N_974);
nor U3747 (N_3747,N_1520,N_712);
nand U3748 (N_3748,N_1809,N_930);
nand U3749 (N_3749,N_1780,N_1344);
or U3750 (N_3750,N_1657,N_526);
and U3751 (N_3751,N_2064,N_840);
and U3752 (N_3752,N_2210,N_274);
nand U3753 (N_3753,N_2169,N_1893);
and U3754 (N_3754,N_1218,N_1811);
and U3755 (N_3755,N_1448,N_1191);
and U3756 (N_3756,N_36,N_1780);
xor U3757 (N_3757,N_969,N_2001);
and U3758 (N_3758,N_2472,N_1260);
or U3759 (N_3759,N_1706,N_379);
and U3760 (N_3760,N_574,N_588);
or U3761 (N_3761,N_1302,N_1065);
or U3762 (N_3762,N_1650,N_1697);
nand U3763 (N_3763,N_74,N_2108);
nand U3764 (N_3764,N_1220,N_1527);
and U3765 (N_3765,N_1445,N_1355);
nor U3766 (N_3766,N_868,N_966);
nand U3767 (N_3767,N_936,N_1445);
nand U3768 (N_3768,N_963,N_534);
or U3769 (N_3769,N_984,N_1847);
or U3770 (N_3770,N_1873,N_2356);
nand U3771 (N_3771,N_568,N_1357);
and U3772 (N_3772,N_1449,N_1547);
nor U3773 (N_3773,N_480,N_1432);
or U3774 (N_3774,N_2205,N_765);
nor U3775 (N_3775,N_1749,N_809);
and U3776 (N_3776,N_1945,N_1700);
and U3777 (N_3777,N_1939,N_386);
nor U3778 (N_3778,N_1018,N_2140);
nor U3779 (N_3779,N_2336,N_689);
nand U3780 (N_3780,N_1473,N_645);
nor U3781 (N_3781,N_307,N_637);
nand U3782 (N_3782,N_878,N_938);
nand U3783 (N_3783,N_5,N_634);
or U3784 (N_3784,N_235,N_2395);
nor U3785 (N_3785,N_2183,N_941);
nand U3786 (N_3786,N_638,N_420);
nor U3787 (N_3787,N_787,N_2242);
or U3788 (N_3788,N_1061,N_1234);
nor U3789 (N_3789,N_1568,N_2448);
or U3790 (N_3790,N_861,N_882);
nand U3791 (N_3791,N_714,N_725);
and U3792 (N_3792,N_136,N_1065);
or U3793 (N_3793,N_2149,N_314);
nand U3794 (N_3794,N_1396,N_303);
or U3795 (N_3795,N_1736,N_879);
and U3796 (N_3796,N_1065,N_2341);
nand U3797 (N_3797,N_1161,N_46);
nand U3798 (N_3798,N_1020,N_777);
or U3799 (N_3799,N_2048,N_2422);
xor U3800 (N_3800,N_820,N_2443);
and U3801 (N_3801,N_2240,N_1204);
and U3802 (N_3802,N_2178,N_189);
nand U3803 (N_3803,N_2106,N_2002);
or U3804 (N_3804,N_1019,N_1056);
nor U3805 (N_3805,N_68,N_2466);
xor U3806 (N_3806,N_1411,N_280);
nand U3807 (N_3807,N_1964,N_2112);
nor U3808 (N_3808,N_246,N_1847);
nor U3809 (N_3809,N_2246,N_1760);
and U3810 (N_3810,N_1203,N_1284);
nand U3811 (N_3811,N_1032,N_355);
nand U3812 (N_3812,N_315,N_1699);
and U3813 (N_3813,N_1989,N_1837);
and U3814 (N_3814,N_121,N_1250);
nor U3815 (N_3815,N_1653,N_1725);
nor U3816 (N_3816,N_1861,N_443);
xnor U3817 (N_3817,N_2373,N_950);
xor U3818 (N_3818,N_1039,N_2079);
nand U3819 (N_3819,N_1610,N_364);
or U3820 (N_3820,N_310,N_1703);
or U3821 (N_3821,N_2271,N_1778);
or U3822 (N_3822,N_764,N_6);
nor U3823 (N_3823,N_1795,N_470);
or U3824 (N_3824,N_878,N_2080);
and U3825 (N_3825,N_1915,N_298);
and U3826 (N_3826,N_1184,N_1637);
and U3827 (N_3827,N_2381,N_475);
nand U3828 (N_3828,N_80,N_460);
or U3829 (N_3829,N_1615,N_2328);
nand U3830 (N_3830,N_53,N_1086);
or U3831 (N_3831,N_249,N_177);
nand U3832 (N_3832,N_2200,N_1207);
or U3833 (N_3833,N_1674,N_1082);
or U3834 (N_3834,N_1963,N_2047);
or U3835 (N_3835,N_1153,N_1363);
nand U3836 (N_3836,N_250,N_665);
or U3837 (N_3837,N_2348,N_886);
nand U3838 (N_3838,N_1906,N_2181);
and U3839 (N_3839,N_2120,N_660);
nand U3840 (N_3840,N_2025,N_1965);
and U3841 (N_3841,N_1294,N_1696);
nand U3842 (N_3842,N_846,N_1790);
and U3843 (N_3843,N_1109,N_2402);
nor U3844 (N_3844,N_537,N_1387);
nor U3845 (N_3845,N_1915,N_2337);
and U3846 (N_3846,N_2078,N_529);
or U3847 (N_3847,N_2223,N_1813);
and U3848 (N_3848,N_210,N_512);
nand U3849 (N_3849,N_2249,N_574);
or U3850 (N_3850,N_1180,N_1908);
or U3851 (N_3851,N_2370,N_1408);
nor U3852 (N_3852,N_114,N_621);
nand U3853 (N_3853,N_1714,N_2179);
nor U3854 (N_3854,N_1813,N_2101);
nand U3855 (N_3855,N_1871,N_669);
nor U3856 (N_3856,N_2335,N_2325);
nor U3857 (N_3857,N_66,N_173);
and U3858 (N_3858,N_1447,N_2140);
and U3859 (N_3859,N_1117,N_32);
or U3860 (N_3860,N_1717,N_971);
or U3861 (N_3861,N_77,N_1975);
nor U3862 (N_3862,N_868,N_901);
nand U3863 (N_3863,N_603,N_36);
or U3864 (N_3864,N_1331,N_1608);
nand U3865 (N_3865,N_107,N_1574);
nand U3866 (N_3866,N_10,N_305);
nor U3867 (N_3867,N_1345,N_47);
nand U3868 (N_3868,N_955,N_162);
nor U3869 (N_3869,N_2127,N_1667);
and U3870 (N_3870,N_133,N_968);
nand U3871 (N_3871,N_1590,N_144);
or U3872 (N_3872,N_1461,N_528);
and U3873 (N_3873,N_1154,N_1194);
or U3874 (N_3874,N_1772,N_2456);
and U3875 (N_3875,N_1491,N_1312);
and U3876 (N_3876,N_895,N_2474);
nor U3877 (N_3877,N_483,N_2481);
nor U3878 (N_3878,N_1232,N_2426);
xor U3879 (N_3879,N_1368,N_852);
and U3880 (N_3880,N_1201,N_783);
nor U3881 (N_3881,N_1546,N_263);
nand U3882 (N_3882,N_2379,N_1214);
and U3883 (N_3883,N_959,N_2282);
or U3884 (N_3884,N_2331,N_845);
or U3885 (N_3885,N_2488,N_333);
nor U3886 (N_3886,N_784,N_321);
nor U3887 (N_3887,N_951,N_1323);
nand U3888 (N_3888,N_443,N_1325);
and U3889 (N_3889,N_407,N_931);
and U3890 (N_3890,N_979,N_1577);
or U3891 (N_3891,N_581,N_2307);
and U3892 (N_3892,N_1023,N_114);
nor U3893 (N_3893,N_2275,N_821);
nand U3894 (N_3894,N_778,N_1183);
and U3895 (N_3895,N_962,N_495);
and U3896 (N_3896,N_1691,N_1823);
and U3897 (N_3897,N_1919,N_1065);
nand U3898 (N_3898,N_1217,N_2491);
nor U3899 (N_3899,N_284,N_2348);
and U3900 (N_3900,N_1669,N_1688);
nand U3901 (N_3901,N_594,N_104);
nand U3902 (N_3902,N_1513,N_2405);
and U3903 (N_3903,N_482,N_1600);
and U3904 (N_3904,N_486,N_1835);
nor U3905 (N_3905,N_1326,N_2412);
and U3906 (N_3906,N_2329,N_1543);
nand U3907 (N_3907,N_680,N_1246);
or U3908 (N_3908,N_677,N_1833);
and U3909 (N_3909,N_184,N_1491);
nand U3910 (N_3910,N_2345,N_2455);
or U3911 (N_3911,N_674,N_1583);
and U3912 (N_3912,N_1075,N_1374);
or U3913 (N_3913,N_2227,N_2202);
nand U3914 (N_3914,N_1662,N_2402);
nor U3915 (N_3915,N_314,N_1665);
and U3916 (N_3916,N_551,N_1792);
and U3917 (N_3917,N_1561,N_229);
and U3918 (N_3918,N_1661,N_2481);
nand U3919 (N_3919,N_1182,N_5);
nor U3920 (N_3920,N_300,N_721);
and U3921 (N_3921,N_1311,N_1573);
nand U3922 (N_3922,N_2400,N_1853);
and U3923 (N_3923,N_1386,N_1205);
nor U3924 (N_3924,N_746,N_1460);
and U3925 (N_3925,N_629,N_986);
or U3926 (N_3926,N_1350,N_1319);
nor U3927 (N_3927,N_2090,N_483);
nor U3928 (N_3928,N_1603,N_206);
and U3929 (N_3929,N_1674,N_2037);
nand U3930 (N_3930,N_1793,N_2432);
nand U3931 (N_3931,N_1045,N_306);
nor U3932 (N_3932,N_1966,N_2480);
or U3933 (N_3933,N_1793,N_1218);
or U3934 (N_3934,N_391,N_327);
nor U3935 (N_3935,N_1319,N_809);
nand U3936 (N_3936,N_1368,N_1863);
nor U3937 (N_3937,N_1053,N_826);
or U3938 (N_3938,N_1691,N_2338);
nor U3939 (N_3939,N_1730,N_282);
nand U3940 (N_3940,N_2282,N_1512);
nand U3941 (N_3941,N_1704,N_2318);
and U3942 (N_3942,N_288,N_1896);
nor U3943 (N_3943,N_544,N_744);
nor U3944 (N_3944,N_1096,N_1545);
or U3945 (N_3945,N_2031,N_2164);
nor U3946 (N_3946,N_501,N_2028);
nand U3947 (N_3947,N_558,N_1254);
and U3948 (N_3948,N_2420,N_1896);
nor U3949 (N_3949,N_1342,N_964);
or U3950 (N_3950,N_872,N_1608);
and U3951 (N_3951,N_2102,N_488);
nor U3952 (N_3952,N_1663,N_2360);
and U3953 (N_3953,N_1192,N_795);
nor U3954 (N_3954,N_2202,N_107);
nand U3955 (N_3955,N_777,N_1806);
nand U3956 (N_3956,N_2178,N_532);
or U3957 (N_3957,N_1200,N_342);
nand U3958 (N_3958,N_1919,N_315);
nand U3959 (N_3959,N_579,N_600);
nor U3960 (N_3960,N_1362,N_2100);
and U3961 (N_3961,N_2362,N_396);
and U3962 (N_3962,N_1965,N_2448);
or U3963 (N_3963,N_1302,N_1788);
or U3964 (N_3964,N_1302,N_1160);
and U3965 (N_3965,N_2112,N_197);
or U3966 (N_3966,N_879,N_2372);
or U3967 (N_3967,N_668,N_448);
nand U3968 (N_3968,N_1332,N_1787);
nand U3969 (N_3969,N_1151,N_719);
nand U3970 (N_3970,N_1740,N_429);
or U3971 (N_3971,N_1662,N_33);
and U3972 (N_3972,N_37,N_831);
nor U3973 (N_3973,N_660,N_2186);
or U3974 (N_3974,N_1744,N_399);
and U3975 (N_3975,N_2330,N_629);
or U3976 (N_3976,N_459,N_1172);
nor U3977 (N_3977,N_2474,N_1330);
nor U3978 (N_3978,N_1271,N_942);
nand U3979 (N_3979,N_642,N_2346);
or U3980 (N_3980,N_1736,N_385);
or U3981 (N_3981,N_404,N_1549);
nor U3982 (N_3982,N_2354,N_1681);
nor U3983 (N_3983,N_2023,N_575);
nor U3984 (N_3984,N_323,N_642);
nor U3985 (N_3985,N_1988,N_110);
or U3986 (N_3986,N_716,N_2176);
nor U3987 (N_3987,N_952,N_1731);
and U3988 (N_3988,N_737,N_283);
nor U3989 (N_3989,N_415,N_2185);
nor U3990 (N_3990,N_272,N_1520);
or U3991 (N_3991,N_462,N_1168);
and U3992 (N_3992,N_1598,N_1813);
nand U3993 (N_3993,N_1437,N_2135);
nor U3994 (N_3994,N_147,N_2076);
nor U3995 (N_3995,N_2074,N_385);
nor U3996 (N_3996,N_889,N_1132);
or U3997 (N_3997,N_268,N_1063);
or U3998 (N_3998,N_2449,N_973);
nor U3999 (N_3999,N_1345,N_1888);
or U4000 (N_4000,N_1016,N_124);
nor U4001 (N_4001,N_1703,N_157);
and U4002 (N_4002,N_1430,N_1929);
and U4003 (N_4003,N_820,N_1403);
or U4004 (N_4004,N_1857,N_155);
or U4005 (N_4005,N_2473,N_763);
nor U4006 (N_4006,N_636,N_1799);
or U4007 (N_4007,N_325,N_837);
nand U4008 (N_4008,N_1881,N_2158);
or U4009 (N_4009,N_237,N_2462);
nor U4010 (N_4010,N_2032,N_919);
nor U4011 (N_4011,N_14,N_1036);
and U4012 (N_4012,N_400,N_1480);
or U4013 (N_4013,N_305,N_1152);
nand U4014 (N_4014,N_0,N_627);
and U4015 (N_4015,N_390,N_2411);
nor U4016 (N_4016,N_2093,N_560);
nor U4017 (N_4017,N_140,N_1777);
nand U4018 (N_4018,N_1147,N_758);
nand U4019 (N_4019,N_1991,N_567);
nor U4020 (N_4020,N_2381,N_1281);
or U4021 (N_4021,N_1775,N_1841);
and U4022 (N_4022,N_1997,N_1785);
and U4023 (N_4023,N_1274,N_2426);
nand U4024 (N_4024,N_2164,N_602);
and U4025 (N_4025,N_818,N_904);
and U4026 (N_4026,N_97,N_1739);
nand U4027 (N_4027,N_1529,N_2081);
or U4028 (N_4028,N_334,N_778);
or U4029 (N_4029,N_5,N_1419);
xor U4030 (N_4030,N_1540,N_2340);
nor U4031 (N_4031,N_1743,N_862);
nor U4032 (N_4032,N_172,N_1085);
and U4033 (N_4033,N_866,N_859);
nor U4034 (N_4034,N_1449,N_320);
and U4035 (N_4035,N_1573,N_185);
nor U4036 (N_4036,N_2475,N_2092);
nand U4037 (N_4037,N_2230,N_1218);
and U4038 (N_4038,N_1486,N_268);
nand U4039 (N_4039,N_258,N_1479);
nand U4040 (N_4040,N_211,N_1872);
nand U4041 (N_4041,N_1485,N_2220);
nor U4042 (N_4042,N_241,N_1146);
nand U4043 (N_4043,N_555,N_1596);
nor U4044 (N_4044,N_2370,N_1606);
and U4045 (N_4045,N_2002,N_781);
nand U4046 (N_4046,N_849,N_496);
and U4047 (N_4047,N_418,N_1836);
nand U4048 (N_4048,N_972,N_1561);
nor U4049 (N_4049,N_1132,N_2420);
nand U4050 (N_4050,N_775,N_675);
or U4051 (N_4051,N_1787,N_2118);
and U4052 (N_4052,N_1655,N_1839);
and U4053 (N_4053,N_1326,N_374);
and U4054 (N_4054,N_1136,N_1241);
and U4055 (N_4055,N_306,N_684);
nand U4056 (N_4056,N_1479,N_748);
or U4057 (N_4057,N_1980,N_867);
or U4058 (N_4058,N_574,N_381);
nand U4059 (N_4059,N_1388,N_906);
nand U4060 (N_4060,N_601,N_646);
nand U4061 (N_4061,N_1441,N_1684);
nand U4062 (N_4062,N_2142,N_2231);
nor U4063 (N_4063,N_339,N_491);
nor U4064 (N_4064,N_1738,N_1680);
nor U4065 (N_4065,N_1974,N_125);
or U4066 (N_4066,N_2339,N_1127);
and U4067 (N_4067,N_565,N_1674);
nand U4068 (N_4068,N_129,N_1039);
and U4069 (N_4069,N_1664,N_26);
nand U4070 (N_4070,N_1680,N_573);
and U4071 (N_4071,N_677,N_1290);
and U4072 (N_4072,N_356,N_1336);
or U4073 (N_4073,N_1461,N_625);
or U4074 (N_4074,N_2158,N_1937);
and U4075 (N_4075,N_2241,N_1170);
and U4076 (N_4076,N_1932,N_2298);
or U4077 (N_4077,N_2075,N_865);
nand U4078 (N_4078,N_1819,N_18);
or U4079 (N_4079,N_1707,N_265);
nor U4080 (N_4080,N_1884,N_1888);
nor U4081 (N_4081,N_384,N_1860);
nand U4082 (N_4082,N_1705,N_183);
and U4083 (N_4083,N_1508,N_158);
nand U4084 (N_4084,N_489,N_110);
xor U4085 (N_4085,N_2279,N_1735);
or U4086 (N_4086,N_2308,N_2465);
nor U4087 (N_4087,N_535,N_551);
nand U4088 (N_4088,N_1426,N_216);
or U4089 (N_4089,N_221,N_1984);
nand U4090 (N_4090,N_1440,N_1471);
nand U4091 (N_4091,N_948,N_2295);
nand U4092 (N_4092,N_737,N_850);
nor U4093 (N_4093,N_1858,N_610);
nand U4094 (N_4094,N_226,N_1179);
nand U4095 (N_4095,N_1705,N_1196);
and U4096 (N_4096,N_945,N_901);
or U4097 (N_4097,N_322,N_2472);
nand U4098 (N_4098,N_1733,N_1434);
or U4099 (N_4099,N_1874,N_1882);
xor U4100 (N_4100,N_380,N_687);
nor U4101 (N_4101,N_846,N_835);
nand U4102 (N_4102,N_870,N_2142);
nor U4103 (N_4103,N_1103,N_2222);
nor U4104 (N_4104,N_2022,N_1240);
nand U4105 (N_4105,N_1706,N_887);
nor U4106 (N_4106,N_767,N_2393);
nand U4107 (N_4107,N_1974,N_841);
nand U4108 (N_4108,N_1187,N_37);
or U4109 (N_4109,N_1763,N_1762);
nand U4110 (N_4110,N_695,N_835);
xor U4111 (N_4111,N_952,N_237);
or U4112 (N_4112,N_2058,N_2441);
or U4113 (N_4113,N_257,N_567);
and U4114 (N_4114,N_1482,N_927);
nand U4115 (N_4115,N_1562,N_1785);
xor U4116 (N_4116,N_648,N_449);
nor U4117 (N_4117,N_2300,N_2167);
and U4118 (N_4118,N_746,N_1599);
nand U4119 (N_4119,N_2352,N_579);
and U4120 (N_4120,N_324,N_1379);
or U4121 (N_4121,N_456,N_1353);
nor U4122 (N_4122,N_2073,N_183);
nand U4123 (N_4123,N_2129,N_1027);
or U4124 (N_4124,N_2000,N_2426);
nand U4125 (N_4125,N_1937,N_874);
and U4126 (N_4126,N_817,N_2344);
or U4127 (N_4127,N_2266,N_1314);
and U4128 (N_4128,N_1556,N_496);
or U4129 (N_4129,N_837,N_1521);
and U4130 (N_4130,N_1163,N_1247);
and U4131 (N_4131,N_248,N_270);
nand U4132 (N_4132,N_1714,N_2468);
nor U4133 (N_4133,N_1767,N_586);
and U4134 (N_4134,N_356,N_1384);
nor U4135 (N_4135,N_1858,N_2436);
and U4136 (N_4136,N_2326,N_607);
nand U4137 (N_4137,N_882,N_665);
or U4138 (N_4138,N_602,N_143);
and U4139 (N_4139,N_551,N_2368);
nand U4140 (N_4140,N_1463,N_2105);
nand U4141 (N_4141,N_1873,N_1841);
and U4142 (N_4142,N_1321,N_322);
nor U4143 (N_4143,N_824,N_603);
or U4144 (N_4144,N_602,N_1040);
or U4145 (N_4145,N_463,N_1341);
nor U4146 (N_4146,N_1249,N_416);
nor U4147 (N_4147,N_2264,N_939);
and U4148 (N_4148,N_1446,N_442);
or U4149 (N_4149,N_111,N_2024);
nand U4150 (N_4150,N_554,N_1034);
or U4151 (N_4151,N_1312,N_1757);
and U4152 (N_4152,N_2148,N_2049);
nor U4153 (N_4153,N_2234,N_86);
or U4154 (N_4154,N_2311,N_1535);
and U4155 (N_4155,N_2493,N_662);
and U4156 (N_4156,N_2011,N_959);
nand U4157 (N_4157,N_504,N_766);
or U4158 (N_4158,N_1437,N_702);
nand U4159 (N_4159,N_465,N_1528);
nor U4160 (N_4160,N_145,N_1052);
and U4161 (N_4161,N_54,N_881);
xor U4162 (N_4162,N_1994,N_1121);
or U4163 (N_4163,N_1495,N_442);
nor U4164 (N_4164,N_326,N_761);
nand U4165 (N_4165,N_2286,N_1390);
or U4166 (N_4166,N_241,N_2054);
nor U4167 (N_4167,N_1859,N_1438);
and U4168 (N_4168,N_1147,N_734);
and U4169 (N_4169,N_1005,N_855);
nand U4170 (N_4170,N_1905,N_1087);
nor U4171 (N_4171,N_375,N_1670);
and U4172 (N_4172,N_938,N_2289);
nor U4173 (N_4173,N_2136,N_2383);
and U4174 (N_4174,N_951,N_695);
or U4175 (N_4175,N_2094,N_831);
and U4176 (N_4176,N_282,N_822);
nor U4177 (N_4177,N_340,N_429);
nand U4178 (N_4178,N_363,N_729);
nor U4179 (N_4179,N_2350,N_1026);
and U4180 (N_4180,N_2493,N_418);
or U4181 (N_4181,N_255,N_970);
or U4182 (N_4182,N_853,N_532);
nor U4183 (N_4183,N_1687,N_1843);
nor U4184 (N_4184,N_654,N_1433);
nor U4185 (N_4185,N_1791,N_353);
xor U4186 (N_4186,N_1227,N_2355);
nor U4187 (N_4187,N_1337,N_1029);
nand U4188 (N_4188,N_1221,N_922);
or U4189 (N_4189,N_534,N_63);
nand U4190 (N_4190,N_1352,N_1032);
and U4191 (N_4191,N_1184,N_1281);
nand U4192 (N_4192,N_43,N_665);
nor U4193 (N_4193,N_1927,N_1962);
or U4194 (N_4194,N_2167,N_1364);
or U4195 (N_4195,N_460,N_1370);
and U4196 (N_4196,N_141,N_1087);
xnor U4197 (N_4197,N_2225,N_2023);
and U4198 (N_4198,N_1656,N_2221);
or U4199 (N_4199,N_213,N_1776);
nor U4200 (N_4200,N_1567,N_1029);
or U4201 (N_4201,N_1398,N_1943);
nand U4202 (N_4202,N_1309,N_1991);
or U4203 (N_4203,N_2481,N_672);
nor U4204 (N_4204,N_2347,N_216);
nand U4205 (N_4205,N_1419,N_1887);
nand U4206 (N_4206,N_639,N_570);
nor U4207 (N_4207,N_53,N_2343);
and U4208 (N_4208,N_2119,N_163);
or U4209 (N_4209,N_190,N_607);
and U4210 (N_4210,N_1342,N_94);
nand U4211 (N_4211,N_383,N_285);
and U4212 (N_4212,N_2499,N_411);
xnor U4213 (N_4213,N_2490,N_1681);
or U4214 (N_4214,N_2002,N_670);
nor U4215 (N_4215,N_2082,N_434);
and U4216 (N_4216,N_498,N_1576);
and U4217 (N_4217,N_2270,N_1009);
or U4218 (N_4218,N_2211,N_31);
xor U4219 (N_4219,N_269,N_1198);
nand U4220 (N_4220,N_1055,N_1771);
or U4221 (N_4221,N_1587,N_1303);
or U4222 (N_4222,N_843,N_1991);
nand U4223 (N_4223,N_303,N_2110);
or U4224 (N_4224,N_2238,N_839);
or U4225 (N_4225,N_1715,N_2204);
and U4226 (N_4226,N_1803,N_50);
and U4227 (N_4227,N_1664,N_2065);
nand U4228 (N_4228,N_623,N_2069);
nor U4229 (N_4229,N_1994,N_97);
and U4230 (N_4230,N_262,N_2456);
and U4231 (N_4231,N_1558,N_1157);
nor U4232 (N_4232,N_1973,N_1902);
and U4233 (N_4233,N_35,N_9);
nor U4234 (N_4234,N_568,N_610);
nand U4235 (N_4235,N_2372,N_1281);
or U4236 (N_4236,N_1064,N_2487);
nor U4237 (N_4237,N_719,N_2266);
or U4238 (N_4238,N_1538,N_1126);
nor U4239 (N_4239,N_264,N_806);
and U4240 (N_4240,N_885,N_911);
nor U4241 (N_4241,N_978,N_1856);
and U4242 (N_4242,N_1319,N_251);
nor U4243 (N_4243,N_2034,N_1854);
and U4244 (N_4244,N_2477,N_1991);
and U4245 (N_4245,N_926,N_2348);
nor U4246 (N_4246,N_243,N_1327);
and U4247 (N_4247,N_14,N_1478);
or U4248 (N_4248,N_1492,N_961);
or U4249 (N_4249,N_917,N_315);
or U4250 (N_4250,N_453,N_2362);
and U4251 (N_4251,N_1167,N_1369);
nor U4252 (N_4252,N_2325,N_16);
nor U4253 (N_4253,N_879,N_2406);
and U4254 (N_4254,N_1501,N_1039);
nor U4255 (N_4255,N_530,N_213);
or U4256 (N_4256,N_2474,N_802);
nand U4257 (N_4257,N_1516,N_1654);
and U4258 (N_4258,N_2018,N_387);
nor U4259 (N_4259,N_236,N_325);
and U4260 (N_4260,N_1859,N_2458);
and U4261 (N_4261,N_793,N_2366);
and U4262 (N_4262,N_2096,N_1841);
nand U4263 (N_4263,N_1113,N_675);
xnor U4264 (N_4264,N_1455,N_966);
nand U4265 (N_4265,N_1444,N_1803);
nand U4266 (N_4266,N_2019,N_1800);
nand U4267 (N_4267,N_317,N_2395);
nor U4268 (N_4268,N_508,N_1035);
or U4269 (N_4269,N_2149,N_1546);
and U4270 (N_4270,N_887,N_324);
nor U4271 (N_4271,N_914,N_134);
nand U4272 (N_4272,N_649,N_1510);
nand U4273 (N_4273,N_1046,N_2198);
and U4274 (N_4274,N_467,N_536);
and U4275 (N_4275,N_201,N_1192);
and U4276 (N_4276,N_204,N_391);
nand U4277 (N_4277,N_134,N_1671);
or U4278 (N_4278,N_1265,N_2418);
nand U4279 (N_4279,N_1050,N_1688);
nor U4280 (N_4280,N_113,N_1944);
nor U4281 (N_4281,N_651,N_1120);
and U4282 (N_4282,N_368,N_2010);
or U4283 (N_4283,N_1180,N_234);
or U4284 (N_4284,N_1237,N_1936);
and U4285 (N_4285,N_1902,N_2336);
nor U4286 (N_4286,N_140,N_1550);
or U4287 (N_4287,N_604,N_2201);
or U4288 (N_4288,N_2261,N_1357);
nor U4289 (N_4289,N_664,N_2084);
nand U4290 (N_4290,N_1594,N_239);
nor U4291 (N_4291,N_1021,N_1104);
nor U4292 (N_4292,N_2325,N_609);
or U4293 (N_4293,N_485,N_549);
and U4294 (N_4294,N_1237,N_380);
or U4295 (N_4295,N_100,N_1657);
and U4296 (N_4296,N_382,N_1502);
and U4297 (N_4297,N_1405,N_1166);
and U4298 (N_4298,N_1043,N_1227);
or U4299 (N_4299,N_1842,N_316);
or U4300 (N_4300,N_1452,N_737);
and U4301 (N_4301,N_506,N_1606);
and U4302 (N_4302,N_2159,N_794);
nor U4303 (N_4303,N_2362,N_2205);
and U4304 (N_4304,N_2086,N_2022);
nor U4305 (N_4305,N_1034,N_645);
nand U4306 (N_4306,N_364,N_193);
or U4307 (N_4307,N_441,N_2070);
xor U4308 (N_4308,N_1436,N_449);
nand U4309 (N_4309,N_1239,N_1230);
nor U4310 (N_4310,N_1310,N_1232);
or U4311 (N_4311,N_1562,N_2021);
nor U4312 (N_4312,N_1525,N_1612);
xor U4313 (N_4313,N_1641,N_1599);
or U4314 (N_4314,N_1077,N_1855);
nand U4315 (N_4315,N_230,N_1156);
nand U4316 (N_4316,N_2404,N_2482);
or U4317 (N_4317,N_423,N_766);
or U4318 (N_4318,N_1328,N_1500);
or U4319 (N_4319,N_750,N_292);
xnor U4320 (N_4320,N_2334,N_2408);
xor U4321 (N_4321,N_1160,N_873);
nor U4322 (N_4322,N_1861,N_464);
nand U4323 (N_4323,N_1328,N_112);
or U4324 (N_4324,N_2157,N_1506);
or U4325 (N_4325,N_88,N_2325);
nor U4326 (N_4326,N_508,N_603);
and U4327 (N_4327,N_2455,N_1260);
nor U4328 (N_4328,N_2424,N_94);
nand U4329 (N_4329,N_724,N_1199);
and U4330 (N_4330,N_1185,N_918);
nor U4331 (N_4331,N_1221,N_1745);
and U4332 (N_4332,N_2452,N_2039);
nor U4333 (N_4333,N_385,N_1248);
or U4334 (N_4334,N_878,N_395);
or U4335 (N_4335,N_431,N_1406);
or U4336 (N_4336,N_1445,N_2432);
nand U4337 (N_4337,N_440,N_2155);
nor U4338 (N_4338,N_999,N_1912);
and U4339 (N_4339,N_2371,N_2453);
and U4340 (N_4340,N_518,N_465);
nand U4341 (N_4341,N_1371,N_1945);
and U4342 (N_4342,N_1609,N_1864);
or U4343 (N_4343,N_247,N_1057);
nand U4344 (N_4344,N_701,N_1216);
nor U4345 (N_4345,N_762,N_1371);
or U4346 (N_4346,N_839,N_2409);
nand U4347 (N_4347,N_2127,N_727);
nor U4348 (N_4348,N_1046,N_1601);
nor U4349 (N_4349,N_1972,N_1204);
or U4350 (N_4350,N_233,N_1786);
and U4351 (N_4351,N_1140,N_103);
or U4352 (N_4352,N_94,N_1395);
nand U4353 (N_4353,N_1476,N_1079);
nor U4354 (N_4354,N_1668,N_63);
or U4355 (N_4355,N_247,N_1957);
xor U4356 (N_4356,N_1808,N_2346);
and U4357 (N_4357,N_875,N_607);
or U4358 (N_4358,N_62,N_771);
nand U4359 (N_4359,N_721,N_274);
or U4360 (N_4360,N_1517,N_1834);
nor U4361 (N_4361,N_1534,N_1779);
nand U4362 (N_4362,N_1996,N_682);
or U4363 (N_4363,N_816,N_739);
nand U4364 (N_4364,N_2103,N_0);
nand U4365 (N_4365,N_2361,N_1498);
nand U4366 (N_4366,N_1121,N_1031);
and U4367 (N_4367,N_1034,N_166);
nor U4368 (N_4368,N_939,N_1463);
or U4369 (N_4369,N_1330,N_1326);
and U4370 (N_4370,N_812,N_291);
or U4371 (N_4371,N_2135,N_1033);
or U4372 (N_4372,N_280,N_991);
or U4373 (N_4373,N_2215,N_287);
or U4374 (N_4374,N_1940,N_2212);
nand U4375 (N_4375,N_2380,N_1302);
or U4376 (N_4376,N_2295,N_279);
and U4377 (N_4377,N_2472,N_1394);
nand U4378 (N_4378,N_398,N_2208);
nand U4379 (N_4379,N_372,N_195);
or U4380 (N_4380,N_228,N_2082);
nand U4381 (N_4381,N_327,N_562);
nand U4382 (N_4382,N_1921,N_764);
nand U4383 (N_4383,N_2379,N_1210);
nand U4384 (N_4384,N_2032,N_714);
or U4385 (N_4385,N_522,N_2350);
or U4386 (N_4386,N_1943,N_1867);
xnor U4387 (N_4387,N_2487,N_2396);
and U4388 (N_4388,N_1996,N_687);
or U4389 (N_4389,N_224,N_2165);
and U4390 (N_4390,N_198,N_1999);
nand U4391 (N_4391,N_862,N_332);
nor U4392 (N_4392,N_346,N_2491);
nand U4393 (N_4393,N_1985,N_511);
nor U4394 (N_4394,N_1401,N_912);
or U4395 (N_4395,N_1796,N_143);
and U4396 (N_4396,N_289,N_1743);
nand U4397 (N_4397,N_481,N_965);
nand U4398 (N_4398,N_160,N_528);
or U4399 (N_4399,N_1914,N_939);
and U4400 (N_4400,N_1471,N_879);
nor U4401 (N_4401,N_494,N_1801);
and U4402 (N_4402,N_1208,N_956);
nor U4403 (N_4403,N_1574,N_1192);
xor U4404 (N_4404,N_277,N_612);
and U4405 (N_4405,N_53,N_1234);
nand U4406 (N_4406,N_2073,N_1162);
nor U4407 (N_4407,N_557,N_1624);
nand U4408 (N_4408,N_629,N_848);
nand U4409 (N_4409,N_665,N_2092);
or U4410 (N_4410,N_2492,N_299);
and U4411 (N_4411,N_2332,N_1573);
or U4412 (N_4412,N_1135,N_2187);
and U4413 (N_4413,N_1481,N_1008);
and U4414 (N_4414,N_1591,N_1156);
and U4415 (N_4415,N_1250,N_1337);
nand U4416 (N_4416,N_395,N_1962);
nand U4417 (N_4417,N_2116,N_1016);
nor U4418 (N_4418,N_272,N_81);
nor U4419 (N_4419,N_260,N_2494);
or U4420 (N_4420,N_154,N_1737);
nor U4421 (N_4421,N_74,N_519);
and U4422 (N_4422,N_1549,N_1890);
nand U4423 (N_4423,N_2401,N_1495);
nand U4424 (N_4424,N_2265,N_1136);
nand U4425 (N_4425,N_180,N_713);
xor U4426 (N_4426,N_1908,N_448);
nor U4427 (N_4427,N_412,N_2434);
and U4428 (N_4428,N_2239,N_32);
nand U4429 (N_4429,N_2225,N_2489);
or U4430 (N_4430,N_1737,N_1178);
or U4431 (N_4431,N_1822,N_1450);
or U4432 (N_4432,N_427,N_440);
and U4433 (N_4433,N_953,N_1190);
nand U4434 (N_4434,N_985,N_1650);
nand U4435 (N_4435,N_1356,N_356);
nor U4436 (N_4436,N_1310,N_2068);
nor U4437 (N_4437,N_272,N_502);
or U4438 (N_4438,N_357,N_2045);
nor U4439 (N_4439,N_248,N_859);
or U4440 (N_4440,N_413,N_1562);
or U4441 (N_4441,N_1582,N_2316);
and U4442 (N_4442,N_414,N_814);
nand U4443 (N_4443,N_2309,N_1149);
nor U4444 (N_4444,N_1161,N_1278);
nand U4445 (N_4445,N_902,N_2283);
or U4446 (N_4446,N_1878,N_2436);
and U4447 (N_4447,N_1490,N_1665);
or U4448 (N_4448,N_388,N_847);
nor U4449 (N_4449,N_562,N_2107);
nor U4450 (N_4450,N_798,N_38);
nand U4451 (N_4451,N_2312,N_249);
nand U4452 (N_4452,N_2244,N_2336);
nand U4453 (N_4453,N_1255,N_433);
nand U4454 (N_4454,N_1128,N_503);
nand U4455 (N_4455,N_903,N_694);
nand U4456 (N_4456,N_502,N_617);
or U4457 (N_4457,N_1197,N_102);
or U4458 (N_4458,N_2277,N_785);
nor U4459 (N_4459,N_2204,N_371);
or U4460 (N_4460,N_1784,N_303);
and U4461 (N_4461,N_185,N_457);
nor U4462 (N_4462,N_1673,N_599);
xor U4463 (N_4463,N_982,N_1993);
nor U4464 (N_4464,N_2016,N_1669);
or U4465 (N_4465,N_741,N_1605);
nor U4466 (N_4466,N_563,N_1665);
or U4467 (N_4467,N_1629,N_1359);
xor U4468 (N_4468,N_1722,N_1023);
and U4469 (N_4469,N_2080,N_708);
nand U4470 (N_4470,N_742,N_2070);
nand U4471 (N_4471,N_1038,N_99);
or U4472 (N_4472,N_56,N_1103);
or U4473 (N_4473,N_339,N_207);
xor U4474 (N_4474,N_221,N_163);
and U4475 (N_4475,N_1972,N_1878);
nand U4476 (N_4476,N_1922,N_267);
or U4477 (N_4477,N_1936,N_2196);
nor U4478 (N_4478,N_68,N_97);
and U4479 (N_4479,N_368,N_1221);
and U4480 (N_4480,N_1174,N_535);
or U4481 (N_4481,N_76,N_1399);
nor U4482 (N_4482,N_109,N_792);
nand U4483 (N_4483,N_734,N_2242);
nor U4484 (N_4484,N_2302,N_2491);
nor U4485 (N_4485,N_1373,N_1359);
and U4486 (N_4486,N_1688,N_1763);
xnor U4487 (N_4487,N_1643,N_2407);
xnor U4488 (N_4488,N_779,N_2458);
nand U4489 (N_4489,N_1612,N_643);
nand U4490 (N_4490,N_528,N_1832);
or U4491 (N_4491,N_1147,N_1220);
xnor U4492 (N_4492,N_1160,N_2439);
nor U4493 (N_4493,N_918,N_875);
and U4494 (N_4494,N_1736,N_1473);
xor U4495 (N_4495,N_325,N_826);
or U4496 (N_4496,N_968,N_2407);
and U4497 (N_4497,N_139,N_285);
nor U4498 (N_4498,N_279,N_700);
nand U4499 (N_4499,N_238,N_894);
or U4500 (N_4500,N_421,N_194);
and U4501 (N_4501,N_1013,N_502);
nand U4502 (N_4502,N_653,N_1855);
or U4503 (N_4503,N_1946,N_27);
and U4504 (N_4504,N_241,N_1566);
and U4505 (N_4505,N_975,N_806);
nor U4506 (N_4506,N_1872,N_2338);
or U4507 (N_4507,N_1282,N_2490);
nand U4508 (N_4508,N_164,N_909);
nor U4509 (N_4509,N_2182,N_1643);
nand U4510 (N_4510,N_2269,N_1192);
nor U4511 (N_4511,N_1637,N_2411);
or U4512 (N_4512,N_1853,N_998);
or U4513 (N_4513,N_541,N_457);
nor U4514 (N_4514,N_842,N_272);
or U4515 (N_4515,N_1650,N_2498);
nand U4516 (N_4516,N_1617,N_927);
nand U4517 (N_4517,N_911,N_1110);
nand U4518 (N_4518,N_2214,N_1413);
or U4519 (N_4519,N_2178,N_78);
nor U4520 (N_4520,N_1529,N_556);
or U4521 (N_4521,N_327,N_466);
nor U4522 (N_4522,N_714,N_1196);
nor U4523 (N_4523,N_1141,N_273);
nand U4524 (N_4524,N_162,N_1808);
or U4525 (N_4525,N_326,N_1062);
and U4526 (N_4526,N_205,N_1250);
or U4527 (N_4527,N_2474,N_447);
nor U4528 (N_4528,N_2226,N_2051);
and U4529 (N_4529,N_1933,N_1979);
nor U4530 (N_4530,N_2319,N_2340);
nor U4531 (N_4531,N_2391,N_722);
and U4532 (N_4532,N_521,N_918);
nor U4533 (N_4533,N_1968,N_2083);
and U4534 (N_4534,N_2357,N_1321);
and U4535 (N_4535,N_608,N_1054);
or U4536 (N_4536,N_923,N_2446);
or U4537 (N_4537,N_1889,N_519);
or U4538 (N_4538,N_1042,N_1315);
nor U4539 (N_4539,N_1247,N_22);
nand U4540 (N_4540,N_1149,N_1479);
and U4541 (N_4541,N_2045,N_747);
and U4542 (N_4542,N_163,N_2486);
and U4543 (N_4543,N_2322,N_1903);
and U4544 (N_4544,N_54,N_1614);
nor U4545 (N_4545,N_887,N_2162);
xnor U4546 (N_4546,N_2438,N_1779);
and U4547 (N_4547,N_176,N_1152);
nand U4548 (N_4548,N_260,N_953);
or U4549 (N_4549,N_900,N_5);
nor U4550 (N_4550,N_1661,N_2268);
and U4551 (N_4551,N_451,N_1306);
nor U4552 (N_4552,N_498,N_2095);
and U4553 (N_4553,N_556,N_2132);
and U4554 (N_4554,N_615,N_1934);
nor U4555 (N_4555,N_2056,N_683);
or U4556 (N_4556,N_502,N_889);
and U4557 (N_4557,N_1197,N_380);
and U4558 (N_4558,N_2057,N_546);
nand U4559 (N_4559,N_849,N_176);
and U4560 (N_4560,N_2004,N_1681);
xor U4561 (N_4561,N_2405,N_14);
nand U4562 (N_4562,N_248,N_267);
and U4563 (N_4563,N_2481,N_2421);
and U4564 (N_4564,N_1992,N_1523);
nand U4565 (N_4565,N_1780,N_378);
nor U4566 (N_4566,N_1710,N_573);
or U4567 (N_4567,N_30,N_3);
and U4568 (N_4568,N_2376,N_1647);
or U4569 (N_4569,N_1784,N_1857);
nand U4570 (N_4570,N_1358,N_377);
nand U4571 (N_4571,N_1381,N_21);
and U4572 (N_4572,N_1880,N_1713);
xor U4573 (N_4573,N_1155,N_143);
or U4574 (N_4574,N_2173,N_888);
or U4575 (N_4575,N_468,N_2282);
nor U4576 (N_4576,N_1353,N_879);
or U4577 (N_4577,N_763,N_1077);
and U4578 (N_4578,N_1403,N_133);
or U4579 (N_4579,N_1141,N_1397);
xor U4580 (N_4580,N_2408,N_1120);
nand U4581 (N_4581,N_1278,N_327);
nor U4582 (N_4582,N_156,N_1336);
xor U4583 (N_4583,N_1593,N_1054);
or U4584 (N_4584,N_1942,N_80);
and U4585 (N_4585,N_293,N_55);
xor U4586 (N_4586,N_578,N_2221);
nand U4587 (N_4587,N_1725,N_2386);
nor U4588 (N_4588,N_207,N_1007);
nand U4589 (N_4589,N_567,N_1039);
nand U4590 (N_4590,N_1312,N_958);
and U4591 (N_4591,N_2319,N_2145);
nor U4592 (N_4592,N_228,N_544);
or U4593 (N_4593,N_1950,N_1937);
nor U4594 (N_4594,N_1262,N_48);
or U4595 (N_4595,N_521,N_316);
nand U4596 (N_4596,N_293,N_739);
nand U4597 (N_4597,N_1816,N_1698);
and U4598 (N_4598,N_1074,N_1362);
or U4599 (N_4599,N_1506,N_1684);
nor U4600 (N_4600,N_2001,N_2027);
and U4601 (N_4601,N_1203,N_1055);
nor U4602 (N_4602,N_1003,N_2096);
nor U4603 (N_4603,N_1076,N_2463);
and U4604 (N_4604,N_561,N_1657);
xor U4605 (N_4605,N_1353,N_328);
and U4606 (N_4606,N_2323,N_22);
or U4607 (N_4607,N_772,N_1571);
or U4608 (N_4608,N_2199,N_2065);
nand U4609 (N_4609,N_1115,N_394);
or U4610 (N_4610,N_1853,N_1176);
or U4611 (N_4611,N_1353,N_1202);
nand U4612 (N_4612,N_1346,N_1510);
or U4613 (N_4613,N_2406,N_1235);
and U4614 (N_4614,N_123,N_1216);
nor U4615 (N_4615,N_323,N_2382);
and U4616 (N_4616,N_2487,N_1039);
nand U4617 (N_4617,N_1346,N_2096);
or U4618 (N_4618,N_2485,N_1392);
nand U4619 (N_4619,N_2316,N_1462);
or U4620 (N_4620,N_2307,N_942);
nor U4621 (N_4621,N_1560,N_134);
or U4622 (N_4622,N_610,N_597);
and U4623 (N_4623,N_1755,N_1508);
nor U4624 (N_4624,N_266,N_776);
or U4625 (N_4625,N_1266,N_664);
or U4626 (N_4626,N_291,N_2223);
or U4627 (N_4627,N_2137,N_164);
or U4628 (N_4628,N_16,N_1179);
xnor U4629 (N_4629,N_1079,N_1581);
and U4630 (N_4630,N_153,N_1614);
and U4631 (N_4631,N_1277,N_1211);
and U4632 (N_4632,N_2177,N_1908);
and U4633 (N_4633,N_672,N_883);
nor U4634 (N_4634,N_2361,N_2234);
and U4635 (N_4635,N_1105,N_1985);
nand U4636 (N_4636,N_2389,N_705);
nand U4637 (N_4637,N_789,N_2035);
or U4638 (N_4638,N_1627,N_17);
or U4639 (N_4639,N_1052,N_612);
xnor U4640 (N_4640,N_2026,N_849);
and U4641 (N_4641,N_663,N_2246);
or U4642 (N_4642,N_2260,N_2132);
nand U4643 (N_4643,N_2130,N_858);
and U4644 (N_4644,N_176,N_1838);
and U4645 (N_4645,N_1217,N_1679);
and U4646 (N_4646,N_1843,N_257);
nor U4647 (N_4647,N_1839,N_2471);
and U4648 (N_4648,N_1054,N_1444);
or U4649 (N_4649,N_1824,N_110);
nor U4650 (N_4650,N_950,N_43);
nand U4651 (N_4651,N_1332,N_548);
and U4652 (N_4652,N_1716,N_1004);
nand U4653 (N_4653,N_1706,N_2439);
nand U4654 (N_4654,N_724,N_1045);
nor U4655 (N_4655,N_841,N_1586);
or U4656 (N_4656,N_1503,N_510);
nand U4657 (N_4657,N_1883,N_1262);
nor U4658 (N_4658,N_1546,N_1341);
nor U4659 (N_4659,N_446,N_1149);
nand U4660 (N_4660,N_103,N_1388);
nor U4661 (N_4661,N_400,N_343);
nand U4662 (N_4662,N_1734,N_2401);
and U4663 (N_4663,N_1228,N_2144);
or U4664 (N_4664,N_943,N_319);
or U4665 (N_4665,N_1289,N_2012);
nand U4666 (N_4666,N_865,N_17);
xnor U4667 (N_4667,N_1786,N_1230);
and U4668 (N_4668,N_820,N_480);
or U4669 (N_4669,N_625,N_439);
nor U4670 (N_4670,N_2298,N_2402);
nor U4671 (N_4671,N_1309,N_763);
nand U4672 (N_4672,N_2050,N_407);
nand U4673 (N_4673,N_226,N_1715);
or U4674 (N_4674,N_1368,N_108);
or U4675 (N_4675,N_404,N_2483);
nor U4676 (N_4676,N_488,N_1364);
or U4677 (N_4677,N_2498,N_2386);
or U4678 (N_4678,N_1101,N_1178);
nand U4679 (N_4679,N_2323,N_2310);
nand U4680 (N_4680,N_14,N_1798);
nand U4681 (N_4681,N_2011,N_864);
or U4682 (N_4682,N_604,N_2265);
and U4683 (N_4683,N_2457,N_1315);
nor U4684 (N_4684,N_1026,N_1526);
nor U4685 (N_4685,N_1232,N_2008);
nor U4686 (N_4686,N_568,N_523);
nor U4687 (N_4687,N_1846,N_2435);
or U4688 (N_4688,N_2086,N_1155);
and U4689 (N_4689,N_1950,N_335);
and U4690 (N_4690,N_2197,N_1118);
and U4691 (N_4691,N_1649,N_2238);
nor U4692 (N_4692,N_81,N_1925);
nand U4693 (N_4693,N_1381,N_685);
and U4694 (N_4694,N_765,N_1328);
or U4695 (N_4695,N_1073,N_932);
or U4696 (N_4696,N_103,N_1112);
and U4697 (N_4697,N_2297,N_1773);
nand U4698 (N_4698,N_1045,N_54);
or U4699 (N_4699,N_1749,N_61);
and U4700 (N_4700,N_1371,N_750);
nor U4701 (N_4701,N_701,N_577);
nor U4702 (N_4702,N_274,N_502);
nand U4703 (N_4703,N_308,N_1413);
nor U4704 (N_4704,N_2196,N_2043);
or U4705 (N_4705,N_1306,N_865);
or U4706 (N_4706,N_235,N_652);
and U4707 (N_4707,N_46,N_240);
nand U4708 (N_4708,N_1199,N_1693);
or U4709 (N_4709,N_484,N_2135);
or U4710 (N_4710,N_633,N_491);
nor U4711 (N_4711,N_2211,N_950);
xnor U4712 (N_4712,N_1766,N_765);
nor U4713 (N_4713,N_782,N_1627);
nand U4714 (N_4714,N_1310,N_2404);
nand U4715 (N_4715,N_2475,N_409);
or U4716 (N_4716,N_39,N_57);
or U4717 (N_4717,N_1897,N_1530);
nand U4718 (N_4718,N_498,N_1080);
or U4719 (N_4719,N_1120,N_294);
or U4720 (N_4720,N_352,N_1157);
and U4721 (N_4721,N_2124,N_462);
or U4722 (N_4722,N_1875,N_2321);
nand U4723 (N_4723,N_1746,N_288);
and U4724 (N_4724,N_1163,N_1039);
nor U4725 (N_4725,N_527,N_2217);
and U4726 (N_4726,N_472,N_2375);
and U4727 (N_4727,N_719,N_222);
nor U4728 (N_4728,N_1993,N_851);
or U4729 (N_4729,N_2384,N_1936);
or U4730 (N_4730,N_1414,N_836);
nor U4731 (N_4731,N_2315,N_792);
nand U4732 (N_4732,N_1481,N_1963);
nand U4733 (N_4733,N_1041,N_1460);
or U4734 (N_4734,N_674,N_978);
nand U4735 (N_4735,N_1370,N_2213);
xor U4736 (N_4736,N_2230,N_17);
or U4737 (N_4737,N_411,N_1759);
and U4738 (N_4738,N_1559,N_2291);
nor U4739 (N_4739,N_1998,N_1258);
and U4740 (N_4740,N_1379,N_2350);
and U4741 (N_4741,N_1065,N_830);
or U4742 (N_4742,N_2464,N_1361);
nand U4743 (N_4743,N_1911,N_1876);
nor U4744 (N_4744,N_1073,N_228);
nand U4745 (N_4745,N_320,N_1368);
xor U4746 (N_4746,N_245,N_502);
nor U4747 (N_4747,N_1281,N_4);
or U4748 (N_4748,N_690,N_1655);
nor U4749 (N_4749,N_2189,N_2483);
nand U4750 (N_4750,N_1721,N_484);
or U4751 (N_4751,N_1680,N_1658);
nand U4752 (N_4752,N_1621,N_1289);
or U4753 (N_4753,N_176,N_1310);
xor U4754 (N_4754,N_193,N_1771);
xor U4755 (N_4755,N_2152,N_173);
nor U4756 (N_4756,N_1648,N_1132);
or U4757 (N_4757,N_1395,N_1138);
or U4758 (N_4758,N_1994,N_1133);
or U4759 (N_4759,N_2009,N_641);
or U4760 (N_4760,N_2294,N_1798);
nor U4761 (N_4761,N_639,N_263);
or U4762 (N_4762,N_2105,N_43);
and U4763 (N_4763,N_1275,N_852);
and U4764 (N_4764,N_1243,N_997);
and U4765 (N_4765,N_2056,N_1926);
or U4766 (N_4766,N_1915,N_1793);
xnor U4767 (N_4767,N_2428,N_1656);
nand U4768 (N_4768,N_2343,N_599);
or U4769 (N_4769,N_1049,N_745);
and U4770 (N_4770,N_911,N_609);
nor U4771 (N_4771,N_1281,N_363);
and U4772 (N_4772,N_1439,N_1387);
nor U4773 (N_4773,N_2279,N_1612);
and U4774 (N_4774,N_840,N_1781);
or U4775 (N_4775,N_822,N_460);
and U4776 (N_4776,N_2159,N_887);
and U4777 (N_4777,N_2050,N_1623);
nor U4778 (N_4778,N_2364,N_894);
nand U4779 (N_4779,N_448,N_1030);
xor U4780 (N_4780,N_2055,N_811);
or U4781 (N_4781,N_1703,N_890);
and U4782 (N_4782,N_849,N_829);
nand U4783 (N_4783,N_206,N_1978);
and U4784 (N_4784,N_2152,N_627);
nor U4785 (N_4785,N_84,N_125);
or U4786 (N_4786,N_1598,N_1811);
nor U4787 (N_4787,N_285,N_322);
nand U4788 (N_4788,N_1617,N_370);
nor U4789 (N_4789,N_1839,N_1753);
nor U4790 (N_4790,N_1422,N_579);
nand U4791 (N_4791,N_1977,N_2283);
or U4792 (N_4792,N_1008,N_507);
nand U4793 (N_4793,N_1926,N_207);
and U4794 (N_4794,N_1015,N_1535);
nor U4795 (N_4795,N_2358,N_2081);
nand U4796 (N_4796,N_2102,N_1637);
nand U4797 (N_4797,N_1482,N_2390);
or U4798 (N_4798,N_798,N_490);
nand U4799 (N_4799,N_1073,N_110);
or U4800 (N_4800,N_1996,N_2369);
or U4801 (N_4801,N_2373,N_220);
and U4802 (N_4802,N_140,N_2113);
nand U4803 (N_4803,N_1584,N_855);
and U4804 (N_4804,N_2322,N_547);
and U4805 (N_4805,N_576,N_1337);
and U4806 (N_4806,N_1025,N_1371);
or U4807 (N_4807,N_518,N_254);
nor U4808 (N_4808,N_819,N_1340);
nand U4809 (N_4809,N_467,N_2107);
nand U4810 (N_4810,N_677,N_240);
nor U4811 (N_4811,N_871,N_923);
nor U4812 (N_4812,N_583,N_405);
nand U4813 (N_4813,N_653,N_777);
and U4814 (N_4814,N_2006,N_1851);
or U4815 (N_4815,N_702,N_1241);
or U4816 (N_4816,N_1184,N_1621);
and U4817 (N_4817,N_1097,N_1812);
or U4818 (N_4818,N_236,N_2268);
or U4819 (N_4819,N_2148,N_1780);
nand U4820 (N_4820,N_1295,N_1183);
nand U4821 (N_4821,N_1881,N_1756);
nand U4822 (N_4822,N_2408,N_2489);
nand U4823 (N_4823,N_1685,N_1989);
nand U4824 (N_4824,N_283,N_733);
or U4825 (N_4825,N_171,N_1837);
nor U4826 (N_4826,N_1038,N_597);
nand U4827 (N_4827,N_1166,N_1750);
and U4828 (N_4828,N_1031,N_1021);
nor U4829 (N_4829,N_1295,N_516);
nor U4830 (N_4830,N_169,N_662);
and U4831 (N_4831,N_1589,N_115);
xnor U4832 (N_4832,N_1780,N_2414);
nand U4833 (N_4833,N_2401,N_17);
nor U4834 (N_4834,N_908,N_733);
nand U4835 (N_4835,N_2087,N_2210);
and U4836 (N_4836,N_368,N_1563);
or U4837 (N_4837,N_1497,N_701);
nor U4838 (N_4838,N_51,N_769);
nand U4839 (N_4839,N_1144,N_769);
or U4840 (N_4840,N_2239,N_679);
nor U4841 (N_4841,N_1761,N_1668);
nand U4842 (N_4842,N_2103,N_1304);
nand U4843 (N_4843,N_952,N_62);
nand U4844 (N_4844,N_1933,N_2048);
nor U4845 (N_4845,N_2167,N_2319);
or U4846 (N_4846,N_326,N_1069);
nand U4847 (N_4847,N_261,N_292);
nor U4848 (N_4848,N_1621,N_2010);
nor U4849 (N_4849,N_988,N_1665);
nand U4850 (N_4850,N_2195,N_1733);
or U4851 (N_4851,N_305,N_1821);
and U4852 (N_4852,N_778,N_740);
nor U4853 (N_4853,N_1924,N_1132);
and U4854 (N_4854,N_1152,N_2320);
nor U4855 (N_4855,N_1755,N_472);
and U4856 (N_4856,N_814,N_712);
nand U4857 (N_4857,N_692,N_2243);
and U4858 (N_4858,N_1480,N_909);
nand U4859 (N_4859,N_1982,N_218);
and U4860 (N_4860,N_1238,N_221);
nor U4861 (N_4861,N_263,N_768);
nor U4862 (N_4862,N_530,N_470);
nor U4863 (N_4863,N_1630,N_2090);
or U4864 (N_4864,N_2015,N_2184);
nand U4865 (N_4865,N_2114,N_859);
and U4866 (N_4866,N_808,N_1685);
nand U4867 (N_4867,N_639,N_344);
or U4868 (N_4868,N_1588,N_2461);
or U4869 (N_4869,N_1943,N_1410);
and U4870 (N_4870,N_1603,N_2337);
or U4871 (N_4871,N_1359,N_1166);
nand U4872 (N_4872,N_2367,N_249);
nor U4873 (N_4873,N_1962,N_1726);
and U4874 (N_4874,N_1933,N_1842);
nor U4875 (N_4875,N_1094,N_375);
and U4876 (N_4876,N_797,N_1051);
nand U4877 (N_4877,N_1648,N_2123);
or U4878 (N_4878,N_562,N_900);
nand U4879 (N_4879,N_2244,N_1696);
or U4880 (N_4880,N_907,N_668);
or U4881 (N_4881,N_1937,N_1612);
nand U4882 (N_4882,N_1152,N_1047);
nand U4883 (N_4883,N_342,N_1530);
or U4884 (N_4884,N_1077,N_1257);
and U4885 (N_4885,N_1360,N_2401);
nand U4886 (N_4886,N_1037,N_1080);
nand U4887 (N_4887,N_445,N_1648);
nand U4888 (N_4888,N_2486,N_770);
nand U4889 (N_4889,N_1406,N_897);
nor U4890 (N_4890,N_239,N_26);
nor U4891 (N_4891,N_860,N_2218);
nand U4892 (N_4892,N_339,N_2164);
and U4893 (N_4893,N_1214,N_1788);
nor U4894 (N_4894,N_2386,N_508);
or U4895 (N_4895,N_2212,N_2354);
or U4896 (N_4896,N_878,N_1064);
nor U4897 (N_4897,N_1221,N_1162);
nor U4898 (N_4898,N_965,N_636);
or U4899 (N_4899,N_1148,N_350);
or U4900 (N_4900,N_97,N_1265);
nor U4901 (N_4901,N_833,N_584);
and U4902 (N_4902,N_1722,N_1969);
nand U4903 (N_4903,N_2318,N_172);
nand U4904 (N_4904,N_1645,N_1292);
nor U4905 (N_4905,N_2488,N_1317);
and U4906 (N_4906,N_725,N_696);
nor U4907 (N_4907,N_1011,N_1266);
nand U4908 (N_4908,N_2462,N_1290);
nand U4909 (N_4909,N_2493,N_527);
nand U4910 (N_4910,N_2257,N_1537);
nand U4911 (N_4911,N_863,N_134);
nand U4912 (N_4912,N_363,N_1411);
or U4913 (N_4913,N_1035,N_1214);
or U4914 (N_4914,N_962,N_1554);
nor U4915 (N_4915,N_389,N_1054);
nor U4916 (N_4916,N_1035,N_2252);
and U4917 (N_4917,N_850,N_379);
nor U4918 (N_4918,N_2125,N_496);
nand U4919 (N_4919,N_1398,N_1949);
and U4920 (N_4920,N_301,N_1396);
or U4921 (N_4921,N_1131,N_157);
nand U4922 (N_4922,N_925,N_1505);
or U4923 (N_4923,N_652,N_622);
or U4924 (N_4924,N_1024,N_2047);
or U4925 (N_4925,N_2392,N_2175);
nor U4926 (N_4926,N_255,N_2007);
nor U4927 (N_4927,N_2372,N_1537);
nor U4928 (N_4928,N_279,N_1221);
nor U4929 (N_4929,N_2425,N_2439);
nor U4930 (N_4930,N_335,N_1672);
or U4931 (N_4931,N_1800,N_347);
and U4932 (N_4932,N_901,N_1762);
and U4933 (N_4933,N_2427,N_146);
or U4934 (N_4934,N_1288,N_637);
nand U4935 (N_4935,N_1806,N_650);
and U4936 (N_4936,N_156,N_2163);
nor U4937 (N_4937,N_2375,N_1955);
nand U4938 (N_4938,N_841,N_2104);
nand U4939 (N_4939,N_1604,N_1907);
or U4940 (N_4940,N_751,N_1064);
or U4941 (N_4941,N_2421,N_1712);
and U4942 (N_4942,N_135,N_1889);
or U4943 (N_4943,N_1404,N_810);
or U4944 (N_4944,N_1551,N_1468);
nand U4945 (N_4945,N_77,N_1534);
nor U4946 (N_4946,N_1742,N_229);
and U4947 (N_4947,N_1296,N_0);
or U4948 (N_4948,N_1348,N_1565);
or U4949 (N_4949,N_2125,N_1765);
nand U4950 (N_4950,N_1360,N_1847);
and U4951 (N_4951,N_1351,N_291);
and U4952 (N_4952,N_828,N_938);
nor U4953 (N_4953,N_1057,N_710);
nor U4954 (N_4954,N_1729,N_1676);
nand U4955 (N_4955,N_1008,N_1982);
nor U4956 (N_4956,N_972,N_1228);
or U4957 (N_4957,N_1680,N_1386);
nand U4958 (N_4958,N_125,N_2066);
nand U4959 (N_4959,N_1641,N_1004);
xnor U4960 (N_4960,N_127,N_1539);
nor U4961 (N_4961,N_1844,N_1793);
or U4962 (N_4962,N_1825,N_1833);
or U4963 (N_4963,N_1616,N_1486);
nand U4964 (N_4964,N_446,N_1065);
nand U4965 (N_4965,N_2314,N_929);
nor U4966 (N_4966,N_2450,N_1272);
and U4967 (N_4967,N_3,N_206);
nand U4968 (N_4968,N_1702,N_470);
and U4969 (N_4969,N_478,N_1679);
or U4970 (N_4970,N_1087,N_887);
and U4971 (N_4971,N_970,N_721);
nor U4972 (N_4972,N_769,N_2027);
nand U4973 (N_4973,N_2397,N_2085);
nand U4974 (N_4974,N_777,N_208);
nor U4975 (N_4975,N_1977,N_946);
nand U4976 (N_4976,N_2220,N_1314);
and U4977 (N_4977,N_752,N_980);
or U4978 (N_4978,N_2152,N_1665);
nand U4979 (N_4979,N_2411,N_1789);
nor U4980 (N_4980,N_1063,N_2065);
or U4981 (N_4981,N_1443,N_1627);
nor U4982 (N_4982,N_1370,N_962);
and U4983 (N_4983,N_341,N_2084);
nor U4984 (N_4984,N_56,N_1143);
nor U4985 (N_4985,N_1396,N_1117);
or U4986 (N_4986,N_220,N_825);
or U4987 (N_4987,N_1972,N_2131);
and U4988 (N_4988,N_180,N_511);
or U4989 (N_4989,N_472,N_616);
nor U4990 (N_4990,N_393,N_1035);
or U4991 (N_4991,N_611,N_1679);
nand U4992 (N_4992,N_2489,N_598);
nand U4993 (N_4993,N_1159,N_1587);
nor U4994 (N_4994,N_1171,N_1200);
nor U4995 (N_4995,N_1689,N_513);
or U4996 (N_4996,N_136,N_1499);
and U4997 (N_4997,N_151,N_2110);
nand U4998 (N_4998,N_9,N_381);
xnor U4999 (N_4999,N_1703,N_97);
or U5000 (N_5000,N_2800,N_3791);
and U5001 (N_5001,N_3758,N_2998);
nand U5002 (N_5002,N_3393,N_4102);
nand U5003 (N_5003,N_4621,N_4875);
and U5004 (N_5004,N_3987,N_3961);
and U5005 (N_5005,N_3755,N_3965);
or U5006 (N_5006,N_3578,N_4497);
nor U5007 (N_5007,N_4629,N_4751);
or U5008 (N_5008,N_4563,N_4492);
and U5009 (N_5009,N_4516,N_3364);
nand U5010 (N_5010,N_3597,N_4351);
nor U5011 (N_5011,N_4525,N_4521);
nor U5012 (N_5012,N_4661,N_4366);
or U5013 (N_5013,N_3512,N_3410);
or U5014 (N_5014,N_3291,N_3833);
nor U5015 (N_5015,N_3341,N_4717);
nand U5016 (N_5016,N_4644,N_4152);
or U5017 (N_5017,N_4568,N_3325);
nand U5018 (N_5018,N_4474,N_4550);
and U5019 (N_5019,N_4197,N_4898);
xor U5020 (N_5020,N_4647,N_4071);
nor U5021 (N_5021,N_3979,N_2944);
or U5022 (N_5022,N_3228,N_3124);
nand U5023 (N_5023,N_4515,N_4211);
and U5024 (N_5024,N_4358,N_2730);
and U5025 (N_5025,N_4893,N_4559);
xnor U5026 (N_5026,N_4467,N_2544);
or U5027 (N_5027,N_3395,N_4592);
and U5028 (N_5028,N_3792,N_3397);
nor U5029 (N_5029,N_3862,N_2665);
nand U5030 (N_5030,N_4763,N_2719);
nand U5031 (N_5031,N_3194,N_3760);
or U5032 (N_5032,N_4498,N_3317);
nor U5033 (N_5033,N_4458,N_4291);
or U5034 (N_5034,N_4546,N_3158);
and U5035 (N_5035,N_2969,N_3136);
and U5036 (N_5036,N_2811,N_2554);
and U5037 (N_5037,N_4585,N_4596);
nor U5038 (N_5038,N_2648,N_2988);
and U5039 (N_5039,N_4586,N_2832);
and U5040 (N_5040,N_4134,N_4948);
and U5041 (N_5041,N_3593,N_4496);
nor U5042 (N_5042,N_4506,N_4942);
nand U5043 (N_5043,N_3037,N_4398);
nand U5044 (N_5044,N_4907,N_3362);
nand U5045 (N_5045,N_3730,N_2706);
nand U5046 (N_5046,N_3352,N_4173);
nor U5047 (N_5047,N_2760,N_2804);
and U5048 (N_5048,N_4535,N_4547);
nand U5049 (N_5049,N_4713,N_4182);
nor U5050 (N_5050,N_4040,N_4016);
nand U5051 (N_5051,N_4029,N_3371);
nand U5052 (N_5052,N_4681,N_3957);
nor U5053 (N_5053,N_3480,N_4840);
or U5054 (N_5054,N_3763,N_3648);
or U5055 (N_5055,N_4817,N_4979);
or U5056 (N_5056,N_4962,N_3592);
or U5057 (N_5057,N_4815,N_4143);
and U5058 (N_5058,N_3129,N_4400);
or U5059 (N_5059,N_4368,N_4131);
nor U5060 (N_5060,N_2866,N_3335);
nor U5061 (N_5061,N_4880,N_3923);
nand U5062 (N_5062,N_4154,N_2593);
xnor U5063 (N_5063,N_2623,N_3048);
nand U5064 (N_5064,N_2978,N_4419);
nor U5065 (N_5065,N_4047,N_4045);
nor U5066 (N_5066,N_4825,N_3983);
nor U5067 (N_5067,N_3798,N_4561);
xnor U5068 (N_5068,N_4830,N_2683);
nor U5069 (N_5069,N_4837,N_4660);
and U5070 (N_5070,N_3533,N_4532);
nor U5071 (N_5071,N_2555,N_4334);
nand U5072 (N_5072,N_3296,N_3333);
and U5073 (N_5073,N_2870,N_3265);
or U5074 (N_5074,N_2673,N_4350);
or U5075 (N_5075,N_4427,N_2518);
nand U5076 (N_5076,N_3693,N_4557);
and U5077 (N_5077,N_3458,N_4487);
and U5078 (N_5078,N_3354,N_3982);
xnor U5079 (N_5079,N_3985,N_4059);
nand U5080 (N_5080,N_3163,N_3249);
nor U5081 (N_5081,N_2604,N_3051);
and U5082 (N_5082,N_3407,N_3677);
and U5083 (N_5083,N_2505,N_4000);
and U5084 (N_5084,N_4638,N_3479);
or U5085 (N_5085,N_3485,N_3161);
xor U5086 (N_5086,N_3142,N_2887);
and U5087 (N_5087,N_3771,N_2512);
or U5088 (N_5088,N_4193,N_3254);
nand U5089 (N_5089,N_3858,N_3277);
or U5090 (N_5090,N_3890,N_3524);
nand U5091 (N_5091,N_4931,N_2976);
nand U5092 (N_5092,N_3525,N_4798);
and U5093 (N_5093,N_3422,N_4331);
or U5094 (N_5094,N_4337,N_3306);
and U5095 (N_5095,N_3856,N_3756);
or U5096 (N_5096,N_3276,N_2680);
and U5097 (N_5097,N_4773,N_4578);
and U5098 (N_5098,N_4604,N_3537);
nand U5099 (N_5099,N_3218,N_3319);
and U5100 (N_5100,N_4064,N_3505);
and U5101 (N_5101,N_2594,N_3391);
nand U5102 (N_5102,N_4272,N_4949);
and U5103 (N_5103,N_3871,N_3713);
nand U5104 (N_5104,N_4453,N_2956);
nor U5105 (N_5105,N_4223,N_3717);
nand U5106 (N_5106,N_3247,N_4758);
or U5107 (N_5107,N_4821,N_2628);
or U5108 (N_5108,N_2696,N_3409);
nand U5109 (N_5109,N_4121,N_4411);
and U5110 (N_5110,N_3206,N_2773);
or U5111 (N_5111,N_3672,N_3554);
nand U5112 (N_5112,N_4999,N_4285);
and U5113 (N_5113,N_4150,N_4384);
xor U5114 (N_5114,N_4764,N_3788);
or U5115 (N_5115,N_3171,N_2578);
and U5116 (N_5116,N_2500,N_3849);
nand U5117 (N_5117,N_4021,N_2691);
and U5118 (N_5118,N_3112,N_3236);
nand U5119 (N_5119,N_3618,N_3326);
or U5120 (N_5120,N_2847,N_4381);
or U5121 (N_5121,N_2888,N_3538);
nor U5122 (N_5122,N_4194,N_4116);
and U5123 (N_5123,N_3470,N_2961);
nand U5124 (N_5124,N_2589,N_4097);
nor U5125 (N_5125,N_2983,N_3483);
and U5126 (N_5126,N_2861,N_3387);
nand U5127 (N_5127,N_4756,N_4290);
or U5128 (N_5128,N_4281,N_4611);
nor U5129 (N_5129,N_3603,N_3684);
nand U5130 (N_5130,N_3655,N_2975);
and U5131 (N_5131,N_3845,N_4663);
or U5132 (N_5132,N_2645,N_4551);
or U5133 (N_5133,N_3912,N_3619);
or U5134 (N_5134,N_4365,N_3383);
and U5135 (N_5135,N_4712,N_3570);
xnor U5136 (N_5136,N_4231,N_3068);
and U5137 (N_5137,N_3318,N_3567);
or U5138 (N_5138,N_4299,N_2559);
nand U5139 (N_5139,N_4235,N_3239);
nor U5140 (N_5140,N_3049,N_3436);
and U5141 (N_5141,N_4389,N_4273);
nand U5142 (N_5142,N_3356,N_4617);
or U5143 (N_5143,N_4656,N_4424);
and U5144 (N_5144,N_3621,N_3038);
and U5145 (N_5145,N_2721,N_2729);
and U5146 (N_5146,N_4108,N_3565);
nand U5147 (N_5147,N_4011,N_4459);
and U5148 (N_5148,N_4239,N_3959);
or U5149 (N_5149,N_2560,N_2957);
nor U5150 (N_5150,N_2783,N_4715);
nor U5151 (N_5151,N_2584,N_2611);
and U5152 (N_5152,N_4205,N_4128);
or U5153 (N_5153,N_4106,N_4510);
nor U5154 (N_5154,N_3951,N_2855);
xnor U5155 (N_5155,N_3696,N_4049);
nand U5156 (N_5156,N_4704,N_3465);
and U5157 (N_5157,N_3885,N_4399);
nor U5158 (N_5158,N_3581,N_3240);
or U5159 (N_5159,N_3650,N_4544);
nor U5160 (N_5160,N_2826,N_4031);
xnor U5161 (N_5161,N_4484,N_4328);
nand U5162 (N_5162,N_3147,N_3992);
or U5163 (N_5163,N_3935,N_4144);
nor U5164 (N_5164,N_3761,N_3767);
nor U5165 (N_5165,N_2769,N_4086);
nor U5166 (N_5166,N_4813,N_4500);
nand U5167 (N_5167,N_2600,N_4556);
nand U5168 (N_5168,N_2885,N_4125);
or U5169 (N_5169,N_2960,N_3309);
nand U5170 (N_5170,N_2917,N_4085);
nand U5171 (N_5171,N_4930,N_2839);
nor U5172 (N_5172,N_3423,N_4548);
nand U5173 (N_5173,N_4985,N_4870);
and U5174 (N_5174,N_2844,N_4669);
nand U5175 (N_5175,N_2601,N_3904);
nand U5176 (N_5176,N_4362,N_3210);
nand U5177 (N_5177,N_3338,N_4853);
or U5178 (N_5178,N_3886,N_3521);
nor U5179 (N_5179,N_4781,N_4402);
nand U5180 (N_5180,N_4140,N_3063);
and U5181 (N_5181,N_2525,N_3810);
and U5182 (N_5182,N_3934,N_3852);
nor U5183 (N_5183,N_4294,N_2881);
and U5184 (N_5184,N_3750,N_3739);
nor U5185 (N_5185,N_4412,N_3579);
nor U5186 (N_5186,N_4593,N_3360);
nand U5187 (N_5187,N_4444,N_4543);
nand U5188 (N_5188,N_4785,N_3057);
or U5189 (N_5189,N_4303,N_3462);
nor U5190 (N_5190,N_4302,N_4729);
nor U5191 (N_5191,N_4320,N_4927);
nand U5192 (N_5192,N_4565,N_2949);
nor U5193 (N_5193,N_4918,N_3117);
and U5194 (N_5194,N_3549,N_4808);
or U5195 (N_5195,N_4483,N_4261);
and U5196 (N_5196,N_4939,N_4020);
nor U5197 (N_5197,N_4854,N_4843);
nand U5198 (N_5198,N_3144,N_4124);
or U5199 (N_5199,N_4195,N_4008);
nand U5200 (N_5200,N_3146,N_4324);
and U5201 (N_5201,N_4944,N_4508);
or U5202 (N_5202,N_3825,N_3346);
or U5203 (N_5203,N_4142,N_3006);
nand U5204 (N_5204,N_4452,N_4456);
and U5205 (N_5205,N_3310,N_2892);
or U5206 (N_5206,N_2583,N_3154);
nor U5207 (N_5207,N_3607,N_4101);
or U5208 (N_5208,N_3072,N_3999);
nor U5209 (N_5209,N_2527,N_4397);
nand U5210 (N_5210,N_3417,N_4673);
and U5211 (N_5211,N_2767,N_3751);
xnor U5212 (N_5212,N_2869,N_4860);
and U5213 (N_5213,N_4014,N_4185);
nor U5214 (N_5214,N_4626,N_4706);
and U5215 (N_5215,N_4753,N_3198);
and U5216 (N_5216,N_3754,N_2842);
nand U5217 (N_5217,N_3520,N_3111);
or U5218 (N_5218,N_4623,N_3910);
and U5219 (N_5219,N_2548,N_4845);
or U5220 (N_5220,N_4080,N_3237);
nand U5221 (N_5221,N_3938,N_3324);
nor U5222 (N_5222,N_3009,N_3686);
nand U5223 (N_5223,N_2854,N_3671);
nand U5224 (N_5224,N_2935,N_3615);
nand U5225 (N_5225,N_2533,N_2794);
nor U5226 (N_5226,N_4494,N_4030);
or U5227 (N_5227,N_3109,N_4972);
nand U5228 (N_5228,N_3605,N_4316);
nand U5229 (N_5229,N_3811,N_4718);
or U5230 (N_5230,N_4913,N_3971);
and U5231 (N_5231,N_3365,N_4742);
and U5232 (N_5232,N_3019,N_3190);
or U5233 (N_5233,N_2558,N_3883);
and U5234 (N_5234,N_4890,N_3468);
and U5235 (N_5235,N_4344,N_3114);
and U5236 (N_5236,N_3864,N_3793);
nor U5237 (N_5237,N_3973,N_4759);
nor U5238 (N_5238,N_3839,N_4341);
xor U5239 (N_5239,N_2521,N_4364);
nor U5240 (N_5240,N_4929,N_3424);
and U5241 (N_5241,N_3900,N_3683);
or U5242 (N_5242,N_3489,N_4639);
nand U5243 (N_5243,N_2681,N_2751);
and U5244 (N_5244,N_4372,N_2971);
or U5245 (N_5245,N_2856,N_3252);
and U5246 (N_5246,N_4079,N_3242);
nand U5247 (N_5247,N_4852,N_3921);
nand U5248 (N_5248,N_2660,N_2724);
nand U5249 (N_5249,N_2549,N_4735);
or U5250 (N_5250,N_2543,N_3818);
or U5251 (N_5251,N_4834,N_4856);
and U5252 (N_5252,N_4158,N_4478);
nor U5253 (N_5253,N_4827,N_3588);
or U5254 (N_5254,N_4187,N_3661);
nor U5255 (N_5255,N_3840,N_2891);
or U5256 (N_5256,N_4092,N_3975);
or U5257 (N_5257,N_2734,N_2625);
nand U5258 (N_5258,N_3083,N_4635);
nor U5259 (N_5259,N_2801,N_4450);
and U5260 (N_5260,N_2556,N_2713);
or U5261 (N_5261,N_3281,N_4004);
nor U5262 (N_5262,N_4876,N_3466);
or U5263 (N_5263,N_3413,N_4694);
nor U5264 (N_5264,N_2984,N_3427);
nor U5265 (N_5265,N_3953,N_4081);
nor U5266 (N_5266,N_2662,N_4333);
nor U5267 (N_5267,N_3636,N_4096);
nand U5268 (N_5268,N_4903,N_3969);
nand U5269 (N_5269,N_2757,N_3843);
and U5270 (N_5270,N_2727,N_4468);
nand U5271 (N_5271,N_3402,N_3404);
nand U5272 (N_5272,N_4265,N_4664);
and U5273 (N_5273,N_4693,N_2868);
and U5274 (N_5274,N_4413,N_3574);
nand U5275 (N_5275,N_2725,N_4159);
or U5276 (N_5276,N_4541,N_3189);
or U5277 (N_5277,N_4218,N_4019);
and U5278 (N_5278,N_2745,N_2828);
nor U5279 (N_5279,N_3966,N_3630);
nand U5280 (N_5280,N_4191,N_4373);
and U5281 (N_5281,N_3685,N_3344);
nand U5282 (N_5282,N_3080,N_4325);
nand U5283 (N_5283,N_4935,N_4613);
or U5284 (N_5284,N_3243,N_4275);
and U5285 (N_5285,N_4990,N_3530);
nor U5286 (N_5286,N_3816,N_2676);
nand U5287 (N_5287,N_3414,N_3742);
and U5288 (N_5288,N_2749,N_3244);
nand U5289 (N_5289,N_4371,N_4915);
and U5290 (N_5290,N_3687,N_4212);
or U5291 (N_5291,N_2596,N_3174);
and U5292 (N_5292,N_2802,N_3909);
or U5293 (N_5293,N_3780,N_3151);
nand U5294 (N_5294,N_4480,N_3017);
or U5295 (N_5295,N_2924,N_3855);
and U5296 (N_5296,N_4858,N_2797);
and U5297 (N_5297,N_2571,N_4038);
or U5298 (N_5298,N_3664,N_2520);
or U5299 (N_5299,N_3178,N_4714);
or U5300 (N_5300,N_4039,N_4301);
nor U5301 (N_5301,N_4957,N_3451);
and U5302 (N_5302,N_4940,N_4387);
nor U5303 (N_5303,N_3370,N_3692);
nand U5304 (N_5304,N_4680,N_3493);
nor U5305 (N_5305,N_2831,N_3203);
nand U5306 (N_5306,N_3842,N_3127);
and U5307 (N_5307,N_4968,N_4479);
nor U5308 (N_5308,N_4417,N_3998);
nor U5309 (N_5309,N_3042,N_2718);
and U5310 (N_5310,N_4287,N_3478);
or U5311 (N_5311,N_4282,N_4820);
nand U5312 (N_5312,N_3859,N_2912);
and U5313 (N_5313,N_4863,N_4309);
and U5314 (N_5314,N_2863,N_2710);
nor U5315 (N_5315,N_2882,N_4104);
nor U5316 (N_5316,N_2789,N_3180);
or U5317 (N_5317,N_3786,N_4594);
nand U5318 (N_5318,N_2954,N_4636);
nor U5319 (N_5319,N_3484,N_4702);
and U5320 (N_5320,N_4010,N_3508);
or U5321 (N_5321,N_3216,N_2570);
nor U5322 (N_5322,N_4296,N_4002);
nand U5323 (N_5323,N_4105,N_4743);
or U5324 (N_5324,N_4583,N_4449);
nand U5325 (N_5325,N_4477,N_3944);
nand U5326 (N_5326,N_4229,N_3749);
nand U5327 (N_5327,N_4530,N_3379);
and U5328 (N_5328,N_3195,N_3459);
nor U5329 (N_5329,N_3928,N_4677);
or U5330 (N_5330,N_4066,N_3990);
nand U5331 (N_5331,N_4679,N_2968);
or U5332 (N_5332,N_2874,N_4920);
and U5333 (N_5333,N_4975,N_3746);
and U5334 (N_5334,N_4848,N_3775);
and U5335 (N_5335,N_4986,N_3293);
or U5336 (N_5336,N_3170,N_3822);
or U5337 (N_5337,N_4847,N_2654);
nor U5338 (N_5338,N_4236,N_2952);
nor U5339 (N_5339,N_3528,N_4386);
nor U5340 (N_5340,N_3962,N_3507);
and U5341 (N_5341,N_2809,N_3014);
or U5342 (N_5342,N_2646,N_3942);
and U5343 (N_5343,N_3429,N_4326);
xnor U5344 (N_5344,N_2784,N_2945);
nor U5345 (N_5345,N_2851,N_3384);
and U5346 (N_5346,N_3782,N_4074);
or U5347 (N_5347,N_3801,N_4090);
and U5348 (N_5348,N_3272,N_2889);
and U5349 (N_5349,N_3817,N_4818);
nor U5350 (N_5350,N_3644,N_2698);
and U5351 (N_5351,N_2865,N_4279);
or U5352 (N_5352,N_2587,N_2682);
or U5353 (N_5353,N_3366,N_3079);
and U5354 (N_5354,N_3821,N_4099);
nor U5355 (N_5355,N_3590,N_2739);
nor U5356 (N_5356,N_3898,N_4132);
nor U5357 (N_5357,N_4761,N_4186);
and U5358 (N_5358,N_4857,N_4491);
nor U5359 (N_5359,N_3629,N_3740);
nor U5360 (N_5360,N_4741,N_4201);
or U5361 (N_5361,N_3369,N_3523);
nor U5362 (N_5362,N_3303,N_3441);
nor U5363 (N_5363,N_2788,N_3967);
nand U5364 (N_5364,N_4938,N_2852);
and U5365 (N_5365,N_2772,N_4652);
nand U5366 (N_5366,N_4200,N_3421);
nor U5367 (N_5367,N_2720,N_3916);
nand U5368 (N_5368,N_4046,N_3926);
and U5369 (N_5369,N_3262,N_4357);
nor U5370 (N_5370,N_2686,N_2685);
and U5371 (N_5371,N_4256,N_3986);
nand U5372 (N_5372,N_4244,N_4601);
or U5373 (N_5373,N_2904,N_2667);
nand U5374 (N_5374,N_2890,N_3645);
and U5375 (N_5375,N_3774,N_4595);
nor U5376 (N_5376,N_2823,N_4199);
or U5377 (N_5377,N_4075,N_2938);
or U5378 (N_5378,N_2753,N_2810);
or U5379 (N_5379,N_3678,N_3908);
or U5380 (N_5380,N_3994,N_3620);
nand U5381 (N_5381,N_4149,N_3669);
or U5382 (N_5382,N_4198,N_4001);
and U5383 (N_5383,N_4514,N_4851);
or U5384 (N_5384,N_4425,N_4057);
nand U5385 (N_5385,N_4674,N_3301);
nor U5386 (N_5386,N_4502,N_4100);
xnor U5387 (N_5387,N_4599,N_2886);
or U5388 (N_5388,N_4499,N_4094);
nor U5389 (N_5389,N_2764,N_4526);
nand U5390 (N_5390,N_3450,N_3232);
and U5391 (N_5391,N_3679,N_3492);
nand U5392 (N_5392,N_4312,N_3694);
nand U5393 (N_5393,N_3777,N_4118);
nor U5394 (N_5394,N_4887,N_4462);
nand U5395 (N_5395,N_4575,N_3226);
nor U5396 (N_5396,N_4012,N_2922);
and U5397 (N_5397,N_3718,N_2965);
nand U5398 (N_5398,N_4338,N_3841);
or U5399 (N_5399,N_2607,N_3453);
nor U5400 (N_5400,N_4165,N_2837);
xor U5401 (N_5401,N_3133,N_2655);
nor U5402 (N_5402,N_3295,N_4087);
nand U5403 (N_5403,N_3400,N_2781);
nor U5404 (N_5404,N_2825,N_3930);
or U5405 (N_5405,N_3534,N_4527);
and U5406 (N_5406,N_2782,N_4609);
or U5407 (N_5407,N_4612,N_3457);
or U5408 (N_5408,N_3700,N_4597);
xnor U5409 (N_5409,N_3209,N_3110);
xor U5410 (N_5410,N_4422,N_4598);
or U5411 (N_5411,N_2736,N_2511);
and U5412 (N_5412,N_2818,N_4367);
and U5413 (N_5413,N_3285,N_3974);
and U5414 (N_5414,N_3269,N_2668);
and U5415 (N_5415,N_4616,N_3116);
and U5416 (N_5416,N_4724,N_4649);
nor U5417 (N_5417,N_4906,N_4603);
and U5418 (N_5418,N_3380,N_4405);
nor U5419 (N_5419,N_2977,N_2641);
xnor U5420 (N_5420,N_4088,N_4571);
or U5421 (N_5421,N_3545,N_4760);
nand U5422 (N_5422,N_4572,N_4025);
or U5423 (N_5423,N_4782,N_3207);
nand U5424 (N_5424,N_3572,N_3869);
or U5425 (N_5425,N_2714,N_2858);
nand U5426 (N_5426,N_4879,N_3772);
and U5427 (N_5427,N_3455,N_2914);
nand U5428 (N_5428,N_3490,N_4917);
or U5429 (N_5429,N_2859,N_3220);
and U5430 (N_5430,N_4869,N_4528);
or U5431 (N_5431,N_4207,N_3005);
nand U5432 (N_5432,N_3280,N_4923);
nor U5433 (N_5433,N_3861,N_3197);
nor U5434 (N_5434,N_3461,N_2996);
nor U5435 (N_5435,N_4657,N_3613);
or U5436 (N_5436,N_4441,N_4787);
nor U5437 (N_5437,N_2678,N_3150);
nand U5438 (N_5438,N_3770,N_2848);
and U5439 (N_5439,N_4866,N_3571);
or U5440 (N_5440,N_3988,N_2808);
nor U5441 (N_5441,N_2750,N_3382);
nor U5442 (N_5442,N_2535,N_3225);
or U5443 (N_5443,N_2539,N_2950);
or U5444 (N_5444,N_4163,N_4545);
nand U5445 (N_5445,N_3271,N_4313);
nand U5446 (N_5446,N_4050,N_4306);
or U5447 (N_5447,N_3001,N_4469);
and U5448 (N_5448,N_3018,N_3826);
nor U5449 (N_5449,N_3405,N_3625);
and U5450 (N_5450,N_2923,N_4378);
and U5451 (N_5451,N_3323,N_4454);
nor U5452 (N_5452,N_4709,N_4552);
nor U5453 (N_5453,N_3828,N_3430);
or U5454 (N_5454,N_4114,N_3070);
and U5455 (N_5455,N_4802,N_2744);
nor U5456 (N_5456,N_2840,N_3997);
and U5457 (N_5457,N_3115,N_4878);
and U5458 (N_5458,N_3846,N_3632);
or U5459 (N_5459,N_3073,N_3690);
xnor U5460 (N_5460,N_4574,N_3932);
and U5461 (N_5461,N_3358,N_3292);
nor U5462 (N_5462,N_4383,N_4914);
nand U5463 (N_5463,N_4631,N_4699);
and U5464 (N_5464,N_4024,N_4461);
or U5465 (N_5465,N_3652,N_4439);
nand U5466 (N_5466,N_4130,N_3302);
and U5467 (N_5467,N_3355,N_2973);
and U5468 (N_5468,N_2761,N_2829);
or U5469 (N_5469,N_4241,N_2759);
nor U5470 (N_5470,N_2542,N_3497);
nand U5471 (N_5471,N_4327,N_2805);
or U5472 (N_5472,N_4928,N_4844);
nand U5473 (N_5473,N_2516,N_2806);
and U5474 (N_5474,N_3100,N_3546);
nor U5475 (N_5475,N_3963,N_2790);
or U5476 (N_5476,N_3991,N_3710);
nor U5477 (N_5477,N_3901,N_3311);
or U5478 (N_5478,N_3604,N_3182);
nor U5479 (N_5479,N_3175,N_3097);
and U5480 (N_5480,N_2843,N_3741);
nor U5481 (N_5481,N_3569,N_3223);
or U5482 (N_5482,N_4188,N_4446);
nor U5483 (N_5483,N_3606,N_4909);
nand U5484 (N_5484,N_3212,N_3865);
nand U5485 (N_5485,N_2872,N_4676);
or U5486 (N_5486,N_3555,N_4691);
and U5487 (N_5487,N_2576,N_4776);
or U5488 (N_5488,N_4481,N_3820);
nand U5489 (N_5489,N_4954,N_3045);
nor U5490 (N_5490,N_4540,N_4242);
and U5491 (N_5491,N_4747,N_2709);
and U5492 (N_5492,N_2931,N_3540);
or U5493 (N_5493,N_4642,N_3654);
or U5494 (N_5494,N_4181,N_3394);
and U5495 (N_5495,N_4767,N_3887);
and U5496 (N_5496,N_4916,N_2684);
nand U5497 (N_5497,N_4960,N_3179);
nand U5498 (N_5498,N_3010,N_2633);
and U5499 (N_5499,N_4888,N_3917);
nor U5500 (N_5500,N_3105,N_2964);
or U5501 (N_5501,N_2591,N_2878);
nor U5502 (N_5502,N_3547,N_3800);
nor U5503 (N_5503,N_4539,N_2906);
and U5504 (N_5504,N_2746,N_4896);
and U5505 (N_5505,N_3797,N_4668);
or U5506 (N_5506,N_4925,N_4396);
nor U5507 (N_5507,N_3008,N_3829);
xor U5508 (N_5508,N_3809,N_3681);
or U5509 (N_5509,N_2529,N_3487);
xnor U5510 (N_5510,N_3876,N_4356);
or U5511 (N_5511,N_3108,N_2884);
and U5512 (N_5512,N_4126,N_4055);
and U5513 (N_5513,N_2763,N_3082);
and U5514 (N_5514,N_3106,N_4471);
and U5515 (N_5515,N_2702,N_4007);
or U5516 (N_5516,N_2771,N_4434);
nand U5517 (N_5517,N_2656,N_2639);
nor U5518 (N_5518,N_3359,N_4053);
and U5519 (N_5519,N_3434,N_3711);
nand U5520 (N_5520,N_4945,N_3511);
or U5521 (N_5521,N_2943,N_4009);
nor U5522 (N_5522,N_4346,N_4068);
nor U5523 (N_5523,N_4690,N_4359);
or U5524 (N_5524,N_4251,N_3260);
or U5525 (N_5525,N_2896,N_3177);
or U5526 (N_5526,N_2928,N_2880);
or U5527 (N_5527,N_3428,N_3217);
and U5528 (N_5528,N_3738,N_4697);
and U5529 (N_5529,N_4736,N_4385);
and U5530 (N_5530,N_3851,N_3256);
nor U5531 (N_5531,N_4005,N_4093);
or U5532 (N_5532,N_3764,N_3074);
nor U5533 (N_5533,N_2613,N_3585);
nor U5534 (N_5534,N_3726,N_3078);
or U5535 (N_5535,N_3550,N_3258);
and U5536 (N_5536,N_2770,N_2834);
nand U5537 (N_5537,N_4922,N_4951);
and U5538 (N_5538,N_3647,N_3789);
or U5539 (N_5539,N_4978,N_4329);
nand U5540 (N_5540,N_2562,N_4822);
and U5541 (N_5541,N_2700,N_4070);
nor U5542 (N_5542,N_4947,N_3753);
nor U5543 (N_5543,N_4625,N_3090);
or U5544 (N_5544,N_3704,N_3808);
or U5545 (N_5545,N_3165,N_3844);
or U5546 (N_5546,N_3835,N_4192);
and U5547 (N_5547,N_3463,N_2688);
nand U5548 (N_5548,N_3783,N_3649);
nand U5549 (N_5549,N_3176,N_4682);
nand U5550 (N_5550,N_3066,N_4804);
or U5551 (N_5551,N_4641,N_4463);
nor U5552 (N_5552,N_3187,N_3385);
or U5553 (N_5553,N_4643,N_3674);
nor U5554 (N_5554,N_3035,N_3213);
and U5555 (N_5555,N_3640,N_4308);
nor U5556 (N_5556,N_4849,N_4900);
nor U5557 (N_5557,N_2614,N_3399);
and U5558 (N_5558,N_2540,N_4722);
and U5559 (N_5559,N_4790,N_3367);
or U5560 (N_5560,N_4662,N_3897);
and U5561 (N_5561,N_3744,N_3680);
and U5562 (N_5562,N_3733,N_3275);
xor U5563 (N_5563,N_3202,N_3481);
nor U5564 (N_5564,N_2597,N_3927);
nand U5565 (N_5565,N_3125,N_3250);
nor U5566 (N_5566,N_2907,N_3548);
and U5567 (N_5567,N_4569,N_2552);
nor U5568 (N_5568,N_3591,N_4513);
nand U5569 (N_5569,N_3449,N_4587);
or U5570 (N_5570,N_4666,N_4015);
or U5571 (N_5571,N_3331,N_3536);
and U5572 (N_5572,N_3201,N_3308);
nor U5573 (N_5573,N_2827,N_3092);
nor U5574 (N_5574,N_2778,N_4675);
or U5575 (N_5575,N_3631,N_4994);
xnor U5576 (N_5576,N_3627,N_2921);
nand U5577 (N_5577,N_2824,N_4745);
xnor U5578 (N_5578,N_2679,N_2567);
nor U5579 (N_5579,N_4728,N_2946);
nand U5580 (N_5580,N_3743,N_2708);
or U5581 (N_5581,N_4864,N_2999);
nor U5582 (N_5582,N_3334,N_4196);
and U5583 (N_5583,N_4671,N_4868);
nor U5584 (N_5584,N_3184,N_4651);
nor U5585 (N_5585,N_3204,N_3012);
or U5586 (N_5586,N_2572,N_3568);
nor U5587 (N_5587,N_4352,N_4801);
nor U5588 (N_5588,N_3535,N_4321);
or U5589 (N_5589,N_2553,N_4110);
or U5590 (N_5590,N_4992,N_4460);
nor U5591 (N_5591,N_3119,N_3586);
or U5592 (N_5592,N_2786,N_3386);
nor U5593 (N_5593,N_4103,N_3670);
nand U5594 (N_5594,N_3279,N_4964);
and U5595 (N_5595,N_2913,N_4067);
nor U5596 (N_5596,N_3781,N_2942);
nand U5597 (N_5597,N_2503,N_4162);
or U5598 (N_5598,N_4716,N_4209);
nor U5599 (N_5599,N_4245,N_3662);
nor U5600 (N_5600,N_4214,N_4659);
nor U5601 (N_5601,N_3940,N_3960);
nor U5602 (N_5602,N_2616,N_4379);
nand U5603 (N_5603,N_2820,N_3444);
and U5604 (N_5604,N_4330,N_2803);
nand U5605 (N_5605,N_3388,N_3130);
or U5606 (N_5606,N_3193,N_4051);
or U5607 (N_5607,N_2979,N_3141);
or U5608 (N_5608,N_2541,N_2672);
xor U5609 (N_5609,N_3259,N_4475);
and U5610 (N_5610,N_4769,N_4311);
xnor U5611 (N_5611,N_3349,N_4044);
and U5612 (N_5612,N_4348,N_2707);
nor U5613 (N_5613,N_2528,N_3719);
nor U5614 (N_5614,N_4926,N_4423);
nor U5615 (N_5615,N_2510,N_3476);
nor U5616 (N_5616,N_4377,N_4447);
nand U5617 (N_5617,N_4180,N_2732);
or U5618 (N_5618,N_3267,N_2893);
nand U5619 (N_5619,N_2635,N_3562);
xor U5620 (N_5620,N_2776,N_3278);
or U5621 (N_5621,N_4109,N_4482);
or U5622 (N_5622,N_4872,N_2617);
and U5623 (N_5623,N_3494,N_4084);
or U5624 (N_5624,N_2550,N_2514);
nor U5625 (N_5625,N_4157,N_3509);
nor U5626 (N_5626,N_3257,N_4120);
and U5627 (N_5627,N_3768,N_2612);
nand U5628 (N_5628,N_4304,N_4037);
nor U5629 (N_5629,N_2780,N_2524);
or U5630 (N_5630,N_3342,N_3946);
and U5631 (N_5631,N_3542,N_2862);
or U5632 (N_5632,N_3827,N_4054);
and U5633 (N_5633,N_4995,N_2622);
or U5634 (N_5634,N_2974,N_2926);
nor U5635 (N_5635,N_2930,N_2910);
and U5636 (N_5636,N_4314,N_4805);
nand U5637 (N_5637,N_3558,N_4730);
nand U5638 (N_5638,N_3731,N_2671);
and U5639 (N_5639,N_3437,N_4278);
nor U5640 (N_5640,N_3941,N_2666);
nor U5641 (N_5641,N_4354,N_2937);
nor U5642 (N_5642,N_4969,N_3426);
and U5643 (N_5643,N_2689,N_3582);
and U5644 (N_5644,N_3381,N_4654);
nor U5645 (N_5645,N_3721,N_3378);
nand U5646 (N_5646,N_4943,N_4560);
nand U5647 (N_5647,N_4215,N_4048);
nand U5648 (N_5648,N_3205,N_3657);
nand U5649 (N_5649,N_4762,N_4789);
and U5650 (N_5650,N_3769,N_3499);
nand U5651 (N_5651,N_3188,N_3911);
nor U5652 (N_5652,N_4179,N_3735);
or U5653 (N_5653,N_2664,N_2608);
nor U5654 (N_5654,N_4605,N_3819);
or U5655 (N_5655,N_3411,N_3868);
and U5656 (N_5656,N_4961,N_4139);
xnor U5657 (N_5657,N_4155,N_3047);
or U5658 (N_5658,N_2569,N_4028);
nand U5659 (N_5659,N_2853,N_4300);
or U5660 (N_5660,N_3069,N_2636);
nor U5661 (N_5661,N_3504,N_4393);
nand U5662 (N_5662,N_4846,N_2658);
nand U5663 (N_5663,N_4127,N_2835);
or U5664 (N_5664,N_3804,N_4141);
or U5665 (N_5665,N_3031,N_4343);
and U5666 (N_5666,N_4203,N_4564);
nand U5667 (N_5667,N_3183,N_2916);
nand U5668 (N_5668,N_4089,N_4737);
nand U5669 (N_5669,N_2743,N_4298);
and U5670 (N_5670,N_3392,N_2687);
nand U5671 (N_5671,N_4984,N_4268);
and U5672 (N_5672,N_3007,N_3149);
nor U5673 (N_5673,N_2595,N_3899);
nand U5674 (N_5674,N_2701,N_3191);
and U5675 (N_5675,N_2993,N_3779);
nand U5676 (N_5676,N_4146,N_3706);
nor U5677 (N_5677,N_4058,N_3646);
and U5678 (N_5678,N_4486,N_4271);
nor U5679 (N_5679,N_2561,N_3375);
or U5680 (N_5680,N_2796,N_3970);
or U5681 (N_5681,N_3838,N_3919);
or U5682 (N_5682,N_4435,N_3996);
or U5683 (N_5683,N_4683,N_4855);
nor U5684 (N_5684,N_4176,N_4336);
xnor U5685 (N_5685,N_2532,N_4755);
and U5686 (N_5686,N_2845,N_4672);
and U5687 (N_5687,N_2755,N_3233);
or U5688 (N_5688,N_4098,N_3506);
nand U5689 (N_5689,N_2501,N_3219);
nor U5690 (N_5690,N_2661,N_3329);
nor U5691 (N_5691,N_4842,N_2657);
nand U5692 (N_5692,N_2901,N_3737);
and U5693 (N_5693,N_4226,N_3651);
nor U5694 (N_5694,N_4430,N_3440);
nand U5695 (N_5695,N_3778,N_2502);
nor U5696 (N_5696,N_4952,N_4216);
and U5697 (N_5697,N_4780,N_4809);
nor U5698 (N_5698,N_3796,N_4065);
or U5699 (N_5699,N_3094,N_4361);
and U5700 (N_5700,N_4958,N_3526);
and U5701 (N_5701,N_3431,N_3123);
nor U5702 (N_5702,N_4225,N_4443);
nor U5703 (N_5703,N_4164,N_4493);
or U5704 (N_5704,N_3091,N_4520);
and U5705 (N_5705,N_2740,N_3230);
and U5706 (N_5706,N_2581,N_3831);
nand U5707 (N_5707,N_4522,N_3408);
or U5708 (N_5708,N_2741,N_3027);
or U5709 (N_5709,N_4248,N_2620);
or U5710 (N_5710,N_4832,N_3925);
nor U5711 (N_5711,N_4841,N_4246);
and U5712 (N_5712,N_3030,N_2677);
or U5713 (N_5713,N_3245,N_2723);
or U5714 (N_5714,N_3289,N_3266);
xnor U5715 (N_5715,N_4284,N_4901);
or U5716 (N_5716,N_3668,N_2627);
nand U5717 (N_5717,N_4013,N_3140);
nor U5718 (N_5718,N_4726,N_4784);
or U5719 (N_5719,N_4701,N_3255);
or U5720 (N_5720,N_3251,N_2526);
or U5721 (N_5721,N_3439,N_3939);
nor U5722 (N_5722,N_2911,N_3446);
nor U5723 (N_5723,N_3734,N_4775);
nand U5724 (N_5724,N_3878,N_2592);
and U5725 (N_5725,N_4018,N_4777);
nand U5726 (N_5726,N_4826,N_3516);
and U5727 (N_5727,N_3473,N_4171);
nor U5728 (N_5728,N_4517,N_4369);
nor U5729 (N_5729,N_3660,N_2900);
and U5730 (N_5730,N_3874,N_2506);
nor U5731 (N_5731,N_4703,N_4573);
and U5732 (N_5732,N_4395,N_2624);
nor U5733 (N_5733,N_4210,N_3101);
and U5734 (N_5734,N_2777,N_4262);
nand U5735 (N_5735,N_3241,N_4689);
nor U5736 (N_5736,N_2940,N_3145);
and U5737 (N_5737,N_4732,N_3950);
or U5738 (N_5738,N_2659,N_3948);
nand U5739 (N_5739,N_3784,N_3502);
or U5740 (N_5740,N_3015,N_3004);
nand U5741 (N_5741,N_3121,N_3025);
nor U5742 (N_5742,N_4891,N_3920);
nand U5743 (N_5743,N_4495,N_4519);
or U5744 (N_5744,N_3616,N_4250);
or U5745 (N_5745,N_4558,N_4062);
or U5746 (N_5746,N_4529,N_3491);
xnor U5747 (N_5747,N_2929,N_4796);
nand U5748 (N_5748,N_3284,N_3043);
nor U5749 (N_5749,N_3795,N_4027);
nand U5750 (N_5750,N_4511,N_3166);
or U5751 (N_5751,N_4950,N_3725);
nand U5752 (N_5752,N_3438,N_4700);
nor U5753 (N_5753,N_3299,N_4317);
and U5754 (N_5754,N_4274,N_2897);
or U5755 (N_5755,N_2813,N_3673);
nand U5756 (N_5756,N_2565,N_4615);
and U5757 (N_5757,N_2798,N_2985);
nand U5758 (N_5758,N_4628,N_3098);
and U5759 (N_5759,N_3729,N_3747);
and U5760 (N_5760,N_3936,N_4485);
nand U5761 (N_5761,N_3854,N_4734);
or U5762 (N_5762,N_4111,N_2598);
and U5763 (N_5763,N_3877,N_2517);
nand U5764 (N_5764,N_2568,N_3698);
or U5765 (N_5765,N_3088,N_3238);
or U5766 (N_5766,N_2747,N_4895);
nand U5767 (N_5767,N_4280,N_2812);
nor U5768 (N_5768,N_4882,N_4345);
and U5769 (N_5769,N_3062,N_2711);
xnor U5770 (N_5770,N_3863,N_2925);
and U5771 (N_5771,N_4752,N_3656);
nand U5772 (N_5772,N_4632,N_4562);
or U5773 (N_5773,N_2564,N_3328);
nand U5774 (N_5774,N_3227,N_3891);
or U5775 (N_5775,N_3137,N_2908);
and U5776 (N_5776,N_4230,N_4723);
and U5777 (N_5777,N_3442,N_4190);
nor U5778 (N_5778,N_2909,N_4305);
nand U5779 (N_5779,N_3896,N_4977);
and U5780 (N_5780,N_4222,N_2915);
or U5781 (N_5781,N_3639,N_4812);
and U5782 (N_5782,N_3714,N_2758);
and U5783 (N_5783,N_4791,N_4036);
and U5784 (N_5784,N_4172,N_2523);
and U5785 (N_5785,N_3608,N_4117);
nor U5786 (N_5786,N_4426,N_4374);
nor U5787 (N_5787,N_3155,N_3002);
or U5788 (N_5788,N_4220,N_3952);
or U5789 (N_5789,N_3748,N_3153);
nand U5790 (N_5790,N_2838,N_4489);
nor U5791 (N_5791,N_4360,N_3872);
and U5792 (N_5792,N_2695,N_3675);
and U5793 (N_5793,N_4885,N_3515);
and U5794 (N_5794,N_4505,N_3288);
nand U5795 (N_5795,N_4082,N_3185);
nand U5796 (N_5796,N_3853,N_3039);
or U5797 (N_5797,N_4342,N_2631);
nand U5798 (N_5798,N_4420,N_3699);
nand U5799 (N_5799,N_4156,N_4684);
nor U5800 (N_5800,N_4289,N_4332);
nand U5801 (N_5801,N_3085,N_4708);
nor U5802 (N_5802,N_4136,N_4221);
xor U5803 (N_5803,N_3498,N_2643);
and U5804 (N_5804,N_3968,N_3134);
and U5805 (N_5805,N_4227,N_4455);
and U5806 (N_5806,N_2955,N_3587);
or U5807 (N_5807,N_3790,N_3720);
nor U5808 (N_5808,N_3443,N_3561);
nand U5809 (N_5809,N_4589,N_4137);
nor U5810 (N_5810,N_3337,N_3553);
or U5811 (N_5811,N_2860,N_4286);
or U5812 (N_5812,N_3246,N_3638);
nor U5813 (N_5813,N_2793,N_2642);
or U5814 (N_5814,N_3022,N_3024);
nand U5815 (N_5815,N_4160,N_3026);
and U5816 (N_5816,N_4233,N_4476);
and U5817 (N_5817,N_2531,N_3635);
nand U5818 (N_5818,N_4448,N_4107);
nand U5819 (N_5819,N_2605,N_3403);
or U5820 (N_5820,N_4608,N_3041);
nor U5821 (N_5821,N_3889,N_3880);
and U5822 (N_5822,N_2959,N_3398);
or U5823 (N_5823,N_3736,N_3208);
nor U5824 (N_5824,N_4056,N_3304);
nor U5825 (N_5825,N_4069,N_2647);
nor U5826 (N_5826,N_2807,N_3067);
nand U5827 (N_5827,N_4970,N_3330);
and U5828 (N_5828,N_2610,N_3947);
and U5829 (N_5829,N_3374,N_2815);
and U5830 (N_5830,N_4989,N_4740);
or U5831 (N_5831,N_4240,N_4765);
nand U5832 (N_5832,N_4536,N_4133);
and U5833 (N_5833,N_4584,N_4871);
nand U5834 (N_5834,N_4307,N_3860);
nand U5835 (N_5835,N_3059,N_2919);
nor U5836 (N_5836,N_3617,N_2903);
and U5837 (N_5837,N_4980,N_2590);
nor U5838 (N_5838,N_3224,N_4243);
xnor U5839 (N_5839,N_4686,N_4794);
or U5840 (N_5840,N_3682,N_3766);
nor U5841 (N_5841,N_3892,N_2534);
nand U5842 (N_5842,N_4258,N_3802);
nor U5843 (N_5843,N_4655,N_4738);
nand U5844 (N_5844,N_4566,N_4270);
nor U5845 (N_5845,N_3894,N_3785);
nand U5846 (N_5846,N_4376,N_3624);
nor U5847 (N_5847,N_3514,N_4228);
xnor U5848 (N_5848,N_2958,N_4733);
and U5849 (N_5849,N_2836,N_4473);
or U5850 (N_5850,N_2995,N_4658);
nand U5851 (N_5851,N_3529,N_4627);
nand U5852 (N_5852,N_3075,N_2972);
nand U5853 (N_5853,N_4749,N_3727);
or U5854 (N_5854,N_4810,N_4355);
nor U5855 (N_5855,N_4750,N_3321);
nand U5856 (N_5856,N_4772,N_2987);
nand U5857 (N_5857,N_4823,N_3044);
and U5858 (N_5858,N_3902,N_4646);
nor U5859 (N_5859,N_3913,N_2537);
nor U5860 (N_5860,N_4178,N_2649);
or U5861 (N_5861,N_3274,N_2867);
nand U5862 (N_5862,N_4873,N_3050);
or U5863 (N_5863,N_2742,N_3666);
nor U5864 (N_5864,N_4607,N_4023);
or U5865 (N_5865,N_3401,N_4488);
nand U5866 (N_5866,N_4814,N_2947);
and U5867 (N_5867,N_4183,N_4911);
and U5868 (N_5868,N_3046,N_4670);
nand U5869 (N_5869,N_2877,N_2690);
or U5870 (N_5870,N_4624,N_2966);
and U5871 (N_5871,N_3552,N_3297);
nor U5872 (N_5872,N_3200,N_4816);
xnor U5873 (N_5873,N_4523,N_4757);
nand U5874 (N_5874,N_4555,N_2515);
or U5875 (N_5875,N_2509,N_2967);
nor U5876 (N_5876,N_4620,N_2822);
and U5877 (N_5877,N_2816,N_2920);
nor U5878 (N_5878,N_3474,N_3028);
nand U5879 (N_5879,N_4257,N_3695);
or U5880 (N_5880,N_4838,N_2650);
and U5881 (N_5881,N_3709,N_4247);
nor U5882 (N_5882,N_2791,N_3931);
nor U5883 (N_5883,N_2970,N_3488);
nor U5884 (N_5884,N_4464,N_2754);
or U5885 (N_5885,N_4189,N_3600);
or U5886 (N_5886,N_4988,N_3875);
or U5887 (N_5887,N_4292,N_3541);
and U5888 (N_5888,N_3396,N_4166);
nor U5889 (N_5889,N_3622,N_4974);
nand U5890 (N_5890,N_4912,N_3634);
and U5891 (N_5891,N_2992,N_2615);
nand U5892 (N_5892,N_3300,N_2821);
nor U5893 (N_5893,N_4518,N_3313);
and U5894 (N_5894,N_3799,N_2864);
and U5895 (N_5895,N_3532,N_4249);
nand U5896 (N_5896,N_3984,N_4237);
nand U5897 (N_5897,N_3327,N_3943);
nor U5898 (N_5898,N_4382,N_3120);
nor U5899 (N_5899,N_4034,N_4707);
xnor U5900 (N_5900,N_3995,N_4799);
and U5901 (N_5901,N_4432,N_3467);
nor U5902 (N_5902,N_4754,N_4797);
nand U5903 (N_5903,N_3283,N_2775);
nor U5904 (N_5904,N_3447,N_2588);
or U5905 (N_5905,N_3013,N_4688);
and U5906 (N_5906,N_4335,N_4622);
and U5907 (N_5907,N_3583,N_3034);
and U5908 (N_5908,N_4946,N_4537);
or U5909 (N_5909,N_3715,N_3376);
nor U5910 (N_5910,N_3976,N_3544);
nor U5911 (N_5911,N_2586,N_4401);
nor U5912 (N_5912,N_4836,N_3023);
and U5913 (N_5913,N_3823,N_3350);
nor U5914 (N_5914,N_2953,N_4534);
nor U5915 (N_5915,N_2898,N_4695);
nand U5916 (N_5916,N_4259,N_4129);
nor U5917 (N_5917,N_3732,N_3168);
nor U5918 (N_5918,N_4428,N_2989);
and U5919 (N_5919,N_3814,N_4727);
nor U5920 (N_5920,N_3584,N_4168);
nor U5921 (N_5921,N_3589,N_2603);
or U5922 (N_5922,N_3305,N_2640);
nor U5923 (N_5923,N_4353,N_3152);
or U5924 (N_5924,N_2948,N_3406);
and U5925 (N_5925,N_3559,N_3128);
and U5926 (N_5926,N_4746,N_2573);
or U5927 (N_5927,N_4470,N_3234);
nand U5928 (N_5928,N_2712,N_4554);
nor U5929 (N_5929,N_2653,N_3162);
or U5930 (N_5930,N_4322,N_4807);
nand U5931 (N_5931,N_3156,N_4908);
nand U5932 (N_5932,N_2557,N_4409);
nand U5933 (N_5933,N_2731,N_3566);
and U5934 (N_5934,N_3903,N_4148);
and U5935 (N_5935,N_4819,N_4881);
nand U5936 (N_5936,N_4266,N_4083);
or U5937 (N_5937,N_2694,N_4963);
or U5938 (N_5938,N_2507,N_2819);
or U5939 (N_5939,N_4263,N_2675);
nor U5940 (N_5940,N_3316,N_4698);
nand U5941 (N_5941,N_3503,N_3496);
nor U5942 (N_5942,N_3522,N_4725);
nand U5943 (N_5943,N_2674,N_4370);
nand U5944 (N_5944,N_3752,N_2833);
nand U5945 (N_5945,N_3611,N_3728);
or U5946 (N_5946,N_3312,N_4829);
and U5947 (N_5947,N_4403,N_3173);
and U5948 (N_5948,N_3556,N_3412);
or U5949 (N_5949,N_3486,N_4161);
or U5950 (N_5950,N_2669,N_4921);
and U5951 (N_5951,N_4602,N_3832);
nor U5952 (N_5952,N_4645,N_2895);
or U5953 (N_5953,N_4692,N_2774);
nand U5954 (N_5954,N_3065,N_3879);
nand U5955 (N_5955,N_3095,N_4897);
or U5956 (N_5956,N_4924,N_4288);
and U5957 (N_5957,N_4319,N_3290);
and U5958 (N_5958,N_2626,N_2905);
or U5959 (N_5959,N_2817,N_3701);
or U5960 (N_5960,N_3003,N_2652);
nor U5961 (N_5961,N_3222,N_3924);
nor U5962 (N_5962,N_4380,N_4490);
and U5963 (N_5963,N_3339,N_4283);
nand U5964 (N_5964,N_3495,N_2530);
or U5965 (N_5965,N_3363,N_3456);
xnor U5966 (N_5966,N_3543,N_3445);
and U5967 (N_5967,N_4472,N_3836);
nor U5968 (N_5968,N_2538,N_3659);
or U5969 (N_5969,N_4138,N_3580);
or U5970 (N_5970,N_3712,N_2609);
or U5971 (N_5971,N_4835,N_4202);
or U5972 (N_5972,N_3425,N_2566);
and U5973 (N_5973,N_3089,N_2697);
nor U5974 (N_5974,N_3131,N_3773);
or U5975 (N_5975,N_3667,N_3118);
or U5976 (N_5976,N_3061,N_2765);
nand U5977 (N_5977,N_3527,N_3164);
nand U5978 (N_5978,N_4042,N_3054);
or U5979 (N_5979,N_3286,N_4600);
or U5980 (N_5980,N_3419,N_4580);
or U5981 (N_5981,N_4766,N_4934);
nor U5982 (N_5982,N_3881,N_4619);
and U5983 (N_5983,N_2982,N_3977);
and U5984 (N_5984,N_2752,N_4862);
and U5985 (N_5985,N_2768,N_4976);
nor U5986 (N_5986,N_4169,N_2962);
nor U5987 (N_5987,N_3058,N_3933);
nand U5988 (N_5988,N_3641,N_4981);
nor U5989 (N_5989,N_4060,N_4955);
nand U5990 (N_5990,N_2692,N_4184);
nor U5991 (N_5991,N_4650,N_3813);
and U5992 (N_5992,N_3702,N_2875);
nand U5993 (N_5993,N_2795,N_2599);
xor U5994 (N_5994,N_3368,N_4033);
or U5995 (N_5995,N_2737,N_4771);
and U5996 (N_5996,N_4828,N_3757);
nor U5997 (N_5997,N_3390,N_3418);
or U5998 (N_5998,N_4696,N_3192);
and U5999 (N_5999,N_4503,N_4252);
or U6000 (N_6000,N_3626,N_3596);
and U6001 (N_6001,N_4052,N_4590);
and U6002 (N_6002,N_2990,N_4318);
and U6003 (N_6003,N_3598,N_3181);
and U6004 (N_6004,N_4531,N_3806);
and U6005 (N_6005,N_3676,N_3169);
nor U6006 (N_6006,N_3135,N_3978);
nand U6007 (N_6007,N_4151,N_2619);
nor U6008 (N_6008,N_3955,N_4063);
or U6009 (N_6009,N_3787,N_3221);
nand U6010 (N_6010,N_2849,N_3268);
or U6011 (N_6011,N_4721,N_3139);
and U6012 (N_6012,N_3776,N_3307);
nor U6013 (N_6013,N_3989,N_2846);
or U6014 (N_6014,N_3107,N_3893);
and U6015 (N_6015,N_3373,N_3980);
or U6016 (N_6016,N_4966,N_3084);
and U6017 (N_6017,N_4022,N_2726);
nor U6018 (N_6018,N_4267,N_4219);
nor U6019 (N_6019,N_3501,N_2879);
xor U6020 (N_6020,N_2602,N_4606);
and U6021 (N_6021,N_3104,N_4570);
nand U6022 (N_6022,N_3914,N_4937);
and U6023 (N_6023,N_3857,N_4685);
nor U6024 (N_6024,N_4884,N_3707);
nor U6025 (N_6025,N_3471,N_4445);
or U6026 (N_6026,N_3614,N_4414);
nor U6027 (N_6027,N_4122,N_3560);
nor U6028 (N_6028,N_3475,N_2756);
or U6029 (N_6029,N_4406,N_4418);
nor U6030 (N_6030,N_2981,N_3815);
xnor U6031 (N_6031,N_4577,N_3138);
nand U6032 (N_6032,N_2779,N_4440);
nor U6033 (N_6033,N_4983,N_3126);
nor U6034 (N_6034,N_4206,N_4687);
or U6035 (N_6035,N_3345,N_2704);
and U6036 (N_6036,N_2894,N_3895);
or U6037 (N_6037,N_4438,N_4582);
nor U6038 (N_6038,N_4408,N_4113);
nand U6039 (N_6039,N_4744,N_3332);
nor U6040 (N_6040,N_3688,N_2504);
xor U6041 (N_6041,N_3261,N_3361);
or U6042 (N_6042,N_3609,N_4095);
nand U6043 (N_6043,N_3513,N_4833);
nor U6044 (N_6044,N_3575,N_4507);
and U6045 (N_6045,N_3517,N_3011);
nand U6046 (N_6046,N_3599,N_4175);
nand U6047 (N_6047,N_2733,N_2934);
nor U6048 (N_6048,N_4610,N_3945);
nor U6049 (N_6049,N_3745,N_3000);
and U6050 (N_6050,N_2762,N_3132);
or U6051 (N_6051,N_3628,N_4026);
or U6052 (N_6052,N_2933,N_4997);
xor U6053 (N_6053,N_4770,N_4429);
nand U6054 (N_6054,N_3196,N_3954);
nor U6055 (N_6055,N_3348,N_3812);
or U6056 (N_6056,N_4431,N_4293);
and U6057 (N_6057,N_4634,N_2630);
or U6058 (N_6058,N_2871,N_4768);
and U6059 (N_6059,N_4295,N_2663);
or U6060 (N_6060,N_3958,N_3703);
or U6061 (N_6061,N_2632,N_3157);
and U6062 (N_6062,N_4576,N_4254);
nor U6063 (N_6063,N_4653,N_4982);
or U6064 (N_6064,N_4404,N_2963);
xnor U6065 (N_6065,N_3697,N_2873);
and U6066 (N_6066,N_3199,N_3643);
and U6067 (N_6067,N_3866,N_3020);
nor U6068 (N_6068,N_4859,N_2876);
nand U6069 (N_6069,N_3873,N_2585);
or U6070 (N_6070,N_3663,N_4648);
and U6071 (N_6071,N_4451,N_3322);
and U6072 (N_6072,N_3389,N_4410);
nand U6073 (N_6073,N_3964,N_4416);
nor U6074 (N_6074,N_4112,N_3081);
xor U6075 (N_6075,N_3708,N_4739);
nor U6076 (N_6076,N_2748,N_3435);
and U6077 (N_6077,N_4665,N_4224);
and U6078 (N_6078,N_3564,N_3372);
xor U6079 (N_6079,N_3637,N_2951);
or U6080 (N_6080,N_3972,N_2986);
or U6081 (N_6081,N_2547,N_3077);
or U6082 (N_6082,N_4779,N_4174);
or U6083 (N_6083,N_4933,N_4553);
nand U6084 (N_6084,N_3531,N_3122);
and U6085 (N_6085,N_3922,N_4874);
and U6086 (N_6086,N_2582,N_3103);
nor U6087 (N_6087,N_3803,N_4315);
nand U6088 (N_6088,N_4032,N_4710);
nand U6089 (N_6089,N_4217,N_4421);
and U6090 (N_6090,N_2638,N_3099);
and U6091 (N_6091,N_3377,N_3248);
nand U6092 (N_6092,N_3867,N_4208);
nor U6093 (N_6093,N_3353,N_3060);
and U6094 (N_6094,N_3029,N_4678);
nor U6095 (N_6095,N_4061,N_3231);
and U6096 (N_6096,N_2606,N_4415);
or U6097 (N_6097,N_4437,N_4407);
or U6098 (N_6098,N_3102,N_4987);
and U6099 (N_6099,N_4865,N_2850);
and U6100 (N_6100,N_4041,N_4786);
nand U6101 (N_6101,N_2980,N_2629);
and U6102 (N_6102,N_4800,N_4788);
nand U6103 (N_6103,N_4533,N_4806);
or U6104 (N_6104,N_4465,N_3805);
nand U6105 (N_6105,N_3040,N_3055);
nand U6106 (N_6106,N_3472,N_2787);
nor U6107 (N_6107,N_3519,N_4965);
or U6108 (N_6108,N_4792,N_4783);
nand U6109 (N_6109,N_4310,N_4936);
nor U6110 (N_6110,N_4442,N_3053);
nor U6111 (N_6111,N_3577,N_3021);
or U6112 (N_6112,N_3016,N_4719);
nor U6113 (N_6113,N_4803,N_3510);
or U6114 (N_6114,N_3273,N_4640);
and U6115 (N_6115,N_4839,N_3093);
and U6116 (N_6116,N_3351,N_4297);
and U6117 (N_6117,N_2792,N_4504);
nor U6118 (N_6118,N_2634,N_2722);
nand U6119 (N_6119,N_2991,N_4959);
or U6120 (N_6120,N_3633,N_3563);
nand U6121 (N_6121,N_4867,N_2932);
nand U6122 (N_6122,N_4466,N_4017);
and U6123 (N_6123,N_4971,N_2785);
and U6124 (N_6124,N_4232,N_4260);
nand U6125 (N_6125,N_4076,N_3723);
or U6126 (N_6126,N_3500,N_4902);
nand U6127 (N_6127,N_3454,N_2899);
xnor U6128 (N_6128,N_3794,N_2902);
or U6129 (N_6129,N_4996,N_3884);
nor U6130 (N_6130,N_2728,N_3850);
nand U6131 (N_6131,N_3336,N_4630);
nor U6132 (N_6132,N_3573,N_3830);
or U6133 (N_6133,N_2577,N_3076);
and U6134 (N_6134,N_3113,N_3595);
nor U6135 (N_6135,N_4119,N_2651);
or U6136 (N_6136,N_3167,N_3314);
nand U6137 (N_6137,N_2580,N_4091);
nor U6138 (N_6138,N_3658,N_4793);
nand U6139 (N_6139,N_4795,N_3320);
or U6140 (N_6140,N_4363,N_2519);
nor U6141 (N_6141,N_3460,N_4213);
and U6142 (N_6142,N_3807,N_4861);
nor U6143 (N_6143,N_4392,N_4538);
or U6144 (N_6144,N_3477,N_3464);
nor U6145 (N_6145,N_3452,N_4904);
and U6146 (N_6146,N_2551,N_3765);
or U6147 (N_6147,N_4238,N_2670);
and U6148 (N_6148,N_3214,N_4905);
and U6149 (N_6149,N_3282,N_4077);
nand U6150 (N_6150,N_4614,N_3602);
nand U6151 (N_6151,N_4941,N_3610);
and U6152 (N_6152,N_4953,N_2766);
nand U6153 (N_6153,N_3594,N_3518);
and U6154 (N_6154,N_2545,N_4998);
xnor U6155 (N_6155,N_4003,N_3837);
nor U6156 (N_6156,N_2997,N_4390);
or U6157 (N_6157,N_3870,N_4347);
and U6158 (N_6158,N_3539,N_4512);
nand U6159 (N_6159,N_2508,N_3601);
nand U6160 (N_6160,N_4277,N_4883);
nand U6161 (N_6161,N_2716,N_3263);
nand U6162 (N_6162,N_4549,N_3551);
and U6163 (N_6163,N_4255,N_4388);
and U6164 (N_6164,N_4886,N_3064);
nand U6165 (N_6165,N_4349,N_4899);
and U6166 (N_6166,N_3882,N_3689);
or U6167 (N_6167,N_2814,N_2918);
nor U6168 (N_6168,N_3253,N_2738);
nand U6169 (N_6169,N_3160,N_3433);
or U6170 (N_6170,N_3086,N_4043);
or U6171 (N_6171,N_3888,N_3623);
and U6172 (N_6172,N_2841,N_4391);
xor U6173 (N_6173,N_2513,N_3033);
or U6174 (N_6174,N_4167,N_4436);
or U6175 (N_6175,N_3642,N_3264);
nand U6176 (N_6176,N_4850,N_2715);
nand U6177 (N_6177,N_3722,N_4711);
nand U6178 (N_6178,N_4340,N_4269);
and U6179 (N_6179,N_4276,N_2857);
or U6180 (N_6180,N_4567,N_4618);
nor U6181 (N_6181,N_4253,N_4509);
and U6182 (N_6182,N_2939,N_3071);
or U6183 (N_6183,N_4831,N_3759);
and U6184 (N_6184,N_2618,N_3287);
and U6185 (N_6185,N_4323,N_3724);
nand U6186 (N_6186,N_4339,N_4177);
xnor U6187 (N_6187,N_2705,N_4991);
or U6188 (N_6188,N_2936,N_3705);
and U6189 (N_6189,N_2637,N_3087);
or U6190 (N_6190,N_4524,N_2927);
and U6191 (N_6191,N_4123,N_3143);
nor U6192 (N_6192,N_4073,N_3907);
nand U6193 (N_6193,N_4170,N_2830);
nand U6194 (N_6194,N_4778,N_4633);
or U6195 (N_6195,N_2883,N_3036);
or U6196 (N_6196,N_3448,N_3469);
or U6197 (N_6197,N_3918,N_4705);
and U6198 (N_6198,N_3148,N_4973);
or U6199 (N_6199,N_3211,N_3993);
or U6200 (N_6200,N_3557,N_4145);
nor U6201 (N_6201,N_3716,N_4264);
and U6202 (N_6202,N_3229,N_4375);
nor U6203 (N_6203,N_4877,N_2579);
nor U6204 (N_6204,N_4956,N_4919);
xnor U6205 (N_6205,N_2717,N_3315);
nor U6206 (N_6206,N_4204,N_3905);
and U6207 (N_6207,N_4394,N_3824);
or U6208 (N_6208,N_4993,N_2574);
nor U6209 (N_6209,N_4894,N_3949);
nand U6210 (N_6210,N_4542,N_4072);
and U6211 (N_6211,N_4932,N_4147);
or U6212 (N_6212,N_3956,N_3415);
or U6213 (N_6213,N_3159,N_2735);
and U6214 (N_6214,N_4720,N_4006);
or U6215 (N_6215,N_2536,N_3906);
nor U6216 (N_6216,N_2799,N_3343);
nand U6217 (N_6217,N_3052,N_4967);
nor U6218 (N_6218,N_4115,N_3294);
xor U6219 (N_6219,N_2703,N_4234);
or U6220 (N_6220,N_3762,N_3416);
or U6221 (N_6221,N_3186,N_3653);
nor U6222 (N_6222,N_3298,N_4591);
and U6223 (N_6223,N_3420,N_2941);
nor U6224 (N_6224,N_3432,N_4892);
or U6225 (N_6225,N_4581,N_4889);
nand U6226 (N_6226,N_2994,N_3847);
nand U6227 (N_6227,N_4731,N_3032);
and U6228 (N_6228,N_4457,N_3576);
nor U6229 (N_6229,N_4153,N_4910);
and U6230 (N_6230,N_3340,N_4135);
nor U6231 (N_6231,N_4637,N_4824);
and U6232 (N_6232,N_4774,N_4078);
nor U6233 (N_6233,N_3665,N_3929);
or U6234 (N_6234,N_2575,N_3834);
and U6235 (N_6235,N_4035,N_3612);
and U6236 (N_6236,N_4501,N_3937);
nor U6237 (N_6237,N_2693,N_3915);
and U6238 (N_6238,N_2522,N_4433);
nand U6239 (N_6239,N_4667,N_4811);
nand U6240 (N_6240,N_3270,N_3357);
nor U6241 (N_6241,N_3235,N_3096);
nand U6242 (N_6242,N_3347,N_2621);
or U6243 (N_6243,N_4579,N_3981);
or U6244 (N_6244,N_3691,N_3215);
xor U6245 (N_6245,N_2563,N_2699);
nand U6246 (N_6246,N_3482,N_2546);
nor U6247 (N_6247,N_4748,N_3848);
nor U6248 (N_6248,N_3056,N_4588);
nor U6249 (N_6249,N_3172,N_2644);
nor U6250 (N_6250,N_3554,N_4754);
nor U6251 (N_6251,N_2826,N_3891);
and U6252 (N_6252,N_3053,N_3096);
and U6253 (N_6253,N_2605,N_4575);
nor U6254 (N_6254,N_3571,N_4345);
and U6255 (N_6255,N_4010,N_3914);
and U6256 (N_6256,N_4688,N_2539);
xor U6257 (N_6257,N_3147,N_4455);
or U6258 (N_6258,N_3570,N_4860);
nor U6259 (N_6259,N_3272,N_2861);
nor U6260 (N_6260,N_2769,N_2598);
and U6261 (N_6261,N_3785,N_2960);
nand U6262 (N_6262,N_3004,N_3697);
or U6263 (N_6263,N_2903,N_3180);
and U6264 (N_6264,N_4515,N_2695);
nor U6265 (N_6265,N_3092,N_4822);
nor U6266 (N_6266,N_4554,N_4150);
nor U6267 (N_6267,N_4939,N_3464);
nand U6268 (N_6268,N_4893,N_3778);
nand U6269 (N_6269,N_3910,N_4149);
nor U6270 (N_6270,N_3489,N_4091);
and U6271 (N_6271,N_4025,N_2527);
nand U6272 (N_6272,N_3868,N_4059);
or U6273 (N_6273,N_3957,N_4639);
nor U6274 (N_6274,N_3199,N_4941);
nor U6275 (N_6275,N_2577,N_3095);
xnor U6276 (N_6276,N_4947,N_4775);
and U6277 (N_6277,N_3193,N_3544);
or U6278 (N_6278,N_4359,N_4880);
nor U6279 (N_6279,N_3969,N_3771);
or U6280 (N_6280,N_3517,N_2943);
nor U6281 (N_6281,N_2918,N_2669);
and U6282 (N_6282,N_4446,N_4284);
nand U6283 (N_6283,N_4750,N_4918);
nand U6284 (N_6284,N_2641,N_4555);
nand U6285 (N_6285,N_3072,N_2919);
nand U6286 (N_6286,N_4957,N_4821);
nand U6287 (N_6287,N_4778,N_4513);
nor U6288 (N_6288,N_4200,N_4686);
nor U6289 (N_6289,N_3936,N_3659);
or U6290 (N_6290,N_3980,N_3847);
and U6291 (N_6291,N_3331,N_3549);
nand U6292 (N_6292,N_4949,N_4043);
or U6293 (N_6293,N_4778,N_4376);
and U6294 (N_6294,N_3242,N_3507);
nor U6295 (N_6295,N_4736,N_4933);
or U6296 (N_6296,N_3593,N_4668);
nand U6297 (N_6297,N_3399,N_4741);
nand U6298 (N_6298,N_4829,N_4945);
xor U6299 (N_6299,N_4311,N_3681);
nor U6300 (N_6300,N_4550,N_2988);
or U6301 (N_6301,N_2792,N_4382);
and U6302 (N_6302,N_3948,N_4644);
nand U6303 (N_6303,N_4068,N_4485);
and U6304 (N_6304,N_3494,N_4437);
or U6305 (N_6305,N_2606,N_2944);
or U6306 (N_6306,N_2661,N_4905);
or U6307 (N_6307,N_3431,N_4446);
nand U6308 (N_6308,N_3798,N_4201);
nand U6309 (N_6309,N_4630,N_3806);
or U6310 (N_6310,N_2590,N_3817);
or U6311 (N_6311,N_2911,N_3342);
nor U6312 (N_6312,N_2856,N_3734);
or U6313 (N_6313,N_3253,N_3885);
nor U6314 (N_6314,N_4668,N_3400);
nor U6315 (N_6315,N_4870,N_3202);
nand U6316 (N_6316,N_3812,N_4864);
and U6317 (N_6317,N_2602,N_2899);
nor U6318 (N_6318,N_2946,N_2549);
nor U6319 (N_6319,N_3960,N_3458);
nand U6320 (N_6320,N_4433,N_3076);
and U6321 (N_6321,N_2769,N_3123);
and U6322 (N_6322,N_4825,N_2881);
or U6323 (N_6323,N_3508,N_3684);
or U6324 (N_6324,N_2713,N_2813);
nor U6325 (N_6325,N_4107,N_3877);
nor U6326 (N_6326,N_4157,N_3218);
and U6327 (N_6327,N_3025,N_4587);
nor U6328 (N_6328,N_4707,N_3344);
and U6329 (N_6329,N_2922,N_3478);
nand U6330 (N_6330,N_4827,N_2993);
nand U6331 (N_6331,N_4156,N_3334);
nor U6332 (N_6332,N_4561,N_3260);
nand U6333 (N_6333,N_2973,N_4821);
or U6334 (N_6334,N_4790,N_3842);
nand U6335 (N_6335,N_3700,N_3462);
and U6336 (N_6336,N_3957,N_4375);
or U6337 (N_6337,N_3855,N_4163);
nand U6338 (N_6338,N_2925,N_3168);
nand U6339 (N_6339,N_2814,N_2790);
nand U6340 (N_6340,N_3977,N_4440);
nand U6341 (N_6341,N_4896,N_4198);
or U6342 (N_6342,N_4658,N_3212);
and U6343 (N_6343,N_4825,N_2690);
and U6344 (N_6344,N_4366,N_4095);
nor U6345 (N_6345,N_2857,N_4863);
nor U6346 (N_6346,N_3193,N_4811);
nand U6347 (N_6347,N_3094,N_3643);
or U6348 (N_6348,N_2782,N_4942);
and U6349 (N_6349,N_4237,N_2753);
nand U6350 (N_6350,N_4321,N_4463);
nor U6351 (N_6351,N_3957,N_4296);
and U6352 (N_6352,N_4899,N_2948);
and U6353 (N_6353,N_2675,N_3673);
nand U6354 (N_6354,N_2967,N_2506);
or U6355 (N_6355,N_3064,N_4139);
nand U6356 (N_6356,N_2693,N_3159);
or U6357 (N_6357,N_4017,N_4205);
nand U6358 (N_6358,N_3417,N_4307);
nand U6359 (N_6359,N_3436,N_3628);
nor U6360 (N_6360,N_4759,N_4068);
or U6361 (N_6361,N_2588,N_4203);
nand U6362 (N_6362,N_3758,N_4331);
and U6363 (N_6363,N_2549,N_4169);
or U6364 (N_6364,N_3405,N_4245);
nor U6365 (N_6365,N_3732,N_4388);
or U6366 (N_6366,N_4506,N_3248);
and U6367 (N_6367,N_2626,N_4133);
and U6368 (N_6368,N_4709,N_2569);
or U6369 (N_6369,N_3421,N_4967);
nand U6370 (N_6370,N_2805,N_4975);
nor U6371 (N_6371,N_4044,N_3475);
nand U6372 (N_6372,N_3678,N_4566);
nand U6373 (N_6373,N_3320,N_4067);
or U6374 (N_6374,N_2523,N_3507);
and U6375 (N_6375,N_4145,N_4948);
or U6376 (N_6376,N_4563,N_4131);
or U6377 (N_6377,N_3895,N_3832);
nand U6378 (N_6378,N_3068,N_4116);
nor U6379 (N_6379,N_3272,N_3343);
nand U6380 (N_6380,N_2720,N_4574);
and U6381 (N_6381,N_2806,N_3944);
xor U6382 (N_6382,N_3731,N_2891);
nor U6383 (N_6383,N_2552,N_2598);
nor U6384 (N_6384,N_3373,N_3845);
or U6385 (N_6385,N_4545,N_3858);
nand U6386 (N_6386,N_3128,N_3342);
and U6387 (N_6387,N_3300,N_4428);
and U6388 (N_6388,N_2852,N_3787);
or U6389 (N_6389,N_4041,N_3814);
and U6390 (N_6390,N_2813,N_4339);
nand U6391 (N_6391,N_3030,N_2536);
nor U6392 (N_6392,N_4983,N_3563);
or U6393 (N_6393,N_3801,N_4158);
or U6394 (N_6394,N_2980,N_4566);
nor U6395 (N_6395,N_4140,N_3636);
and U6396 (N_6396,N_3105,N_4613);
and U6397 (N_6397,N_3284,N_4750);
nor U6398 (N_6398,N_2836,N_4783);
and U6399 (N_6399,N_3339,N_4572);
and U6400 (N_6400,N_4455,N_2665);
and U6401 (N_6401,N_3873,N_3413);
nor U6402 (N_6402,N_2930,N_4197);
nor U6403 (N_6403,N_3835,N_3542);
nor U6404 (N_6404,N_4508,N_4275);
nand U6405 (N_6405,N_3755,N_2899);
nand U6406 (N_6406,N_4108,N_3367);
nor U6407 (N_6407,N_3339,N_4376);
and U6408 (N_6408,N_2766,N_2748);
and U6409 (N_6409,N_3761,N_3114);
nand U6410 (N_6410,N_2563,N_2947);
or U6411 (N_6411,N_4440,N_3121);
and U6412 (N_6412,N_3002,N_3917);
or U6413 (N_6413,N_4487,N_4706);
nor U6414 (N_6414,N_2691,N_2531);
nand U6415 (N_6415,N_4757,N_3122);
nand U6416 (N_6416,N_2720,N_2869);
or U6417 (N_6417,N_4716,N_3782);
and U6418 (N_6418,N_2832,N_4614);
nand U6419 (N_6419,N_3866,N_3992);
or U6420 (N_6420,N_4094,N_2557);
and U6421 (N_6421,N_4405,N_3214);
nand U6422 (N_6422,N_3944,N_3931);
and U6423 (N_6423,N_4140,N_4575);
or U6424 (N_6424,N_3454,N_2738);
and U6425 (N_6425,N_3972,N_3440);
nor U6426 (N_6426,N_4293,N_4904);
or U6427 (N_6427,N_2824,N_3591);
and U6428 (N_6428,N_3175,N_3904);
xnor U6429 (N_6429,N_2700,N_4154);
xnor U6430 (N_6430,N_4980,N_3574);
nand U6431 (N_6431,N_3897,N_4601);
and U6432 (N_6432,N_3509,N_3471);
and U6433 (N_6433,N_4586,N_4744);
and U6434 (N_6434,N_4562,N_4075);
nand U6435 (N_6435,N_4253,N_4868);
and U6436 (N_6436,N_3126,N_3263);
or U6437 (N_6437,N_2778,N_4350);
or U6438 (N_6438,N_4331,N_4807);
and U6439 (N_6439,N_4806,N_4739);
or U6440 (N_6440,N_2634,N_2702);
nand U6441 (N_6441,N_3557,N_3699);
nand U6442 (N_6442,N_2531,N_3860);
xor U6443 (N_6443,N_4331,N_2793);
and U6444 (N_6444,N_4345,N_4306);
xor U6445 (N_6445,N_4693,N_3682);
and U6446 (N_6446,N_4648,N_3148);
or U6447 (N_6447,N_4614,N_4475);
nor U6448 (N_6448,N_4290,N_4015);
nor U6449 (N_6449,N_4646,N_4141);
nor U6450 (N_6450,N_4248,N_4527);
or U6451 (N_6451,N_4395,N_4971);
and U6452 (N_6452,N_4593,N_3007);
nor U6453 (N_6453,N_3227,N_3712);
and U6454 (N_6454,N_4822,N_2939);
and U6455 (N_6455,N_3307,N_3900);
or U6456 (N_6456,N_4386,N_2772);
or U6457 (N_6457,N_4139,N_2809);
xnor U6458 (N_6458,N_4927,N_3176);
or U6459 (N_6459,N_3863,N_4707);
or U6460 (N_6460,N_3637,N_3131);
nand U6461 (N_6461,N_3049,N_2826);
nand U6462 (N_6462,N_3963,N_4879);
nor U6463 (N_6463,N_3721,N_3463);
or U6464 (N_6464,N_3246,N_4248);
nor U6465 (N_6465,N_3475,N_4776);
nor U6466 (N_6466,N_3148,N_2914);
and U6467 (N_6467,N_4405,N_4824);
or U6468 (N_6468,N_4873,N_3568);
or U6469 (N_6469,N_4903,N_3925);
or U6470 (N_6470,N_4534,N_4526);
nand U6471 (N_6471,N_2856,N_4753);
nand U6472 (N_6472,N_3526,N_3061);
or U6473 (N_6473,N_4077,N_4852);
or U6474 (N_6474,N_3432,N_4342);
and U6475 (N_6475,N_4923,N_4519);
nor U6476 (N_6476,N_4294,N_3924);
and U6477 (N_6477,N_3706,N_2773);
nand U6478 (N_6478,N_3868,N_4233);
and U6479 (N_6479,N_4188,N_4540);
nor U6480 (N_6480,N_2955,N_3856);
nand U6481 (N_6481,N_4496,N_2610);
nor U6482 (N_6482,N_2690,N_3032);
xnor U6483 (N_6483,N_3598,N_3414);
nor U6484 (N_6484,N_3326,N_4032);
and U6485 (N_6485,N_3619,N_3131);
nand U6486 (N_6486,N_4371,N_4070);
nand U6487 (N_6487,N_4077,N_3817);
and U6488 (N_6488,N_3027,N_2627);
nor U6489 (N_6489,N_3441,N_3823);
nand U6490 (N_6490,N_4013,N_3668);
and U6491 (N_6491,N_4310,N_3113);
nor U6492 (N_6492,N_3575,N_2539);
and U6493 (N_6493,N_2799,N_2814);
and U6494 (N_6494,N_4911,N_2630);
nand U6495 (N_6495,N_3624,N_2698);
and U6496 (N_6496,N_4544,N_4914);
and U6497 (N_6497,N_2768,N_4979);
nor U6498 (N_6498,N_3265,N_3472);
or U6499 (N_6499,N_4375,N_4891);
nor U6500 (N_6500,N_3074,N_3030);
nor U6501 (N_6501,N_2952,N_4859);
or U6502 (N_6502,N_4925,N_4640);
nand U6503 (N_6503,N_3110,N_4962);
nand U6504 (N_6504,N_4216,N_4631);
nor U6505 (N_6505,N_2881,N_4471);
nor U6506 (N_6506,N_3265,N_4199);
nor U6507 (N_6507,N_2865,N_3443);
and U6508 (N_6508,N_3979,N_2589);
nand U6509 (N_6509,N_3677,N_4998);
nand U6510 (N_6510,N_3459,N_4014);
xnor U6511 (N_6511,N_2823,N_2688);
or U6512 (N_6512,N_3659,N_2897);
or U6513 (N_6513,N_4428,N_2845);
nand U6514 (N_6514,N_2763,N_4026);
and U6515 (N_6515,N_2777,N_3398);
nand U6516 (N_6516,N_3739,N_4321);
and U6517 (N_6517,N_3102,N_4766);
or U6518 (N_6518,N_3593,N_4542);
and U6519 (N_6519,N_3702,N_4291);
and U6520 (N_6520,N_4136,N_3603);
nor U6521 (N_6521,N_3216,N_4255);
or U6522 (N_6522,N_4150,N_3336);
nor U6523 (N_6523,N_3881,N_2851);
nor U6524 (N_6524,N_2861,N_4887);
or U6525 (N_6525,N_2646,N_3050);
and U6526 (N_6526,N_4682,N_4997);
nand U6527 (N_6527,N_4322,N_3303);
nand U6528 (N_6528,N_2540,N_3916);
xor U6529 (N_6529,N_2537,N_4784);
nand U6530 (N_6530,N_3268,N_4953);
or U6531 (N_6531,N_4597,N_3755);
nand U6532 (N_6532,N_3357,N_3295);
and U6533 (N_6533,N_4408,N_4208);
nand U6534 (N_6534,N_4089,N_2885);
nor U6535 (N_6535,N_3834,N_3167);
or U6536 (N_6536,N_4745,N_2654);
and U6537 (N_6537,N_2651,N_3854);
or U6538 (N_6538,N_3510,N_4971);
or U6539 (N_6539,N_3065,N_4166);
nor U6540 (N_6540,N_4453,N_4259);
nor U6541 (N_6541,N_3412,N_2878);
or U6542 (N_6542,N_4692,N_3120);
and U6543 (N_6543,N_4357,N_2782);
nor U6544 (N_6544,N_4225,N_4783);
and U6545 (N_6545,N_2562,N_3988);
nand U6546 (N_6546,N_3673,N_3134);
or U6547 (N_6547,N_3055,N_4943);
or U6548 (N_6548,N_4220,N_4981);
or U6549 (N_6549,N_3959,N_3044);
or U6550 (N_6550,N_2545,N_3097);
nand U6551 (N_6551,N_2519,N_3031);
and U6552 (N_6552,N_2659,N_4058);
and U6553 (N_6553,N_4065,N_3873);
nor U6554 (N_6554,N_4189,N_4342);
nand U6555 (N_6555,N_4502,N_4614);
nor U6556 (N_6556,N_3700,N_2723);
or U6557 (N_6557,N_4608,N_4453);
nor U6558 (N_6558,N_4751,N_4017);
or U6559 (N_6559,N_4713,N_2607);
nor U6560 (N_6560,N_4828,N_3194);
nor U6561 (N_6561,N_3271,N_2888);
nor U6562 (N_6562,N_2570,N_3267);
nand U6563 (N_6563,N_4424,N_3773);
and U6564 (N_6564,N_4218,N_4056);
nand U6565 (N_6565,N_2967,N_4472);
or U6566 (N_6566,N_4390,N_3251);
nand U6567 (N_6567,N_2963,N_3996);
and U6568 (N_6568,N_4872,N_3365);
nor U6569 (N_6569,N_3734,N_4721);
or U6570 (N_6570,N_2650,N_3356);
nand U6571 (N_6571,N_4154,N_3086);
nand U6572 (N_6572,N_3258,N_4937);
nand U6573 (N_6573,N_4425,N_3271);
and U6574 (N_6574,N_2883,N_4579);
nand U6575 (N_6575,N_4616,N_2516);
nand U6576 (N_6576,N_4037,N_3039);
nand U6577 (N_6577,N_4084,N_3444);
or U6578 (N_6578,N_3200,N_3293);
or U6579 (N_6579,N_2858,N_2633);
and U6580 (N_6580,N_2505,N_4394);
or U6581 (N_6581,N_2889,N_3114);
and U6582 (N_6582,N_4317,N_2848);
nand U6583 (N_6583,N_2530,N_3746);
or U6584 (N_6584,N_2961,N_3959);
xor U6585 (N_6585,N_2723,N_3549);
nor U6586 (N_6586,N_4808,N_4706);
nor U6587 (N_6587,N_3062,N_3337);
and U6588 (N_6588,N_3365,N_4306);
nor U6589 (N_6589,N_3996,N_4730);
nand U6590 (N_6590,N_2594,N_3540);
and U6591 (N_6591,N_3472,N_3300);
nand U6592 (N_6592,N_3988,N_4282);
nand U6593 (N_6593,N_4720,N_2566);
nand U6594 (N_6594,N_3675,N_2512);
xor U6595 (N_6595,N_3113,N_4812);
nand U6596 (N_6596,N_3484,N_3470);
nand U6597 (N_6597,N_3909,N_3646);
or U6598 (N_6598,N_2869,N_3904);
nor U6599 (N_6599,N_2734,N_3922);
and U6600 (N_6600,N_4585,N_3850);
nand U6601 (N_6601,N_3295,N_4466);
nand U6602 (N_6602,N_4323,N_3108);
nand U6603 (N_6603,N_3212,N_3143);
nor U6604 (N_6604,N_3904,N_2620);
nor U6605 (N_6605,N_2952,N_3010);
nor U6606 (N_6606,N_4249,N_4597);
or U6607 (N_6607,N_4651,N_4857);
nor U6608 (N_6608,N_4003,N_4886);
nand U6609 (N_6609,N_4144,N_3492);
nor U6610 (N_6610,N_4568,N_4567);
nand U6611 (N_6611,N_4083,N_4865);
nand U6612 (N_6612,N_2810,N_3326);
nor U6613 (N_6613,N_3837,N_4231);
nor U6614 (N_6614,N_4714,N_3578);
nor U6615 (N_6615,N_4321,N_4478);
and U6616 (N_6616,N_4247,N_2967);
or U6617 (N_6617,N_4560,N_2590);
and U6618 (N_6618,N_3597,N_3868);
or U6619 (N_6619,N_4139,N_3856);
and U6620 (N_6620,N_3658,N_3460);
nor U6621 (N_6621,N_3505,N_2937);
and U6622 (N_6622,N_3520,N_2512);
nor U6623 (N_6623,N_4078,N_4566);
nor U6624 (N_6624,N_4313,N_3509);
and U6625 (N_6625,N_2699,N_4601);
nand U6626 (N_6626,N_2795,N_3154);
nor U6627 (N_6627,N_2502,N_3890);
nor U6628 (N_6628,N_3996,N_3770);
nor U6629 (N_6629,N_3318,N_3860);
or U6630 (N_6630,N_2637,N_3725);
xor U6631 (N_6631,N_4711,N_2534);
or U6632 (N_6632,N_4833,N_4232);
or U6633 (N_6633,N_4049,N_3474);
and U6634 (N_6634,N_3692,N_3119);
nor U6635 (N_6635,N_4152,N_3104);
or U6636 (N_6636,N_3935,N_4871);
nor U6637 (N_6637,N_2597,N_3538);
xnor U6638 (N_6638,N_4274,N_3638);
or U6639 (N_6639,N_3155,N_2519);
and U6640 (N_6640,N_3954,N_4268);
and U6641 (N_6641,N_4499,N_3440);
nand U6642 (N_6642,N_3685,N_2788);
and U6643 (N_6643,N_4963,N_4416);
nand U6644 (N_6644,N_2995,N_4708);
and U6645 (N_6645,N_3737,N_3293);
nand U6646 (N_6646,N_3572,N_3462);
nor U6647 (N_6647,N_4836,N_3669);
and U6648 (N_6648,N_3523,N_4116);
nand U6649 (N_6649,N_4442,N_2953);
nand U6650 (N_6650,N_2835,N_3128);
xnor U6651 (N_6651,N_4157,N_4420);
nand U6652 (N_6652,N_3744,N_3813);
or U6653 (N_6653,N_4495,N_3868);
or U6654 (N_6654,N_4880,N_3518);
nor U6655 (N_6655,N_4760,N_3963);
nand U6656 (N_6656,N_3305,N_3394);
xor U6657 (N_6657,N_4019,N_2960);
and U6658 (N_6658,N_4662,N_4694);
xnor U6659 (N_6659,N_3878,N_4134);
nor U6660 (N_6660,N_3618,N_2605);
nand U6661 (N_6661,N_3181,N_3302);
nor U6662 (N_6662,N_3629,N_4401);
and U6663 (N_6663,N_3416,N_3604);
and U6664 (N_6664,N_4792,N_3934);
or U6665 (N_6665,N_4273,N_3742);
nand U6666 (N_6666,N_4448,N_2652);
nor U6667 (N_6667,N_4502,N_3982);
nand U6668 (N_6668,N_4795,N_3644);
or U6669 (N_6669,N_4856,N_4747);
and U6670 (N_6670,N_4285,N_4078);
and U6671 (N_6671,N_3834,N_3975);
nor U6672 (N_6672,N_3656,N_4337);
and U6673 (N_6673,N_4196,N_4331);
and U6674 (N_6674,N_4834,N_2989);
nor U6675 (N_6675,N_3718,N_4156);
nand U6676 (N_6676,N_2897,N_4599);
and U6677 (N_6677,N_3833,N_3668);
or U6678 (N_6678,N_4176,N_3853);
or U6679 (N_6679,N_2966,N_4575);
or U6680 (N_6680,N_4818,N_3155);
nand U6681 (N_6681,N_4496,N_4778);
nand U6682 (N_6682,N_4389,N_2669);
and U6683 (N_6683,N_3933,N_3768);
xor U6684 (N_6684,N_2673,N_3726);
or U6685 (N_6685,N_4623,N_4319);
nand U6686 (N_6686,N_2897,N_3942);
nand U6687 (N_6687,N_2762,N_3158);
nor U6688 (N_6688,N_4104,N_2707);
nor U6689 (N_6689,N_4446,N_4610);
xor U6690 (N_6690,N_3684,N_4276);
nand U6691 (N_6691,N_4728,N_3082);
or U6692 (N_6692,N_4318,N_3563);
and U6693 (N_6693,N_4191,N_2984);
nor U6694 (N_6694,N_4171,N_3984);
nand U6695 (N_6695,N_4516,N_2790);
nor U6696 (N_6696,N_3754,N_3672);
and U6697 (N_6697,N_4362,N_3061);
nor U6698 (N_6698,N_2879,N_3134);
or U6699 (N_6699,N_3233,N_3493);
or U6700 (N_6700,N_4702,N_4302);
nor U6701 (N_6701,N_4415,N_4086);
nand U6702 (N_6702,N_2862,N_4051);
or U6703 (N_6703,N_3551,N_4607);
nand U6704 (N_6704,N_4254,N_2950);
and U6705 (N_6705,N_4790,N_3673);
and U6706 (N_6706,N_4622,N_4441);
or U6707 (N_6707,N_2506,N_3644);
or U6708 (N_6708,N_3634,N_4853);
xor U6709 (N_6709,N_2767,N_2928);
and U6710 (N_6710,N_3855,N_3047);
nand U6711 (N_6711,N_2918,N_3344);
nand U6712 (N_6712,N_4262,N_4556);
nand U6713 (N_6713,N_4286,N_3132);
nor U6714 (N_6714,N_3070,N_2804);
nor U6715 (N_6715,N_2971,N_3318);
or U6716 (N_6716,N_3566,N_3839);
and U6717 (N_6717,N_3007,N_3364);
xnor U6718 (N_6718,N_3397,N_4128);
nand U6719 (N_6719,N_2633,N_4479);
or U6720 (N_6720,N_4804,N_3337);
and U6721 (N_6721,N_3066,N_4070);
xor U6722 (N_6722,N_3781,N_3171);
and U6723 (N_6723,N_4665,N_2505);
nor U6724 (N_6724,N_4854,N_3681);
nand U6725 (N_6725,N_4869,N_4113);
nor U6726 (N_6726,N_4577,N_2974);
nand U6727 (N_6727,N_4912,N_3394);
nor U6728 (N_6728,N_4268,N_4507);
or U6729 (N_6729,N_3208,N_4218);
and U6730 (N_6730,N_4385,N_4619);
nor U6731 (N_6731,N_2970,N_4969);
and U6732 (N_6732,N_3533,N_4070);
or U6733 (N_6733,N_2847,N_2917);
and U6734 (N_6734,N_4756,N_4473);
and U6735 (N_6735,N_3979,N_2720);
or U6736 (N_6736,N_4006,N_2963);
and U6737 (N_6737,N_4036,N_2951);
or U6738 (N_6738,N_3123,N_2629);
or U6739 (N_6739,N_3319,N_3410);
nand U6740 (N_6740,N_3401,N_3353);
nor U6741 (N_6741,N_3021,N_2546);
or U6742 (N_6742,N_2582,N_4478);
and U6743 (N_6743,N_4142,N_2503);
or U6744 (N_6744,N_3539,N_4473);
and U6745 (N_6745,N_4234,N_4889);
or U6746 (N_6746,N_4409,N_2825);
or U6747 (N_6747,N_4802,N_3567);
nand U6748 (N_6748,N_4266,N_2521);
and U6749 (N_6749,N_3962,N_4769);
or U6750 (N_6750,N_3445,N_4255);
and U6751 (N_6751,N_4905,N_4086);
and U6752 (N_6752,N_2940,N_4706);
nor U6753 (N_6753,N_3572,N_3615);
or U6754 (N_6754,N_2988,N_2627);
nand U6755 (N_6755,N_4815,N_3772);
or U6756 (N_6756,N_4317,N_4762);
and U6757 (N_6757,N_4979,N_4004);
nor U6758 (N_6758,N_3795,N_3159);
or U6759 (N_6759,N_4495,N_4741);
or U6760 (N_6760,N_4024,N_4957);
nand U6761 (N_6761,N_2945,N_2605);
and U6762 (N_6762,N_2712,N_2875);
or U6763 (N_6763,N_3690,N_2611);
and U6764 (N_6764,N_2642,N_4788);
nand U6765 (N_6765,N_4891,N_3390);
and U6766 (N_6766,N_3649,N_2813);
and U6767 (N_6767,N_3630,N_3925);
and U6768 (N_6768,N_3228,N_4489);
nand U6769 (N_6769,N_3170,N_3603);
nor U6770 (N_6770,N_2798,N_2650);
xnor U6771 (N_6771,N_4395,N_4019);
or U6772 (N_6772,N_4387,N_3984);
xnor U6773 (N_6773,N_3130,N_2548);
nand U6774 (N_6774,N_3185,N_2991);
or U6775 (N_6775,N_4744,N_2872);
or U6776 (N_6776,N_4876,N_4116);
nand U6777 (N_6777,N_4417,N_4946);
or U6778 (N_6778,N_3943,N_2531);
xor U6779 (N_6779,N_4818,N_4355);
nand U6780 (N_6780,N_3937,N_2894);
or U6781 (N_6781,N_3495,N_2849);
or U6782 (N_6782,N_4127,N_4287);
nor U6783 (N_6783,N_4969,N_4123);
nor U6784 (N_6784,N_2846,N_4681);
xnor U6785 (N_6785,N_4445,N_4904);
or U6786 (N_6786,N_4069,N_3702);
nor U6787 (N_6787,N_4914,N_4656);
nor U6788 (N_6788,N_4453,N_3281);
nand U6789 (N_6789,N_3970,N_4441);
nor U6790 (N_6790,N_4238,N_4685);
nor U6791 (N_6791,N_4860,N_2746);
and U6792 (N_6792,N_4404,N_3628);
nor U6793 (N_6793,N_3702,N_4682);
xor U6794 (N_6794,N_3884,N_2658);
nor U6795 (N_6795,N_3547,N_2850);
nor U6796 (N_6796,N_2510,N_2821);
or U6797 (N_6797,N_2999,N_4128);
and U6798 (N_6798,N_3861,N_4209);
and U6799 (N_6799,N_3036,N_4804);
nand U6800 (N_6800,N_3601,N_2798);
nor U6801 (N_6801,N_2510,N_4911);
nand U6802 (N_6802,N_4777,N_4652);
nor U6803 (N_6803,N_4807,N_4003);
and U6804 (N_6804,N_2568,N_4739);
nor U6805 (N_6805,N_3635,N_2900);
nor U6806 (N_6806,N_3607,N_2563);
nor U6807 (N_6807,N_2691,N_3858);
and U6808 (N_6808,N_2727,N_4794);
nand U6809 (N_6809,N_3002,N_2715);
nor U6810 (N_6810,N_3085,N_3947);
nand U6811 (N_6811,N_4880,N_3205);
nand U6812 (N_6812,N_4090,N_3661);
xor U6813 (N_6813,N_3565,N_2752);
nand U6814 (N_6814,N_2642,N_3680);
nand U6815 (N_6815,N_3637,N_4120);
nand U6816 (N_6816,N_4356,N_3155);
and U6817 (N_6817,N_4033,N_4799);
or U6818 (N_6818,N_2903,N_4122);
nor U6819 (N_6819,N_3704,N_4646);
or U6820 (N_6820,N_3738,N_2651);
nor U6821 (N_6821,N_4668,N_3017);
and U6822 (N_6822,N_3267,N_4041);
and U6823 (N_6823,N_2583,N_4928);
or U6824 (N_6824,N_4408,N_4055);
nor U6825 (N_6825,N_4122,N_4825);
and U6826 (N_6826,N_3109,N_3031);
and U6827 (N_6827,N_2527,N_3035);
nand U6828 (N_6828,N_3442,N_3637);
nand U6829 (N_6829,N_2721,N_4017);
nand U6830 (N_6830,N_4928,N_3733);
nand U6831 (N_6831,N_4709,N_3722);
nor U6832 (N_6832,N_4880,N_4490);
or U6833 (N_6833,N_3026,N_4152);
or U6834 (N_6834,N_3148,N_4019);
nor U6835 (N_6835,N_3023,N_4972);
and U6836 (N_6836,N_2612,N_3645);
and U6837 (N_6837,N_2811,N_3451);
and U6838 (N_6838,N_2597,N_3702);
and U6839 (N_6839,N_3395,N_2568);
or U6840 (N_6840,N_4743,N_3658);
and U6841 (N_6841,N_3668,N_3239);
nor U6842 (N_6842,N_3538,N_3359);
or U6843 (N_6843,N_3516,N_4627);
nand U6844 (N_6844,N_2715,N_4828);
or U6845 (N_6845,N_4853,N_4974);
nand U6846 (N_6846,N_4345,N_4686);
or U6847 (N_6847,N_2885,N_2952);
nand U6848 (N_6848,N_4754,N_3551);
nor U6849 (N_6849,N_3519,N_3548);
xnor U6850 (N_6850,N_4006,N_3629);
nor U6851 (N_6851,N_4977,N_4535);
nor U6852 (N_6852,N_2614,N_2914);
or U6853 (N_6853,N_4039,N_4234);
nor U6854 (N_6854,N_4507,N_2843);
or U6855 (N_6855,N_2513,N_3383);
or U6856 (N_6856,N_3781,N_4361);
or U6857 (N_6857,N_3570,N_4405);
nor U6858 (N_6858,N_3909,N_4328);
nand U6859 (N_6859,N_2525,N_4476);
nand U6860 (N_6860,N_4042,N_2939);
or U6861 (N_6861,N_2870,N_3648);
or U6862 (N_6862,N_3264,N_3077);
and U6863 (N_6863,N_2509,N_4800);
and U6864 (N_6864,N_4664,N_3243);
nand U6865 (N_6865,N_3821,N_2685);
and U6866 (N_6866,N_2982,N_3703);
xor U6867 (N_6867,N_2661,N_4757);
nor U6868 (N_6868,N_2866,N_3864);
or U6869 (N_6869,N_2640,N_4833);
nor U6870 (N_6870,N_3082,N_3614);
or U6871 (N_6871,N_4325,N_3421);
or U6872 (N_6872,N_4330,N_3767);
and U6873 (N_6873,N_3679,N_4796);
nand U6874 (N_6874,N_2826,N_4259);
or U6875 (N_6875,N_3795,N_4322);
or U6876 (N_6876,N_3298,N_3961);
xnor U6877 (N_6877,N_4693,N_2573);
and U6878 (N_6878,N_4343,N_3802);
nor U6879 (N_6879,N_4577,N_4329);
nor U6880 (N_6880,N_2656,N_3765);
and U6881 (N_6881,N_3773,N_3128);
and U6882 (N_6882,N_4124,N_4277);
nor U6883 (N_6883,N_2529,N_3131);
nor U6884 (N_6884,N_3010,N_2543);
nor U6885 (N_6885,N_3893,N_3125);
nor U6886 (N_6886,N_2568,N_4580);
or U6887 (N_6887,N_3061,N_4213);
and U6888 (N_6888,N_2574,N_4162);
and U6889 (N_6889,N_2667,N_3916);
nand U6890 (N_6890,N_3237,N_4404);
nor U6891 (N_6891,N_3699,N_2948);
nand U6892 (N_6892,N_2562,N_3087);
or U6893 (N_6893,N_4435,N_4897);
nor U6894 (N_6894,N_3016,N_2626);
nand U6895 (N_6895,N_2837,N_4484);
or U6896 (N_6896,N_4138,N_4625);
nor U6897 (N_6897,N_4926,N_3632);
or U6898 (N_6898,N_3504,N_3545);
and U6899 (N_6899,N_4442,N_4070);
nor U6900 (N_6900,N_3354,N_2582);
and U6901 (N_6901,N_4033,N_3091);
or U6902 (N_6902,N_4075,N_3351);
and U6903 (N_6903,N_3659,N_4087);
nand U6904 (N_6904,N_4594,N_4994);
nand U6905 (N_6905,N_2542,N_3878);
nand U6906 (N_6906,N_3743,N_4752);
and U6907 (N_6907,N_2990,N_4167);
nand U6908 (N_6908,N_3556,N_4710);
or U6909 (N_6909,N_4120,N_3288);
or U6910 (N_6910,N_4703,N_3824);
nand U6911 (N_6911,N_2863,N_4524);
nand U6912 (N_6912,N_3842,N_2570);
nand U6913 (N_6913,N_3212,N_2840);
nor U6914 (N_6914,N_2607,N_3430);
nand U6915 (N_6915,N_4719,N_4365);
nand U6916 (N_6916,N_4114,N_4249);
and U6917 (N_6917,N_3294,N_3623);
or U6918 (N_6918,N_3225,N_3476);
nor U6919 (N_6919,N_3625,N_2863);
nor U6920 (N_6920,N_4163,N_3188);
nand U6921 (N_6921,N_3367,N_4617);
nand U6922 (N_6922,N_4647,N_4974);
or U6923 (N_6923,N_3981,N_3940);
and U6924 (N_6924,N_3840,N_4447);
and U6925 (N_6925,N_4449,N_4565);
and U6926 (N_6926,N_3840,N_4478);
nand U6927 (N_6927,N_4788,N_4041);
or U6928 (N_6928,N_3355,N_2804);
nor U6929 (N_6929,N_4822,N_4461);
or U6930 (N_6930,N_2647,N_3915);
nand U6931 (N_6931,N_3688,N_2734);
or U6932 (N_6932,N_3061,N_3798);
and U6933 (N_6933,N_3533,N_3723);
nor U6934 (N_6934,N_3416,N_4367);
or U6935 (N_6935,N_4938,N_4513);
or U6936 (N_6936,N_3364,N_4353);
or U6937 (N_6937,N_2919,N_4788);
or U6938 (N_6938,N_2757,N_3935);
nor U6939 (N_6939,N_3007,N_4955);
nand U6940 (N_6940,N_4248,N_2687);
nor U6941 (N_6941,N_3016,N_2973);
nand U6942 (N_6942,N_3785,N_3507);
nor U6943 (N_6943,N_3484,N_4938);
nor U6944 (N_6944,N_3278,N_3780);
nand U6945 (N_6945,N_4079,N_2597);
or U6946 (N_6946,N_3940,N_4256);
nor U6947 (N_6947,N_3983,N_4643);
and U6948 (N_6948,N_2848,N_2782);
or U6949 (N_6949,N_3657,N_3050);
nand U6950 (N_6950,N_3950,N_3407);
and U6951 (N_6951,N_3559,N_4296);
or U6952 (N_6952,N_3765,N_3946);
or U6953 (N_6953,N_4816,N_4313);
nand U6954 (N_6954,N_3748,N_4760);
nor U6955 (N_6955,N_2538,N_2776);
nor U6956 (N_6956,N_3011,N_2669);
nor U6957 (N_6957,N_3963,N_4794);
and U6958 (N_6958,N_3262,N_3603);
nor U6959 (N_6959,N_3012,N_4581);
nand U6960 (N_6960,N_3715,N_4403);
nor U6961 (N_6961,N_2937,N_4389);
nor U6962 (N_6962,N_2740,N_3223);
and U6963 (N_6963,N_3562,N_2711);
and U6964 (N_6964,N_4819,N_4650);
nor U6965 (N_6965,N_3598,N_3706);
or U6966 (N_6966,N_3605,N_2523);
xnor U6967 (N_6967,N_3674,N_4456);
or U6968 (N_6968,N_3616,N_4873);
nand U6969 (N_6969,N_3557,N_3951);
nor U6970 (N_6970,N_3426,N_4978);
nor U6971 (N_6971,N_4345,N_4240);
or U6972 (N_6972,N_3651,N_3068);
nand U6973 (N_6973,N_3711,N_4622);
or U6974 (N_6974,N_3373,N_3667);
nand U6975 (N_6975,N_3618,N_4850);
or U6976 (N_6976,N_4717,N_3305);
and U6977 (N_6977,N_3397,N_2765);
or U6978 (N_6978,N_3094,N_4809);
and U6979 (N_6979,N_4320,N_3863);
nor U6980 (N_6980,N_3661,N_4172);
nand U6981 (N_6981,N_4578,N_2866);
or U6982 (N_6982,N_2555,N_4957);
nand U6983 (N_6983,N_2618,N_4641);
nor U6984 (N_6984,N_3366,N_4011);
and U6985 (N_6985,N_4779,N_2698);
nor U6986 (N_6986,N_4225,N_4938);
nor U6987 (N_6987,N_3826,N_4372);
nor U6988 (N_6988,N_4042,N_4954);
and U6989 (N_6989,N_3669,N_4942);
and U6990 (N_6990,N_4031,N_3864);
nor U6991 (N_6991,N_4512,N_3619);
and U6992 (N_6992,N_2993,N_2615);
or U6993 (N_6993,N_4926,N_2550);
nor U6994 (N_6994,N_4053,N_3573);
nor U6995 (N_6995,N_4159,N_4242);
nor U6996 (N_6996,N_4769,N_2524);
xnor U6997 (N_6997,N_4823,N_4449);
and U6998 (N_6998,N_3936,N_2544);
and U6999 (N_6999,N_2745,N_3453);
or U7000 (N_7000,N_4667,N_3285);
or U7001 (N_7001,N_4472,N_4145);
nand U7002 (N_7002,N_3144,N_2908);
nor U7003 (N_7003,N_4151,N_4916);
nand U7004 (N_7004,N_3546,N_4012);
nand U7005 (N_7005,N_3781,N_3816);
nor U7006 (N_7006,N_2938,N_4019);
and U7007 (N_7007,N_2556,N_3416);
and U7008 (N_7008,N_4328,N_3576);
and U7009 (N_7009,N_2663,N_4588);
and U7010 (N_7010,N_3897,N_4670);
and U7011 (N_7011,N_4159,N_3289);
or U7012 (N_7012,N_3056,N_4677);
nor U7013 (N_7013,N_3883,N_2689);
nand U7014 (N_7014,N_2727,N_4183);
nand U7015 (N_7015,N_3432,N_2742);
or U7016 (N_7016,N_2905,N_4515);
nor U7017 (N_7017,N_4171,N_4568);
or U7018 (N_7018,N_3448,N_3318);
nor U7019 (N_7019,N_3706,N_2677);
nor U7020 (N_7020,N_2849,N_4572);
nor U7021 (N_7021,N_3164,N_3148);
nand U7022 (N_7022,N_3903,N_3294);
or U7023 (N_7023,N_4879,N_4800);
and U7024 (N_7024,N_3863,N_3945);
or U7025 (N_7025,N_2710,N_4784);
or U7026 (N_7026,N_2964,N_4678);
nor U7027 (N_7027,N_3873,N_4683);
or U7028 (N_7028,N_3595,N_4695);
nor U7029 (N_7029,N_3344,N_4772);
nor U7030 (N_7030,N_4077,N_3645);
nand U7031 (N_7031,N_3172,N_3545);
nand U7032 (N_7032,N_3123,N_3714);
and U7033 (N_7033,N_4148,N_4440);
nand U7034 (N_7034,N_3512,N_4880);
or U7035 (N_7035,N_4982,N_2648);
nand U7036 (N_7036,N_4582,N_3331);
nor U7037 (N_7037,N_3642,N_3057);
nor U7038 (N_7038,N_4700,N_2620);
or U7039 (N_7039,N_2622,N_2767);
nand U7040 (N_7040,N_3766,N_4899);
nor U7041 (N_7041,N_3323,N_3013);
or U7042 (N_7042,N_3259,N_3948);
nand U7043 (N_7043,N_4822,N_4601);
and U7044 (N_7044,N_4781,N_4577);
and U7045 (N_7045,N_2668,N_4233);
or U7046 (N_7046,N_3296,N_2775);
or U7047 (N_7047,N_4923,N_4241);
or U7048 (N_7048,N_3502,N_4881);
nand U7049 (N_7049,N_3567,N_4274);
or U7050 (N_7050,N_3990,N_4534);
or U7051 (N_7051,N_2585,N_4384);
nand U7052 (N_7052,N_3307,N_4700);
nand U7053 (N_7053,N_4822,N_4295);
and U7054 (N_7054,N_4849,N_2717);
and U7055 (N_7055,N_2856,N_4629);
or U7056 (N_7056,N_4171,N_4781);
and U7057 (N_7057,N_3341,N_3140);
nand U7058 (N_7058,N_3685,N_2632);
nor U7059 (N_7059,N_3476,N_3296);
nor U7060 (N_7060,N_2930,N_2724);
and U7061 (N_7061,N_2985,N_4923);
and U7062 (N_7062,N_2809,N_4540);
nand U7063 (N_7063,N_3771,N_3702);
and U7064 (N_7064,N_3607,N_4520);
or U7065 (N_7065,N_3693,N_3316);
nand U7066 (N_7066,N_3250,N_3397);
and U7067 (N_7067,N_4368,N_4967);
and U7068 (N_7068,N_3856,N_4433);
and U7069 (N_7069,N_3328,N_2524);
and U7070 (N_7070,N_2615,N_4855);
nor U7071 (N_7071,N_3024,N_2943);
or U7072 (N_7072,N_3499,N_3100);
nor U7073 (N_7073,N_4526,N_3772);
nand U7074 (N_7074,N_4867,N_4053);
nand U7075 (N_7075,N_4517,N_3234);
and U7076 (N_7076,N_3568,N_3105);
nor U7077 (N_7077,N_3899,N_4876);
nand U7078 (N_7078,N_2721,N_4870);
nor U7079 (N_7079,N_4359,N_4076);
or U7080 (N_7080,N_4583,N_4488);
and U7081 (N_7081,N_2532,N_3548);
nand U7082 (N_7082,N_4742,N_2952);
nand U7083 (N_7083,N_4923,N_3341);
nor U7084 (N_7084,N_3959,N_4588);
and U7085 (N_7085,N_4649,N_3311);
nand U7086 (N_7086,N_2767,N_2575);
nand U7087 (N_7087,N_3095,N_3470);
or U7088 (N_7088,N_2642,N_4952);
nand U7089 (N_7089,N_4392,N_2884);
and U7090 (N_7090,N_2597,N_4736);
nand U7091 (N_7091,N_2617,N_4741);
nor U7092 (N_7092,N_3138,N_4711);
nor U7093 (N_7093,N_4649,N_4443);
or U7094 (N_7094,N_3292,N_3191);
nand U7095 (N_7095,N_3661,N_3428);
and U7096 (N_7096,N_3395,N_2787);
and U7097 (N_7097,N_2960,N_2907);
or U7098 (N_7098,N_3288,N_3277);
and U7099 (N_7099,N_4712,N_3125);
and U7100 (N_7100,N_3330,N_3340);
nor U7101 (N_7101,N_3430,N_2892);
or U7102 (N_7102,N_3059,N_4363);
nor U7103 (N_7103,N_3940,N_3211);
and U7104 (N_7104,N_3297,N_3546);
and U7105 (N_7105,N_2941,N_3101);
nand U7106 (N_7106,N_2872,N_3716);
nor U7107 (N_7107,N_3190,N_2711);
and U7108 (N_7108,N_3182,N_3795);
nand U7109 (N_7109,N_3023,N_3873);
nand U7110 (N_7110,N_2873,N_3462);
nor U7111 (N_7111,N_2809,N_4445);
nand U7112 (N_7112,N_4899,N_4912);
and U7113 (N_7113,N_3035,N_3236);
or U7114 (N_7114,N_4695,N_3419);
nor U7115 (N_7115,N_4822,N_3037);
and U7116 (N_7116,N_4061,N_3586);
and U7117 (N_7117,N_4810,N_4188);
xnor U7118 (N_7118,N_4215,N_4435);
nand U7119 (N_7119,N_3825,N_2833);
and U7120 (N_7120,N_3312,N_3190);
nor U7121 (N_7121,N_2811,N_3419);
xnor U7122 (N_7122,N_2779,N_4586);
or U7123 (N_7123,N_3038,N_3053);
or U7124 (N_7124,N_4253,N_3896);
or U7125 (N_7125,N_3528,N_3251);
or U7126 (N_7126,N_4734,N_4396);
nor U7127 (N_7127,N_3311,N_2926);
or U7128 (N_7128,N_4952,N_2668);
and U7129 (N_7129,N_3180,N_2881);
or U7130 (N_7130,N_3560,N_2608);
or U7131 (N_7131,N_3543,N_4964);
nand U7132 (N_7132,N_2792,N_4948);
and U7133 (N_7133,N_3839,N_3939);
nor U7134 (N_7134,N_4898,N_2583);
and U7135 (N_7135,N_4522,N_3954);
and U7136 (N_7136,N_4349,N_3671);
nor U7137 (N_7137,N_3561,N_4975);
or U7138 (N_7138,N_4991,N_4913);
nand U7139 (N_7139,N_4335,N_2699);
nor U7140 (N_7140,N_4367,N_3853);
nor U7141 (N_7141,N_4950,N_3173);
xor U7142 (N_7142,N_3866,N_2851);
nor U7143 (N_7143,N_4260,N_4287);
nor U7144 (N_7144,N_4475,N_2530);
xnor U7145 (N_7145,N_4963,N_4419);
or U7146 (N_7146,N_4238,N_3445);
and U7147 (N_7147,N_2556,N_2670);
or U7148 (N_7148,N_3332,N_3018);
nor U7149 (N_7149,N_3614,N_3046);
nor U7150 (N_7150,N_3189,N_4797);
and U7151 (N_7151,N_3459,N_3426);
and U7152 (N_7152,N_4855,N_4440);
nor U7153 (N_7153,N_4545,N_3386);
nand U7154 (N_7154,N_2544,N_3099);
nand U7155 (N_7155,N_3196,N_4578);
nor U7156 (N_7156,N_3587,N_4027);
or U7157 (N_7157,N_2633,N_4690);
nand U7158 (N_7158,N_2577,N_2596);
nor U7159 (N_7159,N_3519,N_3813);
and U7160 (N_7160,N_3177,N_4133);
or U7161 (N_7161,N_4787,N_2812);
nor U7162 (N_7162,N_2576,N_4347);
nor U7163 (N_7163,N_2831,N_4806);
and U7164 (N_7164,N_3283,N_3373);
nand U7165 (N_7165,N_2834,N_4780);
or U7166 (N_7166,N_3653,N_2507);
nor U7167 (N_7167,N_2619,N_2524);
nor U7168 (N_7168,N_4347,N_2734);
nor U7169 (N_7169,N_3758,N_3294);
and U7170 (N_7170,N_2622,N_2706);
or U7171 (N_7171,N_3882,N_4932);
and U7172 (N_7172,N_4187,N_4515);
and U7173 (N_7173,N_4754,N_3049);
and U7174 (N_7174,N_4205,N_4963);
and U7175 (N_7175,N_3854,N_4154);
nor U7176 (N_7176,N_3930,N_4666);
and U7177 (N_7177,N_3060,N_2640);
or U7178 (N_7178,N_2810,N_4772);
or U7179 (N_7179,N_2601,N_4359);
nand U7180 (N_7180,N_2742,N_2781);
nor U7181 (N_7181,N_3559,N_3169);
and U7182 (N_7182,N_4624,N_2842);
or U7183 (N_7183,N_3371,N_3214);
nor U7184 (N_7184,N_4131,N_4094);
nand U7185 (N_7185,N_2839,N_4534);
or U7186 (N_7186,N_4913,N_3898);
nor U7187 (N_7187,N_3895,N_4805);
nor U7188 (N_7188,N_3343,N_4555);
or U7189 (N_7189,N_3153,N_3958);
xnor U7190 (N_7190,N_4046,N_3433);
or U7191 (N_7191,N_3654,N_4487);
and U7192 (N_7192,N_3893,N_4133);
nor U7193 (N_7193,N_4451,N_4275);
nor U7194 (N_7194,N_4277,N_3495);
nand U7195 (N_7195,N_3620,N_3711);
nor U7196 (N_7196,N_3048,N_4251);
nor U7197 (N_7197,N_3290,N_3015);
and U7198 (N_7198,N_3886,N_4966);
and U7199 (N_7199,N_3933,N_3254);
nor U7200 (N_7200,N_4435,N_2669);
xor U7201 (N_7201,N_4778,N_3789);
nor U7202 (N_7202,N_4943,N_3072);
nor U7203 (N_7203,N_3247,N_4395);
nor U7204 (N_7204,N_3413,N_3748);
or U7205 (N_7205,N_3539,N_4984);
nand U7206 (N_7206,N_3153,N_4419);
nor U7207 (N_7207,N_3946,N_2755);
and U7208 (N_7208,N_3058,N_4328);
nor U7209 (N_7209,N_3520,N_2754);
or U7210 (N_7210,N_4807,N_4597);
or U7211 (N_7211,N_2740,N_4357);
or U7212 (N_7212,N_4782,N_2721);
and U7213 (N_7213,N_3871,N_3217);
nor U7214 (N_7214,N_4805,N_3359);
nor U7215 (N_7215,N_3840,N_4318);
and U7216 (N_7216,N_3089,N_4727);
and U7217 (N_7217,N_4798,N_3335);
nand U7218 (N_7218,N_4379,N_3555);
nor U7219 (N_7219,N_2640,N_4853);
and U7220 (N_7220,N_4636,N_4621);
nor U7221 (N_7221,N_4342,N_2686);
nor U7222 (N_7222,N_2999,N_3601);
or U7223 (N_7223,N_3531,N_2640);
nand U7224 (N_7224,N_4837,N_4171);
nand U7225 (N_7225,N_3726,N_3170);
or U7226 (N_7226,N_4778,N_2512);
and U7227 (N_7227,N_2768,N_4575);
nor U7228 (N_7228,N_3347,N_2728);
and U7229 (N_7229,N_4513,N_4038);
nor U7230 (N_7230,N_2621,N_4639);
or U7231 (N_7231,N_3249,N_3143);
nand U7232 (N_7232,N_3435,N_3734);
or U7233 (N_7233,N_3349,N_3690);
nor U7234 (N_7234,N_3355,N_3805);
or U7235 (N_7235,N_3919,N_3713);
nor U7236 (N_7236,N_4821,N_2950);
nor U7237 (N_7237,N_3249,N_2751);
nor U7238 (N_7238,N_4887,N_2687);
nand U7239 (N_7239,N_4352,N_3885);
and U7240 (N_7240,N_3407,N_4993);
and U7241 (N_7241,N_2970,N_2525);
nand U7242 (N_7242,N_4974,N_3539);
nor U7243 (N_7243,N_3127,N_3335);
and U7244 (N_7244,N_3169,N_3866);
or U7245 (N_7245,N_4787,N_4449);
or U7246 (N_7246,N_4128,N_3184);
nor U7247 (N_7247,N_2516,N_4726);
and U7248 (N_7248,N_3365,N_4957);
nand U7249 (N_7249,N_3512,N_4797);
and U7250 (N_7250,N_4494,N_4407);
or U7251 (N_7251,N_4760,N_2702);
and U7252 (N_7252,N_2743,N_2624);
nor U7253 (N_7253,N_4001,N_4675);
or U7254 (N_7254,N_3970,N_3613);
and U7255 (N_7255,N_3645,N_3983);
or U7256 (N_7256,N_3985,N_3755);
and U7257 (N_7257,N_3606,N_2544);
and U7258 (N_7258,N_4410,N_3532);
xor U7259 (N_7259,N_4213,N_3773);
nand U7260 (N_7260,N_3000,N_3214);
and U7261 (N_7261,N_4665,N_2729);
and U7262 (N_7262,N_4392,N_4591);
and U7263 (N_7263,N_2928,N_3950);
or U7264 (N_7264,N_3953,N_3961);
or U7265 (N_7265,N_3573,N_3755);
or U7266 (N_7266,N_4317,N_3460);
nand U7267 (N_7267,N_3277,N_2699);
nor U7268 (N_7268,N_4258,N_4854);
or U7269 (N_7269,N_4529,N_2589);
nand U7270 (N_7270,N_3957,N_4914);
nor U7271 (N_7271,N_3182,N_3972);
and U7272 (N_7272,N_2649,N_3883);
nand U7273 (N_7273,N_3095,N_3646);
nor U7274 (N_7274,N_4972,N_3315);
and U7275 (N_7275,N_4140,N_4385);
nand U7276 (N_7276,N_4745,N_4997);
nand U7277 (N_7277,N_4522,N_4687);
nor U7278 (N_7278,N_3838,N_3410);
nand U7279 (N_7279,N_2960,N_3722);
nand U7280 (N_7280,N_3847,N_3718);
and U7281 (N_7281,N_2577,N_4599);
nor U7282 (N_7282,N_4841,N_4868);
or U7283 (N_7283,N_3758,N_2852);
and U7284 (N_7284,N_3536,N_4598);
xnor U7285 (N_7285,N_3889,N_4744);
nor U7286 (N_7286,N_3364,N_3844);
nor U7287 (N_7287,N_2754,N_3253);
nor U7288 (N_7288,N_3111,N_3126);
nor U7289 (N_7289,N_4830,N_2794);
nand U7290 (N_7290,N_4225,N_3857);
and U7291 (N_7291,N_4583,N_4431);
and U7292 (N_7292,N_3925,N_3576);
and U7293 (N_7293,N_2625,N_2522);
or U7294 (N_7294,N_2973,N_3289);
or U7295 (N_7295,N_4206,N_4924);
or U7296 (N_7296,N_2841,N_2545);
or U7297 (N_7297,N_4556,N_4016);
and U7298 (N_7298,N_3608,N_4546);
nor U7299 (N_7299,N_4045,N_4159);
nor U7300 (N_7300,N_3167,N_3348);
and U7301 (N_7301,N_2727,N_3213);
or U7302 (N_7302,N_4463,N_2513);
or U7303 (N_7303,N_3023,N_4231);
nor U7304 (N_7304,N_4709,N_3461);
nand U7305 (N_7305,N_3273,N_3670);
xor U7306 (N_7306,N_4025,N_4072);
and U7307 (N_7307,N_4716,N_4707);
nand U7308 (N_7308,N_4846,N_3007);
and U7309 (N_7309,N_4106,N_2843);
nand U7310 (N_7310,N_4050,N_3924);
nor U7311 (N_7311,N_4632,N_3562);
nor U7312 (N_7312,N_3106,N_4864);
and U7313 (N_7313,N_2841,N_3038);
nand U7314 (N_7314,N_3126,N_3808);
nand U7315 (N_7315,N_2817,N_3687);
nor U7316 (N_7316,N_2633,N_2588);
nand U7317 (N_7317,N_4935,N_3813);
nand U7318 (N_7318,N_3267,N_4137);
nor U7319 (N_7319,N_4122,N_2757);
or U7320 (N_7320,N_3762,N_2927);
xor U7321 (N_7321,N_3738,N_4528);
or U7322 (N_7322,N_4513,N_4250);
and U7323 (N_7323,N_3371,N_4587);
nand U7324 (N_7324,N_3870,N_4566);
nor U7325 (N_7325,N_3751,N_3739);
nor U7326 (N_7326,N_3075,N_2871);
nand U7327 (N_7327,N_4959,N_4771);
nor U7328 (N_7328,N_4984,N_4027);
nor U7329 (N_7329,N_3967,N_4124);
or U7330 (N_7330,N_4105,N_4167);
nor U7331 (N_7331,N_3456,N_4383);
and U7332 (N_7332,N_4786,N_4523);
nand U7333 (N_7333,N_2933,N_4739);
nor U7334 (N_7334,N_3009,N_4903);
nor U7335 (N_7335,N_2853,N_3135);
nor U7336 (N_7336,N_3360,N_4754);
nand U7337 (N_7337,N_4853,N_3638);
nand U7338 (N_7338,N_4002,N_4930);
or U7339 (N_7339,N_2893,N_4201);
or U7340 (N_7340,N_4947,N_4475);
nand U7341 (N_7341,N_4520,N_3849);
nand U7342 (N_7342,N_3644,N_4309);
nand U7343 (N_7343,N_4368,N_4599);
nand U7344 (N_7344,N_3090,N_4513);
nor U7345 (N_7345,N_4478,N_3196);
nor U7346 (N_7346,N_2765,N_3799);
and U7347 (N_7347,N_4226,N_4828);
xor U7348 (N_7348,N_3520,N_3525);
nor U7349 (N_7349,N_2782,N_4244);
nor U7350 (N_7350,N_3353,N_3982);
nor U7351 (N_7351,N_3508,N_2636);
nand U7352 (N_7352,N_2521,N_2662);
and U7353 (N_7353,N_3641,N_2918);
and U7354 (N_7354,N_3144,N_4306);
nor U7355 (N_7355,N_3770,N_4611);
nand U7356 (N_7356,N_3550,N_4645);
or U7357 (N_7357,N_3993,N_3074);
nand U7358 (N_7358,N_3574,N_2751);
and U7359 (N_7359,N_2770,N_4586);
or U7360 (N_7360,N_4965,N_4458);
nor U7361 (N_7361,N_4248,N_3829);
or U7362 (N_7362,N_3381,N_3168);
or U7363 (N_7363,N_4715,N_3800);
or U7364 (N_7364,N_4699,N_3471);
and U7365 (N_7365,N_2543,N_2566);
and U7366 (N_7366,N_4960,N_3182);
nand U7367 (N_7367,N_3505,N_4285);
nand U7368 (N_7368,N_4267,N_2931);
or U7369 (N_7369,N_4042,N_3006);
nor U7370 (N_7370,N_4858,N_3758);
or U7371 (N_7371,N_2870,N_4898);
and U7372 (N_7372,N_3699,N_3810);
nor U7373 (N_7373,N_2708,N_2539);
nor U7374 (N_7374,N_4857,N_3578);
or U7375 (N_7375,N_3866,N_3681);
and U7376 (N_7376,N_3424,N_4091);
nor U7377 (N_7377,N_4903,N_3417);
or U7378 (N_7378,N_3144,N_2691);
and U7379 (N_7379,N_3250,N_4159);
and U7380 (N_7380,N_2534,N_4292);
or U7381 (N_7381,N_3800,N_4479);
and U7382 (N_7382,N_4669,N_4907);
and U7383 (N_7383,N_3139,N_3922);
and U7384 (N_7384,N_3179,N_3443);
and U7385 (N_7385,N_3867,N_4319);
nand U7386 (N_7386,N_3758,N_4724);
nor U7387 (N_7387,N_4902,N_4164);
nor U7388 (N_7388,N_4430,N_2783);
nor U7389 (N_7389,N_4381,N_3357);
nor U7390 (N_7390,N_2751,N_4448);
and U7391 (N_7391,N_4110,N_3426);
or U7392 (N_7392,N_3958,N_2823);
and U7393 (N_7393,N_4829,N_4217);
and U7394 (N_7394,N_4398,N_2957);
nor U7395 (N_7395,N_4224,N_2807);
nand U7396 (N_7396,N_3962,N_3887);
or U7397 (N_7397,N_3965,N_2541);
nand U7398 (N_7398,N_2910,N_3168);
or U7399 (N_7399,N_3341,N_3101);
and U7400 (N_7400,N_2605,N_3320);
and U7401 (N_7401,N_3042,N_3399);
or U7402 (N_7402,N_3321,N_3737);
nand U7403 (N_7403,N_2513,N_4571);
nor U7404 (N_7404,N_2528,N_3783);
xor U7405 (N_7405,N_4064,N_4729);
xnor U7406 (N_7406,N_4692,N_4216);
or U7407 (N_7407,N_3123,N_4583);
or U7408 (N_7408,N_2638,N_3035);
and U7409 (N_7409,N_4643,N_3183);
and U7410 (N_7410,N_3076,N_4050);
and U7411 (N_7411,N_4263,N_3217);
and U7412 (N_7412,N_3396,N_3824);
nand U7413 (N_7413,N_2834,N_2745);
or U7414 (N_7414,N_4770,N_3896);
nor U7415 (N_7415,N_4090,N_4956);
xor U7416 (N_7416,N_4728,N_2587);
and U7417 (N_7417,N_4294,N_2600);
nor U7418 (N_7418,N_3405,N_3062);
or U7419 (N_7419,N_2730,N_4830);
nand U7420 (N_7420,N_3721,N_3765);
nand U7421 (N_7421,N_2764,N_4837);
nand U7422 (N_7422,N_4830,N_3711);
or U7423 (N_7423,N_3298,N_3523);
nand U7424 (N_7424,N_3530,N_3636);
nand U7425 (N_7425,N_3895,N_4531);
nor U7426 (N_7426,N_3092,N_2967);
or U7427 (N_7427,N_3856,N_2637);
nor U7428 (N_7428,N_2959,N_3788);
and U7429 (N_7429,N_3752,N_4190);
and U7430 (N_7430,N_3023,N_4860);
nor U7431 (N_7431,N_3494,N_4149);
or U7432 (N_7432,N_2689,N_3711);
or U7433 (N_7433,N_4945,N_4120);
or U7434 (N_7434,N_3321,N_4689);
nand U7435 (N_7435,N_4447,N_4399);
or U7436 (N_7436,N_4781,N_4217);
or U7437 (N_7437,N_2515,N_4114);
nand U7438 (N_7438,N_2917,N_4410);
or U7439 (N_7439,N_2947,N_2587);
nor U7440 (N_7440,N_3909,N_4559);
and U7441 (N_7441,N_4237,N_3689);
nand U7442 (N_7442,N_3121,N_3562);
and U7443 (N_7443,N_4479,N_2924);
or U7444 (N_7444,N_2520,N_2807);
and U7445 (N_7445,N_4929,N_4518);
nand U7446 (N_7446,N_3833,N_3945);
or U7447 (N_7447,N_2838,N_2532);
or U7448 (N_7448,N_3469,N_4811);
and U7449 (N_7449,N_3096,N_3003);
and U7450 (N_7450,N_3580,N_4653);
nand U7451 (N_7451,N_2666,N_3533);
and U7452 (N_7452,N_2926,N_3168);
nor U7453 (N_7453,N_4159,N_2828);
or U7454 (N_7454,N_3579,N_4738);
nor U7455 (N_7455,N_3316,N_4388);
nor U7456 (N_7456,N_4243,N_3116);
or U7457 (N_7457,N_2670,N_3059);
nor U7458 (N_7458,N_2818,N_3427);
or U7459 (N_7459,N_4208,N_3635);
or U7460 (N_7460,N_2813,N_3021);
and U7461 (N_7461,N_4300,N_4894);
nand U7462 (N_7462,N_4570,N_4210);
and U7463 (N_7463,N_3273,N_3052);
and U7464 (N_7464,N_3969,N_4827);
and U7465 (N_7465,N_3683,N_3564);
nand U7466 (N_7466,N_4470,N_2928);
nand U7467 (N_7467,N_3841,N_4991);
nor U7468 (N_7468,N_3583,N_3398);
nand U7469 (N_7469,N_3967,N_3350);
nand U7470 (N_7470,N_3656,N_3688);
nor U7471 (N_7471,N_2599,N_2610);
or U7472 (N_7472,N_4177,N_3933);
or U7473 (N_7473,N_3664,N_3150);
or U7474 (N_7474,N_4138,N_4948);
nand U7475 (N_7475,N_3349,N_3830);
nand U7476 (N_7476,N_4070,N_3561);
and U7477 (N_7477,N_3001,N_4850);
or U7478 (N_7478,N_4967,N_3209);
or U7479 (N_7479,N_4809,N_3473);
or U7480 (N_7480,N_4358,N_2519);
and U7481 (N_7481,N_4287,N_2506);
and U7482 (N_7482,N_3075,N_3753);
and U7483 (N_7483,N_2583,N_4341);
nand U7484 (N_7484,N_2509,N_4182);
nor U7485 (N_7485,N_3126,N_3412);
and U7486 (N_7486,N_3796,N_4230);
or U7487 (N_7487,N_4561,N_4633);
nand U7488 (N_7488,N_3287,N_3261);
and U7489 (N_7489,N_2921,N_3177);
and U7490 (N_7490,N_3533,N_3938);
and U7491 (N_7491,N_4525,N_2888);
or U7492 (N_7492,N_4169,N_3999);
and U7493 (N_7493,N_2649,N_4477);
nand U7494 (N_7494,N_4560,N_4312);
nor U7495 (N_7495,N_2662,N_3625);
or U7496 (N_7496,N_3949,N_2870);
and U7497 (N_7497,N_2555,N_3629);
nand U7498 (N_7498,N_2650,N_3012);
nor U7499 (N_7499,N_3395,N_2817);
or U7500 (N_7500,N_6209,N_5303);
nand U7501 (N_7501,N_6720,N_7260);
or U7502 (N_7502,N_5321,N_7092);
or U7503 (N_7503,N_6300,N_6432);
nand U7504 (N_7504,N_6415,N_6368);
nand U7505 (N_7505,N_6750,N_6408);
nand U7506 (N_7506,N_5731,N_5344);
or U7507 (N_7507,N_6542,N_5103);
or U7508 (N_7508,N_7202,N_5665);
or U7509 (N_7509,N_6439,N_5526);
nor U7510 (N_7510,N_6983,N_6955);
and U7511 (N_7511,N_5500,N_6605);
or U7512 (N_7512,N_5358,N_5166);
nand U7513 (N_7513,N_6562,N_6360);
nand U7514 (N_7514,N_5946,N_6261);
or U7515 (N_7515,N_5318,N_7127);
and U7516 (N_7516,N_5858,N_5035);
nor U7517 (N_7517,N_5814,N_7125);
or U7518 (N_7518,N_6323,N_6664);
and U7519 (N_7519,N_6317,N_7041);
or U7520 (N_7520,N_6397,N_7131);
or U7521 (N_7521,N_5393,N_7227);
nor U7522 (N_7522,N_5610,N_5425);
nand U7523 (N_7523,N_5597,N_6172);
and U7524 (N_7524,N_7012,N_6784);
and U7525 (N_7525,N_6221,N_7451);
nor U7526 (N_7526,N_7339,N_5109);
and U7527 (N_7527,N_7289,N_5983);
or U7528 (N_7528,N_7374,N_7393);
nor U7529 (N_7529,N_5199,N_7257);
or U7530 (N_7530,N_5911,N_7252);
and U7531 (N_7531,N_7259,N_5867);
nand U7532 (N_7532,N_7347,N_6019);
and U7533 (N_7533,N_5095,N_5666);
nor U7534 (N_7534,N_7377,N_6100);
and U7535 (N_7535,N_5609,N_5599);
nand U7536 (N_7536,N_7460,N_6339);
or U7537 (N_7537,N_7258,N_5114);
and U7538 (N_7538,N_5053,N_6251);
nand U7539 (N_7539,N_5022,N_7022);
nand U7540 (N_7540,N_7416,N_7140);
or U7541 (N_7541,N_6770,N_6066);
and U7542 (N_7542,N_6158,N_7098);
nand U7543 (N_7543,N_6441,N_6508);
nand U7544 (N_7544,N_7061,N_7219);
nor U7545 (N_7545,N_6632,N_6090);
xnor U7546 (N_7546,N_6450,N_6622);
nor U7547 (N_7547,N_7471,N_7344);
nor U7548 (N_7548,N_6776,N_6695);
or U7549 (N_7549,N_5144,N_6222);
nor U7550 (N_7550,N_6073,N_5213);
or U7551 (N_7551,N_7062,N_6585);
nor U7552 (N_7552,N_5210,N_5941);
and U7553 (N_7553,N_6617,N_6858);
and U7554 (N_7554,N_6686,N_7182);
nor U7555 (N_7555,N_5119,N_5269);
nand U7556 (N_7556,N_6016,N_7267);
nor U7557 (N_7557,N_6823,N_5904);
and U7558 (N_7558,N_6520,N_6410);
and U7559 (N_7559,N_6655,N_6097);
or U7560 (N_7560,N_7063,N_6546);
nor U7561 (N_7561,N_5945,N_6581);
or U7562 (N_7562,N_7058,N_6281);
or U7563 (N_7563,N_5080,N_7086);
or U7564 (N_7564,N_5395,N_5973);
and U7565 (N_7565,N_6236,N_7466);
and U7566 (N_7566,N_6773,N_5376);
or U7567 (N_7567,N_6496,N_6824);
nand U7568 (N_7568,N_5850,N_5219);
nand U7569 (N_7569,N_5214,N_6952);
or U7570 (N_7570,N_5564,N_5504);
and U7571 (N_7571,N_5137,N_7019);
nand U7572 (N_7572,N_6467,N_5441);
or U7573 (N_7573,N_7372,N_6991);
and U7574 (N_7574,N_5200,N_5203);
and U7575 (N_7575,N_6126,N_6110);
nor U7576 (N_7576,N_7053,N_6525);
nand U7577 (N_7577,N_5511,N_6091);
nand U7578 (N_7578,N_6836,N_5592);
nand U7579 (N_7579,N_5872,N_6917);
and U7580 (N_7580,N_5679,N_5031);
and U7581 (N_7581,N_5548,N_6280);
nand U7582 (N_7582,N_7494,N_7121);
or U7583 (N_7583,N_5189,N_6088);
nand U7584 (N_7584,N_5366,N_6111);
xor U7585 (N_7585,N_6700,N_7176);
nor U7586 (N_7586,N_7271,N_5832);
xnor U7587 (N_7587,N_6697,N_5228);
nor U7588 (N_7588,N_5322,N_6850);
and U7589 (N_7589,N_6744,N_6143);
nor U7590 (N_7590,N_6215,N_6906);
nor U7591 (N_7591,N_7417,N_6396);
or U7592 (N_7592,N_5554,N_5929);
or U7593 (N_7593,N_7395,N_5796);
or U7594 (N_7594,N_6780,N_6514);
nand U7595 (N_7595,N_6272,N_6404);
and U7596 (N_7596,N_5662,N_6925);
nand U7597 (N_7597,N_5217,N_5400);
or U7598 (N_7598,N_6354,N_6376);
nand U7599 (N_7599,N_7065,N_6682);
nor U7600 (N_7600,N_5543,N_5473);
nor U7601 (N_7601,N_5834,N_6528);
and U7602 (N_7602,N_6247,N_5996);
and U7603 (N_7603,N_7305,N_6296);
nor U7604 (N_7604,N_6896,N_5444);
xnor U7605 (N_7605,N_7264,N_7123);
nor U7606 (N_7606,N_7263,N_6041);
and U7607 (N_7607,N_6549,N_5990);
and U7608 (N_7608,N_6973,N_6327);
or U7609 (N_7609,N_7486,N_5994);
nand U7610 (N_7610,N_5813,N_6616);
or U7611 (N_7611,N_6321,N_5222);
and U7612 (N_7612,N_6954,N_6839);
nand U7613 (N_7613,N_5306,N_5681);
nand U7614 (N_7614,N_5244,N_5678);
or U7615 (N_7615,N_5497,N_7438);
nor U7616 (N_7616,N_5073,N_5353);
or U7617 (N_7617,N_6861,N_6948);
nand U7618 (N_7618,N_5803,N_6085);
or U7619 (N_7619,N_5374,N_5055);
nor U7620 (N_7620,N_6976,N_6208);
and U7621 (N_7621,N_5593,N_6586);
or U7622 (N_7622,N_6003,N_5894);
nand U7623 (N_7623,N_5237,N_6014);
nor U7624 (N_7624,N_6036,N_5216);
and U7625 (N_7625,N_5236,N_7241);
nand U7626 (N_7626,N_5557,N_6465);
and U7627 (N_7627,N_7101,N_6464);
and U7628 (N_7628,N_6289,N_5633);
nand U7629 (N_7629,N_6042,N_6064);
and U7630 (N_7630,N_6060,N_5628);
nand U7631 (N_7631,N_5312,N_5041);
nor U7632 (N_7632,N_6517,N_6507);
nand U7633 (N_7633,N_5392,N_5367);
and U7634 (N_7634,N_5205,N_5157);
and U7635 (N_7635,N_5383,N_5350);
nor U7636 (N_7636,N_6595,N_7413);
nor U7637 (N_7637,N_5925,N_6388);
and U7638 (N_7638,N_5962,N_6257);
xnor U7639 (N_7639,N_5487,N_6862);
and U7640 (N_7640,N_5076,N_7371);
nor U7641 (N_7641,N_6648,N_6718);
and U7642 (N_7642,N_5057,N_7407);
and U7643 (N_7643,N_5278,N_7095);
or U7644 (N_7644,N_6455,N_7013);
and U7645 (N_7645,N_6270,N_5719);
nand U7646 (N_7646,N_5579,N_6480);
or U7647 (N_7647,N_6913,N_5506);
nand U7648 (N_7648,N_5470,N_6214);
and U7649 (N_7649,N_6969,N_5617);
nand U7650 (N_7650,N_6030,N_5281);
or U7651 (N_7651,N_5958,N_6055);
or U7652 (N_7652,N_7448,N_6637);
or U7653 (N_7653,N_6411,N_7387);
and U7654 (N_7654,N_6279,N_7352);
and U7655 (N_7655,N_5775,N_6890);
and U7656 (N_7656,N_5711,N_5771);
nand U7657 (N_7657,N_6371,N_7007);
and U7658 (N_7658,N_6628,N_5355);
and U7659 (N_7659,N_5865,N_6844);
nand U7660 (N_7660,N_7298,N_6361);
or U7661 (N_7661,N_7214,N_6384);
nor U7662 (N_7662,N_5536,N_5721);
nor U7663 (N_7663,N_6136,N_7453);
or U7664 (N_7664,N_5625,N_7401);
or U7665 (N_7665,N_5459,N_6802);
or U7666 (N_7666,N_5739,N_6867);
nand U7667 (N_7667,N_5408,N_6774);
nand U7668 (N_7668,N_6422,N_6212);
and U7669 (N_7669,N_6592,N_7035);
nand U7670 (N_7670,N_6988,N_7358);
or U7671 (N_7671,N_6963,N_5452);
nor U7672 (N_7672,N_6102,N_6031);
or U7673 (N_7673,N_6054,N_6125);
and U7674 (N_7674,N_5466,N_5952);
nor U7675 (N_7675,N_7415,N_6928);
and U7676 (N_7676,N_6083,N_5156);
nor U7677 (N_7677,N_5177,N_5265);
or U7678 (N_7678,N_5328,N_7248);
xor U7679 (N_7679,N_7126,N_5718);
and U7680 (N_7680,N_6240,N_6606);
or U7681 (N_7681,N_5063,N_5453);
nand U7682 (N_7682,N_7034,N_6044);
or U7683 (N_7683,N_6936,N_6334);
nor U7684 (N_7684,N_5496,N_7188);
and U7685 (N_7685,N_6337,N_6702);
nor U7686 (N_7686,N_7002,N_5810);
nor U7687 (N_7687,N_5493,N_5825);
nand U7688 (N_7688,N_6128,N_7112);
and U7689 (N_7689,N_5180,N_6828);
or U7690 (N_7690,N_5622,N_7097);
and U7691 (N_7691,N_5720,N_6551);
nor U7692 (N_7692,N_6650,N_6488);
nand U7693 (N_7693,N_7194,N_5456);
nand U7694 (N_7694,N_6293,N_5451);
nand U7695 (N_7695,N_7164,N_5113);
nand U7696 (N_7696,N_6949,N_5785);
nand U7697 (N_7697,N_5017,N_5623);
xor U7698 (N_7698,N_6196,N_6149);
nand U7699 (N_7699,N_5507,N_6608);
or U7700 (N_7700,N_5188,N_6275);
nand U7701 (N_7701,N_6736,N_6071);
and U7702 (N_7702,N_6957,N_5870);
nand U7703 (N_7703,N_6856,N_7147);
nand U7704 (N_7704,N_6364,N_6587);
nor U7705 (N_7705,N_6444,N_5435);
nor U7706 (N_7706,N_6959,N_7273);
nor U7707 (N_7707,N_6479,N_5152);
nand U7708 (N_7708,N_5651,N_7403);
nor U7709 (N_7709,N_6059,N_7433);
nor U7710 (N_7710,N_5852,N_5263);
nand U7711 (N_7711,N_6712,N_5676);
and U7712 (N_7712,N_6918,N_6927);
nor U7713 (N_7713,N_5656,N_5715);
and U7714 (N_7714,N_6375,N_7026);
nand U7715 (N_7715,N_6937,N_5737);
nor U7716 (N_7716,N_5970,N_5067);
nand U7717 (N_7717,N_7286,N_5296);
and U7718 (N_7718,N_5158,N_6502);
nand U7719 (N_7719,N_7011,N_5066);
nand U7720 (N_7720,N_6420,N_7354);
nor U7721 (N_7721,N_7047,N_5967);
or U7722 (N_7722,N_5752,N_5999);
xor U7723 (N_7723,N_5283,N_7447);
or U7724 (N_7724,N_5964,N_5495);
nand U7725 (N_7725,N_5551,N_6755);
xnor U7726 (N_7726,N_6521,N_5713);
and U7727 (N_7727,N_5133,N_5956);
xor U7728 (N_7728,N_6344,N_7443);
nand U7729 (N_7729,N_5123,N_5920);
nor U7730 (N_7730,N_6716,N_7238);
nand U7731 (N_7731,N_6678,N_6288);
nor U7732 (N_7732,N_6714,N_5880);
and U7733 (N_7733,N_7315,N_6006);
and U7734 (N_7734,N_7322,N_7021);
and U7735 (N_7735,N_6241,N_6843);
nand U7736 (N_7736,N_7069,N_6934);
xnor U7737 (N_7737,N_5172,N_6685);
nor U7738 (N_7738,N_7146,N_5347);
nand U7739 (N_7739,N_5330,N_5749);
or U7740 (N_7740,N_6942,N_7275);
nor U7741 (N_7741,N_6846,N_6571);
xor U7742 (N_7742,N_5710,N_6096);
xnor U7743 (N_7743,N_5699,N_5257);
or U7744 (N_7744,N_5437,N_5221);
nor U7745 (N_7745,N_7262,N_5953);
nand U7746 (N_7746,N_5815,N_7349);
nand U7747 (N_7747,N_5225,N_6476);
and U7748 (N_7748,N_7308,N_5000);
nand U7749 (N_7749,N_6421,N_6228);
or U7750 (N_7750,N_6558,N_7279);
nand U7751 (N_7751,N_6638,N_7190);
and U7752 (N_7752,N_5051,N_5805);
nand U7753 (N_7753,N_5782,N_5369);
and U7754 (N_7754,N_5307,N_6553);
and U7755 (N_7755,N_7096,N_6458);
nor U7756 (N_7756,N_5838,N_5837);
nand U7757 (N_7757,N_7199,N_5800);
nor U7758 (N_7758,N_5842,N_7060);
and U7759 (N_7759,N_6137,N_5434);
nor U7760 (N_7760,N_7309,N_6944);
xnor U7761 (N_7761,N_5270,N_5256);
and U7762 (N_7762,N_6821,N_6238);
and U7763 (N_7763,N_6310,N_6000);
or U7764 (N_7764,N_6911,N_7091);
and U7765 (N_7765,N_6472,N_5424);
nand U7766 (N_7766,N_5845,N_7225);
nor U7767 (N_7767,N_6218,N_5044);
nand U7768 (N_7768,N_7468,N_5988);
and U7769 (N_7769,N_7142,N_5012);
or U7770 (N_7770,N_6207,N_5407);
nor U7771 (N_7771,N_6416,N_6295);
nand U7772 (N_7772,N_5575,N_5345);
nand U7773 (N_7773,N_6095,N_6387);
nor U7774 (N_7774,N_5758,N_5950);
and U7775 (N_7775,N_5847,N_6227);
nor U7776 (N_7776,N_6484,N_6004);
or U7777 (N_7777,N_5913,N_7470);
or U7778 (N_7778,N_6081,N_7191);
or U7779 (N_7779,N_5528,N_5280);
or U7780 (N_7780,N_5140,N_6604);
or U7781 (N_7781,N_5115,N_5914);
or U7782 (N_7782,N_5129,N_6367);
or U7783 (N_7783,N_7467,N_7427);
or U7784 (N_7784,N_5045,N_5191);
or U7785 (N_7785,N_7392,N_5039);
nor U7786 (N_7786,N_6121,N_5589);
and U7787 (N_7787,N_6267,N_6038);
nor U7788 (N_7788,N_6056,N_7281);
nor U7789 (N_7789,N_6947,N_6769);
nand U7790 (N_7790,N_5846,N_6181);
nor U7791 (N_7791,N_5272,N_5241);
or U7792 (N_7792,N_6008,N_5671);
or U7793 (N_7793,N_6148,N_6303);
and U7794 (N_7794,N_5294,N_6366);
or U7795 (N_7795,N_6609,N_7244);
nand U7796 (N_7796,N_5448,N_6061);
nor U7797 (N_7797,N_7228,N_6298);
or U7798 (N_7798,N_6199,N_6242);
nor U7799 (N_7799,N_7333,N_7155);
and U7800 (N_7800,N_5398,N_5650);
or U7801 (N_7801,N_5293,N_6735);
nor U7802 (N_7802,N_7030,N_6533);
or U7803 (N_7803,N_5429,N_7066);
nor U7804 (N_7804,N_6803,N_7111);
nor U7805 (N_7805,N_6929,N_5149);
or U7806 (N_7806,N_6576,N_5480);
nor U7807 (N_7807,N_6989,N_5433);
or U7808 (N_7808,N_6167,N_5816);
nand U7809 (N_7809,N_6899,N_5636);
nand U7810 (N_7810,N_5975,N_6249);
nand U7811 (N_7811,N_5336,N_6941);
nor U7812 (N_7812,N_5895,N_6547);
or U7813 (N_7813,N_7362,N_6347);
nand U7814 (N_7814,N_6194,N_6400);
and U7815 (N_7815,N_5488,N_5744);
and U7816 (N_7816,N_5323,N_6732);
nand U7817 (N_7817,N_6322,N_7221);
or U7818 (N_7818,N_5583,N_5447);
or U7819 (N_7819,N_7226,N_5394);
nand U7820 (N_7820,N_6406,N_7074);
and U7821 (N_7821,N_6179,N_6490);
or U7822 (N_7822,N_6010,N_7269);
and U7823 (N_7823,N_5181,N_5326);
nor U7824 (N_7824,N_5741,N_6916);
and U7825 (N_7825,N_5742,N_6103);
nand U7826 (N_7826,N_7493,N_7004);
and U7827 (N_7827,N_5049,N_7028);
nand U7828 (N_7828,N_7280,N_5750);
and U7829 (N_7829,N_5624,N_6244);
nor U7830 (N_7830,N_6140,N_5827);
nor U7831 (N_7831,N_5889,N_5851);
and U7832 (N_7832,N_6738,N_7446);
or U7833 (N_7833,N_5111,N_7032);
nor U7834 (N_7834,N_5260,N_6013);
and U7835 (N_7835,N_6186,N_6779);
xnor U7836 (N_7836,N_6094,N_6037);
nor U7837 (N_7837,N_5254,N_5783);
or U7838 (N_7838,N_7180,N_6523);
nor U7839 (N_7839,N_6302,N_7306);
or U7840 (N_7840,N_7031,N_6990);
nand U7841 (N_7841,N_7463,N_6499);
and U7842 (N_7842,N_5716,N_5768);
and U7843 (N_7843,N_5584,N_5933);
nor U7844 (N_7844,N_5841,N_6975);
or U7845 (N_7845,N_6982,N_6707);
nand U7846 (N_7846,N_6751,N_5462);
nand U7847 (N_7847,N_5627,N_5764);
or U7848 (N_7848,N_6104,N_5036);
or U7849 (N_7849,N_6579,N_6264);
nand U7850 (N_7850,N_6427,N_6793);
and U7851 (N_7851,N_6224,N_6837);
and U7852 (N_7852,N_5823,N_5023);
nor U7853 (N_7853,N_6342,N_5763);
nor U7854 (N_7854,N_5559,N_5364);
nand U7855 (N_7855,N_5161,N_6356);
and U7856 (N_7856,N_7179,N_5591);
and U7857 (N_7857,N_5324,N_6204);
or U7858 (N_7858,N_6825,N_6854);
nand U7859 (N_7859,N_5982,N_6092);
nor U7860 (N_7860,N_5082,N_7181);
or U7861 (N_7861,N_7391,N_7476);
or U7862 (N_7862,N_7234,N_5160);
nor U7863 (N_7863,N_5995,N_6184);
and U7864 (N_7864,N_6559,N_5380);
nor U7865 (N_7865,N_5010,N_6745);
or U7866 (N_7866,N_6883,N_5690);
or U7867 (N_7867,N_7249,N_6058);
nand U7868 (N_7868,N_6902,N_5853);
nand U7869 (N_7869,N_5302,N_6070);
and U7870 (N_7870,N_6552,N_5682);
nand U7871 (N_7871,N_7108,N_5709);
nor U7872 (N_7872,N_6974,N_5352);
and U7873 (N_7873,N_6329,N_5342);
and U7874 (N_7874,N_7014,N_6806);
nand U7875 (N_7875,N_6357,N_6150);
nor U7876 (N_7876,N_7198,N_7473);
or U7877 (N_7877,N_6398,N_6893);
or U7878 (N_7878,N_5648,N_5885);
nor U7879 (N_7879,N_5375,N_5091);
and U7880 (N_7880,N_6381,N_7268);
or U7881 (N_7881,N_5518,N_5164);
nor U7882 (N_7882,N_6333,N_7441);
nand U7883 (N_7883,N_6067,N_5926);
or U7884 (N_7884,N_5391,N_5949);
nor U7885 (N_7885,N_6938,N_6946);
and U7886 (N_7886,N_5547,N_7410);
or U7887 (N_7887,N_6764,N_6574);
nand U7888 (N_7888,N_6739,N_7492);
or U7889 (N_7889,N_5986,N_5505);
nor U7890 (N_7890,N_5381,N_6453);
nor U7891 (N_7891,N_7003,N_6461);
and U7892 (N_7892,N_7076,N_6516);
nand U7893 (N_7893,N_5315,N_7288);
nand U7894 (N_7894,N_5420,N_5596);
nor U7895 (N_7895,N_7364,N_6414);
or U7896 (N_7896,N_5708,N_5879);
nor U7897 (N_7897,N_5276,N_5234);
nand U7898 (N_7898,N_6001,N_5977);
or U7899 (N_7899,N_6636,N_5338);
and U7900 (N_7900,N_6258,N_7052);
nand U7901 (N_7901,N_6762,N_7114);
and U7902 (N_7902,N_5093,N_6266);
nand U7903 (N_7903,N_6152,N_6176);
or U7904 (N_7904,N_6129,N_5252);
nor U7905 (N_7905,N_6193,N_7158);
nor U7906 (N_7906,N_6112,N_6498);
and U7907 (N_7907,N_6869,N_5555);
and U7908 (N_7908,N_5074,N_7431);
or U7909 (N_7909,N_5226,N_5106);
and U7910 (N_7910,N_5359,N_5242);
nand U7911 (N_7911,N_7499,N_6188);
or U7912 (N_7912,N_6513,N_5427);
and U7913 (N_7913,N_6940,N_6195);
and U7914 (N_7914,N_6358,N_6076);
nor U7915 (N_7915,N_5397,N_5569);
or U7916 (N_7916,N_6120,N_5725);
and U7917 (N_7917,N_5849,N_5415);
nand U7918 (N_7918,N_7336,N_5498);
and U7919 (N_7919,N_7018,N_5279);
and U7920 (N_7920,N_6319,N_5766);
nand U7921 (N_7921,N_5450,N_5961);
and U7922 (N_7922,N_7067,N_6130);
or U7923 (N_7923,N_7345,N_6807);
nand U7924 (N_7924,N_5478,N_7046);
nor U7925 (N_7925,N_5207,N_6652);
or U7926 (N_7926,N_7218,N_5292);
nor U7927 (N_7927,N_7209,N_7385);
and U7928 (N_7928,N_6331,N_5966);
nor U7929 (N_7929,N_6492,N_5806);
nand U7930 (N_7930,N_7171,N_6679);
nor U7931 (N_7931,N_5386,N_5406);
nand U7932 (N_7932,N_5740,N_7200);
nor U7933 (N_7933,N_5009,N_5064);
nor U7934 (N_7934,N_7016,N_5175);
nor U7935 (N_7935,N_5038,N_6246);
nand U7936 (N_7936,N_6022,N_6572);
nor U7937 (N_7937,N_5818,N_5378);
or U7938 (N_7938,N_6489,N_5343);
or U7939 (N_7939,N_6101,N_6248);
or U7940 (N_7940,N_5635,N_7153);
nor U7941 (N_7941,N_6313,N_6437);
nor U7942 (N_7942,N_7350,N_7231);
or U7943 (N_7943,N_6646,N_6425);
nand U7944 (N_7944,N_6029,N_5833);
or U7945 (N_7945,N_6430,N_6252);
and U7946 (N_7946,N_6185,N_5687);
or U7947 (N_7947,N_6442,N_5614);
or U7948 (N_7948,N_7000,N_5972);
nand U7949 (N_7949,N_6201,N_5086);
or U7950 (N_7950,N_6978,N_6894);
nor U7951 (N_7951,N_5934,N_6448);
and U7952 (N_7952,N_7220,N_5522);
nand U7953 (N_7953,N_6229,N_5138);
or U7954 (N_7954,N_6007,N_5245);
nand U7955 (N_7955,N_5629,N_6132);
and U7956 (N_7956,N_5096,N_5788);
and U7957 (N_7957,N_5524,N_6506);
or U7958 (N_7958,N_7477,N_5215);
and U7959 (N_7959,N_5637,N_7029);
nand U7960 (N_7960,N_7055,N_7085);
nand U7961 (N_7961,N_5923,N_5700);
nand U7962 (N_7962,N_6688,N_6668);
or U7963 (N_7963,N_6932,N_5431);
and U7964 (N_7964,N_5382,N_5034);
nand U7965 (N_7965,N_5954,N_5249);
nand U7966 (N_7966,N_5198,N_6098);
or U7967 (N_7967,N_6138,N_5061);
nor U7968 (N_7968,N_6673,N_6747);
nand U7969 (N_7969,N_7254,N_5413);
and U7970 (N_7970,N_7452,N_5791);
or U7971 (N_7971,N_6124,N_7109);
nand U7972 (N_7972,N_6984,N_6588);
nor U7973 (N_7973,N_6203,N_5033);
nand U7974 (N_7974,N_5918,N_7278);
nor U7975 (N_7975,N_5541,N_6666);
or U7976 (N_7976,N_5826,N_5230);
nor U7977 (N_7977,N_5150,N_5620);
and U7978 (N_7978,N_5464,N_5601);
and U7979 (N_7979,N_6282,N_5099);
or U7980 (N_7980,N_5606,N_5131);
nor U7981 (N_7981,N_5804,N_6383);
and U7982 (N_7982,N_5285,N_5736);
nor U7983 (N_7983,N_5795,N_5331);
nand U7984 (N_7984,N_5947,N_5942);
or U7985 (N_7985,N_6259,N_7359);
or U7986 (N_7986,N_5660,N_6749);
or U7987 (N_7987,N_6378,N_7484);
or U7988 (N_7988,N_6535,N_5348);
or U7989 (N_7989,N_5419,N_6391);
nor U7990 (N_7990,N_6601,N_6213);
or U7991 (N_7991,N_6080,N_5550);
nor U7992 (N_7992,N_6596,N_7009);
nor U7993 (N_7993,N_5955,N_5971);
or U7994 (N_7994,N_5631,N_7247);
and U7995 (N_7995,N_7398,N_5032);
or U7996 (N_7996,N_5011,N_5563);
or U7997 (N_7997,N_6706,N_7368);
or U7998 (N_7998,N_6879,N_6877);
and U7999 (N_7999,N_7090,N_5717);
nor U8000 (N_8000,N_6276,N_7329);
or U8001 (N_8001,N_5006,N_6237);
nor U8002 (N_8002,N_5590,N_5615);
nor U8003 (N_8003,N_5417,N_5078);
nand U8004 (N_8004,N_7023,N_6473);
or U8005 (N_8005,N_6343,N_5240);
and U8006 (N_8006,N_6722,N_6443);
nor U8007 (N_8007,N_6832,N_6621);
nor U8008 (N_8008,N_5284,N_6833);
nor U8009 (N_8009,N_7456,N_6166);
or U8010 (N_8010,N_6324,N_6827);
and U8011 (N_8011,N_5578,N_6274);
nand U8012 (N_8012,N_5612,N_7307);
nand U8013 (N_8013,N_5287,N_6555);
and U8014 (N_8014,N_7157,N_7287);
and U8015 (N_8015,N_7242,N_7434);
nor U8016 (N_8016,N_6311,N_5645);
xnor U8017 (N_8017,N_6299,N_6992);
nand U8018 (N_8018,N_7464,N_5680);
nor U8019 (N_8019,N_5110,N_5515);
and U8020 (N_8020,N_7103,N_6012);
or U8021 (N_8021,N_7064,N_6495);
and U8022 (N_8022,N_6791,N_5871);
nor U8023 (N_8023,N_6859,N_6910);
nand U8024 (N_8024,N_5025,N_6767);
xor U8025 (N_8025,N_6089,N_6466);
nor U8026 (N_8026,N_5685,N_5295);
and U8027 (N_8027,N_6446,N_6336);
nor U8028 (N_8028,N_5054,N_5316);
or U8029 (N_8029,N_7040,N_7166);
or U8030 (N_8030,N_5251,N_6623);
and U8031 (N_8031,N_6024,N_5751);
nor U8032 (N_8032,N_6557,N_5714);
and U8033 (N_8033,N_6034,N_5960);
nor U8034 (N_8034,N_5368,N_6139);
nand U8035 (N_8035,N_5183,N_6284);
nor U8036 (N_8036,N_6109,N_5521);
or U8037 (N_8037,N_5235,N_5185);
or U8038 (N_8038,N_6729,N_5171);
and U8039 (N_8039,N_6122,N_5537);
xnor U8040 (N_8040,N_5282,N_7050);
and U8041 (N_8041,N_6169,N_5694);
nand U8042 (N_8042,N_6160,N_7318);
nor U8043 (N_8043,N_7409,N_6717);
nand U8044 (N_8044,N_5517,N_7310);
nand U8045 (N_8045,N_7457,N_5414);
nor U8046 (N_8046,N_6560,N_5258);
nor U8047 (N_8047,N_5001,N_5360);
or U8048 (N_8048,N_6459,N_6799);
nor U8049 (N_8049,N_5361,N_7421);
nand U8050 (N_8050,N_7462,N_6503);
and U8051 (N_8051,N_6301,N_6980);
nand U8052 (N_8052,N_6470,N_5979);
or U8053 (N_8053,N_6161,N_5145);
nand U8054 (N_8054,N_5357,N_6842);
and U8055 (N_8055,N_7075,N_5723);
nor U8056 (N_8056,N_5600,N_5937);
nand U8057 (N_8057,N_5206,N_5985);
and U8058 (N_8058,N_6561,N_6788);
or U8059 (N_8059,N_7272,N_5856);
nor U8060 (N_8060,N_7373,N_6915);
or U8061 (N_8061,N_5978,N_6841);
and U8062 (N_8062,N_5399,N_6996);
nand U8063 (N_8063,N_7324,N_6599);
nand U8064 (N_8064,N_6463,N_5046);
and U8065 (N_8065,N_5289,N_6566);
and U8066 (N_8066,N_6487,N_6332);
or U8067 (N_8067,N_6908,N_6897);
and U8068 (N_8068,N_6117,N_5116);
nand U8069 (N_8069,N_6223,N_7104);
and U8070 (N_8070,N_5503,N_7480);
nor U8071 (N_8071,N_5250,N_6285);
and U8072 (N_8072,N_6914,N_7328);
nand U8073 (N_8073,N_7178,N_5644);
or U8074 (N_8074,N_7192,N_6509);
nand U8075 (N_8075,N_5616,N_7478);
and U8076 (N_8076,N_5641,N_5863);
or U8077 (N_8077,N_5905,N_7335);
and U8078 (N_8078,N_6543,N_6074);
nor U8079 (N_8079,N_5440,N_7189);
nor U8080 (N_8080,N_6315,N_6451);
nand U8081 (N_8081,N_5778,N_6979);
or U8082 (N_8082,N_6447,N_5523);
nor U8083 (N_8083,N_5855,N_5105);
nor U8084 (N_8084,N_5886,N_5349);
nand U8085 (N_8085,N_5436,N_5401);
nor U8086 (N_8086,N_7474,N_5377);
or U8087 (N_8087,N_7071,N_6607);
nand U8088 (N_8088,N_6286,N_7496);
nor U8089 (N_8089,N_6197,N_5820);
and U8090 (N_8090,N_6817,N_5179);
nand U8091 (N_8091,N_6891,N_5081);
or U8092 (N_8092,N_5789,N_6895);
or U8093 (N_8093,N_7341,N_5799);
and U8094 (N_8094,N_6772,N_6538);
nand U8095 (N_8095,N_6025,N_7488);
nand U8096 (N_8096,N_5890,N_7162);
nor U8097 (N_8097,N_5062,N_6187);
and U8098 (N_8098,N_5844,N_7139);
and U8099 (N_8099,N_6522,N_5707);
and U8100 (N_8100,N_6144,N_5801);
and U8101 (N_8101,N_6701,N_6829);
nor U8102 (N_8102,N_5730,N_5917);
nand U8103 (N_8103,N_6625,N_6431);
or U8104 (N_8104,N_6380,N_6454);
nor U8105 (N_8105,N_6812,N_6225);
and U8106 (N_8106,N_7212,N_7423);
nor U8107 (N_8107,N_6704,N_7348);
and U8108 (N_8108,N_5028,N_5421);
nand U8109 (N_8109,N_6011,N_7319);
or U8110 (N_8110,N_6584,N_5194);
nand U8111 (N_8111,N_5574,N_5822);
and U8112 (N_8112,N_7426,N_5747);
nor U8113 (N_8113,N_5980,N_5182);
or U8114 (N_8114,N_6105,N_5108);
nor U8115 (N_8115,N_5097,N_6785);
and U8116 (N_8116,N_5491,N_6870);
nor U8117 (N_8117,N_6880,N_5897);
nand U8118 (N_8118,N_5611,N_6602);
and U8119 (N_8119,N_5233,N_6068);
nor U8120 (N_8120,N_5412,N_7386);
or U8121 (N_8121,N_7455,N_5570);
nor U8122 (N_8122,N_5190,N_6407);
or U8123 (N_8123,N_6260,N_7388);
nand U8124 (N_8124,N_6875,N_7138);
nor U8125 (N_8125,N_7079,N_5371);
and U8126 (N_8126,N_5657,N_6171);
and U8127 (N_8127,N_5339,N_7435);
and U8128 (N_8128,N_5697,N_7355);
and U8129 (N_8129,N_7383,N_6527);
or U8130 (N_8130,N_5117,N_5124);
nor U8131 (N_8131,N_5664,N_5626);
or U8132 (N_8132,N_6532,N_5050);
or U8133 (N_8133,N_6567,N_6254);
nand U8134 (N_8134,N_5860,N_5652);
or U8135 (N_8135,N_6715,N_6577);
nor U8136 (N_8136,N_6872,N_7084);
and U8137 (N_8137,N_5461,N_5704);
nor U8138 (N_8138,N_7363,N_6972);
and U8139 (N_8139,N_6481,N_6809);
and U8140 (N_8140,N_5127,N_5405);
or U8141 (N_8141,N_5388,N_5535);
nor U8142 (N_8142,N_7497,N_5259);
nor U8143 (N_8143,N_6536,N_5598);
and U8144 (N_8144,N_7206,N_5015);
nor U8145 (N_8145,N_6598,N_7049);
or U8146 (N_8146,N_6290,N_6419);
xor U8147 (N_8147,N_6226,N_5308);
or U8148 (N_8148,N_6436,N_6497);
or U8149 (N_8149,N_6757,N_5831);
nand U8150 (N_8150,N_5232,N_7428);
nor U8151 (N_8151,N_6795,N_5533);
nand U8152 (N_8152,N_6093,N_5212);
and U8153 (N_8153,N_7135,N_5007);
nand U8154 (N_8154,N_6849,N_6782);
or U8155 (N_8155,N_6263,N_6309);
and U8156 (N_8156,N_6154,N_6804);
or U8157 (N_8157,N_5273,N_7251);
or U8158 (N_8158,N_6834,N_5703);
nand U8159 (N_8159,N_5075,N_6728);
nand U8160 (N_8160,N_7332,N_6783);
nand U8161 (N_8161,N_7312,N_6116);
nor U8162 (N_8162,N_6292,N_5571);
nor U8163 (N_8163,N_7353,N_7080);
nor U8164 (N_8164,N_5774,N_5797);
nor U8165 (N_8165,N_5489,N_6512);
nor U8166 (N_8166,N_5173,N_5689);
nand U8167 (N_8167,N_6047,N_5196);
or U8168 (N_8168,N_6550,N_5544);
or U8169 (N_8169,N_7295,N_6866);
and U8170 (N_8170,N_5568,N_6075);
and U8171 (N_8171,N_5426,N_7119);
nand U8172 (N_8172,N_5223,N_7232);
nand U8173 (N_8173,N_6405,N_5486);
or U8174 (N_8174,N_6661,N_5428);
and U8175 (N_8175,N_5888,N_5683);
xnor U8176 (N_8176,N_7056,N_7404);
or U8177 (N_8177,N_6603,N_7303);
nand U8178 (N_8178,N_7400,N_7450);
and U8179 (N_8179,N_6457,N_6801);
and U8180 (N_8180,N_7357,N_6900);
nor U8181 (N_8181,N_5224,N_6857);
nor U8182 (N_8182,N_5479,N_5661);
nor U8183 (N_8183,N_6743,N_6758);
and U8184 (N_8184,N_6155,N_6052);
nor U8185 (N_8185,N_6569,N_7150);
or U8186 (N_8186,N_5812,N_6200);
nor U8187 (N_8187,N_6173,N_6863);
nor U8188 (N_8188,N_7314,N_6708);
nand U8189 (N_8189,N_5083,N_5184);
or U8190 (N_8190,N_5696,N_6346);
nand U8191 (N_8191,N_5085,N_5220);
nand U8192 (N_8192,N_6848,N_5337);
nor U8193 (N_8193,N_6192,N_7444);
nand U8194 (N_8194,N_5476,N_6591);
or U8195 (N_8195,N_7205,N_5154);
nand U8196 (N_8196,N_7270,N_6220);
nor U8197 (N_8197,N_5209,N_6647);
nand U8198 (N_8198,N_5102,N_6777);
nand U8199 (N_8199,N_7293,N_6395);
nor U8200 (N_8200,N_6696,N_7311);
or U8201 (N_8201,N_6438,N_6106);
or U8202 (N_8202,N_6190,N_6676);
and U8203 (N_8203,N_6433,N_5354);
nand U8204 (N_8204,N_5301,N_7436);
and U8205 (N_8205,N_5780,N_5238);
nand U8206 (N_8206,N_7414,N_6564);
nor U8207 (N_8207,N_6501,N_5069);
nor U8208 (N_8208,N_7051,N_5193);
nor U8209 (N_8209,N_6255,N_5304);
nand U8210 (N_8210,N_5670,N_6341);
nand U8211 (N_8211,N_5781,N_5168);
or U8212 (N_8212,N_5900,N_6219);
nor U8213 (N_8213,N_6230,N_7418);
nor U8214 (N_8214,N_7334,N_7025);
nor U8215 (N_8215,N_6995,N_6178);
nand U8216 (N_8216,N_7169,N_6705);
and U8217 (N_8217,N_7360,N_5014);
nor U8218 (N_8218,N_5147,N_7406);
nand U8219 (N_8219,N_5165,N_6962);
nor U8220 (N_8220,N_5532,N_6568);
or U8221 (N_8221,N_7343,N_7208);
nand U8222 (N_8222,N_7184,N_5643);
nor U8223 (N_8223,N_7081,N_5135);
and U8224 (N_8224,N_5883,N_7472);
nand U8225 (N_8225,N_5510,N_6907);
nand U8226 (N_8226,N_5132,N_6386);
and U8227 (N_8227,N_5909,N_6049);
xor U8228 (N_8228,N_6681,N_5756);
and U8229 (N_8229,N_5153,N_6669);
nand U8230 (N_8230,N_5247,N_7282);
nand U8231 (N_8231,N_7317,N_7037);
nand U8232 (N_8232,N_5065,N_5829);
nand U8233 (N_8233,N_7005,N_6864);
nand U8234 (N_8234,N_6374,N_5072);
and U8235 (N_8235,N_7132,N_6614);
or U8236 (N_8236,N_5262,N_6662);
or U8237 (N_8237,N_7207,N_6175);
and U8238 (N_8238,N_6250,N_7001);
nor U8239 (N_8239,N_5728,N_6721);
nand U8240 (N_8240,N_5577,N_5530);
nand U8241 (N_8241,N_7361,N_6924);
xor U8242 (N_8242,N_7172,N_7442);
or U8243 (N_8243,N_7384,N_5211);
and U8244 (N_8244,N_5602,N_7183);
nor U8245 (N_8245,N_5271,N_5621);
or U8246 (N_8246,N_6202,N_6233);
nor U8247 (N_8247,N_5792,N_6320);
nor U8248 (N_8248,N_6644,N_6753);
and U8249 (N_8249,N_5317,N_5777);
nand U8250 (N_8250,N_6811,N_7203);
or U8251 (N_8251,N_6394,N_6530);
nand U8252 (N_8252,N_6919,N_7346);
nor U8253 (N_8253,N_7491,N_6667);
or U8254 (N_8254,N_7429,N_7115);
nand U8255 (N_8255,N_6423,N_5743);
or U8256 (N_8256,N_6435,N_7083);
nand U8257 (N_8257,N_6796,N_6768);
nor U8258 (N_8258,N_6691,N_7291);
nor U8259 (N_8259,N_5765,N_5335);
nor U8260 (N_8260,N_5141,N_6756);
and U8261 (N_8261,N_6740,N_6505);
nor U8262 (N_8262,N_5794,N_6912);
or U8263 (N_8263,N_5474,N_6164);
nand U8264 (N_8264,N_6794,N_6627);
or U8265 (N_8265,N_7424,N_5325);
nor U8266 (N_8266,N_6573,N_6540);
nor U8267 (N_8267,N_6726,N_5432);
nor U8268 (N_8268,N_5416,N_6519);
and U8269 (N_8269,N_5891,N_6884);
nand U8270 (N_8270,N_6511,N_5924);
nand U8271 (N_8271,N_6790,N_6960);
nand U8272 (N_8272,N_7340,N_6671);
and U8273 (N_8273,N_5987,N_5594);
nand U8274 (N_8274,N_6998,N_5346);
and U8275 (N_8275,N_6986,N_6316);
or U8276 (N_8276,N_5126,N_5919);
and U8277 (N_8277,N_7237,N_5939);
or U8278 (N_8278,N_5762,N_6147);
nand U8279 (N_8279,N_6539,N_5446);
nand U8280 (N_8280,N_5118,N_5835);
and U8281 (N_8281,N_5748,N_5058);
nand U8282 (N_8282,N_6151,N_6278);
or U8283 (N_8283,N_6565,N_5638);
nand U8284 (N_8284,N_5089,N_6294);
or U8285 (N_8285,N_6967,N_5455);
or U8286 (N_8286,N_7122,N_6537);
and U8287 (N_8287,N_6905,N_5068);
and U8288 (N_8288,N_7107,N_6634);
and U8289 (N_8289,N_5494,N_5663);
nand U8290 (N_8290,N_6970,N_5422);
nand U8291 (N_8291,N_5724,N_7070);
and U8292 (N_8292,N_6057,N_6633);
nor U8293 (N_8293,N_6939,N_5549);
nand U8294 (N_8294,N_6402,N_6611);
or U8295 (N_8295,N_5861,N_5458);
nor U8296 (N_8296,N_7283,N_5878);
nand U8297 (N_8297,N_6630,N_5332);
or U8298 (N_8298,N_5587,N_6043);
nand U8299 (N_8299,N_5122,N_5079);
nand U8300 (N_8300,N_6428,N_7440);
nor U8301 (N_8301,N_5439,N_6635);
and U8302 (N_8302,N_6231,N_5735);
and U8303 (N_8303,N_7236,N_6876);
or U8304 (N_8304,N_5253,N_7454);
nor U8305 (N_8305,N_6399,N_5373);
nor U8306 (N_8306,N_6330,N_5603);
and U8307 (N_8307,N_7143,N_7133);
and U8308 (N_8308,N_5745,N_5481);
and U8309 (N_8309,N_6909,N_5760);
nor U8310 (N_8310,N_7038,N_5516);
nor U8311 (N_8311,N_5492,N_6615);
and U8312 (N_8312,N_6820,N_5457);
nor U8313 (N_8313,N_7177,N_7425);
nor U8314 (N_8314,N_5060,N_5396);
and U8315 (N_8315,N_5379,N_6589);
nor U8316 (N_8316,N_5163,N_5605);
and U8317 (N_8317,N_6771,N_7323);
and U8318 (N_8318,N_7482,N_7054);
and U8319 (N_8319,N_6816,N_6684);
and U8320 (N_8320,N_7487,N_6062);
and U8321 (N_8321,N_5705,N_5582);
or U8322 (N_8322,N_7489,N_6370);
and U8323 (N_8323,N_6474,N_6177);
or U8324 (N_8324,N_6886,N_5798);
or U8325 (N_8325,N_6818,N_6312);
nor U8326 (N_8326,N_6069,N_6142);
and U8327 (N_8327,N_5513,N_5387);
and U8328 (N_8328,N_6524,N_6401);
nand U8329 (N_8329,N_5454,N_5204);
nand U8330 (N_8330,N_7130,N_5423);
or U8331 (N_8331,N_5729,N_5767);
and U8332 (N_8332,N_7145,N_6385);
or U8333 (N_8333,N_7285,N_6742);
and U8334 (N_8334,N_7412,N_6805);
and U8335 (N_8335,N_5030,N_6440);
or U8336 (N_8336,N_6510,N_5310);
nor U8337 (N_8337,N_6504,N_5468);
nand U8338 (N_8338,N_6493,N_6923);
nor U8339 (N_8339,N_5981,N_6326);
or U8340 (N_8340,N_5667,N_5418);
nand U8341 (N_8341,N_5921,N_7498);
or U8342 (N_8342,N_6922,N_6198);
nand U8343 (N_8343,N_7224,N_5757);
nor U8344 (N_8344,N_6352,N_7394);
nor U8345 (N_8345,N_6482,N_6131);
and U8346 (N_8346,N_6649,N_6390);
and U8347 (N_8347,N_5588,N_7445);
or U8348 (N_8348,N_7378,N_6999);
nand U8349 (N_8349,N_6216,N_6483);
and U8350 (N_8350,N_5561,N_6021);
nand U8351 (N_8351,N_6471,N_6926);
nand U8352 (N_8352,N_6733,N_6362);
nand U8353 (N_8353,N_6491,N_6789);
and U8354 (N_8354,N_7481,N_7089);
and U8355 (N_8355,N_5773,N_6153);
nand U8356 (N_8356,N_6518,N_6382);
nor U8357 (N_8357,N_5893,N_6351);
xnor U8358 (N_8358,N_7389,N_6724);
nor U8359 (N_8359,N_6654,N_7379);
nor U8360 (N_8360,N_5839,N_7163);
nor U8361 (N_8361,N_7256,N_5691);
or U8362 (N_8362,N_6269,N_6781);
or U8363 (N_8363,N_7327,N_6211);
and U8364 (N_8364,N_6624,N_5143);
and U8365 (N_8365,N_7137,N_6663);
or U8366 (N_8366,N_5056,N_5268);
nand U8367 (N_8367,N_5508,N_5876);
nand U8368 (N_8368,N_5363,N_6141);
or U8369 (N_8369,N_5901,N_5639);
nor U8370 (N_8370,N_5026,N_5438);
or U8371 (N_8371,N_6350,N_5881);
or U8372 (N_8372,N_7170,N_6719);
or U8373 (N_8373,N_7072,N_6026);
nor U8374 (N_8374,N_6526,N_6951);
nor U8375 (N_8375,N_5887,N_5793);
and U8376 (N_8376,N_5340,N_6145);
and U8377 (N_8377,N_7197,N_5959);
nand U8378 (N_8378,N_5993,N_6020);
or U8379 (N_8379,N_6763,N_7461);
nor U8380 (N_8380,N_5229,N_6039);
nor U8381 (N_8381,N_6873,N_6027);
nand U8382 (N_8382,N_7380,N_5021);
and U8383 (N_8383,N_5467,N_5475);
and U8384 (N_8384,N_7129,N_6672);
and U8385 (N_8385,N_6424,N_6348);
nor U8386 (N_8386,N_5389,N_6575);
or U8387 (N_8387,N_7255,N_7106);
and U8388 (N_8388,N_6017,N_6698);
or U8389 (N_8389,N_7144,N_7304);
nor U8390 (N_8390,N_5807,N_5040);
and U8391 (N_8391,N_7326,N_5869);
nand U8392 (N_8392,N_7045,N_5754);
nor U8393 (N_8393,N_7316,N_7175);
or U8394 (N_8394,N_6494,N_6583);
nor U8395 (N_8395,N_7365,N_6958);
and U8396 (N_8396,N_7342,N_6355);
and U8397 (N_8397,N_6746,N_5092);
nor U8398 (N_8398,N_6778,N_5402);
nand U8399 (N_8399,N_5534,N_6040);
xor U8400 (N_8400,N_7369,N_6847);
nor U8401 (N_8401,N_5275,N_5581);
or U8402 (N_8402,N_7331,N_6620);
nand U8403 (N_8403,N_6741,N_6308);
xor U8404 (N_8404,N_7396,N_6245);
and U8405 (N_8405,N_5734,N_6931);
and U8406 (N_8406,N_7124,N_5686);
or U8407 (N_8407,N_5519,N_5932);
nor U8408 (N_8408,N_5802,N_6851);
nand U8409 (N_8409,N_6545,N_7195);
and U8410 (N_8410,N_5120,N_5896);
nand U8411 (N_8411,N_5540,N_5854);
or U8412 (N_8412,N_6159,N_5646);
nor U8413 (N_8413,N_5912,N_6968);
nand U8414 (N_8414,N_6594,N_6898);
and U8415 (N_8415,N_6610,N_5948);
nand U8416 (N_8416,N_7261,N_6477);
and U8417 (N_8417,N_7419,N_5828);
or U8418 (N_8418,N_5936,N_5553);
or U8419 (N_8419,N_6534,N_6045);
nand U8420 (N_8420,N_5176,N_6418);
nand U8421 (N_8421,N_6920,N_6865);
nand U8422 (N_8422,N_6262,N_5125);
and U8423 (N_8423,N_6871,N_5013);
and U8424 (N_8424,N_5824,N_5542);
and U8425 (N_8425,N_5864,N_6840);
xor U8426 (N_8426,N_7301,N_6692);
and U8427 (N_8427,N_5830,N_6426);
and U8428 (N_8428,N_6082,N_5566);
and U8429 (N_8429,N_5170,N_7043);
or U8430 (N_8430,N_6660,N_5836);
and U8431 (N_8431,N_7370,N_7266);
or U8432 (N_8432,N_5018,N_5134);
and U8433 (N_8433,N_6035,N_6478);
and U8434 (N_8434,N_6904,N_7082);
nor U8435 (N_8435,N_6639,N_7216);
nand U8436 (N_8436,N_7102,N_7201);
or U8437 (N_8437,N_7375,N_5019);
nor U8438 (N_8438,N_5016,N_5197);
and U8439 (N_8439,N_6734,N_5562);
nand U8440 (N_8440,N_5266,N_6363);
and U8441 (N_8441,N_6028,N_5677);
nand U8442 (N_8442,N_6921,N_7156);
nor U8443 (N_8443,N_7284,N_5529);
or U8444 (N_8444,N_5538,N_6393);
and U8445 (N_8445,N_6086,N_6590);
nand U8446 (N_8446,N_7495,N_6271);
nor U8447 (N_8447,N_5351,N_5333);
or U8448 (N_8448,N_5927,N_5755);
nand U8449 (N_8449,N_6462,N_5341);
and U8450 (N_8450,N_5770,N_5640);
or U8451 (N_8451,N_5430,N_5580);
and U8452 (N_8452,N_6050,N_5100);
nand U8453 (N_8453,N_5255,N_5943);
or U8454 (N_8454,N_5776,N_5940);
nor U8455 (N_8455,N_6901,N_6709);
and U8456 (N_8456,N_6429,N_5790);
nor U8457 (N_8457,N_7087,N_6469);
xor U8458 (N_8458,N_6349,N_6168);
and U8459 (N_8459,N_5037,N_6256);
nand U8460 (N_8460,N_7033,N_6365);
nor U8461 (N_8461,N_6183,N_5465);
and U8462 (N_8462,N_6690,N_6797);
nor U8463 (N_8463,N_7113,N_6703);
nor U8464 (N_8464,N_5998,N_5277);
nand U8465 (N_8465,N_7276,N_6760);
nor U8466 (N_8466,N_6710,N_6878);
nand U8467 (N_8467,N_5136,N_6930);
nor U8468 (N_8468,N_7057,N_6830);
nand U8469 (N_8469,N_6340,N_6297);
nand U8470 (N_8470,N_7020,N_7093);
and U8471 (N_8471,N_6452,N_6853);
nand U8472 (N_8472,N_5227,N_6174);
and U8473 (N_8473,N_5202,N_6731);
nor U8474 (N_8474,N_6657,N_7405);
or U8475 (N_8475,N_7277,N_5654);
and U8476 (N_8476,N_7250,N_5698);
and U8477 (N_8477,N_5761,N_5819);
nor U8478 (N_8478,N_5695,N_5884);
nor U8479 (N_8479,N_7039,N_5047);
or U8480 (N_8480,N_7243,N_6475);
nand U8481 (N_8481,N_7422,N_6456);
nor U8482 (N_8482,N_7094,N_5922);
nand U8483 (N_8483,N_6956,N_5546);
nor U8484 (N_8484,N_6971,N_6210);
nor U8485 (N_8485,N_6205,N_5974);
and U8486 (N_8486,N_5655,N_6831);
and U8487 (N_8487,N_7217,N_5738);
and U8488 (N_8488,N_5311,N_5390);
nor U8489 (N_8489,N_6127,N_6460);
nor U8490 (N_8490,N_6108,N_6277);
nor U8491 (N_8491,N_6373,N_7465);
nand U8492 (N_8492,N_5090,N_5404);
and U8493 (N_8493,N_6766,N_5327);
nand U8494 (N_8494,N_5976,N_5298);
nand U8495 (N_8495,N_5042,N_7134);
nor U8496 (N_8496,N_6953,N_6659);
and U8497 (N_8497,N_6656,N_5471);
nor U8498 (N_8498,N_5087,N_6157);
xor U8499 (N_8499,N_6965,N_5501);
nand U8500 (N_8500,N_5052,N_5048);
nor U8501 (N_8501,N_5733,N_6881);
and U8502 (N_8502,N_7240,N_5162);
nand U8503 (N_8503,N_5309,N_5320);
or U8504 (N_8504,N_5024,N_5873);
or U8505 (N_8505,N_6556,N_5630);
or U8506 (N_8506,N_5297,N_6808);
or U8507 (N_8507,N_6033,N_5104);
and U8508 (N_8508,N_7411,N_5356);
nand U8509 (N_8509,N_5821,N_6680);
xnor U8510 (N_8510,N_6888,N_6306);
or U8511 (N_8511,N_6217,N_5460);
and U8512 (N_8512,N_5862,N_7077);
or U8513 (N_8513,N_5365,N_5231);
xor U8514 (N_8514,N_6165,N_7320);
nor U8515 (N_8515,N_5059,N_5572);
nor U8516 (N_8516,N_5618,N_5642);
and U8517 (N_8517,N_6018,N_6903);
or U8518 (N_8518,N_6485,N_5159);
nor U8519 (N_8519,N_5722,N_5445);
nand U8520 (N_8520,N_6593,N_6613);
nand U8521 (N_8521,N_5586,N_5002);
nor U8522 (N_8522,N_5552,N_7233);
nor U8523 (N_8523,N_6239,N_7420);
nand U8524 (N_8524,N_7210,N_6580);
nand U8525 (N_8525,N_5585,N_5187);
nand U8526 (N_8526,N_7230,N_7449);
nand U8527 (N_8527,N_6651,N_6162);
or U8528 (N_8528,N_5008,N_7165);
and U8529 (N_8529,N_7167,N_6619);
and U8530 (N_8530,N_5938,N_6123);
and U8531 (N_8531,N_6981,N_5499);
or U8532 (N_8532,N_7299,N_5192);
and U8533 (N_8533,N_7430,N_5313);
nand U8534 (N_8534,N_6835,N_6268);
nand U8535 (N_8535,N_6683,N_7222);
nand U8536 (N_8536,N_5706,N_6868);
or U8537 (N_8537,N_6775,N_6265);
nand U8538 (N_8538,N_5668,N_7325);
or U8539 (N_8539,N_6815,N_5779);
or U8540 (N_8540,N_7099,N_7117);
or U8541 (N_8541,N_7367,N_5264);
nor U8542 (N_8542,N_6359,N_5565);
and U8543 (N_8543,N_7296,N_7215);
nand U8544 (N_8544,N_5246,N_5469);
and U8545 (N_8545,N_6950,N_5608);
nand U8546 (N_8546,N_5477,N_7168);
and U8547 (N_8547,N_6051,N_5319);
nand U8548 (N_8548,N_6798,N_7338);
nand U8549 (N_8549,N_5693,N_5003);
nand U8550 (N_8550,N_5576,N_7229);
and U8551 (N_8551,N_5514,N_7120);
or U8552 (N_8552,N_5930,N_6002);
and U8553 (N_8553,N_6737,N_5688);
or U8554 (N_8554,N_5604,N_5362);
nor U8555 (N_8555,N_6761,N_5701);
nor U8556 (N_8556,N_5239,N_5619);
and U8557 (N_8557,N_7408,N_6345);
nor U8558 (N_8558,N_6417,N_6335);
nor U8559 (N_8559,N_6997,N_5906);
xor U8560 (N_8560,N_5443,N_5649);
or U8561 (N_8561,N_5931,N_6015);
nor U8562 (N_8562,N_6135,N_5148);
and U8563 (N_8563,N_6641,N_5840);
nand U8564 (N_8564,N_5857,N_5531);
or U8565 (N_8565,N_5410,N_5674);
nor U8566 (N_8566,N_5300,N_6307);
nor U8567 (N_8567,N_5372,N_7187);
or U8568 (N_8568,N_5509,N_5201);
xnor U8569 (N_8569,N_5107,N_5672);
or U8570 (N_8570,N_6305,N_7196);
and U8571 (N_8571,N_6372,N_6889);
nor U8572 (N_8572,N_7382,N_7173);
and U8573 (N_8573,N_7141,N_6009);
or U8574 (N_8574,N_5903,N_6541);
nand U8575 (N_8575,N_7105,N_5442);
and U8576 (N_8576,N_6675,N_5525);
or U8577 (N_8577,N_7469,N_5112);
or U8578 (N_8578,N_7128,N_6687);
nor U8579 (N_8579,N_7402,N_6653);
nor U8580 (N_8580,N_5142,N_6338);
and U8581 (N_8581,N_6693,N_6612);
nor U8582 (N_8582,N_6935,N_6235);
nand U8583 (N_8583,N_6369,N_7186);
nor U8584 (N_8584,N_6291,N_5146);
and U8585 (N_8585,N_7485,N_5935);
nand U8586 (N_8586,N_5370,N_7246);
nand U8587 (N_8587,N_6943,N_5595);
or U8588 (N_8588,N_5727,N_6892);
and U8589 (N_8589,N_6813,N_5968);
or U8590 (N_8590,N_5753,N_6855);
nand U8591 (N_8591,N_6065,N_5769);
and U8592 (N_8592,N_6819,N_6618);
and U8593 (N_8593,N_5634,N_7223);
nor U8594 (N_8594,N_5702,N_5128);
and U8595 (N_8595,N_6084,N_6500);
nor U8596 (N_8596,N_7042,N_7110);
or U8597 (N_8597,N_5243,N_6994);
nor U8598 (N_8598,N_7265,N_7010);
and U8599 (N_8599,N_5951,N_5669);
nand U8600 (N_8600,N_6754,N_5963);
and U8601 (N_8601,N_5908,N_5928);
nand U8602 (N_8602,N_6434,N_5290);
nor U8603 (N_8603,N_6600,N_5334);
and U8604 (N_8604,N_7439,N_6206);
xor U8605 (N_8605,N_5329,N_7136);
nor U8606 (N_8606,N_7193,N_7152);
nand U8607 (N_8607,N_5409,N_6232);
or U8608 (N_8608,N_5490,N_7294);
and U8609 (N_8609,N_5005,N_6786);
or U8610 (N_8610,N_6689,N_7015);
or U8611 (N_8611,N_6445,N_6677);
and U8612 (N_8612,N_6730,N_5997);
nor U8613 (N_8613,N_6845,N_5248);
nor U8614 (N_8614,N_5746,N_5101);
nand U8615 (N_8615,N_7036,N_5658);
nor U8616 (N_8616,N_7399,N_7490);
nand U8617 (N_8617,N_6658,N_6287);
or U8618 (N_8618,N_7479,N_5984);
or U8619 (N_8619,N_5174,N_6046);
nand U8620 (N_8620,N_5916,N_5151);
nor U8621 (N_8621,N_5299,N_5020);
and U8622 (N_8622,N_6887,N_6643);
nor U8623 (N_8623,N_7159,N_6563);
or U8624 (N_8624,N_5463,N_7239);
or U8625 (N_8625,N_6063,N_7174);
or U8626 (N_8626,N_6852,N_6993);
and U8627 (N_8627,N_7381,N_5907);
or U8628 (N_8628,N_6987,N_7154);
nand U8629 (N_8629,N_5484,N_6665);
nand U8630 (N_8630,N_5004,N_6243);
and U8631 (N_8631,N_6072,N_6642);
nand U8632 (N_8632,N_7116,N_7088);
nand U8633 (N_8633,N_5613,N_6353);
xor U8634 (N_8634,N_6725,N_5684);
or U8635 (N_8635,N_7483,N_5811);
and U8636 (N_8636,N_5868,N_7356);
nand U8637 (N_8637,N_5195,N_6403);
or U8638 (N_8638,N_6191,N_6328);
or U8639 (N_8639,N_7458,N_5944);
nand U8640 (N_8640,N_5527,N_5898);
or U8641 (N_8641,N_5560,N_6048);
nor U8642 (N_8642,N_6787,N_5288);
and U8643 (N_8643,N_6713,N_6626);
and U8644 (N_8644,N_5875,N_6597);
or U8645 (N_8645,N_6945,N_5573);
nor U8646 (N_8646,N_6578,N_6723);
nor U8647 (N_8647,N_5874,N_5084);
nor U8648 (N_8648,N_5088,N_7390);
nor U8649 (N_8649,N_5305,N_6170);
xnor U8650 (N_8650,N_6005,N_5991);
nor U8651 (N_8651,N_7321,N_5130);
nor U8652 (N_8652,N_6182,N_7149);
nor U8653 (N_8653,N_6515,N_5659);
and U8654 (N_8654,N_6966,N_5726);
nand U8655 (N_8655,N_7017,N_7245);
nor U8656 (N_8656,N_7148,N_6053);
or U8657 (N_8657,N_5186,N_5877);
nor U8658 (N_8658,N_5607,N_5384);
and U8659 (N_8659,N_6409,N_7292);
nor U8660 (N_8660,N_6119,N_5483);
nand U8661 (N_8661,N_5675,N_6234);
or U8662 (N_8662,N_6882,N_5098);
nor U8663 (N_8663,N_7290,N_5261);
and U8664 (N_8664,N_7008,N_6156);
nand U8665 (N_8665,N_6670,N_5899);
or U8666 (N_8666,N_6468,N_5915);
nand U8667 (N_8667,N_6180,N_5892);
nand U8668 (N_8668,N_7302,N_6629);
nor U8669 (N_8669,N_7151,N_5071);
or U8670 (N_8670,N_7160,N_6765);
and U8671 (N_8671,N_6077,N_5286);
and U8672 (N_8672,N_5567,N_6389);
nand U8673 (N_8673,N_6582,N_7397);
nand U8674 (N_8674,N_5545,N_6099);
or U8675 (N_8675,N_5208,N_5902);
or U8676 (N_8676,N_5784,N_5029);
or U8677 (N_8677,N_7330,N_7274);
nand U8678 (N_8678,N_6377,N_6114);
or U8679 (N_8679,N_5692,N_5787);
or U8680 (N_8680,N_5808,N_6115);
or U8681 (N_8681,N_5759,N_5411);
and U8682 (N_8682,N_5632,N_5859);
or U8683 (N_8683,N_6645,N_7351);
or U8684 (N_8684,N_5910,N_6163);
and U8685 (N_8685,N_5848,N_6113);
nor U8686 (N_8686,N_5653,N_7297);
or U8687 (N_8687,N_5539,N_6146);
nand U8688 (N_8688,N_6079,N_5167);
and U8689 (N_8689,N_5647,N_6392);
nor U8690 (N_8690,N_6023,N_6107);
and U8691 (N_8691,N_5449,N_7044);
nand U8692 (N_8692,N_5772,N_5403);
xnor U8693 (N_8693,N_6838,N_5957);
or U8694 (N_8694,N_5992,N_7006);
and U8695 (N_8695,N_6860,N_5556);
and U8696 (N_8696,N_7253,N_5472);
or U8697 (N_8697,N_5673,N_7048);
nor U8698 (N_8698,N_7337,N_6699);
and U8699 (N_8699,N_6253,N_5155);
nand U8700 (N_8700,N_6318,N_5732);
or U8701 (N_8701,N_6379,N_6449);
nor U8702 (N_8702,N_5094,N_6078);
or U8703 (N_8703,N_6977,N_6748);
and U8704 (N_8704,N_5866,N_6874);
nor U8705 (N_8705,N_6283,N_5558);
and U8706 (N_8706,N_5121,N_5485);
or U8707 (N_8707,N_6792,N_6548);
nor U8708 (N_8708,N_5786,N_5043);
nor U8709 (N_8709,N_6759,N_7185);
nand U8710 (N_8710,N_7300,N_5314);
or U8711 (N_8711,N_7213,N_6826);
nand U8712 (N_8712,N_6032,N_6554);
and U8713 (N_8713,N_5070,N_7376);
and U8714 (N_8714,N_6531,N_6711);
nor U8715 (N_8715,N_7100,N_6640);
nor U8716 (N_8716,N_6694,N_7024);
nand U8717 (N_8717,N_6961,N_7313);
or U8718 (N_8718,N_6118,N_5712);
xor U8719 (N_8719,N_6570,N_6964);
or U8720 (N_8720,N_6985,N_5520);
and U8721 (N_8721,N_6314,N_6814);
nor U8722 (N_8722,N_6486,N_5965);
nor U8723 (N_8723,N_7068,N_5385);
or U8724 (N_8724,N_5027,N_5482);
nor U8725 (N_8725,N_6674,N_7059);
nor U8726 (N_8726,N_5969,N_6087);
nor U8727 (N_8727,N_6885,N_7211);
nor U8728 (N_8728,N_7118,N_6189);
and U8729 (N_8729,N_7161,N_7078);
nor U8730 (N_8730,N_6413,N_5512);
nor U8731 (N_8731,N_7027,N_6822);
nand U8732 (N_8732,N_7073,N_6727);
or U8733 (N_8733,N_6304,N_7437);
nor U8734 (N_8734,N_6631,N_5809);
and U8735 (N_8735,N_6134,N_7432);
or U8736 (N_8736,N_5882,N_6133);
or U8737 (N_8737,N_5274,N_7204);
nor U8738 (N_8738,N_5139,N_5218);
or U8739 (N_8739,N_5502,N_6412);
xor U8740 (N_8740,N_5989,N_5267);
nand U8741 (N_8741,N_5817,N_7475);
and U8742 (N_8742,N_6933,N_6810);
and U8743 (N_8743,N_6800,N_7235);
and U8744 (N_8744,N_7366,N_5178);
nand U8745 (N_8745,N_6273,N_7459);
nand U8746 (N_8746,N_6325,N_6544);
nor U8747 (N_8747,N_5169,N_5077);
and U8748 (N_8748,N_5843,N_6752);
or U8749 (N_8749,N_5291,N_6529);
nand U8750 (N_8750,N_5252,N_5141);
nor U8751 (N_8751,N_5957,N_5809);
and U8752 (N_8752,N_5056,N_7304);
and U8753 (N_8753,N_7137,N_6054);
nor U8754 (N_8754,N_5755,N_6328);
and U8755 (N_8755,N_7270,N_6692);
nor U8756 (N_8756,N_5897,N_6965);
nand U8757 (N_8757,N_6252,N_5726);
nand U8758 (N_8758,N_6107,N_5848);
or U8759 (N_8759,N_6034,N_5359);
nor U8760 (N_8760,N_7286,N_5092);
and U8761 (N_8761,N_6795,N_7154);
nor U8762 (N_8762,N_6136,N_5078);
and U8763 (N_8763,N_5056,N_6625);
xor U8764 (N_8764,N_5675,N_5571);
nor U8765 (N_8765,N_5862,N_5954);
nor U8766 (N_8766,N_5922,N_5661);
xor U8767 (N_8767,N_7478,N_5013);
nand U8768 (N_8768,N_6311,N_5181);
xnor U8769 (N_8769,N_5088,N_6212);
or U8770 (N_8770,N_6562,N_5593);
nor U8771 (N_8771,N_5486,N_6089);
or U8772 (N_8772,N_5224,N_6581);
nor U8773 (N_8773,N_5639,N_5336);
and U8774 (N_8774,N_5689,N_6694);
nand U8775 (N_8775,N_7020,N_5795);
nand U8776 (N_8776,N_7131,N_7127);
and U8777 (N_8777,N_5739,N_6846);
nor U8778 (N_8778,N_5554,N_5948);
nor U8779 (N_8779,N_5728,N_7285);
nand U8780 (N_8780,N_6347,N_5892);
nor U8781 (N_8781,N_7213,N_5805);
nor U8782 (N_8782,N_6635,N_5547);
or U8783 (N_8783,N_7357,N_5556);
nand U8784 (N_8784,N_7076,N_6405);
nor U8785 (N_8785,N_6029,N_5807);
or U8786 (N_8786,N_7222,N_5760);
and U8787 (N_8787,N_6780,N_6618);
and U8788 (N_8788,N_5235,N_5817);
xnor U8789 (N_8789,N_7120,N_5774);
xor U8790 (N_8790,N_7362,N_7302);
nor U8791 (N_8791,N_6849,N_6382);
nor U8792 (N_8792,N_7178,N_7186);
nor U8793 (N_8793,N_5702,N_6225);
or U8794 (N_8794,N_7370,N_7268);
and U8795 (N_8795,N_5286,N_6370);
nand U8796 (N_8796,N_5730,N_5850);
or U8797 (N_8797,N_6435,N_6803);
nor U8798 (N_8798,N_5697,N_7405);
and U8799 (N_8799,N_5010,N_6757);
nand U8800 (N_8800,N_5259,N_6099);
and U8801 (N_8801,N_6274,N_6995);
xnor U8802 (N_8802,N_7371,N_5106);
and U8803 (N_8803,N_5818,N_6405);
nor U8804 (N_8804,N_5489,N_7117);
nand U8805 (N_8805,N_5628,N_6940);
and U8806 (N_8806,N_5204,N_7012);
or U8807 (N_8807,N_6389,N_5406);
and U8808 (N_8808,N_5147,N_5179);
or U8809 (N_8809,N_5706,N_6669);
or U8810 (N_8810,N_6516,N_5267);
nand U8811 (N_8811,N_5941,N_5153);
and U8812 (N_8812,N_6385,N_6036);
nor U8813 (N_8813,N_6803,N_6613);
or U8814 (N_8814,N_6678,N_5481);
nor U8815 (N_8815,N_7296,N_6562);
or U8816 (N_8816,N_5381,N_6130);
or U8817 (N_8817,N_5802,N_5366);
nor U8818 (N_8818,N_6453,N_7396);
or U8819 (N_8819,N_6145,N_6606);
nor U8820 (N_8820,N_7495,N_5214);
nor U8821 (N_8821,N_5267,N_6504);
and U8822 (N_8822,N_6541,N_7233);
xnor U8823 (N_8823,N_5592,N_7140);
nor U8824 (N_8824,N_6567,N_5140);
nand U8825 (N_8825,N_7342,N_6383);
and U8826 (N_8826,N_5398,N_6840);
nand U8827 (N_8827,N_6286,N_5568);
nor U8828 (N_8828,N_5844,N_6722);
and U8829 (N_8829,N_5452,N_7423);
or U8830 (N_8830,N_7311,N_6911);
nor U8831 (N_8831,N_6782,N_5900);
and U8832 (N_8832,N_5062,N_7016);
or U8833 (N_8833,N_6360,N_7057);
and U8834 (N_8834,N_6785,N_7084);
nor U8835 (N_8835,N_6711,N_6919);
nand U8836 (N_8836,N_5636,N_6863);
or U8837 (N_8837,N_5060,N_5240);
or U8838 (N_8838,N_5545,N_5425);
xor U8839 (N_8839,N_5825,N_5513);
nand U8840 (N_8840,N_7145,N_5803);
nand U8841 (N_8841,N_6761,N_7072);
nor U8842 (N_8842,N_6573,N_5617);
and U8843 (N_8843,N_6223,N_7471);
nor U8844 (N_8844,N_6388,N_5667);
or U8845 (N_8845,N_6631,N_6448);
nor U8846 (N_8846,N_6117,N_6537);
nand U8847 (N_8847,N_6762,N_6633);
nor U8848 (N_8848,N_6793,N_7310);
and U8849 (N_8849,N_6336,N_6192);
or U8850 (N_8850,N_5931,N_5696);
or U8851 (N_8851,N_5383,N_6164);
nor U8852 (N_8852,N_6649,N_6113);
and U8853 (N_8853,N_5064,N_7107);
nor U8854 (N_8854,N_7260,N_6182);
nor U8855 (N_8855,N_6345,N_6538);
nor U8856 (N_8856,N_5284,N_5131);
nor U8857 (N_8857,N_7138,N_5715);
xnor U8858 (N_8858,N_6508,N_6662);
or U8859 (N_8859,N_6382,N_5712);
and U8860 (N_8860,N_5612,N_5034);
nand U8861 (N_8861,N_5496,N_7407);
or U8862 (N_8862,N_5677,N_5940);
nor U8863 (N_8863,N_6971,N_7440);
and U8864 (N_8864,N_6914,N_7451);
and U8865 (N_8865,N_6606,N_6585);
nand U8866 (N_8866,N_6736,N_6564);
or U8867 (N_8867,N_7159,N_7033);
nor U8868 (N_8868,N_5278,N_7346);
nand U8869 (N_8869,N_6483,N_5473);
or U8870 (N_8870,N_5509,N_5008);
nand U8871 (N_8871,N_7476,N_5867);
nand U8872 (N_8872,N_6663,N_5712);
or U8873 (N_8873,N_6018,N_5846);
nor U8874 (N_8874,N_6550,N_6299);
and U8875 (N_8875,N_6468,N_6251);
nand U8876 (N_8876,N_7059,N_6881);
nand U8877 (N_8877,N_7279,N_5718);
and U8878 (N_8878,N_5353,N_5262);
nor U8879 (N_8879,N_6343,N_5866);
and U8880 (N_8880,N_6256,N_5604);
or U8881 (N_8881,N_6889,N_6494);
or U8882 (N_8882,N_5562,N_6500);
and U8883 (N_8883,N_7475,N_5669);
nor U8884 (N_8884,N_6713,N_7186);
and U8885 (N_8885,N_5862,N_5428);
or U8886 (N_8886,N_6421,N_6892);
and U8887 (N_8887,N_7235,N_6698);
or U8888 (N_8888,N_5137,N_6762);
or U8889 (N_8889,N_6422,N_6906);
or U8890 (N_8890,N_5384,N_6560);
or U8891 (N_8891,N_5910,N_5831);
or U8892 (N_8892,N_6808,N_6642);
nor U8893 (N_8893,N_6957,N_7213);
nand U8894 (N_8894,N_6270,N_6418);
or U8895 (N_8895,N_5875,N_6116);
or U8896 (N_8896,N_6452,N_5298);
nor U8897 (N_8897,N_5684,N_6943);
nand U8898 (N_8898,N_6746,N_6738);
nand U8899 (N_8899,N_5717,N_6253);
nor U8900 (N_8900,N_6068,N_7005);
or U8901 (N_8901,N_6058,N_5559);
nand U8902 (N_8902,N_7050,N_6531);
and U8903 (N_8903,N_5195,N_6454);
or U8904 (N_8904,N_6730,N_5798);
and U8905 (N_8905,N_6071,N_5975);
nor U8906 (N_8906,N_5051,N_6638);
or U8907 (N_8907,N_5508,N_5093);
nand U8908 (N_8908,N_7434,N_6284);
and U8909 (N_8909,N_6818,N_7426);
nor U8910 (N_8910,N_7494,N_7079);
nand U8911 (N_8911,N_6828,N_5467);
or U8912 (N_8912,N_5634,N_5272);
or U8913 (N_8913,N_7199,N_5775);
nor U8914 (N_8914,N_6593,N_7144);
or U8915 (N_8915,N_5160,N_5225);
or U8916 (N_8916,N_5339,N_7256);
nor U8917 (N_8917,N_7108,N_6270);
nor U8918 (N_8918,N_5627,N_5942);
nor U8919 (N_8919,N_5458,N_6020);
nor U8920 (N_8920,N_5263,N_7047);
xnor U8921 (N_8921,N_7477,N_6295);
nand U8922 (N_8922,N_5273,N_6136);
or U8923 (N_8923,N_5076,N_5489);
and U8924 (N_8924,N_5881,N_5799);
and U8925 (N_8925,N_6851,N_7138);
nand U8926 (N_8926,N_6085,N_5469);
or U8927 (N_8927,N_5928,N_7298);
nor U8928 (N_8928,N_6326,N_5845);
and U8929 (N_8929,N_6489,N_6180);
nand U8930 (N_8930,N_7384,N_6417);
nor U8931 (N_8931,N_5227,N_5016);
xnor U8932 (N_8932,N_6250,N_5640);
nand U8933 (N_8933,N_6542,N_5515);
or U8934 (N_8934,N_5063,N_6189);
nor U8935 (N_8935,N_7272,N_5706);
and U8936 (N_8936,N_6211,N_5541);
nand U8937 (N_8937,N_6254,N_6341);
or U8938 (N_8938,N_7009,N_5948);
and U8939 (N_8939,N_5435,N_7039);
and U8940 (N_8940,N_6159,N_7073);
nand U8941 (N_8941,N_5694,N_6971);
nor U8942 (N_8942,N_5372,N_5374);
nor U8943 (N_8943,N_7444,N_7092);
nand U8944 (N_8944,N_6342,N_6412);
or U8945 (N_8945,N_6722,N_5416);
nor U8946 (N_8946,N_6799,N_6028);
nand U8947 (N_8947,N_7299,N_5333);
or U8948 (N_8948,N_5733,N_6308);
nand U8949 (N_8949,N_6679,N_7175);
and U8950 (N_8950,N_5685,N_7230);
and U8951 (N_8951,N_6403,N_6877);
nor U8952 (N_8952,N_7028,N_5420);
or U8953 (N_8953,N_7228,N_5906);
nor U8954 (N_8954,N_5030,N_5735);
nand U8955 (N_8955,N_7224,N_6865);
nand U8956 (N_8956,N_7495,N_6464);
and U8957 (N_8957,N_6827,N_6571);
nand U8958 (N_8958,N_6441,N_7421);
or U8959 (N_8959,N_6787,N_5501);
and U8960 (N_8960,N_5760,N_6120);
nand U8961 (N_8961,N_5659,N_7024);
nand U8962 (N_8962,N_6486,N_7032);
and U8963 (N_8963,N_5676,N_6517);
or U8964 (N_8964,N_5331,N_6845);
and U8965 (N_8965,N_5533,N_7250);
and U8966 (N_8966,N_5246,N_5759);
nand U8967 (N_8967,N_6383,N_5933);
nor U8968 (N_8968,N_6607,N_5568);
nand U8969 (N_8969,N_6590,N_6770);
xnor U8970 (N_8970,N_5275,N_6185);
nor U8971 (N_8971,N_7157,N_6224);
or U8972 (N_8972,N_7217,N_5480);
and U8973 (N_8973,N_5500,N_5797);
nand U8974 (N_8974,N_5836,N_5134);
and U8975 (N_8975,N_7431,N_5651);
xnor U8976 (N_8976,N_5362,N_6697);
nor U8977 (N_8977,N_7311,N_5361);
nand U8978 (N_8978,N_6367,N_5550);
or U8979 (N_8979,N_6678,N_7258);
or U8980 (N_8980,N_7228,N_6882);
and U8981 (N_8981,N_5210,N_5243);
and U8982 (N_8982,N_7204,N_6664);
nand U8983 (N_8983,N_5244,N_5298);
or U8984 (N_8984,N_5308,N_5803);
nor U8985 (N_8985,N_6783,N_6340);
nor U8986 (N_8986,N_7218,N_5521);
or U8987 (N_8987,N_5280,N_6895);
nand U8988 (N_8988,N_6776,N_6775);
nand U8989 (N_8989,N_7071,N_5385);
nand U8990 (N_8990,N_5714,N_5220);
nor U8991 (N_8991,N_5727,N_7189);
nor U8992 (N_8992,N_5582,N_7032);
xor U8993 (N_8993,N_6113,N_6375);
nor U8994 (N_8994,N_6504,N_6728);
nor U8995 (N_8995,N_6065,N_6924);
and U8996 (N_8996,N_5203,N_7286);
and U8997 (N_8997,N_5854,N_7032);
and U8998 (N_8998,N_6441,N_5552);
or U8999 (N_8999,N_5286,N_6389);
nor U9000 (N_9000,N_6687,N_7204);
or U9001 (N_9001,N_6040,N_5434);
and U9002 (N_9002,N_6724,N_5670);
or U9003 (N_9003,N_5057,N_6391);
or U9004 (N_9004,N_5415,N_7218);
or U9005 (N_9005,N_5122,N_5996);
or U9006 (N_9006,N_5131,N_6418);
and U9007 (N_9007,N_5777,N_5601);
nand U9008 (N_9008,N_5836,N_6824);
or U9009 (N_9009,N_5203,N_6634);
nand U9010 (N_9010,N_7058,N_5045);
nand U9011 (N_9011,N_5177,N_6500);
and U9012 (N_9012,N_5432,N_6444);
nand U9013 (N_9013,N_5384,N_5237);
nor U9014 (N_9014,N_6611,N_6647);
and U9015 (N_9015,N_5743,N_5666);
and U9016 (N_9016,N_5000,N_5263);
nor U9017 (N_9017,N_5758,N_5630);
and U9018 (N_9018,N_5910,N_6267);
nand U9019 (N_9019,N_5481,N_7492);
nand U9020 (N_9020,N_5272,N_5436);
and U9021 (N_9021,N_6821,N_5053);
nand U9022 (N_9022,N_6601,N_7372);
or U9023 (N_9023,N_7071,N_5702);
and U9024 (N_9024,N_7124,N_5957);
or U9025 (N_9025,N_6105,N_5129);
nor U9026 (N_9026,N_6631,N_5610);
nor U9027 (N_9027,N_6126,N_5152);
or U9028 (N_9028,N_5526,N_6626);
and U9029 (N_9029,N_7356,N_6994);
nor U9030 (N_9030,N_7038,N_7004);
xor U9031 (N_9031,N_7468,N_7166);
nor U9032 (N_9032,N_6252,N_5405);
nand U9033 (N_9033,N_5680,N_5229);
nor U9034 (N_9034,N_6644,N_5505);
nand U9035 (N_9035,N_6617,N_7451);
xnor U9036 (N_9036,N_5631,N_6074);
nand U9037 (N_9037,N_5059,N_5614);
nand U9038 (N_9038,N_5042,N_7148);
and U9039 (N_9039,N_7446,N_6410);
or U9040 (N_9040,N_6777,N_6875);
nand U9041 (N_9041,N_5577,N_5144);
nor U9042 (N_9042,N_6515,N_6781);
xor U9043 (N_9043,N_5362,N_7125);
nor U9044 (N_9044,N_7402,N_6942);
and U9045 (N_9045,N_7148,N_5012);
nor U9046 (N_9046,N_6243,N_7190);
and U9047 (N_9047,N_7395,N_7490);
nor U9048 (N_9048,N_5863,N_6221);
and U9049 (N_9049,N_5641,N_7359);
xnor U9050 (N_9050,N_5505,N_6425);
or U9051 (N_9051,N_6350,N_7156);
nor U9052 (N_9052,N_6132,N_7343);
and U9053 (N_9053,N_6729,N_6579);
nor U9054 (N_9054,N_7361,N_5521);
or U9055 (N_9055,N_7191,N_6405);
nand U9056 (N_9056,N_6054,N_6601);
nand U9057 (N_9057,N_5957,N_5687);
and U9058 (N_9058,N_5126,N_5356);
nor U9059 (N_9059,N_7135,N_5861);
or U9060 (N_9060,N_5871,N_5647);
and U9061 (N_9061,N_6075,N_5061);
nor U9062 (N_9062,N_6053,N_6202);
nor U9063 (N_9063,N_6688,N_6154);
nand U9064 (N_9064,N_7256,N_5919);
and U9065 (N_9065,N_5054,N_7442);
nor U9066 (N_9066,N_5551,N_6817);
and U9067 (N_9067,N_5086,N_7079);
nor U9068 (N_9068,N_7155,N_5031);
nand U9069 (N_9069,N_5441,N_5014);
and U9070 (N_9070,N_5572,N_6970);
or U9071 (N_9071,N_6069,N_6014);
or U9072 (N_9072,N_6566,N_7331);
and U9073 (N_9073,N_7281,N_7448);
or U9074 (N_9074,N_5133,N_6288);
nand U9075 (N_9075,N_6187,N_5929);
and U9076 (N_9076,N_7461,N_5268);
or U9077 (N_9077,N_7191,N_7342);
or U9078 (N_9078,N_5874,N_7202);
nand U9079 (N_9079,N_5512,N_6628);
nand U9080 (N_9080,N_6599,N_5145);
or U9081 (N_9081,N_6974,N_5528);
nor U9082 (N_9082,N_6874,N_6269);
or U9083 (N_9083,N_6518,N_5204);
nand U9084 (N_9084,N_7381,N_5279);
and U9085 (N_9085,N_5785,N_5134);
nand U9086 (N_9086,N_6495,N_5688);
nand U9087 (N_9087,N_6821,N_7233);
and U9088 (N_9088,N_5203,N_5057);
nor U9089 (N_9089,N_7071,N_5656);
nor U9090 (N_9090,N_6669,N_6498);
or U9091 (N_9091,N_7282,N_5238);
nand U9092 (N_9092,N_6436,N_6961);
nor U9093 (N_9093,N_7026,N_7143);
nand U9094 (N_9094,N_5575,N_7223);
nand U9095 (N_9095,N_7108,N_5796);
or U9096 (N_9096,N_5566,N_5406);
and U9097 (N_9097,N_5281,N_7105);
and U9098 (N_9098,N_6952,N_5696);
nor U9099 (N_9099,N_7332,N_5197);
and U9100 (N_9100,N_7037,N_7181);
or U9101 (N_9101,N_5488,N_7352);
or U9102 (N_9102,N_5441,N_6009);
xnor U9103 (N_9103,N_7251,N_5848);
or U9104 (N_9104,N_7422,N_5582);
nor U9105 (N_9105,N_6995,N_6456);
nor U9106 (N_9106,N_6785,N_6714);
nand U9107 (N_9107,N_7117,N_5633);
nand U9108 (N_9108,N_6788,N_6177);
xor U9109 (N_9109,N_5126,N_6303);
nand U9110 (N_9110,N_6769,N_6307);
nor U9111 (N_9111,N_5004,N_6157);
nor U9112 (N_9112,N_5554,N_6360);
nand U9113 (N_9113,N_5682,N_7047);
and U9114 (N_9114,N_5964,N_6106);
or U9115 (N_9115,N_6517,N_6259);
nor U9116 (N_9116,N_5840,N_5731);
nand U9117 (N_9117,N_6172,N_6029);
nor U9118 (N_9118,N_5762,N_7317);
or U9119 (N_9119,N_5698,N_6274);
nor U9120 (N_9120,N_5978,N_6706);
and U9121 (N_9121,N_6660,N_5474);
or U9122 (N_9122,N_6759,N_7460);
nand U9123 (N_9123,N_5850,N_6648);
or U9124 (N_9124,N_5195,N_6515);
nand U9125 (N_9125,N_6108,N_5444);
and U9126 (N_9126,N_6299,N_6077);
nand U9127 (N_9127,N_6971,N_7375);
nand U9128 (N_9128,N_6373,N_7031);
or U9129 (N_9129,N_6257,N_7395);
and U9130 (N_9130,N_5208,N_5525);
and U9131 (N_9131,N_5052,N_6196);
and U9132 (N_9132,N_6906,N_6908);
nand U9133 (N_9133,N_5165,N_5030);
or U9134 (N_9134,N_6022,N_6272);
and U9135 (N_9135,N_5380,N_5844);
nand U9136 (N_9136,N_5777,N_6705);
nor U9137 (N_9137,N_7219,N_5728);
and U9138 (N_9138,N_5151,N_7386);
and U9139 (N_9139,N_5976,N_5146);
or U9140 (N_9140,N_5831,N_7001);
nand U9141 (N_9141,N_5420,N_5850);
nor U9142 (N_9142,N_6255,N_5786);
nand U9143 (N_9143,N_5808,N_5947);
nor U9144 (N_9144,N_5960,N_5008);
nor U9145 (N_9145,N_7339,N_6992);
nand U9146 (N_9146,N_7246,N_5060);
and U9147 (N_9147,N_6896,N_6596);
or U9148 (N_9148,N_6756,N_6659);
nor U9149 (N_9149,N_5150,N_6740);
or U9150 (N_9150,N_6922,N_6967);
and U9151 (N_9151,N_6705,N_6713);
or U9152 (N_9152,N_7243,N_7275);
and U9153 (N_9153,N_6085,N_7177);
nor U9154 (N_9154,N_6528,N_7349);
nand U9155 (N_9155,N_6524,N_5554);
nand U9156 (N_9156,N_5334,N_6960);
or U9157 (N_9157,N_5725,N_6977);
nand U9158 (N_9158,N_7273,N_6349);
nand U9159 (N_9159,N_5976,N_6550);
xor U9160 (N_9160,N_5861,N_7439);
nor U9161 (N_9161,N_6214,N_5243);
nor U9162 (N_9162,N_7343,N_5015);
nand U9163 (N_9163,N_7359,N_7000);
nor U9164 (N_9164,N_7241,N_5563);
or U9165 (N_9165,N_7296,N_6596);
nand U9166 (N_9166,N_5575,N_5998);
nand U9167 (N_9167,N_5913,N_7018);
or U9168 (N_9168,N_7243,N_6693);
nor U9169 (N_9169,N_5389,N_6303);
nor U9170 (N_9170,N_7481,N_7459);
or U9171 (N_9171,N_6312,N_5226);
nand U9172 (N_9172,N_5473,N_6991);
and U9173 (N_9173,N_5794,N_7127);
and U9174 (N_9174,N_5771,N_5712);
nand U9175 (N_9175,N_5456,N_7477);
nand U9176 (N_9176,N_7249,N_6104);
and U9177 (N_9177,N_6164,N_5150);
and U9178 (N_9178,N_5525,N_5032);
xnor U9179 (N_9179,N_6931,N_5184);
and U9180 (N_9180,N_6142,N_6318);
or U9181 (N_9181,N_6210,N_5531);
and U9182 (N_9182,N_7356,N_6419);
and U9183 (N_9183,N_6211,N_5152);
and U9184 (N_9184,N_6391,N_5708);
and U9185 (N_9185,N_6928,N_5232);
and U9186 (N_9186,N_6191,N_5569);
and U9187 (N_9187,N_5049,N_5548);
and U9188 (N_9188,N_7295,N_6105);
and U9189 (N_9189,N_6185,N_5005);
and U9190 (N_9190,N_6219,N_6106);
and U9191 (N_9191,N_5177,N_6968);
nor U9192 (N_9192,N_6357,N_6162);
or U9193 (N_9193,N_7480,N_5814);
nor U9194 (N_9194,N_5209,N_6248);
and U9195 (N_9195,N_7318,N_7334);
nor U9196 (N_9196,N_5822,N_5565);
nand U9197 (N_9197,N_6393,N_6780);
and U9198 (N_9198,N_6390,N_5800);
or U9199 (N_9199,N_7191,N_5284);
nand U9200 (N_9200,N_5734,N_6867);
nor U9201 (N_9201,N_5224,N_5396);
nor U9202 (N_9202,N_6650,N_7438);
nand U9203 (N_9203,N_6940,N_5621);
and U9204 (N_9204,N_5560,N_5186);
nand U9205 (N_9205,N_6488,N_7060);
and U9206 (N_9206,N_5655,N_5264);
nand U9207 (N_9207,N_6060,N_6336);
nand U9208 (N_9208,N_6516,N_6608);
nand U9209 (N_9209,N_5969,N_6596);
nand U9210 (N_9210,N_6652,N_5156);
nor U9211 (N_9211,N_7042,N_5692);
nand U9212 (N_9212,N_6447,N_7495);
or U9213 (N_9213,N_7133,N_6360);
and U9214 (N_9214,N_5676,N_7197);
nor U9215 (N_9215,N_5150,N_5879);
nor U9216 (N_9216,N_6204,N_6405);
nor U9217 (N_9217,N_5270,N_5945);
and U9218 (N_9218,N_5407,N_6049);
nand U9219 (N_9219,N_5685,N_5083);
nand U9220 (N_9220,N_7380,N_5153);
or U9221 (N_9221,N_7476,N_5695);
nor U9222 (N_9222,N_5216,N_5131);
nor U9223 (N_9223,N_5266,N_5165);
and U9224 (N_9224,N_5148,N_5510);
and U9225 (N_9225,N_6281,N_5320);
nor U9226 (N_9226,N_5592,N_5356);
nand U9227 (N_9227,N_6508,N_6434);
or U9228 (N_9228,N_6927,N_7316);
or U9229 (N_9229,N_6875,N_5633);
nand U9230 (N_9230,N_7446,N_6755);
or U9231 (N_9231,N_7360,N_7359);
and U9232 (N_9232,N_6794,N_7216);
and U9233 (N_9233,N_5781,N_5816);
nor U9234 (N_9234,N_6349,N_6799);
or U9235 (N_9235,N_5069,N_5850);
nand U9236 (N_9236,N_6855,N_6994);
xor U9237 (N_9237,N_6488,N_6285);
or U9238 (N_9238,N_6402,N_5552);
or U9239 (N_9239,N_5029,N_6814);
or U9240 (N_9240,N_5460,N_5755);
or U9241 (N_9241,N_5857,N_7080);
and U9242 (N_9242,N_6607,N_6531);
nand U9243 (N_9243,N_6188,N_7055);
nor U9244 (N_9244,N_6548,N_5902);
and U9245 (N_9245,N_7005,N_6277);
or U9246 (N_9246,N_7480,N_6882);
and U9247 (N_9247,N_6725,N_6479);
and U9248 (N_9248,N_7153,N_6393);
nand U9249 (N_9249,N_5542,N_6474);
nor U9250 (N_9250,N_5234,N_6109);
or U9251 (N_9251,N_7003,N_7026);
or U9252 (N_9252,N_6296,N_6752);
nand U9253 (N_9253,N_7426,N_5849);
nand U9254 (N_9254,N_6558,N_6655);
and U9255 (N_9255,N_5495,N_7337);
or U9256 (N_9256,N_6557,N_6964);
or U9257 (N_9257,N_5269,N_6292);
and U9258 (N_9258,N_6012,N_6042);
and U9259 (N_9259,N_7270,N_5915);
and U9260 (N_9260,N_6010,N_5447);
nor U9261 (N_9261,N_7490,N_6457);
nor U9262 (N_9262,N_5134,N_7065);
nor U9263 (N_9263,N_6855,N_5790);
or U9264 (N_9264,N_6834,N_6059);
nand U9265 (N_9265,N_5586,N_6870);
nor U9266 (N_9266,N_5279,N_6053);
xnor U9267 (N_9267,N_5919,N_7184);
and U9268 (N_9268,N_7136,N_6026);
and U9269 (N_9269,N_6470,N_7114);
or U9270 (N_9270,N_6721,N_7113);
or U9271 (N_9271,N_6931,N_5152);
or U9272 (N_9272,N_6057,N_6370);
nand U9273 (N_9273,N_6302,N_6161);
nor U9274 (N_9274,N_6476,N_6387);
nor U9275 (N_9275,N_5153,N_5015);
nand U9276 (N_9276,N_6722,N_5342);
nand U9277 (N_9277,N_7461,N_5587);
and U9278 (N_9278,N_6280,N_6230);
or U9279 (N_9279,N_6217,N_6772);
and U9280 (N_9280,N_7358,N_6314);
or U9281 (N_9281,N_6753,N_6081);
and U9282 (N_9282,N_5031,N_5439);
nand U9283 (N_9283,N_5630,N_7304);
and U9284 (N_9284,N_6714,N_5701);
nor U9285 (N_9285,N_5914,N_5726);
or U9286 (N_9286,N_6383,N_5595);
nand U9287 (N_9287,N_6850,N_6916);
or U9288 (N_9288,N_5062,N_6716);
xor U9289 (N_9289,N_5681,N_7295);
xnor U9290 (N_9290,N_6520,N_6984);
or U9291 (N_9291,N_6596,N_7409);
nor U9292 (N_9292,N_5808,N_6297);
nand U9293 (N_9293,N_5076,N_6783);
or U9294 (N_9294,N_5001,N_6131);
and U9295 (N_9295,N_5530,N_6483);
and U9296 (N_9296,N_6137,N_6980);
xnor U9297 (N_9297,N_7172,N_5831);
nor U9298 (N_9298,N_6098,N_6113);
or U9299 (N_9299,N_5255,N_7162);
and U9300 (N_9300,N_6293,N_5726);
or U9301 (N_9301,N_6045,N_6618);
and U9302 (N_9302,N_5898,N_6352);
nand U9303 (N_9303,N_6689,N_5558);
nand U9304 (N_9304,N_6339,N_6503);
and U9305 (N_9305,N_6323,N_7046);
and U9306 (N_9306,N_6566,N_6231);
and U9307 (N_9307,N_6567,N_5885);
nand U9308 (N_9308,N_6789,N_6656);
nor U9309 (N_9309,N_6339,N_6078);
nor U9310 (N_9310,N_6457,N_6011);
and U9311 (N_9311,N_6799,N_5502);
and U9312 (N_9312,N_6993,N_6027);
nand U9313 (N_9313,N_7258,N_7421);
nor U9314 (N_9314,N_7258,N_6452);
nand U9315 (N_9315,N_5853,N_7259);
or U9316 (N_9316,N_6887,N_5056);
and U9317 (N_9317,N_7436,N_6393);
nand U9318 (N_9318,N_5291,N_6795);
nor U9319 (N_9319,N_6665,N_7407);
or U9320 (N_9320,N_6480,N_5020);
and U9321 (N_9321,N_6322,N_6768);
and U9322 (N_9322,N_5248,N_6715);
nand U9323 (N_9323,N_5377,N_5205);
and U9324 (N_9324,N_6711,N_6039);
or U9325 (N_9325,N_5476,N_6325);
nor U9326 (N_9326,N_6899,N_7438);
nor U9327 (N_9327,N_6710,N_6506);
nor U9328 (N_9328,N_5284,N_6900);
and U9329 (N_9329,N_5988,N_5234);
or U9330 (N_9330,N_7309,N_7361);
nand U9331 (N_9331,N_6110,N_5148);
and U9332 (N_9332,N_6425,N_5426);
nor U9333 (N_9333,N_5100,N_6361);
nor U9334 (N_9334,N_7126,N_7010);
nor U9335 (N_9335,N_6986,N_5787);
and U9336 (N_9336,N_5999,N_7152);
and U9337 (N_9337,N_6612,N_6751);
nand U9338 (N_9338,N_5479,N_6862);
and U9339 (N_9339,N_7133,N_5044);
or U9340 (N_9340,N_6194,N_7025);
nor U9341 (N_9341,N_5957,N_6027);
nor U9342 (N_9342,N_7021,N_6568);
nand U9343 (N_9343,N_5211,N_7342);
or U9344 (N_9344,N_5640,N_5553);
or U9345 (N_9345,N_5749,N_5540);
or U9346 (N_9346,N_6823,N_5747);
nand U9347 (N_9347,N_5553,N_5907);
nand U9348 (N_9348,N_5631,N_7410);
nand U9349 (N_9349,N_6709,N_5595);
nor U9350 (N_9350,N_7241,N_6462);
nand U9351 (N_9351,N_5973,N_6569);
or U9352 (N_9352,N_5030,N_7328);
nand U9353 (N_9353,N_5952,N_5634);
and U9354 (N_9354,N_6865,N_6668);
and U9355 (N_9355,N_5295,N_6985);
nand U9356 (N_9356,N_6092,N_5959);
and U9357 (N_9357,N_7192,N_5053);
or U9358 (N_9358,N_6033,N_7211);
or U9359 (N_9359,N_5701,N_7461);
nand U9360 (N_9360,N_6470,N_5123);
or U9361 (N_9361,N_5639,N_7051);
nand U9362 (N_9362,N_5613,N_5464);
nor U9363 (N_9363,N_6920,N_7034);
nand U9364 (N_9364,N_6320,N_5818);
and U9365 (N_9365,N_5337,N_5771);
or U9366 (N_9366,N_6135,N_6859);
and U9367 (N_9367,N_7221,N_6417);
xor U9368 (N_9368,N_5341,N_5119);
or U9369 (N_9369,N_6124,N_7117);
or U9370 (N_9370,N_5011,N_5377);
or U9371 (N_9371,N_6091,N_6877);
or U9372 (N_9372,N_5011,N_5280);
nand U9373 (N_9373,N_7198,N_6557);
nor U9374 (N_9374,N_6142,N_7253);
xnor U9375 (N_9375,N_6314,N_7050);
and U9376 (N_9376,N_5075,N_5489);
and U9377 (N_9377,N_5246,N_5548);
and U9378 (N_9378,N_6551,N_5861);
nor U9379 (N_9379,N_6061,N_5597);
nand U9380 (N_9380,N_7228,N_5120);
nor U9381 (N_9381,N_5937,N_6003);
or U9382 (N_9382,N_5520,N_5325);
nor U9383 (N_9383,N_6261,N_7441);
nor U9384 (N_9384,N_5772,N_5981);
nand U9385 (N_9385,N_6800,N_5365);
nand U9386 (N_9386,N_5087,N_6428);
and U9387 (N_9387,N_6774,N_6500);
or U9388 (N_9388,N_5662,N_6367);
and U9389 (N_9389,N_6251,N_6709);
nor U9390 (N_9390,N_6411,N_5989);
or U9391 (N_9391,N_6751,N_6355);
and U9392 (N_9392,N_6682,N_6182);
or U9393 (N_9393,N_6586,N_6298);
or U9394 (N_9394,N_6881,N_7188);
or U9395 (N_9395,N_6580,N_7165);
nor U9396 (N_9396,N_5725,N_7040);
or U9397 (N_9397,N_5412,N_5660);
nor U9398 (N_9398,N_5466,N_7270);
nor U9399 (N_9399,N_5434,N_6601);
nor U9400 (N_9400,N_7077,N_5438);
and U9401 (N_9401,N_7457,N_5515);
or U9402 (N_9402,N_5717,N_6843);
or U9403 (N_9403,N_5757,N_7493);
nor U9404 (N_9404,N_5422,N_5321);
or U9405 (N_9405,N_6660,N_6562);
nor U9406 (N_9406,N_5613,N_7321);
nand U9407 (N_9407,N_5704,N_7194);
nand U9408 (N_9408,N_6836,N_5763);
nor U9409 (N_9409,N_7161,N_7369);
nor U9410 (N_9410,N_5952,N_6056);
nand U9411 (N_9411,N_6360,N_6681);
xnor U9412 (N_9412,N_5743,N_6171);
and U9413 (N_9413,N_6302,N_7185);
and U9414 (N_9414,N_5368,N_5302);
nor U9415 (N_9415,N_6023,N_7007);
nor U9416 (N_9416,N_5382,N_5165);
nor U9417 (N_9417,N_5094,N_5341);
or U9418 (N_9418,N_5537,N_5911);
or U9419 (N_9419,N_6398,N_5556);
nand U9420 (N_9420,N_7264,N_5086);
or U9421 (N_9421,N_7429,N_6083);
nor U9422 (N_9422,N_5295,N_5562);
nand U9423 (N_9423,N_5476,N_7478);
and U9424 (N_9424,N_7149,N_7407);
and U9425 (N_9425,N_7188,N_5730);
nand U9426 (N_9426,N_7110,N_5923);
or U9427 (N_9427,N_6485,N_6828);
xor U9428 (N_9428,N_5692,N_7440);
and U9429 (N_9429,N_6645,N_5153);
nand U9430 (N_9430,N_7110,N_5134);
and U9431 (N_9431,N_6084,N_7134);
and U9432 (N_9432,N_6247,N_7415);
nor U9433 (N_9433,N_7126,N_5161);
or U9434 (N_9434,N_5664,N_6887);
nor U9435 (N_9435,N_5447,N_6417);
nand U9436 (N_9436,N_5517,N_5379);
or U9437 (N_9437,N_6783,N_7076);
and U9438 (N_9438,N_7177,N_5848);
nand U9439 (N_9439,N_7308,N_6408);
or U9440 (N_9440,N_7054,N_6630);
nand U9441 (N_9441,N_6136,N_6489);
nand U9442 (N_9442,N_7479,N_7206);
nand U9443 (N_9443,N_6867,N_6587);
nor U9444 (N_9444,N_7280,N_6839);
xnor U9445 (N_9445,N_5516,N_5601);
and U9446 (N_9446,N_7409,N_5528);
or U9447 (N_9447,N_7205,N_5219);
nand U9448 (N_9448,N_7112,N_7236);
or U9449 (N_9449,N_6506,N_5443);
and U9450 (N_9450,N_6508,N_6952);
and U9451 (N_9451,N_7357,N_5743);
nor U9452 (N_9452,N_7075,N_7082);
or U9453 (N_9453,N_7204,N_6287);
or U9454 (N_9454,N_7281,N_6152);
nor U9455 (N_9455,N_5535,N_5500);
nor U9456 (N_9456,N_7146,N_6807);
nand U9457 (N_9457,N_6153,N_6841);
nand U9458 (N_9458,N_5542,N_6742);
nor U9459 (N_9459,N_5701,N_5758);
and U9460 (N_9460,N_6876,N_6874);
or U9461 (N_9461,N_6871,N_5705);
and U9462 (N_9462,N_5949,N_7026);
and U9463 (N_9463,N_5683,N_5872);
nand U9464 (N_9464,N_7313,N_6021);
nor U9465 (N_9465,N_5110,N_5760);
nor U9466 (N_9466,N_6785,N_6170);
nor U9467 (N_9467,N_6008,N_6862);
nor U9468 (N_9468,N_6372,N_7475);
nor U9469 (N_9469,N_6381,N_6549);
or U9470 (N_9470,N_6521,N_6010);
or U9471 (N_9471,N_5118,N_5993);
or U9472 (N_9472,N_7490,N_6340);
and U9473 (N_9473,N_5266,N_5622);
nand U9474 (N_9474,N_6726,N_5466);
or U9475 (N_9475,N_7028,N_6502);
nor U9476 (N_9476,N_5704,N_6623);
or U9477 (N_9477,N_5588,N_5323);
nor U9478 (N_9478,N_5066,N_6534);
or U9479 (N_9479,N_7001,N_7399);
nor U9480 (N_9480,N_7348,N_6155);
or U9481 (N_9481,N_5607,N_5928);
xor U9482 (N_9482,N_5318,N_7041);
nand U9483 (N_9483,N_5977,N_6650);
xnor U9484 (N_9484,N_5103,N_6441);
and U9485 (N_9485,N_5072,N_6493);
nand U9486 (N_9486,N_5455,N_5650);
and U9487 (N_9487,N_5719,N_7190);
or U9488 (N_9488,N_5132,N_7035);
xnor U9489 (N_9489,N_6642,N_5479);
and U9490 (N_9490,N_5565,N_7289);
and U9491 (N_9491,N_5861,N_6446);
or U9492 (N_9492,N_5234,N_6502);
or U9493 (N_9493,N_5603,N_5417);
and U9494 (N_9494,N_7372,N_7115);
nor U9495 (N_9495,N_6310,N_5840);
nand U9496 (N_9496,N_7385,N_7140);
and U9497 (N_9497,N_6579,N_7392);
or U9498 (N_9498,N_6979,N_6011);
nor U9499 (N_9499,N_5245,N_7367);
nor U9500 (N_9500,N_6014,N_5090);
xnor U9501 (N_9501,N_7123,N_6536);
or U9502 (N_9502,N_7424,N_6019);
nor U9503 (N_9503,N_7121,N_5250);
nand U9504 (N_9504,N_6766,N_6307);
nor U9505 (N_9505,N_5960,N_6718);
nor U9506 (N_9506,N_6684,N_7336);
or U9507 (N_9507,N_5350,N_7057);
and U9508 (N_9508,N_6663,N_5969);
nor U9509 (N_9509,N_7430,N_5064);
or U9510 (N_9510,N_5940,N_6768);
nor U9511 (N_9511,N_6700,N_7077);
nand U9512 (N_9512,N_6478,N_5294);
and U9513 (N_9513,N_7053,N_7101);
nand U9514 (N_9514,N_6433,N_6851);
nor U9515 (N_9515,N_6052,N_7069);
and U9516 (N_9516,N_7341,N_7497);
or U9517 (N_9517,N_6393,N_5186);
nor U9518 (N_9518,N_6017,N_5170);
and U9519 (N_9519,N_7449,N_7095);
nor U9520 (N_9520,N_6453,N_7255);
nand U9521 (N_9521,N_5700,N_6680);
nor U9522 (N_9522,N_6656,N_5041);
nand U9523 (N_9523,N_7347,N_5908);
nor U9524 (N_9524,N_5228,N_5397);
nor U9525 (N_9525,N_6997,N_6662);
nand U9526 (N_9526,N_5306,N_7270);
nor U9527 (N_9527,N_7001,N_7111);
and U9528 (N_9528,N_5783,N_6687);
and U9529 (N_9529,N_6580,N_6708);
or U9530 (N_9530,N_7155,N_6250);
or U9531 (N_9531,N_6375,N_6749);
and U9532 (N_9532,N_5488,N_5483);
and U9533 (N_9533,N_7465,N_5748);
and U9534 (N_9534,N_7036,N_6282);
and U9535 (N_9535,N_6317,N_7161);
nand U9536 (N_9536,N_6350,N_6149);
and U9537 (N_9537,N_5072,N_6173);
nor U9538 (N_9538,N_6849,N_6072);
nand U9539 (N_9539,N_5572,N_5881);
nand U9540 (N_9540,N_6263,N_6988);
nand U9541 (N_9541,N_7143,N_6460);
and U9542 (N_9542,N_6203,N_6053);
nor U9543 (N_9543,N_7252,N_5554);
or U9544 (N_9544,N_6552,N_7425);
or U9545 (N_9545,N_5170,N_5811);
and U9546 (N_9546,N_6690,N_5770);
nand U9547 (N_9547,N_5716,N_7120);
nand U9548 (N_9548,N_6880,N_5763);
nor U9549 (N_9549,N_6139,N_5128);
and U9550 (N_9550,N_5961,N_7336);
nor U9551 (N_9551,N_5342,N_5749);
nor U9552 (N_9552,N_6683,N_5389);
and U9553 (N_9553,N_7056,N_7297);
nand U9554 (N_9554,N_6578,N_6135);
or U9555 (N_9555,N_5791,N_6334);
nor U9556 (N_9556,N_7041,N_7277);
or U9557 (N_9557,N_5413,N_5393);
or U9558 (N_9558,N_5786,N_6792);
nor U9559 (N_9559,N_7170,N_6976);
or U9560 (N_9560,N_5860,N_7434);
nand U9561 (N_9561,N_6678,N_6612);
or U9562 (N_9562,N_5540,N_6921);
and U9563 (N_9563,N_5966,N_6392);
nor U9564 (N_9564,N_5967,N_6386);
and U9565 (N_9565,N_5278,N_6108);
xnor U9566 (N_9566,N_5616,N_6703);
and U9567 (N_9567,N_5905,N_6048);
nor U9568 (N_9568,N_6402,N_7104);
nand U9569 (N_9569,N_7213,N_6714);
and U9570 (N_9570,N_5145,N_5857);
nand U9571 (N_9571,N_6088,N_5638);
or U9572 (N_9572,N_7300,N_5150);
nand U9573 (N_9573,N_7124,N_6402);
nor U9574 (N_9574,N_6819,N_6239);
or U9575 (N_9575,N_5468,N_6825);
nor U9576 (N_9576,N_5162,N_6123);
nand U9577 (N_9577,N_7142,N_5970);
nor U9578 (N_9578,N_6737,N_7379);
nor U9579 (N_9579,N_5403,N_5604);
nand U9580 (N_9580,N_6127,N_7019);
nand U9581 (N_9581,N_6206,N_6411);
or U9582 (N_9582,N_6265,N_7218);
or U9583 (N_9583,N_5251,N_6945);
or U9584 (N_9584,N_5138,N_5659);
nor U9585 (N_9585,N_5851,N_6782);
or U9586 (N_9586,N_5434,N_6091);
or U9587 (N_9587,N_5849,N_6957);
nand U9588 (N_9588,N_7203,N_5398);
nand U9589 (N_9589,N_6181,N_7073);
nand U9590 (N_9590,N_6514,N_6201);
or U9591 (N_9591,N_7007,N_5778);
and U9592 (N_9592,N_7232,N_6710);
and U9593 (N_9593,N_5237,N_6087);
nand U9594 (N_9594,N_6221,N_5954);
nor U9595 (N_9595,N_6431,N_7113);
nor U9596 (N_9596,N_6876,N_6985);
and U9597 (N_9597,N_6247,N_6681);
or U9598 (N_9598,N_5649,N_5640);
and U9599 (N_9599,N_6608,N_6089);
and U9600 (N_9600,N_7360,N_5129);
or U9601 (N_9601,N_6597,N_5581);
nor U9602 (N_9602,N_5793,N_5587);
nor U9603 (N_9603,N_6691,N_7241);
and U9604 (N_9604,N_6108,N_7281);
nand U9605 (N_9605,N_5064,N_5561);
or U9606 (N_9606,N_7118,N_6436);
and U9607 (N_9607,N_5302,N_5454);
nor U9608 (N_9608,N_6277,N_5866);
nand U9609 (N_9609,N_5120,N_6450);
nand U9610 (N_9610,N_6429,N_5824);
and U9611 (N_9611,N_6157,N_5897);
or U9612 (N_9612,N_6140,N_5768);
or U9613 (N_9613,N_6132,N_7497);
nand U9614 (N_9614,N_7213,N_7480);
nor U9615 (N_9615,N_6763,N_7440);
or U9616 (N_9616,N_7059,N_7471);
or U9617 (N_9617,N_7007,N_6602);
or U9618 (N_9618,N_5004,N_6884);
and U9619 (N_9619,N_7063,N_6768);
nor U9620 (N_9620,N_6774,N_7465);
or U9621 (N_9621,N_5774,N_5072);
and U9622 (N_9622,N_5286,N_5927);
or U9623 (N_9623,N_5829,N_6686);
nand U9624 (N_9624,N_6764,N_6384);
nand U9625 (N_9625,N_5026,N_5431);
and U9626 (N_9626,N_7079,N_6885);
or U9627 (N_9627,N_5735,N_6566);
and U9628 (N_9628,N_7498,N_6007);
nor U9629 (N_9629,N_6169,N_6746);
nand U9630 (N_9630,N_5173,N_6907);
nor U9631 (N_9631,N_6884,N_6293);
nor U9632 (N_9632,N_5223,N_5026);
and U9633 (N_9633,N_5303,N_6331);
nor U9634 (N_9634,N_7001,N_5365);
xor U9635 (N_9635,N_5952,N_5860);
or U9636 (N_9636,N_5552,N_5368);
nor U9637 (N_9637,N_6208,N_6196);
and U9638 (N_9638,N_5911,N_6390);
nand U9639 (N_9639,N_7307,N_6281);
nand U9640 (N_9640,N_7100,N_6572);
xor U9641 (N_9641,N_5075,N_6197);
nand U9642 (N_9642,N_6754,N_6977);
or U9643 (N_9643,N_5934,N_7076);
nor U9644 (N_9644,N_6419,N_6812);
and U9645 (N_9645,N_5609,N_5150);
or U9646 (N_9646,N_6847,N_6264);
xnor U9647 (N_9647,N_6419,N_5973);
nor U9648 (N_9648,N_6872,N_5850);
nand U9649 (N_9649,N_6476,N_6587);
nor U9650 (N_9650,N_5055,N_6169);
nand U9651 (N_9651,N_6948,N_7157);
or U9652 (N_9652,N_5524,N_5604);
nand U9653 (N_9653,N_7423,N_6792);
and U9654 (N_9654,N_6125,N_6181);
or U9655 (N_9655,N_7314,N_6924);
or U9656 (N_9656,N_7461,N_7350);
nor U9657 (N_9657,N_7489,N_5319);
or U9658 (N_9658,N_5089,N_5555);
or U9659 (N_9659,N_5358,N_6300);
nor U9660 (N_9660,N_6855,N_5177);
and U9661 (N_9661,N_5918,N_5037);
or U9662 (N_9662,N_5070,N_6380);
and U9663 (N_9663,N_7175,N_5057);
and U9664 (N_9664,N_6522,N_7315);
xnor U9665 (N_9665,N_5035,N_5579);
nand U9666 (N_9666,N_7036,N_7168);
nand U9667 (N_9667,N_5464,N_6873);
nand U9668 (N_9668,N_7270,N_7034);
and U9669 (N_9669,N_5822,N_6323);
or U9670 (N_9670,N_7446,N_5255);
or U9671 (N_9671,N_6620,N_7304);
and U9672 (N_9672,N_5872,N_5726);
or U9673 (N_9673,N_6369,N_5318);
or U9674 (N_9674,N_5878,N_6784);
nand U9675 (N_9675,N_5224,N_7387);
and U9676 (N_9676,N_5499,N_5248);
and U9677 (N_9677,N_6573,N_6798);
or U9678 (N_9678,N_6312,N_6360);
or U9679 (N_9679,N_5490,N_7288);
nand U9680 (N_9680,N_6123,N_5688);
and U9681 (N_9681,N_5774,N_6476);
nor U9682 (N_9682,N_5228,N_6235);
nor U9683 (N_9683,N_5718,N_7168);
nor U9684 (N_9684,N_5297,N_6500);
nor U9685 (N_9685,N_6383,N_6927);
nor U9686 (N_9686,N_5120,N_6777);
and U9687 (N_9687,N_6954,N_5537);
and U9688 (N_9688,N_5062,N_6189);
and U9689 (N_9689,N_5235,N_7452);
nor U9690 (N_9690,N_6794,N_5761);
and U9691 (N_9691,N_7436,N_6152);
or U9692 (N_9692,N_6968,N_7444);
or U9693 (N_9693,N_6444,N_7303);
nor U9694 (N_9694,N_7308,N_6333);
nand U9695 (N_9695,N_6790,N_5832);
nor U9696 (N_9696,N_5644,N_6292);
or U9697 (N_9697,N_6121,N_5745);
and U9698 (N_9698,N_6413,N_6768);
and U9699 (N_9699,N_6484,N_5599);
nor U9700 (N_9700,N_6660,N_7436);
nand U9701 (N_9701,N_6956,N_5605);
nand U9702 (N_9702,N_5974,N_7484);
nor U9703 (N_9703,N_6794,N_5703);
nor U9704 (N_9704,N_6055,N_5072);
nor U9705 (N_9705,N_6892,N_5235);
xor U9706 (N_9706,N_5423,N_5279);
or U9707 (N_9707,N_6007,N_6799);
nand U9708 (N_9708,N_6412,N_6462);
xnor U9709 (N_9709,N_6732,N_5729);
or U9710 (N_9710,N_5871,N_5094);
and U9711 (N_9711,N_7157,N_6987);
or U9712 (N_9712,N_5707,N_5477);
or U9713 (N_9713,N_7143,N_5480);
nor U9714 (N_9714,N_6995,N_6407);
and U9715 (N_9715,N_7364,N_7025);
and U9716 (N_9716,N_5610,N_7349);
nand U9717 (N_9717,N_6263,N_5656);
or U9718 (N_9718,N_5545,N_5250);
nor U9719 (N_9719,N_5530,N_5811);
or U9720 (N_9720,N_6694,N_5457);
and U9721 (N_9721,N_6949,N_6552);
nand U9722 (N_9722,N_6048,N_6686);
nor U9723 (N_9723,N_5562,N_7150);
nand U9724 (N_9724,N_5802,N_5725);
and U9725 (N_9725,N_6737,N_5175);
nor U9726 (N_9726,N_6903,N_6253);
or U9727 (N_9727,N_5849,N_6003);
and U9728 (N_9728,N_5835,N_5159);
or U9729 (N_9729,N_7056,N_7177);
nand U9730 (N_9730,N_6840,N_6434);
or U9731 (N_9731,N_7201,N_6525);
nand U9732 (N_9732,N_5943,N_5940);
nand U9733 (N_9733,N_6134,N_5820);
or U9734 (N_9734,N_5599,N_7409);
or U9735 (N_9735,N_6099,N_7116);
and U9736 (N_9736,N_5079,N_6258);
nand U9737 (N_9737,N_5262,N_6404);
and U9738 (N_9738,N_5780,N_7252);
or U9739 (N_9739,N_6694,N_6148);
or U9740 (N_9740,N_5971,N_5498);
nor U9741 (N_9741,N_6669,N_6534);
nor U9742 (N_9742,N_6411,N_6190);
and U9743 (N_9743,N_5842,N_6704);
and U9744 (N_9744,N_6362,N_7151);
and U9745 (N_9745,N_5838,N_5893);
nand U9746 (N_9746,N_5696,N_5697);
nor U9747 (N_9747,N_5013,N_7051);
or U9748 (N_9748,N_5986,N_5221);
xnor U9749 (N_9749,N_6225,N_6577);
nor U9750 (N_9750,N_5205,N_7086);
or U9751 (N_9751,N_7110,N_6205);
or U9752 (N_9752,N_6801,N_7044);
nand U9753 (N_9753,N_5895,N_5690);
xor U9754 (N_9754,N_7065,N_7323);
xor U9755 (N_9755,N_5299,N_6629);
or U9756 (N_9756,N_5065,N_5327);
nor U9757 (N_9757,N_5959,N_5389);
nor U9758 (N_9758,N_5270,N_5254);
nor U9759 (N_9759,N_7137,N_7286);
or U9760 (N_9760,N_7350,N_6457);
nand U9761 (N_9761,N_5038,N_5995);
nor U9762 (N_9762,N_5489,N_7265);
or U9763 (N_9763,N_6147,N_7033);
nor U9764 (N_9764,N_5170,N_6538);
or U9765 (N_9765,N_6314,N_6537);
and U9766 (N_9766,N_5218,N_5142);
xnor U9767 (N_9767,N_5524,N_7299);
nor U9768 (N_9768,N_6892,N_6995);
nand U9769 (N_9769,N_5971,N_6078);
or U9770 (N_9770,N_5646,N_6400);
and U9771 (N_9771,N_7219,N_6265);
or U9772 (N_9772,N_5855,N_5752);
and U9773 (N_9773,N_6642,N_5392);
nand U9774 (N_9774,N_7338,N_6128);
and U9775 (N_9775,N_5636,N_7411);
and U9776 (N_9776,N_6049,N_5097);
and U9777 (N_9777,N_6228,N_5566);
nand U9778 (N_9778,N_5347,N_6912);
and U9779 (N_9779,N_6065,N_6034);
nand U9780 (N_9780,N_5877,N_6663);
or U9781 (N_9781,N_6019,N_6693);
nand U9782 (N_9782,N_5093,N_6516);
and U9783 (N_9783,N_6141,N_7199);
or U9784 (N_9784,N_5191,N_7476);
nor U9785 (N_9785,N_5002,N_6745);
or U9786 (N_9786,N_6758,N_6818);
nand U9787 (N_9787,N_6504,N_6875);
nand U9788 (N_9788,N_7268,N_6358);
or U9789 (N_9789,N_5918,N_5314);
nor U9790 (N_9790,N_5197,N_6120);
xnor U9791 (N_9791,N_6217,N_7120);
and U9792 (N_9792,N_6090,N_5626);
or U9793 (N_9793,N_5252,N_6084);
or U9794 (N_9794,N_6390,N_6737);
nand U9795 (N_9795,N_5385,N_6384);
nand U9796 (N_9796,N_7093,N_6660);
and U9797 (N_9797,N_5747,N_6951);
and U9798 (N_9798,N_6134,N_5718);
or U9799 (N_9799,N_7041,N_5983);
nor U9800 (N_9800,N_7240,N_6529);
or U9801 (N_9801,N_5955,N_5340);
nor U9802 (N_9802,N_7127,N_5188);
and U9803 (N_9803,N_5422,N_6583);
xnor U9804 (N_9804,N_5290,N_5592);
or U9805 (N_9805,N_6146,N_6379);
nand U9806 (N_9806,N_5960,N_6223);
and U9807 (N_9807,N_6313,N_7415);
nor U9808 (N_9808,N_7468,N_6633);
nand U9809 (N_9809,N_5891,N_5079);
nand U9810 (N_9810,N_5976,N_5868);
nor U9811 (N_9811,N_6604,N_6011);
or U9812 (N_9812,N_5081,N_5550);
and U9813 (N_9813,N_5471,N_5793);
or U9814 (N_9814,N_7276,N_6598);
nor U9815 (N_9815,N_6246,N_6476);
or U9816 (N_9816,N_6804,N_6935);
and U9817 (N_9817,N_6038,N_7265);
nor U9818 (N_9818,N_5811,N_6141);
nand U9819 (N_9819,N_5857,N_5283);
or U9820 (N_9820,N_5691,N_6567);
or U9821 (N_9821,N_5281,N_7372);
and U9822 (N_9822,N_5872,N_5742);
nand U9823 (N_9823,N_6045,N_6392);
and U9824 (N_9824,N_5407,N_5608);
nor U9825 (N_9825,N_7283,N_6523);
or U9826 (N_9826,N_5838,N_5660);
nand U9827 (N_9827,N_6579,N_7428);
nand U9828 (N_9828,N_6495,N_6793);
nand U9829 (N_9829,N_6722,N_6831);
and U9830 (N_9830,N_6179,N_6532);
and U9831 (N_9831,N_6330,N_6218);
xor U9832 (N_9832,N_6750,N_6699);
or U9833 (N_9833,N_5655,N_6641);
or U9834 (N_9834,N_7176,N_6089);
nor U9835 (N_9835,N_6271,N_7234);
or U9836 (N_9836,N_6442,N_7380);
or U9837 (N_9837,N_5161,N_6469);
and U9838 (N_9838,N_6672,N_6668);
nand U9839 (N_9839,N_7459,N_5830);
or U9840 (N_9840,N_6428,N_5269);
nor U9841 (N_9841,N_7171,N_6288);
or U9842 (N_9842,N_6884,N_6116);
nor U9843 (N_9843,N_6901,N_5237);
nor U9844 (N_9844,N_5244,N_7235);
nand U9845 (N_9845,N_6913,N_5657);
nand U9846 (N_9846,N_6702,N_6841);
nand U9847 (N_9847,N_7224,N_7356);
nand U9848 (N_9848,N_6956,N_6011);
or U9849 (N_9849,N_5784,N_5000);
nor U9850 (N_9850,N_5943,N_7174);
nor U9851 (N_9851,N_7127,N_5057);
or U9852 (N_9852,N_6074,N_6757);
and U9853 (N_9853,N_6872,N_5206);
nor U9854 (N_9854,N_6532,N_6619);
nand U9855 (N_9855,N_7003,N_5902);
and U9856 (N_9856,N_5697,N_5787);
and U9857 (N_9857,N_5378,N_6578);
nand U9858 (N_9858,N_6845,N_5010);
and U9859 (N_9859,N_5312,N_7131);
nor U9860 (N_9860,N_6731,N_5047);
and U9861 (N_9861,N_7305,N_5696);
nor U9862 (N_9862,N_7269,N_5254);
or U9863 (N_9863,N_5510,N_6520);
or U9864 (N_9864,N_6351,N_5550);
nor U9865 (N_9865,N_5123,N_5565);
xor U9866 (N_9866,N_5413,N_6770);
and U9867 (N_9867,N_7026,N_5958);
or U9868 (N_9868,N_5395,N_7335);
xor U9869 (N_9869,N_7293,N_5924);
nor U9870 (N_9870,N_5153,N_6175);
nor U9871 (N_9871,N_5855,N_5218);
and U9872 (N_9872,N_7215,N_6918);
or U9873 (N_9873,N_5658,N_7349);
nor U9874 (N_9874,N_7355,N_7028);
nand U9875 (N_9875,N_5830,N_7102);
nor U9876 (N_9876,N_7187,N_5765);
or U9877 (N_9877,N_6029,N_5309);
and U9878 (N_9878,N_7058,N_5781);
and U9879 (N_9879,N_7290,N_7107);
nand U9880 (N_9880,N_5687,N_5913);
and U9881 (N_9881,N_6383,N_5861);
and U9882 (N_9882,N_7347,N_5069);
or U9883 (N_9883,N_6687,N_5851);
or U9884 (N_9884,N_6319,N_7377);
nand U9885 (N_9885,N_5257,N_7079);
nand U9886 (N_9886,N_7310,N_6601);
or U9887 (N_9887,N_6390,N_7104);
and U9888 (N_9888,N_6773,N_6960);
nor U9889 (N_9889,N_6652,N_6349);
and U9890 (N_9890,N_6487,N_6114);
and U9891 (N_9891,N_5230,N_6870);
nor U9892 (N_9892,N_6755,N_5080);
nor U9893 (N_9893,N_7132,N_7351);
and U9894 (N_9894,N_7047,N_7164);
nand U9895 (N_9895,N_6924,N_5822);
or U9896 (N_9896,N_6733,N_6774);
and U9897 (N_9897,N_5269,N_5040);
and U9898 (N_9898,N_6449,N_7329);
nand U9899 (N_9899,N_6952,N_5643);
nor U9900 (N_9900,N_6666,N_5549);
nand U9901 (N_9901,N_5715,N_6365);
and U9902 (N_9902,N_6124,N_5197);
or U9903 (N_9903,N_6575,N_7066);
nand U9904 (N_9904,N_5220,N_6267);
xnor U9905 (N_9905,N_5465,N_5652);
or U9906 (N_9906,N_6623,N_5325);
xnor U9907 (N_9907,N_5738,N_6339);
nor U9908 (N_9908,N_5241,N_5112);
nand U9909 (N_9909,N_6154,N_6834);
nand U9910 (N_9910,N_5959,N_5869);
and U9911 (N_9911,N_6212,N_6219);
or U9912 (N_9912,N_5647,N_7284);
or U9913 (N_9913,N_5178,N_7346);
nand U9914 (N_9914,N_6945,N_6645);
nor U9915 (N_9915,N_7259,N_5916);
xor U9916 (N_9916,N_5138,N_5351);
and U9917 (N_9917,N_6548,N_5884);
and U9918 (N_9918,N_6289,N_7086);
or U9919 (N_9919,N_6442,N_5427);
or U9920 (N_9920,N_6020,N_7368);
nor U9921 (N_9921,N_5377,N_5130);
or U9922 (N_9922,N_6316,N_6204);
or U9923 (N_9923,N_6658,N_5491);
and U9924 (N_9924,N_6334,N_5442);
nor U9925 (N_9925,N_5141,N_5571);
and U9926 (N_9926,N_6558,N_6356);
nand U9927 (N_9927,N_5316,N_6377);
and U9928 (N_9928,N_5193,N_6178);
or U9929 (N_9929,N_7369,N_5208);
or U9930 (N_9930,N_5263,N_5534);
or U9931 (N_9931,N_5039,N_6657);
and U9932 (N_9932,N_7007,N_5597);
nand U9933 (N_9933,N_5715,N_6670);
or U9934 (N_9934,N_5366,N_5159);
nand U9935 (N_9935,N_6979,N_7033);
and U9936 (N_9936,N_5590,N_6025);
and U9937 (N_9937,N_5997,N_6563);
nor U9938 (N_9938,N_6737,N_6445);
nand U9939 (N_9939,N_5913,N_5112);
nor U9940 (N_9940,N_5617,N_5962);
or U9941 (N_9941,N_5764,N_7223);
nor U9942 (N_9942,N_6338,N_5500);
or U9943 (N_9943,N_5130,N_7413);
nand U9944 (N_9944,N_6456,N_6096);
or U9945 (N_9945,N_7017,N_7147);
or U9946 (N_9946,N_7053,N_6972);
nor U9947 (N_9947,N_5758,N_5102);
xor U9948 (N_9948,N_6189,N_7286);
and U9949 (N_9949,N_5179,N_6169);
nor U9950 (N_9950,N_5274,N_6827);
nor U9951 (N_9951,N_5367,N_6757);
and U9952 (N_9952,N_6206,N_6445);
nor U9953 (N_9953,N_5417,N_6471);
nor U9954 (N_9954,N_5805,N_6113);
nand U9955 (N_9955,N_5903,N_6896);
and U9956 (N_9956,N_6763,N_6457);
or U9957 (N_9957,N_6426,N_6731);
nor U9958 (N_9958,N_6927,N_7400);
or U9959 (N_9959,N_6287,N_5741);
nand U9960 (N_9960,N_6854,N_5412);
nor U9961 (N_9961,N_5403,N_7370);
nand U9962 (N_9962,N_7237,N_5256);
nor U9963 (N_9963,N_5750,N_6036);
nand U9964 (N_9964,N_5637,N_5432);
or U9965 (N_9965,N_6725,N_5394);
nor U9966 (N_9966,N_6846,N_7483);
nor U9967 (N_9967,N_6355,N_6547);
or U9968 (N_9968,N_7055,N_6971);
or U9969 (N_9969,N_6010,N_7343);
and U9970 (N_9970,N_6617,N_5294);
nand U9971 (N_9971,N_7307,N_7110);
nand U9972 (N_9972,N_6386,N_6548);
nand U9973 (N_9973,N_7398,N_6827);
nand U9974 (N_9974,N_5867,N_6813);
nor U9975 (N_9975,N_7137,N_5187);
nand U9976 (N_9976,N_6776,N_6391);
nor U9977 (N_9977,N_6358,N_6332);
nor U9978 (N_9978,N_6746,N_6788);
or U9979 (N_9979,N_6651,N_6968);
nor U9980 (N_9980,N_5409,N_5784);
and U9981 (N_9981,N_7486,N_5338);
nand U9982 (N_9982,N_6848,N_7057);
or U9983 (N_9983,N_6241,N_7071);
or U9984 (N_9984,N_6279,N_6636);
and U9985 (N_9985,N_5728,N_5920);
xnor U9986 (N_9986,N_5225,N_6407);
and U9987 (N_9987,N_5370,N_6818);
nand U9988 (N_9988,N_5102,N_7323);
and U9989 (N_9989,N_6477,N_6302);
nand U9990 (N_9990,N_6634,N_5697);
or U9991 (N_9991,N_7310,N_6470);
and U9992 (N_9992,N_5429,N_5946);
nor U9993 (N_9993,N_5839,N_6419);
nand U9994 (N_9994,N_6118,N_6036);
or U9995 (N_9995,N_5828,N_6467);
nor U9996 (N_9996,N_6330,N_5214);
or U9997 (N_9997,N_5671,N_5101);
and U9998 (N_9998,N_5041,N_5574);
nand U9999 (N_9999,N_5479,N_6738);
or UO_0 (O_0,N_7962,N_8433);
nand UO_1 (O_1,N_9268,N_8408);
nor UO_2 (O_2,N_8125,N_8723);
nand UO_3 (O_3,N_7700,N_8384);
nand UO_4 (O_4,N_9640,N_8077);
and UO_5 (O_5,N_9600,N_8176);
nand UO_6 (O_6,N_8698,N_8790);
xnor UO_7 (O_7,N_8170,N_9708);
or UO_8 (O_8,N_8796,N_8775);
and UO_9 (O_9,N_8245,N_8058);
and UO_10 (O_10,N_8270,N_9248);
nand UO_11 (O_11,N_9283,N_8541);
or UO_12 (O_12,N_9701,N_7793);
nor UO_13 (O_13,N_8223,N_9187);
nor UO_14 (O_14,N_8745,N_9931);
nor UO_15 (O_15,N_9364,N_8147);
nor UO_16 (O_16,N_9919,N_9506);
and UO_17 (O_17,N_7605,N_9448);
nor UO_18 (O_18,N_9397,N_9146);
nor UO_19 (O_19,N_8478,N_7666);
and UO_20 (O_20,N_8192,N_9532);
nand UO_21 (O_21,N_8039,N_7881);
xnor UO_22 (O_22,N_7902,N_8087);
nor UO_23 (O_23,N_9104,N_8117);
nor UO_24 (O_24,N_8654,N_8590);
and UO_25 (O_25,N_9550,N_8203);
nor UO_26 (O_26,N_9790,N_8878);
or UO_27 (O_27,N_8500,N_7609);
nor UO_28 (O_28,N_9110,N_8581);
or UO_29 (O_29,N_9086,N_7848);
and UO_30 (O_30,N_8778,N_9686);
and UO_31 (O_31,N_8962,N_9244);
nand UO_32 (O_32,N_9592,N_7556);
xor UO_33 (O_33,N_8286,N_9040);
or UO_34 (O_34,N_7724,N_9261);
xnor UO_35 (O_35,N_9196,N_9973);
nor UO_36 (O_36,N_9336,N_8678);
nor UO_37 (O_37,N_7736,N_7882);
and UO_38 (O_38,N_8091,N_9420);
or UO_39 (O_39,N_9533,N_8266);
and UO_40 (O_40,N_9875,N_9867);
nor UO_41 (O_41,N_8320,N_9656);
nand UO_42 (O_42,N_9025,N_8481);
and UO_43 (O_43,N_9451,N_8934);
nand UO_44 (O_44,N_9596,N_8637);
or UO_45 (O_45,N_8886,N_8565);
and UO_46 (O_46,N_8363,N_9045);
nor UO_47 (O_47,N_8785,N_8052);
nor UO_48 (O_48,N_8564,N_8927);
and UO_49 (O_49,N_9015,N_7948);
nand UO_50 (O_50,N_9957,N_9907);
nand UO_51 (O_51,N_9180,N_9116);
and UO_52 (O_52,N_8197,N_8332);
nor UO_53 (O_53,N_8402,N_8587);
nand UO_54 (O_54,N_8630,N_8917);
nor UO_55 (O_55,N_9432,N_8706);
nor UO_56 (O_56,N_9011,N_9812);
xor UO_57 (O_57,N_9636,N_8764);
or UO_58 (O_58,N_8167,N_9270);
nand UO_59 (O_59,N_9682,N_7581);
nand UO_60 (O_60,N_7553,N_7812);
or UO_61 (O_61,N_8652,N_8939);
and UO_62 (O_62,N_9933,N_9173);
and UO_63 (O_63,N_8022,N_8949);
nor UO_64 (O_64,N_8891,N_8644);
nor UO_65 (O_65,N_9737,N_9013);
or UO_66 (O_66,N_8161,N_7791);
and UO_67 (O_67,N_9249,N_9413);
nand UO_68 (O_68,N_8748,N_9410);
nor UO_69 (O_69,N_9658,N_9746);
nor UO_70 (O_70,N_8633,N_7953);
nor UO_71 (O_71,N_7939,N_9387);
or UO_72 (O_72,N_7878,N_8726);
and UO_73 (O_73,N_7608,N_8829);
or UO_74 (O_74,N_8208,N_8072);
and UO_75 (O_75,N_8471,N_9102);
or UO_76 (O_76,N_7715,N_8997);
nand UO_77 (O_77,N_7831,N_9170);
and UO_78 (O_78,N_7932,N_9051);
and UO_79 (O_79,N_9767,N_8733);
nand UO_80 (O_80,N_7935,N_9510);
nand UO_81 (O_81,N_9172,N_7596);
nor UO_82 (O_82,N_9845,N_9329);
or UO_83 (O_83,N_7846,N_7680);
nor UO_84 (O_84,N_8018,N_9954);
nand UO_85 (O_85,N_7858,N_9368);
and UO_86 (O_86,N_9998,N_9624);
nor UO_87 (O_87,N_7699,N_8298);
and UO_88 (O_88,N_9318,N_8033);
nand UO_89 (O_89,N_7655,N_9811);
and UO_90 (O_90,N_8114,N_8529);
nand UO_91 (O_91,N_9833,N_8538);
or UO_92 (O_92,N_8101,N_8497);
nor UO_93 (O_93,N_7803,N_8990);
nand UO_94 (O_94,N_9393,N_9406);
and UO_95 (O_95,N_9455,N_9588);
and UO_96 (O_96,N_8913,N_8430);
xor UO_97 (O_97,N_8322,N_9466);
or UO_98 (O_98,N_9101,N_8936);
and UO_99 (O_99,N_8687,N_9788);
or UO_100 (O_100,N_8132,N_8234);
nand UO_101 (O_101,N_8046,N_8124);
or UO_102 (O_102,N_9956,N_9513);
nand UO_103 (O_103,N_9317,N_7901);
nor UO_104 (O_104,N_9552,N_7507);
xnor UO_105 (O_105,N_9348,N_8912);
nor UO_106 (O_106,N_8342,N_9810);
nor UO_107 (O_107,N_7915,N_9257);
nor UO_108 (O_108,N_9141,N_8391);
nor UO_109 (O_109,N_7573,N_7565);
nor UO_110 (O_110,N_9523,N_9351);
nor UO_111 (O_111,N_9654,N_7806);
nor UO_112 (O_112,N_7644,N_9326);
nand UO_113 (O_113,N_8404,N_7899);
nand UO_114 (O_114,N_8054,N_8274);
or UO_115 (O_115,N_9797,N_9107);
or UO_116 (O_116,N_9475,N_9117);
nor UO_117 (O_117,N_8434,N_8346);
nand UO_118 (O_118,N_9302,N_8051);
and UO_119 (O_119,N_9852,N_8691);
and UO_120 (O_120,N_7575,N_8100);
and UO_121 (O_121,N_7636,N_8888);
and UO_122 (O_122,N_9256,N_9203);
or UO_123 (O_123,N_8089,N_9255);
or UO_124 (O_124,N_8789,N_8506);
nor UO_125 (O_125,N_9704,N_9434);
or UO_126 (O_126,N_9356,N_9665);
nor UO_127 (O_127,N_8001,N_8589);
nand UO_128 (O_128,N_8436,N_9723);
and UO_129 (O_129,N_8839,N_8470);
nand UO_130 (O_130,N_9186,N_8923);
or UO_131 (O_131,N_8284,N_8961);
nor UO_132 (O_132,N_9539,N_9820);
nand UO_133 (O_133,N_7933,N_9199);
nor UO_134 (O_134,N_8112,N_8777);
nor UO_135 (O_135,N_8666,N_8884);
xnor UO_136 (O_136,N_8827,N_8216);
nor UO_137 (O_137,N_7892,N_8043);
nand UO_138 (O_138,N_7929,N_8562);
nand UO_139 (O_139,N_8915,N_8896);
or UO_140 (O_140,N_9238,N_7684);
or UO_141 (O_141,N_8289,N_7748);
nand UO_142 (O_142,N_7987,N_8853);
nand UO_143 (O_143,N_7864,N_8660);
nand UO_144 (O_144,N_8528,N_8304);
or UO_145 (O_145,N_9358,N_8452);
nor UO_146 (O_146,N_8484,N_8215);
and UO_147 (O_147,N_8754,N_8048);
and UO_148 (O_148,N_7629,N_8686);
nor UO_149 (O_149,N_9094,N_9328);
nor UO_150 (O_150,N_9923,N_8293);
nand UO_151 (O_151,N_9498,N_8211);
or UO_152 (O_152,N_8307,N_7865);
or UO_153 (O_153,N_7545,N_8258);
nor UO_154 (O_154,N_9716,N_8956);
nor UO_155 (O_155,N_7794,N_9740);
nand UO_156 (O_156,N_8979,N_8151);
nor UO_157 (O_157,N_8443,N_9603);
nand UO_158 (O_158,N_9555,N_9572);
and UO_159 (O_159,N_8584,N_9517);
nor UO_160 (O_160,N_8297,N_9285);
nor UO_161 (O_161,N_8537,N_9787);
and UO_162 (O_162,N_8422,N_9191);
nand UO_163 (O_163,N_8895,N_9727);
and UO_164 (O_164,N_7819,N_7652);
xnor UO_165 (O_165,N_9688,N_9304);
xor UO_166 (O_166,N_9939,N_7722);
and UO_167 (O_167,N_7702,N_9985);
xor UO_168 (O_168,N_9885,N_8805);
and UO_169 (O_169,N_7613,N_9216);
nor UO_170 (O_170,N_8916,N_9240);
and UO_171 (O_171,N_8393,N_7628);
nor UO_172 (O_172,N_7754,N_7975);
or UO_173 (O_173,N_8392,N_8467);
or UO_174 (O_174,N_7610,N_7895);
and UO_175 (O_175,N_9404,N_9075);
nand UO_176 (O_176,N_8677,N_8141);
nand UO_177 (O_177,N_8505,N_9394);
or UO_178 (O_178,N_7714,N_9158);
nor UO_179 (O_179,N_8664,N_9872);
or UO_180 (O_180,N_7734,N_9910);
or UO_181 (O_181,N_9766,N_9278);
and UO_182 (O_182,N_9068,N_7520);
or UO_183 (O_183,N_8116,N_9971);
or UO_184 (O_184,N_8327,N_9381);
nand UO_185 (O_185,N_9694,N_8194);
or UO_186 (O_186,N_8428,N_8256);
and UO_187 (O_187,N_9019,N_9211);
nor UO_188 (O_188,N_8974,N_8597);
nor UO_189 (O_189,N_9380,N_8948);
nand UO_190 (O_190,N_8239,N_8804);
nand UO_191 (O_191,N_9782,N_9021);
or UO_192 (O_192,N_7549,N_9604);
nor UO_193 (O_193,N_9222,N_9690);
and UO_194 (O_194,N_9259,N_7623);
xnor UO_195 (O_195,N_8069,N_8640);
nor UO_196 (O_196,N_8808,N_9389);
or UO_197 (O_197,N_8305,N_8591);
nor UO_198 (O_198,N_7822,N_8473);
nor UO_199 (O_199,N_8411,N_8740);
nor UO_200 (O_200,N_8746,N_8291);
xnor UO_201 (O_201,N_8155,N_8798);
nor UO_202 (O_202,N_8771,N_8094);
or UO_203 (O_203,N_7983,N_8314);
nand UO_204 (O_204,N_7993,N_9773);
or UO_205 (O_205,N_7536,N_7562);
and UO_206 (O_206,N_9247,N_9152);
and UO_207 (O_207,N_7578,N_8407);
nand UO_208 (O_208,N_7761,N_7758);
or UO_209 (O_209,N_8469,N_9728);
or UO_210 (O_210,N_9385,N_8819);
nand UO_211 (O_211,N_9783,N_7522);
or UO_212 (O_212,N_8079,N_7606);
nor UO_213 (O_213,N_8366,N_9722);
xor UO_214 (O_214,N_9936,N_7570);
nand UO_215 (O_215,N_9745,N_8813);
or UO_216 (O_216,N_8549,N_7688);
or UO_217 (O_217,N_8029,N_9006);
nand UO_218 (O_218,N_8930,N_7548);
nand UO_219 (O_219,N_9889,N_9043);
or UO_220 (O_220,N_9871,N_7701);
nand UO_221 (O_221,N_7537,N_8975);
and UO_222 (O_222,N_8011,N_8037);
nor UO_223 (O_223,N_8929,N_8960);
nor UO_224 (O_224,N_9135,N_9072);
nor UO_225 (O_225,N_8950,N_9534);
and UO_226 (O_226,N_9841,N_9252);
nand UO_227 (O_227,N_7946,N_9299);
and UO_228 (O_228,N_9946,N_8493);
xnor UO_229 (O_229,N_8440,N_9312);
or UO_230 (O_230,N_7571,N_9674);
or UO_231 (O_231,N_9613,N_9855);
nand UO_232 (O_232,N_7880,N_7854);
or UO_233 (O_233,N_7642,N_8999);
nand UO_234 (O_234,N_9288,N_9582);
nor UO_235 (O_235,N_9542,N_9258);
nor UO_236 (O_236,N_9402,N_8680);
and UO_237 (O_237,N_9932,N_7853);
and UO_238 (O_238,N_8350,N_8450);
or UO_239 (O_239,N_8665,N_9225);
or UO_240 (O_240,N_9725,N_7957);
nor UO_241 (O_241,N_7926,N_8833);
nor UO_242 (O_242,N_8889,N_9602);
or UO_243 (O_243,N_9770,N_8683);
nor UO_244 (O_244,N_8328,N_8026);
nor UO_245 (O_245,N_9494,N_9464);
and UO_246 (O_246,N_8892,N_8521);
nand UO_247 (O_247,N_7792,N_8871);
and UO_248 (O_248,N_8187,N_9063);
nor UO_249 (O_249,N_7810,N_9363);
or UO_250 (O_250,N_9961,N_7814);
or UO_251 (O_251,N_9324,N_9093);
and UO_252 (O_252,N_9501,N_8277);
and UO_253 (O_253,N_7723,N_8598);
nand UO_254 (O_254,N_9059,N_9357);
nor UO_255 (O_255,N_9988,N_9527);
nand UO_256 (O_256,N_8028,N_7826);
nor UO_257 (O_257,N_9468,N_8019);
nand UO_258 (O_258,N_8104,N_8514);
and UO_259 (O_259,N_9847,N_9126);
or UO_260 (O_260,N_7862,N_9729);
or UO_261 (O_261,N_9132,N_9755);
or UO_262 (O_262,N_9097,N_7569);
nand UO_263 (O_263,N_8682,N_8031);
or UO_264 (O_264,N_8618,N_7563);
nand UO_265 (O_265,N_9496,N_7801);
or UO_266 (O_266,N_7733,N_8164);
or UO_267 (O_267,N_8841,N_9091);
nor UO_268 (O_268,N_9470,N_8414);
or UO_269 (O_269,N_9499,N_8752);
nand UO_270 (O_270,N_8074,N_9497);
or UO_271 (O_271,N_9339,N_7711);
or UO_272 (O_272,N_9095,N_9689);
nand UO_273 (O_273,N_9515,N_9753);
nand UO_274 (O_274,N_8636,N_7572);
nand UO_275 (O_275,N_9041,N_9193);
nor UO_276 (O_276,N_9806,N_8449);
nand UO_277 (O_277,N_9298,N_9994);
or UO_278 (O_278,N_8082,N_9207);
or UO_279 (O_279,N_7779,N_8511);
nor UO_280 (O_280,N_7614,N_9700);
and UO_281 (O_281,N_7798,N_9712);
or UO_282 (O_282,N_9585,N_8247);
nor UO_283 (O_283,N_8042,N_8869);
xnor UO_284 (O_284,N_7739,N_9012);
and UO_285 (O_285,N_8045,N_9421);
nor UO_286 (O_286,N_9106,N_8204);
nand UO_287 (O_287,N_7682,N_8801);
and UO_288 (O_288,N_9438,N_9219);
and UO_289 (O_289,N_7675,N_7890);
or UO_290 (O_290,N_9149,N_7783);
or UO_291 (O_291,N_8476,N_8134);
or UO_292 (O_292,N_9112,N_8571);
or UO_293 (O_293,N_8122,N_8719);
or UO_294 (O_294,N_9154,N_9962);
or UO_295 (O_295,N_7799,N_8717);
or UO_296 (O_296,N_8133,N_8588);
nor UO_297 (O_297,N_7967,N_7938);
xor UO_298 (O_298,N_9004,N_7710);
nand UO_299 (O_299,N_8231,N_8238);
nor UO_300 (O_300,N_9853,N_8381);
and UO_301 (O_301,N_8842,N_8942);
and UO_302 (O_302,N_9379,N_7863);
and UO_303 (O_303,N_9566,N_9103);
nor UO_304 (O_304,N_9130,N_9964);
nand UO_305 (O_305,N_9284,N_9334);
or UO_306 (O_306,N_8338,N_9148);
or UO_307 (O_307,N_8527,N_8498);
nand UO_308 (O_308,N_9221,N_9802);
nand UO_309 (O_309,N_7871,N_8925);
nor UO_310 (O_310,N_8090,N_9338);
nand UO_311 (O_311,N_7960,N_7752);
or UO_312 (O_312,N_8820,N_7589);
and UO_313 (O_313,N_9245,N_9611);
and UO_314 (O_314,N_8821,N_8668);
nor UO_315 (O_315,N_9373,N_8697);
nor UO_316 (O_316,N_9442,N_9229);
nand UO_317 (O_317,N_8757,N_8799);
or UO_318 (O_318,N_7620,N_9975);
and UO_319 (O_319,N_8919,N_9064);
nand UO_320 (O_320,N_7557,N_8020);
nor UO_321 (O_321,N_8980,N_7961);
nand UO_322 (O_322,N_8149,N_8526);
and UO_323 (O_323,N_9017,N_7651);
nor UO_324 (O_324,N_9504,N_9078);
nor UO_325 (O_325,N_8670,N_9267);
nand UO_326 (O_326,N_8628,N_8749);
xor UO_327 (O_327,N_8202,N_8188);
nand UO_328 (O_328,N_8809,N_8490);
nor UO_329 (O_329,N_7927,N_9327);
nand UO_330 (O_330,N_8236,N_8047);
and UO_331 (O_331,N_9703,N_8814);
or UO_332 (O_332,N_9641,N_9441);
or UO_333 (O_333,N_8860,N_7603);
nor UO_334 (O_334,N_8978,N_8085);
and UO_335 (O_335,N_8106,N_7870);
or UO_336 (O_336,N_9092,N_9349);
and UO_337 (O_337,N_9220,N_9874);
or UO_338 (O_338,N_8403,N_9607);
or UO_339 (O_339,N_9558,N_9950);
nand UO_340 (O_340,N_7877,N_8863);
nor UO_341 (O_341,N_7698,N_9159);
nor UO_342 (O_342,N_8333,N_9809);
and UO_343 (O_343,N_9553,N_8413);
xor UO_344 (O_344,N_8520,N_9067);
and UO_345 (O_345,N_9991,N_7869);
nor UO_346 (O_346,N_8292,N_8845);
nor UO_347 (O_347,N_7815,N_9167);
nand UO_348 (O_348,N_8377,N_8220);
nor UO_349 (O_349,N_9635,N_7523);
xor UO_350 (O_350,N_8772,N_8463);
nand UO_351 (O_351,N_9129,N_8958);
nand UO_352 (O_352,N_8744,N_9065);
nand UO_353 (O_353,N_7668,N_8712);
and UO_354 (O_354,N_8575,N_9398);
and UO_355 (O_355,N_9807,N_7998);
or UO_356 (O_356,N_8613,N_7516);
nor UO_357 (O_357,N_8663,N_7588);
nor UO_358 (O_358,N_9821,N_7551);
or UO_359 (O_359,N_9291,N_7830);
nor UO_360 (O_360,N_8861,N_9374);
and UO_361 (O_361,N_7911,N_7958);
or UO_362 (O_362,N_8987,N_7641);
nor UO_363 (O_363,N_7705,N_7506);
or UO_364 (O_364,N_7991,N_8688);
or UO_365 (O_365,N_7847,N_7944);
nand UO_366 (O_366,N_9595,N_9835);
and UO_367 (O_367,N_9390,N_8225);
nor UO_368 (O_368,N_7740,N_7616);
nand UO_369 (O_369,N_8313,N_9754);
nor UO_370 (O_370,N_7823,N_8099);
nand UO_371 (O_371,N_9228,N_9431);
or UO_372 (O_372,N_8337,N_9137);
nor UO_373 (O_373,N_9779,N_8240);
or UO_374 (O_374,N_9382,N_8823);
and UO_375 (O_375,N_9408,N_8183);
nand UO_376 (O_376,N_8175,N_7727);
nor UO_377 (O_377,N_9726,N_9551);
nor UO_378 (O_378,N_7850,N_7693);
or UO_379 (O_379,N_9734,N_7947);
and UO_380 (O_380,N_9488,N_8868);
nor UO_381 (O_381,N_9647,N_9145);
nand UO_382 (O_382,N_9188,N_9519);
or UO_383 (O_383,N_9403,N_9756);
or UO_384 (O_384,N_8675,N_7787);
nand UO_385 (O_385,N_9540,N_9803);
or UO_386 (O_386,N_8097,N_8874);
or UO_387 (O_387,N_9623,N_7540);
or UO_388 (O_388,N_9058,N_9236);
nor UO_389 (O_389,N_9880,N_7832);
nand UO_390 (O_390,N_9644,N_7972);
nor UO_391 (O_391,N_8480,N_8570);
nand UO_392 (O_392,N_8992,N_9795);
and UO_393 (O_393,N_9090,N_8922);
or UO_394 (O_394,N_9630,N_7542);
or UO_395 (O_395,N_9346,N_9776);
and UO_396 (O_396,N_8872,N_8522);
or UO_397 (O_397,N_9929,N_8611);
nor UO_398 (O_398,N_9953,N_9817);
or UO_399 (O_399,N_8838,N_8770);
and UO_400 (O_400,N_8574,N_9436);
nand UO_401 (O_401,N_9096,N_9714);
and UO_402 (O_402,N_9127,N_8879);
nor UO_403 (O_403,N_9272,N_8062);
nand UO_404 (O_404,N_9054,N_9483);
or UO_405 (O_405,N_7839,N_9282);
nand UO_406 (O_406,N_7868,N_8120);
and UO_407 (O_407,N_7820,N_9921);
nor UO_408 (O_408,N_9634,N_8540);
nand UO_409 (O_409,N_7986,N_8271);
or UO_410 (O_410,N_7505,N_8750);
nor UO_411 (O_411,N_9616,N_8642);
xnor UO_412 (O_412,N_9952,N_7977);
nand UO_413 (O_413,N_9955,N_8931);
xor UO_414 (O_414,N_8139,N_8154);
or UO_415 (O_415,N_8646,N_9109);
nand UO_416 (O_416,N_9702,N_7866);
nor UO_417 (O_417,N_9347,N_7517);
nor UO_418 (O_418,N_9799,N_9968);
and UO_419 (O_419,N_8616,N_8013);
nand UO_420 (O_420,N_8601,N_8299);
or UO_421 (O_421,N_9560,N_7500);
or UO_422 (O_422,N_8780,N_9863);
nor UO_423 (O_423,N_7861,N_9816);
nand UO_424 (O_424,N_8036,N_7531);
or UO_425 (O_425,N_8453,N_7829);
xnor UO_426 (O_426,N_9509,N_8705);
nand UO_427 (O_427,N_9711,N_9705);
nor UO_428 (O_428,N_8951,N_8966);
or UO_429 (O_429,N_8907,N_8981);
nand UO_430 (O_430,N_8890,N_9586);
nand UO_431 (O_431,N_9650,N_9618);
and UO_432 (O_432,N_9485,N_9648);
and UO_433 (O_433,N_9206,N_9877);
and UO_434 (O_434,N_9111,N_9706);
nor UO_435 (O_435,N_9061,N_9492);
nand UO_436 (O_436,N_7679,N_8412);
and UO_437 (O_437,N_7547,N_8280);
or UO_438 (O_438,N_7757,N_8217);
and UO_439 (O_439,N_7844,N_9699);
nand UO_440 (O_440,N_8519,N_7533);
nor UO_441 (O_441,N_8315,N_8968);
nor UO_442 (O_442,N_7965,N_9502);
or UO_443 (O_443,N_8093,N_8765);
and UO_444 (O_444,N_8608,N_8118);
and UO_445 (O_445,N_9887,N_9342);
or UO_446 (O_446,N_8825,N_8834);
nor UO_447 (O_447,N_8437,N_9227);
nand UO_448 (O_448,N_8676,N_8472);
or UO_449 (O_449,N_8272,N_9030);
nand UO_450 (O_450,N_7851,N_9424);
nor UO_451 (O_451,N_9185,N_9049);
nand UO_452 (O_452,N_8083,N_9947);
nor UO_453 (O_453,N_8995,N_9233);
or UO_454 (O_454,N_9562,N_8973);
nand UO_455 (O_455,N_8615,N_8250);
or UO_456 (O_456,N_8397,N_8854);
nor UO_457 (O_457,N_9738,N_8877);
nand UO_458 (O_458,N_8938,N_9925);
and UO_459 (O_459,N_9984,N_9447);
or UO_460 (O_460,N_9565,N_8301);
nor UO_461 (O_461,N_9898,N_9995);
and UO_462 (O_462,N_8184,N_9399);
and UO_463 (O_463,N_9904,N_9698);
nand UO_464 (O_464,N_9815,N_9693);
or UO_465 (O_465,N_8483,N_8559);
and UO_466 (O_466,N_9440,N_8727);
and UO_467 (O_467,N_8002,N_7955);
nor UO_468 (O_468,N_8679,N_8901);
nor UO_469 (O_469,N_7692,N_7503);
or UO_470 (O_470,N_8362,N_8041);
or UO_471 (O_471,N_9578,N_8880);
nor UO_472 (O_472,N_8068,N_8131);
nor UO_473 (O_473,N_9166,N_9563);
nand UO_474 (O_474,N_7708,N_9200);
or UO_475 (O_475,N_7790,N_9123);
or UO_476 (O_476,N_8783,N_7514);
nor UO_477 (O_477,N_9575,N_7704);
nor UO_478 (O_478,N_9490,N_7583);
nor UO_479 (O_479,N_9281,N_8578);
nand UO_480 (O_480,N_7735,N_8228);
and UO_481 (O_481,N_8398,N_9718);
and UO_482 (O_482,N_7689,N_8351);
nand UO_483 (O_483,N_9361,N_8056);
nor UO_484 (O_484,N_9307,N_8319);
nand UO_485 (O_485,N_8507,N_8410);
nand UO_486 (O_486,N_8409,N_7974);
nor UO_487 (O_487,N_7501,N_8067);
nor UO_488 (O_488,N_8635,N_9290);
or UO_489 (O_489,N_8445,N_7905);
xnor UO_490 (O_490,N_9036,N_8826);
and UO_491 (O_491,N_7900,N_8699);
or UO_492 (O_492,N_7561,N_8572);
nor UO_493 (O_493,N_8004,N_9365);
and UO_494 (O_494,N_8797,N_8209);
nor UO_495 (O_495,N_8899,N_8283);
or UO_496 (O_496,N_9516,N_9453);
or UO_497 (O_497,N_8367,N_9444);
nand UO_498 (O_498,N_9423,N_9869);
or UO_499 (O_499,N_8257,N_9157);
nand UO_500 (O_500,N_8800,N_9121);
and UO_501 (O_501,N_9484,N_8906);
nand UO_502 (O_502,N_8510,N_9400);
or UO_503 (O_503,N_7867,N_8495);
nor UO_504 (O_504,N_7773,N_8386);
nand UO_505 (O_505,N_8693,N_8504);
nor UO_506 (O_506,N_9567,N_8290);
nand UO_507 (O_507,N_7622,N_8534);
nand UO_508 (O_508,N_7697,N_9246);
nor UO_509 (O_509,N_7802,N_9762);
or UO_510 (O_510,N_9114,N_7535);
xor UO_511 (O_511,N_9744,N_8760);
nor UO_512 (O_512,N_7836,N_8535);
or UO_513 (O_513,N_7769,N_7888);
and UO_514 (O_514,N_9024,N_8405);
or UO_515 (O_515,N_7889,N_8253);
nand UO_516 (O_516,N_8837,N_9987);
and UO_517 (O_517,N_7995,N_8904);
nor UO_518 (O_518,N_9183,N_9264);
and UO_519 (O_519,N_8025,N_9720);
or UO_520 (O_520,N_9859,N_9370);
nor UO_521 (O_521,N_7872,N_9664);
or UO_522 (O_522,N_8279,N_8784);
xor UO_523 (O_523,N_9824,N_8954);
or UO_524 (O_524,N_9164,N_9916);
and UO_525 (O_525,N_8459,N_9886);
or UO_526 (O_526,N_7604,N_9344);
and UO_527 (O_527,N_9591,N_7577);
and UO_528 (O_528,N_9162,N_7558);
and UO_529 (O_529,N_9028,N_7931);
nor UO_530 (O_530,N_9707,N_9868);
and UO_531 (O_531,N_9176,N_7539);
nor UO_532 (O_532,N_8200,N_8779);
or UO_533 (O_533,N_9633,N_7530);
nand UO_534 (O_534,N_8885,N_9174);
and UO_535 (O_535,N_9425,N_9412);
or UO_536 (O_536,N_9798,N_8150);
or UO_537 (O_537,N_9840,N_9360);
or UO_538 (O_538,N_8583,N_8650);
or UO_539 (O_539,N_7653,N_8840);
or UO_540 (O_540,N_7763,N_8689);
or UO_541 (O_541,N_8831,N_8457);
xor UO_542 (O_542,N_7716,N_8010);
and UO_543 (O_543,N_7560,N_9082);
and UO_544 (O_544,N_8364,N_8275);
and UO_545 (O_545,N_8791,N_8368);
nand UO_546 (O_546,N_7781,N_8373);
or UO_547 (O_547,N_7525,N_7592);
nor UO_548 (O_548,N_7904,N_7910);
nor UO_549 (O_549,N_8592,N_7941);
and UO_550 (O_550,N_9639,N_9894);
nand UO_551 (O_551,N_8621,N_8639);
and UO_552 (O_552,N_9593,N_8281);
nor UO_553 (O_553,N_8488,N_9352);
nand UO_554 (O_554,N_7743,N_9657);
or UO_555 (O_555,N_9179,N_7664);
and UO_556 (O_556,N_9771,N_9321);
nor UO_557 (O_557,N_9775,N_9056);
nor UO_558 (O_558,N_8985,N_9212);
nor UO_559 (O_559,N_7504,N_8172);
nor UO_560 (O_560,N_9917,N_9181);
or UO_561 (O_561,N_9764,N_9457);
or UO_562 (O_562,N_9153,N_8084);
or UO_563 (O_563,N_9266,N_8078);
nor UO_564 (O_564,N_7759,N_9308);
or UO_565 (O_565,N_9543,N_8802);
nand UO_566 (O_566,N_9669,N_9920);
and UO_567 (O_567,N_8517,N_8224);
and UO_568 (O_568,N_8066,N_8107);
or UO_569 (O_569,N_8810,N_7678);
nor UO_570 (O_570,N_8415,N_9459);
nor UO_571 (O_571,N_8695,N_8439);
nor UO_572 (O_572,N_9601,N_7738);
and UO_573 (O_573,N_9128,N_9142);
and UO_574 (O_574,N_7841,N_9621);
nand UO_575 (O_575,N_9763,N_8545);
or UO_576 (O_576,N_9758,N_9014);
and UO_577 (O_577,N_7981,N_8851);
and UO_578 (O_578,N_7766,N_8905);
and UO_579 (O_579,N_9508,N_8448);
xor UO_580 (O_580,N_8053,N_9277);
nand UO_581 (O_581,N_9751,N_9866);
xnor UO_582 (O_582,N_9202,N_9330);
nand UO_583 (O_583,N_9311,N_7663);
or UO_584 (O_584,N_7875,N_9922);
or UO_585 (O_585,N_9310,N_8921);
nand UO_586 (O_586,N_9651,N_7963);
nand UO_587 (O_587,N_9832,N_9343);
and UO_588 (O_588,N_8201,N_9411);
nand UO_589 (O_589,N_8694,N_9341);
and UO_590 (O_590,N_7706,N_8977);
or UO_591 (O_591,N_8474,N_7994);
and UO_592 (O_592,N_9271,N_7707);
nor UO_593 (O_593,N_8651,N_9032);
nand UO_594 (O_594,N_9739,N_7528);
nor UO_595 (O_595,N_9557,N_7951);
nor UO_596 (O_596,N_9990,N_8515);
and UO_597 (O_597,N_9967,N_9760);
and UO_598 (O_598,N_7665,N_9009);
nor UO_599 (O_599,N_9778,N_7891);
and UO_600 (O_600,N_7681,N_9541);
or UO_601 (O_601,N_8243,N_9736);
and UO_602 (O_602,N_7835,N_8909);
or UO_603 (O_603,N_7751,N_9668);
nor UO_604 (O_604,N_7750,N_9827);
nand UO_605 (O_605,N_8003,N_8395);
or UO_606 (O_606,N_8370,N_8662);
and UO_607 (O_607,N_8725,N_9934);
nand UO_608 (O_608,N_9804,N_9050);
and UO_609 (O_609,N_9377,N_8959);
nand UO_610 (O_610,N_8876,N_8123);
nor UO_611 (O_611,N_8898,N_7840);
nor UO_612 (O_612,N_9081,N_8858);
nor UO_613 (O_613,N_9823,N_7937);
nor UO_614 (O_614,N_9405,N_9375);
nor UO_615 (O_615,N_8494,N_8586);
and UO_616 (O_616,N_9914,N_9443);
nor UO_617 (O_617,N_9896,N_8806);
nor UO_618 (O_618,N_9481,N_9881);
nand UO_619 (O_619,N_8603,N_7550);
and UO_620 (O_620,N_9978,N_8612);
or UO_621 (O_621,N_8014,N_8811);
or UO_622 (O_622,N_7997,N_9655);
nand UO_623 (O_623,N_8599,N_9151);
and UO_624 (O_624,N_8702,N_8110);
nand UO_625 (O_625,N_9080,N_8617);
and UO_626 (O_626,N_8730,N_7767);
and UO_627 (O_627,N_9856,N_8873);
or UO_628 (O_628,N_9046,N_9752);
and UO_629 (O_629,N_7546,N_8701);
nand UO_630 (O_630,N_8070,N_8910);
nor UO_631 (O_631,N_9721,N_8994);
nor UO_632 (O_632,N_8012,N_7618);
or UO_633 (O_633,N_8465,N_9888);
and UO_634 (O_634,N_8169,N_9192);
and UO_635 (O_635,N_9430,N_9619);
and UO_636 (O_636,N_9645,N_7874);
nand UO_637 (O_637,N_9489,N_9482);
nand UO_638 (O_638,N_7909,N_7923);
and UO_639 (O_639,N_8918,N_9241);
nand UO_640 (O_640,N_7821,N_9479);
and UO_641 (O_641,N_9276,N_9301);
and UO_642 (O_642,N_9296,N_9610);
nand UO_643 (O_643,N_8179,N_8625);
nor UO_644 (O_644,N_7591,N_7541);
nand UO_645 (O_645,N_8944,N_7534);
and UO_646 (O_646,N_8967,N_7597);
nor UO_647 (O_647,N_9445,N_7725);
or UO_648 (O_648,N_7928,N_7670);
or UO_649 (O_649,N_8432,N_7796);
nand UO_650 (O_650,N_8551,N_8265);
or UO_651 (O_651,N_8729,N_9691);
and UO_652 (O_652,N_7656,N_8866);
nor UO_653 (O_653,N_8920,N_9825);
and UO_654 (O_654,N_7593,N_8554);
or UO_655 (O_655,N_8207,N_9449);
and UO_656 (O_656,N_9757,N_9458);
or UO_657 (O_657,N_9230,N_8242);
xnor UO_658 (O_658,N_9911,N_8807);
and UO_659 (O_659,N_8218,N_9437);
or UO_660 (O_660,N_8191,N_8524);
nand UO_661 (O_661,N_9662,N_8311);
and UO_662 (O_662,N_9982,N_8316);
or UO_663 (O_663,N_8181,N_9966);
nand UO_664 (O_664,N_8330,N_7524);
nor UO_665 (O_665,N_8902,N_8953);
nand UO_666 (O_666,N_8160,N_9275);
or UO_667 (O_667,N_8720,N_9055);
nand UO_668 (O_668,N_9500,N_9396);
or UO_669 (O_669,N_8627,N_8148);
nor UO_670 (O_670,N_9195,N_9367);
or UO_671 (O_671,N_7988,N_7619);
or UO_672 (O_672,N_9719,N_9609);
or UO_673 (O_673,N_8007,N_7753);
nor UO_674 (O_674,N_9355,N_9008);
nand UO_675 (O_675,N_9573,N_8848);
and UO_676 (O_676,N_9454,N_7934);
nor UO_677 (O_677,N_9478,N_8940);
or UO_678 (O_678,N_9253,N_9631);
nand UO_679 (O_679,N_8788,N_9568);
nand UO_680 (O_680,N_8552,N_7876);
nor UO_681 (O_681,N_9893,N_7607);
nand UO_682 (O_682,N_9687,N_8372);
nand UO_683 (O_683,N_9709,N_8882);
and UO_684 (O_684,N_8986,N_9676);
or UO_685 (O_685,N_9077,N_9608);
and UO_686 (O_686,N_8092,N_9020);
nor UO_687 (O_687,N_9133,N_7755);
and UO_688 (O_688,N_9401,N_8555);
and UO_689 (O_689,N_9125,N_8857);
and UO_690 (O_690,N_8832,N_8356);
or UO_691 (O_691,N_8105,N_8935);
nand UO_692 (O_692,N_8619,N_8263);
and UO_693 (O_693,N_9474,N_8251);
or UO_694 (O_694,N_9884,N_8976);
and UO_695 (O_695,N_8893,N_9452);
nand UO_696 (O_696,N_7859,N_8491);
nand UO_697 (O_697,N_7966,N_9819);
nand UO_698 (O_698,N_8331,N_7584);
nand UO_699 (O_699,N_8794,N_9140);
nor UO_700 (O_700,N_8163,N_8349);
nand UO_701 (O_701,N_9115,N_7837);
nor UO_702 (O_702,N_9122,N_9743);
nor UO_703 (O_703,N_8991,N_9559);
nor UO_704 (O_704,N_8344,N_8136);
nor UO_705 (O_705,N_9938,N_8246);
xnor UO_706 (O_706,N_8715,N_8850);
nor UO_707 (O_707,N_9912,N_8846);
nor UO_708 (O_708,N_7626,N_8768);
nor UO_709 (O_709,N_8908,N_8399);
and UO_710 (O_710,N_7729,N_8482);
nor UO_711 (O_711,N_9395,N_8401);
and UO_712 (O_712,N_8847,N_8875);
nor UO_713 (O_713,N_8566,N_8456);
nand UO_714 (O_714,N_9584,N_9581);
and UO_715 (O_715,N_7788,N_7741);
nor UO_716 (O_716,N_8460,N_7952);
and UO_717 (O_717,N_8631,N_7580);
nor UO_718 (O_718,N_8365,N_7599);
nand UO_719 (O_719,N_8387,N_7713);
nand UO_720 (O_720,N_8696,N_9100);
or UO_721 (O_721,N_8162,N_8946);
nor UO_722 (O_722,N_7638,N_9548);
nor UO_723 (O_723,N_8475,N_7612);
nor UO_724 (O_724,N_7646,N_8728);
and UO_725 (O_725,N_8911,N_8761);
nand UO_726 (O_726,N_7718,N_9201);
nand UO_727 (O_727,N_9861,N_8964);
or UO_728 (O_728,N_8605,N_8468);
nand UO_729 (O_729,N_8222,N_7717);
nor UO_730 (O_730,N_9322,N_9579);
and UO_731 (O_731,N_7985,N_9316);
or UO_732 (O_732,N_8034,N_7945);
or UO_733 (O_733,N_8516,N_7843);
or UO_734 (O_734,N_8230,N_7956);
or UO_735 (O_735,N_8166,N_7611);
or UO_736 (O_736,N_9465,N_9838);
nand UO_737 (O_737,N_9386,N_9035);
and UO_738 (O_738,N_7816,N_7598);
nor UO_739 (O_739,N_8751,N_9197);
and UO_740 (O_740,N_7756,N_9155);
or UO_741 (O_741,N_8221,N_9750);
nor UO_742 (O_742,N_9605,N_8455);
nor UO_743 (O_743,N_9683,N_7508);
or UO_744 (O_744,N_8803,N_8000);
and UO_745 (O_745,N_9890,N_8021);
and UO_746 (O_746,N_9315,N_8383);
nand UO_747 (O_747,N_9435,N_9416);
or UO_748 (O_748,N_9681,N_7778);
or UO_749 (O_749,N_9857,N_8418);
and UO_750 (O_750,N_9511,N_7567);
nor UO_751 (O_751,N_9801,N_9320);
nand UO_752 (O_752,N_7776,N_8512);
nand UO_753 (O_753,N_8431,N_9834);
or UO_754 (O_754,N_7852,N_9818);
or UO_755 (O_755,N_7509,N_9378);
nand UO_756 (O_756,N_9088,N_7659);
or UO_757 (O_757,N_9526,N_8732);
nand UO_758 (O_758,N_8196,N_9493);
nor UO_759 (O_759,N_7690,N_9168);
and UO_760 (O_760,N_7555,N_8487);
and UO_761 (O_761,N_9171,N_8157);
and UO_762 (O_762,N_7744,N_9844);
nor UO_763 (O_763,N_9554,N_8609);
and UO_764 (O_764,N_8641,N_8193);
or UO_765 (O_765,N_9476,N_9570);
xnor UO_766 (O_766,N_8674,N_7883);
nor UO_767 (O_767,N_7674,N_9977);
nand UO_768 (O_768,N_9429,N_9175);
nor UO_769 (O_769,N_8523,N_8576);
nand UO_770 (O_770,N_9908,N_9184);
or UO_771 (O_771,N_7726,N_9909);
nand UO_772 (O_772,N_9808,N_7807);
and UO_773 (O_773,N_9792,N_9362);
or UO_774 (O_774,N_8419,N_9214);
and UO_775 (O_775,N_9407,N_8427);
and UO_776 (O_776,N_7903,N_9765);
nand UO_777 (O_777,N_8969,N_9292);
and UO_778 (O_778,N_8897,N_8249);
or UO_779 (O_779,N_8038,N_8792);
or UO_780 (O_780,N_9848,N_9002);
nor UO_781 (O_781,N_7838,N_7709);
nor UO_782 (O_782,N_8632,N_7521);
or UO_783 (O_783,N_7694,N_7519);
nand UO_784 (O_784,N_8171,N_8489);
nor UO_785 (O_785,N_9450,N_8016);
nor UO_786 (O_786,N_9260,N_7654);
nand UO_787 (O_787,N_9314,N_7574);
nand UO_788 (O_788,N_9232,N_7980);
and UO_789 (O_789,N_9899,N_9461);
and UO_790 (O_790,N_8610,N_9371);
nor UO_791 (O_791,N_8126,N_8485);
nand UO_792 (O_792,N_9895,N_9085);
or UO_793 (O_793,N_9663,N_8561);
nand UO_794 (O_794,N_9741,N_7855);
nand UO_795 (O_795,N_8672,N_7797);
or UO_796 (O_796,N_7633,N_9518);
nor UO_797 (O_797,N_8008,N_8015);
or UO_798 (O_798,N_9243,N_9161);
or UO_799 (O_799,N_7703,N_9839);
and UO_800 (O_800,N_8624,N_9594);
nor UO_801 (O_801,N_7631,N_9235);
nand UO_802 (O_802,N_7720,N_8379);
or UO_803 (O_803,N_9587,N_9480);
nor UO_804 (O_804,N_9612,N_9018);
nand UO_805 (O_805,N_9678,N_9675);
nand UO_806 (O_806,N_8060,N_8195);
or UO_807 (O_807,N_8998,N_8032);
nor UO_808 (O_808,N_9460,N_9156);
and UO_809 (O_809,N_9969,N_7990);
and UO_810 (O_810,N_8759,N_8212);
nor UO_811 (O_811,N_9079,N_9622);
and UO_812 (O_812,N_8295,N_8098);
and UO_813 (O_813,N_7529,N_9794);
and UO_814 (O_814,N_8096,N_7842);
and UO_815 (O_815,N_9935,N_9124);
nor UO_816 (O_816,N_9627,N_9670);
and UO_817 (O_817,N_8531,N_8580);
nor UO_818 (O_818,N_9439,N_9785);
or UO_819 (O_819,N_9580,N_7999);
xor UO_820 (O_820,N_8335,N_8620);
and UO_821 (O_821,N_9525,N_9796);
nor UO_822 (O_822,N_9564,N_8657);
or UO_823 (O_823,N_9057,N_9666);
nor UO_824 (O_824,N_9590,N_9279);
and UO_825 (O_825,N_7824,N_8345);
nor UO_826 (O_826,N_7833,N_8734);
and UO_827 (O_827,N_7760,N_9940);
nor UO_828 (O_828,N_8185,N_8887);
nand UO_829 (O_829,N_8747,N_9083);
xor UO_830 (O_830,N_9671,N_7742);
xnor UO_831 (O_831,N_7804,N_9462);
nand UO_832 (O_832,N_9319,N_8260);
nor UO_833 (O_833,N_8709,N_7964);
or UO_834 (O_834,N_8816,N_8156);
nor UO_835 (O_835,N_7625,N_9960);
nand UO_836 (O_836,N_7749,N_8049);
or UO_837 (O_837,N_9697,N_8525);
and UO_838 (O_838,N_9544,N_8557);
nand UO_839 (O_839,N_8259,N_9118);
and UO_840 (O_840,N_9979,N_8774);
nand UO_841 (O_841,N_9959,N_7768);
nor UO_842 (O_842,N_8614,N_9569);
and UO_843 (O_843,N_8830,N_7908);
or UO_844 (O_844,N_7582,N_9426);
and UO_845 (O_845,N_9262,N_8982);
and UO_846 (O_846,N_9829,N_9027);
nand UO_847 (O_847,N_8237,N_9854);
nand UO_848 (O_848,N_9732,N_8343);
nor UO_849 (O_849,N_9672,N_9422);
and UO_850 (O_850,N_8380,N_8278);
nor UO_851 (O_851,N_7730,N_8543);
nand UO_852 (O_852,N_9177,N_8153);
and UO_853 (O_853,N_8812,N_8862);
and UO_854 (O_854,N_8758,N_8352);
or UO_855 (O_855,N_8458,N_8138);
nor UO_856 (O_856,N_7921,N_8262);
nor UO_857 (O_857,N_9287,N_9034);
and UO_858 (O_858,N_9948,N_9951);
or UO_859 (O_859,N_9473,N_9528);
nand UO_860 (O_860,N_9747,N_7686);
or UO_861 (O_861,N_7992,N_8057);
nor UO_862 (O_862,N_9108,N_9208);
nand UO_863 (O_863,N_8645,N_9507);
nor UO_864 (O_864,N_7950,N_7856);
or UO_865 (O_865,N_9696,N_8268);
and UO_866 (O_866,N_8119,N_7979);
nor UO_867 (O_867,N_8241,N_8205);
and UO_868 (O_868,N_8669,N_7913);
nand UO_869 (O_869,N_8903,N_9297);
and UO_870 (O_870,N_8198,N_7673);
nor UO_871 (O_871,N_8382,N_8933);
or UO_872 (O_872,N_8129,N_8795);
and UO_873 (O_873,N_9001,N_9026);
nor UO_874 (O_874,N_7772,N_7647);
or UO_875 (O_875,N_9680,N_8499);
or UO_876 (O_876,N_9918,N_7894);
or UO_877 (O_877,N_9409,N_8369);
and UO_878 (O_878,N_9073,N_9016);
nand UO_879 (O_879,N_9937,N_9883);
or UO_880 (O_880,N_9044,N_9606);
nor UO_881 (O_881,N_8681,N_9822);
and UO_882 (O_882,N_9902,N_9814);
nand UO_883 (O_883,N_8718,N_7634);
and UO_884 (O_884,N_7630,N_9837);
or UO_885 (O_885,N_9944,N_8030);
or UO_886 (O_886,N_8753,N_9529);
nand UO_887 (O_887,N_8182,N_8086);
nand UO_888 (O_888,N_8690,N_9384);
nand UO_889 (O_889,N_9303,N_9333);
nand UO_890 (O_890,N_8996,N_8040);
nand UO_891 (O_891,N_9274,N_9223);
nor UO_892 (O_892,N_9226,N_8835);
nand UO_893 (O_893,N_7667,N_9667);
nand UO_894 (O_894,N_8648,N_7637);
nand UO_895 (O_895,N_8340,N_9945);
and UO_896 (O_896,N_9620,N_7825);
or UO_897 (O_897,N_7936,N_8984);
nand UO_898 (O_898,N_8359,N_9769);
and UO_899 (O_899,N_8109,N_7887);
nor UO_900 (O_900,N_8423,N_8883);
and UO_901 (O_901,N_7879,N_8406);
nand UO_902 (O_902,N_8623,N_7687);
nand UO_903 (O_903,N_8424,N_8971);
or UO_904 (O_904,N_9428,N_9392);
or UO_905 (O_905,N_7512,N_7552);
nor UO_906 (O_906,N_9391,N_7527);
or UO_907 (O_907,N_9661,N_8102);
nor UO_908 (O_908,N_8108,N_9735);
nor UO_909 (O_909,N_7918,N_7639);
nor UO_910 (O_910,N_9524,N_8255);
and UO_911 (O_911,N_8993,N_8288);
nand UO_912 (O_912,N_8711,N_8317);
nor UO_913 (O_913,N_9642,N_8867);
nor UO_914 (O_914,N_8075,N_9242);
nor UO_915 (O_915,N_9224,N_9649);
and UO_916 (O_916,N_7513,N_9843);
and UO_917 (O_917,N_9637,N_8357);
nand UO_918 (O_918,N_8607,N_9724);
nor UO_919 (O_919,N_9836,N_9891);
nand UO_920 (O_920,N_9561,N_9074);
or UO_921 (O_921,N_9521,N_8513);
nor UO_922 (O_922,N_9038,N_9858);
and UO_923 (O_923,N_9150,N_7968);
and UO_924 (O_924,N_8739,N_9294);
nor UO_925 (O_925,N_9194,N_8708);
nand UO_926 (O_926,N_8115,N_9069);
nand UO_927 (O_927,N_9643,N_9846);
nor UO_928 (O_928,N_9331,N_7845);
nand UO_929 (O_929,N_8302,N_8130);
nand UO_930 (O_930,N_9210,N_8065);
nand UO_931 (O_931,N_8376,N_8773);
nand UO_932 (O_932,N_9419,N_9949);
or UO_933 (O_933,N_9066,N_7943);
or UO_934 (O_934,N_7989,N_7721);
and UO_935 (O_935,N_9695,N_8137);
and UO_936 (O_936,N_7982,N_8140);
nand UO_937 (O_937,N_9383,N_7595);
nor UO_938 (O_938,N_8685,N_8661);
and UO_939 (O_939,N_8941,N_9325);
or UO_940 (O_940,N_8312,N_7621);
or UO_941 (O_941,N_8568,N_8210);
nand UO_942 (O_942,N_9269,N_8721);
nor UO_943 (O_943,N_8963,N_9217);
or UO_944 (O_944,N_8518,N_8159);
nor UO_945 (O_945,N_8214,N_9306);
or UO_946 (O_946,N_8178,N_9415);
nor UO_947 (O_947,N_8174,N_8937);
or UO_948 (O_948,N_8310,N_7897);
or UO_949 (O_949,N_8264,N_9335);
nor UO_950 (O_950,N_8849,N_9427);
nand UO_951 (O_951,N_8190,N_8658);
nor UO_952 (O_952,N_9289,N_8707);
or UO_953 (O_953,N_8955,N_8128);
and UO_954 (O_954,N_7912,N_9060);
nand UO_955 (O_955,N_8815,N_8553);
or UO_956 (O_956,N_8671,N_8731);
and UO_957 (O_957,N_8080,N_7789);
and UO_958 (O_958,N_7954,N_9793);
nand UO_959 (O_959,N_8569,N_9062);
nand UO_960 (O_960,N_9571,N_7885);
and UO_961 (O_961,N_8444,N_8146);
or UO_962 (O_962,N_8546,N_9512);
and UO_963 (O_963,N_8005,N_9350);
nand UO_964 (O_964,N_9472,N_8856);
or UO_965 (O_965,N_9547,N_9372);
or UO_966 (O_966,N_9039,N_9731);
nand UO_967 (O_967,N_8273,N_9250);
or UO_968 (O_968,N_8378,N_9927);
or UO_969 (O_969,N_8285,N_8582);
nor UO_970 (O_970,N_8325,N_7615);
and UO_971 (O_971,N_7919,N_8318);
or UO_972 (O_972,N_9295,N_9029);
nand UO_973 (O_973,N_9878,N_8111);
and UO_974 (O_974,N_9313,N_8818);
nor UO_975 (O_975,N_9906,N_7774);
and UO_976 (O_976,N_9537,N_9549);
or UO_977 (O_977,N_9000,N_8451);
or UO_978 (O_978,N_9433,N_7526);
and UO_979 (O_979,N_8076,N_7683);
and UO_980 (O_980,N_8213,N_8303);
nand UO_981 (O_981,N_8604,N_9087);
and UO_982 (O_982,N_8595,N_8972);
nor UO_983 (O_983,N_7942,N_8550);
nand UO_984 (O_984,N_8502,N_8324);
and UO_985 (O_985,N_9237,N_9628);
nand UO_986 (O_986,N_7811,N_8429);
or UO_987 (O_987,N_7800,N_9471);
or UO_988 (O_988,N_8466,N_7566);
or UO_989 (O_989,N_9099,N_9842);
or UO_990 (O_990,N_7970,N_8061);
or UO_991 (O_991,N_7728,N_9781);
and UO_992 (O_992,N_8653,N_8339);
nand UO_993 (O_993,N_7662,N_7643);
nand UO_994 (O_994,N_8742,N_8769);
or UO_995 (O_995,N_8714,N_8396);
or UO_996 (O_996,N_9713,N_7924);
and UO_997 (O_997,N_9928,N_8308);
nor UO_998 (O_998,N_8441,N_8113);
and UO_999 (O_999,N_9981,N_7896);
or UO_1000 (O_1000,N_8782,N_9505);
or UO_1001 (O_1001,N_7920,N_9418);
nor UO_1002 (O_1002,N_7515,N_7917);
and UO_1003 (O_1003,N_8044,N_9048);
nand UO_1004 (O_1004,N_9996,N_8988);
and UO_1005 (O_1005,N_8673,N_8165);
nor UO_1006 (O_1006,N_8957,N_8287);
nand UO_1007 (O_1007,N_7930,N_8542);
nand UO_1008 (O_1008,N_9556,N_8716);
nand UO_1009 (O_1009,N_9986,N_8928);
and UO_1010 (O_1010,N_8269,N_9417);
and UO_1011 (O_1011,N_7671,N_9042);
nand UO_1012 (O_1012,N_8276,N_8756);
and UO_1013 (O_1013,N_8649,N_7518);
xor UO_1014 (O_1014,N_8596,N_7969);
nor UO_1015 (O_1015,N_8509,N_9487);
nor UO_1016 (O_1016,N_7747,N_9198);
or UO_1017 (O_1017,N_9491,N_7922);
nor UO_1018 (O_1018,N_8006,N_9997);
nand UO_1019 (O_1019,N_7696,N_8643);
or UO_1020 (O_1020,N_9254,N_9828);
nor UO_1021 (O_1021,N_7914,N_9323);
xor UO_1022 (O_1022,N_9305,N_9007);
nand UO_1023 (O_1023,N_8244,N_8755);
nor UO_1024 (O_1024,N_8371,N_8844);
or UO_1025 (O_1025,N_7916,N_8232);
nor UO_1026 (O_1026,N_7996,N_8121);
nor UO_1027 (O_1027,N_8703,N_8594);
and UO_1028 (O_1028,N_9538,N_8943);
or UO_1029 (O_1029,N_8722,N_7672);
or UO_1030 (O_1030,N_7818,N_8659);
nor UO_1031 (O_1031,N_9742,N_8656);
or UO_1032 (O_1032,N_9629,N_7857);
or UO_1033 (O_1033,N_9677,N_9800);
nand UO_1034 (O_1034,N_8144,N_8142);
or UO_1035 (O_1035,N_9178,N_8334);
nand UO_1036 (O_1036,N_9768,N_9414);
nand UO_1037 (O_1037,N_8508,N_7640);
or UO_1038 (O_1038,N_9646,N_9989);
nor UO_1039 (O_1039,N_8063,N_8477);
nor UO_1040 (O_1040,N_8438,N_9865);
and UO_1041 (O_1041,N_7978,N_9169);
nor UO_1042 (O_1042,N_8306,N_7658);
nand UO_1043 (O_1043,N_7971,N_8323);
and UO_1044 (O_1044,N_9280,N_9189);
and UO_1045 (O_1045,N_8563,N_9999);
xnor UO_1046 (O_1046,N_8446,N_8127);
nand UO_1047 (O_1047,N_9332,N_8965);
and UO_1048 (O_1048,N_7886,N_7594);
and UO_1049 (O_1049,N_8309,N_9879);
nor UO_1050 (O_1050,N_8186,N_7737);
or UO_1051 (O_1051,N_7586,N_7632);
and UO_1052 (O_1052,N_9638,N_9577);
nand UO_1053 (O_1053,N_8983,N_7732);
and UO_1054 (O_1054,N_7510,N_8738);
or UO_1055 (O_1055,N_9786,N_7600);
nor UO_1056 (O_1056,N_8704,N_9265);
nand UO_1057 (O_1057,N_8647,N_9514);
or UO_1058 (O_1058,N_9876,N_9780);
nand UO_1059 (O_1059,N_8233,N_7559);
nand UO_1060 (O_1060,N_9251,N_8388);
nand UO_1061 (O_1061,N_9924,N_8462);
or UO_1062 (O_1062,N_8881,N_8533);
nand UO_1063 (O_1063,N_9503,N_8435);
or UO_1064 (O_1064,N_8655,N_9182);
nor UO_1065 (O_1065,N_8763,N_8035);
nor UO_1066 (O_1066,N_9830,N_9761);
or UO_1067 (O_1067,N_9805,N_9530);
nor UO_1068 (O_1068,N_8824,N_9772);
xnor UO_1069 (O_1069,N_8600,N_8634);
and UO_1070 (O_1070,N_9138,N_9531);
nor UO_1071 (O_1071,N_8454,N_7695);
nor UO_1072 (O_1072,N_9851,N_9882);
and UO_1073 (O_1073,N_9353,N_8952);
or UO_1074 (O_1074,N_8737,N_9826);
nor UO_1075 (O_1075,N_8743,N_9345);
and UO_1076 (O_1076,N_7691,N_9469);
nor UO_1077 (O_1077,N_8023,N_8180);
nor UO_1078 (O_1078,N_8321,N_9495);
and UO_1079 (O_1079,N_9119,N_9231);
nor UO_1080 (O_1080,N_9589,N_8294);
nand UO_1081 (O_1081,N_9748,N_9930);
or UO_1082 (O_1082,N_9071,N_9205);
nor UO_1083 (O_1083,N_7925,N_9733);
nand UO_1084 (O_1084,N_7669,N_9749);
and UO_1085 (O_1085,N_8817,N_9023);
or UO_1086 (O_1086,N_8852,N_9113);
nand UO_1087 (O_1087,N_9897,N_9905);
and UO_1088 (O_1088,N_8055,N_9831);
and UO_1089 (O_1089,N_8300,N_9576);
or UO_1090 (O_1090,N_9467,N_8088);
nand UO_1091 (O_1091,N_9915,N_9120);
nor UO_1092 (O_1092,N_9536,N_8787);
nand UO_1093 (O_1093,N_7940,N_8261);
or UO_1094 (O_1094,N_8447,N_8579);
or UO_1095 (O_1095,N_9147,N_9913);
nand UO_1096 (O_1096,N_8024,N_9037);
nand UO_1097 (O_1097,N_7677,N_8135);
nor UO_1098 (O_1098,N_8606,N_8282);
and UO_1099 (O_1099,N_7762,N_9134);
nand UO_1100 (O_1100,N_9993,N_9165);
nor UO_1101 (O_1101,N_8227,N_7775);
and UO_1102 (O_1102,N_8168,N_8173);
nand UO_1103 (O_1103,N_8385,N_9903);
and UO_1104 (O_1104,N_9789,N_9900);
or UO_1105 (O_1105,N_8989,N_7764);
nand UO_1106 (O_1106,N_9862,N_7786);
nor UO_1107 (O_1107,N_7601,N_8544);
and UO_1108 (O_1108,N_9974,N_9263);
nand UO_1109 (O_1109,N_9053,N_9653);
nor UO_1110 (O_1110,N_9583,N_9983);
and UO_1111 (O_1111,N_9163,N_8865);
or UO_1112 (O_1112,N_8793,N_9359);
nand UO_1113 (O_1113,N_9293,N_8479);
and UO_1114 (O_1114,N_8864,N_9234);
and UO_1115 (O_1115,N_9340,N_8235);
and UO_1116 (O_1116,N_9047,N_8776);
or UO_1117 (O_1117,N_7554,N_9715);
nand UO_1118 (O_1118,N_9777,N_7645);
nand UO_1119 (O_1119,N_9546,N_9477);
nor UO_1120 (O_1120,N_7782,N_7543);
and UO_1121 (O_1121,N_9076,N_8389);
nor UO_1122 (O_1122,N_7780,N_9717);
or UO_1123 (O_1123,N_7765,N_9943);
and UO_1124 (O_1124,N_7795,N_9366);
xor UO_1125 (O_1125,N_8638,N_8073);
and UO_1126 (O_1126,N_8158,N_7564);
nand UO_1127 (O_1127,N_9992,N_7834);
nand UO_1128 (O_1128,N_8420,N_8461);
nor UO_1129 (O_1129,N_9965,N_9144);
or UO_1130 (O_1130,N_9679,N_9901);
nand UO_1131 (O_1131,N_8558,N_8219);
and UO_1132 (O_1132,N_9574,N_8700);
nor UO_1133 (O_1133,N_8828,N_8464);
nand UO_1134 (O_1134,N_9005,N_9052);
nor UO_1135 (O_1135,N_8692,N_9209);
or UO_1136 (O_1136,N_8767,N_9870);
and UO_1137 (O_1137,N_7544,N_8486);
and UO_1138 (O_1138,N_7568,N_9131);
nand UO_1139 (O_1139,N_9213,N_8017);
and UO_1140 (O_1140,N_7770,N_7949);
nand UO_1141 (O_1141,N_8347,N_9942);
nor UO_1142 (O_1142,N_8425,N_7828);
nor UO_1143 (O_1143,N_7893,N_9849);
nor UO_1144 (O_1144,N_8348,N_9599);
nor UO_1145 (O_1145,N_7746,N_8547);
nor UO_1146 (O_1146,N_7712,N_9660);
and UO_1147 (O_1147,N_9010,N_7771);
and UO_1148 (O_1148,N_9520,N_8360);
or UO_1149 (O_1149,N_8602,N_9376);
and UO_1150 (O_1150,N_8766,N_9033);
or UO_1151 (O_1151,N_8836,N_9273);
and UO_1152 (O_1152,N_8593,N_9139);
or UO_1153 (O_1153,N_8496,N_9652);
or UO_1154 (O_1154,N_8924,N_9813);
and UO_1155 (O_1155,N_8573,N_8926);
nor UO_1156 (O_1156,N_9617,N_8532);
nand UO_1157 (O_1157,N_7976,N_8354);
nand UO_1158 (O_1158,N_8252,N_8855);
nand UO_1159 (O_1159,N_7617,N_8417);
nor UO_1160 (O_1160,N_8358,N_9286);
and UO_1161 (O_1161,N_8710,N_9976);
nand UO_1162 (O_1162,N_7635,N_8741);
nand UO_1163 (O_1163,N_8859,N_8567);
nand UO_1164 (O_1164,N_7731,N_9597);
nor UO_1165 (O_1165,N_9215,N_8713);
nand UO_1166 (O_1166,N_8254,N_9926);
or UO_1167 (O_1167,N_8199,N_7898);
and UO_1168 (O_1168,N_9892,N_7984);
or UO_1169 (O_1169,N_8059,N_8667);
and UO_1170 (O_1170,N_9337,N_7511);
or UO_1171 (O_1171,N_8914,N_9239);
or UO_1172 (O_1172,N_8442,N_9958);
and UO_1173 (O_1173,N_9759,N_7809);
xor UO_1174 (O_1174,N_8536,N_8932);
nor UO_1175 (O_1175,N_8095,N_7502);
or UO_1176 (O_1176,N_8145,N_7906);
or UO_1177 (O_1177,N_9309,N_9160);
and UO_1178 (O_1178,N_9598,N_9486);
nor UO_1179 (O_1179,N_9626,N_7576);
or UO_1180 (O_1180,N_7860,N_7805);
or UO_1181 (O_1181,N_8539,N_7884);
or UO_1182 (O_1182,N_7784,N_7777);
nand UO_1183 (O_1183,N_8416,N_8009);
nor UO_1184 (O_1184,N_8189,N_7585);
nand UO_1185 (O_1185,N_9970,N_9941);
nand UO_1186 (O_1186,N_9522,N_9615);
and UO_1187 (O_1187,N_8735,N_8870);
and UO_1188 (O_1188,N_7590,N_8081);
or UO_1189 (O_1189,N_9136,N_9873);
nor UO_1190 (O_1190,N_7973,N_8822);
or UO_1191 (O_1191,N_8336,N_8375);
and UO_1192 (O_1192,N_8786,N_8355);
or UO_1193 (O_1193,N_9084,N_8361);
and UO_1194 (O_1194,N_7538,N_8296);
or UO_1195 (O_1195,N_9730,N_8341);
or UO_1196 (O_1196,N_9190,N_7649);
and UO_1197 (O_1197,N_8206,N_8152);
nor UO_1198 (O_1198,N_9850,N_8071);
or UO_1199 (O_1199,N_8426,N_9774);
and UO_1200 (O_1200,N_8143,N_7579);
nand UO_1201 (O_1201,N_8894,N_7719);
nand UO_1202 (O_1202,N_9864,N_8626);
or UO_1203 (O_1203,N_9625,N_8900);
nand UO_1204 (O_1204,N_7602,N_8762);
or UO_1205 (O_1205,N_9963,N_8781);
nand UO_1206 (O_1206,N_8585,N_8622);
or UO_1207 (O_1207,N_9098,N_7745);
or UO_1208 (O_1208,N_9692,N_9456);
or UO_1209 (O_1209,N_8503,N_9659);
and UO_1210 (O_1210,N_8329,N_7650);
and UO_1211 (O_1211,N_8400,N_9105);
nor UO_1212 (O_1212,N_8843,N_8492);
nor UO_1213 (O_1213,N_9446,N_8970);
or UO_1214 (O_1214,N_9972,N_8064);
xor UO_1215 (O_1215,N_8736,N_9614);
or UO_1216 (O_1216,N_7676,N_7624);
nor UO_1217 (O_1217,N_7627,N_8390);
and UO_1218 (O_1218,N_8326,N_7685);
and UO_1219 (O_1219,N_8629,N_7849);
nand UO_1220 (O_1220,N_8530,N_9143);
nand UO_1221 (O_1221,N_9218,N_8947);
and UO_1222 (O_1222,N_7813,N_7817);
nand UO_1223 (O_1223,N_7827,N_9300);
nor UO_1224 (O_1224,N_9784,N_8945);
or UO_1225 (O_1225,N_8421,N_7873);
or UO_1226 (O_1226,N_8501,N_9710);
nand UO_1227 (O_1227,N_8226,N_8560);
xnor UO_1228 (O_1228,N_7657,N_8556);
and UO_1229 (O_1229,N_8684,N_8027);
or UO_1230 (O_1230,N_8267,N_9632);
nor UO_1231 (O_1231,N_7587,N_9070);
nor UO_1232 (O_1232,N_8548,N_9673);
or UO_1233 (O_1233,N_9003,N_8050);
nor UO_1234 (O_1234,N_7648,N_7661);
and UO_1235 (O_1235,N_9980,N_8229);
and UO_1236 (O_1236,N_9685,N_9545);
xnor UO_1237 (O_1237,N_9204,N_7907);
nand UO_1238 (O_1238,N_9791,N_8577);
xor UO_1239 (O_1239,N_7532,N_9860);
nand UO_1240 (O_1240,N_7808,N_8394);
and UO_1241 (O_1241,N_7785,N_7959);
and UO_1242 (O_1242,N_9369,N_9022);
nand UO_1243 (O_1243,N_9354,N_9684);
nand UO_1244 (O_1244,N_9089,N_8177);
nor UO_1245 (O_1245,N_9463,N_9031);
or UO_1246 (O_1246,N_7660,N_8724);
nand UO_1247 (O_1247,N_9388,N_8374);
and UO_1248 (O_1248,N_8353,N_9535);
and UO_1249 (O_1249,N_8103,N_8248);
and UO_1250 (O_1250,N_9570,N_9974);
or UO_1251 (O_1251,N_9263,N_7964);
nor UO_1252 (O_1252,N_7546,N_8973);
nor UO_1253 (O_1253,N_8023,N_8712);
nor UO_1254 (O_1254,N_7586,N_7637);
and UO_1255 (O_1255,N_9388,N_9842);
nand UO_1256 (O_1256,N_8289,N_7826);
nand UO_1257 (O_1257,N_8881,N_9626);
nand UO_1258 (O_1258,N_9541,N_8242);
or UO_1259 (O_1259,N_9402,N_9933);
and UO_1260 (O_1260,N_9579,N_7982);
and UO_1261 (O_1261,N_8592,N_7697);
nand UO_1262 (O_1262,N_7978,N_7981);
nor UO_1263 (O_1263,N_8952,N_9050);
or UO_1264 (O_1264,N_8334,N_9735);
nor UO_1265 (O_1265,N_7647,N_9299);
and UO_1266 (O_1266,N_9804,N_9232);
nor UO_1267 (O_1267,N_9389,N_8299);
and UO_1268 (O_1268,N_9064,N_9027);
or UO_1269 (O_1269,N_9417,N_8735);
nand UO_1270 (O_1270,N_7519,N_9224);
or UO_1271 (O_1271,N_8576,N_9332);
and UO_1272 (O_1272,N_9089,N_8852);
nand UO_1273 (O_1273,N_8067,N_9805);
or UO_1274 (O_1274,N_7524,N_9600);
nand UO_1275 (O_1275,N_9933,N_8838);
nand UO_1276 (O_1276,N_8890,N_7838);
nand UO_1277 (O_1277,N_7807,N_8850);
and UO_1278 (O_1278,N_9908,N_9159);
nand UO_1279 (O_1279,N_9597,N_7583);
or UO_1280 (O_1280,N_9002,N_8655);
and UO_1281 (O_1281,N_9016,N_8082);
and UO_1282 (O_1282,N_8407,N_9980);
nor UO_1283 (O_1283,N_9265,N_7766);
and UO_1284 (O_1284,N_7664,N_9462);
or UO_1285 (O_1285,N_9344,N_7877);
and UO_1286 (O_1286,N_9787,N_8631);
xnor UO_1287 (O_1287,N_7994,N_8111);
nand UO_1288 (O_1288,N_7766,N_8535);
and UO_1289 (O_1289,N_7613,N_9464);
and UO_1290 (O_1290,N_9973,N_9390);
and UO_1291 (O_1291,N_8880,N_8240);
and UO_1292 (O_1292,N_7531,N_9963);
nand UO_1293 (O_1293,N_7847,N_7727);
nor UO_1294 (O_1294,N_8778,N_8341);
or UO_1295 (O_1295,N_8193,N_8146);
nor UO_1296 (O_1296,N_7759,N_7609);
nor UO_1297 (O_1297,N_9094,N_8625);
and UO_1298 (O_1298,N_9643,N_9515);
and UO_1299 (O_1299,N_7546,N_9770);
nor UO_1300 (O_1300,N_8155,N_7754);
nor UO_1301 (O_1301,N_9220,N_9486);
nand UO_1302 (O_1302,N_9061,N_8455);
nand UO_1303 (O_1303,N_7804,N_9017);
nor UO_1304 (O_1304,N_9152,N_8550);
and UO_1305 (O_1305,N_8646,N_8134);
xor UO_1306 (O_1306,N_8241,N_8646);
and UO_1307 (O_1307,N_8009,N_9122);
or UO_1308 (O_1308,N_7822,N_9684);
or UO_1309 (O_1309,N_9443,N_8827);
and UO_1310 (O_1310,N_9355,N_7802);
and UO_1311 (O_1311,N_7602,N_8371);
or UO_1312 (O_1312,N_8958,N_8507);
nor UO_1313 (O_1313,N_8109,N_8462);
and UO_1314 (O_1314,N_8252,N_9179);
or UO_1315 (O_1315,N_8101,N_9691);
or UO_1316 (O_1316,N_8086,N_9467);
nor UO_1317 (O_1317,N_8769,N_9058);
or UO_1318 (O_1318,N_8634,N_8091);
or UO_1319 (O_1319,N_8485,N_7955);
xor UO_1320 (O_1320,N_9754,N_8876);
nor UO_1321 (O_1321,N_9137,N_8217);
and UO_1322 (O_1322,N_8851,N_8173);
nor UO_1323 (O_1323,N_8835,N_8008);
or UO_1324 (O_1324,N_8975,N_9647);
nor UO_1325 (O_1325,N_8546,N_8968);
or UO_1326 (O_1326,N_9523,N_9530);
nor UO_1327 (O_1327,N_9258,N_9298);
or UO_1328 (O_1328,N_9003,N_8022);
nor UO_1329 (O_1329,N_9504,N_9487);
or UO_1330 (O_1330,N_8652,N_8471);
nor UO_1331 (O_1331,N_8779,N_9737);
and UO_1332 (O_1332,N_7854,N_8689);
and UO_1333 (O_1333,N_9667,N_8933);
nand UO_1334 (O_1334,N_7925,N_7588);
or UO_1335 (O_1335,N_7505,N_8358);
and UO_1336 (O_1336,N_8094,N_8577);
and UO_1337 (O_1337,N_9671,N_9595);
nand UO_1338 (O_1338,N_9887,N_8079);
nor UO_1339 (O_1339,N_8491,N_7842);
and UO_1340 (O_1340,N_8700,N_8828);
xor UO_1341 (O_1341,N_9624,N_9917);
nor UO_1342 (O_1342,N_9697,N_9295);
nand UO_1343 (O_1343,N_9900,N_8030);
nand UO_1344 (O_1344,N_8199,N_8821);
nor UO_1345 (O_1345,N_8221,N_9009);
and UO_1346 (O_1346,N_9677,N_9358);
nand UO_1347 (O_1347,N_7834,N_9320);
and UO_1348 (O_1348,N_7791,N_9257);
and UO_1349 (O_1349,N_8735,N_9914);
and UO_1350 (O_1350,N_8050,N_7579);
and UO_1351 (O_1351,N_8597,N_8863);
and UO_1352 (O_1352,N_9474,N_7940);
or UO_1353 (O_1353,N_9942,N_7570);
nand UO_1354 (O_1354,N_7941,N_9385);
or UO_1355 (O_1355,N_9467,N_9209);
and UO_1356 (O_1356,N_8695,N_8927);
or UO_1357 (O_1357,N_7885,N_8585);
xnor UO_1358 (O_1358,N_8035,N_8848);
xor UO_1359 (O_1359,N_7814,N_7556);
nand UO_1360 (O_1360,N_8615,N_9224);
and UO_1361 (O_1361,N_8651,N_8577);
nand UO_1362 (O_1362,N_8416,N_8614);
nor UO_1363 (O_1363,N_7688,N_8110);
nand UO_1364 (O_1364,N_8682,N_7983);
or UO_1365 (O_1365,N_9680,N_9418);
nand UO_1366 (O_1366,N_9719,N_8222);
and UO_1367 (O_1367,N_7550,N_9071);
and UO_1368 (O_1368,N_8606,N_9762);
and UO_1369 (O_1369,N_8604,N_9897);
or UO_1370 (O_1370,N_7879,N_7984);
and UO_1371 (O_1371,N_7689,N_8930);
or UO_1372 (O_1372,N_8740,N_9168);
and UO_1373 (O_1373,N_8536,N_9186);
nor UO_1374 (O_1374,N_9570,N_9148);
and UO_1375 (O_1375,N_8512,N_9211);
and UO_1376 (O_1376,N_9699,N_7814);
nor UO_1377 (O_1377,N_8721,N_8060);
or UO_1378 (O_1378,N_7946,N_7855);
nand UO_1379 (O_1379,N_9466,N_9901);
nor UO_1380 (O_1380,N_9376,N_8903);
and UO_1381 (O_1381,N_9570,N_8699);
or UO_1382 (O_1382,N_9932,N_8596);
or UO_1383 (O_1383,N_9619,N_8782);
nor UO_1384 (O_1384,N_8771,N_9405);
nand UO_1385 (O_1385,N_8667,N_8357);
nand UO_1386 (O_1386,N_7678,N_8620);
and UO_1387 (O_1387,N_7568,N_7519);
nand UO_1388 (O_1388,N_9408,N_7601);
or UO_1389 (O_1389,N_8825,N_8118);
and UO_1390 (O_1390,N_7767,N_9043);
nand UO_1391 (O_1391,N_8731,N_8353);
nand UO_1392 (O_1392,N_9842,N_9421);
nor UO_1393 (O_1393,N_7955,N_8678);
or UO_1394 (O_1394,N_8575,N_9186);
or UO_1395 (O_1395,N_9967,N_9567);
and UO_1396 (O_1396,N_7759,N_9867);
or UO_1397 (O_1397,N_7695,N_9603);
and UO_1398 (O_1398,N_9993,N_8615);
or UO_1399 (O_1399,N_9490,N_9085);
and UO_1400 (O_1400,N_7954,N_7845);
xor UO_1401 (O_1401,N_7820,N_8869);
nand UO_1402 (O_1402,N_9386,N_7945);
or UO_1403 (O_1403,N_9760,N_9526);
xor UO_1404 (O_1404,N_9443,N_7855);
nand UO_1405 (O_1405,N_7573,N_8513);
or UO_1406 (O_1406,N_9692,N_9084);
nor UO_1407 (O_1407,N_8052,N_8846);
nor UO_1408 (O_1408,N_8482,N_9164);
nor UO_1409 (O_1409,N_8877,N_7694);
nand UO_1410 (O_1410,N_8895,N_8432);
and UO_1411 (O_1411,N_9212,N_8132);
and UO_1412 (O_1412,N_8592,N_9627);
nand UO_1413 (O_1413,N_9397,N_9732);
and UO_1414 (O_1414,N_8406,N_7620);
or UO_1415 (O_1415,N_8742,N_8199);
or UO_1416 (O_1416,N_9792,N_9932);
or UO_1417 (O_1417,N_8258,N_9034);
or UO_1418 (O_1418,N_8130,N_9965);
and UO_1419 (O_1419,N_7929,N_7862);
nor UO_1420 (O_1420,N_8750,N_8883);
or UO_1421 (O_1421,N_8739,N_8211);
nand UO_1422 (O_1422,N_9968,N_9168);
or UO_1423 (O_1423,N_9364,N_8977);
and UO_1424 (O_1424,N_8021,N_8719);
or UO_1425 (O_1425,N_9529,N_7639);
and UO_1426 (O_1426,N_7740,N_7545);
or UO_1427 (O_1427,N_8902,N_9704);
and UO_1428 (O_1428,N_8609,N_8936);
nor UO_1429 (O_1429,N_9466,N_8268);
nor UO_1430 (O_1430,N_8081,N_8974);
nor UO_1431 (O_1431,N_9807,N_8514);
and UO_1432 (O_1432,N_9636,N_9009);
or UO_1433 (O_1433,N_8845,N_8794);
nand UO_1434 (O_1434,N_9677,N_9157);
and UO_1435 (O_1435,N_8242,N_8875);
or UO_1436 (O_1436,N_9965,N_8299);
nand UO_1437 (O_1437,N_9740,N_8419);
nand UO_1438 (O_1438,N_8606,N_9295);
or UO_1439 (O_1439,N_8525,N_8081);
nand UO_1440 (O_1440,N_8674,N_8817);
or UO_1441 (O_1441,N_9218,N_9913);
nand UO_1442 (O_1442,N_7601,N_7879);
and UO_1443 (O_1443,N_7960,N_8540);
nor UO_1444 (O_1444,N_7902,N_8948);
nand UO_1445 (O_1445,N_8068,N_8772);
nor UO_1446 (O_1446,N_7582,N_8059);
and UO_1447 (O_1447,N_7649,N_9268);
nor UO_1448 (O_1448,N_8448,N_7768);
or UO_1449 (O_1449,N_8239,N_8856);
or UO_1450 (O_1450,N_9261,N_8606);
and UO_1451 (O_1451,N_9675,N_8849);
nor UO_1452 (O_1452,N_8741,N_9004);
and UO_1453 (O_1453,N_8396,N_8809);
and UO_1454 (O_1454,N_8379,N_8971);
and UO_1455 (O_1455,N_7612,N_9130);
xnor UO_1456 (O_1456,N_9511,N_8122);
nor UO_1457 (O_1457,N_9705,N_9419);
and UO_1458 (O_1458,N_9449,N_9497);
and UO_1459 (O_1459,N_9457,N_9672);
and UO_1460 (O_1460,N_9338,N_7733);
nor UO_1461 (O_1461,N_8233,N_8516);
and UO_1462 (O_1462,N_9761,N_9850);
or UO_1463 (O_1463,N_8187,N_8649);
nand UO_1464 (O_1464,N_8514,N_7744);
or UO_1465 (O_1465,N_8229,N_7552);
and UO_1466 (O_1466,N_9767,N_7821);
nor UO_1467 (O_1467,N_8883,N_8449);
nor UO_1468 (O_1468,N_9932,N_8166);
or UO_1469 (O_1469,N_8521,N_9553);
or UO_1470 (O_1470,N_8825,N_8098);
nor UO_1471 (O_1471,N_9522,N_8991);
nand UO_1472 (O_1472,N_7838,N_9377);
nor UO_1473 (O_1473,N_8704,N_9596);
nor UO_1474 (O_1474,N_8583,N_9704);
nand UO_1475 (O_1475,N_7782,N_8595);
or UO_1476 (O_1476,N_8066,N_8022);
and UO_1477 (O_1477,N_9921,N_9458);
nor UO_1478 (O_1478,N_7711,N_8284);
nor UO_1479 (O_1479,N_9295,N_8933);
nand UO_1480 (O_1480,N_8096,N_7520);
or UO_1481 (O_1481,N_7653,N_9742);
nor UO_1482 (O_1482,N_7837,N_8832);
or UO_1483 (O_1483,N_9619,N_8450);
and UO_1484 (O_1484,N_8873,N_8500);
nand UO_1485 (O_1485,N_8369,N_9145);
and UO_1486 (O_1486,N_8694,N_8021);
or UO_1487 (O_1487,N_8697,N_9081);
and UO_1488 (O_1488,N_9164,N_9975);
or UO_1489 (O_1489,N_8541,N_8561);
nor UO_1490 (O_1490,N_9139,N_9690);
nand UO_1491 (O_1491,N_7816,N_9515);
nand UO_1492 (O_1492,N_7655,N_8199);
nor UO_1493 (O_1493,N_9522,N_8565);
nand UO_1494 (O_1494,N_9672,N_7719);
nand UO_1495 (O_1495,N_8247,N_9631);
and UO_1496 (O_1496,N_8377,N_9438);
nor UO_1497 (O_1497,N_9213,N_8164);
nor UO_1498 (O_1498,N_8359,N_8003);
and UO_1499 (O_1499,N_9504,N_9127);
endmodule