module basic_500_3000_500_50_levels_2xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_133,In_367);
and U1 (N_1,In_372,In_78);
nand U2 (N_2,In_432,In_400);
nor U3 (N_3,In_20,In_131);
nand U4 (N_4,In_61,In_88);
or U5 (N_5,In_220,In_363);
or U6 (N_6,In_34,In_163);
nand U7 (N_7,In_129,In_484);
nand U8 (N_8,In_461,In_257);
or U9 (N_9,In_409,In_355);
xor U10 (N_10,In_240,In_354);
nor U11 (N_11,In_251,In_307);
and U12 (N_12,In_419,In_105);
nand U13 (N_13,In_237,In_35);
and U14 (N_14,In_384,In_150);
or U15 (N_15,In_118,In_315);
xor U16 (N_16,In_36,In_197);
xnor U17 (N_17,In_42,In_290);
nor U18 (N_18,In_256,In_438);
nor U19 (N_19,In_296,In_292);
nor U20 (N_20,In_134,In_71);
and U21 (N_21,In_450,In_176);
xnor U22 (N_22,In_491,In_120);
nand U23 (N_23,In_386,In_281);
or U24 (N_24,In_459,In_286);
nand U25 (N_25,In_229,In_404);
or U26 (N_26,In_244,In_454);
or U27 (N_27,In_322,In_106);
nand U28 (N_28,In_216,In_53);
and U29 (N_29,In_250,In_184);
or U30 (N_30,In_275,In_164);
or U31 (N_31,In_331,In_142);
nor U32 (N_32,In_98,In_239);
and U33 (N_33,In_127,In_73);
nor U34 (N_34,In_55,In_72);
and U35 (N_35,In_125,In_447);
nor U36 (N_36,In_300,In_249);
and U37 (N_37,In_497,In_448);
or U38 (N_38,In_429,In_130);
and U39 (N_39,In_80,In_190);
nor U40 (N_40,In_375,In_117);
nand U41 (N_41,In_264,In_314);
or U42 (N_42,In_340,In_136);
nor U43 (N_43,In_43,In_68);
or U44 (N_44,In_449,In_19);
and U45 (N_45,In_310,In_319);
nand U46 (N_46,In_496,In_308);
nand U47 (N_47,In_199,In_94);
and U48 (N_48,In_223,In_172);
nor U49 (N_49,In_65,In_205);
nand U50 (N_50,In_393,In_316);
nor U51 (N_51,In_111,In_417);
or U52 (N_52,In_392,In_334);
or U53 (N_53,In_152,In_396);
and U54 (N_54,In_420,In_69);
nor U55 (N_55,In_58,In_489);
and U56 (N_56,In_138,In_347);
and U57 (N_57,In_299,In_3);
nand U58 (N_58,In_439,In_265);
nand U59 (N_59,In_301,In_132);
nand U60 (N_60,In_415,In_14);
or U61 (N_61,In_82,In_26);
nand U62 (N_62,In_333,In_276);
and U63 (N_63,In_233,In_102);
nand U64 (N_64,In_227,In_294);
nor U65 (N_65,In_371,In_402);
or U66 (N_66,In_104,In_303);
nand U67 (N_67,In_85,N_48);
xnor U68 (N_68,In_262,In_66);
and U69 (N_69,In_173,In_270);
nor U70 (N_70,N_36,In_206);
or U71 (N_71,In_293,In_304);
or U72 (N_72,In_200,In_4);
and U73 (N_73,In_477,In_469);
nand U74 (N_74,In_215,In_39);
or U75 (N_75,In_253,In_346);
nor U76 (N_76,N_39,In_312);
and U77 (N_77,In_122,In_178);
nand U78 (N_78,In_271,In_466);
and U79 (N_79,In_428,In_370);
or U80 (N_80,In_350,In_70);
nor U81 (N_81,In_268,In_202);
nand U82 (N_82,In_252,In_311);
nand U83 (N_83,In_101,In_12);
nand U84 (N_84,In_187,In_156);
xor U85 (N_85,In_362,In_0);
and U86 (N_86,N_47,In_189);
nor U87 (N_87,In_493,In_425);
and U88 (N_88,In_284,In_395);
and U89 (N_89,N_37,In_388);
nand U90 (N_90,N_40,N_0);
nor U91 (N_91,In_295,In_435);
nor U92 (N_92,In_481,In_24);
nor U93 (N_93,In_325,N_18);
or U94 (N_94,In_231,In_47);
and U95 (N_95,In_398,In_441);
nor U96 (N_96,In_499,In_259);
nor U97 (N_97,In_46,In_280);
nor U98 (N_98,N_21,N_29);
or U99 (N_99,In_203,In_91);
or U100 (N_100,In_475,In_326);
nand U101 (N_101,In_234,In_298);
nand U102 (N_102,In_40,In_451);
or U103 (N_103,N_53,N_44);
or U104 (N_104,In_146,In_309);
nand U105 (N_105,In_29,In_181);
nand U106 (N_106,In_490,N_34);
nor U107 (N_107,In_140,In_457);
and U108 (N_108,In_198,In_107);
and U109 (N_109,In_153,In_443);
or U110 (N_110,In_471,In_54);
or U111 (N_111,N_19,In_179);
nor U112 (N_112,In_480,In_336);
or U113 (N_113,In_149,In_483);
or U114 (N_114,In_147,N_58);
nor U115 (N_115,In_313,In_405);
nand U116 (N_116,In_28,In_135);
nor U117 (N_117,In_278,In_210);
and U118 (N_118,In_25,In_341);
nand U119 (N_119,In_317,In_247);
nand U120 (N_120,In_380,In_182);
or U121 (N_121,In_267,In_460);
and U122 (N_122,In_38,N_38);
or U123 (N_123,In_11,N_15);
or U124 (N_124,N_88,In_273);
or U125 (N_125,In_95,In_279);
nand U126 (N_126,In_175,In_403);
nand U127 (N_127,In_30,In_49);
nor U128 (N_128,In_196,N_90);
or U129 (N_129,In_414,In_285);
or U130 (N_130,In_476,N_13);
and U131 (N_131,In_155,N_25);
nor U132 (N_132,In_166,N_108);
nor U133 (N_133,In_387,In_306);
nor U134 (N_134,N_2,In_406);
and U135 (N_135,In_114,In_389);
nand U136 (N_136,In_62,In_385);
or U137 (N_137,In_453,N_30);
nand U138 (N_138,In_201,In_174);
nor U139 (N_139,N_85,N_57);
nor U140 (N_140,In_288,In_151);
or U141 (N_141,In_359,N_63);
nor U142 (N_142,In_494,In_245);
nor U143 (N_143,In_467,In_472);
nor U144 (N_144,N_72,N_7);
and U145 (N_145,In_15,In_431);
and U146 (N_146,In_446,In_186);
nand U147 (N_147,In_373,In_8);
and U148 (N_148,In_32,In_185);
or U149 (N_149,N_32,In_368);
and U150 (N_150,N_22,In_23);
or U151 (N_151,In_59,In_337);
nor U152 (N_152,N_42,In_241);
nand U153 (N_153,In_492,In_243);
nand U154 (N_154,N_106,In_16);
nor U155 (N_155,N_95,In_144);
or U156 (N_156,In_486,N_50);
nand U157 (N_157,N_113,In_327);
nand U158 (N_158,N_55,In_67);
and U159 (N_159,In_44,N_8);
or U160 (N_160,N_45,In_260);
and U161 (N_161,In_209,In_413);
nor U162 (N_162,In_440,In_90);
nor U163 (N_163,N_119,In_407);
nor U164 (N_164,In_103,In_180);
or U165 (N_165,In_169,N_114);
or U166 (N_166,In_269,In_2);
and U167 (N_167,In_328,In_320);
nor U168 (N_168,In_305,In_57);
nand U169 (N_169,In_342,N_60);
nor U170 (N_170,N_20,N_71);
nand U171 (N_171,In_128,In_485);
and U172 (N_172,In_408,In_246);
nor U173 (N_173,In_226,In_109);
and U174 (N_174,In_33,In_100);
nand U175 (N_175,N_78,In_21);
nand U176 (N_176,In_365,In_235);
or U177 (N_177,In_302,In_52);
nor U178 (N_178,In_424,In_255);
and U179 (N_179,In_86,In_361);
nand U180 (N_180,In_455,In_258);
nor U181 (N_181,N_16,N_173);
nor U182 (N_182,In_79,N_152);
or U183 (N_183,N_143,In_50);
nor U184 (N_184,In_412,In_277);
nor U185 (N_185,In_498,N_74);
nand U186 (N_186,N_70,In_126);
nor U187 (N_187,N_137,In_148);
nor U188 (N_188,In_157,In_391);
and U189 (N_189,In_442,N_89);
nor U190 (N_190,In_353,In_390);
and U191 (N_191,In_113,N_91);
nand U192 (N_192,N_132,N_122);
and U193 (N_193,N_124,In_445);
nand U194 (N_194,N_100,In_115);
nand U195 (N_195,In_323,In_339);
nand U196 (N_196,In_397,In_369);
nand U197 (N_197,In_158,In_236);
or U198 (N_198,In_364,N_35);
and U199 (N_199,N_160,In_465);
and U200 (N_200,In_427,N_134);
nor U201 (N_201,N_116,In_145);
nand U202 (N_202,N_144,N_176);
nor U203 (N_203,N_129,In_356);
and U204 (N_204,N_145,N_107);
or U205 (N_205,N_125,In_96);
or U206 (N_206,In_474,N_17);
nor U207 (N_207,N_76,In_470);
and U208 (N_208,In_165,N_49);
and U209 (N_209,N_140,N_66);
and U210 (N_210,In_45,In_211);
and U211 (N_211,N_87,In_5);
and U212 (N_212,N_120,In_214);
nand U213 (N_213,N_142,N_177);
and U214 (N_214,N_178,In_338);
and U215 (N_215,In_382,In_160);
nor U216 (N_216,In_159,N_10);
nor U217 (N_217,N_175,In_64);
nor U218 (N_218,N_67,N_31);
nor U219 (N_219,N_98,In_458);
nand U220 (N_220,N_112,In_183);
nand U221 (N_221,In_463,N_59);
and U222 (N_222,In_495,N_61);
nor U223 (N_223,In_421,N_84);
or U224 (N_224,In_6,In_487);
and U225 (N_225,N_136,N_164);
and U226 (N_226,N_69,N_179);
nand U227 (N_227,N_135,In_191);
and U228 (N_228,In_426,In_330);
nand U229 (N_229,N_127,In_230);
or U230 (N_230,In_171,N_62);
or U231 (N_231,In_444,In_381);
and U232 (N_232,In_394,In_112);
or U233 (N_233,N_46,In_75);
or U234 (N_234,N_126,N_83);
and U235 (N_235,N_9,N_118);
nand U236 (N_236,N_154,In_208);
nor U237 (N_237,N_86,N_157);
and U238 (N_238,In_482,In_366);
and U239 (N_239,In_9,N_79);
nor U240 (N_240,N_191,In_41);
nor U241 (N_241,In_108,In_254);
and U242 (N_242,N_198,In_248);
and U243 (N_243,In_479,In_274);
and U244 (N_244,In_358,In_219);
nand U245 (N_245,In_224,N_186);
nand U246 (N_246,N_218,In_462);
and U247 (N_247,N_216,N_213);
or U248 (N_248,In_399,N_148);
nor U249 (N_249,N_155,In_221);
nor U250 (N_250,In_116,N_26);
nand U251 (N_251,In_349,In_204);
nor U252 (N_252,N_223,In_324);
nand U253 (N_253,In_352,N_12);
nor U254 (N_254,N_156,In_139);
nand U255 (N_255,N_131,In_376);
and U256 (N_256,N_162,In_81);
or U257 (N_257,N_215,In_360);
nor U258 (N_258,N_68,N_210);
nor U259 (N_259,N_185,N_237);
or U260 (N_260,N_105,In_13);
or U261 (N_261,In_22,In_92);
nor U262 (N_262,In_89,N_227);
or U263 (N_263,In_141,In_348);
or U264 (N_264,N_77,In_434);
and U265 (N_265,N_6,N_28);
nand U266 (N_266,N_139,N_109);
or U267 (N_267,N_221,N_123);
nand U268 (N_268,N_110,In_238);
nor U269 (N_269,N_200,N_141);
nand U270 (N_270,In_289,In_261);
or U271 (N_271,N_203,N_174);
nor U272 (N_272,In_263,N_189);
or U273 (N_273,N_230,In_192);
nor U274 (N_274,N_151,In_436);
xor U275 (N_275,In_344,N_188);
and U276 (N_276,In_242,N_65);
nor U277 (N_277,In_162,N_196);
or U278 (N_278,In_121,In_212);
nand U279 (N_279,N_239,N_33);
or U280 (N_280,In_63,In_10);
or U281 (N_281,In_74,N_111);
nor U282 (N_282,In_468,N_209);
nor U283 (N_283,N_92,In_218);
nand U284 (N_284,N_171,N_5);
nor U285 (N_285,N_93,N_23);
and U286 (N_286,N_225,In_194);
xnor U287 (N_287,In_374,N_219);
nand U288 (N_288,In_464,N_130);
nor U289 (N_289,In_287,N_94);
nor U290 (N_290,In_83,N_54);
or U291 (N_291,In_207,In_93);
xor U292 (N_292,N_194,In_110);
xnor U293 (N_293,In_418,N_133);
and U294 (N_294,In_456,N_51);
nor U295 (N_295,In_488,In_332);
nand U296 (N_296,In_7,In_51);
or U297 (N_297,N_222,N_73);
nor U298 (N_298,N_3,N_1);
or U299 (N_299,In_411,N_199);
nor U300 (N_300,N_260,In_170);
nand U301 (N_301,N_172,In_87);
nand U302 (N_302,N_246,N_138);
nor U303 (N_303,N_217,In_193);
and U304 (N_304,N_241,In_266);
nand U305 (N_305,In_430,N_80);
nand U306 (N_306,N_190,N_279);
nor U307 (N_307,In_213,In_232);
and U308 (N_308,In_410,N_245);
nor U309 (N_309,N_182,N_290);
nand U310 (N_310,In_48,N_204);
and U311 (N_311,N_274,In_437);
nand U312 (N_312,N_150,N_261);
nand U313 (N_313,N_249,N_297);
nor U314 (N_314,N_4,N_238);
nand U315 (N_315,N_229,In_222);
nand U316 (N_316,N_235,In_378);
nor U317 (N_317,N_275,N_287);
or U318 (N_318,N_81,In_283);
nand U319 (N_319,N_27,N_272);
or U320 (N_320,N_273,N_159);
nand U321 (N_321,N_250,In_379);
or U322 (N_322,N_244,N_262);
nand U323 (N_323,In_343,N_234);
and U324 (N_324,N_146,N_153);
nand U325 (N_325,N_233,N_293);
nor U326 (N_326,N_14,N_294);
or U327 (N_327,In_31,N_242);
nor U328 (N_328,N_247,N_258);
nand U329 (N_329,N_282,N_103);
and U330 (N_330,In_76,N_266);
and U331 (N_331,N_267,N_231);
nor U332 (N_332,N_255,N_295);
nor U333 (N_333,N_251,N_170);
nor U334 (N_334,N_254,N_128);
nor U335 (N_335,N_240,N_207);
and U336 (N_336,In_17,N_212);
nand U337 (N_337,N_163,In_345);
and U338 (N_338,N_226,N_224);
nor U339 (N_339,In_143,N_286);
or U340 (N_340,In_124,N_276);
and U341 (N_341,N_232,N_248);
nand U342 (N_342,N_269,In_195);
nand U343 (N_343,In_119,N_180);
xnor U344 (N_344,N_202,In_27);
and U345 (N_345,N_166,N_64);
or U346 (N_346,In_351,In_217);
nor U347 (N_347,In_416,In_168);
and U348 (N_348,In_318,In_272);
or U349 (N_349,In_401,N_115);
nor U350 (N_350,In_18,N_289);
nor U351 (N_351,In_99,In_433);
nor U352 (N_352,In_357,N_291);
and U353 (N_353,N_270,N_256);
and U354 (N_354,N_82,In_282);
or U355 (N_355,In_1,N_284);
nor U356 (N_356,N_265,In_473);
nor U357 (N_357,N_104,In_60);
and U358 (N_358,N_271,N_263);
or U359 (N_359,N_280,N_158);
or U360 (N_360,In_37,N_327);
or U361 (N_361,N_315,N_352);
and U362 (N_362,N_205,N_313);
nor U363 (N_363,N_181,N_165);
xnor U364 (N_364,N_328,In_167);
nand U365 (N_365,N_357,N_220);
nor U366 (N_366,In_77,N_52);
nor U367 (N_367,N_321,N_43);
nand U368 (N_368,N_350,N_319);
nand U369 (N_369,N_332,N_345);
or U370 (N_370,N_193,N_149);
nor U371 (N_371,N_296,N_184);
nand U372 (N_372,N_102,N_337);
nand U373 (N_373,N_306,N_351);
nor U374 (N_374,In_452,N_302);
nand U375 (N_375,N_236,N_121);
nor U376 (N_376,N_341,N_309);
nor U377 (N_377,N_147,N_336);
and U378 (N_378,N_292,In_321);
and U379 (N_379,N_41,N_281);
nor U380 (N_380,In_161,N_11);
and U381 (N_381,N_96,N_299);
or U382 (N_382,In_177,N_322);
or U383 (N_383,In_297,N_333);
and U384 (N_384,In_188,N_97);
or U385 (N_385,N_307,N_316);
or U386 (N_386,N_268,N_342);
and U387 (N_387,In_56,N_168);
or U388 (N_388,N_298,In_383);
and U389 (N_389,N_303,N_320);
and U390 (N_390,N_201,N_183);
and U391 (N_391,N_101,N_325);
and U392 (N_392,N_278,In_423);
and U393 (N_393,N_344,N_192);
and U394 (N_394,N_308,N_169);
and U395 (N_395,In_228,N_348);
or U396 (N_396,N_330,N_161);
and U397 (N_397,In_422,In_329);
or U398 (N_398,N_253,N_326);
or U399 (N_399,N_277,N_323);
nor U400 (N_400,N_75,In_137);
nor U401 (N_401,N_24,N_304);
nand U402 (N_402,N_211,N_329);
nor U403 (N_403,N_346,In_377);
nand U404 (N_404,N_335,In_478);
nor U405 (N_405,N_358,N_318);
or U406 (N_406,N_288,N_324);
nand U407 (N_407,N_259,N_208);
nand U408 (N_408,N_257,N_300);
nand U409 (N_409,N_334,N_343);
and U410 (N_410,N_355,N_340);
nand U411 (N_411,N_206,N_197);
nand U412 (N_412,N_356,N_283);
or U413 (N_413,N_214,In_97);
and U414 (N_414,N_187,N_285);
nand U415 (N_415,N_117,N_359);
and U416 (N_416,N_243,In_154);
or U417 (N_417,N_312,In_123);
nor U418 (N_418,N_317,N_347);
nand U419 (N_419,N_339,N_99);
or U420 (N_420,N_264,N_353);
nand U421 (N_421,N_386,In_291);
or U422 (N_422,N_414,N_362);
or U423 (N_423,N_405,N_409);
and U424 (N_424,N_395,N_415);
and U425 (N_425,N_407,N_396);
nor U426 (N_426,N_367,N_314);
and U427 (N_427,N_416,N_417);
nand U428 (N_428,N_399,N_380);
and U429 (N_429,N_413,In_335);
and U430 (N_430,N_373,N_361);
xnor U431 (N_431,N_331,N_371);
or U432 (N_432,N_311,N_384);
nand U433 (N_433,N_377,N_385);
and U434 (N_434,N_419,N_349);
and U435 (N_435,N_389,N_390);
xor U436 (N_436,N_305,N_391);
nor U437 (N_437,N_388,N_408);
and U438 (N_438,N_406,N_364);
nor U439 (N_439,N_368,N_354);
or U440 (N_440,N_374,N_412);
nor U441 (N_441,N_372,N_418);
nor U442 (N_442,N_252,N_392);
or U443 (N_443,N_195,N_378);
nand U444 (N_444,N_56,N_310);
or U445 (N_445,N_394,In_225);
and U446 (N_446,N_398,N_370);
nand U447 (N_447,N_167,N_381);
and U448 (N_448,N_369,N_411);
nor U449 (N_449,N_387,N_403);
nor U450 (N_450,N_397,N_366);
or U451 (N_451,N_338,N_365);
or U452 (N_452,In_84,N_376);
nand U453 (N_453,N_360,N_393);
or U454 (N_454,N_379,N_410);
or U455 (N_455,N_382,N_375);
nand U456 (N_456,N_402,N_301);
nand U457 (N_457,N_401,N_404);
nor U458 (N_458,N_383,N_363);
nand U459 (N_459,N_400,N_228);
or U460 (N_460,N_408,N_363);
and U461 (N_461,N_365,N_419);
xnor U462 (N_462,N_56,N_388);
or U463 (N_463,In_225,N_399);
and U464 (N_464,N_392,N_408);
nand U465 (N_465,N_383,N_409);
nor U466 (N_466,N_362,N_374);
xor U467 (N_467,N_402,N_390);
nor U468 (N_468,N_407,N_390);
and U469 (N_469,In_84,N_366);
or U470 (N_470,N_354,N_399);
or U471 (N_471,N_305,N_367);
or U472 (N_472,N_398,N_404);
nand U473 (N_473,N_354,N_378);
or U474 (N_474,N_353,N_408);
nor U475 (N_475,N_395,N_410);
or U476 (N_476,N_228,N_384);
and U477 (N_477,N_410,N_397);
and U478 (N_478,N_375,In_291);
xor U479 (N_479,N_368,N_404);
nor U480 (N_480,N_439,N_445);
nor U481 (N_481,N_478,N_452);
or U482 (N_482,N_426,N_456);
nor U483 (N_483,N_435,N_475);
nand U484 (N_484,N_436,N_430);
and U485 (N_485,N_465,N_477);
or U486 (N_486,N_472,N_461);
nor U487 (N_487,N_425,N_454);
nor U488 (N_488,N_432,N_442);
and U489 (N_489,N_458,N_451);
nor U490 (N_490,N_438,N_453);
and U491 (N_491,N_447,N_473);
nand U492 (N_492,N_459,N_471);
and U493 (N_493,N_474,N_428);
or U494 (N_494,N_467,N_460);
nand U495 (N_495,N_427,N_464);
nand U496 (N_496,N_421,N_429);
or U497 (N_497,N_455,N_424);
or U498 (N_498,N_470,N_434);
or U499 (N_499,N_444,N_422);
or U500 (N_500,N_437,N_462);
or U501 (N_501,N_450,N_469);
nor U502 (N_502,N_433,N_448);
nand U503 (N_503,N_431,N_423);
or U504 (N_504,N_446,N_479);
and U505 (N_505,N_468,N_457);
and U506 (N_506,N_463,N_476);
or U507 (N_507,N_443,N_449);
and U508 (N_508,N_441,N_440);
nor U509 (N_509,N_420,N_466);
or U510 (N_510,N_474,N_420);
nand U511 (N_511,N_424,N_461);
and U512 (N_512,N_433,N_427);
nand U513 (N_513,N_463,N_457);
and U514 (N_514,N_454,N_449);
and U515 (N_515,N_473,N_479);
nand U516 (N_516,N_436,N_469);
and U517 (N_517,N_456,N_435);
nor U518 (N_518,N_429,N_424);
nand U519 (N_519,N_439,N_463);
nand U520 (N_520,N_449,N_450);
nor U521 (N_521,N_422,N_442);
nand U522 (N_522,N_430,N_420);
nor U523 (N_523,N_467,N_452);
or U524 (N_524,N_468,N_472);
or U525 (N_525,N_456,N_448);
nand U526 (N_526,N_464,N_426);
or U527 (N_527,N_449,N_455);
nand U528 (N_528,N_441,N_428);
nand U529 (N_529,N_473,N_429);
or U530 (N_530,N_450,N_435);
nor U531 (N_531,N_475,N_442);
nor U532 (N_532,N_432,N_440);
and U533 (N_533,N_470,N_427);
and U534 (N_534,N_421,N_450);
and U535 (N_535,N_435,N_425);
nand U536 (N_536,N_425,N_468);
nor U537 (N_537,N_460,N_436);
nand U538 (N_538,N_447,N_441);
or U539 (N_539,N_449,N_421);
nand U540 (N_540,N_488,N_531);
nor U541 (N_541,N_530,N_498);
xor U542 (N_542,N_482,N_483);
and U543 (N_543,N_526,N_532);
and U544 (N_544,N_512,N_481);
nand U545 (N_545,N_535,N_506);
nor U546 (N_546,N_492,N_520);
nor U547 (N_547,N_487,N_490);
nor U548 (N_548,N_523,N_484);
or U549 (N_549,N_534,N_521);
nand U550 (N_550,N_500,N_513);
nor U551 (N_551,N_486,N_511);
nand U552 (N_552,N_537,N_529);
nand U553 (N_553,N_491,N_517);
nand U554 (N_554,N_515,N_524);
and U555 (N_555,N_516,N_505);
or U556 (N_556,N_495,N_514);
nand U557 (N_557,N_527,N_518);
or U558 (N_558,N_502,N_519);
and U559 (N_559,N_489,N_494);
and U560 (N_560,N_493,N_480);
nor U561 (N_561,N_522,N_528);
or U562 (N_562,N_497,N_507);
or U563 (N_563,N_538,N_508);
nor U564 (N_564,N_510,N_496);
or U565 (N_565,N_501,N_533);
or U566 (N_566,N_539,N_525);
nor U567 (N_567,N_485,N_503);
or U568 (N_568,N_536,N_499);
nor U569 (N_569,N_509,N_504);
or U570 (N_570,N_484,N_502);
and U571 (N_571,N_517,N_509);
or U572 (N_572,N_528,N_525);
nor U573 (N_573,N_523,N_537);
nand U574 (N_574,N_486,N_490);
nand U575 (N_575,N_491,N_482);
or U576 (N_576,N_495,N_525);
nor U577 (N_577,N_529,N_527);
or U578 (N_578,N_499,N_492);
nand U579 (N_579,N_501,N_526);
or U580 (N_580,N_484,N_493);
nor U581 (N_581,N_520,N_538);
or U582 (N_582,N_514,N_491);
nor U583 (N_583,N_485,N_531);
nor U584 (N_584,N_511,N_514);
and U585 (N_585,N_509,N_503);
or U586 (N_586,N_526,N_508);
and U587 (N_587,N_502,N_493);
or U588 (N_588,N_480,N_525);
or U589 (N_589,N_508,N_481);
nand U590 (N_590,N_494,N_500);
and U591 (N_591,N_507,N_502);
or U592 (N_592,N_507,N_523);
nand U593 (N_593,N_539,N_489);
and U594 (N_594,N_515,N_521);
and U595 (N_595,N_488,N_503);
and U596 (N_596,N_537,N_484);
nor U597 (N_597,N_486,N_539);
or U598 (N_598,N_517,N_537);
nand U599 (N_599,N_537,N_528);
nor U600 (N_600,N_573,N_585);
xnor U601 (N_601,N_576,N_586);
or U602 (N_602,N_596,N_551);
nor U603 (N_603,N_577,N_574);
nand U604 (N_604,N_597,N_569);
or U605 (N_605,N_589,N_595);
nand U606 (N_606,N_555,N_571);
nor U607 (N_607,N_546,N_552);
nor U608 (N_608,N_547,N_590);
nor U609 (N_609,N_560,N_557);
and U610 (N_610,N_561,N_592);
nand U611 (N_611,N_562,N_564);
or U612 (N_612,N_565,N_588);
nand U613 (N_613,N_579,N_554);
and U614 (N_614,N_598,N_580);
nand U615 (N_615,N_541,N_578);
or U616 (N_616,N_545,N_542);
nor U617 (N_617,N_599,N_563);
or U618 (N_618,N_567,N_556);
nor U619 (N_619,N_575,N_543);
nand U620 (N_620,N_594,N_593);
and U621 (N_621,N_584,N_548);
and U622 (N_622,N_582,N_587);
and U623 (N_623,N_572,N_540);
and U624 (N_624,N_550,N_570);
xor U625 (N_625,N_549,N_568);
xor U626 (N_626,N_591,N_559);
nor U627 (N_627,N_553,N_583);
and U628 (N_628,N_581,N_566);
and U629 (N_629,N_558,N_544);
nand U630 (N_630,N_581,N_555);
nor U631 (N_631,N_584,N_599);
and U632 (N_632,N_569,N_545);
nor U633 (N_633,N_564,N_543);
nor U634 (N_634,N_551,N_570);
nor U635 (N_635,N_569,N_577);
nor U636 (N_636,N_542,N_550);
nor U637 (N_637,N_540,N_555);
and U638 (N_638,N_579,N_561);
nand U639 (N_639,N_547,N_571);
nor U640 (N_640,N_597,N_553);
or U641 (N_641,N_590,N_597);
nand U642 (N_642,N_593,N_567);
and U643 (N_643,N_552,N_567);
and U644 (N_644,N_584,N_568);
or U645 (N_645,N_579,N_596);
and U646 (N_646,N_593,N_597);
and U647 (N_647,N_589,N_573);
nor U648 (N_648,N_571,N_546);
nor U649 (N_649,N_594,N_591);
nor U650 (N_650,N_559,N_574);
or U651 (N_651,N_583,N_560);
or U652 (N_652,N_584,N_558);
nor U653 (N_653,N_561,N_585);
nand U654 (N_654,N_581,N_545);
xor U655 (N_655,N_599,N_552);
nand U656 (N_656,N_556,N_549);
nor U657 (N_657,N_566,N_549);
nand U658 (N_658,N_569,N_592);
or U659 (N_659,N_561,N_589);
nand U660 (N_660,N_654,N_659);
nor U661 (N_661,N_604,N_620);
nand U662 (N_662,N_614,N_610);
and U663 (N_663,N_602,N_658);
nor U664 (N_664,N_606,N_657);
nand U665 (N_665,N_626,N_618);
and U666 (N_666,N_638,N_632);
or U667 (N_667,N_649,N_648);
or U668 (N_668,N_643,N_612);
nand U669 (N_669,N_600,N_630);
and U670 (N_670,N_642,N_624);
nand U671 (N_671,N_652,N_631);
nand U672 (N_672,N_636,N_629);
nand U673 (N_673,N_627,N_635);
nor U674 (N_674,N_645,N_619);
nand U675 (N_675,N_605,N_653);
nor U676 (N_676,N_613,N_639);
or U677 (N_677,N_621,N_603);
nor U678 (N_678,N_608,N_601);
nand U679 (N_679,N_650,N_641);
xnor U680 (N_680,N_625,N_616);
and U681 (N_681,N_623,N_644);
nor U682 (N_682,N_651,N_633);
and U683 (N_683,N_611,N_609);
and U684 (N_684,N_655,N_637);
nand U685 (N_685,N_628,N_634);
nor U686 (N_686,N_646,N_622);
and U687 (N_687,N_615,N_607);
nor U688 (N_688,N_647,N_656);
nand U689 (N_689,N_640,N_617);
and U690 (N_690,N_602,N_653);
nand U691 (N_691,N_658,N_659);
or U692 (N_692,N_640,N_615);
or U693 (N_693,N_618,N_655);
and U694 (N_694,N_611,N_628);
and U695 (N_695,N_620,N_625);
nand U696 (N_696,N_605,N_601);
and U697 (N_697,N_619,N_601);
nand U698 (N_698,N_611,N_652);
nand U699 (N_699,N_645,N_607);
nor U700 (N_700,N_628,N_636);
nand U701 (N_701,N_600,N_619);
and U702 (N_702,N_650,N_632);
and U703 (N_703,N_630,N_620);
and U704 (N_704,N_621,N_657);
or U705 (N_705,N_620,N_611);
or U706 (N_706,N_653,N_647);
nor U707 (N_707,N_628,N_618);
nor U708 (N_708,N_651,N_645);
nand U709 (N_709,N_641,N_605);
or U710 (N_710,N_634,N_630);
or U711 (N_711,N_642,N_611);
nor U712 (N_712,N_633,N_621);
and U713 (N_713,N_633,N_638);
nor U714 (N_714,N_638,N_611);
nor U715 (N_715,N_651,N_600);
or U716 (N_716,N_615,N_646);
nor U717 (N_717,N_640,N_603);
nand U718 (N_718,N_619,N_648);
or U719 (N_719,N_649,N_626);
and U720 (N_720,N_710,N_690);
or U721 (N_721,N_700,N_713);
and U722 (N_722,N_687,N_684);
nand U723 (N_723,N_716,N_696);
nand U724 (N_724,N_667,N_685);
xor U725 (N_725,N_670,N_683);
nand U726 (N_726,N_679,N_707);
nand U727 (N_727,N_689,N_692);
nand U728 (N_728,N_676,N_662);
or U729 (N_729,N_715,N_708);
nand U730 (N_730,N_672,N_680);
or U731 (N_731,N_668,N_674);
nor U732 (N_732,N_704,N_686);
nor U733 (N_733,N_694,N_665);
nand U734 (N_734,N_666,N_705);
nand U735 (N_735,N_699,N_660);
nor U736 (N_736,N_703,N_664);
or U737 (N_737,N_673,N_663);
and U738 (N_738,N_718,N_669);
and U739 (N_739,N_671,N_677);
and U740 (N_740,N_693,N_717);
nand U741 (N_741,N_678,N_695);
or U742 (N_742,N_714,N_661);
and U743 (N_743,N_709,N_711);
nor U744 (N_744,N_697,N_681);
and U745 (N_745,N_698,N_675);
nand U746 (N_746,N_688,N_712);
and U747 (N_747,N_706,N_702);
nand U748 (N_748,N_701,N_682);
nand U749 (N_749,N_691,N_719);
and U750 (N_750,N_686,N_702);
xor U751 (N_751,N_664,N_690);
nand U752 (N_752,N_664,N_718);
xnor U753 (N_753,N_713,N_679);
and U754 (N_754,N_689,N_703);
nand U755 (N_755,N_661,N_692);
nor U756 (N_756,N_718,N_693);
nor U757 (N_757,N_683,N_675);
nand U758 (N_758,N_678,N_711);
and U759 (N_759,N_667,N_719);
nand U760 (N_760,N_716,N_691);
nand U761 (N_761,N_711,N_667);
nand U762 (N_762,N_715,N_718);
and U763 (N_763,N_713,N_705);
nor U764 (N_764,N_705,N_668);
nand U765 (N_765,N_682,N_702);
or U766 (N_766,N_668,N_667);
nand U767 (N_767,N_677,N_683);
nor U768 (N_768,N_698,N_709);
nand U769 (N_769,N_679,N_674);
nand U770 (N_770,N_706,N_683);
nand U771 (N_771,N_670,N_696);
nand U772 (N_772,N_694,N_711);
nand U773 (N_773,N_687,N_688);
nand U774 (N_774,N_685,N_671);
and U775 (N_775,N_680,N_707);
nor U776 (N_776,N_714,N_692);
and U777 (N_777,N_663,N_672);
nor U778 (N_778,N_675,N_708);
or U779 (N_779,N_673,N_711);
or U780 (N_780,N_730,N_771);
and U781 (N_781,N_731,N_740);
nand U782 (N_782,N_754,N_762);
and U783 (N_783,N_755,N_750);
or U784 (N_784,N_735,N_761);
nor U785 (N_785,N_778,N_747);
nand U786 (N_786,N_732,N_779);
nor U787 (N_787,N_739,N_727);
or U788 (N_788,N_721,N_737);
or U789 (N_789,N_758,N_752);
or U790 (N_790,N_734,N_733);
and U791 (N_791,N_769,N_720);
or U792 (N_792,N_741,N_772);
and U793 (N_793,N_728,N_773);
nor U794 (N_794,N_777,N_724);
or U795 (N_795,N_722,N_753);
nor U796 (N_796,N_723,N_757);
nor U797 (N_797,N_743,N_748);
nor U798 (N_798,N_756,N_742);
nor U799 (N_799,N_745,N_776);
nor U800 (N_800,N_770,N_746);
nor U801 (N_801,N_765,N_736);
and U802 (N_802,N_768,N_749);
nor U803 (N_803,N_775,N_759);
nor U804 (N_804,N_725,N_744);
nand U805 (N_805,N_774,N_763);
xnor U806 (N_806,N_760,N_767);
and U807 (N_807,N_729,N_751);
and U808 (N_808,N_726,N_738);
and U809 (N_809,N_766,N_764);
nor U810 (N_810,N_733,N_732);
nor U811 (N_811,N_727,N_763);
and U812 (N_812,N_741,N_748);
or U813 (N_813,N_720,N_779);
or U814 (N_814,N_775,N_764);
and U815 (N_815,N_732,N_773);
nor U816 (N_816,N_736,N_760);
nor U817 (N_817,N_726,N_746);
and U818 (N_818,N_779,N_729);
or U819 (N_819,N_750,N_763);
nor U820 (N_820,N_748,N_721);
and U821 (N_821,N_778,N_729);
or U822 (N_822,N_777,N_774);
or U823 (N_823,N_749,N_729);
or U824 (N_824,N_721,N_777);
or U825 (N_825,N_768,N_732);
nor U826 (N_826,N_722,N_765);
and U827 (N_827,N_738,N_763);
and U828 (N_828,N_726,N_768);
nor U829 (N_829,N_767,N_773);
and U830 (N_830,N_736,N_754);
nand U831 (N_831,N_722,N_764);
or U832 (N_832,N_775,N_744);
and U833 (N_833,N_773,N_763);
nor U834 (N_834,N_757,N_756);
or U835 (N_835,N_730,N_734);
or U836 (N_836,N_756,N_728);
or U837 (N_837,N_774,N_755);
nor U838 (N_838,N_727,N_753);
nand U839 (N_839,N_760,N_761);
nand U840 (N_840,N_817,N_812);
nor U841 (N_841,N_839,N_808);
or U842 (N_842,N_804,N_800);
nor U843 (N_843,N_823,N_786);
nand U844 (N_844,N_802,N_819);
and U845 (N_845,N_810,N_818);
or U846 (N_846,N_801,N_788);
or U847 (N_847,N_826,N_789);
nand U848 (N_848,N_797,N_781);
nand U849 (N_849,N_824,N_793);
or U850 (N_850,N_830,N_805);
and U851 (N_851,N_798,N_822);
or U852 (N_852,N_782,N_827);
or U853 (N_853,N_832,N_813);
nand U854 (N_854,N_785,N_799);
xnor U855 (N_855,N_831,N_790);
nand U856 (N_856,N_792,N_820);
nand U857 (N_857,N_807,N_821);
and U858 (N_858,N_829,N_783);
nor U859 (N_859,N_787,N_838);
and U860 (N_860,N_809,N_811);
nor U861 (N_861,N_828,N_796);
and U862 (N_862,N_834,N_836);
nand U863 (N_863,N_780,N_814);
and U864 (N_864,N_784,N_795);
nand U865 (N_865,N_835,N_816);
or U866 (N_866,N_833,N_791);
and U867 (N_867,N_837,N_803);
nand U868 (N_868,N_806,N_794);
nand U869 (N_869,N_825,N_815);
and U870 (N_870,N_798,N_800);
nand U871 (N_871,N_788,N_822);
nor U872 (N_872,N_827,N_836);
or U873 (N_873,N_792,N_827);
and U874 (N_874,N_811,N_795);
and U875 (N_875,N_811,N_818);
nor U876 (N_876,N_839,N_794);
nand U877 (N_877,N_791,N_836);
nand U878 (N_878,N_780,N_785);
nor U879 (N_879,N_798,N_791);
nand U880 (N_880,N_783,N_832);
nand U881 (N_881,N_795,N_786);
or U882 (N_882,N_796,N_835);
nor U883 (N_883,N_784,N_828);
nand U884 (N_884,N_807,N_801);
and U885 (N_885,N_837,N_814);
and U886 (N_886,N_791,N_816);
nand U887 (N_887,N_825,N_830);
nor U888 (N_888,N_812,N_790);
nor U889 (N_889,N_798,N_827);
and U890 (N_890,N_818,N_819);
or U891 (N_891,N_808,N_823);
nand U892 (N_892,N_801,N_799);
or U893 (N_893,N_823,N_838);
and U894 (N_894,N_813,N_806);
and U895 (N_895,N_784,N_791);
and U896 (N_896,N_815,N_796);
nand U897 (N_897,N_800,N_824);
or U898 (N_898,N_817,N_835);
nand U899 (N_899,N_828,N_804);
and U900 (N_900,N_869,N_859);
or U901 (N_901,N_873,N_872);
or U902 (N_902,N_898,N_890);
or U903 (N_903,N_861,N_896);
nand U904 (N_904,N_851,N_847);
and U905 (N_905,N_886,N_850);
nor U906 (N_906,N_860,N_874);
nand U907 (N_907,N_866,N_846);
or U908 (N_908,N_867,N_843);
nand U909 (N_909,N_871,N_855);
or U910 (N_910,N_875,N_852);
nand U911 (N_911,N_856,N_889);
or U912 (N_912,N_840,N_897);
or U913 (N_913,N_877,N_862);
nand U914 (N_914,N_891,N_882);
and U915 (N_915,N_881,N_854);
nor U916 (N_916,N_879,N_878);
and U917 (N_917,N_849,N_895);
nor U918 (N_918,N_893,N_865);
or U919 (N_919,N_899,N_863);
nor U920 (N_920,N_876,N_845);
nor U921 (N_921,N_864,N_884);
xnor U922 (N_922,N_842,N_892);
nand U923 (N_923,N_880,N_887);
nor U924 (N_924,N_858,N_885);
nand U925 (N_925,N_868,N_844);
or U926 (N_926,N_870,N_857);
and U927 (N_927,N_883,N_853);
or U928 (N_928,N_841,N_888);
nand U929 (N_929,N_848,N_894);
or U930 (N_930,N_887,N_892);
nand U931 (N_931,N_871,N_848);
nand U932 (N_932,N_887,N_876);
nand U933 (N_933,N_850,N_856);
nor U934 (N_934,N_866,N_840);
and U935 (N_935,N_855,N_848);
nand U936 (N_936,N_896,N_892);
and U937 (N_937,N_870,N_841);
and U938 (N_938,N_852,N_854);
nand U939 (N_939,N_851,N_877);
xnor U940 (N_940,N_849,N_857);
and U941 (N_941,N_861,N_850);
nand U942 (N_942,N_856,N_847);
nor U943 (N_943,N_858,N_870);
nor U944 (N_944,N_882,N_889);
nor U945 (N_945,N_880,N_858);
nand U946 (N_946,N_850,N_878);
or U947 (N_947,N_867,N_893);
or U948 (N_948,N_848,N_844);
or U949 (N_949,N_846,N_878);
and U950 (N_950,N_879,N_886);
or U951 (N_951,N_869,N_856);
nand U952 (N_952,N_881,N_867);
nor U953 (N_953,N_897,N_855);
nand U954 (N_954,N_867,N_879);
and U955 (N_955,N_896,N_884);
and U956 (N_956,N_846,N_889);
nor U957 (N_957,N_884,N_889);
nor U958 (N_958,N_850,N_873);
nor U959 (N_959,N_884,N_897);
and U960 (N_960,N_934,N_904);
nor U961 (N_961,N_901,N_949);
or U962 (N_962,N_935,N_933);
nand U963 (N_963,N_918,N_915);
or U964 (N_964,N_948,N_939);
nor U965 (N_965,N_911,N_947);
nand U966 (N_966,N_914,N_945);
and U967 (N_967,N_926,N_946);
xor U968 (N_968,N_936,N_923);
or U969 (N_969,N_957,N_919);
nor U970 (N_970,N_951,N_913);
and U971 (N_971,N_925,N_944);
nor U972 (N_972,N_921,N_910);
or U973 (N_973,N_912,N_937);
nor U974 (N_974,N_930,N_909);
and U975 (N_975,N_954,N_941);
nand U976 (N_976,N_943,N_942);
and U977 (N_977,N_924,N_906);
or U978 (N_978,N_952,N_905);
nor U979 (N_979,N_916,N_928);
xor U980 (N_980,N_922,N_953);
xor U981 (N_981,N_920,N_900);
nand U982 (N_982,N_927,N_903);
nor U983 (N_983,N_956,N_959);
and U984 (N_984,N_955,N_902);
or U985 (N_985,N_938,N_917);
nor U986 (N_986,N_950,N_958);
or U987 (N_987,N_940,N_932);
or U988 (N_988,N_908,N_907);
nor U989 (N_989,N_931,N_929);
or U990 (N_990,N_924,N_950);
nand U991 (N_991,N_915,N_927);
nand U992 (N_992,N_915,N_933);
nor U993 (N_993,N_906,N_905);
and U994 (N_994,N_956,N_936);
or U995 (N_995,N_940,N_915);
or U996 (N_996,N_918,N_905);
or U997 (N_997,N_926,N_945);
nand U998 (N_998,N_929,N_941);
and U999 (N_999,N_953,N_900);
nor U1000 (N_1000,N_940,N_943);
and U1001 (N_1001,N_937,N_923);
and U1002 (N_1002,N_948,N_958);
nor U1003 (N_1003,N_924,N_943);
nand U1004 (N_1004,N_900,N_950);
or U1005 (N_1005,N_903,N_947);
or U1006 (N_1006,N_929,N_922);
nor U1007 (N_1007,N_901,N_914);
xnor U1008 (N_1008,N_957,N_904);
and U1009 (N_1009,N_928,N_932);
nand U1010 (N_1010,N_954,N_915);
nor U1011 (N_1011,N_905,N_941);
nor U1012 (N_1012,N_910,N_912);
and U1013 (N_1013,N_945,N_927);
nand U1014 (N_1014,N_922,N_926);
nor U1015 (N_1015,N_914,N_942);
nor U1016 (N_1016,N_914,N_958);
and U1017 (N_1017,N_950,N_920);
nor U1018 (N_1018,N_921,N_955);
and U1019 (N_1019,N_904,N_951);
nand U1020 (N_1020,N_968,N_1004);
or U1021 (N_1021,N_999,N_1011);
or U1022 (N_1022,N_1009,N_992);
or U1023 (N_1023,N_964,N_965);
nand U1024 (N_1024,N_981,N_983);
nor U1025 (N_1025,N_989,N_963);
and U1026 (N_1026,N_1007,N_994);
or U1027 (N_1027,N_1019,N_966);
nand U1028 (N_1028,N_1001,N_961);
or U1029 (N_1029,N_974,N_976);
or U1030 (N_1030,N_1003,N_1015);
nor U1031 (N_1031,N_967,N_986);
nor U1032 (N_1032,N_1002,N_998);
and U1033 (N_1033,N_996,N_1000);
or U1034 (N_1034,N_1014,N_969);
nand U1035 (N_1035,N_970,N_1006);
or U1036 (N_1036,N_987,N_977);
and U1037 (N_1037,N_962,N_985);
nand U1038 (N_1038,N_978,N_971);
nor U1039 (N_1039,N_1005,N_979);
and U1040 (N_1040,N_982,N_995);
nor U1041 (N_1041,N_1017,N_1012);
nand U1042 (N_1042,N_980,N_988);
nand U1043 (N_1043,N_1018,N_1013);
xnor U1044 (N_1044,N_1016,N_993);
nor U1045 (N_1045,N_990,N_1008);
or U1046 (N_1046,N_1010,N_991);
nand U1047 (N_1047,N_960,N_975);
nor U1048 (N_1048,N_973,N_997);
or U1049 (N_1049,N_984,N_972);
or U1050 (N_1050,N_963,N_982);
nor U1051 (N_1051,N_1014,N_1005);
or U1052 (N_1052,N_960,N_963);
nand U1053 (N_1053,N_974,N_975);
or U1054 (N_1054,N_961,N_998);
or U1055 (N_1055,N_999,N_1010);
nand U1056 (N_1056,N_976,N_965);
nor U1057 (N_1057,N_1002,N_972);
xor U1058 (N_1058,N_966,N_969);
and U1059 (N_1059,N_965,N_963);
or U1060 (N_1060,N_969,N_1011);
nor U1061 (N_1061,N_1009,N_1014);
nand U1062 (N_1062,N_964,N_1008);
xor U1063 (N_1063,N_995,N_996);
or U1064 (N_1064,N_1014,N_985);
nor U1065 (N_1065,N_1018,N_984);
or U1066 (N_1066,N_968,N_1017);
and U1067 (N_1067,N_1012,N_1019);
nand U1068 (N_1068,N_964,N_980);
nor U1069 (N_1069,N_1002,N_980);
and U1070 (N_1070,N_989,N_988);
nor U1071 (N_1071,N_1008,N_993);
or U1072 (N_1072,N_1018,N_1008);
or U1073 (N_1073,N_972,N_997);
or U1074 (N_1074,N_1008,N_1002);
and U1075 (N_1075,N_990,N_1016);
nor U1076 (N_1076,N_1017,N_1004);
nand U1077 (N_1077,N_1013,N_961);
or U1078 (N_1078,N_973,N_991);
and U1079 (N_1079,N_982,N_992);
and U1080 (N_1080,N_1042,N_1061);
or U1081 (N_1081,N_1062,N_1064);
nand U1082 (N_1082,N_1053,N_1076);
and U1083 (N_1083,N_1045,N_1040);
or U1084 (N_1084,N_1072,N_1033);
nor U1085 (N_1085,N_1070,N_1059);
or U1086 (N_1086,N_1071,N_1065);
and U1087 (N_1087,N_1074,N_1060);
or U1088 (N_1088,N_1063,N_1020);
nor U1089 (N_1089,N_1024,N_1075);
and U1090 (N_1090,N_1077,N_1030);
nand U1091 (N_1091,N_1044,N_1058);
nand U1092 (N_1092,N_1029,N_1027);
and U1093 (N_1093,N_1022,N_1069);
and U1094 (N_1094,N_1057,N_1026);
nor U1095 (N_1095,N_1025,N_1036);
nand U1096 (N_1096,N_1037,N_1031);
nor U1097 (N_1097,N_1047,N_1043);
nor U1098 (N_1098,N_1052,N_1054);
nand U1099 (N_1099,N_1023,N_1041);
and U1100 (N_1100,N_1034,N_1021);
and U1101 (N_1101,N_1051,N_1032);
or U1102 (N_1102,N_1028,N_1035);
nor U1103 (N_1103,N_1046,N_1078);
or U1104 (N_1104,N_1068,N_1073);
or U1105 (N_1105,N_1067,N_1049);
xor U1106 (N_1106,N_1066,N_1039);
and U1107 (N_1107,N_1055,N_1056);
nor U1108 (N_1108,N_1048,N_1038);
or U1109 (N_1109,N_1050,N_1079);
nor U1110 (N_1110,N_1036,N_1049);
or U1111 (N_1111,N_1028,N_1032);
nand U1112 (N_1112,N_1033,N_1078);
nor U1113 (N_1113,N_1065,N_1037);
and U1114 (N_1114,N_1074,N_1064);
nor U1115 (N_1115,N_1048,N_1044);
and U1116 (N_1116,N_1033,N_1062);
or U1117 (N_1117,N_1038,N_1033);
xor U1118 (N_1118,N_1054,N_1035);
and U1119 (N_1119,N_1051,N_1044);
nand U1120 (N_1120,N_1032,N_1061);
or U1121 (N_1121,N_1030,N_1024);
or U1122 (N_1122,N_1052,N_1063);
and U1123 (N_1123,N_1064,N_1076);
nand U1124 (N_1124,N_1060,N_1034);
xnor U1125 (N_1125,N_1061,N_1064);
nand U1126 (N_1126,N_1079,N_1074);
or U1127 (N_1127,N_1029,N_1064);
nor U1128 (N_1128,N_1024,N_1022);
nor U1129 (N_1129,N_1064,N_1035);
or U1130 (N_1130,N_1055,N_1022);
nand U1131 (N_1131,N_1028,N_1053);
or U1132 (N_1132,N_1072,N_1029);
nand U1133 (N_1133,N_1075,N_1029);
nor U1134 (N_1134,N_1057,N_1042);
nor U1135 (N_1135,N_1059,N_1074);
and U1136 (N_1136,N_1046,N_1069);
nand U1137 (N_1137,N_1056,N_1043);
and U1138 (N_1138,N_1027,N_1061);
nor U1139 (N_1139,N_1043,N_1076);
or U1140 (N_1140,N_1105,N_1117);
nor U1141 (N_1141,N_1139,N_1138);
nor U1142 (N_1142,N_1125,N_1135);
and U1143 (N_1143,N_1100,N_1095);
and U1144 (N_1144,N_1103,N_1092);
nor U1145 (N_1145,N_1093,N_1082);
nor U1146 (N_1146,N_1124,N_1118);
and U1147 (N_1147,N_1097,N_1119);
or U1148 (N_1148,N_1113,N_1123);
or U1149 (N_1149,N_1112,N_1104);
and U1150 (N_1150,N_1107,N_1130);
or U1151 (N_1151,N_1090,N_1127);
and U1152 (N_1152,N_1106,N_1120);
xor U1153 (N_1153,N_1129,N_1116);
nor U1154 (N_1154,N_1083,N_1088);
nor U1155 (N_1155,N_1101,N_1084);
or U1156 (N_1156,N_1108,N_1137);
nor U1157 (N_1157,N_1121,N_1098);
nor U1158 (N_1158,N_1128,N_1081);
nor U1159 (N_1159,N_1114,N_1109);
or U1160 (N_1160,N_1131,N_1085);
and U1161 (N_1161,N_1122,N_1102);
or U1162 (N_1162,N_1111,N_1132);
nand U1163 (N_1163,N_1087,N_1089);
nor U1164 (N_1164,N_1115,N_1136);
or U1165 (N_1165,N_1096,N_1080);
and U1166 (N_1166,N_1133,N_1094);
and U1167 (N_1167,N_1126,N_1134);
or U1168 (N_1168,N_1091,N_1110);
nand U1169 (N_1169,N_1099,N_1086);
or U1170 (N_1170,N_1108,N_1133);
nor U1171 (N_1171,N_1131,N_1092);
and U1172 (N_1172,N_1099,N_1118);
or U1173 (N_1173,N_1137,N_1094);
or U1174 (N_1174,N_1093,N_1089);
and U1175 (N_1175,N_1099,N_1130);
and U1176 (N_1176,N_1097,N_1100);
and U1177 (N_1177,N_1135,N_1097);
nand U1178 (N_1178,N_1127,N_1134);
nor U1179 (N_1179,N_1106,N_1136);
nand U1180 (N_1180,N_1116,N_1132);
nand U1181 (N_1181,N_1100,N_1112);
nor U1182 (N_1182,N_1118,N_1103);
and U1183 (N_1183,N_1095,N_1101);
nand U1184 (N_1184,N_1108,N_1117);
or U1185 (N_1185,N_1090,N_1102);
nor U1186 (N_1186,N_1080,N_1105);
and U1187 (N_1187,N_1115,N_1116);
or U1188 (N_1188,N_1090,N_1110);
or U1189 (N_1189,N_1110,N_1120);
nand U1190 (N_1190,N_1137,N_1132);
or U1191 (N_1191,N_1098,N_1085);
or U1192 (N_1192,N_1096,N_1130);
nor U1193 (N_1193,N_1112,N_1136);
and U1194 (N_1194,N_1109,N_1089);
or U1195 (N_1195,N_1124,N_1139);
nor U1196 (N_1196,N_1097,N_1109);
and U1197 (N_1197,N_1098,N_1129);
nor U1198 (N_1198,N_1088,N_1080);
and U1199 (N_1199,N_1114,N_1101);
nor U1200 (N_1200,N_1165,N_1155);
or U1201 (N_1201,N_1148,N_1140);
nand U1202 (N_1202,N_1183,N_1167);
and U1203 (N_1203,N_1141,N_1196);
and U1204 (N_1204,N_1195,N_1170);
nand U1205 (N_1205,N_1144,N_1166);
nor U1206 (N_1206,N_1176,N_1178);
nand U1207 (N_1207,N_1186,N_1162);
and U1208 (N_1208,N_1145,N_1184);
or U1209 (N_1209,N_1173,N_1197);
nand U1210 (N_1210,N_1181,N_1163);
and U1211 (N_1211,N_1193,N_1191);
or U1212 (N_1212,N_1168,N_1199);
nand U1213 (N_1213,N_1158,N_1151);
nand U1214 (N_1214,N_1152,N_1142);
or U1215 (N_1215,N_1194,N_1171);
nand U1216 (N_1216,N_1179,N_1192);
nor U1217 (N_1217,N_1182,N_1177);
and U1218 (N_1218,N_1180,N_1147);
and U1219 (N_1219,N_1185,N_1175);
nand U1220 (N_1220,N_1160,N_1164);
nand U1221 (N_1221,N_1174,N_1156);
and U1222 (N_1222,N_1150,N_1146);
and U1223 (N_1223,N_1172,N_1157);
nand U1224 (N_1224,N_1149,N_1161);
nor U1225 (N_1225,N_1188,N_1153);
and U1226 (N_1226,N_1159,N_1187);
nand U1227 (N_1227,N_1189,N_1143);
and U1228 (N_1228,N_1198,N_1190);
and U1229 (N_1229,N_1169,N_1154);
nor U1230 (N_1230,N_1186,N_1189);
nor U1231 (N_1231,N_1151,N_1145);
or U1232 (N_1232,N_1195,N_1173);
or U1233 (N_1233,N_1162,N_1152);
or U1234 (N_1234,N_1165,N_1192);
nor U1235 (N_1235,N_1190,N_1199);
xnor U1236 (N_1236,N_1143,N_1177);
or U1237 (N_1237,N_1184,N_1152);
nand U1238 (N_1238,N_1154,N_1146);
nor U1239 (N_1239,N_1189,N_1188);
nor U1240 (N_1240,N_1175,N_1156);
or U1241 (N_1241,N_1174,N_1185);
or U1242 (N_1242,N_1172,N_1184);
or U1243 (N_1243,N_1152,N_1156);
nand U1244 (N_1244,N_1193,N_1173);
and U1245 (N_1245,N_1178,N_1197);
nand U1246 (N_1246,N_1141,N_1182);
or U1247 (N_1247,N_1180,N_1175);
nor U1248 (N_1248,N_1193,N_1163);
nor U1249 (N_1249,N_1153,N_1154);
or U1250 (N_1250,N_1165,N_1145);
nor U1251 (N_1251,N_1191,N_1197);
nand U1252 (N_1252,N_1183,N_1146);
nor U1253 (N_1253,N_1182,N_1158);
or U1254 (N_1254,N_1145,N_1154);
nor U1255 (N_1255,N_1160,N_1177);
and U1256 (N_1256,N_1187,N_1161);
or U1257 (N_1257,N_1144,N_1183);
or U1258 (N_1258,N_1155,N_1183);
nand U1259 (N_1259,N_1188,N_1192);
nor U1260 (N_1260,N_1231,N_1244);
xor U1261 (N_1261,N_1224,N_1241);
and U1262 (N_1262,N_1201,N_1233);
and U1263 (N_1263,N_1254,N_1226);
or U1264 (N_1264,N_1242,N_1210);
nor U1265 (N_1265,N_1209,N_1225);
nand U1266 (N_1266,N_1248,N_1255);
nor U1267 (N_1267,N_1216,N_1202);
xnor U1268 (N_1268,N_1221,N_1227);
nand U1269 (N_1269,N_1200,N_1211);
nor U1270 (N_1270,N_1240,N_1203);
nor U1271 (N_1271,N_1218,N_1229);
or U1272 (N_1272,N_1230,N_1258);
or U1273 (N_1273,N_1236,N_1213);
nor U1274 (N_1274,N_1235,N_1219);
nor U1275 (N_1275,N_1232,N_1252);
nand U1276 (N_1276,N_1206,N_1238);
and U1277 (N_1277,N_1212,N_1204);
or U1278 (N_1278,N_1253,N_1228);
nand U1279 (N_1279,N_1246,N_1251);
and U1280 (N_1280,N_1239,N_1205);
nor U1281 (N_1281,N_1259,N_1256);
nor U1282 (N_1282,N_1208,N_1249);
or U1283 (N_1283,N_1214,N_1215);
and U1284 (N_1284,N_1247,N_1237);
and U1285 (N_1285,N_1223,N_1234);
or U1286 (N_1286,N_1250,N_1243);
and U1287 (N_1287,N_1207,N_1257);
or U1288 (N_1288,N_1217,N_1222);
or U1289 (N_1289,N_1220,N_1245);
nor U1290 (N_1290,N_1223,N_1241);
or U1291 (N_1291,N_1241,N_1214);
or U1292 (N_1292,N_1252,N_1214);
nand U1293 (N_1293,N_1201,N_1208);
nand U1294 (N_1294,N_1229,N_1220);
or U1295 (N_1295,N_1213,N_1231);
and U1296 (N_1296,N_1246,N_1255);
nor U1297 (N_1297,N_1256,N_1230);
and U1298 (N_1298,N_1206,N_1218);
and U1299 (N_1299,N_1241,N_1218);
and U1300 (N_1300,N_1244,N_1226);
and U1301 (N_1301,N_1208,N_1248);
and U1302 (N_1302,N_1226,N_1255);
nor U1303 (N_1303,N_1227,N_1239);
or U1304 (N_1304,N_1222,N_1208);
nand U1305 (N_1305,N_1233,N_1227);
or U1306 (N_1306,N_1215,N_1233);
and U1307 (N_1307,N_1234,N_1250);
or U1308 (N_1308,N_1225,N_1244);
and U1309 (N_1309,N_1243,N_1236);
or U1310 (N_1310,N_1214,N_1235);
nor U1311 (N_1311,N_1209,N_1226);
and U1312 (N_1312,N_1247,N_1241);
or U1313 (N_1313,N_1256,N_1251);
and U1314 (N_1314,N_1207,N_1223);
nand U1315 (N_1315,N_1230,N_1225);
xnor U1316 (N_1316,N_1230,N_1245);
or U1317 (N_1317,N_1233,N_1252);
nand U1318 (N_1318,N_1212,N_1205);
nand U1319 (N_1319,N_1234,N_1257);
nand U1320 (N_1320,N_1271,N_1278);
and U1321 (N_1321,N_1296,N_1314);
nand U1322 (N_1322,N_1313,N_1301);
or U1323 (N_1323,N_1309,N_1269);
and U1324 (N_1324,N_1290,N_1306);
and U1325 (N_1325,N_1293,N_1265);
nand U1326 (N_1326,N_1274,N_1282);
or U1327 (N_1327,N_1304,N_1312);
nor U1328 (N_1328,N_1267,N_1268);
and U1329 (N_1329,N_1273,N_1264);
nor U1330 (N_1330,N_1275,N_1310);
nand U1331 (N_1331,N_1300,N_1302);
nand U1332 (N_1332,N_1308,N_1298);
and U1333 (N_1333,N_1279,N_1283);
or U1334 (N_1334,N_1292,N_1263);
nand U1335 (N_1335,N_1291,N_1277);
and U1336 (N_1336,N_1288,N_1311);
nand U1337 (N_1337,N_1295,N_1272);
nor U1338 (N_1338,N_1270,N_1260);
xor U1339 (N_1339,N_1266,N_1294);
nor U1340 (N_1340,N_1287,N_1297);
and U1341 (N_1341,N_1285,N_1276);
and U1342 (N_1342,N_1316,N_1317);
or U1343 (N_1343,N_1303,N_1281);
nand U1344 (N_1344,N_1318,N_1299);
nor U1345 (N_1345,N_1261,N_1305);
nor U1346 (N_1346,N_1319,N_1284);
or U1347 (N_1347,N_1315,N_1289);
or U1348 (N_1348,N_1262,N_1286);
nor U1349 (N_1349,N_1280,N_1307);
or U1350 (N_1350,N_1271,N_1314);
and U1351 (N_1351,N_1270,N_1316);
xnor U1352 (N_1352,N_1307,N_1313);
and U1353 (N_1353,N_1295,N_1294);
nor U1354 (N_1354,N_1270,N_1303);
and U1355 (N_1355,N_1301,N_1307);
nor U1356 (N_1356,N_1266,N_1316);
or U1357 (N_1357,N_1266,N_1295);
and U1358 (N_1358,N_1292,N_1306);
and U1359 (N_1359,N_1291,N_1274);
and U1360 (N_1360,N_1270,N_1276);
or U1361 (N_1361,N_1280,N_1317);
or U1362 (N_1362,N_1306,N_1264);
or U1363 (N_1363,N_1309,N_1312);
and U1364 (N_1364,N_1319,N_1294);
and U1365 (N_1365,N_1264,N_1272);
and U1366 (N_1366,N_1296,N_1290);
and U1367 (N_1367,N_1297,N_1307);
nand U1368 (N_1368,N_1300,N_1280);
nor U1369 (N_1369,N_1319,N_1305);
nand U1370 (N_1370,N_1276,N_1279);
or U1371 (N_1371,N_1295,N_1319);
nand U1372 (N_1372,N_1295,N_1307);
nor U1373 (N_1373,N_1309,N_1291);
and U1374 (N_1374,N_1297,N_1266);
and U1375 (N_1375,N_1293,N_1303);
nand U1376 (N_1376,N_1318,N_1312);
nor U1377 (N_1377,N_1295,N_1270);
or U1378 (N_1378,N_1312,N_1294);
and U1379 (N_1379,N_1291,N_1295);
and U1380 (N_1380,N_1357,N_1378);
and U1381 (N_1381,N_1363,N_1328);
and U1382 (N_1382,N_1375,N_1359);
nand U1383 (N_1383,N_1331,N_1338);
nand U1384 (N_1384,N_1335,N_1372);
and U1385 (N_1385,N_1368,N_1330);
nand U1386 (N_1386,N_1370,N_1358);
or U1387 (N_1387,N_1348,N_1326);
nand U1388 (N_1388,N_1329,N_1356);
nand U1389 (N_1389,N_1340,N_1325);
nor U1390 (N_1390,N_1322,N_1367);
or U1391 (N_1391,N_1349,N_1361);
and U1392 (N_1392,N_1353,N_1341);
or U1393 (N_1393,N_1339,N_1327);
and U1394 (N_1394,N_1351,N_1343);
nand U1395 (N_1395,N_1334,N_1323);
nor U1396 (N_1396,N_1379,N_1354);
nand U1397 (N_1397,N_1369,N_1352);
or U1398 (N_1398,N_1362,N_1360);
and U1399 (N_1399,N_1344,N_1333);
xnor U1400 (N_1400,N_1365,N_1366);
nand U1401 (N_1401,N_1324,N_1345);
or U1402 (N_1402,N_1355,N_1332);
nor U1403 (N_1403,N_1336,N_1364);
and U1404 (N_1404,N_1376,N_1373);
xor U1405 (N_1405,N_1337,N_1320);
nand U1406 (N_1406,N_1374,N_1347);
nand U1407 (N_1407,N_1377,N_1342);
and U1408 (N_1408,N_1321,N_1346);
or U1409 (N_1409,N_1350,N_1371);
nand U1410 (N_1410,N_1355,N_1379);
nand U1411 (N_1411,N_1360,N_1340);
nand U1412 (N_1412,N_1347,N_1345);
nor U1413 (N_1413,N_1349,N_1324);
nand U1414 (N_1414,N_1320,N_1326);
and U1415 (N_1415,N_1341,N_1337);
nand U1416 (N_1416,N_1378,N_1365);
and U1417 (N_1417,N_1358,N_1321);
and U1418 (N_1418,N_1320,N_1343);
nand U1419 (N_1419,N_1349,N_1373);
and U1420 (N_1420,N_1347,N_1331);
nand U1421 (N_1421,N_1349,N_1366);
or U1422 (N_1422,N_1336,N_1329);
nor U1423 (N_1423,N_1322,N_1337);
nand U1424 (N_1424,N_1379,N_1378);
or U1425 (N_1425,N_1346,N_1347);
or U1426 (N_1426,N_1338,N_1323);
xnor U1427 (N_1427,N_1360,N_1354);
or U1428 (N_1428,N_1376,N_1343);
nor U1429 (N_1429,N_1349,N_1343);
or U1430 (N_1430,N_1371,N_1347);
nand U1431 (N_1431,N_1332,N_1374);
and U1432 (N_1432,N_1359,N_1349);
nor U1433 (N_1433,N_1325,N_1324);
and U1434 (N_1434,N_1378,N_1356);
and U1435 (N_1435,N_1333,N_1377);
nor U1436 (N_1436,N_1349,N_1371);
nand U1437 (N_1437,N_1321,N_1351);
or U1438 (N_1438,N_1378,N_1376);
nor U1439 (N_1439,N_1326,N_1372);
xor U1440 (N_1440,N_1403,N_1386);
or U1441 (N_1441,N_1389,N_1427);
nand U1442 (N_1442,N_1400,N_1384);
and U1443 (N_1443,N_1430,N_1435);
and U1444 (N_1444,N_1397,N_1438);
and U1445 (N_1445,N_1422,N_1396);
nand U1446 (N_1446,N_1417,N_1433);
nand U1447 (N_1447,N_1434,N_1405);
or U1448 (N_1448,N_1410,N_1426);
xnor U1449 (N_1449,N_1391,N_1431);
nand U1450 (N_1450,N_1432,N_1413);
nand U1451 (N_1451,N_1388,N_1392);
or U1452 (N_1452,N_1423,N_1424);
nand U1453 (N_1453,N_1383,N_1412);
or U1454 (N_1454,N_1420,N_1429);
nand U1455 (N_1455,N_1439,N_1382);
nor U1456 (N_1456,N_1404,N_1406);
and U1457 (N_1457,N_1402,N_1387);
nand U1458 (N_1458,N_1428,N_1411);
and U1459 (N_1459,N_1415,N_1398);
or U1460 (N_1460,N_1385,N_1401);
xor U1461 (N_1461,N_1380,N_1414);
and U1462 (N_1462,N_1425,N_1437);
nor U1463 (N_1463,N_1407,N_1409);
nand U1464 (N_1464,N_1419,N_1421);
nor U1465 (N_1465,N_1399,N_1390);
nand U1466 (N_1466,N_1418,N_1408);
and U1467 (N_1467,N_1416,N_1395);
nand U1468 (N_1468,N_1393,N_1381);
or U1469 (N_1469,N_1436,N_1394);
and U1470 (N_1470,N_1402,N_1412);
nor U1471 (N_1471,N_1427,N_1437);
and U1472 (N_1472,N_1412,N_1429);
or U1473 (N_1473,N_1431,N_1424);
nor U1474 (N_1474,N_1408,N_1415);
nand U1475 (N_1475,N_1427,N_1388);
nor U1476 (N_1476,N_1432,N_1414);
nand U1477 (N_1477,N_1427,N_1383);
nand U1478 (N_1478,N_1430,N_1439);
xor U1479 (N_1479,N_1422,N_1400);
or U1480 (N_1480,N_1422,N_1417);
nand U1481 (N_1481,N_1417,N_1395);
nor U1482 (N_1482,N_1383,N_1408);
nand U1483 (N_1483,N_1412,N_1394);
nand U1484 (N_1484,N_1388,N_1389);
and U1485 (N_1485,N_1422,N_1413);
nand U1486 (N_1486,N_1418,N_1411);
nor U1487 (N_1487,N_1392,N_1409);
and U1488 (N_1488,N_1435,N_1399);
or U1489 (N_1489,N_1403,N_1411);
or U1490 (N_1490,N_1385,N_1391);
nor U1491 (N_1491,N_1390,N_1431);
or U1492 (N_1492,N_1414,N_1410);
or U1493 (N_1493,N_1389,N_1415);
nand U1494 (N_1494,N_1402,N_1383);
nand U1495 (N_1495,N_1434,N_1407);
nand U1496 (N_1496,N_1421,N_1433);
nand U1497 (N_1497,N_1402,N_1398);
and U1498 (N_1498,N_1382,N_1402);
nor U1499 (N_1499,N_1434,N_1384);
nor U1500 (N_1500,N_1466,N_1475);
nand U1501 (N_1501,N_1477,N_1463);
and U1502 (N_1502,N_1479,N_1489);
and U1503 (N_1503,N_1495,N_1481);
xor U1504 (N_1504,N_1488,N_1451);
nor U1505 (N_1505,N_1453,N_1450);
nand U1506 (N_1506,N_1473,N_1491);
nand U1507 (N_1507,N_1483,N_1458);
nor U1508 (N_1508,N_1442,N_1460);
nand U1509 (N_1509,N_1447,N_1494);
nor U1510 (N_1510,N_1482,N_1454);
and U1511 (N_1511,N_1446,N_1484);
and U1512 (N_1512,N_1468,N_1480);
nand U1513 (N_1513,N_1496,N_1492);
and U1514 (N_1514,N_1464,N_1493);
nand U1515 (N_1515,N_1471,N_1490);
nand U1516 (N_1516,N_1485,N_1465);
xnor U1517 (N_1517,N_1467,N_1457);
or U1518 (N_1518,N_1472,N_1459);
or U1519 (N_1519,N_1462,N_1498);
nand U1520 (N_1520,N_1455,N_1476);
nand U1521 (N_1521,N_1441,N_1444);
nand U1522 (N_1522,N_1497,N_1445);
and U1523 (N_1523,N_1470,N_1440);
nand U1524 (N_1524,N_1474,N_1456);
nand U1525 (N_1525,N_1478,N_1449);
nand U1526 (N_1526,N_1487,N_1448);
nand U1527 (N_1527,N_1443,N_1499);
and U1528 (N_1528,N_1452,N_1486);
nand U1529 (N_1529,N_1461,N_1469);
nor U1530 (N_1530,N_1480,N_1446);
nor U1531 (N_1531,N_1488,N_1484);
or U1532 (N_1532,N_1486,N_1440);
and U1533 (N_1533,N_1476,N_1463);
nor U1534 (N_1534,N_1440,N_1460);
or U1535 (N_1535,N_1470,N_1451);
and U1536 (N_1536,N_1445,N_1461);
nand U1537 (N_1537,N_1469,N_1447);
and U1538 (N_1538,N_1467,N_1452);
or U1539 (N_1539,N_1481,N_1471);
or U1540 (N_1540,N_1498,N_1464);
nand U1541 (N_1541,N_1487,N_1453);
or U1542 (N_1542,N_1442,N_1492);
and U1543 (N_1543,N_1455,N_1489);
nand U1544 (N_1544,N_1457,N_1459);
nor U1545 (N_1545,N_1460,N_1483);
and U1546 (N_1546,N_1487,N_1497);
and U1547 (N_1547,N_1476,N_1473);
and U1548 (N_1548,N_1453,N_1463);
nor U1549 (N_1549,N_1462,N_1441);
or U1550 (N_1550,N_1454,N_1445);
nand U1551 (N_1551,N_1471,N_1465);
nand U1552 (N_1552,N_1480,N_1494);
and U1553 (N_1553,N_1492,N_1448);
xnor U1554 (N_1554,N_1466,N_1443);
xor U1555 (N_1555,N_1488,N_1494);
nand U1556 (N_1556,N_1493,N_1451);
or U1557 (N_1557,N_1480,N_1461);
nand U1558 (N_1558,N_1465,N_1480);
or U1559 (N_1559,N_1471,N_1442);
nand U1560 (N_1560,N_1511,N_1517);
nand U1561 (N_1561,N_1527,N_1536);
and U1562 (N_1562,N_1507,N_1552);
nand U1563 (N_1563,N_1550,N_1542);
nor U1564 (N_1564,N_1540,N_1522);
nor U1565 (N_1565,N_1541,N_1516);
and U1566 (N_1566,N_1512,N_1543);
nor U1567 (N_1567,N_1520,N_1558);
nand U1568 (N_1568,N_1519,N_1523);
nor U1569 (N_1569,N_1508,N_1529);
nand U1570 (N_1570,N_1515,N_1525);
nand U1571 (N_1571,N_1533,N_1524);
and U1572 (N_1572,N_1551,N_1534);
nand U1573 (N_1573,N_1500,N_1518);
nand U1574 (N_1574,N_1547,N_1531);
nor U1575 (N_1575,N_1549,N_1528);
nand U1576 (N_1576,N_1546,N_1538);
or U1577 (N_1577,N_1501,N_1537);
nand U1578 (N_1578,N_1557,N_1532);
and U1579 (N_1579,N_1554,N_1556);
nor U1580 (N_1580,N_1509,N_1530);
nand U1581 (N_1581,N_1502,N_1514);
nor U1582 (N_1582,N_1521,N_1555);
or U1583 (N_1583,N_1559,N_1539);
nand U1584 (N_1584,N_1548,N_1510);
and U1585 (N_1585,N_1513,N_1505);
and U1586 (N_1586,N_1506,N_1526);
or U1587 (N_1587,N_1545,N_1504);
or U1588 (N_1588,N_1535,N_1544);
or U1589 (N_1589,N_1503,N_1553);
and U1590 (N_1590,N_1512,N_1556);
and U1591 (N_1591,N_1552,N_1508);
and U1592 (N_1592,N_1527,N_1513);
nand U1593 (N_1593,N_1525,N_1502);
and U1594 (N_1594,N_1507,N_1553);
nand U1595 (N_1595,N_1540,N_1546);
and U1596 (N_1596,N_1537,N_1553);
nand U1597 (N_1597,N_1500,N_1525);
or U1598 (N_1598,N_1525,N_1532);
and U1599 (N_1599,N_1512,N_1520);
nor U1600 (N_1600,N_1505,N_1508);
and U1601 (N_1601,N_1544,N_1552);
or U1602 (N_1602,N_1531,N_1520);
and U1603 (N_1603,N_1542,N_1523);
nand U1604 (N_1604,N_1524,N_1510);
and U1605 (N_1605,N_1539,N_1509);
nor U1606 (N_1606,N_1540,N_1536);
nor U1607 (N_1607,N_1525,N_1519);
xnor U1608 (N_1608,N_1517,N_1515);
nor U1609 (N_1609,N_1535,N_1511);
nor U1610 (N_1610,N_1502,N_1555);
and U1611 (N_1611,N_1557,N_1539);
nand U1612 (N_1612,N_1546,N_1522);
nand U1613 (N_1613,N_1520,N_1508);
nand U1614 (N_1614,N_1549,N_1548);
nand U1615 (N_1615,N_1509,N_1550);
nor U1616 (N_1616,N_1559,N_1516);
nor U1617 (N_1617,N_1548,N_1541);
nor U1618 (N_1618,N_1559,N_1558);
xnor U1619 (N_1619,N_1550,N_1548);
nand U1620 (N_1620,N_1607,N_1600);
nand U1621 (N_1621,N_1603,N_1598);
or U1622 (N_1622,N_1578,N_1599);
nor U1623 (N_1623,N_1573,N_1592);
nand U1624 (N_1624,N_1585,N_1589);
nor U1625 (N_1625,N_1560,N_1584);
or U1626 (N_1626,N_1619,N_1591);
nor U1627 (N_1627,N_1618,N_1569);
and U1628 (N_1628,N_1568,N_1608);
and U1629 (N_1629,N_1576,N_1613);
nor U1630 (N_1630,N_1561,N_1581);
nor U1631 (N_1631,N_1604,N_1580);
nand U1632 (N_1632,N_1577,N_1597);
nor U1633 (N_1633,N_1617,N_1609);
nand U1634 (N_1634,N_1571,N_1586);
or U1635 (N_1635,N_1593,N_1601);
nor U1636 (N_1636,N_1574,N_1583);
nand U1637 (N_1637,N_1611,N_1575);
and U1638 (N_1638,N_1579,N_1590);
or U1639 (N_1639,N_1587,N_1563);
nand U1640 (N_1640,N_1562,N_1570);
and U1641 (N_1641,N_1566,N_1596);
and U1642 (N_1642,N_1582,N_1612);
nor U1643 (N_1643,N_1567,N_1605);
and U1644 (N_1644,N_1564,N_1606);
nor U1645 (N_1645,N_1565,N_1616);
nand U1646 (N_1646,N_1614,N_1615);
nor U1647 (N_1647,N_1602,N_1594);
or U1648 (N_1648,N_1572,N_1610);
and U1649 (N_1649,N_1588,N_1595);
or U1650 (N_1650,N_1596,N_1565);
nand U1651 (N_1651,N_1580,N_1608);
or U1652 (N_1652,N_1598,N_1573);
nand U1653 (N_1653,N_1610,N_1598);
xor U1654 (N_1654,N_1600,N_1614);
nand U1655 (N_1655,N_1571,N_1572);
nor U1656 (N_1656,N_1576,N_1561);
or U1657 (N_1657,N_1571,N_1589);
or U1658 (N_1658,N_1607,N_1611);
xor U1659 (N_1659,N_1619,N_1563);
nand U1660 (N_1660,N_1576,N_1604);
or U1661 (N_1661,N_1563,N_1588);
nor U1662 (N_1662,N_1577,N_1565);
nand U1663 (N_1663,N_1567,N_1565);
or U1664 (N_1664,N_1579,N_1603);
and U1665 (N_1665,N_1567,N_1583);
or U1666 (N_1666,N_1560,N_1607);
and U1667 (N_1667,N_1573,N_1564);
or U1668 (N_1668,N_1601,N_1606);
and U1669 (N_1669,N_1585,N_1617);
nor U1670 (N_1670,N_1579,N_1604);
nor U1671 (N_1671,N_1574,N_1594);
nor U1672 (N_1672,N_1617,N_1593);
or U1673 (N_1673,N_1617,N_1586);
and U1674 (N_1674,N_1576,N_1617);
nor U1675 (N_1675,N_1612,N_1589);
xnor U1676 (N_1676,N_1604,N_1569);
nand U1677 (N_1677,N_1579,N_1586);
nand U1678 (N_1678,N_1580,N_1617);
nand U1679 (N_1679,N_1609,N_1597);
or U1680 (N_1680,N_1623,N_1639);
and U1681 (N_1681,N_1674,N_1649);
nand U1682 (N_1682,N_1651,N_1648);
or U1683 (N_1683,N_1634,N_1668);
nor U1684 (N_1684,N_1679,N_1663);
or U1685 (N_1685,N_1666,N_1660);
or U1686 (N_1686,N_1636,N_1667);
nor U1687 (N_1687,N_1676,N_1632);
and U1688 (N_1688,N_1630,N_1646);
or U1689 (N_1689,N_1661,N_1635);
nor U1690 (N_1690,N_1629,N_1625);
nor U1691 (N_1691,N_1653,N_1627);
nor U1692 (N_1692,N_1673,N_1624);
and U1693 (N_1693,N_1670,N_1672);
nor U1694 (N_1694,N_1647,N_1654);
nand U1695 (N_1695,N_1638,N_1658);
nor U1696 (N_1696,N_1652,N_1664);
nand U1697 (N_1697,N_1671,N_1656);
nand U1698 (N_1698,N_1677,N_1644);
and U1699 (N_1699,N_1622,N_1669);
nor U1700 (N_1700,N_1650,N_1640);
nand U1701 (N_1701,N_1628,N_1626);
nand U1702 (N_1702,N_1675,N_1643);
nand U1703 (N_1703,N_1665,N_1657);
and U1704 (N_1704,N_1678,N_1645);
or U1705 (N_1705,N_1631,N_1662);
nor U1706 (N_1706,N_1620,N_1633);
and U1707 (N_1707,N_1641,N_1637);
and U1708 (N_1708,N_1642,N_1659);
nor U1709 (N_1709,N_1655,N_1621);
nand U1710 (N_1710,N_1657,N_1633);
nor U1711 (N_1711,N_1657,N_1647);
and U1712 (N_1712,N_1663,N_1646);
or U1713 (N_1713,N_1627,N_1665);
nor U1714 (N_1714,N_1661,N_1633);
or U1715 (N_1715,N_1624,N_1644);
nor U1716 (N_1716,N_1622,N_1621);
nor U1717 (N_1717,N_1666,N_1641);
or U1718 (N_1718,N_1631,N_1675);
nor U1719 (N_1719,N_1636,N_1624);
and U1720 (N_1720,N_1666,N_1655);
and U1721 (N_1721,N_1641,N_1668);
nand U1722 (N_1722,N_1664,N_1627);
and U1723 (N_1723,N_1622,N_1662);
or U1724 (N_1724,N_1678,N_1657);
and U1725 (N_1725,N_1654,N_1637);
nand U1726 (N_1726,N_1637,N_1667);
nor U1727 (N_1727,N_1634,N_1666);
or U1728 (N_1728,N_1661,N_1662);
and U1729 (N_1729,N_1637,N_1622);
or U1730 (N_1730,N_1627,N_1644);
nor U1731 (N_1731,N_1659,N_1665);
nor U1732 (N_1732,N_1675,N_1670);
and U1733 (N_1733,N_1670,N_1657);
and U1734 (N_1734,N_1629,N_1678);
or U1735 (N_1735,N_1672,N_1657);
and U1736 (N_1736,N_1642,N_1676);
nor U1737 (N_1737,N_1679,N_1669);
nor U1738 (N_1738,N_1646,N_1666);
nor U1739 (N_1739,N_1642,N_1658);
nand U1740 (N_1740,N_1733,N_1729);
nor U1741 (N_1741,N_1685,N_1739);
and U1742 (N_1742,N_1702,N_1720);
or U1743 (N_1743,N_1736,N_1711);
nand U1744 (N_1744,N_1689,N_1701);
or U1745 (N_1745,N_1693,N_1691);
or U1746 (N_1746,N_1687,N_1683);
nor U1747 (N_1747,N_1680,N_1715);
nor U1748 (N_1748,N_1707,N_1704);
nand U1749 (N_1749,N_1703,N_1725);
or U1750 (N_1750,N_1686,N_1726);
and U1751 (N_1751,N_1708,N_1738);
or U1752 (N_1752,N_1716,N_1695);
nand U1753 (N_1753,N_1718,N_1727);
nand U1754 (N_1754,N_1697,N_1728);
and U1755 (N_1755,N_1696,N_1698);
nor U1756 (N_1756,N_1684,N_1717);
nand U1757 (N_1757,N_1719,N_1722);
or U1758 (N_1758,N_1723,N_1692);
and U1759 (N_1759,N_1731,N_1705);
nand U1760 (N_1760,N_1713,N_1681);
and U1761 (N_1761,N_1712,N_1732);
nand U1762 (N_1762,N_1724,N_1721);
or U1763 (N_1763,N_1730,N_1700);
or U1764 (N_1764,N_1734,N_1699);
xor U1765 (N_1765,N_1706,N_1714);
and U1766 (N_1766,N_1682,N_1737);
and U1767 (N_1767,N_1709,N_1690);
nor U1768 (N_1768,N_1694,N_1735);
nor U1769 (N_1769,N_1688,N_1710);
nor U1770 (N_1770,N_1686,N_1681);
nand U1771 (N_1771,N_1705,N_1681);
and U1772 (N_1772,N_1728,N_1713);
nor U1773 (N_1773,N_1687,N_1698);
nand U1774 (N_1774,N_1685,N_1703);
nor U1775 (N_1775,N_1687,N_1680);
and U1776 (N_1776,N_1736,N_1698);
nand U1777 (N_1777,N_1688,N_1714);
and U1778 (N_1778,N_1695,N_1723);
nor U1779 (N_1779,N_1701,N_1714);
and U1780 (N_1780,N_1693,N_1721);
and U1781 (N_1781,N_1724,N_1701);
and U1782 (N_1782,N_1732,N_1724);
and U1783 (N_1783,N_1719,N_1723);
nand U1784 (N_1784,N_1697,N_1684);
and U1785 (N_1785,N_1682,N_1694);
or U1786 (N_1786,N_1720,N_1736);
nand U1787 (N_1787,N_1697,N_1733);
nand U1788 (N_1788,N_1718,N_1698);
nor U1789 (N_1789,N_1684,N_1714);
and U1790 (N_1790,N_1721,N_1739);
or U1791 (N_1791,N_1702,N_1684);
and U1792 (N_1792,N_1719,N_1739);
nor U1793 (N_1793,N_1716,N_1709);
nand U1794 (N_1794,N_1733,N_1738);
nor U1795 (N_1795,N_1681,N_1696);
or U1796 (N_1796,N_1686,N_1689);
or U1797 (N_1797,N_1735,N_1722);
and U1798 (N_1798,N_1721,N_1685);
nor U1799 (N_1799,N_1710,N_1690);
nor U1800 (N_1800,N_1756,N_1743);
or U1801 (N_1801,N_1776,N_1767);
and U1802 (N_1802,N_1788,N_1786);
nor U1803 (N_1803,N_1772,N_1759);
or U1804 (N_1804,N_1751,N_1762);
or U1805 (N_1805,N_1766,N_1758);
nor U1806 (N_1806,N_1777,N_1785);
and U1807 (N_1807,N_1768,N_1773);
and U1808 (N_1808,N_1791,N_1761);
and U1809 (N_1809,N_1798,N_1754);
and U1810 (N_1810,N_1790,N_1775);
and U1811 (N_1811,N_1760,N_1765);
and U1812 (N_1812,N_1755,N_1770);
nor U1813 (N_1813,N_1769,N_1764);
and U1814 (N_1814,N_1742,N_1797);
or U1815 (N_1815,N_1781,N_1763);
nor U1816 (N_1816,N_1753,N_1741);
nand U1817 (N_1817,N_1748,N_1771);
nand U1818 (N_1818,N_1778,N_1793);
and U1819 (N_1819,N_1752,N_1787);
nand U1820 (N_1820,N_1779,N_1750);
and U1821 (N_1821,N_1792,N_1789);
or U1822 (N_1822,N_1774,N_1782);
and U1823 (N_1823,N_1795,N_1747);
nand U1824 (N_1824,N_1740,N_1799);
and U1825 (N_1825,N_1784,N_1744);
nor U1826 (N_1826,N_1796,N_1794);
nand U1827 (N_1827,N_1757,N_1783);
nor U1828 (N_1828,N_1749,N_1780);
nand U1829 (N_1829,N_1746,N_1745);
nand U1830 (N_1830,N_1796,N_1745);
and U1831 (N_1831,N_1776,N_1763);
nand U1832 (N_1832,N_1787,N_1756);
nand U1833 (N_1833,N_1747,N_1744);
nor U1834 (N_1834,N_1785,N_1765);
and U1835 (N_1835,N_1744,N_1771);
nor U1836 (N_1836,N_1794,N_1760);
nand U1837 (N_1837,N_1792,N_1750);
nand U1838 (N_1838,N_1797,N_1786);
nand U1839 (N_1839,N_1781,N_1785);
and U1840 (N_1840,N_1791,N_1798);
nand U1841 (N_1841,N_1742,N_1753);
nor U1842 (N_1842,N_1751,N_1743);
and U1843 (N_1843,N_1781,N_1754);
nand U1844 (N_1844,N_1793,N_1747);
nor U1845 (N_1845,N_1795,N_1753);
and U1846 (N_1846,N_1790,N_1779);
and U1847 (N_1847,N_1764,N_1780);
and U1848 (N_1848,N_1741,N_1758);
or U1849 (N_1849,N_1798,N_1771);
and U1850 (N_1850,N_1786,N_1750);
nand U1851 (N_1851,N_1759,N_1751);
nand U1852 (N_1852,N_1791,N_1779);
nand U1853 (N_1853,N_1797,N_1778);
nand U1854 (N_1854,N_1799,N_1754);
and U1855 (N_1855,N_1754,N_1760);
or U1856 (N_1856,N_1779,N_1740);
or U1857 (N_1857,N_1792,N_1766);
nand U1858 (N_1858,N_1768,N_1746);
nand U1859 (N_1859,N_1758,N_1788);
nor U1860 (N_1860,N_1859,N_1811);
and U1861 (N_1861,N_1843,N_1840);
nand U1862 (N_1862,N_1827,N_1848);
nand U1863 (N_1863,N_1836,N_1832);
and U1864 (N_1864,N_1807,N_1841);
nand U1865 (N_1865,N_1801,N_1802);
and U1866 (N_1866,N_1847,N_1817);
or U1867 (N_1867,N_1854,N_1808);
and U1868 (N_1868,N_1838,N_1835);
or U1869 (N_1869,N_1844,N_1824);
nand U1870 (N_1870,N_1856,N_1833);
or U1871 (N_1871,N_1809,N_1821);
nand U1872 (N_1872,N_1837,N_1834);
or U1873 (N_1873,N_1855,N_1829);
or U1874 (N_1874,N_1839,N_1815);
nor U1875 (N_1875,N_1830,N_1825);
and U1876 (N_1876,N_1819,N_1812);
nor U1877 (N_1877,N_1831,N_1853);
or U1878 (N_1878,N_1803,N_1828);
nor U1879 (N_1879,N_1804,N_1816);
nand U1880 (N_1880,N_1818,N_1813);
or U1881 (N_1881,N_1842,N_1851);
and U1882 (N_1882,N_1806,N_1850);
xor U1883 (N_1883,N_1805,N_1810);
and U1884 (N_1884,N_1857,N_1846);
nor U1885 (N_1885,N_1849,N_1814);
nand U1886 (N_1886,N_1820,N_1826);
nand U1887 (N_1887,N_1845,N_1858);
nor U1888 (N_1888,N_1823,N_1822);
xor U1889 (N_1889,N_1852,N_1800);
nor U1890 (N_1890,N_1806,N_1844);
nand U1891 (N_1891,N_1851,N_1843);
and U1892 (N_1892,N_1845,N_1842);
and U1893 (N_1893,N_1854,N_1848);
nor U1894 (N_1894,N_1810,N_1852);
or U1895 (N_1895,N_1833,N_1830);
and U1896 (N_1896,N_1841,N_1805);
nor U1897 (N_1897,N_1851,N_1821);
nor U1898 (N_1898,N_1826,N_1836);
nor U1899 (N_1899,N_1820,N_1827);
and U1900 (N_1900,N_1842,N_1810);
nand U1901 (N_1901,N_1801,N_1842);
nand U1902 (N_1902,N_1807,N_1854);
and U1903 (N_1903,N_1847,N_1815);
or U1904 (N_1904,N_1856,N_1851);
or U1905 (N_1905,N_1856,N_1827);
or U1906 (N_1906,N_1804,N_1827);
or U1907 (N_1907,N_1824,N_1842);
nor U1908 (N_1908,N_1807,N_1805);
and U1909 (N_1909,N_1824,N_1813);
or U1910 (N_1910,N_1848,N_1836);
xnor U1911 (N_1911,N_1842,N_1806);
nand U1912 (N_1912,N_1855,N_1854);
nand U1913 (N_1913,N_1830,N_1808);
or U1914 (N_1914,N_1821,N_1839);
nor U1915 (N_1915,N_1816,N_1820);
nand U1916 (N_1916,N_1834,N_1822);
or U1917 (N_1917,N_1828,N_1804);
xor U1918 (N_1918,N_1821,N_1802);
and U1919 (N_1919,N_1828,N_1833);
and U1920 (N_1920,N_1893,N_1891);
nor U1921 (N_1921,N_1865,N_1884);
or U1922 (N_1922,N_1898,N_1919);
and U1923 (N_1923,N_1904,N_1903);
nand U1924 (N_1924,N_1917,N_1886);
nor U1925 (N_1925,N_1914,N_1864);
and U1926 (N_1926,N_1870,N_1866);
nand U1927 (N_1927,N_1913,N_1890);
nand U1928 (N_1928,N_1908,N_1900);
or U1929 (N_1929,N_1869,N_1905);
nand U1930 (N_1930,N_1863,N_1899);
or U1931 (N_1931,N_1868,N_1877);
nand U1932 (N_1932,N_1876,N_1872);
nor U1933 (N_1933,N_1874,N_1867);
nor U1934 (N_1934,N_1897,N_1882);
nand U1935 (N_1935,N_1909,N_1883);
or U1936 (N_1936,N_1918,N_1894);
and U1937 (N_1937,N_1901,N_1880);
nand U1938 (N_1938,N_1889,N_1887);
nand U1939 (N_1939,N_1911,N_1906);
nor U1940 (N_1940,N_1878,N_1888);
or U1941 (N_1941,N_1875,N_1881);
nand U1942 (N_1942,N_1895,N_1892);
nor U1943 (N_1943,N_1916,N_1879);
nand U1944 (N_1944,N_1885,N_1862);
nor U1945 (N_1945,N_1871,N_1915);
nand U1946 (N_1946,N_1912,N_1896);
nor U1947 (N_1947,N_1902,N_1910);
and U1948 (N_1948,N_1861,N_1907);
and U1949 (N_1949,N_1860,N_1873);
or U1950 (N_1950,N_1885,N_1893);
nor U1951 (N_1951,N_1866,N_1861);
nor U1952 (N_1952,N_1910,N_1899);
or U1953 (N_1953,N_1899,N_1897);
nor U1954 (N_1954,N_1893,N_1882);
and U1955 (N_1955,N_1906,N_1896);
and U1956 (N_1956,N_1878,N_1915);
and U1957 (N_1957,N_1898,N_1891);
or U1958 (N_1958,N_1915,N_1904);
nand U1959 (N_1959,N_1869,N_1895);
nor U1960 (N_1960,N_1885,N_1875);
nor U1961 (N_1961,N_1866,N_1875);
nor U1962 (N_1962,N_1894,N_1905);
xor U1963 (N_1963,N_1875,N_1887);
nand U1964 (N_1964,N_1916,N_1887);
nor U1965 (N_1965,N_1910,N_1882);
or U1966 (N_1966,N_1862,N_1907);
xnor U1967 (N_1967,N_1864,N_1912);
or U1968 (N_1968,N_1890,N_1903);
and U1969 (N_1969,N_1863,N_1867);
nand U1970 (N_1970,N_1890,N_1885);
or U1971 (N_1971,N_1891,N_1897);
and U1972 (N_1972,N_1903,N_1889);
or U1973 (N_1973,N_1896,N_1918);
nor U1974 (N_1974,N_1863,N_1896);
or U1975 (N_1975,N_1861,N_1916);
and U1976 (N_1976,N_1891,N_1894);
nor U1977 (N_1977,N_1870,N_1874);
and U1978 (N_1978,N_1916,N_1876);
and U1979 (N_1979,N_1860,N_1919);
or U1980 (N_1980,N_1941,N_1951);
or U1981 (N_1981,N_1943,N_1940);
nor U1982 (N_1982,N_1965,N_1959);
nor U1983 (N_1983,N_1928,N_1974);
and U1984 (N_1984,N_1977,N_1953);
and U1985 (N_1985,N_1927,N_1939);
and U1986 (N_1986,N_1933,N_1957);
xnor U1987 (N_1987,N_1969,N_1948);
nand U1988 (N_1988,N_1963,N_1950);
and U1989 (N_1989,N_1960,N_1952);
nor U1990 (N_1990,N_1945,N_1935);
or U1991 (N_1991,N_1934,N_1973);
nor U1992 (N_1992,N_1938,N_1922);
nor U1993 (N_1993,N_1970,N_1942);
and U1994 (N_1994,N_1923,N_1937);
nand U1995 (N_1995,N_1921,N_1971);
nor U1996 (N_1996,N_1932,N_1956);
and U1997 (N_1997,N_1925,N_1949);
xnor U1998 (N_1998,N_1931,N_1967);
nor U1999 (N_1999,N_1968,N_1924);
or U2000 (N_2000,N_1930,N_1961);
and U2001 (N_2001,N_1946,N_1978);
xor U2002 (N_2002,N_1976,N_1975);
or U2003 (N_2003,N_1936,N_1964);
nand U2004 (N_2004,N_1979,N_1972);
and U2005 (N_2005,N_1920,N_1954);
or U2006 (N_2006,N_1955,N_1966);
nand U2007 (N_2007,N_1962,N_1929);
and U2008 (N_2008,N_1947,N_1926);
nor U2009 (N_2009,N_1958,N_1944);
nor U2010 (N_2010,N_1962,N_1947);
nor U2011 (N_2011,N_1925,N_1976);
nand U2012 (N_2012,N_1974,N_1949);
and U2013 (N_2013,N_1964,N_1958);
and U2014 (N_2014,N_1967,N_1963);
or U2015 (N_2015,N_1965,N_1949);
or U2016 (N_2016,N_1944,N_1963);
nor U2017 (N_2017,N_1966,N_1930);
and U2018 (N_2018,N_1966,N_1978);
and U2019 (N_2019,N_1978,N_1926);
nand U2020 (N_2020,N_1973,N_1945);
or U2021 (N_2021,N_1977,N_1965);
nor U2022 (N_2022,N_1932,N_1923);
and U2023 (N_2023,N_1921,N_1953);
or U2024 (N_2024,N_1922,N_1923);
nand U2025 (N_2025,N_1957,N_1935);
or U2026 (N_2026,N_1962,N_1936);
or U2027 (N_2027,N_1924,N_1941);
or U2028 (N_2028,N_1930,N_1942);
or U2029 (N_2029,N_1938,N_1970);
nor U2030 (N_2030,N_1944,N_1953);
or U2031 (N_2031,N_1965,N_1961);
nor U2032 (N_2032,N_1978,N_1920);
nand U2033 (N_2033,N_1959,N_1937);
and U2034 (N_2034,N_1922,N_1973);
nor U2035 (N_2035,N_1924,N_1979);
nor U2036 (N_2036,N_1925,N_1958);
or U2037 (N_2037,N_1925,N_1933);
nand U2038 (N_2038,N_1967,N_1955);
nand U2039 (N_2039,N_1968,N_1955);
xnor U2040 (N_2040,N_2028,N_2004);
nand U2041 (N_2041,N_2015,N_2012);
nand U2042 (N_2042,N_2003,N_1989);
and U2043 (N_2043,N_2036,N_1985);
or U2044 (N_2044,N_2039,N_2030);
nand U2045 (N_2045,N_1984,N_2019);
nor U2046 (N_2046,N_2025,N_2024);
and U2047 (N_2047,N_2007,N_1999);
or U2048 (N_2048,N_2000,N_2021);
nor U2049 (N_2049,N_1994,N_2033);
or U2050 (N_2050,N_1995,N_1996);
or U2051 (N_2051,N_2011,N_2013);
or U2052 (N_2052,N_1987,N_2022);
or U2053 (N_2053,N_2034,N_2035);
or U2054 (N_2054,N_2037,N_1982);
and U2055 (N_2055,N_2032,N_2031);
and U2056 (N_2056,N_2017,N_1988);
nand U2057 (N_2057,N_2023,N_2026);
nand U2058 (N_2058,N_2029,N_2008);
nand U2059 (N_2059,N_2038,N_1991);
or U2060 (N_2060,N_1990,N_2005);
or U2061 (N_2061,N_1986,N_1998);
or U2062 (N_2062,N_2016,N_1981);
xnor U2063 (N_2063,N_2002,N_2020);
nand U2064 (N_2064,N_1983,N_2001);
nor U2065 (N_2065,N_1980,N_2009);
nand U2066 (N_2066,N_2027,N_1992);
and U2067 (N_2067,N_1997,N_2018);
nand U2068 (N_2068,N_1993,N_2010);
nand U2069 (N_2069,N_2014,N_2006);
or U2070 (N_2070,N_1983,N_1980);
or U2071 (N_2071,N_2033,N_1999);
or U2072 (N_2072,N_2002,N_2023);
or U2073 (N_2073,N_2024,N_2020);
nand U2074 (N_2074,N_2016,N_2001);
or U2075 (N_2075,N_1991,N_2009);
nor U2076 (N_2076,N_2004,N_2021);
or U2077 (N_2077,N_2017,N_2002);
nand U2078 (N_2078,N_2011,N_2001);
nor U2079 (N_2079,N_1982,N_2026);
and U2080 (N_2080,N_1981,N_2007);
nand U2081 (N_2081,N_2032,N_2002);
and U2082 (N_2082,N_2019,N_2008);
or U2083 (N_2083,N_2033,N_2032);
nand U2084 (N_2084,N_2013,N_1981);
nand U2085 (N_2085,N_2005,N_2033);
nand U2086 (N_2086,N_2005,N_2039);
or U2087 (N_2087,N_2015,N_2001);
nor U2088 (N_2088,N_2031,N_2009);
nand U2089 (N_2089,N_2002,N_1986);
nand U2090 (N_2090,N_1988,N_2000);
and U2091 (N_2091,N_2000,N_2007);
and U2092 (N_2092,N_2030,N_2026);
and U2093 (N_2093,N_2036,N_2009);
and U2094 (N_2094,N_2023,N_1997);
and U2095 (N_2095,N_2017,N_2015);
nand U2096 (N_2096,N_2028,N_1999);
and U2097 (N_2097,N_1985,N_2002);
nand U2098 (N_2098,N_1992,N_2009);
or U2099 (N_2099,N_2015,N_1994);
or U2100 (N_2100,N_2083,N_2098);
xor U2101 (N_2101,N_2070,N_2063);
or U2102 (N_2102,N_2045,N_2066);
nand U2103 (N_2103,N_2075,N_2041);
and U2104 (N_2104,N_2061,N_2093);
nor U2105 (N_2105,N_2085,N_2052);
or U2106 (N_2106,N_2065,N_2071);
or U2107 (N_2107,N_2054,N_2096);
nand U2108 (N_2108,N_2055,N_2046);
nor U2109 (N_2109,N_2076,N_2072);
xor U2110 (N_2110,N_2049,N_2094);
and U2111 (N_2111,N_2086,N_2077);
nand U2112 (N_2112,N_2058,N_2068);
nor U2113 (N_2113,N_2089,N_2040);
or U2114 (N_2114,N_2050,N_2087);
and U2115 (N_2115,N_2091,N_2095);
nor U2116 (N_2116,N_2090,N_2059);
nand U2117 (N_2117,N_2080,N_2060);
nand U2118 (N_2118,N_2042,N_2069);
nand U2119 (N_2119,N_2078,N_2079);
nor U2120 (N_2120,N_2082,N_2067);
nand U2121 (N_2121,N_2053,N_2081);
or U2122 (N_2122,N_2088,N_2064);
or U2123 (N_2123,N_2043,N_2074);
nand U2124 (N_2124,N_2084,N_2057);
nor U2125 (N_2125,N_2097,N_2092);
and U2126 (N_2126,N_2051,N_2062);
or U2127 (N_2127,N_2048,N_2073);
or U2128 (N_2128,N_2056,N_2047);
nand U2129 (N_2129,N_2044,N_2099);
and U2130 (N_2130,N_2070,N_2044);
nand U2131 (N_2131,N_2068,N_2071);
or U2132 (N_2132,N_2075,N_2057);
and U2133 (N_2133,N_2061,N_2074);
nor U2134 (N_2134,N_2078,N_2049);
nand U2135 (N_2135,N_2042,N_2049);
nor U2136 (N_2136,N_2046,N_2090);
or U2137 (N_2137,N_2099,N_2045);
nand U2138 (N_2138,N_2047,N_2055);
or U2139 (N_2139,N_2060,N_2049);
nand U2140 (N_2140,N_2085,N_2086);
or U2141 (N_2141,N_2087,N_2040);
nand U2142 (N_2142,N_2096,N_2045);
nand U2143 (N_2143,N_2045,N_2061);
or U2144 (N_2144,N_2055,N_2067);
nand U2145 (N_2145,N_2055,N_2057);
nor U2146 (N_2146,N_2061,N_2095);
and U2147 (N_2147,N_2059,N_2069);
nand U2148 (N_2148,N_2050,N_2067);
and U2149 (N_2149,N_2056,N_2063);
or U2150 (N_2150,N_2064,N_2068);
or U2151 (N_2151,N_2088,N_2092);
and U2152 (N_2152,N_2091,N_2071);
and U2153 (N_2153,N_2052,N_2072);
and U2154 (N_2154,N_2059,N_2045);
and U2155 (N_2155,N_2077,N_2044);
or U2156 (N_2156,N_2083,N_2093);
nand U2157 (N_2157,N_2063,N_2078);
and U2158 (N_2158,N_2098,N_2061);
or U2159 (N_2159,N_2094,N_2046);
and U2160 (N_2160,N_2130,N_2152);
nor U2161 (N_2161,N_2121,N_2103);
or U2162 (N_2162,N_2134,N_2140);
and U2163 (N_2163,N_2149,N_2126);
or U2164 (N_2164,N_2110,N_2154);
nand U2165 (N_2165,N_2104,N_2114);
and U2166 (N_2166,N_2138,N_2111);
nand U2167 (N_2167,N_2113,N_2137);
and U2168 (N_2168,N_2142,N_2141);
nor U2169 (N_2169,N_2136,N_2151);
and U2170 (N_2170,N_2112,N_2120);
nand U2171 (N_2171,N_2123,N_2117);
nand U2172 (N_2172,N_2100,N_2105);
and U2173 (N_2173,N_2124,N_2139);
and U2174 (N_2174,N_2122,N_2158);
and U2175 (N_2175,N_2155,N_2146);
or U2176 (N_2176,N_2156,N_2127);
and U2177 (N_2177,N_2129,N_2109);
and U2178 (N_2178,N_2115,N_2143);
nand U2179 (N_2179,N_2132,N_2102);
nand U2180 (N_2180,N_2116,N_2107);
nand U2181 (N_2181,N_2133,N_2144);
or U2182 (N_2182,N_2128,N_2125);
or U2183 (N_2183,N_2148,N_2101);
and U2184 (N_2184,N_2131,N_2118);
nor U2185 (N_2185,N_2108,N_2150);
nand U2186 (N_2186,N_2106,N_2157);
or U2187 (N_2187,N_2135,N_2153);
or U2188 (N_2188,N_2119,N_2147);
and U2189 (N_2189,N_2145,N_2159);
and U2190 (N_2190,N_2101,N_2149);
nand U2191 (N_2191,N_2121,N_2128);
nor U2192 (N_2192,N_2142,N_2115);
or U2193 (N_2193,N_2155,N_2101);
or U2194 (N_2194,N_2116,N_2154);
nor U2195 (N_2195,N_2139,N_2108);
or U2196 (N_2196,N_2154,N_2114);
nand U2197 (N_2197,N_2149,N_2128);
nor U2198 (N_2198,N_2156,N_2123);
or U2199 (N_2199,N_2151,N_2152);
nand U2200 (N_2200,N_2139,N_2121);
nor U2201 (N_2201,N_2122,N_2127);
or U2202 (N_2202,N_2145,N_2107);
or U2203 (N_2203,N_2134,N_2104);
nand U2204 (N_2204,N_2111,N_2148);
and U2205 (N_2205,N_2130,N_2116);
xnor U2206 (N_2206,N_2121,N_2129);
and U2207 (N_2207,N_2127,N_2140);
or U2208 (N_2208,N_2126,N_2145);
and U2209 (N_2209,N_2156,N_2131);
nor U2210 (N_2210,N_2136,N_2150);
and U2211 (N_2211,N_2154,N_2155);
xnor U2212 (N_2212,N_2156,N_2132);
or U2213 (N_2213,N_2130,N_2132);
nand U2214 (N_2214,N_2102,N_2124);
and U2215 (N_2215,N_2127,N_2141);
nor U2216 (N_2216,N_2129,N_2150);
and U2217 (N_2217,N_2118,N_2139);
nand U2218 (N_2218,N_2145,N_2112);
nor U2219 (N_2219,N_2111,N_2114);
nor U2220 (N_2220,N_2199,N_2195);
nand U2221 (N_2221,N_2200,N_2217);
nor U2222 (N_2222,N_2171,N_2178);
and U2223 (N_2223,N_2219,N_2190);
or U2224 (N_2224,N_2167,N_2164);
or U2225 (N_2225,N_2175,N_2210);
and U2226 (N_2226,N_2204,N_2194);
or U2227 (N_2227,N_2163,N_2177);
nand U2228 (N_2228,N_2172,N_2188);
or U2229 (N_2229,N_2180,N_2198);
nor U2230 (N_2230,N_2173,N_2170);
nor U2231 (N_2231,N_2213,N_2166);
or U2232 (N_2232,N_2207,N_2176);
nor U2233 (N_2233,N_2181,N_2183);
and U2234 (N_2234,N_2160,N_2168);
or U2235 (N_2235,N_2218,N_2209);
nand U2236 (N_2236,N_2186,N_2205);
nor U2237 (N_2237,N_2206,N_2196);
or U2238 (N_2238,N_2165,N_2215);
nand U2239 (N_2239,N_2202,N_2197);
and U2240 (N_2240,N_2216,N_2191);
and U2241 (N_2241,N_2193,N_2184);
and U2242 (N_2242,N_2187,N_2174);
nor U2243 (N_2243,N_2214,N_2189);
nor U2244 (N_2244,N_2208,N_2169);
or U2245 (N_2245,N_2203,N_2162);
nor U2246 (N_2246,N_2182,N_2161);
and U2247 (N_2247,N_2201,N_2179);
nand U2248 (N_2248,N_2211,N_2192);
nand U2249 (N_2249,N_2212,N_2185);
nor U2250 (N_2250,N_2197,N_2162);
or U2251 (N_2251,N_2207,N_2191);
nand U2252 (N_2252,N_2179,N_2168);
or U2253 (N_2253,N_2202,N_2170);
or U2254 (N_2254,N_2176,N_2177);
nor U2255 (N_2255,N_2205,N_2217);
nand U2256 (N_2256,N_2211,N_2218);
and U2257 (N_2257,N_2204,N_2167);
or U2258 (N_2258,N_2206,N_2171);
nand U2259 (N_2259,N_2202,N_2206);
nor U2260 (N_2260,N_2197,N_2163);
and U2261 (N_2261,N_2200,N_2203);
or U2262 (N_2262,N_2212,N_2201);
or U2263 (N_2263,N_2200,N_2189);
and U2264 (N_2264,N_2171,N_2176);
nor U2265 (N_2265,N_2185,N_2180);
or U2266 (N_2266,N_2187,N_2164);
nand U2267 (N_2267,N_2209,N_2207);
nand U2268 (N_2268,N_2207,N_2170);
nand U2269 (N_2269,N_2167,N_2172);
or U2270 (N_2270,N_2170,N_2218);
and U2271 (N_2271,N_2169,N_2196);
nor U2272 (N_2272,N_2161,N_2174);
or U2273 (N_2273,N_2162,N_2172);
nand U2274 (N_2274,N_2164,N_2163);
and U2275 (N_2275,N_2164,N_2199);
nand U2276 (N_2276,N_2166,N_2172);
nand U2277 (N_2277,N_2183,N_2172);
nand U2278 (N_2278,N_2173,N_2167);
nor U2279 (N_2279,N_2201,N_2197);
or U2280 (N_2280,N_2232,N_2238);
nor U2281 (N_2281,N_2220,N_2241);
nor U2282 (N_2282,N_2275,N_2265);
nand U2283 (N_2283,N_2221,N_2237);
nand U2284 (N_2284,N_2260,N_2240);
nand U2285 (N_2285,N_2231,N_2252);
nor U2286 (N_2286,N_2268,N_2222);
or U2287 (N_2287,N_2274,N_2242);
and U2288 (N_2288,N_2228,N_2226);
or U2289 (N_2289,N_2277,N_2225);
nand U2290 (N_2290,N_2273,N_2269);
and U2291 (N_2291,N_2227,N_2239);
nor U2292 (N_2292,N_2246,N_2247);
and U2293 (N_2293,N_2278,N_2243);
or U2294 (N_2294,N_2270,N_2230);
nor U2295 (N_2295,N_2276,N_2250);
nand U2296 (N_2296,N_2248,N_2236);
nand U2297 (N_2297,N_2251,N_2235);
nor U2298 (N_2298,N_2272,N_2259);
or U2299 (N_2299,N_2234,N_2253);
and U2300 (N_2300,N_2258,N_2244);
or U2301 (N_2301,N_2257,N_2255);
xnor U2302 (N_2302,N_2254,N_2264);
nand U2303 (N_2303,N_2249,N_2229);
and U2304 (N_2304,N_2266,N_2262);
nand U2305 (N_2305,N_2267,N_2223);
nand U2306 (N_2306,N_2279,N_2245);
nand U2307 (N_2307,N_2233,N_2256);
nand U2308 (N_2308,N_2261,N_2224);
nor U2309 (N_2309,N_2271,N_2263);
or U2310 (N_2310,N_2241,N_2244);
and U2311 (N_2311,N_2260,N_2252);
nand U2312 (N_2312,N_2237,N_2223);
nand U2313 (N_2313,N_2254,N_2231);
nand U2314 (N_2314,N_2269,N_2257);
nor U2315 (N_2315,N_2272,N_2270);
nand U2316 (N_2316,N_2264,N_2277);
nor U2317 (N_2317,N_2225,N_2242);
nor U2318 (N_2318,N_2228,N_2224);
or U2319 (N_2319,N_2263,N_2257);
and U2320 (N_2320,N_2235,N_2272);
and U2321 (N_2321,N_2232,N_2254);
nor U2322 (N_2322,N_2234,N_2269);
and U2323 (N_2323,N_2256,N_2242);
nand U2324 (N_2324,N_2227,N_2271);
and U2325 (N_2325,N_2264,N_2228);
nand U2326 (N_2326,N_2235,N_2259);
nand U2327 (N_2327,N_2244,N_2248);
nor U2328 (N_2328,N_2274,N_2260);
nand U2329 (N_2329,N_2258,N_2261);
nor U2330 (N_2330,N_2266,N_2264);
or U2331 (N_2331,N_2227,N_2240);
and U2332 (N_2332,N_2229,N_2257);
or U2333 (N_2333,N_2269,N_2264);
nand U2334 (N_2334,N_2228,N_2274);
nand U2335 (N_2335,N_2222,N_2234);
or U2336 (N_2336,N_2259,N_2253);
or U2337 (N_2337,N_2256,N_2244);
and U2338 (N_2338,N_2248,N_2243);
nor U2339 (N_2339,N_2234,N_2244);
or U2340 (N_2340,N_2290,N_2336);
or U2341 (N_2341,N_2331,N_2321);
or U2342 (N_2342,N_2329,N_2281);
or U2343 (N_2343,N_2289,N_2325);
nand U2344 (N_2344,N_2307,N_2303);
and U2345 (N_2345,N_2296,N_2334);
and U2346 (N_2346,N_2291,N_2309);
xor U2347 (N_2347,N_2311,N_2292);
or U2348 (N_2348,N_2322,N_2335);
nor U2349 (N_2349,N_2282,N_2315);
and U2350 (N_2350,N_2337,N_2320);
nor U2351 (N_2351,N_2304,N_2283);
nand U2352 (N_2352,N_2287,N_2288);
nor U2353 (N_2353,N_2318,N_2293);
nand U2354 (N_2354,N_2302,N_2297);
or U2355 (N_2355,N_2280,N_2295);
and U2356 (N_2356,N_2314,N_2323);
nand U2357 (N_2357,N_2326,N_2310);
and U2358 (N_2358,N_2313,N_2338);
nand U2359 (N_2359,N_2330,N_2300);
nor U2360 (N_2360,N_2298,N_2306);
nand U2361 (N_2361,N_2317,N_2324);
nand U2362 (N_2362,N_2284,N_2299);
nand U2363 (N_2363,N_2308,N_2332);
xnor U2364 (N_2364,N_2333,N_2327);
and U2365 (N_2365,N_2294,N_2301);
or U2366 (N_2366,N_2339,N_2319);
nor U2367 (N_2367,N_2285,N_2286);
nand U2368 (N_2368,N_2312,N_2316);
and U2369 (N_2369,N_2328,N_2305);
nand U2370 (N_2370,N_2284,N_2338);
nand U2371 (N_2371,N_2314,N_2289);
nor U2372 (N_2372,N_2292,N_2325);
nor U2373 (N_2373,N_2304,N_2335);
nand U2374 (N_2374,N_2321,N_2305);
nor U2375 (N_2375,N_2287,N_2292);
nand U2376 (N_2376,N_2311,N_2326);
and U2377 (N_2377,N_2287,N_2286);
nand U2378 (N_2378,N_2295,N_2328);
and U2379 (N_2379,N_2329,N_2286);
nand U2380 (N_2380,N_2317,N_2318);
or U2381 (N_2381,N_2338,N_2329);
nand U2382 (N_2382,N_2303,N_2321);
nor U2383 (N_2383,N_2280,N_2310);
nor U2384 (N_2384,N_2311,N_2300);
nand U2385 (N_2385,N_2282,N_2332);
nor U2386 (N_2386,N_2303,N_2330);
and U2387 (N_2387,N_2290,N_2332);
nor U2388 (N_2388,N_2312,N_2298);
and U2389 (N_2389,N_2295,N_2290);
nand U2390 (N_2390,N_2297,N_2325);
or U2391 (N_2391,N_2328,N_2333);
or U2392 (N_2392,N_2338,N_2280);
and U2393 (N_2393,N_2326,N_2283);
nor U2394 (N_2394,N_2319,N_2286);
or U2395 (N_2395,N_2314,N_2290);
nor U2396 (N_2396,N_2287,N_2336);
and U2397 (N_2397,N_2331,N_2337);
nand U2398 (N_2398,N_2326,N_2294);
nand U2399 (N_2399,N_2288,N_2310);
and U2400 (N_2400,N_2374,N_2384);
and U2401 (N_2401,N_2394,N_2354);
and U2402 (N_2402,N_2376,N_2389);
nand U2403 (N_2403,N_2398,N_2379);
nand U2404 (N_2404,N_2358,N_2348);
nor U2405 (N_2405,N_2365,N_2390);
or U2406 (N_2406,N_2350,N_2349);
nor U2407 (N_2407,N_2363,N_2399);
and U2408 (N_2408,N_2367,N_2345);
nor U2409 (N_2409,N_2382,N_2385);
and U2410 (N_2410,N_2364,N_2359);
nor U2411 (N_2411,N_2395,N_2396);
or U2412 (N_2412,N_2388,N_2386);
and U2413 (N_2413,N_2352,N_2380);
nand U2414 (N_2414,N_2387,N_2375);
nand U2415 (N_2415,N_2351,N_2397);
or U2416 (N_2416,N_2360,N_2346);
nand U2417 (N_2417,N_2362,N_2391);
nand U2418 (N_2418,N_2371,N_2383);
nor U2419 (N_2419,N_2341,N_2347);
and U2420 (N_2420,N_2373,N_2355);
nand U2421 (N_2421,N_2343,N_2353);
and U2422 (N_2422,N_2361,N_2356);
xor U2423 (N_2423,N_2377,N_2368);
and U2424 (N_2424,N_2378,N_2366);
nand U2425 (N_2425,N_2344,N_2370);
and U2426 (N_2426,N_2392,N_2340);
nor U2427 (N_2427,N_2357,N_2381);
and U2428 (N_2428,N_2369,N_2372);
nor U2429 (N_2429,N_2342,N_2393);
and U2430 (N_2430,N_2368,N_2367);
and U2431 (N_2431,N_2393,N_2383);
nor U2432 (N_2432,N_2350,N_2368);
or U2433 (N_2433,N_2344,N_2392);
and U2434 (N_2434,N_2376,N_2384);
xor U2435 (N_2435,N_2377,N_2360);
or U2436 (N_2436,N_2362,N_2346);
nand U2437 (N_2437,N_2396,N_2361);
nand U2438 (N_2438,N_2390,N_2346);
nor U2439 (N_2439,N_2373,N_2362);
and U2440 (N_2440,N_2379,N_2343);
or U2441 (N_2441,N_2373,N_2375);
and U2442 (N_2442,N_2392,N_2385);
nand U2443 (N_2443,N_2356,N_2378);
and U2444 (N_2444,N_2347,N_2362);
or U2445 (N_2445,N_2346,N_2388);
xor U2446 (N_2446,N_2366,N_2368);
and U2447 (N_2447,N_2364,N_2390);
or U2448 (N_2448,N_2396,N_2369);
nor U2449 (N_2449,N_2379,N_2354);
and U2450 (N_2450,N_2353,N_2395);
and U2451 (N_2451,N_2350,N_2375);
and U2452 (N_2452,N_2362,N_2376);
nand U2453 (N_2453,N_2342,N_2379);
nand U2454 (N_2454,N_2382,N_2392);
nor U2455 (N_2455,N_2369,N_2389);
or U2456 (N_2456,N_2377,N_2341);
or U2457 (N_2457,N_2368,N_2357);
or U2458 (N_2458,N_2362,N_2381);
and U2459 (N_2459,N_2380,N_2360);
nand U2460 (N_2460,N_2442,N_2449);
nand U2461 (N_2461,N_2445,N_2427);
nand U2462 (N_2462,N_2459,N_2436);
and U2463 (N_2463,N_2454,N_2455);
and U2464 (N_2464,N_2440,N_2431);
or U2465 (N_2465,N_2418,N_2450);
or U2466 (N_2466,N_2441,N_2435);
nor U2467 (N_2467,N_2430,N_2428);
nor U2468 (N_2468,N_2410,N_2412);
and U2469 (N_2469,N_2452,N_2420);
nor U2470 (N_2470,N_2408,N_2407);
and U2471 (N_2471,N_2409,N_2451);
nand U2472 (N_2472,N_2426,N_2425);
nand U2473 (N_2473,N_2453,N_2456);
nand U2474 (N_2474,N_2415,N_2447);
nand U2475 (N_2475,N_2423,N_2419);
and U2476 (N_2476,N_2458,N_2443);
nor U2477 (N_2477,N_2448,N_2446);
nand U2478 (N_2478,N_2457,N_2405);
nand U2479 (N_2479,N_2417,N_2414);
nand U2480 (N_2480,N_2401,N_2444);
and U2481 (N_2481,N_2439,N_2438);
and U2482 (N_2482,N_2424,N_2402);
and U2483 (N_2483,N_2437,N_2422);
and U2484 (N_2484,N_2429,N_2403);
nand U2485 (N_2485,N_2411,N_2434);
or U2486 (N_2486,N_2433,N_2400);
nand U2487 (N_2487,N_2404,N_2416);
nor U2488 (N_2488,N_2432,N_2421);
and U2489 (N_2489,N_2406,N_2413);
and U2490 (N_2490,N_2440,N_2414);
or U2491 (N_2491,N_2441,N_2444);
and U2492 (N_2492,N_2447,N_2423);
or U2493 (N_2493,N_2412,N_2430);
or U2494 (N_2494,N_2435,N_2405);
or U2495 (N_2495,N_2407,N_2450);
or U2496 (N_2496,N_2423,N_2451);
nor U2497 (N_2497,N_2421,N_2448);
and U2498 (N_2498,N_2439,N_2448);
or U2499 (N_2499,N_2458,N_2412);
nand U2500 (N_2500,N_2412,N_2422);
or U2501 (N_2501,N_2440,N_2438);
and U2502 (N_2502,N_2414,N_2448);
or U2503 (N_2503,N_2431,N_2407);
nand U2504 (N_2504,N_2457,N_2450);
or U2505 (N_2505,N_2429,N_2401);
nor U2506 (N_2506,N_2435,N_2428);
and U2507 (N_2507,N_2416,N_2417);
and U2508 (N_2508,N_2405,N_2421);
xnor U2509 (N_2509,N_2429,N_2409);
nand U2510 (N_2510,N_2426,N_2410);
and U2511 (N_2511,N_2458,N_2414);
nor U2512 (N_2512,N_2424,N_2457);
nand U2513 (N_2513,N_2438,N_2455);
or U2514 (N_2514,N_2447,N_2451);
or U2515 (N_2515,N_2443,N_2403);
nand U2516 (N_2516,N_2450,N_2455);
nor U2517 (N_2517,N_2438,N_2408);
or U2518 (N_2518,N_2428,N_2420);
or U2519 (N_2519,N_2459,N_2423);
and U2520 (N_2520,N_2504,N_2503);
and U2521 (N_2521,N_2515,N_2494);
nor U2522 (N_2522,N_2478,N_2518);
nor U2523 (N_2523,N_2500,N_2517);
nor U2524 (N_2524,N_2476,N_2491);
nand U2525 (N_2525,N_2486,N_2475);
or U2526 (N_2526,N_2513,N_2510);
and U2527 (N_2527,N_2482,N_2472);
or U2528 (N_2528,N_2489,N_2481);
and U2529 (N_2529,N_2509,N_2483);
and U2530 (N_2530,N_2480,N_2511);
nor U2531 (N_2531,N_2463,N_2465);
or U2532 (N_2532,N_2496,N_2501);
and U2533 (N_2533,N_2516,N_2493);
nor U2534 (N_2534,N_2502,N_2477);
nand U2535 (N_2535,N_2497,N_2473);
nor U2536 (N_2536,N_2470,N_2514);
nor U2537 (N_2537,N_2461,N_2488);
or U2538 (N_2538,N_2462,N_2519);
nand U2539 (N_2539,N_2460,N_2505);
and U2540 (N_2540,N_2474,N_2507);
or U2541 (N_2541,N_2479,N_2498);
or U2542 (N_2542,N_2468,N_2487);
nand U2543 (N_2543,N_2495,N_2484);
and U2544 (N_2544,N_2467,N_2492);
nand U2545 (N_2545,N_2499,N_2508);
or U2546 (N_2546,N_2490,N_2466);
nor U2547 (N_2547,N_2471,N_2506);
nor U2548 (N_2548,N_2469,N_2464);
and U2549 (N_2549,N_2512,N_2485);
nor U2550 (N_2550,N_2480,N_2501);
and U2551 (N_2551,N_2514,N_2493);
nand U2552 (N_2552,N_2481,N_2480);
nand U2553 (N_2553,N_2501,N_2461);
and U2554 (N_2554,N_2466,N_2472);
and U2555 (N_2555,N_2463,N_2484);
or U2556 (N_2556,N_2512,N_2489);
and U2557 (N_2557,N_2464,N_2494);
nand U2558 (N_2558,N_2464,N_2493);
or U2559 (N_2559,N_2504,N_2490);
nand U2560 (N_2560,N_2508,N_2461);
and U2561 (N_2561,N_2509,N_2479);
and U2562 (N_2562,N_2515,N_2462);
nand U2563 (N_2563,N_2491,N_2518);
nor U2564 (N_2564,N_2481,N_2492);
and U2565 (N_2565,N_2496,N_2485);
nand U2566 (N_2566,N_2514,N_2461);
nand U2567 (N_2567,N_2515,N_2490);
nand U2568 (N_2568,N_2516,N_2515);
nand U2569 (N_2569,N_2482,N_2497);
nand U2570 (N_2570,N_2472,N_2504);
nand U2571 (N_2571,N_2474,N_2489);
or U2572 (N_2572,N_2501,N_2513);
nand U2573 (N_2573,N_2515,N_2472);
and U2574 (N_2574,N_2510,N_2499);
nor U2575 (N_2575,N_2515,N_2467);
and U2576 (N_2576,N_2498,N_2492);
and U2577 (N_2577,N_2511,N_2517);
nand U2578 (N_2578,N_2514,N_2467);
or U2579 (N_2579,N_2510,N_2478);
nand U2580 (N_2580,N_2537,N_2535);
nor U2581 (N_2581,N_2571,N_2543);
nand U2582 (N_2582,N_2536,N_2523);
nor U2583 (N_2583,N_2549,N_2550);
or U2584 (N_2584,N_2579,N_2522);
and U2585 (N_2585,N_2578,N_2561);
nand U2586 (N_2586,N_2533,N_2567);
and U2587 (N_2587,N_2541,N_2524);
or U2588 (N_2588,N_2570,N_2564);
and U2589 (N_2589,N_2553,N_2525);
nand U2590 (N_2590,N_2573,N_2526);
xor U2591 (N_2591,N_2558,N_2540);
nor U2592 (N_2592,N_2521,N_2560);
nand U2593 (N_2593,N_2574,N_2539);
or U2594 (N_2594,N_2531,N_2542);
and U2595 (N_2595,N_2545,N_2520);
nor U2596 (N_2596,N_2548,N_2547);
nor U2597 (N_2597,N_2527,N_2532);
nand U2598 (N_2598,N_2563,N_2555);
and U2599 (N_2599,N_2577,N_2552);
and U2600 (N_2600,N_2575,N_2538);
or U2601 (N_2601,N_2528,N_2562);
nor U2602 (N_2602,N_2569,N_2529);
nand U2603 (N_2603,N_2530,N_2566);
nor U2604 (N_2604,N_2546,N_2534);
and U2605 (N_2605,N_2551,N_2572);
or U2606 (N_2606,N_2554,N_2576);
or U2607 (N_2607,N_2544,N_2568);
and U2608 (N_2608,N_2557,N_2556);
or U2609 (N_2609,N_2559,N_2565);
or U2610 (N_2610,N_2571,N_2534);
or U2611 (N_2611,N_2578,N_2575);
xor U2612 (N_2612,N_2570,N_2549);
and U2613 (N_2613,N_2560,N_2557);
nand U2614 (N_2614,N_2524,N_2544);
or U2615 (N_2615,N_2566,N_2550);
and U2616 (N_2616,N_2579,N_2530);
or U2617 (N_2617,N_2556,N_2553);
and U2618 (N_2618,N_2529,N_2531);
and U2619 (N_2619,N_2549,N_2565);
nor U2620 (N_2620,N_2549,N_2532);
or U2621 (N_2621,N_2546,N_2571);
nor U2622 (N_2622,N_2542,N_2520);
nand U2623 (N_2623,N_2570,N_2535);
nor U2624 (N_2624,N_2533,N_2543);
xor U2625 (N_2625,N_2556,N_2572);
nand U2626 (N_2626,N_2532,N_2566);
nand U2627 (N_2627,N_2551,N_2520);
nand U2628 (N_2628,N_2532,N_2571);
nand U2629 (N_2629,N_2522,N_2533);
nand U2630 (N_2630,N_2559,N_2521);
and U2631 (N_2631,N_2567,N_2542);
xnor U2632 (N_2632,N_2577,N_2545);
and U2633 (N_2633,N_2523,N_2545);
or U2634 (N_2634,N_2573,N_2570);
nor U2635 (N_2635,N_2567,N_2520);
and U2636 (N_2636,N_2533,N_2559);
and U2637 (N_2637,N_2579,N_2564);
nand U2638 (N_2638,N_2553,N_2560);
nand U2639 (N_2639,N_2541,N_2534);
and U2640 (N_2640,N_2591,N_2583);
and U2641 (N_2641,N_2586,N_2600);
or U2642 (N_2642,N_2623,N_2597);
and U2643 (N_2643,N_2622,N_2590);
and U2644 (N_2644,N_2629,N_2606);
nand U2645 (N_2645,N_2621,N_2588);
nor U2646 (N_2646,N_2627,N_2637);
nand U2647 (N_2647,N_2595,N_2584);
nor U2648 (N_2648,N_2592,N_2620);
or U2649 (N_2649,N_2609,N_2602);
or U2650 (N_2650,N_2596,N_2581);
nand U2651 (N_2651,N_2612,N_2585);
nor U2652 (N_2652,N_2626,N_2605);
and U2653 (N_2653,N_2619,N_2625);
nor U2654 (N_2654,N_2601,N_2598);
nor U2655 (N_2655,N_2589,N_2593);
and U2656 (N_2656,N_2613,N_2638);
nor U2657 (N_2657,N_2610,N_2580);
and U2658 (N_2658,N_2587,N_2632);
nor U2659 (N_2659,N_2628,N_2604);
nor U2660 (N_2660,N_2615,N_2630);
and U2661 (N_2661,N_2599,N_2624);
or U2662 (N_2662,N_2633,N_2635);
nand U2663 (N_2663,N_2616,N_2618);
or U2664 (N_2664,N_2614,N_2639);
and U2665 (N_2665,N_2636,N_2617);
or U2666 (N_2666,N_2594,N_2582);
and U2667 (N_2667,N_2603,N_2607);
and U2668 (N_2668,N_2631,N_2611);
nor U2669 (N_2669,N_2608,N_2634);
nand U2670 (N_2670,N_2619,N_2637);
nand U2671 (N_2671,N_2583,N_2621);
nand U2672 (N_2672,N_2604,N_2619);
nor U2673 (N_2673,N_2617,N_2611);
and U2674 (N_2674,N_2623,N_2581);
and U2675 (N_2675,N_2592,N_2608);
or U2676 (N_2676,N_2582,N_2587);
nand U2677 (N_2677,N_2608,N_2593);
nand U2678 (N_2678,N_2623,N_2621);
nor U2679 (N_2679,N_2630,N_2582);
and U2680 (N_2680,N_2629,N_2620);
xor U2681 (N_2681,N_2590,N_2632);
nor U2682 (N_2682,N_2634,N_2583);
nor U2683 (N_2683,N_2615,N_2598);
or U2684 (N_2684,N_2626,N_2623);
and U2685 (N_2685,N_2636,N_2614);
nand U2686 (N_2686,N_2611,N_2636);
nand U2687 (N_2687,N_2628,N_2596);
nor U2688 (N_2688,N_2589,N_2631);
and U2689 (N_2689,N_2602,N_2588);
nor U2690 (N_2690,N_2596,N_2607);
or U2691 (N_2691,N_2608,N_2580);
nand U2692 (N_2692,N_2589,N_2582);
nor U2693 (N_2693,N_2616,N_2592);
and U2694 (N_2694,N_2637,N_2613);
or U2695 (N_2695,N_2610,N_2622);
nor U2696 (N_2696,N_2604,N_2584);
nand U2697 (N_2697,N_2628,N_2626);
and U2698 (N_2698,N_2630,N_2597);
nor U2699 (N_2699,N_2631,N_2608);
nand U2700 (N_2700,N_2673,N_2696);
nand U2701 (N_2701,N_2694,N_2663);
nand U2702 (N_2702,N_2693,N_2650);
and U2703 (N_2703,N_2689,N_2671);
and U2704 (N_2704,N_2666,N_2658);
nor U2705 (N_2705,N_2695,N_2661);
xnor U2706 (N_2706,N_2675,N_2667);
nand U2707 (N_2707,N_2690,N_2657);
or U2708 (N_2708,N_2686,N_2679);
xor U2709 (N_2709,N_2677,N_2648);
or U2710 (N_2710,N_2681,N_2698);
and U2711 (N_2711,N_2670,N_2662);
nor U2712 (N_2712,N_2678,N_2688);
or U2713 (N_2713,N_2691,N_2655);
nor U2714 (N_2714,N_2644,N_2664);
or U2715 (N_2715,N_2676,N_2699);
nand U2716 (N_2716,N_2646,N_2672);
and U2717 (N_2717,N_2653,N_2665);
nand U2718 (N_2718,N_2697,N_2669);
nor U2719 (N_2719,N_2659,N_2651);
nand U2720 (N_2720,N_2684,N_2645);
and U2721 (N_2721,N_2682,N_2668);
and U2722 (N_2722,N_2656,N_2660);
xnor U2723 (N_2723,N_2647,N_2640);
and U2724 (N_2724,N_2642,N_2674);
nor U2725 (N_2725,N_2687,N_2685);
nor U2726 (N_2726,N_2680,N_2652);
and U2727 (N_2727,N_2641,N_2692);
nor U2728 (N_2728,N_2683,N_2649);
and U2729 (N_2729,N_2643,N_2654);
and U2730 (N_2730,N_2685,N_2677);
or U2731 (N_2731,N_2687,N_2644);
and U2732 (N_2732,N_2671,N_2672);
nor U2733 (N_2733,N_2688,N_2645);
nand U2734 (N_2734,N_2650,N_2669);
nor U2735 (N_2735,N_2657,N_2669);
and U2736 (N_2736,N_2649,N_2644);
nor U2737 (N_2737,N_2693,N_2672);
nand U2738 (N_2738,N_2644,N_2671);
and U2739 (N_2739,N_2695,N_2687);
nand U2740 (N_2740,N_2647,N_2685);
nor U2741 (N_2741,N_2674,N_2699);
and U2742 (N_2742,N_2657,N_2662);
or U2743 (N_2743,N_2656,N_2684);
nor U2744 (N_2744,N_2672,N_2681);
or U2745 (N_2745,N_2668,N_2687);
or U2746 (N_2746,N_2671,N_2679);
nor U2747 (N_2747,N_2684,N_2654);
nand U2748 (N_2748,N_2662,N_2690);
nand U2749 (N_2749,N_2699,N_2649);
or U2750 (N_2750,N_2657,N_2697);
nor U2751 (N_2751,N_2652,N_2653);
nor U2752 (N_2752,N_2684,N_2672);
and U2753 (N_2753,N_2653,N_2697);
nor U2754 (N_2754,N_2658,N_2661);
nand U2755 (N_2755,N_2679,N_2685);
xor U2756 (N_2756,N_2661,N_2670);
or U2757 (N_2757,N_2664,N_2659);
nor U2758 (N_2758,N_2658,N_2671);
or U2759 (N_2759,N_2694,N_2675);
nand U2760 (N_2760,N_2726,N_2722);
nor U2761 (N_2761,N_2728,N_2719);
nand U2762 (N_2762,N_2718,N_2756);
and U2763 (N_2763,N_2725,N_2729);
nor U2764 (N_2764,N_2702,N_2731);
or U2765 (N_2765,N_2710,N_2704);
xnor U2766 (N_2766,N_2752,N_2734);
or U2767 (N_2767,N_2724,N_2737);
nand U2768 (N_2768,N_2759,N_2732);
nor U2769 (N_2769,N_2708,N_2720);
or U2770 (N_2770,N_2730,N_2715);
nor U2771 (N_2771,N_2711,N_2735);
or U2772 (N_2772,N_2745,N_2712);
or U2773 (N_2773,N_2705,N_2703);
and U2774 (N_2774,N_2717,N_2709);
nor U2775 (N_2775,N_2738,N_2733);
or U2776 (N_2776,N_2714,N_2706);
nor U2777 (N_2777,N_2723,N_2751);
nand U2778 (N_2778,N_2755,N_2749);
nand U2779 (N_2779,N_2739,N_2707);
and U2780 (N_2780,N_2750,N_2713);
or U2781 (N_2781,N_2742,N_2741);
nand U2782 (N_2782,N_2736,N_2757);
nand U2783 (N_2783,N_2753,N_2700);
nor U2784 (N_2784,N_2746,N_2701);
nor U2785 (N_2785,N_2748,N_2747);
nand U2786 (N_2786,N_2744,N_2716);
nor U2787 (N_2787,N_2727,N_2743);
and U2788 (N_2788,N_2740,N_2721);
and U2789 (N_2789,N_2754,N_2758);
and U2790 (N_2790,N_2712,N_2758);
or U2791 (N_2791,N_2724,N_2705);
nand U2792 (N_2792,N_2759,N_2746);
and U2793 (N_2793,N_2752,N_2712);
and U2794 (N_2794,N_2708,N_2723);
and U2795 (N_2795,N_2739,N_2754);
or U2796 (N_2796,N_2739,N_2745);
or U2797 (N_2797,N_2706,N_2755);
and U2798 (N_2798,N_2747,N_2704);
or U2799 (N_2799,N_2711,N_2748);
nor U2800 (N_2800,N_2704,N_2753);
nand U2801 (N_2801,N_2751,N_2717);
nand U2802 (N_2802,N_2748,N_2722);
or U2803 (N_2803,N_2737,N_2732);
nor U2804 (N_2804,N_2757,N_2702);
xor U2805 (N_2805,N_2734,N_2722);
and U2806 (N_2806,N_2703,N_2711);
nor U2807 (N_2807,N_2709,N_2732);
nor U2808 (N_2808,N_2743,N_2713);
and U2809 (N_2809,N_2736,N_2709);
or U2810 (N_2810,N_2727,N_2748);
nor U2811 (N_2811,N_2711,N_2704);
or U2812 (N_2812,N_2741,N_2739);
nor U2813 (N_2813,N_2715,N_2735);
or U2814 (N_2814,N_2721,N_2702);
nand U2815 (N_2815,N_2714,N_2710);
and U2816 (N_2816,N_2719,N_2732);
or U2817 (N_2817,N_2735,N_2754);
nand U2818 (N_2818,N_2713,N_2749);
nor U2819 (N_2819,N_2714,N_2753);
or U2820 (N_2820,N_2797,N_2761);
or U2821 (N_2821,N_2765,N_2808);
nand U2822 (N_2822,N_2795,N_2784);
or U2823 (N_2823,N_2767,N_2774);
xnor U2824 (N_2824,N_2769,N_2811);
and U2825 (N_2825,N_2790,N_2816);
nor U2826 (N_2826,N_2799,N_2813);
xnor U2827 (N_2827,N_2789,N_2760);
and U2828 (N_2828,N_2776,N_2794);
or U2829 (N_2829,N_2764,N_2815);
xor U2830 (N_2830,N_2768,N_2818);
nand U2831 (N_2831,N_2788,N_2806);
nor U2832 (N_2832,N_2773,N_2819);
nand U2833 (N_2833,N_2775,N_2785);
nor U2834 (N_2834,N_2772,N_2762);
nand U2835 (N_2835,N_2781,N_2771);
or U2836 (N_2836,N_2804,N_2792);
nand U2837 (N_2837,N_2779,N_2809);
and U2838 (N_2838,N_2777,N_2805);
or U2839 (N_2839,N_2817,N_2791);
nor U2840 (N_2840,N_2778,N_2798);
and U2841 (N_2841,N_2770,N_2814);
or U2842 (N_2842,N_2793,N_2807);
or U2843 (N_2843,N_2783,N_2796);
nand U2844 (N_2844,N_2800,N_2812);
nand U2845 (N_2845,N_2802,N_2787);
nor U2846 (N_2846,N_2786,N_2766);
and U2847 (N_2847,N_2803,N_2810);
nand U2848 (N_2848,N_2780,N_2782);
and U2849 (N_2849,N_2763,N_2801);
or U2850 (N_2850,N_2785,N_2788);
nand U2851 (N_2851,N_2785,N_2770);
and U2852 (N_2852,N_2771,N_2795);
and U2853 (N_2853,N_2794,N_2790);
nand U2854 (N_2854,N_2792,N_2809);
or U2855 (N_2855,N_2817,N_2803);
or U2856 (N_2856,N_2780,N_2794);
nor U2857 (N_2857,N_2792,N_2786);
and U2858 (N_2858,N_2760,N_2768);
and U2859 (N_2859,N_2790,N_2786);
nand U2860 (N_2860,N_2771,N_2773);
nand U2861 (N_2861,N_2819,N_2797);
or U2862 (N_2862,N_2766,N_2797);
and U2863 (N_2863,N_2764,N_2793);
nor U2864 (N_2864,N_2788,N_2767);
nor U2865 (N_2865,N_2811,N_2772);
nor U2866 (N_2866,N_2763,N_2762);
nor U2867 (N_2867,N_2774,N_2810);
and U2868 (N_2868,N_2774,N_2769);
nor U2869 (N_2869,N_2783,N_2792);
nand U2870 (N_2870,N_2800,N_2775);
nand U2871 (N_2871,N_2761,N_2763);
or U2872 (N_2872,N_2790,N_2769);
or U2873 (N_2873,N_2766,N_2793);
xnor U2874 (N_2874,N_2809,N_2781);
nand U2875 (N_2875,N_2798,N_2811);
nor U2876 (N_2876,N_2819,N_2817);
nand U2877 (N_2877,N_2779,N_2799);
xor U2878 (N_2878,N_2786,N_2777);
xor U2879 (N_2879,N_2775,N_2811);
and U2880 (N_2880,N_2829,N_2824);
and U2881 (N_2881,N_2867,N_2827);
or U2882 (N_2882,N_2865,N_2838);
nor U2883 (N_2883,N_2848,N_2851);
nor U2884 (N_2884,N_2861,N_2855);
nor U2885 (N_2885,N_2871,N_2847);
and U2886 (N_2886,N_2868,N_2879);
or U2887 (N_2887,N_2832,N_2856);
nand U2888 (N_2888,N_2821,N_2872);
and U2889 (N_2889,N_2876,N_2869);
nand U2890 (N_2890,N_2870,N_2839);
nor U2891 (N_2891,N_2852,N_2822);
and U2892 (N_2892,N_2860,N_2874);
or U2893 (N_2893,N_2875,N_2825);
nor U2894 (N_2894,N_2842,N_2828);
or U2895 (N_2895,N_2830,N_2864);
nor U2896 (N_2896,N_2853,N_2849);
nor U2897 (N_2897,N_2857,N_2863);
and U2898 (N_2898,N_2854,N_2844);
and U2899 (N_2899,N_2820,N_2834);
and U2900 (N_2900,N_2878,N_2877);
nor U2901 (N_2901,N_2833,N_2850);
or U2902 (N_2902,N_2873,N_2826);
nor U2903 (N_2903,N_2835,N_2836);
nand U2904 (N_2904,N_2866,N_2845);
nor U2905 (N_2905,N_2846,N_2823);
and U2906 (N_2906,N_2843,N_2831);
nor U2907 (N_2907,N_2840,N_2837);
and U2908 (N_2908,N_2862,N_2841);
nor U2909 (N_2909,N_2858,N_2859);
and U2910 (N_2910,N_2839,N_2822);
nor U2911 (N_2911,N_2835,N_2876);
and U2912 (N_2912,N_2830,N_2877);
or U2913 (N_2913,N_2840,N_2875);
nor U2914 (N_2914,N_2842,N_2836);
or U2915 (N_2915,N_2839,N_2844);
and U2916 (N_2916,N_2874,N_2873);
nand U2917 (N_2917,N_2871,N_2858);
nor U2918 (N_2918,N_2875,N_2830);
or U2919 (N_2919,N_2852,N_2845);
nor U2920 (N_2920,N_2857,N_2830);
nor U2921 (N_2921,N_2878,N_2828);
or U2922 (N_2922,N_2870,N_2875);
or U2923 (N_2923,N_2834,N_2824);
or U2924 (N_2924,N_2864,N_2878);
and U2925 (N_2925,N_2839,N_2832);
and U2926 (N_2926,N_2865,N_2866);
xnor U2927 (N_2927,N_2836,N_2877);
nor U2928 (N_2928,N_2851,N_2841);
and U2929 (N_2929,N_2830,N_2860);
or U2930 (N_2930,N_2855,N_2839);
or U2931 (N_2931,N_2823,N_2824);
nor U2932 (N_2932,N_2857,N_2843);
and U2933 (N_2933,N_2851,N_2867);
or U2934 (N_2934,N_2879,N_2823);
and U2935 (N_2935,N_2839,N_2858);
xor U2936 (N_2936,N_2827,N_2835);
nor U2937 (N_2937,N_2830,N_2835);
or U2938 (N_2938,N_2845,N_2862);
nor U2939 (N_2939,N_2863,N_2870);
nor U2940 (N_2940,N_2906,N_2935);
and U2941 (N_2941,N_2890,N_2910);
and U2942 (N_2942,N_2908,N_2916);
xnor U2943 (N_2943,N_2907,N_2887);
and U2944 (N_2944,N_2882,N_2900);
nand U2945 (N_2945,N_2903,N_2893);
and U2946 (N_2946,N_2939,N_2904);
nor U2947 (N_2947,N_2923,N_2920);
or U2948 (N_2948,N_2886,N_2896);
or U2949 (N_2949,N_2924,N_2926);
and U2950 (N_2950,N_2913,N_2899);
and U2951 (N_2951,N_2883,N_2929);
xor U2952 (N_2952,N_2921,N_2925);
nand U2953 (N_2953,N_2889,N_2895);
and U2954 (N_2954,N_2909,N_2898);
or U2955 (N_2955,N_2880,N_2905);
or U2956 (N_2956,N_2902,N_2881);
or U2957 (N_2957,N_2938,N_2930);
or U2958 (N_2958,N_2927,N_2892);
or U2959 (N_2959,N_2922,N_2936);
nand U2960 (N_2960,N_2928,N_2937);
nor U2961 (N_2961,N_2931,N_2911);
and U2962 (N_2962,N_2919,N_2885);
nor U2963 (N_2963,N_2917,N_2891);
or U2964 (N_2964,N_2901,N_2934);
nand U2965 (N_2965,N_2912,N_2918);
and U2966 (N_2966,N_2884,N_2933);
nor U2967 (N_2967,N_2932,N_2888);
or U2968 (N_2968,N_2897,N_2915);
and U2969 (N_2969,N_2914,N_2894);
and U2970 (N_2970,N_2932,N_2904);
nand U2971 (N_2971,N_2884,N_2901);
nor U2972 (N_2972,N_2902,N_2915);
nor U2973 (N_2973,N_2881,N_2899);
or U2974 (N_2974,N_2922,N_2905);
nand U2975 (N_2975,N_2893,N_2928);
or U2976 (N_2976,N_2881,N_2916);
nand U2977 (N_2977,N_2905,N_2914);
and U2978 (N_2978,N_2921,N_2916);
or U2979 (N_2979,N_2927,N_2897);
and U2980 (N_2980,N_2931,N_2916);
nor U2981 (N_2981,N_2910,N_2884);
or U2982 (N_2982,N_2939,N_2889);
and U2983 (N_2983,N_2919,N_2908);
and U2984 (N_2984,N_2925,N_2937);
or U2985 (N_2985,N_2889,N_2899);
nor U2986 (N_2986,N_2935,N_2903);
nand U2987 (N_2987,N_2896,N_2931);
nor U2988 (N_2988,N_2930,N_2886);
or U2989 (N_2989,N_2909,N_2923);
and U2990 (N_2990,N_2888,N_2924);
nand U2991 (N_2991,N_2924,N_2936);
nand U2992 (N_2992,N_2936,N_2930);
nor U2993 (N_2993,N_2883,N_2934);
nor U2994 (N_2994,N_2893,N_2897);
and U2995 (N_2995,N_2906,N_2883);
nand U2996 (N_2996,N_2912,N_2900);
nor U2997 (N_2997,N_2911,N_2909);
nor U2998 (N_2998,N_2892,N_2915);
nand U2999 (N_2999,N_2923,N_2933);
nand UO_0 (O_0,N_2966,N_2970);
and UO_1 (O_1,N_2993,N_2995);
nand UO_2 (O_2,N_2945,N_2941);
nor UO_3 (O_3,N_2991,N_2997);
or UO_4 (O_4,N_2949,N_2983);
or UO_5 (O_5,N_2984,N_2990);
and UO_6 (O_6,N_2994,N_2962);
nor UO_7 (O_7,N_2959,N_2987);
nor UO_8 (O_8,N_2940,N_2960);
nor UO_9 (O_9,N_2974,N_2971);
nand UO_10 (O_10,N_2948,N_2986);
or UO_11 (O_11,N_2968,N_2982);
and UO_12 (O_12,N_2975,N_2957);
nor UO_13 (O_13,N_2951,N_2965);
or UO_14 (O_14,N_2950,N_2953);
nand UO_15 (O_15,N_2978,N_2947);
and UO_16 (O_16,N_2967,N_2980);
nand UO_17 (O_17,N_2943,N_2979);
or UO_18 (O_18,N_2973,N_2976);
or UO_19 (O_19,N_2996,N_2998);
and UO_20 (O_20,N_2946,N_2954);
nor UO_21 (O_21,N_2989,N_2958);
or UO_22 (O_22,N_2942,N_2964);
or UO_23 (O_23,N_2963,N_2952);
nand UO_24 (O_24,N_2961,N_2977);
and UO_25 (O_25,N_2944,N_2985);
and UO_26 (O_26,N_2969,N_2999);
nand UO_27 (O_27,N_2955,N_2972);
nor UO_28 (O_28,N_2988,N_2981);
nor UO_29 (O_29,N_2956,N_2992);
nand UO_30 (O_30,N_2984,N_2974);
or UO_31 (O_31,N_2995,N_2957);
and UO_32 (O_32,N_2969,N_2973);
nand UO_33 (O_33,N_2952,N_2993);
or UO_34 (O_34,N_2988,N_2954);
nor UO_35 (O_35,N_2947,N_2977);
or UO_36 (O_36,N_2949,N_2977);
nand UO_37 (O_37,N_2973,N_2943);
or UO_38 (O_38,N_2985,N_2983);
nor UO_39 (O_39,N_2951,N_2981);
nand UO_40 (O_40,N_2972,N_2968);
and UO_41 (O_41,N_2987,N_2993);
and UO_42 (O_42,N_2951,N_2966);
xor UO_43 (O_43,N_2979,N_2972);
and UO_44 (O_44,N_2954,N_2999);
nor UO_45 (O_45,N_2980,N_2992);
or UO_46 (O_46,N_2967,N_2969);
and UO_47 (O_47,N_2966,N_2964);
or UO_48 (O_48,N_2995,N_2965);
and UO_49 (O_49,N_2967,N_2965);
nor UO_50 (O_50,N_2998,N_2990);
and UO_51 (O_51,N_2982,N_2944);
and UO_52 (O_52,N_2980,N_2987);
and UO_53 (O_53,N_2976,N_2968);
or UO_54 (O_54,N_2987,N_2978);
or UO_55 (O_55,N_2967,N_2951);
and UO_56 (O_56,N_2972,N_2993);
or UO_57 (O_57,N_2961,N_2955);
nand UO_58 (O_58,N_2976,N_2979);
or UO_59 (O_59,N_2977,N_2972);
and UO_60 (O_60,N_2992,N_2970);
and UO_61 (O_61,N_2943,N_2974);
nor UO_62 (O_62,N_2945,N_2948);
or UO_63 (O_63,N_2997,N_2979);
nand UO_64 (O_64,N_2978,N_2988);
or UO_65 (O_65,N_2978,N_2994);
nor UO_66 (O_66,N_2975,N_2996);
nor UO_67 (O_67,N_2988,N_2947);
and UO_68 (O_68,N_2986,N_2983);
and UO_69 (O_69,N_2941,N_2975);
and UO_70 (O_70,N_2950,N_2958);
nor UO_71 (O_71,N_2997,N_2944);
nor UO_72 (O_72,N_2993,N_2965);
and UO_73 (O_73,N_2980,N_2963);
or UO_74 (O_74,N_2994,N_2965);
or UO_75 (O_75,N_2946,N_2966);
nand UO_76 (O_76,N_2943,N_2982);
nand UO_77 (O_77,N_2990,N_2969);
or UO_78 (O_78,N_2964,N_2994);
or UO_79 (O_79,N_2957,N_2973);
and UO_80 (O_80,N_2963,N_2970);
nand UO_81 (O_81,N_2960,N_2982);
nor UO_82 (O_82,N_2989,N_2991);
or UO_83 (O_83,N_2955,N_2950);
and UO_84 (O_84,N_2997,N_2972);
nand UO_85 (O_85,N_2968,N_2998);
nor UO_86 (O_86,N_2958,N_2966);
or UO_87 (O_87,N_2970,N_2942);
or UO_88 (O_88,N_2983,N_2989);
nor UO_89 (O_89,N_2959,N_2949);
and UO_90 (O_90,N_2994,N_2942);
and UO_91 (O_91,N_2956,N_2978);
nand UO_92 (O_92,N_2940,N_2955);
and UO_93 (O_93,N_2999,N_2995);
nand UO_94 (O_94,N_2989,N_2942);
and UO_95 (O_95,N_2965,N_2952);
nand UO_96 (O_96,N_2949,N_2958);
xnor UO_97 (O_97,N_2974,N_2996);
or UO_98 (O_98,N_2958,N_2975);
and UO_99 (O_99,N_2948,N_2953);
or UO_100 (O_100,N_2962,N_2947);
or UO_101 (O_101,N_2985,N_2941);
and UO_102 (O_102,N_2963,N_2981);
or UO_103 (O_103,N_2947,N_2967);
and UO_104 (O_104,N_2950,N_2956);
or UO_105 (O_105,N_2954,N_2995);
nor UO_106 (O_106,N_2981,N_2994);
nor UO_107 (O_107,N_2960,N_2958);
or UO_108 (O_108,N_2943,N_2950);
and UO_109 (O_109,N_2989,N_2975);
nor UO_110 (O_110,N_2946,N_2982);
nand UO_111 (O_111,N_2989,N_2998);
or UO_112 (O_112,N_2957,N_2960);
and UO_113 (O_113,N_2990,N_2989);
nand UO_114 (O_114,N_2980,N_2983);
nand UO_115 (O_115,N_2970,N_2973);
nor UO_116 (O_116,N_2989,N_2951);
nor UO_117 (O_117,N_2999,N_2993);
nor UO_118 (O_118,N_2994,N_2941);
or UO_119 (O_119,N_2946,N_2969);
nand UO_120 (O_120,N_2975,N_2976);
nand UO_121 (O_121,N_2950,N_2980);
or UO_122 (O_122,N_2975,N_2970);
nor UO_123 (O_123,N_2951,N_2952);
or UO_124 (O_124,N_2957,N_2976);
nor UO_125 (O_125,N_2998,N_2977);
or UO_126 (O_126,N_2963,N_2999);
or UO_127 (O_127,N_2945,N_2962);
nor UO_128 (O_128,N_2950,N_2962);
and UO_129 (O_129,N_2980,N_2974);
nand UO_130 (O_130,N_2954,N_2945);
nor UO_131 (O_131,N_2980,N_2949);
nor UO_132 (O_132,N_2958,N_2961);
or UO_133 (O_133,N_2952,N_2980);
and UO_134 (O_134,N_2981,N_2968);
and UO_135 (O_135,N_2995,N_2941);
and UO_136 (O_136,N_2980,N_2978);
or UO_137 (O_137,N_2946,N_2989);
nand UO_138 (O_138,N_2959,N_2968);
or UO_139 (O_139,N_2991,N_2980);
and UO_140 (O_140,N_2944,N_2972);
or UO_141 (O_141,N_2990,N_2961);
or UO_142 (O_142,N_2970,N_2987);
nor UO_143 (O_143,N_2975,N_2987);
nand UO_144 (O_144,N_2973,N_2951);
nor UO_145 (O_145,N_2964,N_2973);
nand UO_146 (O_146,N_2978,N_2975);
and UO_147 (O_147,N_2985,N_2950);
nand UO_148 (O_148,N_2965,N_2972);
and UO_149 (O_149,N_2960,N_2971);
nor UO_150 (O_150,N_2985,N_2981);
nor UO_151 (O_151,N_2992,N_2958);
nor UO_152 (O_152,N_2961,N_2947);
or UO_153 (O_153,N_2992,N_2955);
and UO_154 (O_154,N_2979,N_2995);
nor UO_155 (O_155,N_2992,N_2946);
nand UO_156 (O_156,N_2950,N_2998);
nand UO_157 (O_157,N_2980,N_2957);
nor UO_158 (O_158,N_2963,N_2967);
xor UO_159 (O_159,N_2979,N_2954);
nor UO_160 (O_160,N_2954,N_2952);
or UO_161 (O_161,N_2985,N_2971);
or UO_162 (O_162,N_2978,N_2996);
or UO_163 (O_163,N_2969,N_2985);
nand UO_164 (O_164,N_2964,N_2953);
and UO_165 (O_165,N_2946,N_2959);
xnor UO_166 (O_166,N_2979,N_2999);
nand UO_167 (O_167,N_2981,N_2982);
nand UO_168 (O_168,N_2961,N_2978);
and UO_169 (O_169,N_2982,N_2983);
nor UO_170 (O_170,N_2959,N_2952);
nor UO_171 (O_171,N_2997,N_2967);
and UO_172 (O_172,N_2993,N_2986);
and UO_173 (O_173,N_2958,N_2988);
nand UO_174 (O_174,N_2969,N_2963);
nor UO_175 (O_175,N_2960,N_2967);
nor UO_176 (O_176,N_2977,N_2957);
nor UO_177 (O_177,N_2977,N_2973);
nor UO_178 (O_178,N_2965,N_2978);
nor UO_179 (O_179,N_2985,N_2953);
nand UO_180 (O_180,N_2997,N_2955);
or UO_181 (O_181,N_2950,N_2966);
and UO_182 (O_182,N_2998,N_2963);
nor UO_183 (O_183,N_2989,N_2945);
xnor UO_184 (O_184,N_2992,N_2994);
or UO_185 (O_185,N_2989,N_2970);
nand UO_186 (O_186,N_2990,N_2968);
nand UO_187 (O_187,N_2979,N_2969);
nor UO_188 (O_188,N_2948,N_2951);
and UO_189 (O_189,N_2969,N_2960);
and UO_190 (O_190,N_2942,N_2968);
xnor UO_191 (O_191,N_2978,N_2984);
nor UO_192 (O_192,N_2951,N_2959);
nand UO_193 (O_193,N_2990,N_2970);
nand UO_194 (O_194,N_2984,N_2989);
and UO_195 (O_195,N_2962,N_2986);
and UO_196 (O_196,N_2967,N_2994);
nor UO_197 (O_197,N_2977,N_2990);
or UO_198 (O_198,N_2947,N_2970);
and UO_199 (O_199,N_2976,N_2996);
and UO_200 (O_200,N_2958,N_2986);
nand UO_201 (O_201,N_2989,N_2947);
xor UO_202 (O_202,N_2992,N_2940);
or UO_203 (O_203,N_2942,N_2958);
and UO_204 (O_204,N_2987,N_2998);
or UO_205 (O_205,N_2969,N_2943);
or UO_206 (O_206,N_2953,N_2997);
or UO_207 (O_207,N_2990,N_2996);
and UO_208 (O_208,N_2976,N_2944);
and UO_209 (O_209,N_2986,N_2970);
or UO_210 (O_210,N_2986,N_2960);
and UO_211 (O_211,N_2971,N_2973);
or UO_212 (O_212,N_2972,N_2992);
and UO_213 (O_213,N_2983,N_2996);
nand UO_214 (O_214,N_2945,N_2959);
nor UO_215 (O_215,N_2981,N_2970);
nor UO_216 (O_216,N_2956,N_2969);
or UO_217 (O_217,N_2965,N_2962);
or UO_218 (O_218,N_2949,N_2964);
xor UO_219 (O_219,N_2947,N_2951);
nand UO_220 (O_220,N_2941,N_2968);
or UO_221 (O_221,N_2953,N_2965);
and UO_222 (O_222,N_2979,N_2996);
or UO_223 (O_223,N_2963,N_2971);
nand UO_224 (O_224,N_2991,N_2979);
xnor UO_225 (O_225,N_2981,N_2965);
and UO_226 (O_226,N_2997,N_2999);
or UO_227 (O_227,N_2983,N_2977);
or UO_228 (O_228,N_2953,N_2958);
and UO_229 (O_229,N_2982,N_2964);
or UO_230 (O_230,N_2966,N_2957);
nand UO_231 (O_231,N_2995,N_2971);
or UO_232 (O_232,N_2980,N_2990);
nand UO_233 (O_233,N_2988,N_2953);
or UO_234 (O_234,N_2966,N_2995);
nand UO_235 (O_235,N_2977,N_2954);
nor UO_236 (O_236,N_2997,N_2980);
nor UO_237 (O_237,N_2954,N_2982);
nor UO_238 (O_238,N_2956,N_2998);
and UO_239 (O_239,N_2973,N_2978);
or UO_240 (O_240,N_2991,N_2966);
and UO_241 (O_241,N_2976,N_2992);
or UO_242 (O_242,N_2985,N_2948);
xnor UO_243 (O_243,N_2999,N_2972);
or UO_244 (O_244,N_2990,N_2965);
and UO_245 (O_245,N_2996,N_2961);
or UO_246 (O_246,N_2975,N_2993);
nor UO_247 (O_247,N_2979,N_2941);
or UO_248 (O_248,N_2983,N_2940);
and UO_249 (O_249,N_2991,N_2990);
and UO_250 (O_250,N_2996,N_2994);
or UO_251 (O_251,N_2997,N_2983);
nor UO_252 (O_252,N_2964,N_2945);
nand UO_253 (O_253,N_2950,N_2975);
xor UO_254 (O_254,N_2964,N_2971);
and UO_255 (O_255,N_2998,N_2945);
nor UO_256 (O_256,N_2947,N_2941);
and UO_257 (O_257,N_2999,N_2944);
nand UO_258 (O_258,N_2941,N_2967);
nand UO_259 (O_259,N_2990,N_2997);
or UO_260 (O_260,N_2966,N_2963);
and UO_261 (O_261,N_2941,N_2973);
or UO_262 (O_262,N_2990,N_2957);
or UO_263 (O_263,N_2955,N_2981);
nor UO_264 (O_264,N_2993,N_2950);
and UO_265 (O_265,N_2967,N_2999);
and UO_266 (O_266,N_2989,N_2977);
and UO_267 (O_267,N_2945,N_2955);
and UO_268 (O_268,N_2982,N_2973);
and UO_269 (O_269,N_2968,N_2969);
or UO_270 (O_270,N_2997,N_2995);
nor UO_271 (O_271,N_2963,N_2975);
and UO_272 (O_272,N_2948,N_2962);
and UO_273 (O_273,N_2959,N_2984);
and UO_274 (O_274,N_2942,N_2961);
or UO_275 (O_275,N_2993,N_2951);
xor UO_276 (O_276,N_2985,N_2977);
or UO_277 (O_277,N_2984,N_2962);
nor UO_278 (O_278,N_2974,N_2990);
or UO_279 (O_279,N_2956,N_2985);
or UO_280 (O_280,N_2947,N_2994);
or UO_281 (O_281,N_2952,N_2964);
nand UO_282 (O_282,N_2997,N_2975);
and UO_283 (O_283,N_2988,N_2997);
nand UO_284 (O_284,N_2974,N_2960);
nand UO_285 (O_285,N_2956,N_2987);
or UO_286 (O_286,N_2996,N_2949);
or UO_287 (O_287,N_2966,N_2982);
or UO_288 (O_288,N_2988,N_2995);
nor UO_289 (O_289,N_2959,N_2989);
nand UO_290 (O_290,N_2981,N_2993);
or UO_291 (O_291,N_2980,N_2941);
nor UO_292 (O_292,N_2988,N_2960);
and UO_293 (O_293,N_2961,N_2948);
or UO_294 (O_294,N_2978,N_2946);
nand UO_295 (O_295,N_2946,N_2977);
and UO_296 (O_296,N_2991,N_2967);
and UO_297 (O_297,N_2952,N_2957);
or UO_298 (O_298,N_2958,N_2963);
or UO_299 (O_299,N_2956,N_2944);
nor UO_300 (O_300,N_2959,N_2998);
nand UO_301 (O_301,N_2986,N_2992);
nand UO_302 (O_302,N_2995,N_2947);
and UO_303 (O_303,N_2944,N_2967);
nand UO_304 (O_304,N_2978,N_2958);
nand UO_305 (O_305,N_2940,N_2944);
nor UO_306 (O_306,N_2984,N_2993);
nand UO_307 (O_307,N_2993,N_2961);
nand UO_308 (O_308,N_2977,N_2950);
or UO_309 (O_309,N_2985,N_2967);
nor UO_310 (O_310,N_2990,N_2952);
and UO_311 (O_311,N_2963,N_2991);
nor UO_312 (O_312,N_2978,N_2955);
or UO_313 (O_313,N_2961,N_2989);
nor UO_314 (O_314,N_2951,N_2946);
nor UO_315 (O_315,N_2997,N_2964);
and UO_316 (O_316,N_2962,N_2998);
nor UO_317 (O_317,N_2961,N_2988);
xnor UO_318 (O_318,N_2960,N_2959);
nor UO_319 (O_319,N_2982,N_2953);
nor UO_320 (O_320,N_2955,N_2974);
nand UO_321 (O_321,N_2983,N_2970);
or UO_322 (O_322,N_2985,N_2990);
nand UO_323 (O_323,N_2979,N_2955);
nor UO_324 (O_324,N_2959,N_2955);
and UO_325 (O_325,N_2966,N_2968);
nor UO_326 (O_326,N_2947,N_2986);
nor UO_327 (O_327,N_2940,N_2956);
or UO_328 (O_328,N_2950,N_2944);
nand UO_329 (O_329,N_2957,N_2991);
and UO_330 (O_330,N_2976,N_2984);
nand UO_331 (O_331,N_2973,N_2988);
or UO_332 (O_332,N_2943,N_2989);
nand UO_333 (O_333,N_2972,N_2956);
and UO_334 (O_334,N_2972,N_2957);
nor UO_335 (O_335,N_2961,N_2952);
or UO_336 (O_336,N_2977,N_2980);
or UO_337 (O_337,N_2957,N_2988);
and UO_338 (O_338,N_2994,N_2982);
or UO_339 (O_339,N_2981,N_2950);
or UO_340 (O_340,N_2965,N_2947);
nor UO_341 (O_341,N_2987,N_2989);
and UO_342 (O_342,N_2947,N_2950);
nor UO_343 (O_343,N_2990,N_2979);
or UO_344 (O_344,N_2974,N_2978);
or UO_345 (O_345,N_2985,N_2972);
or UO_346 (O_346,N_2967,N_2990);
or UO_347 (O_347,N_2969,N_2952);
or UO_348 (O_348,N_2982,N_2984);
or UO_349 (O_349,N_2981,N_2986);
and UO_350 (O_350,N_2950,N_2969);
nor UO_351 (O_351,N_2956,N_2965);
and UO_352 (O_352,N_2990,N_2999);
and UO_353 (O_353,N_2943,N_2955);
nand UO_354 (O_354,N_2943,N_2970);
xor UO_355 (O_355,N_2999,N_2981);
nor UO_356 (O_356,N_2996,N_2981);
nor UO_357 (O_357,N_2961,N_2986);
nor UO_358 (O_358,N_2943,N_2986);
or UO_359 (O_359,N_2969,N_2962);
or UO_360 (O_360,N_2953,N_2974);
nor UO_361 (O_361,N_2995,N_2951);
and UO_362 (O_362,N_2976,N_2967);
or UO_363 (O_363,N_2958,N_2976);
nor UO_364 (O_364,N_2971,N_2984);
nand UO_365 (O_365,N_2954,N_2949);
nor UO_366 (O_366,N_2984,N_2966);
nor UO_367 (O_367,N_2975,N_2994);
nor UO_368 (O_368,N_2987,N_2957);
and UO_369 (O_369,N_2947,N_2952);
nor UO_370 (O_370,N_2947,N_2946);
nand UO_371 (O_371,N_2969,N_2958);
and UO_372 (O_372,N_2974,N_2986);
or UO_373 (O_373,N_2962,N_2977);
nand UO_374 (O_374,N_2962,N_2941);
or UO_375 (O_375,N_2959,N_2980);
and UO_376 (O_376,N_2989,N_2953);
or UO_377 (O_377,N_2948,N_2987);
nand UO_378 (O_378,N_2946,N_2948);
nor UO_379 (O_379,N_2965,N_2983);
and UO_380 (O_380,N_2965,N_2979);
nand UO_381 (O_381,N_2975,N_2942);
and UO_382 (O_382,N_2954,N_2961);
and UO_383 (O_383,N_2945,N_2975);
nand UO_384 (O_384,N_2955,N_2984);
and UO_385 (O_385,N_2958,N_2993);
nand UO_386 (O_386,N_2974,N_2964);
or UO_387 (O_387,N_2946,N_2974);
nand UO_388 (O_388,N_2950,N_2990);
nor UO_389 (O_389,N_2975,N_2977);
nand UO_390 (O_390,N_2944,N_2979);
nor UO_391 (O_391,N_2950,N_2959);
nor UO_392 (O_392,N_2990,N_2958);
nand UO_393 (O_393,N_2979,N_2992);
and UO_394 (O_394,N_2991,N_2981);
or UO_395 (O_395,N_2984,N_2960);
and UO_396 (O_396,N_2942,N_2996);
xor UO_397 (O_397,N_2993,N_2955);
or UO_398 (O_398,N_2973,N_2966);
or UO_399 (O_399,N_2949,N_2956);
nand UO_400 (O_400,N_2969,N_2976);
nor UO_401 (O_401,N_2959,N_2957);
and UO_402 (O_402,N_2965,N_2943);
nand UO_403 (O_403,N_2979,N_2964);
nand UO_404 (O_404,N_2964,N_2984);
nor UO_405 (O_405,N_2954,N_2950);
nor UO_406 (O_406,N_2957,N_2984);
nor UO_407 (O_407,N_2977,N_2966);
nor UO_408 (O_408,N_2963,N_2940);
nor UO_409 (O_409,N_2967,N_2988);
or UO_410 (O_410,N_2944,N_2984);
or UO_411 (O_411,N_2980,N_2996);
nor UO_412 (O_412,N_2961,N_2979);
nand UO_413 (O_413,N_2941,N_2960);
xor UO_414 (O_414,N_2943,N_2942);
nor UO_415 (O_415,N_2956,N_2963);
and UO_416 (O_416,N_2950,N_2942);
nor UO_417 (O_417,N_2980,N_2995);
nand UO_418 (O_418,N_2980,N_2944);
nor UO_419 (O_419,N_2988,N_2974);
nor UO_420 (O_420,N_2961,N_2994);
and UO_421 (O_421,N_2975,N_2981);
nand UO_422 (O_422,N_2982,N_2978);
or UO_423 (O_423,N_2953,N_2949);
or UO_424 (O_424,N_2982,N_2995);
and UO_425 (O_425,N_2962,N_2956);
and UO_426 (O_426,N_2977,N_2971);
or UO_427 (O_427,N_2952,N_2966);
nand UO_428 (O_428,N_2980,N_2971);
nor UO_429 (O_429,N_2975,N_2982);
and UO_430 (O_430,N_2956,N_2989);
nor UO_431 (O_431,N_2974,N_2951);
or UO_432 (O_432,N_2964,N_2983);
or UO_433 (O_433,N_2996,N_2992);
and UO_434 (O_434,N_2996,N_2946);
nor UO_435 (O_435,N_2996,N_2951);
and UO_436 (O_436,N_2989,N_2944);
nor UO_437 (O_437,N_2998,N_2952);
nand UO_438 (O_438,N_2944,N_2981);
and UO_439 (O_439,N_2975,N_2984);
nor UO_440 (O_440,N_2991,N_2950);
or UO_441 (O_441,N_2968,N_2995);
and UO_442 (O_442,N_2953,N_2952);
nor UO_443 (O_443,N_2980,N_2984);
nor UO_444 (O_444,N_2993,N_2992);
and UO_445 (O_445,N_2948,N_2958);
nor UO_446 (O_446,N_2957,N_2964);
nand UO_447 (O_447,N_2946,N_2945);
nor UO_448 (O_448,N_2984,N_2963);
nor UO_449 (O_449,N_2997,N_2977);
or UO_450 (O_450,N_2992,N_2952);
and UO_451 (O_451,N_2994,N_2957);
nand UO_452 (O_452,N_2961,N_2973);
nand UO_453 (O_453,N_2943,N_2966);
or UO_454 (O_454,N_2975,N_2960);
or UO_455 (O_455,N_2943,N_2957);
and UO_456 (O_456,N_2987,N_2944);
and UO_457 (O_457,N_2991,N_2940);
nand UO_458 (O_458,N_2951,N_2987);
and UO_459 (O_459,N_2952,N_2944);
nor UO_460 (O_460,N_2995,N_2985);
nor UO_461 (O_461,N_2974,N_2957);
nor UO_462 (O_462,N_2989,N_2940);
xor UO_463 (O_463,N_2955,N_2983);
nor UO_464 (O_464,N_2954,N_2970);
nor UO_465 (O_465,N_2945,N_2973);
or UO_466 (O_466,N_2997,N_2992);
and UO_467 (O_467,N_2995,N_2990);
xor UO_468 (O_468,N_2946,N_2993);
or UO_469 (O_469,N_2946,N_2975);
nor UO_470 (O_470,N_2978,N_2940);
nand UO_471 (O_471,N_2954,N_2958);
and UO_472 (O_472,N_2948,N_2955);
or UO_473 (O_473,N_2979,N_2984);
or UO_474 (O_474,N_2996,N_2985);
or UO_475 (O_475,N_2943,N_2961);
nand UO_476 (O_476,N_2979,N_2971);
or UO_477 (O_477,N_2949,N_2948);
nand UO_478 (O_478,N_2949,N_2978);
nand UO_479 (O_479,N_2984,N_2995);
and UO_480 (O_480,N_2958,N_2951);
nand UO_481 (O_481,N_2992,N_2942);
or UO_482 (O_482,N_2968,N_2953);
and UO_483 (O_483,N_2955,N_2980);
nor UO_484 (O_484,N_2976,N_2990);
nor UO_485 (O_485,N_2954,N_2992);
nand UO_486 (O_486,N_2959,N_2994);
and UO_487 (O_487,N_2976,N_2954);
or UO_488 (O_488,N_2986,N_2984);
or UO_489 (O_489,N_2986,N_2997);
or UO_490 (O_490,N_2954,N_2993);
or UO_491 (O_491,N_2960,N_2946);
and UO_492 (O_492,N_2983,N_2959);
or UO_493 (O_493,N_2989,N_2982);
and UO_494 (O_494,N_2964,N_2944);
nor UO_495 (O_495,N_2967,N_2958);
nor UO_496 (O_496,N_2991,N_2970);
and UO_497 (O_497,N_2989,N_2952);
or UO_498 (O_498,N_2943,N_2977);
or UO_499 (O_499,N_2946,N_2957);
endmodule