module basic_750_5000_1000_5_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_422,In_172);
and U1 (N_1,In_290,In_102);
or U2 (N_2,In_433,In_379);
or U3 (N_3,In_157,In_126);
nand U4 (N_4,In_579,In_3);
nand U5 (N_5,In_735,In_174);
nor U6 (N_6,In_437,In_43);
and U7 (N_7,In_501,In_668);
or U8 (N_8,In_477,In_658);
nor U9 (N_9,In_245,In_539);
nand U10 (N_10,In_99,In_572);
nand U11 (N_11,In_693,In_651);
nand U12 (N_12,In_404,In_124);
nand U13 (N_13,In_255,In_131);
or U14 (N_14,In_642,In_465);
nand U15 (N_15,In_81,In_385);
or U16 (N_16,In_732,In_231);
nor U17 (N_17,In_349,In_53);
or U18 (N_18,In_204,In_450);
nand U19 (N_19,In_426,In_652);
or U20 (N_20,In_229,In_549);
xor U21 (N_21,In_462,In_238);
nand U22 (N_22,In_105,In_740);
or U23 (N_23,In_344,In_483);
nand U24 (N_24,In_32,In_27);
or U25 (N_25,In_224,In_354);
and U26 (N_26,In_101,In_506);
and U27 (N_27,In_108,In_79);
or U28 (N_28,In_47,In_235);
or U29 (N_29,In_681,In_534);
and U30 (N_30,In_570,In_4);
nor U31 (N_31,In_340,In_375);
or U32 (N_32,In_689,In_94);
nand U33 (N_33,In_314,In_615);
nand U34 (N_34,In_60,In_466);
nor U35 (N_35,In_300,In_160);
nand U36 (N_36,In_507,In_592);
nor U37 (N_37,In_22,In_562);
nand U38 (N_38,In_621,In_36);
or U39 (N_39,In_352,In_220);
and U40 (N_40,In_631,In_109);
xnor U41 (N_41,In_360,In_414);
xnor U42 (N_42,In_666,In_302);
nand U43 (N_43,In_278,In_331);
nor U44 (N_44,In_698,In_253);
nor U45 (N_45,In_739,In_704);
or U46 (N_46,In_103,In_384);
xor U47 (N_47,In_313,In_107);
nor U48 (N_48,In_590,In_116);
nor U49 (N_49,In_319,In_1);
or U50 (N_50,In_521,In_685);
and U51 (N_51,In_438,In_341);
and U52 (N_52,In_153,In_481);
xnor U53 (N_53,In_70,In_708);
nor U54 (N_54,In_95,In_398);
nand U55 (N_55,In_156,In_96);
or U56 (N_56,In_82,In_171);
or U57 (N_57,In_389,In_476);
nor U58 (N_58,In_610,In_209);
nor U59 (N_59,In_117,In_98);
and U60 (N_60,In_473,In_214);
and U61 (N_61,In_396,In_88);
nand U62 (N_62,In_237,In_273);
nand U63 (N_63,In_46,In_202);
nand U64 (N_64,In_597,In_288);
nand U65 (N_65,In_59,In_742);
and U66 (N_66,In_67,In_97);
or U67 (N_67,In_407,In_147);
nor U68 (N_68,In_111,In_203);
or U69 (N_69,In_645,In_627);
and U70 (N_70,In_464,In_65);
and U71 (N_71,In_439,In_18);
nor U72 (N_72,In_513,In_297);
nand U73 (N_73,In_251,In_206);
or U74 (N_74,In_193,In_62);
or U75 (N_75,In_701,In_596);
and U76 (N_76,In_670,In_730);
and U77 (N_77,In_77,In_716);
or U78 (N_78,In_338,In_227);
nand U79 (N_79,In_57,In_151);
nor U80 (N_80,In_452,In_646);
nor U81 (N_81,In_166,In_680);
nand U82 (N_82,In_6,In_244);
nand U83 (N_83,In_498,In_257);
nand U84 (N_84,In_21,In_205);
and U85 (N_85,In_733,In_576);
nand U86 (N_86,In_91,In_189);
and U87 (N_87,In_170,In_669);
or U88 (N_88,In_408,In_165);
and U89 (N_89,In_537,In_75);
or U90 (N_90,In_359,In_134);
nand U91 (N_91,In_383,In_418);
nand U92 (N_92,In_671,In_120);
nor U93 (N_93,In_162,In_720);
nor U94 (N_94,In_362,In_239);
or U95 (N_95,In_523,In_431);
nand U96 (N_96,In_444,In_9);
or U97 (N_97,In_474,In_516);
or U98 (N_98,In_311,In_718);
nor U99 (N_99,In_115,In_210);
nor U100 (N_100,In_458,In_421);
and U101 (N_101,In_486,In_327);
nor U102 (N_102,In_84,In_640);
nand U103 (N_103,In_342,In_633);
nor U104 (N_104,In_577,In_353);
nor U105 (N_105,In_243,In_390);
and U106 (N_106,In_133,In_571);
or U107 (N_107,In_695,In_283);
or U108 (N_108,In_535,In_451);
or U109 (N_109,In_130,In_86);
and U110 (N_110,In_434,In_589);
nand U111 (N_111,In_137,In_305);
or U112 (N_112,In_482,In_491);
nor U113 (N_113,In_639,In_104);
nand U114 (N_114,In_736,In_54);
and U115 (N_115,In_583,In_217);
nand U116 (N_116,In_580,In_158);
or U117 (N_117,In_643,In_55);
nor U118 (N_118,In_199,In_0);
nor U119 (N_119,In_527,In_405);
or U120 (N_120,In_492,In_269);
nor U121 (N_121,In_365,In_138);
nand U122 (N_122,In_194,In_264);
and U123 (N_123,In_173,In_40);
nand U124 (N_124,In_212,In_457);
and U125 (N_125,In_417,In_598);
and U126 (N_126,In_445,In_167);
and U127 (N_127,In_427,In_508);
or U128 (N_128,In_435,In_606);
nand U129 (N_129,In_68,In_386);
nand U130 (N_130,In_624,In_320);
nor U131 (N_131,In_358,In_279);
nor U132 (N_132,In_554,In_249);
nand U133 (N_133,In_71,In_587);
xnor U134 (N_134,In_650,In_347);
nor U135 (N_135,In_61,In_625);
nor U136 (N_136,In_87,In_282);
nor U137 (N_137,In_677,In_602);
and U138 (N_138,In_242,In_246);
nand U139 (N_139,In_16,In_455);
or U140 (N_140,In_142,In_567);
nor U141 (N_141,In_569,In_560);
and U142 (N_142,In_629,In_588);
nor U143 (N_143,In_73,In_628);
nor U144 (N_144,In_123,In_276);
and U145 (N_145,In_190,In_712);
or U146 (N_146,In_289,In_322);
and U147 (N_147,In_38,In_714);
nor U148 (N_148,In_299,In_315);
or U149 (N_149,In_684,In_710);
or U150 (N_150,In_179,In_494);
or U151 (N_151,In_582,In_8);
and U152 (N_152,In_164,In_292);
or U153 (N_153,In_132,In_89);
nor U154 (N_154,In_328,In_505);
nor U155 (N_155,In_711,In_731);
nand U156 (N_156,In_688,In_28);
nand U157 (N_157,In_557,In_661);
nor U158 (N_158,In_653,In_182);
or U159 (N_159,In_298,In_281);
and U160 (N_160,In_175,In_143);
or U161 (N_161,In_19,In_410);
and U162 (N_162,In_372,In_25);
nand U163 (N_163,In_419,In_613);
nand U164 (N_164,In_412,In_183);
and U165 (N_165,In_530,In_746);
or U166 (N_166,In_363,In_34);
or U167 (N_167,In_659,In_564);
nor U168 (N_168,In_361,In_401);
or U169 (N_169,In_400,In_188);
nor U170 (N_170,In_672,In_442);
or U171 (N_171,In_250,In_163);
or U172 (N_172,In_641,In_339);
and U173 (N_173,In_207,In_424);
and U174 (N_174,In_656,In_346);
or U175 (N_175,In_301,In_180);
or U176 (N_176,In_218,In_308);
or U177 (N_177,In_208,In_44);
nand U178 (N_178,In_168,In_692);
or U179 (N_179,In_186,In_334);
and U180 (N_180,In_11,In_608);
nand U181 (N_181,In_399,In_291);
xor U182 (N_182,In_128,In_420);
and U183 (N_183,In_321,In_377);
and U184 (N_184,In_729,In_460);
and U185 (N_185,In_552,In_617);
or U186 (N_186,In_546,In_490);
xor U187 (N_187,In_665,In_200);
or U188 (N_188,In_488,In_187);
nor U189 (N_189,In_35,In_423);
nand U190 (N_190,In_317,In_578);
nor U191 (N_191,In_333,In_493);
nand U192 (N_192,In_724,In_630);
or U193 (N_193,In_24,In_284);
nand U194 (N_194,In_125,In_679);
and U195 (N_195,In_634,In_268);
nor U196 (N_196,In_441,In_240);
and U197 (N_197,In_357,In_607);
nor U198 (N_198,In_7,In_332);
and U199 (N_199,In_366,In_667);
nor U200 (N_200,In_487,In_80);
and U201 (N_201,In_184,In_324);
nand U202 (N_202,In_416,In_141);
nand U203 (N_203,In_428,In_721);
nor U204 (N_204,In_306,In_371);
nor U205 (N_205,In_48,In_392);
nor U206 (N_206,In_161,In_382);
nand U207 (N_207,In_26,In_635);
nor U208 (N_208,In_17,In_715);
or U209 (N_209,In_644,In_647);
nor U210 (N_210,In_31,In_265);
nor U211 (N_211,In_277,In_745);
or U212 (N_212,In_50,In_456);
nand U213 (N_213,In_565,In_556);
nor U214 (N_214,In_198,In_544);
and U215 (N_215,In_674,In_686);
nand U216 (N_216,In_325,In_63);
nand U217 (N_217,In_127,In_449);
nor U218 (N_218,In_49,In_660);
nor U219 (N_219,In_430,In_550);
nand U220 (N_220,In_485,In_526);
nor U221 (N_221,In_336,In_316);
and U222 (N_222,In_118,In_155);
nand U223 (N_223,In_178,In_515);
and U224 (N_224,In_326,In_738);
nand U225 (N_225,In_558,In_702);
and U226 (N_226,In_397,In_72);
and U227 (N_227,In_555,In_259);
nor U228 (N_228,In_470,In_727);
and U229 (N_229,In_636,In_350);
nor U230 (N_230,In_663,In_637);
nand U231 (N_231,In_113,In_591);
or U232 (N_232,In_743,In_222);
nor U233 (N_233,In_216,In_586);
or U234 (N_234,In_471,In_673);
nand U235 (N_235,In_185,In_30);
or U236 (N_236,In_223,In_37);
and U237 (N_237,In_159,In_748);
or U238 (N_238,In_446,In_532);
and U239 (N_239,In_709,In_304);
or U240 (N_240,In_453,In_318);
and U241 (N_241,In_287,In_266);
and U242 (N_242,In_543,In_149);
or U243 (N_243,In_600,In_723);
nor U244 (N_244,In_52,In_459);
or U245 (N_245,In_626,In_373);
nand U246 (N_246,In_42,In_226);
or U247 (N_247,In_603,In_563);
or U248 (N_248,In_440,In_254);
nor U249 (N_249,In_335,In_475);
or U250 (N_250,In_280,In_376);
or U251 (N_251,In_533,In_119);
or U252 (N_252,In_682,In_585);
nor U253 (N_253,In_737,In_703);
nand U254 (N_254,In_380,In_241);
nor U255 (N_255,In_312,In_525);
or U256 (N_256,In_728,In_690);
nand U257 (N_257,In_262,In_225);
nand U258 (N_258,In_387,In_584);
or U259 (N_259,In_228,In_285);
or U260 (N_260,In_461,In_469);
and U261 (N_261,In_691,In_236);
or U262 (N_262,In_551,In_675);
nand U263 (N_263,In_2,In_56);
nand U264 (N_264,In_413,In_368);
nand U265 (N_265,In_337,In_725);
nand U266 (N_266,In_303,In_76);
or U267 (N_267,In_700,In_744);
and U268 (N_268,In_345,In_15);
nor U269 (N_269,In_609,In_348);
nand U270 (N_270,In_512,In_139);
nor U271 (N_271,In_29,In_545);
and U272 (N_272,In_74,In_694);
and U273 (N_273,In_484,In_406);
and U274 (N_274,In_140,In_500);
or U275 (N_275,In_374,In_136);
or U276 (N_276,In_741,In_370);
nand U277 (N_277,In_529,In_114);
nand U278 (N_278,In_619,In_504);
or U279 (N_279,In_270,In_286);
nor U280 (N_280,In_568,In_467);
and U281 (N_281,In_355,In_649);
nor U282 (N_282,In_497,In_622);
or U283 (N_283,In_154,In_541);
xnor U284 (N_284,In_395,In_201);
nor U285 (N_285,In_454,In_260);
nand U286 (N_286,In_699,In_272);
nand U287 (N_287,In_601,In_391);
nand U288 (N_288,In_330,In_192);
or U289 (N_289,In_267,In_581);
nand U290 (N_290,In_135,In_294);
nor U291 (N_291,In_425,In_664);
xor U292 (N_292,In_12,In_92);
or U293 (N_293,In_14,In_388);
or U294 (N_294,In_181,In_623);
and U295 (N_295,In_51,In_263);
or U296 (N_296,In_542,In_705);
and U297 (N_297,In_478,In_517);
or U298 (N_298,In_66,In_655);
nor U299 (N_299,In_632,In_215);
nand U300 (N_300,In_706,In_747);
nand U301 (N_301,In_69,In_247);
or U302 (N_302,In_150,In_232);
or U303 (N_303,In_447,In_531);
nor U304 (N_304,In_573,In_749);
and U305 (N_305,In_575,In_502);
nand U306 (N_306,In_146,In_112);
xnor U307 (N_307,In_85,In_654);
nor U308 (N_308,In_595,In_605);
and U309 (N_309,In_520,In_616);
nand U310 (N_310,In_381,In_233);
and U311 (N_311,In_122,In_378);
nand U312 (N_312,In_536,In_599);
nor U313 (N_313,In_436,In_191);
nand U314 (N_314,In_93,In_169);
nand U315 (N_315,In_618,In_274);
or U316 (N_316,In_518,In_310);
and U317 (N_317,In_489,In_296);
nand U318 (N_318,In_503,In_211);
xor U319 (N_319,In_468,In_528);
nand U320 (N_320,In_295,In_230);
and U321 (N_321,In_394,In_271);
nand U322 (N_322,In_83,In_100);
nor U323 (N_323,In_261,In_221);
or U324 (N_324,In_522,In_719);
or U325 (N_325,In_726,In_20);
and U326 (N_326,In_356,In_196);
nor U327 (N_327,In_519,In_176);
nor U328 (N_328,In_495,In_393);
or U329 (N_329,In_121,In_566);
nand U330 (N_330,In_678,In_574);
or U331 (N_331,In_33,In_480);
nand U332 (N_332,In_687,In_559);
nand U333 (N_333,In_248,In_547);
and U334 (N_334,In_538,In_45);
or U335 (N_335,In_323,In_5);
nor U336 (N_336,In_329,In_614);
or U337 (N_337,In_479,In_432);
or U338 (N_338,In_90,In_499);
or U339 (N_339,In_364,In_197);
and U340 (N_340,In_145,In_604);
or U341 (N_341,In_152,In_129);
or U342 (N_342,In_612,In_676);
nor U343 (N_343,In_148,In_429);
nand U344 (N_344,In_415,In_593);
and U345 (N_345,In_548,In_293);
nand U346 (N_346,In_402,In_662);
xor U347 (N_347,In_511,In_177);
nand U348 (N_348,In_722,In_697);
and U349 (N_349,In_106,In_275);
or U350 (N_350,In_734,In_369);
or U351 (N_351,In_496,In_41);
or U352 (N_352,In_472,In_463);
and U353 (N_353,In_713,In_252);
nand U354 (N_354,In_648,In_448);
nand U355 (N_355,In_343,In_717);
and U356 (N_356,In_696,In_256);
and U357 (N_357,In_553,In_144);
nand U358 (N_358,In_219,In_443);
nor U359 (N_359,In_23,In_509);
nor U360 (N_360,In_514,In_367);
nor U361 (N_361,In_638,In_110);
or U362 (N_362,In_258,In_594);
nand U363 (N_363,In_213,In_13);
nand U364 (N_364,In_39,In_78);
or U365 (N_365,In_657,In_234);
or U366 (N_366,In_195,In_540);
nand U367 (N_367,In_58,In_409);
xor U368 (N_368,In_64,In_683);
nor U369 (N_369,In_309,In_403);
nor U370 (N_370,In_524,In_411);
and U371 (N_371,In_10,In_351);
nor U372 (N_372,In_707,In_620);
and U373 (N_373,In_307,In_510);
nand U374 (N_374,In_561,In_611);
or U375 (N_375,In_359,In_576);
or U376 (N_376,In_691,In_207);
nor U377 (N_377,In_619,In_386);
nand U378 (N_378,In_471,In_457);
and U379 (N_379,In_442,In_713);
nand U380 (N_380,In_97,In_170);
or U381 (N_381,In_615,In_607);
nand U382 (N_382,In_356,In_143);
or U383 (N_383,In_527,In_623);
nor U384 (N_384,In_480,In_550);
or U385 (N_385,In_349,In_710);
nor U386 (N_386,In_303,In_653);
or U387 (N_387,In_237,In_291);
nor U388 (N_388,In_370,In_435);
or U389 (N_389,In_480,In_504);
or U390 (N_390,In_318,In_71);
nor U391 (N_391,In_634,In_354);
nand U392 (N_392,In_193,In_609);
nand U393 (N_393,In_80,In_519);
and U394 (N_394,In_145,In_50);
or U395 (N_395,In_428,In_675);
nor U396 (N_396,In_169,In_741);
nor U397 (N_397,In_549,In_606);
nand U398 (N_398,In_237,In_349);
or U399 (N_399,In_160,In_452);
and U400 (N_400,In_52,In_44);
nor U401 (N_401,In_344,In_185);
nor U402 (N_402,In_306,In_41);
or U403 (N_403,In_450,In_735);
and U404 (N_404,In_201,In_130);
and U405 (N_405,In_606,In_188);
nor U406 (N_406,In_339,In_428);
and U407 (N_407,In_43,In_569);
or U408 (N_408,In_602,In_299);
nor U409 (N_409,In_156,In_357);
nand U410 (N_410,In_233,In_595);
or U411 (N_411,In_374,In_362);
nand U412 (N_412,In_649,In_345);
and U413 (N_413,In_666,In_288);
or U414 (N_414,In_128,In_501);
or U415 (N_415,In_111,In_698);
and U416 (N_416,In_627,In_617);
and U417 (N_417,In_155,In_703);
nand U418 (N_418,In_442,In_539);
or U419 (N_419,In_477,In_730);
nor U420 (N_420,In_549,In_512);
or U421 (N_421,In_551,In_278);
or U422 (N_422,In_371,In_428);
and U423 (N_423,In_289,In_245);
and U424 (N_424,In_451,In_403);
nand U425 (N_425,In_142,In_719);
or U426 (N_426,In_630,In_292);
and U427 (N_427,In_10,In_576);
and U428 (N_428,In_556,In_153);
nand U429 (N_429,In_247,In_130);
nor U430 (N_430,In_485,In_498);
and U431 (N_431,In_518,In_611);
nand U432 (N_432,In_698,In_137);
nor U433 (N_433,In_213,In_168);
nor U434 (N_434,In_171,In_51);
or U435 (N_435,In_175,In_478);
and U436 (N_436,In_305,In_224);
and U437 (N_437,In_570,In_444);
or U438 (N_438,In_264,In_221);
nor U439 (N_439,In_563,In_73);
nor U440 (N_440,In_236,In_92);
or U441 (N_441,In_130,In_602);
xor U442 (N_442,In_263,In_121);
or U443 (N_443,In_677,In_700);
or U444 (N_444,In_500,In_637);
or U445 (N_445,In_502,In_468);
and U446 (N_446,In_537,In_433);
nand U447 (N_447,In_479,In_476);
nor U448 (N_448,In_599,In_143);
nand U449 (N_449,In_108,In_713);
nor U450 (N_450,In_445,In_530);
and U451 (N_451,In_229,In_231);
and U452 (N_452,In_188,In_573);
and U453 (N_453,In_251,In_416);
nor U454 (N_454,In_200,In_194);
nand U455 (N_455,In_448,In_676);
nor U456 (N_456,In_626,In_594);
and U457 (N_457,In_226,In_582);
or U458 (N_458,In_660,In_340);
and U459 (N_459,In_392,In_600);
or U460 (N_460,In_445,In_335);
and U461 (N_461,In_182,In_209);
and U462 (N_462,In_146,In_551);
nand U463 (N_463,In_739,In_213);
or U464 (N_464,In_568,In_77);
and U465 (N_465,In_450,In_749);
and U466 (N_466,In_407,In_91);
xor U467 (N_467,In_127,In_426);
nor U468 (N_468,In_728,In_672);
nor U469 (N_469,In_391,In_84);
xor U470 (N_470,In_265,In_274);
or U471 (N_471,In_592,In_438);
or U472 (N_472,In_601,In_269);
nor U473 (N_473,In_35,In_725);
and U474 (N_474,In_560,In_391);
nor U475 (N_475,In_283,In_287);
nand U476 (N_476,In_233,In_131);
or U477 (N_477,In_585,In_691);
and U478 (N_478,In_103,In_390);
nor U479 (N_479,In_744,In_333);
nor U480 (N_480,In_168,In_719);
nor U481 (N_481,In_583,In_551);
nor U482 (N_482,In_619,In_524);
and U483 (N_483,In_368,In_590);
nand U484 (N_484,In_283,In_452);
nor U485 (N_485,In_241,In_331);
nor U486 (N_486,In_683,In_53);
and U487 (N_487,In_561,In_643);
and U488 (N_488,In_240,In_436);
xor U489 (N_489,In_688,In_452);
and U490 (N_490,In_516,In_289);
nor U491 (N_491,In_454,In_74);
and U492 (N_492,In_248,In_262);
and U493 (N_493,In_130,In_617);
or U494 (N_494,In_387,In_696);
nand U495 (N_495,In_452,In_417);
and U496 (N_496,In_61,In_297);
nand U497 (N_497,In_392,In_39);
or U498 (N_498,In_243,In_512);
and U499 (N_499,In_496,In_374);
nand U500 (N_500,In_391,In_273);
nand U501 (N_501,In_122,In_738);
or U502 (N_502,In_116,In_438);
and U503 (N_503,In_205,In_424);
and U504 (N_504,In_269,In_262);
or U505 (N_505,In_721,In_622);
or U506 (N_506,In_116,In_466);
nor U507 (N_507,In_481,In_435);
nand U508 (N_508,In_679,In_138);
and U509 (N_509,In_434,In_451);
nor U510 (N_510,In_290,In_275);
xnor U511 (N_511,In_1,In_126);
nor U512 (N_512,In_186,In_120);
or U513 (N_513,In_506,In_234);
or U514 (N_514,In_536,In_343);
nand U515 (N_515,In_674,In_37);
nor U516 (N_516,In_30,In_162);
and U517 (N_517,In_361,In_235);
nand U518 (N_518,In_260,In_145);
nor U519 (N_519,In_595,In_564);
xor U520 (N_520,In_673,In_703);
and U521 (N_521,In_300,In_459);
and U522 (N_522,In_37,In_370);
or U523 (N_523,In_194,In_86);
nor U524 (N_524,In_36,In_38);
or U525 (N_525,In_481,In_453);
and U526 (N_526,In_106,In_46);
or U527 (N_527,In_527,In_274);
and U528 (N_528,In_543,In_70);
or U529 (N_529,In_6,In_222);
nor U530 (N_530,In_83,In_553);
nor U531 (N_531,In_247,In_596);
nor U532 (N_532,In_249,In_318);
or U533 (N_533,In_288,In_533);
nand U534 (N_534,In_714,In_138);
or U535 (N_535,In_598,In_332);
and U536 (N_536,In_494,In_669);
or U537 (N_537,In_0,In_308);
xor U538 (N_538,In_156,In_534);
nand U539 (N_539,In_621,In_131);
and U540 (N_540,In_255,In_607);
or U541 (N_541,In_387,In_410);
nand U542 (N_542,In_561,In_498);
and U543 (N_543,In_190,In_154);
and U544 (N_544,In_85,In_524);
nor U545 (N_545,In_601,In_332);
and U546 (N_546,In_23,In_149);
nor U547 (N_547,In_538,In_415);
and U548 (N_548,In_519,In_81);
xnor U549 (N_549,In_515,In_230);
nor U550 (N_550,In_564,In_334);
xnor U551 (N_551,In_308,In_42);
and U552 (N_552,In_368,In_602);
or U553 (N_553,In_43,In_400);
and U554 (N_554,In_335,In_258);
and U555 (N_555,In_41,In_45);
or U556 (N_556,In_329,In_361);
or U557 (N_557,In_363,In_672);
and U558 (N_558,In_237,In_531);
and U559 (N_559,In_705,In_336);
nor U560 (N_560,In_473,In_749);
nor U561 (N_561,In_297,In_342);
nor U562 (N_562,In_721,In_339);
and U563 (N_563,In_570,In_209);
or U564 (N_564,In_548,In_483);
or U565 (N_565,In_402,In_412);
nand U566 (N_566,In_613,In_324);
nand U567 (N_567,In_164,In_746);
nor U568 (N_568,In_487,In_48);
xnor U569 (N_569,In_301,In_234);
and U570 (N_570,In_527,In_159);
xor U571 (N_571,In_524,In_726);
and U572 (N_572,In_3,In_721);
or U573 (N_573,In_524,In_339);
or U574 (N_574,In_142,In_580);
nand U575 (N_575,In_386,In_106);
nand U576 (N_576,In_561,In_279);
nor U577 (N_577,In_271,In_222);
nor U578 (N_578,In_501,In_172);
and U579 (N_579,In_26,In_325);
or U580 (N_580,In_66,In_283);
and U581 (N_581,In_611,In_33);
nand U582 (N_582,In_593,In_651);
and U583 (N_583,In_730,In_297);
nand U584 (N_584,In_551,In_405);
or U585 (N_585,In_184,In_216);
and U586 (N_586,In_334,In_147);
nand U587 (N_587,In_92,In_552);
or U588 (N_588,In_587,In_556);
nand U589 (N_589,In_535,In_688);
nor U590 (N_590,In_50,In_546);
or U591 (N_591,In_171,In_266);
and U592 (N_592,In_394,In_211);
and U593 (N_593,In_624,In_673);
or U594 (N_594,In_9,In_257);
nand U595 (N_595,In_32,In_30);
and U596 (N_596,In_498,In_18);
nand U597 (N_597,In_740,In_87);
or U598 (N_598,In_716,In_374);
and U599 (N_599,In_587,In_451);
nor U600 (N_600,In_688,In_113);
and U601 (N_601,In_582,In_707);
or U602 (N_602,In_423,In_473);
nor U603 (N_603,In_51,In_177);
or U604 (N_604,In_78,In_504);
and U605 (N_605,In_161,In_176);
and U606 (N_606,In_323,In_482);
and U607 (N_607,In_583,In_113);
nor U608 (N_608,In_5,In_503);
nor U609 (N_609,In_241,In_313);
or U610 (N_610,In_453,In_571);
nor U611 (N_611,In_572,In_657);
nor U612 (N_612,In_540,In_495);
nand U613 (N_613,In_532,In_519);
or U614 (N_614,In_481,In_286);
or U615 (N_615,In_463,In_642);
or U616 (N_616,In_28,In_301);
nor U617 (N_617,In_731,In_603);
nand U618 (N_618,In_200,In_34);
nor U619 (N_619,In_75,In_598);
nand U620 (N_620,In_255,In_478);
nand U621 (N_621,In_147,In_144);
or U622 (N_622,In_168,In_536);
nor U623 (N_623,In_86,In_565);
xor U624 (N_624,In_669,In_64);
or U625 (N_625,In_210,In_5);
or U626 (N_626,In_62,In_536);
and U627 (N_627,In_330,In_293);
or U628 (N_628,In_641,In_620);
nand U629 (N_629,In_357,In_495);
nand U630 (N_630,In_318,In_572);
and U631 (N_631,In_579,In_262);
nand U632 (N_632,In_718,In_18);
nor U633 (N_633,In_699,In_664);
or U634 (N_634,In_522,In_107);
or U635 (N_635,In_369,In_103);
nor U636 (N_636,In_170,In_67);
nor U637 (N_637,In_354,In_727);
nor U638 (N_638,In_2,In_134);
and U639 (N_639,In_148,In_449);
nand U640 (N_640,In_329,In_198);
nor U641 (N_641,In_460,In_557);
and U642 (N_642,In_499,In_183);
or U643 (N_643,In_636,In_310);
nand U644 (N_644,In_108,In_268);
or U645 (N_645,In_550,In_142);
or U646 (N_646,In_94,In_413);
and U647 (N_647,In_480,In_108);
or U648 (N_648,In_485,In_47);
and U649 (N_649,In_30,In_24);
nor U650 (N_650,In_358,In_424);
nor U651 (N_651,In_355,In_448);
and U652 (N_652,In_614,In_657);
or U653 (N_653,In_505,In_108);
and U654 (N_654,In_727,In_521);
nand U655 (N_655,In_676,In_334);
nor U656 (N_656,In_718,In_23);
or U657 (N_657,In_318,In_725);
nand U658 (N_658,In_380,In_127);
and U659 (N_659,In_702,In_163);
and U660 (N_660,In_224,In_309);
nand U661 (N_661,In_504,In_571);
and U662 (N_662,In_37,In_628);
nand U663 (N_663,In_413,In_75);
nor U664 (N_664,In_283,In_456);
or U665 (N_665,In_149,In_20);
nor U666 (N_666,In_653,In_621);
nor U667 (N_667,In_245,In_389);
nand U668 (N_668,In_209,In_534);
nor U669 (N_669,In_635,In_129);
nor U670 (N_670,In_362,In_553);
nor U671 (N_671,In_93,In_431);
nor U672 (N_672,In_210,In_22);
or U673 (N_673,In_621,In_65);
or U674 (N_674,In_119,In_46);
nor U675 (N_675,In_451,In_581);
nor U676 (N_676,In_181,In_226);
and U677 (N_677,In_43,In_647);
nand U678 (N_678,In_374,In_254);
and U679 (N_679,In_240,In_318);
nor U680 (N_680,In_270,In_511);
nor U681 (N_681,In_546,In_579);
nor U682 (N_682,In_659,In_437);
nand U683 (N_683,In_575,In_527);
nand U684 (N_684,In_73,In_65);
nand U685 (N_685,In_464,In_204);
nand U686 (N_686,In_86,In_282);
or U687 (N_687,In_528,In_565);
and U688 (N_688,In_723,In_320);
nand U689 (N_689,In_350,In_382);
and U690 (N_690,In_85,In_142);
and U691 (N_691,In_550,In_472);
or U692 (N_692,In_35,In_686);
and U693 (N_693,In_204,In_445);
nand U694 (N_694,In_565,In_204);
or U695 (N_695,In_7,In_293);
nand U696 (N_696,In_264,In_663);
and U697 (N_697,In_85,In_677);
nor U698 (N_698,In_358,In_187);
xnor U699 (N_699,In_86,In_314);
nand U700 (N_700,In_408,In_217);
nor U701 (N_701,In_274,In_130);
nand U702 (N_702,In_372,In_373);
nand U703 (N_703,In_442,In_406);
and U704 (N_704,In_211,In_411);
nand U705 (N_705,In_442,In_333);
and U706 (N_706,In_506,In_6);
nand U707 (N_707,In_461,In_393);
nor U708 (N_708,In_615,In_664);
nor U709 (N_709,In_271,In_561);
or U710 (N_710,In_209,In_627);
nand U711 (N_711,In_686,In_128);
or U712 (N_712,In_119,In_49);
nand U713 (N_713,In_54,In_384);
or U714 (N_714,In_221,In_470);
or U715 (N_715,In_603,In_467);
nor U716 (N_716,In_689,In_187);
and U717 (N_717,In_408,In_249);
nand U718 (N_718,In_180,In_315);
or U719 (N_719,In_150,In_346);
nand U720 (N_720,In_550,In_542);
nand U721 (N_721,In_688,In_504);
or U722 (N_722,In_592,In_52);
and U723 (N_723,In_381,In_619);
or U724 (N_724,In_475,In_476);
and U725 (N_725,In_444,In_528);
nor U726 (N_726,In_607,In_621);
and U727 (N_727,In_321,In_513);
nand U728 (N_728,In_278,In_372);
or U729 (N_729,In_240,In_742);
nand U730 (N_730,In_278,In_162);
nand U731 (N_731,In_98,In_245);
or U732 (N_732,In_552,In_576);
nor U733 (N_733,In_582,In_122);
nor U734 (N_734,In_537,In_349);
nand U735 (N_735,In_292,In_213);
or U736 (N_736,In_127,In_222);
or U737 (N_737,In_279,In_716);
and U738 (N_738,In_141,In_630);
and U739 (N_739,In_166,In_462);
nor U740 (N_740,In_414,In_126);
nand U741 (N_741,In_148,In_293);
nand U742 (N_742,In_176,In_128);
and U743 (N_743,In_394,In_620);
nand U744 (N_744,In_666,In_615);
or U745 (N_745,In_687,In_139);
or U746 (N_746,In_481,In_75);
nand U747 (N_747,In_2,In_501);
or U748 (N_748,In_144,In_346);
xnor U749 (N_749,In_61,In_526);
xor U750 (N_750,In_274,In_673);
nor U751 (N_751,In_95,In_186);
or U752 (N_752,In_292,In_349);
xor U753 (N_753,In_54,In_446);
nor U754 (N_754,In_200,In_712);
nor U755 (N_755,In_512,In_51);
and U756 (N_756,In_748,In_654);
nor U757 (N_757,In_204,In_504);
or U758 (N_758,In_641,In_138);
and U759 (N_759,In_351,In_182);
nor U760 (N_760,In_374,In_629);
or U761 (N_761,In_345,In_383);
and U762 (N_762,In_337,In_201);
and U763 (N_763,In_90,In_228);
or U764 (N_764,In_564,In_556);
nor U765 (N_765,In_661,In_75);
nor U766 (N_766,In_439,In_92);
or U767 (N_767,In_748,In_596);
nor U768 (N_768,In_518,In_688);
or U769 (N_769,In_451,In_106);
or U770 (N_770,In_220,In_317);
nor U771 (N_771,In_499,In_472);
or U772 (N_772,In_716,In_705);
and U773 (N_773,In_672,In_336);
nor U774 (N_774,In_470,In_628);
nand U775 (N_775,In_430,In_88);
nor U776 (N_776,In_24,In_489);
and U777 (N_777,In_18,In_150);
and U778 (N_778,In_133,In_72);
and U779 (N_779,In_383,In_175);
nand U780 (N_780,In_442,In_525);
nand U781 (N_781,In_529,In_99);
nor U782 (N_782,In_712,In_727);
nor U783 (N_783,In_34,In_381);
nand U784 (N_784,In_446,In_208);
or U785 (N_785,In_489,In_451);
and U786 (N_786,In_430,In_177);
nand U787 (N_787,In_417,In_97);
and U788 (N_788,In_247,In_475);
and U789 (N_789,In_313,In_11);
and U790 (N_790,In_89,In_533);
or U791 (N_791,In_645,In_217);
nor U792 (N_792,In_650,In_420);
or U793 (N_793,In_676,In_243);
or U794 (N_794,In_1,In_712);
nor U795 (N_795,In_332,In_507);
nor U796 (N_796,In_694,In_51);
or U797 (N_797,In_732,In_515);
and U798 (N_798,In_710,In_200);
nand U799 (N_799,In_215,In_527);
nor U800 (N_800,In_629,In_293);
or U801 (N_801,In_197,In_312);
or U802 (N_802,In_599,In_123);
nor U803 (N_803,In_233,In_200);
nand U804 (N_804,In_577,In_540);
or U805 (N_805,In_306,In_203);
nand U806 (N_806,In_187,In_735);
and U807 (N_807,In_18,In_595);
nand U808 (N_808,In_84,In_141);
or U809 (N_809,In_220,In_10);
nor U810 (N_810,In_642,In_74);
and U811 (N_811,In_721,In_79);
or U812 (N_812,In_468,In_271);
and U813 (N_813,In_488,In_673);
nand U814 (N_814,In_496,In_491);
xnor U815 (N_815,In_119,In_266);
and U816 (N_816,In_129,In_58);
and U817 (N_817,In_251,In_447);
or U818 (N_818,In_204,In_393);
and U819 (N_819,In_560,In_158);
and U820 (N_820,In_389,In_254);
nand U821 (N_821,In_239,In_371);
or U822 (N_822,In_486,In_140);
or U823 (N_823,In_464,In_440);
nor U824 (N_824,In_479,In_199);
nand U825 (N_825,In_311,In_140);
or U826 (N_826,In_438,In_598);
nor U827 (N_827,In_694,In_38);
nand U828 (N_828,In_215,In_163);
or U829 (N_829,In_198,In_490);
nor U830 (N_830,In_679,In_275);
or U831 (N_831,In_656,In_245);
and U832 (N_832,In_459,In_712);
or U833 (N_833,In_413,In_81);
nor U834 (N_834,In_340,In_676);
nand U835 (N_835,In_513,In_62);
nor U836 (N_836,In_694,In_268);
nand U837 (N_837,In_499,In_608);
or U838 (N_838,In_467,In_290);
nand U839 (N_839,In_153,In_627);
and U840 (N_840,In_320,In_36);
nor U841 (N_841,In_249,In_211);
nor U842 (N_842,In_101,In_652);
nand U843 (N_843,In_675,In_302);
nor U844 (N_844,In_681,In_585);
nand U845 (N_845,In_338,In_247);
nand U846 (N_846,In_27,In_568);
and U847 (N_847,In_39,In_746);
nand U848 (N_848,In_544,In_233);
and U849 (N_849,In_327,In_584);
nor U850 (N_850,In_207,In_140);
nand U851 (N_851,In_418,In_717);
and U852 (N_852,In_491,In_113);
nor U853 (N_853,In_34,In_407);
nand U854 (N_854,In_67,In_39);
nor U855 (N_855,In_545,In_556);
nor U856 (N_856,In_672,In_595);
or U857 (N_857,In_517,In_742);
and U858 (N_858,In_582,In_670);
and U859 (N_859,In_651,In_560);
nor U860 (N_860,In_737,In_310);
or U861 (N_861,In_155,In_242);
nand U862 (N_862,In_271,In_607);
nor U863 (N_863,In_75,In_423);
and U864 (N_864,In_312,In_370);
nand U865 (N_865,In_472,In_204);
nor U866 (N_866,In_645,In_198);
or U867 (N_867,In_53,In_498);
or U868 (N_868,In_106,In_608);
and U869 (N_869,In_235,In_675);
and U870 (N_870,In_589,In_347);
and U871 (N_871,In_640,In_165);
and U872 (N_872,In_433,In_388);
nor U873 (N_873,In_26,In_604);
and U874 (N_874,In_489,In_27);
nand U875 (N_875,In_736,In_425);
nor U876 (N_876,In_127,In_335);
nand U877 (N_877,In_278,In_306);
nor U878 (N_878,In_258,In_170);
nand U879 (N_879,In_677,In_607);
or U880 (N_880,In_656,In_220);
xnor U881 (N_881,In_11,In_334);
nor U882 (N_882,In_576,In_168);
nor U883 (N_883,In_556,In_697);
nand U884 (N_884,In_654,In_649);
or U885 (N_885,In_83,In_322);
nor U886 (N_886,In_558,In_300);
nand U887 (N_887,In_661,In_398);
nor U888 (N_888,In_61,In_125);
nand U889 (N_889,In_671,In_71);
nand U890 (N_890,In_429,In_409);
and U891 (N_891,In_214,In_283);
nand U892 (N_892,In_362,In_266);
nor U893 (N_893,In_388,In_426);
and U894 (N_894,In_604,In_48);
or U895 (N_895,In_560,In_721);
xnor U896 (N_896,In_66,In_147);
and U897 (N_897,In_567,In_119);
xnor U898 (N_898,In_257,In_304);
or U899 (N_899,In_646,In_440);
or U900 (N_900,In_741,In_283);
and U901 (N_901,In_574,In_226);
nand U902 (N_902,In_62,In_521);
or U903 (N_903,In_748,In_650);
xor U904 (N_904,In_242,In_485);
xnor U905 (N_905,In_329,In_441);
and U906 (N_906,In_497,In_32);
nand U907 (N_907,In_403,In_189);
or U908 (N_908,In_199,In_308);
and U909 (N_909,In_37,In_343);
and U910 (N_910,In_656,In_178);
nor U911 (N_911,In_604,In_616);
nand U912 (N_912,In_351,In_104);
and U913 (N_913,In_462,In_59);
xor U914 (N_914,In_76,In_123);
and U915 (N_915,In_204,In_525);
and U916 (N_916,In_192,In_582);
or U917 (N_917,In_251,In_14);
nand U918 (N_918,In_57,In_633);
nor U919 (N_919,In_448,In_83);
or U920 (N_920,In_100,In_569);
and U921 (N_921,In_400,In_60);
nor U922 (N_922,In_380,In_619);
and U923 (N_923,In_229,In_667);
nand U924 (N_924,In_249,In_160);
or U925 (N_925,In_31,In_599);
or U926 (N_926,In_637,In_218);
nand U927 (N_927,In_214,In_458);
or U928 (N_928,In_196,In_310);
and U929 (N_929,In_233,In_556);
nand U930 (N_930,In_107,In_693);
or U931 (N_931,In_425,In_78);
nor U932 (N_932,In_509,In_313);
and U933 (N_933,In_388,In_76);
nor U934 (N_934,In_722,In_724);
nor U935 (N_935,In_172,In_2);
nor U936 (N_936,In_92,In_604);
and U937 (N_937,In_220,In_681);
nand U938 (N_938,In_677,In_569);
nor U939 (N_939,In_405,In_365);
nand U940 (N_940,In_260,In_135);
and U941 (N_941,In_17,In_99);
nand U942 (N_942,In_534,In_702);
xor U943 (N_943,In_568,In_240);
xor U944 (N_944,In_103,In_360);
or U945 (N_945,In_339,In_27);
nand U946 (N_946,In_211,In_243);
nor U947 (N_947,In_65,In_210);
or U948 (N_948,In_399,In_411);
and U949 (N_949,In_372,In_744);
and U950 (N_950,In_540,In_736);
nand U951 (N_951,In_701,In_290);
nor U952 (N_952,In_208,In_447);
and U953 (N_953,In_143,In_240);
nor U954 (N_954,In_532,In_684);
and U955 (N_955,In_602,In_129);
nor U956 (N_956,In_143,In_168);
or U957 (N_957,In_52,In_77);
nand U958 (N_958,In_178,In_566);
or U959 (N_959,In_57,In_587);
or U960 (N_960,In_738,In_275);
nor U961 (N_961,In_200,In_360);
and U962 (N_962,In_636,In_573);
nand U963 (N_963,In_518,In_20);
or U964 (N_964,In_634,In_558);
and U965 (N_965,In_662,In_122);
nand U966 (N_966,In_68,In_131);
or U967 (N_967,In_16,In_173);
nand U968 (N_968,In_9,In_664);
nand U969 (N_969,In_107,In_518);
or U970 (N_970,In_446,In_165);
nand U971 (N_971,In_748,In_606);
nand U972 (N_972,In_437,In_475);
nand U973 (N_973,In_8,In_550);
or U974 (N_974,In_524,In_468);
or U975 (N_975,In_235,In_584);
nand U976 (N_976,In_196,In_76);
nand U977 (N_977,In_220,In_192);
nand U978 (N_978,In_491,In_648);
and U979 (N_979,In_373,In_652);
or U980 (N_980,In_695,In_39);
or U981 (N_981,In_28,In_572);
or U982 (N_982,In_544,In_206);
nand U983 (N_983,In_10,In_99);
or U984 (N_984,In_707,In_1);
nor U985 (N_985,In_74,In_545);
or U986 (N_986,In_156,In_474);
nand U987 (N_987,In_468,In_663);
or U988 (N_988,In_278,In_327);
nor U989 (N_989,In_437,In_120);
or U990 (N_990,In_728,In_543);
or U991 (N_991,In_570,In_309);
and U992 (N_992,In_140,In_627);
or U993 (N_993,In_49,In_30);
nand U994 (N_994,In_174,In_567);
nor U995 (N_995,In_41,In_77);
and U996 (N_996,In_6,In_276);
or U997 (N_997,In_19,In_233);
nor U998 (N_998,In_716,In_682);
and U999 (N_999,In_98,In_376);
nor U1000 (N_1000,N_44,N_980);
nor U1001 (N_1001,N_342,N_678);
and U1002 (N_1002,N_744,N_358);
xnor U1003 (N_1003,N_430,N_765);
or U1004 (N_1004,N_248,N_572);
nand U1005 (N_1005,N_715,N_783);
nand U1006 (N_1006,N_348,N_285);
and U1007 (N_1007,N_302,N_823);
nand U1008 (N_1008,N_707,N_402);
or U1009 (N_1009,N_301,N_237);
or U1010 (N_1010,N_870,N_610);
or U1011 (N_1011,N_995,N_568);
and U1012 (N_1012,N_520,N_991);
nand U1013 (N_1013,N_68,N_484);
nor U1014 (N_1014,N_762,N_627);
and U1015 (N_1015,N_562,N_999);
nor U1016 (N_1016,N_984,N_888);
or U1017 (N_1017,N_440,N_851);
and U1018 (N_1018,N_625,N_261);
and U1019 (N_1019,N_278,N_263);
or U1020 (N_1020,N_56,N_608);
and U1021 (N_1021,N_48,N_753);
and U1022 (N_1022,N_719,N_446);
or U1023 (N_1023,N_398,N_357);
or U1024 (N_1024,N_677,N_617);
and U1025 (N_1025,N_156,N_733);
xor U1026 (N_1026,N_722,N_815);
nand U1027 (N_1027,N_909,N_307);
and U1028 (N_1028,N_181,N_209);
and U1029 (N_1029,N_464,N_308);
or U1030 (N_1030,N_57,N_604);
or U1031 (N_1031,N_162,N_8);
and U1032 (N_1032,N_894,N_576);
or U1033 (N_1033,N_49,N_921);
nand U1034 (N_1034,N_145,N_16);
and U1035 (N_1035,N_498,N_53);
nand U1036 (N_1036,N_350,N_517);
nand U1037 (N_1037,N_812,N_317);
nor U1038 (N_1038,N_778,N_923);
xor U1039 (N_1039,N_613,N_516);
and U1040 (N_1040,N_533,N_55);
or U1041 (N_1041,N_717,N_501);
nand U1042 (N_1042,N_405,N_238);
or U1043 (N_1043,N_745,N_876);
nand U1044 (N_1044,N_890,N_391);
nor U1045 (N_1045,N_584,N_935);
nor U1046 (N_1046,N_942,N_293);
and U1047 (N_1047,N_754,N_699);
and U1048 (N_1048,N_396,N_370);
and U1049 (N_1049,N_99,N_144);
or U1050 (N_1050,N_970,N_967);
or U1051 (N_1051,N_413,N_406);
and U1052 (N_1052,N_938,N_544);
nand U1053 (N_1053,N_190,N_555);
nor U1054 (N_1054,N_657,N_1);
or U1055 (N_1055,N_690,N_211);
or U1056 (N_1056,N_421,N_708);
nand U1057 (N_1057,N_149,N_705);
nand U1058 (N_1058,N_356,N_19);
nand U1059 (N_1059,N_117,N_454);
xor U1060 (N_1060,N_30,N_362);
or U1061 (N_1061,N_10,N_534);
nand U1062 (N_1062,N_655,N_686);
nor U1063 (N_1063,N_667,N_259);
or U1064 (N_1064,N_133,N_879);
or U1065 (N_1065,N_643,N_456);
nor U1066 (N_1066,N_7,N_485);
or U1067 (N_1067,N_956,N_969);
and U1068 (N_1068,N_96,N_279);
nand U1069 (N_1069,N_164,N_343);
nor U1070 (N_1070,N_877,N_839);
nand U1071 (N_1071,N_423,N_266);
and U1072 (N_1072,N_588,N_509);
and U1073 (N_1073,N_561,N_735);
xor U1074 (N_1074,N_933,N_540);
and U1075 (N_1075,N_861,N_640);
or U1076 (N_1076,N_69,N_341);
nor U1077 (N_1077,N_208,N_602);
nand U1078 (N_1078,N_321,N_739);
nor U1079 (N_1079,N_43,N_168);
and U1080 (N_1080,N_650,N_135);
and U1081 (N_1081,N_775,N_869);
nand U1082 (N_1082,N_789,N_728);
or U1083 (N_1083,N_896,N_893);
nor U1084 (N_1084,N_609,N_510);
or U1085 (N_1085,N_693,N_127);
or U1086 (N_1086,N_521,N_670);
nand U1087 (N_1087,N_236,N_581);
nor U1088 (N_1088,N_74,N_811);
or U1089 (N_1089,N_930,N_571);
nand U1090 (N_1090,N_577,N_37);
nand U1091 (N_1091,N_679,N_442);
nand U1092 (N_1092,N_605,N_788);
and U1093 (N_1093,N_17,N_619);
nand U1094 (N_1094,N_11,N_558);
nor U1095 (N_1095,N_120,N_444);
or U1096 (N_1096,N_629,N_70);
and U1097 (N_1097,N_860,N_689);
nand U1098 (N_1098,N_157,N_926);
or U1099 (N_1099,N_462,N_294);
nand U1100 (N_1100,N_75,N_136);
nand U1101 (N_1101,N_375,N_784);
nor U1102 (N_1102,N_445,N_163);
nor U1103 (N_1103,N_4,N_996);
and U1104 (N_1104,N_770,N_78);
nand U1105 (N_1105,N_473,N_691);
nand U1106 (N_1106,N_505,N_530);
and U1107 (N_1107,N_123,N_184);
nand U1108 (N_1108,N_537,N_915);
and U1109 (N_1109,N_270,N_153);
and U1110 (N_1110,N_207,N_77);
nand U1111 (N_1111,N_185,N_73);
and U1112 (N_1112,N_875,N_541);
nand U1113 (N_1113,N_961,N_697);
or U1114 (N_1114,N_620,N_845);
and U1115 (N_1115,N_47,N_772);
or U1116 (N_1116,N_958,N_333);
or U1117 (N_1117,N_438,N_12);
nand U1118 (N_1118,N_671,N_24);
nand U1119 (N_1119,N_81,N_950);
nor U1120 (N_1120,N_766,N_229);
nand U1121 (N_1121,N_323,N_417);
nand U1122 (N_1122,N_382,N_820);
and U1123 (N_1123,N_871,N_283);
nor U1124 (N_1124,N_886,N_764);
or U1125 (N_1125,N_638,N_489);
and U1126 (N_1126,N_928,N_931);
and U1127 (N_1127,N_666,N_339);
or U1128 (N_1128,N_160,N_425);
or U1129 (N_1129,N_732,N_142);
and U1130 (N_1130,N_734,N_854);
nor U1131 (N_1131,N_660,N_676);
nor U1132 (N_1132,N_175,N_280);
or U1133 (N_1133,N_183,N_431);
and U1134 (N_1134,N_862,N_210);
nor U1135 (N_1135,N_905,N_841);
or U1136 (N_1136,N_553,N_334);
nand U1137 (N_1137,N_101,N_355);
nor U1138 (N_1138,N_380,N_148);
xnor U1139 (N_1139,N_793,N_196);
nor U1140 (N_1140,N_39,N_137);
xor U1141 (N_1141,N_885,N_596);
or U1142 (N_1142,N_64,N_255);
nor U1143 (N_1143,N_222,N_275);
nor U1144 (N_1144,N_347,N_22);
and U1145 (N_1145,N_873,N_177);
and U1146 (N_1146,N_220,N_603);
nand U1147 (N_1147,N_214,N_460);
nand U1148 (N_1148,N_955,N_410);
and U1149 (N_1149,N_597,N_737);
nand U1150 (N_1150,N_412,N_524);
and U1151 (N_1151,N_166,N_791);
nor U1152 (N_1152,N_648,N_892);
nor U1153 (N_1153,N_949,N_178);
and U1154 (N_1154,N_920,N_944);
nand U1155 (N_1155,N_527,N_654);
or U1156 (N_1156,N_554,N_834);
or U1157 (N_1157,N_493,N_636);
or U1158 (N_1158,N_61,N_453);
nor U1159 (N_1159,N_982,N_595);
or U1160 (N_1160,N_763,N_45);
nand U1161 (N_1161,N_467,N_399);
or U1162 (N_1162,N_60,N_752);
nor U1163 (N_1163,N_599,N_774);
xnor U1164 (N_1164,N_212,N_27);
nand U1165 (N_1165,N_36,N_725);
nand U1166 (N_1166,N_107,N_158);
or U1167 (N_1167,N_721,N_750);
xor U1168 (N_1168,N_644,N_231);
and U1169 (N_1169,N_758,N_816);
nor U1170 (N_1170,N_13,N_326);
nor U1171 (N_1171,N_857,N_441);
and U1172 (N_1172,N_977,N_616);
and U1173 (N_1173,N_865,N_390);
nor U1174 (N_1174,N_663,N_476);
nor U1175 (N_1175,N_881,N_374);
and U1176 (N_1176,N_564,N_975);
nand U1177 (N_1177,N_847,N_716);
and U1178 (N_1178,N_151,N_532);
and U1179 (N_1179,N_227,N_639);
or U1180 (N_1180,N_951,N_385);
and U1181 (N_1181,N_428,N_506);
nor U1182 (N_1182,N_429,N_607);
or U1183 (N_1183,N_810,N_563);
xor U1184 (N_1184,N_88,N_548);
nor U1185 (N_1185,N_482,N_288);
nor U1186 (N_1186,N_461,N_940);
nand U1187 (N_1187,N_304,N_269);
nor U1188 (N_1188,N_262,N_914);
xnor U1189 (N_1189,N_726,N_895);
nand U1190 (N_1190,N_466,N_14);
nor U1191 (N_1191,N_418,N_852);
nor U1192 (N_1192,N_5,N_746);
or U1193 (N_1193,N_225,N_161);
nand U1194 (N_1194,N_381,N_880);
or U1195 (N_1195,N_545,N_606);
nand U1196 (N_1196,N_848,N_303);
or U1197 (N_1197,N_974,N_633);
and U1198 (N_1198,N_250,N_511);
or U1199 (N_1199,N_818,N_495);
and U1200 (N_1200,N_863,N_72);
or U1201 (N_1201,N_959,N_249);
nor U1202 (N_1202,N_646,N_528);
xnor U1203 (N_1203,N_388,N_579);
nand U1204 (N_1204,N_305,N_712);
xor U1205 (N_1205,N_853,N_192);
xnor U1206 (N_1206,N_807,N_514);
nor U1207 (N_1207,N_256,N_315);
or U1208 (N_1208,N_169,N_703);
or U1209 (N_1209,N_194,N_138);
xor U1210 (N_1210,N_272,N_546);
and U1211 (N_1211,N_631,N_197);
nor U1212 (N_1212,N_868,N_836);
and U1213 (N_1213,N_59,N_833);
nand U1214 (N_1214,N_883,N_615);
and U1215 (N_1215,N_760,N_580);
and U1216 (N_1216,N_979,N_945);
xnor U1217 (N_1217,N_781,N_206);
or U1218 (N_1218,N_500,N_704);
nand U1219 (N_1219,N_234,N_215);
nand U1220 (N_1220,N_972,N_309);
nor U1221 (N_1221,N_121,N_808);
nor U1222 (N_1222,N_578,N_635);
or U1223 (N_1223,N_379,N_331);
and U1224 (N_1224,N_416,N_573);
and U1225 (N_1225,N_79,N_93);
nand U1226 (N_1226,N_814,N_962);
or U1227 (N_1227,N_394,N_327);
nor U1228 (N_1228,N_46,N_95);
xor U1229 (N_1229,N_832,N_901);
nand U1230 (N_1230,N_939,N_910);
nand U1231 (N_1231,N_235,N_103);
nor U1232 (N_1232,N_219,N_536);
or U1233 (N_1233,N_42,N_366);
or U1234 (N_1234,N_368,N_916);
and U1235 (N_1235,N_66,N_152);
nor U1236 (N_1236,N_276,N_795);
or U1237 (N_1237,N_878,N_965);
nand U1238 (N_1238,N_198,N_634);
and U1239 (N_1239,N_550,N_377);
nand U1240 (N_1240,N_422,N_299);
nor U1241 (N_1241,N_324,N_819);
or U1242 (N_1242,N_943,N_976);
or U1243 (N_1243,N_661,N_993);
or U1244 (N_1244,N_882,N_287);
nor U1245 (N_1245,N_652,N_587);
xnor U1246 (N_1246,N_188,N_300);
or U1247 (N_1247,N_559,N_773);
nand U1248 (N_1248,N_290,N_124);
and U1249 (N_1249,N_34,N_182);
nor U1250 (N_1250,N_224,N_392);
nand U1251 (N_1251,N_415,N_371);
or U1252 (N_1252,N_830,N_365);
or U1253 (N_1253,N_112,N_297);
nor U1254 (N_1254,N_113,N_159);
or U1255 (N_1255,N_556,N_437);
nor U1256 (N_1256,N_384,N_23);
or U1257 (N_1257,N_796,N_903);
and U1258 (N_1258,N_948,N_322);
and U1259 (N_1259,N_451,N_409);
and U1260 (N_1260,N_251,N_585);
nor U1261 (N_1261,N_90,N_228);
and U1262 (N_1262,N_389,N_488);
nor U1263 (N_1263,N_549,N_432);
and U1264 (N_1264,N_286,N_813);
xor U1265 (N_1265,N_240,N_731);
or U1266 (N_1266,N_310,N_340);
nor U1267 (N_1267,N_254,N_264);
or U1268 (N_1268,N_529,N_522);
or U1269 (N_1269,N_681,N_132);
and U1270 (N_1270,N_899,N_87);
nand U1271 (N_1271,N_918,N_768);
or U1272 (N_1272,N_849,N_566);
and U1273 (N_1273,N_929,N_736);
nor U1274 (N_1274,N_363,N_780);
nor U1275 (N_1275,N_565,N_329);
nand U1276 (N_1276,N_260,N_981);
nor U1277 (N_1277,N_217,N_179);
or U1278 (N_1278,N_614,N_167);
and U1279 (N_1279,N_21,N_912);
or U1280 (N_1280,N_176,N_941);
nand U1281 (N_1281,N_724,N_802);
and U1282 (N_1282,N_6,N_419);
and U1283 (N_1283,N_247,N_729);
nor U1284 (N_1284,N_41,N_653);
and U1285 (N_1285,N_111,N_349);
nand U1286 (N_1286,N_470,N_71);
nor U1287 (N_1287,N_471,N_797);
and U1288 (N_1288,N_710,N_557);
and U1289 (N_1289,N_740,N_806);
nor U1290 (N_1290,N_313,N_427);
nor U1291 (N_1291,N_338,N_622);
nand U1292 (N_1292,N_246,N_226);
or U1293 (N_1293,N_325,N_472);
xnor U1294 (N_1294,N_694,N_433);
nand U1295 (N_1295,N_985,N_367);
or U1296 (N_1296,N_492,N_335);
and U1297 (N_1297,N_574,N_515);
nand U1298 (N_1298,N_165,N_267);
xor U1299 (N_1299,N_591,N_512);
or U1300 (N_1300,N_907,N_817);
nor U1301 (N_1301,N_58,N_449);
nand U1302 (N_1302,N_611,N_821);
nor U1303 (N_1303,N_971,N_887);
nand U1304 (N_1304,N_569,N_497);
or U1305 (N_1305,N_477,N_28);
and U1306 (N_1306,N_200,N_487);
nor U1307 (N_1307,N_199,N_665);
or U1308 (N_1308,N_140,N_730);
and U1309 (N_1309,N_128,N_519);
and U1310 (N_1310,N_65,N_526);
or U1311 (N_1311,N_218,N_345);
nor U1312 (N_1312,N_889,N_330);
or U1313 (N_1313,N_682,N_922);
or U1314 (N_1314,N_727,N_786);
nand U1315 (N_1315,N_201,N_193);
or U1316 (N_1316,N_481,N_455);
nand U1317 (N_1317,N_908,N_846);
nor U1318 (N_1318,N_104,N_932);
nand U1319 (N_1319,N_669,N_684);
nand U1320 (N_1320,N_469,N_628);
nand U1321 (N_1321,N_213,N_242);
nand U1322 (N_1322,N_404,N_401);
nand U1323 (N_1323,N_662,N_523);
nand U1324 (N_1324,N_295,N_759);
and U1325 (N_1325,N_129,N_408);
nor U1326 (N_1326,N_826,N_741);
or U1327 (N_1327,N_253,N_593);
nand U1328 (N_1328,N_18,N_289);
or U1329 (N_1329,N_115,N_672);
or U1330 (N_1330,N_244,N_191);
or U1331 (N_1331,N_436,N_296);
nand U1332 (N_1332,N_963,N_361);
or U1333 (N_1333,N_458,N_80);
xor U1334 (N_1334,N_829,N_964);
nand U1335 (N_1335,N_641,N_776);
or U1336 (N_1336,N_491,N_706);
nor U1337 (N_1337,N_656,N_674);
nand U1338 (N_1338,N_479,N_257);
and U1339 (N_1339,N_799,N_531);
nand U1340 (N_1340,N_478,N_673);
nor U1341 (N_1341,N_866,N_292);
or U1342 (N_1342,N_172,N_51);
or U1343 (N_1343,N_989,N_186);
or U1344 (N_1344,N_171,N_114);
xnor U1345 (N_1345,N_62,N_874);
nor U1346 (N_1346,N_538,N_518);
and U1347 (N_1347,N_714,N_67);
or U1348 (N_1348,N_0,N_983);
nor U1349 (N_1349,N_134,N_448);
and U1350 (N_1350,N_503,N_957);
nor U1351 (N_1351,N_998,N_119);
nor U1352 (N_1352,N_2,N_698);
nand U1353 (N_1353,N_867,N_15);
nor U1354 (N_1354,N_452,N_397);
nand U1355 (N_1355,N_52,N_130);
nand U1356 (N_1356,N_205,N_902);
nor U1357 (N_1357,N_369,N_525);
or U1358 (N_1358,N_483,N_475);
xor U1359 (N_1359,N_439,N_583);
nand U1360 (N_1360,N_50,N_651);
and U1361 (N_1361,N_221,N_311);
or U1362 (N_1362,N_490,N_328);
and U1363 (N_1363,N_952,N_97);
and U1364 (N_1364,N_344,N_570);
nor U1365 (N_1365,N_859,N_747);
nand U1366 (N_1366,N_386,N_767);
xor U1367 (N_1367,N_189,N_337);
and U1368 (N_1368,N_232,N_265);
and U1369 (N_1369,N_274,N_803);
or U1370 (N_1370,N_757,N_598);
and U1371 (N_1371,N_897,N_947);
or U1372 (N_1372,N_535,N_29);
nor U1373 (N_1373,N_552,N_755);
or U1374 (N_1374,N_856,N_9);
nand U1375 (N_1375,N_898,N_805);
or U1376 (N_1376,N_761,N_411);
nor U1377 (N_1377,N_284,N_840);
nor U1378 (N_1378,N_116,N_92);
nor U1379 (N_1379,N_98,N_987);
nor U1380 (N_1380,N_364,N_504);
nand U1381 (N_1381,N_838,N_850);
or U1382 (N_1382,N_3,N_316);
nor U1383 (N_1383,N_751,N_804);
nor U1384 (N_1384,N_125,N_695);
or U1385 (N_1385,N_986,N_508);
and U1386 (N_1386,N_911,N_187);
nor U1387 (N_1387,N_794,N_150);
and U1388 (N_1388,N_435,N_630);
and U1389 (N_1389,N_426,N_960);
or U1390 (N_1390,N_319,N_424);
xor U1391 (N_1391,N_925,N_919);
or U1392 (N_1392,N_649,N_154);
xor U1393 (N_1393,N_904,N_913);
nor U1394 (N_1394,N_589,N_659);
and U1395 (N_1395,N_756,N_346);
or U1396 (N_1396,N_837,N_702);
or U1397 (N_1397,N_973,N_314);
nor U1398 (N_1398,N_122,N_383);
nor U1399 (N_1399,N_499,N_202);
nor U1400 (N_1400,N_258,N_828);
xnor U1401 (N_1401,N_687,N_54);
and U1402 (N_1402,N_777,N_954);
or U1403 (N_1403,N_447,N_692);
or U1404 (N_1404,N_170,N_990);
or U1405 (N_1405,N_966,N_216);
and U1406 (N_1406,N_420,N_376);
nand U1407 (N_1407,N_978,N_102);
nor U1408 (N_1408,N_827,N_547);
xor U1409 (N_1409,N_239,N_769);
nand U1410 (N_1410,N_647,N_395);
and U1411 (N_1411,N_594,N_748);
or U1412 (N_1412,N_414,N_601);
or U1413 (N_1413,N_89,N_864);
nor U1414 (N_1414,N_701,N_749);
nand U1415 (N_1415,N_700,N_743);
or U1416 (N_1416,N_988,N_25);
and U1417 (N_1417,N_320,N_675);
nor U1418 (N_1418,N_543,N_233);
nor U1419 (N_1419,N_277,N_373);
nor U1420 (N_1420,N_824,N_32);
and U1421 (N_1421,N_407,N_968);
and U1422 (N_1422,N_474,N_173);
nand U1423 (N_1423,N_801,N_787);
nor U1424 (N_1424,N_612,N_798);
nor U1425 (N_1425,N_91,N_713);
nand U1426 (N_1426,N_855,N_387);
nand U1427 (N_1427,N_884,N_84);
nand U1428 (N_1428,N_680,N_360);
or U1429 (N_1429,N_400,N_291);
or U1430 (N_1430,N_468,N_268);
or U1431 (N_1431,N_906,N_539);
nor U1432 (N_1432,N_496,N_486);
nand U1433 (N_1433,N_443,N_139);
or U1434 (N_1434,N_624,N_621);
and U1435 (N_1435,N_696,N_946);
or U1436 (N_1436,N_720,N_618);
nor U1437 (N_1437,N_480,N_131);
nor U1438 (N_1438,N_664,N_76);
nand U1439 (N_1439,N_822,N_645);
nor U1440 (N_1440,N_953,N_560);
and U1441 (N_1441,N_575,N_118);
nand U1442 (N_1442,N_809,N_372);
nand U1443 (N_1443,N_924,N_800);
and U1444 (N_1444,N_709,N_843);
nor U1445 (N_1445,N_31,N_393);
nand U1446 (N_1446,N_100,N_306);
nor U1447 (N_1447,N_354,N_835);
and U1448 (N_1448,N_35,N_723);
or U1449 (N_1449,N_243,N_245);
and U1450 (N_1450,N_318,N_204);
or U1451 (N_1451,N_779,N_494);
or U1452 (N_1452,N_126,N_203);
nand U1453 (N_1453,N_937,N_685);
and U1454 (N_1454,N_590,N_298);
or U1455 (N_1455,N_450,N_586);
nand U1456 (N_1456,N_891,N_282);
and U1457 (N_1457,N_582,N_86);
and U1458 (N_1458,N_567,N_668);
nor U1459 (N_1459,N_38,N_592);
or U1460 (N_1460,N_825,N_271);
or U1461 (N_1461,N_85,N_223);
nor U1462 (N_1462,N_155,N_792);
or U1463 (N_1463,N_782,N_507);
nand U1464 (N_1464,N_688,N_353);
nor U1465 (N_1465,N_742,N_790);
nor U1466 (N_1466,N_82,N_551);
nand U1467 (N_1467,N_600,N_332);
or U1468 (N_1468,N_63,N_434);
nand U1469 (N_1469,N_542,N_252);
nand U1470 (N_1470,N_997,N_936);
and U1471 (N_1471,N_20,N_312);
nor U1472 (N_1472,N_623,N_502);
nor U1473 (N_1473,N_465,N_33);
nand U1474 (N_1474,N_992,N_459);
and U1475 (N_1475,N_147,N_281);
xnor U1476 (N_1476,N_351,N_642);
or U1477 (N_1477,N_146,N_83);
and U1478 (N_1478,N_463,N_141);
or U1479 (N_1479,N_872,N_180);
nor U1480 (N_1480,N_683,N_738);
nor U1481 (N_1481,N_844,N_457);
and U1482 (N_1482,N_831,N_658);
nor U1483 (N_1483,N_711,N_26);
xnor U1484 (N_1484,N_94,N_626);
or U1485 (N_1485,N_273,N_143);
nor U1486 (N_1486,N_352,N_40);
or U1487 (N_1487,N_632,N_336);
or U1488 (N_1488,N_900,N_771);
xor U1489 (N_1489,N_718,N_359);
and U1490 (N_1490,N_842,N_917);
nand U1491 (N_1491,N_858,N_378);
nor U1492 (N_1492,N_105,N_195);
or U1493 (N_1493,N_109,N_230);
xor U1494 (N_1494,N_241,N_110);
nand U1495 (N_1495,N_994,N_785);
and U1496 (N_1496,N_174,N_106);
and U1497 (N_1497,N_934,N_108);
nor U1498 (N_1498,N_513,N_403);
nor U1499 (N_1499,N_637,N_927);
nor U1500 (N_1500,N_920,N_602);
nand U1501 (N_1501,N_140,N_475);
nor U1502 (N_1502,N_895,N_140);
nor U1503 (N_1503,N_158,N_706);
or U1504 (N_1504,N_969,N_452);
or U1505 (N_1505,N_352,N_148);
or U1506 (N_1506,N_464,N_701);
or U1507 (N_1507,N_628,N_63);
nand U1508 (N_1508,N_495,N_976);
and U1509 (N_1509,N_347,N_316);
nor U1510 (N_1510,N_762,N_704);
nand U1511 (N_1511,N_982,N_960);
nand U1512 (N_1512,N_663,N_148);
nand U1513 (N_1513,N_440,N_178);
nand U1514 (N_1514,N_183,N_562);
or U1515 (N_1515,N_676,N_814);
nand U1516 (N_1516,N_689,N_284);
nand U1517 (N_1517,N_104,N_10);
and U1518 (N_1518,N_529,N_205);
and U1519 (N_1519,N_472,N_666);
and U1520 (N_1520,N_281,N_717);
and U1521 (N_1521,N_28,N_283);
nand U1522 (N_1522,N_109,N_617);
nand U1523 (N_1523,N_10,N_840);
and U1524 (N_1524,N_650,N_903);
or U1525 (N_1525,N_43,N_16);
and U1526 (N_1526,N_925,N_84);
or U1527 (N_1527,N_510,N_653);
nand U1528 (N_1528,N_26,N_577);
nand U1529 (N_1529,N_774,N_747);
nor U1530 (N_1530,N_348,N_193);
or U1531 (N_1531,N_402,N_265);
and U1532 (N_1532,N_838,N_653);
nand U1533 (N_1533,N_673,N_13);
and U1534 (N_1534,N_280,N_405);
nand U1535 (N_1535,N_536,N_319);
xor U1536 (N_1536,N_602,N_441);
nand U1537 (N_1537,N_164,N_488);
or U1538 (N_1538,N_118,N_389);
or U1539 (N_1539,N_212,N_61);
nor U1540 (N_1540,N_968,N_712);
nand U1541 (N_1541,N_731,N_144);
or U1542 (N_1542,N_688,N_9);
and U1543 (N_1543,N_942,N_500);
nand U1544 (N_1544,N_928,N_824);
or U1545 (N_1545,N_637,N_311);
and U1546 (N_1546,N_447,N_603);
and U1547 (N_1547,N_457,N_959);
nor U1548 (N_1548,N_218,N_229);
nand U1549 (N_1549,N_972,N_785);
and U1550 (N_1550,N_939,N_903);
and U1551 (N_1551,N_193,N_272);
nor U1552 (N_1552,N_362,N_478);
and U1553 (N_1553,N_176,N_57);
nor U1554 (N_1554,N_961,N_705);
nor U1555 (N_1555,N_389,N_5);
nand U1556 (N_1556,N_849,N_655);
nand U1557 (N_1557,N_116,N_468);
or U1558 (N_1558,N_672,N_420);
or U1559 (N_1559,N_614,N_506);
nand U1560 (N_1560,N_431,N_713);
nor U1561 (N_1561,N_841,N_164);
nor U1562 (N_1562,N_573,N_71);
or U1563 (N_1563,N_368,N_47);
nand U1564 (N_1564,N_842,N_188);
and U1565 (N_1565,N_501,N_630);
and U1566 (N_1566,N_829,N_554);
and U1567 (N_1567,N_610,N_413);
or U1568 (N_1568,N_48,N_65);
nand U1569 (N_1569,N_47,N_824);
nand U1570 (N_1570,N_767,N_502);
xor U1571 (N_1571,N_664,N_16);
or U1572 (N_1572,N_782,N_24);
and U1573 (N_1573,N_245,N_370);
nand U1574 (N_1574,N_668,N_747);
or U1575 (N_1575,N_584,N_803);
nand U1576 (N_1576,N_279,N_482);
nand U1577 (N_1577,N_666,N_226);
nor U1578 (N_1578,N_676,N_54);
and U1579 (N_1579,N_708,N_276);
nand U1580 (N_1580,N_485,N_680);
nand U1581 (N_1581,N_772,N_212);
nand U1582 (N_1582,N_553,N_800);
or U1583 (N_1583,N_455,N_751);
nand U1584 (N_1584,N_910,N_140);
xnor U1585 (N_1585,N_806,N_15);
and U1586 (N_1586,N_883,N_421);
nand U1587 (N_1587,N_797,N_928);
or U1588 (N_1588,N_816,N_455);
nor U1589 (N_1589,N_892,N_659);
or U1590 (N_1590,N_167,N_246);
and U1591 (N_1591,N_982,N_578);
nand U1592 (N_1592,N_988,N_275);
xor U1593 (N_1593,N_666,N_819);
and U1594 (N_1594,N_85,N_860);
and U1595 (N_1595,N_912,N_394);
and U1596 (N_1596,N_366,N_205);
or U1597 (N_1597,N_732,N_805);
and U1598 (N_1598,N_969,N_337);
or U1599 (N_1599,N_622,N_154);
nor U1600 (N_1600,N_793,N_922);
and U1601 (N_1601,N_861,N_683);
nand U1602 (N_1602,N_190,N_659);
and U1603 (N_1603,N_625,N_3);
or U1604 (N_1604,N_355,N_489);
nor U1605 (N_1605,N_916,N_474);
and U1606 (N_1606,N_655,N_913);
nand U1607 (N_1607,N_192,N_841);
nor U1608 (N_1608,N_514,N_662);
or U1609 (N_1609,N_495,N_234);
and U1610 (N_1610,N_892,N_62);
nand U1611 (N_1611,N_115,N_845);
nor U1612 (N_1612,N_438,N_663);
or U1613 (N_1613,N_386,N_649);
nor U1614 (N_1614,N_523,N_592);
and U1615 (N_1615,N_669,N_759);
nand U1616 (N_1616,N_444,N_674);
and U1617 (N_1617,N_666,N_238);
nor U1618 (N_1618,N_344,N_240);
nor U1619 (N_1619,N_921,N_212);
nor U1620 (N_1620,N_84,N_487);
nand U1621 (N_1621,N_794,N_419);
and U1622 (N_1622,N_438,N_101);
nand U1623 (N_1623,N_658,N_346);
or U1624 (N_1624,N_25,N_731);
or U1625 (N_1625,N_112,N_433);
nand U1626 (N_1626,N_110,N_549);
nor U1627 (N_1627,N_916,N_196);
nand U1628 (N_1628,N_322,N_19);
nor U1629 (N_1629,N_915,N_452);
nor U1630 (N_1630,N_837,N_364);
and U1631 (N_1631,N_367,N_231);
xnor U1632 (N_1632,N_626,N_130);
or U1633 (N_1633,N_780,N_123);
or U1634 (N_1634,N_980,N_665);
nand U1635 (N_1635,N_435,N_917);
xnor U1636 (N_1636,N_7,N_25);
or U1637 (N_1637,N_20,N_619);
or U1638 (N_1638,N_226,N_877);
nand U1639 (N_1639,N_519,N_19);
or U1640 (N_1640,N_888,N_908);
nand U1641 (N_1641,N_770,N_841);
xor U1642 (N_1642,N_949,N_790);
or U1643 (N_1643,N_911,N_384);
or U1644 (N_1644,N_143,N_321);
nor U1645 (N_1645,N_781,N_112);
or U1646 (N_1646,N_395,N_957);
nor U1647 (N_1647,N_101,N_574);
nor U1648 (N_1648,N_880,N_843);
and U1649 (N_1649,N_230,N_119);
nor U1650 (N_1650,N_756,N_14);
nor U1651 (N_1651,N_265,N_464);
nand U1652 (N_1652,N_492,N_885);
nor U1653 (N_1653,N_127,N_102);
nor U1654 (N_1654,N_150,N_138);
and U1655 (N_1655,N_107,N_844);
and U1656 (N_1656,N_655,N_673);
nor U1657 (N_1657,N_685,N_934);
nor U1658 (N_1658,N_320,N_45);
nor U1659 (N_1659,N_157,N_819);
and U1660 (N_1660,N_688,N_166);
and U1661 (N_1661,N_369,N_31);
or U1662 (N_1662,N_405,N_183);
and U1663 (N_1663,N_597,N_369);
nand U1664 (N_1664,N_448,N_806);
or U1665 (N_1665,N_42,N_315);
nor U1666 (N_1666,N_813,N_644);
or U1667 (N_1667,N_646,N_415);
nand U1668 (N_1668,N_441,N_558);
or U1669 (N_1669,N_458,N_885);
or U1670 (N_1670,N_107,N_698);
nor U1671 (N_1671,N_375,N_933);
nor U1672 (N_1672,N_256,N_485);
and U1673 (N_1673,N_149,N_792);
or U1674 (N_1674,N_599,N_146);
and U1675 (N_1675,N_287,N_456);
nor U1676 (N_1676,N_331,N_39);
nand U1677 (N_1677,N_892,N_765);
or U1678 (N_1678,N_986,N_542);
nor U1679 (N_1679,N_636,N_68);
or U1680 (N_1680,N_172,N_210);
and U1681 (N_1681,N_713,N_12);
or U1682 (N_1682,N_926,N_913);
nand U1683 (N_1683,N_28,N_999);
nand U1684 (N_1684,N_850,N_967);
and U1685 (N_1685,N_5,N_541);
xnor U1686 (N_1686,N_716,N_460);
nor U1687 (N_1687,N_18,N_623);
or U1688 (N_1688,N_222,N_142);
nand U1689 (N_1689,N_685,N_553);
nand U1690 (N_1690,N_552,N_48);
nand U1691 (N_1691,N_54,N_743);
and U1692 (N_1692,N_820,N_517);
and U1693 (N_1693,N_573,N_796);
nand U1694 (N_1694,N_298,N_168);
or U1695 (N_1695,N_306,N_338);
and U1696 (N_1696,N_936,N_578);
nand U1697 (N_1697,N_98,N_417);
or U1698 (N_1698,N_176,N_30);
nand U1699 (N_1699,N_629,N_973);
nand U1700 (N_1700,N_920,N_151);
nor U1701 (N_1701,N_403,N_952);
nand U1702 (N_1702,N_427,N_4);
and U1703 (N_1703,N_416,N_292);
and U1704 (N_1704,N_765,N_513);
nor U1705 (N_1705,N_837,N_864);
or U1706 (N_1706,N_93,N_125);
nand U1707 (N_1707,N_956,N_518);
nand U1708 (N_1708,N_806,N_944);
and U1709 (N_1709,N_874,N_144);
nor U1710 (N_1710,N_563,N_287);
or U1711 (N_1711,N_890,N_64);
nand U1712 (N_1712,N_701,N_160);
nor U1713 (N_1713,N_580,N_27);
nor U1714 (N_1714,N_94,N_838);
xor U1715 (N_1715,N_345,N_975);
nor U1716 (N_1716,N_272,N_808);
or U1717 (N_1717,N_334,N_69);
xor U1718 (N_1718,N_74,N_834);
or U1719 (N_1719,N_157,N_82);
nand U1720 (N_1720,N_154,N_715);
nand U1721 (N_1721,N_289,N_977);
and U1722 (N_1722,N_623,N_114);
nand U1723 (N_1723,N_619,N_621);
nor U1724 (N_1724,N_871,N_619);
nor U1725 (N_1725,N_971,N_261);
and U1726 (N_1726,N_36,N_604);
nor U1727 (N_1727,N_897,N_630);
nor U1728 (N_1728,N_333,N_877);
and U1729 (N_1729,N_766,N_912);
nand U1730 (N_1730,N_727,N_822);
and U1731 (N_1731,N_187,N_543);
nand U1732 (N_1732,N_935,N_81);
and U1733 (N_1733,N_776,N_943);
nand U1734 (N_1734,N_476,N_988);
xor U1735 (N_1735,N_866,N_8);
or U1736 (N_1736,N_905,N_148);
or U1737 (N_1737,N_796,N_508);
nor U1738 (N_1738,N_528,N_300);
nor U1739 (N_1739,N_619,N_305);
nand U1740 (N_1740,N_346,N_860);
nor U1741 (N_1741,N_729,N_347);
nor U1742 (N_1742,N_959,N_448);
and U1743 (N_1743,N_499,N_9);
and U1744 (N_1744,N_785,N_932);
and U1745 (N_1745,N_202,N_873);
nand U1746 (N_1746,N_81,N_638);
nand U1747 (N_1747,N_145,N_343);
and U1748 (N_1748,N_681,N_345);
and U1749 (N_1749,N_605,N_798);
and U1750 (N_1750,N_380,N_940);
and U1751 (N_1751,N_335,N_668);
or U1752 (N_1752,N_385,N_901);
nor U1753 (N_1753,N_941,N_52);
and U1754 (N_1754,N_332,N_757);
and U1755 (N_1755,N_318,N_534);
nand U1756 (N_1756,N_761,N_77);
and U1757 (N_1757,N_265,N_817);
and U1758 (N_1758,N_843,N_650);
nor U1759 (N_1759,N_860,N_234);
and U1760 (N_1760,N_183,N_265);
and U1761 (N_1761,N_391,N_813);
and U1762 (N_1762,N_326,N_124);
xnor U1763 (N_1763,N_911,N_897);
nor U1764 (N_1764,N_203,N_328);
nor U1765 (N_1765,N_505,N_761);
and U1766 (N_1766,N_410,N_920);
or U1767 (N_1767,N_565,N_957);
or U1768 (N_1768,N_804,N_453);
or U1769 (N_1769,N_706,N_504);
nand U1770 (N_1770,N_410,N_350);
nor U1771 (N_1771,N_108,N_998);
nor U1772 (N_1772,N_94,N_961);
nor U1773 (N_1773,N_518,N_182);
or U1774 (N_1774,N_141,N_347);
nor U1775 (N_1775,N_363,N_53);
nor U1776 (N_1776,N_745,N_123);
and U1777 (N_1777,N_377,N_732);
nor U1778 (N_1778,N_282,N_513);
nor U1779 (N_1779,N_155,N_819);
nor U1780 (N_1780,N_232,N_920);
or U1781 (N_1781,N_957,N_327);
and U1782 (N_1782,N_595,N_466);
nand U1783 (N_1783,N_5,N_33);
and U1784 (N_1784,N_691,N_60);
or U1785 (N_1785,N_233,N_88);
and U1786 (N_1786,N_420,N_638);
or U1787 (N_1787,N_909,N_561);
xor U1788 (N_1788,N_655,N_235);
nand U1789 (N_1789,N_353,N_103);
or U1790 (N_1790,N_812,N_381);
and U1791 (N_1791,N_264,N_981);
and U1792 (N_1792,N_450,N_28);
or U1793 (N_1793,N_387,N_652);
or U1794 (N_1794,N_410,N_622);
nor U1795 (N_1795,N_948,N_288);
nor U1796 (N_1796,N_730,N_283);
or U1797 (N_1797,N_936,N_750);
nand U1798 (N_1798,N_180,N_928);
nor U1799 (N_1799,N_309,N_483);
nor U1800 (N_1800,N_584,N_856);
nand U1801 (N_1801,N_434,N_86);
nand U1802 (N_1802,N_106,N_454);
and U1803 (N_1803,N_386,N_778);
and U1804 (N_1804,N_116,N_684);
nand U1805 (N_1805,N_141,N_246);
or U1806 (N_1806,N_946,N_748);
or U1807 (N_1807,N_763,N_728);
or U1808 (N_1808,N_620,N_58);
nand U1809 (N_1809,N_33,N_107);
or U1810 (N_1810,N_598,N_515);
or U1811 (N_1811,N_459,N_547);
nor U1812 (N_1812,N_502,N_199);
and U1813 (N_1813,N_317,N_607);
nand U1814 (N_1814,N_719,N_123);
nor U1815 (N_1815,N_552,N_512);
nor U1816 (N_1816,N_572,N_795);
nand U1817 (N_1817,N_531,N_181);
or U1818 (N_1818,N_753,N_462);
nor U1819 (N_1819,N_262,N_342);
or U1820 (N_1820,N_719,N_293);
and U1821 (N_1821,N_27,N_979);
nor U1822 (N_1822,N_97,N_669);
nor U1823 (N_1823,N_929,N_843);
and U1824 (N_1824,N_310,N_501);
xor U1825 (N_1825,N_94,N_218);
and U1826 (N_1826,N_857,N_160);
nor U1827 (N_1827,N_133,N_531);
or U1828 (N_1828,N_93,N_382);
xnor U1829 (N_1829,N_546,N_555);
and U1830 (N_1830,N_85,N_642);
or U1831 (N_1831,N_622,N_383);
nand U1832 (N_1832,N_286,N_271);
or U1833 (N_1833,N_144,N_142);
nand U1834 (N_1834,N_300,N_104);
or U1835 (N_1835,N_150,N_571);
or U1836 (N_1836,N_100,N_909);
nand U1837 (N_1837,N_864,N_153);
nand U1838 (N_1838,N_313,N_505);
nand U1839 (N_1839,N_593,N_974);
nor U1840 (N_1840,N_644,N_722);
or U1841 (N_1841,N_215,N_435);
nand U1842 (N_1842,N_697,N_133);
and U1843 (N_1843,N_428,N_588);
nor U1844 (N_1844,N_817,N_165);
or U1845 (N_1845,N_158,N_698);
nand U1846 (N_1846,N_783,N_2);
nor U1847 (N_1847,N_50,N_993);
nor U1848 (N_1848,N_65,N_752);
or U1849 (N_1849,N_236,N_688);
or U1850 (N_1850,N_369,N_168);
nand U1851 (N_1851,N_789,N_587);
nand U1852 (N_1852,N_793,N_126);
nor U1853 (N_1853,N_987,N_797);
or U1854 (N_1854,N_656,N_777);
or U1855 (N_1855,N_784,N_379);
nand U1856 (N_1856,N_752,N_318);
nor U1857 (N_1857,N_565,N_947);
or U1858 (N_1858,N_552,N_746);
nor U1859 (N_1859,N_621,N_979);
or U1860 (N_1860,N_152,N_389);
or U1861 (N_1861,N_439,N_423);
or U1862 (N_1862,N_87,N_599);
nand U1863 (N_1863,N_879,N_347);
nand U1864 (N_1864,N_721,N_257);
nand U1865 (N_1865,N_106,N_361);
nor U1866 (N_1866,N_398,N_642);
and U1867 (N_1867,N_122,N_981);
or U1868 (N_1868,N_537,N_783);
or U1869 (N_1869,N_616,N_416);
nand U1870 (N_1870,N_316,N_528);
nand U1871 (N_1871,N_309,N_541);
nand U1872 (N_1872,N_424,N_906);
nor U1873 (N_1873,N_642,N_426);
nand U1874 (N_1874,N_566,N_892);
and U1875 (N_1875,N_933,N_795);
nor U1876 (N_1876,N_411,N_386);
or U1877 (N_1877,N_238,N_844);
nand U1878 (N_1878,N_875,N_303);
or U1879 (N_1879,N_348,N_733);
or U1880 (N_1880,N_532,N_548);
nor U1881 (N_1881,N_706,N_56);
nor U1882 (N_1882,N_594,N_798);
or U1883 (N_1883,N_36,N_938);
nor U1884 (N_1884,N_662,N_721);
and U1885 (N_1885,N_864,N_798);
nor U1886 (N_1886,N_528,N_720);
or U1887 (N_1887,N_468,N_477);
and U1888 (N_1888,N_553,N_831);
nor U1889 (N_1889,N_835,N_288);
or U1890 (N_1890,N_710,N_667);
nand U1891 (N_1891,N_835,N_648);
and U1892 (N_1892,N_745,N_35);
nand U1893 (N_1893,N_427,N_471);
nor U1894 (N_1894,N_560,N_33);
or U1895 (N_1895,N_232,N_720);
or U1896 (N_1896,N_719,N_338);
nor U1897 (N_1897,N_388,N_567);
and U1898 (N_1898,N_144,N_276);
nand U1899 (N_1899,N_125,N_55);
nor U1900 (N_1900,N_357,N_690);
and U1901 (N_1901,N_961,N_758);
and U1902 (N_1902,N_88,N_132);
and U1903 (N_1903,N_178,N_631);
and U1904 (N_1904,N_208,N_564);
and U1905 (N_1905,N_439,N_474);
nor U1906 (N_1906,N_684,N_987);
nand U1907 (N_1907,N_125,N_734);
nor U1908 (N_1908,N_107,N_247);
or U1909 (N_1909,N_119,N_77);
or U1910 (N_1910,N_774,N_812);
nand U1911 (N_1911,N_442,N_523);
nand U1912 (N_1912,N_825,N_969);
or U1913 (N_1913,N_620,N_46);
nand U1914 (N_1914,N_636,N_863);
nand U1915 (N_1915,N_905,N_926);
xnor U1916 (N_1916,N_65,N_272);
nand U1917 (N_1917,N_179,N_919);
and U1918 (N_1918,N_830,N_795);
or U1919 (N_1919,N_299,N_976);
nor U1920 (N_1920,N_534,N_470);
nand U1921 (N_1921,N_585,N_384);
nand U1922 (N_1922,N_283,N_960);
nor U1923 (N_1923,N_769,N_763);
and U1924 (N_1924,N_420,N_773);
nand U1925 (N_1925,N_182,N_417);
or U1926 (N_1926,N_935,N_26);
nand U1927 (N_1927,N_310,N_698);
or U1928 (N_1928,N_432,N_928);
and U1929 (N_1929,N_997,N_870);
and U1930 (N_1930,N_885,N_383);
or U1931 (N_1931,N_559,N_655);
and U1932 (N_1932,N_46,N_979);
nor U1933 (N_1933,N_292,N_828);
and U1934 (N_1934,N_332,N_193);
nand U1935 (N_1935,N_983,N_143);
nand U1936 (N_1936,N_753,N_815);
and U1937 (N_1937,N_863,N_216);
nor U1938 (N_1938,N_237,N_924);
xor U1939 (N_1939,N_78,N_4);
nand U1940 (N_1940,N_112,N_379);
nor U1941 (N_1941,N_473,N_524);
and U1942 (N_1942,N_353,N_781);
nor U1943 (N_1943,N_121,N_472);
nor U1944 (N_1944,N_758,N_174);
nand U1945 (N_1945,N_436,N_491);
or U1946 (N_1946,N_535,N_524);
nand U1947 (N_1947,N_769,N_92);
nor U1948 (N_1948,N_317,N_904);
or U1949 (N_1949,N_811,N_126);
and U1950 (N_1950,N_83,N_680);
and U1951 (N_1951,N_669,N_34);
nor U1952 (N_1952,N_129,N_949);
xor U1953 (N_1953,N_66,N_798);
nand U1954 (N_1954,N_420,N_333);
or U1955 (N_1955,N_529,N_894);
or U1956 (N_1956,N_171,N_402);
or U1957 (N_1957,N_945,N_983);
and U1958 (N_1958,N_793,N_177);
and U1959 (N_1959,N_552,N_884);
nor U1960 (N_1960,N_701,N_901);
nand U1961 (N_1961,N_239,N_715);
nand U1962 (N_1962,N_205,N_789);
or U1963 (N_1963,N_622,N_444);
nand U1964 (N_1964,N_629,N_546);
or U1965 (N_1965,N_236,N_250);
or U1966 (N_1966,N_601,N_209);
nand U1967 (N_1967,N_146,N_420);
nor U1968 (N_1968,N_786,N_861);
and U1969 (N_1969,N_31,N_924);
nand U1970 (N_1970,N_385,N_375);
or U1971 (N_1971,N_466,N_171);
or U1972 (N_1972,N_103,N_83);
nand U1973 (N_1973,N_82,N_330);
and U1974 (N_1974,N_634,N_526);
nor U1975 (N_1975,N_598,N_754);
nand U1976 (N_1976,N_121,N_251);
and U1977 (N_1977,N_181,N_567);
or U1978 (N_1978,N_509,N_943);
or U1979 (N_1979,N_643,N_872);
nand U1980 (N_1980,N_585,N_335);
or U1981 (N_1981,N_677,N_526);
nor U1982 (N_1982,N_111,N_506);
or U1983 (N_1983,N_825,N_774);
or U1984 (N_1984,N_481,N_183);
and U1985 (N_1985,N_155,N_740);
nand U1986 (N_1986,N_807,N_227);
nand U1987 (N_1987,N_105,N_28);
nand U1988 (N_1988,N_869,N_139);
or U1989 (N_1989,N_894,N_766);
and U1990 (N_1990,N_203,N_852);
or U1991 (N_1991,N_405,N_402);
nor U1992 (N_1992,N_609,N_345);
nor U1993 (N_1993,N_220,N_408);
or U1994 (N_1994,N_408,N_660);
xnor U1995 (N_1995,N_237,N_191);
nor U1996 (N_1996,N_546,N_264);
nand U1997 (N_1997,N_858,N_431);
xnor U1998 (N_1998,N_393,N_954);
nor U1999 (N_1999,N_363,N_482);
nand U2000 (N_2000,N_1124,N_1071);
nor U2001 (N_2001,N_1588,N_1602);
and U2002 (N_2002,N_1273,N_1385);
nor U2003 (N_2003,N_1682,N_1018);
or U2004 (N_2004,N_1663,N_1313);
nor U2005 (N_2005,N_1964,N_1428);
nand U2006 (N_2006,N_1350,N_1032);
nor U2007 (N_2007,N_1025,N_1337);
nor U2008 (N_2008,N_1779,N_1275);
or U2009 (N_2009,N_1469,N_1811);
or U2010 (N_2010,N_1534,N_1553);
nand U2011 (N_2011,N_1696,N_1103);
nor U2012 (N_2012,N_1339,N_1014);
or U2013 (N_2013,N_1685,N_1919);
nor U2014 (N_2014,N_1826,N_1783);
nand U2015 (N_2015,N_1700,N_1116);
and U2016 (N_2016,N_1804,N_1597);
nand U2017 (N_2017,N_1775,N_1801);
nor U2018 (N_2018,N_1031,N_1105);
or U2019 (N_2019,N_1421,N_1007);
or U2020 (N_2020,N_1211,N_1763);
nand U2021 (N_2021,N_1747,N_1420);
or U2022 (N_2022,N_1302,N_1311);
nor U2023 (N_2023,N_1136,N_1761);
and U2024 (N_2024,N_1147,N_1331);
and U2025 (N_2025,N_1314,N_1830);
xnor U2026 (N_2026,N_1940,N_1265);
nor U2027 (N_2027,N_1338,N_1047);
nand U2028 (N_2028,N_1152,N_1217);
and U2029 (N_2029,N_1299,N_1294);
nor U2030 (N_2030,N_1039,N_1026);
nand U2031 (N_2031,N_1959,N_1794);
nor U2032 (N_2032,N_1080,N_1596);
xor U2033 (N_2033,N_1184,N_1762);
and U2034 (N_2034,N_1507,N_1850);
nand U2035 (N_2035,N_1550,N_1023);
or U2036 (N_2036,N_1442,N_1976);
xnor U2037 (N_2037,N_1626,N_1040);
and U2038 (N_2038,N_1698,N_1849);
nor U2039 (N_2039,N_1030,N_1635);
nand U2040 (N_2040,N_1496,N_1375);
and U2041 (N_2041,N_1423,N_1795);
or U2042 (N_2042,N_1282,N_1713);
and U2043 (N_2043,N_1899,N_1430);
nand U2044 (N_2044,N_1693,N_1893);
or U2045 (N_2045,N_1454,N_1600);
nor U2046 (N_2046,N_1515,N_1812);
nand U2047 (N_2047,N_1360,N_1728);
nor U2048 (N_2048,N_1255,N_1853);
nor U2049 (N_2049,N_1053,N_1814);
and U2050 (N_2050,N_1082,N_1163);
nand U2051 (N_2051,N_1060,N_1409);
nor U2052 (N_2052,N_1611,N_1033);
nand U2053 (N_2053,N_1643,N_1601);
xor U2054 (N_2054,N_1111,N_1154);
or U2055 (N_2055,N_1815,N_1944);
nor U2056 (N_2056,N_1838,N_1495);
or U2057 (N_2057,N_1034,N_1435);
nand U2058 (N_2058,N_1731,N_1400);
and U2059 (N_2059,N_1623,N_1472);
and U2060 (N_2060,N_1908,N_1004);
or U2061 (N_2061,N_1558,N_1022);
nor U2062 (N_2062,N_1340,N_1938);
nand U2063 (N_2063,N_1325,N_1821);
nand U2064 (N_2064,N_1128,N_1739);
nor U2065 (N_2065,N_1113,N_1119);
or U2066 (N_2066,N_1544,N_1721);
and U2067 (N_2067,N_1029,N_1065);
or U2068 (N_2068,N_1538,N_1090);
nand U2069 (N_2069,N_1315,N_1797);
nor U2070 (N_2070,N_1367,N_1536);
nor U2071 (N_2071,N_1993,N_1969);
or U2072 (N_2072,N_1493,N_1453);
or U2073 (N_2073,N_1528,N_1615);
nor U2074 (N_2074,N_1054,N_1517);
nor U2075 (N_2075,N_1010,N_1153);
nor U2076 (N_2076,N_1504,N_1366);
and U2077 (N_2077,N_1992,N_1437);
nor U2078 (N_2078,N_1312,N_1559);
nand U2079 (N_2079,N_1051,N_1260);
nand U2080 (N_2080,N_1569,N_1238);
or U2081 (N_2081,N_1578,N_1896);
and U2082 (N_2082,N_1743,N_1416);
or U2083 (N_2083,N_1048,N_1607);
nor U2084 (N_2084,N_1942,N_1657);
nand U2085 (N_2085,N_1963,N_1310);
nor U2086 (N_2086,N_1017,N_1500);
or U2087 (N_2087,N_1251,N_1669);
nor U2088 (N_2088,N_1316,N_1277);
or U2089 (N_2089,N_1725,N_1870);
nor U2090 (N_2090,N_1603,N_1704);
nor U2091 (N_2091,N_1852,N_1291);
nor U2092 (N_2092,N_1363,N_1433);
nor U2093 (N_2093,N_1929,N_1166);
and U2094 (N_2094,N_1820,N_1901);
nor U2095 (N_2095,N_1408,N_1317);
and U2096 (N_2096,N_1461,N_1372);
or U2097 (N_2097,N_1361,N_1983);
and U2098 (N_2098,N_1407,N_1786);
or U2099 (N_2099,N_1359,N_1921);
and U2100 (N_2100,N_1605,N_1125);
or U2101 (N_2101,N_1126,N_1865);
nor U2102 (N_2102,N_1156,N_1912);
and U2103 (N_2103,N_1191,N_1240);
nand U2104 (N_2104,N_1460,N_1221);
and U2105 (N_2105,N_1527,N_1197);
or U2106 (N_2106,N_1140,N_1646);
nor U2107 (N_2107,N_1494,N_1827);
nor U2108 (N_2108,N_1672,N_1279);
or U2109 (N_2109,N_1190,N_1839);
nand U2110 (N_2110,N_1185,N_1529);
nand U2111 (N_2111,N_1782,N_1982);
and U2112 (N_2112,N_1376,N_1665);
xor U2113 (N_2113,N_1371,N_1522);
xor U2114 (N_2114,N_1264,N_1750);
and U2115 (N_2115,N_1478,N_1381);
nand U2116 (N_2116,N_1560,N_1573);
nor U2117 (N_2117,N_1348,N_1724);
nand U2118 (N_2118,N_1087,N_1104);
or U2119 (N_2119,N_1520,N_1862);
or U2120 (N_2120,N_1131,N_1722);
or U2121 (N_2121,N_1293,N_1514);
nor U2122 (N_2122,N_1357,N_1641);
or U2123 (N_2123,N_1592,N_1470);
nand U2124 (N_2124,N_1229,N_1021);
nor U2125 (N_2125,N_1487,N_1160);
or U2126 (N_2126,N_1146,N_1398);
nor U2127 (N_2127,N_1194,N_1327);
and U2128 (N_2128,N_1482,N_1271);
nor U2129 (N_2129,N_1773,N_1799);
or U2130 (N_2130,N_1076,N_1224);
and U2131 (N_2131,N_1099,N_1633);
nor U2132 (N_2132,N_1521,N_1664);
and U2133 (N_2133,N_1876,N_1412);
and U2134 (N_2134,N_1642,N_1692);
and U2135 (N_2135,N_1044,N_1456);
nand U2136 (N_2136,N_1903,N_1723);
nand U2137 (N_2137,N_1364,N_1123);
nor U2138 (N_2138,N_1297,N_1911);
nor U2139 (N_2139,N_1205,N_1792);
and U2140 (N_2140,N_1178,N_1052);
or U2141 (N_2141,N_1513,N_1415);
and U2142 (N_2142,N_1056,N_1823);
nor U2143 (N_2143,N_1241,N_1502);
or U2144 (N_2144,N_1242,N_1562);
nor U2145 (N_2145,N_1427,N_1736);
or U2146 (N_2146,N_1095,N_1628);
and U2147 (N_2147,N_1943,N_1374);
and U2148 (N_2148,N_1037,N_1443);
nor U2149 (N_2149,N_1622,N_1986);
nor U2150 (N_2150,N_1115,N_1660);
nor U2151 (N_2151,N_1822,N_1898);
or U2152 (N_2152,N_1382,N_1287);
nand U2153 (N_2153,N_1776,N_1842);
nor U2154 (N_2154,N_1377,N_1637);
and U2155 (N_2155,N_1038,N_1064);
or U2156 (N_2156,N_1386,N_1695);
xor U2157 (N_2157,N_1777,N_1595);
nor U2158 (N_2158,N_1614,N_1132);
or U2159 (N_2159,N_1226,N_1995);
or U2160 (N_2160,N_1608,N_1345);
or U2161 (N_2161,N_1329,N_1006);
and U2162 (N_2162,N_1213,N_1844);
nor U2163 (N_2163,N_1247,N_1306);
nor U2164 (N_2164,N_1161,N_1223);
nor U2165 (N_2165,N_1709,N_1196);
nand U2166 (N_2166,N_1059,N_1434);
nand U2167 (N_2167,N_1671,N_1855);
nand U2168 (N_2168,N_1066,N_1636);
nor U2169 (N_2169,N_1403,N_1210);
and U2170 (N_2170,N_1429,N_1965);
nor U2171 (N_2171,N_1174,N_1114);
and U2172 (N_2172,N_1183,N_1148);
nand U2173 (N_2173,N_1106,N_1917);
nor U2174 (N_2174,N_1188,N_1867);
and U2175 (N_2175,N_1518,N_1436);
or U2176 (N_2176,N_1511,N_1118);
and U2177 (N_2177,N_1343,N_1871);
nand U2178 (N_2178,N_1589,N_1680);
or U2179 (N_2179,N_1948,N_1545);
nand U2180 (N_2180,N_1549,N_1181);
and U2181 (N_2181,N_1389,N_1768);
and U2182 (N_2182,N_1117,N_1770);
or U2183 (N_2183,N_1729,N_1180);
nand U2184 (N_2184,N_1767,N_1582);
nor U2185 (N_2185,N_1661,N_1077);
and U2186 (N_2186,N_1571,N_1235);
nor U2187 (N_2187,N_1272,N_1845);
xnor U2188 (N_2188,N_1610,N_1445);
and U2189 (N_2189,N_1172,N_1425);
or U2190 (N_2190,N_1328,N_1539);
or U2191 (N_2191,N_1231,N_1024);
or U2192 (N_2192,N_1414,N_1652);
or U2193 (N_2193,N_1694,N_1543);
nand U2194 (N_2194,N_1309,N_1936);
or U2195 (N_2195,N_1874,N_1249);
or U2196 (N_2196,N_1925,N_1772);
or U2197 (N_2197,N_1653,N_1840);
and U2198 (N_2198,N_1499,N_1846);
nand U2199 (N_2199,N_1927,N_1787);
and U2200 (N_2200,N_1552,N_1028);
nor U2201 (N_2201,N_1324,N_1575);
or U2202 (N_2202,N_1110,N_1624);
nand U2203 (N_2203,N_1887,N_1581);
and U2204 (N_2204,N_1955,N_1800);
and U2205 (N_2205,N_1418,N_1627);
nor U2206 (N_2206,N_1204,N_1753);
and U2207 (N_2207,N_1093,N_1365);
nand U2208 (N_2208,N_1085,N_1996);
nand U2209 (N_2209,N_1236,N_1003);
and U2210 (N_2210,N_1791,N_1263);
and U2211 (N_2211,N_1108,N_1141);
nand U2212 (N_2212,N_1506,N_1404);
nor U2213 (N_2213,N_1662,N_1177);
nor U2214 (N_2214,N_1790,N_1138);
nand U2215 (N_2215,N_1199,N_1764);
or U2216 (N_2216,N_1785,N_1308);
nor U2217 (N_2217,N_1831,N_1321);
or U2218 (N_2218,N_1019,N_1266);
nand U2219 (N_2219,N_1318,N_1426);
and U2220 (N_2220,N_1444,N_1286);
and U2221 (N_2221,N_1091,N_1169);
nor U2222 (N_2222,N_1712,N_1143);
or U2223 (N_2223,N_1462,N_1016);
and U2224 (N_2224,N_1219,N_1906);
xnor U2225 (N_2225,N_1042,N_1058);
nand U2226 (N_2226,N_1278,N_1109);
nand U2227 (N_2227,N_1045,N_1155);
or U2228 (N_2228,N_1203,N_1214);
or U2229 (N_2229,N_1913,N_1285);
nand U2230 (N_2230,N_1904,N_1465);
nor U2231 (N_2231,N_1323,N_1977);
and U2232 (N_2232,N_1561,N_1897);
and U2233 (N_2233,N_1352,N_1910);
or U2234 (N_2234,N_1780,N_1253);
or U2235 (N_2235,N_1304,N_1475);
and U2236 (N_2236,N_1001,N_1533);
nand U2237 (N_2237,N_1926,N_1355);
nor U2238 (N_2238,N_1668,N_1710);
or U2239 (N_2239,N_1145,N_1419);
nand U2240 (N_2240,N_1405,N_1159);
and U2241 (N_2241,N_1130,N_1373);
and U2242 (N_2242,N_1902,N_1707);
and U2243 (N_2243,N_1526,N_1701);
and U2244 (N_2244,N_1836,N_1162);
nand U2245 (N_2245,N_1334,N_1075);
nor U2246 (N_2246,N_1069,N_1617);
nand U2247 (N_2247,N_1686,N_1207);
nand U2248 (N_2248,N_1195,N_1974);
and U2249 (N_2249,N_1956,N_1745);
nor U2250 (N_2250,N_1256,N_1892);
nand U2251 (N_2251,N_1638,N_1049);
nor U2252 (N_2252,N_1730,N_1548);
nor U2253 (N_2253,N_1358,N_1858);
nor U2254 (N_2254,N_1301,N_1630);
and U2255 (N_2255,N_1370,N_1656);
nor U2256 (N_2256,N_1498,N_1555);
nand U2257 (N_2257,N_1735,N_1716);
nand U2258 (N_2258,N_1274,N_1947);
nand U2259 (N_2259,N_1448,N_1688);
or U2260 (N_2260,N_1441,N_1677);
nand U2261 (N_2261,N_1305,N_1503);
and U2262 (N_2262,N_1492,N_1258);
or U2263 (N_2263,N_1179,N_1035);
nand U2264 (N_2264,N_1228,N_1998);
and U2265 (N_2265,N_1990,N_1098);
nor U2266 (N_2266,N_1379,N_1347);
nand U2267 (N_2267,N_1742,N_1399);
nor U2268 (N_2268,N_1000,N_1395);
nand U2269 (N_2269,N_1078,N_1525);
and U2270 (N_2270,N_1864,N_1957);
or U2271 (N_2271,N_1477,N_1915);
nand U2272 (N_2272,N_1580,N_1466);
nand U2273 (N_2273,N_1303,N_1083);
or U2274 (N_2274,N_1684,N_1847);
nand U2275 (N_2275,N_1587,N_1625);
nor U2276 (N_2276,N_1127,N_1289);
nor U2277 (N_2277,N_1733,N_1171);
nand U2278 (N_2278,N_1857,N_1951);
nand U2279 (N_2279,N_1164,N_1916);
nand U2280 (N_2280,N_1793,N_1002);
and U2281 (N_2281,N_1509,N_1268);
nand U2282 (N_2282,N_1781,N_1741);
nand U2283 (N_2283,N_1061,N_1121);
or U2284 (N_2284,N_1288,N_1962);
or U2285 (N_2285,N_1009,N_1819);
or U2286 (N_2286,N_1961,N_1647);
nor U2287 (N_2287,N_1655,N_1089);
nor U2288 (N_2288,N_1640,N_1062);
or U2289 (N_2289,N_1939,N_1576);
or U2290 (N_2290,N_1438,N_1598);
and U2291 (N_2291,N_1391,N_1650);
nand U2292 (N_2292,N_1298,N_1719);
nand U2293 (N_2293,N_1572,N_1206);
and U2294 (N_2294,N_1335,N_1393);
nand U2295 (N_2295,N_1342,N_1057);
or U2296 (N_2296,N_1535,N_1201);
nor U2297 (N_2297,N_1516,N_1005);
or U2298 (N_2298,N_1490,N_1332);
nor U2299 (N_2299,N_1973,N_1250);
nor U2300 (N_2300,N_1248,N_1074);
or U2301 (N_2301,N_1072,N_1150);
nand U2302 (N_2302,N_1817,N_1120);
nand U2303 (N_2303,N_1200,N_1008);
nor U2304 (N_2304,N_1100,N_1193);
and U2305 (N_2305,N_1829,N_1914);
or U2306 (N_2306,N_1067,N_1483);
or U2307 (N_2307,N_1854,N_1952);
nor U2308 (N_2308,N_1991,N_1771);
nor U2309 (N_2309,N_1909,N_1720);
nand U2310 (N_2310,N_1046,N_1501);
and U2311 (N_2311,N_1565,N_1937);
or U2312 (N_2312,N_1765,N_1718);
and U2313 (N_2313,N_1041,N_1810);
nor U2314 (N_2314,N_1877,N_1491);
nand U2315 (N_2315,N_1808,N_1568);
nor U2316 (N_2316,N_1873,N_1209);
and U2317 (N_2317,N_1388,N_1063);
nor U2318 (N_2318,N_1889,N_1036);
nand U2319 (N_2319,N_1907,N_1333);
nor U2320 (N_2320,N_1192,N_1967);
nand U2321 (N_2321,N_1806,N_1632);
and U2322 (N_2322,N_1737,N_1620);
or U2323 (N_2323,N_1928,N_1292);
nor U2324 (N_2324,N_1905,N_1330);
nor U2325 (N_2325,N_1594,N_1122);
nor U2326 (N_2326,N_1380,N_1307);
or U2327 (N_2327,N_1758,N_1243);
nor U2328 (N_2328,N_1674,N_1888);
and U2329 (N_2329,N_1168,N_1922);
nor U2330 (N_2330,N_1689,N_1868);
nand U2331 (N_2331,N_1564,N_1681);
nor U2332 (N_2332,N_1281,N_1542);
nand U2333 (N_2333,N_1740,N_1402);
nand U2334 (N_2334,N_1649,N_1167);
and U2335 (N_2335,N_1994,N_1778);
nand U2336 (N_2336,N_1802,N_1530);
xor U2337 (N_2337,N_1619,N_1459);
or U2338 (N_2338,N_1679,N_1834);
or U2339 (N_2339,N_1218,N_1070);
nand U2340 (N_2340,N_1336,N_1284);
xor U2341 (N_2341,N_1988,N_1583);
nor U2342 (N_2342,N_1699,N_1043);
xnor U2343 (N_2343,N_1451,N_1732);
or U2344 (N_2344,N_1612,N_1866);
or U2345 (N_2345,N_1134,N_1270);
xor U2346 (N_2346,N_1659,N_1424);
and U2347 (N_2347,N_1182,N_1863);
nand U2348 (N_2348,N_1985,N_1691);
nor U2349 (N_2349,N_1252,N_1097);
nand U2350 (N_2350,N_1170,N_1246);
and U2351 (N_2351,N_1081,N_1349);
or U2352 (N_2352,N_1966,N_1841);
nand U2353 (N_2353,N_1702,N_1606);
nor U2354 (N_2354,N_1139,N_1884);
nand U2355 (N_2355,N_1577,N_1411);
nand U2356 (N_2356,N_1708,N_1524);
and U2357 (N_2357,N_1455,N_1259);
nor U2358 (N_2358,N_1439,N_1257);
or U2359 (N_2359,N_1356,N_1267);
or U2360 (N_2360,N_1727,N_1798);
or U2361 (N_2361,N_1984,N_1941);
nor U2362 (N_2362,N_1900,N_1476);
nand U2363 (N_2363,N_1924,N_1978);
nand U2364 (N_2364,N_1970,N_1958);
xnor U2365 (N_2365,N_1697,N_1401);
or U2366 (N_2366,N_1591,N_1746);
or U2367 (N_2367,N_1296,N_1705);
nor U2368 (N_2368,N_1757,N_1930);
nand U2369 (N_2369,N_1519,N_1050);
nor U2370 (N_2370,N_1450,N_1397);
or U2371 (N_2371,N_1809,N_1413);
nor U2372 (N_2372,N_1920,N_1295);
nor U2373 (N_2373,N_1208,N_1923);
xnor U2374 (N_2374,N_1796,N_1351);
nand U2375 (N_2375,N_1621,N_1173);
and U2376 (N_2376,N_1748,N_1566);
or U2377 (N_2377,N_1480,N_1616);
nand U2378 (N_2378,N_1015,N_1934);
or U2379 (N_2379,N_1651,N_1546);
and U2380 (N_2380,N_1457,N_1987);
nor U2381 (N_2381,N_1497,N_1368);
or U2382 (N_2382,N_1755,N_1189);
nand U2383 (N_2383,N_1599,N_1759);
or U2384 (N_2384,N_1676,N_1711);
nand U2385 (N_2385,N_1239,N_1387);
and U2386 (N_2386,N_1648,N_1828);
and U2387 (N_2387,N_1604,N_1157);
or U2388 (N_2388,N_1999,N_1225);
nor U2389 (N_2389,N_1803,N_1754);
xor U2390 (N_2390,N_1890,N_1683);
xnor U2391 (N_2391,N_1432,N_1473);
nor U2392 (N_2392,N_1440,N_1392);
and U2393 (N_2393,N_1354,N_1563);
nor U2394 (N_2394,N_1953,N_1752);
nor U2395 (N_2395,N_1639,N_1202);
or U2396 (N_2396,N_1675,N_1326);
nand U2397 (N_2397,N_1950,N_1678);
nand U2398 (N_2398,N_1715,N_1079);
nand U2399 (N_2399,N_1322,N_1149);
nor U2400 (N_2400,N_1825,N_1112);
nor U2401 (N_2401,N_1458,N_1158);
and U2402 (N_2402,N_1861,N_1234);
nor U2403 (N_2403,N_1133,N_1886);
and U2404 (N_2404,N_1744,N_1135);
or U2405 (N_2405,N_1055,N_1860);
nand U2406 (N_2406,N_1151,N_1756);
and U2407 (N_2407,N_1446,N_1020);
or U2408 (N_2408,N_1980,N_1851);
nand U2409 (N_2409,N_1894,N_1654);
nor U2410 (N_2410,N_1510,N_1262);
or U2411 (N_2411,N_1467,N_1230);
and U2412 (N_2412,N_1816,N_1734);
and U2413 (N_2413,N_1233,N_1590);
nand U2414 (N_2414,N_1137,N_1766);
nand U2415 (N_2415,N_1703,N_1631);
nand U2416 (N_2416,N_1895,N_1644);
nor U2417 (N_2417,N_1872,N_1129);
or U2418 (N_2418,N_1102,N_1975);
and U2419 (N_2419,N_1774,N_1468);
nor U2420 (N_2420,N_1198,N_1186);
or U2421 (N_2421,N_1717,N_1463);
or U2422 (N_2422,N_1751,N_1484);
or U2423 (N_2423,N_1738,N_1879);
nand U2424 (N_2424,N_1673,N_1593);
nor U2425 (N_2425,N_1690,N_1556);
or U2426 (N_2426,N_1749,N_1856);
nand U2427 (N_2427,N_1384,N_1142);
nor U2428 (N_2428,N_1833,N_1394);
and U2429 (N_2429,N_1212,N_1618);
nor U2430 (N_2430,N_1554,N_1486);
or U2431 (N_2431,N_1726,N_1918);
and U2432 (N_2432,N_1222,N_1788);
or U2433 (N_2433,N_1645,N_1613);
nor U2434 (N_2434,N_1237,N_1547);
and U2435 (N_2435,N_1585,N_1290);
nor U2436 (N_2436,N_1931,N_1187);
nand U2437 (N_2437,N_1011,N_1584);
and U2438 (N_2438,N_1935,N_1835);
and U2439 (N_2439,N_1216,N_1068);
nand U2440 (N_2440,N_1574,N_1667);
and U2441 (N_2441,N_1406,N_1997);
nor U2442 (N_2442,N_1396,N_1512);
and U2443 (N_2443,N_1882,N_1878);
nand U2444 (N_2444,N_1471,N_1481);
and U2445 (N_2445,N_1972,N_1474);
nor U2446 (N_2446,N_1505,N_1789);
and U2447 (N_2447,N_1531,N_1875);
nand U2448 (N_2448,N_1232,N_1714);
nand U2449 (N_2449,N_1344,N_1244);
nand U2450 (N_2450,N_1086,N_1586);
or U2451 (N_2451,N_1813,N_1489);
nor U2452 (N_2452,N_1300,N_1946);
nand U2453 (N_2453,N_1848,N_1215);
or U2454 (N_2454,N_1276,N_1687);
or U2455 (N_2455,N_1989,N_1245);
xor U2456 (N_2456,N_1832,N_1784);
or U2457 (N_2457,N_1932,N_1567);
or U2458 (N_2458,N_1532,N_1824);
or U2459 (N_2459,N_1945,N_1013);
and U2460 (N_2460,N_1410,N_1254);
nor U2461 (N_2461,N_1891,N_1088);
or U2462 (N_2462,N_1769,N_1488);
nor U2463 (N_2463,N_1073,N_1869);
and U2464 (N_2464,N_1954,N_1706);
nor U2465 (N_2465,N_1362,N_1557);
nor U2466 (N_2466,N_1390,N_1175);
nand U2467 (N_2467,N_1449,N_1979);
and U2468 (N_2468,N_1319,N_1431);
nor U2469 (N_2469,N_1971,N_1346);
nand U2470 (N_2470,N_1261,N_1859);
nand U2471 (N_2471,N_1479,N_1570);
and U2472 (N_2472,N_1843,N_1107);
nor U2473 (N_2473,N_1320,N_1280);
or U2474 (N_2474,N_1837,N_1369);
nor U2475 (N_2475,N_1269,N_1880);
nand U2476 (N_2476,N_1508,N_1485);
or U2477 (N_2477,N_1949,N_1540);
or U2478 (N_2478,N_1634,N_1658);
or U2479 (N_2479,N_1227,N_1818);
nor U2480 (N_2480,N_1176,N_1541);
and U2481 (N_2481,N_1341,N_1670);
nand U2482 (N_2482,N_1422,N_1537);
nand U2483 (N_2483,N_1144,N_1807);
nand U2484 (N_2484,N_1579,N_1760);
and U2485 (N_2485,N_1609,N_1666);
nor U2486 (N_2486,N_1452,N_1101);
or U2487 (N_2487,N_1968,N_1933);
or U2488 (N_2488,N_1885,N_1447);
and U2489 (N_2489,N_1417,N_1883);
or U2490 (N_2490,N_1220,N_1096);
nor U2491 (N_2491,N_1805,N_1378);
nor U2492 (N_2492,N_1353,N_1981);
xor U2493 (N_2493,N_1283,N_1960);
or U2494 (N_2494,N_1092,N_1881);
or U2495 (N_2495,N_1464,N_1629);
or U2496 (N_2496,N_1012,N_1027);
nor U2497 (N_2497,N_1084,N_1383);
or U2498 (N_2498,N_1165,N_1523);
and U2499 (N_2499,N_1094,N_1551);
nand U2500 (N_2500,N_1949,N_1467);
or U2501 (N_2501,N_1320,N_1702);
and U2502 (N_2502,N_1232,N_1066);
nand U2503 (N_2503,N_1302,N_1904);
nand U2504 (N_2504,N_1594,N_1526);
nor U2505 (N_2505,N_1109,N_1091);
or U2506 (N_2506,N_1911,N_1782);
nor U2507 (N_2507,N_1028,N_1666);
or U2508 (N_2508,N_1947,N_1324);
or U2509 (N_2509,N_1141,N_1583);
nor U2510 (N_2510,N_1929,N_1476);
nand U2511 (N_2511,N_1490,N_1493);
or U2512 (N_2512,N_1875,N_1342);
or U2513 (N_2513,N_1755,N_1577);
nand U2514 (N_2514,N_1095,N_1156);
or U2515 (N_2515,N_1738,N_1561);
nor U2516 (N_2516,N_1538,N_1165);
nor U2517 (N_2517,N_1390,N_1494);
nand U2518 (N_2518,N_1691,N_1802);
and U2519 (N_2519,N_1389,N_1671);
nand U2520 (N_2520,N_1988,N_1464);
and U2521 (N_2521,N_1559,N_1391);
nor U2522 (N_2522,N_1413,N_1032);
nor U2523 (N_2523,N_1205,N_1932);
nand U2524 (N_2524,N_1557,N_1120);
and U2525 (N_2525,N_1311,N_1062);
nor U2526 (N_2526,N_1580,N_1234);
nand U2527 (N_2527,N_1683,N_1378);
nand U2528 (N_2528,N_1521,N_1997);
nor U2529 (N_2529,N_1618,N_1344);
nor U2530 (N_2530,N_1097,N_1899);
nor U2531 (N_2531,N_1636,N_1576);
xnor U2532 (N_2532,N_1346,N_1852);
nor U2533 (N_2533,N_1498,N_1902);
xnor U2534 (N_2534,N_1410,N_1692);
nand U2535 (N_2535,N_1535,N_1661);
or U2536 (N_2536,N_1549,N_1286);
nand U2537 (N_2537,N_1615,N_1896);
nor U2538 (N_2538,N_1964,N_1480);
or U2539 (N_2539,N_1248,N_1563);
nand U2540 (N_2540,N_1917,N_1337);
or U2541 (N_2541,N_1982,N_1712);
nand U2542 (N_2542,N_1415,N_1898);
or U2543 (N_2543,N_1449,N_1524);
nor U2544 (N_2544,N_1611,N_1195);
nor U2545 (N_2545,N_1378,N_1653);
nand U2546 (N_2546,N_1734,N_1912);
nand U2547 (N_2547,N_1586,N_1795);
nor U2548 (N_2548,N_1177,N_1999);
nand U2549 (N_2549,N_1203,N_1048);
and U2550 (N_2550,N_1490,N_1239);
nor U2551 (N_2551,N_1483,N_1697);
nand U2552 (N_2552,N_1624,N_1149);
and U2553 (N_2553,N_1640,N_1812);
and U2554 (N_2554,N_1060,N_1414);
and U2555 (N_2555,N_1376,N_1389);
nand U2556 (N_2556,N_1320,N_1093);
xnor U2557 (N_2557,N_1108,N_1529);
nor U2558 (N_2558,N_1422,N_1645);
nand U2559 (N_2559,N_1653,N_1153);
nor U2560 (N_2560,N_1330,N_1800);
nand U2561 (N_2561,N_1180,N_1924);
or U2562 (N_2562,N_1080,N_1130);
or U2563 (N_2563,N_1631,N_1270);
or U2564 (N_2564,N_1662,N_1991);
and U2565 (N_2565,N_1524,N_1722);
and U2566 (N_2566,N_1714,N_1733);
and U2567 (N_2567,N_1786,N_1176);
xor U2568 (N_2568,N_1124,N_1142);
xor U2569 (N_2569,N_1869,N_1248);
or U2570 (N_2570,N_1975,N_1320);
nand U2571 (N_2571,N_1995,N_1051);
or U2572 (N_2572,N_1331,N_1471);
and U2573 (N_2573,N_1163,N_1625);
and U2574 (N_2574,N_1650,N_1054);
nand U2575 (N_2575,N_1139,N_1720);
and U2576 (N_2576,N_1594,N_1538);
xnor U2577 (N_2577,N_1682,N_1704);
nor U2578 (N_2578,N_1516,N_1244);
nor U2579 (N_2579,N_1964,N_1438);
or U2580 (N_2580,N_1710,N_1744);
and U2581 (N_2581,N_1977,N_1442);
and U2582 (N_2582,N_1769,N_1584);
or U2583 (N_2583,N_1673,N_1904);
nand U2584 (N_2584,N_1149,N_1593);
or U2585 (N_2585,N_1747,N_1421);
nand U2586 (N_2586,N_1874,N_1027);
nor U2587 (N_2587,N_1069,N_1683);
xor U2588 (N_2588,N_1027,N_1753);
nor U2589 (N_2589,N_1781,N_1785);
or U2590 (N_2590,N_1313,N_1589);
nor U2591 (N_2591,N_1678,N_1992);
or U2592 (N_2592,N_1580,N_1261);
or U2593 (N_2593,N_1556,N_1679);
or U2594 (N_2594,N_1078,N_1959);
or U2595 (N_2595,N_1444,N_1526);
or U2596 (N_2596,N_1952,N_1650);
nand U2597 (N_2597,N_1879,N_1019);
nor U2598 (N_2598,N_1646,N_1488);
or U2599 (N_2599,N_1423,N_1858);
or U2600 (N_2600,N_1455,N_1384);
nand U2601 (N_2601,N_1736,N_1101);
or U2602 (N_2602,N_1603,N_1558);
or U2603 (N_2603,N_1259,N_1374);
nor U2604 (N_2604,N_1644,N_1003);
nor U2605 (N_2605,N_1290,N_1940);
nor U2606 (N_2606,N_1809,N_1396);
nand U2607 (N_2607,N_1193,N_1649);
nor U2608 (N_2608,N_1049,N_1407);
or U2609 (N_2609,N_1055,N_1578);
and U2610 (N_2610,N_1780,N_1029);
and U2611 (N_2611,N_1976,N_1361);
or U2612 (N_2612,N_1050,N_1925);
xor U2613 (N_2613,N_1217,N_1266);
nand U2614 (N_2614,N_1256,N_1811);
nor U2615 (N_2615,N_1892,N_1797);
or U2616 (N_2616,N_1196,N_1147);
or U2617 (N_2617,N_1432,N_1923);
nor U2618 (N_2618,N_1089,N_1829);
and U2619 (N_2619,N_1232,N_1506);
nand U2620 (N_2620,N_1977,N_1718);
nand U2621 (N_2621,N_1569,N_1150);
or U2622 (N_2622,N_1879,N_1787);
and U2623 (N_2623,N_1866,N_1723);
nor U2624 (N_2624,N_1454,N_1312);
or U2625 (N_2625,N_1492,N_1823);
nor U2626 (N_2626,N_1298,N_1439);
nand U2627 (N_2627,N_1367,N_1776);
nor U2628 (N_2628,N_1865,N_1667);
nor U2629 (N_2629,N_1262,N_1249);
and U2630 (N_2630,N_1208,N_1823);
nor U2631 (N_2631,N_1196,N_1650);
nand U2632 (N_2632,N_1115,N_1768);
nand U2633 (N_2633,N_1049,N_1156);
and U2634 (N_2634,N_1472,N_1721);
nor U2635 (N_2635,N_1963,N_1308);
nand U2636 (N_2636,N_1839,N_1183);
or U2637 (N_2637,N_1107,N_1667);
or U2638 (N_2638,N_1024,N_1642);
nor U2639 (N_2639,N_1593,N_1979);
nand U2640 (N_2640,N_1036,N_1969);
nor U2641 (N_2641,N_1167,N_1016);
xnor U2642 (N_2642,N_1161,N_1688);
nand U2643 (N_2643,N_1805,N_1108);
and U2644 (N_2644,N_1123,N_1645);
or U2645 (N_2645,N_1912,N_1115);
or U2646 (N_2646,N_1599,N_1163);
xnor U2647 (N_2647,N_1509,N_1434);
nand U2648 (N_2648,N_1246,N_1134);
and U2649 (N_2649,N_1776,N_1894);
and U2650 (N_2650,N_1325,N_1160);
or U2651 (N_2651,N_1806,N_1453);
nand U2652 (N_2652,N_1201,N_1264);
nor U2653 (N_2653,N_1337,N_1226);
and U2654 (N_2654,N_1717,N_1575);
nand U2655 (N_2655,N_1447,N_1040);
nand U2656 (N_2656,N_1679,N_1753);
nand U2657 (N_2657,N_1467,N_1080);
nand U2658 (N_2658,N_1030,N_1993);
nand U2659 (N_2659,N_1752,N_1083);
nor U2660 (N_2660,N_1201,N_1008);
nand U2661 (N_2661,N_1466,N_1759);
xor U2662 (N_2662,N_1647,N_1903);
nand U2663 (N_2663,N_1884,N_1336);
and U2664 (N_2664,N_1530,N_1676);
nor U2665 (N_2665,N_1054,N_1990);
nor U2666 (N_2666,N_1840,N_1579);
or U2667 (N_2667,N_1237,N_1000);
nor U2668 (N_2668,N_1936,N_1288);
or U2669 (N_2669,N_1073,N_1130);
or U2670 (N_2670,N_1277,N_1514);
or U2671 (N_2671,N_1241,N_1692);
nand U2672 (N_2672,N_1053,N_1971);
or U2673 (N_2673,N_1009,N_1270);
nor U2674 (N_2674,N_1127,N_1250);
and U2675 (N_2675,N_1737,N_1970);
nand U2676 (N_2676,N_1705,N_1777);
or U2677 (N_2677,N_1980,N_1913);
or U2678 (N_2678,N_1728,N_1049);
nor U2679 (N_2679,N_1420,N_1766);
nand U2680 (N_2680,N_1737,N_1649);
and U2681 (N_2681,N_1613,N_1993);
nor U2682 (N_2682,N_1599,N_1042);
or U2683 (N_2683,N_1218,N_1738);
nor U2684 (N_2684,N_1346,N_1857);
and U2685 (N_2685,N_1005,N_1654);
or U2686 (N_2686,N_1479,N_1214);
nand U2687 (N_2687,N_1954,N_1043);
nand U2688 (N_2688,N_1453,N_1376);
nor U2689 (N_2689,N_1151,N_1891);
nand U2690 (N_2690,N_1708,N_1195);
or U2691 (N_2691,N_1982,N_1965);
or U2692 (N_2692,N_1390,N_1825);
nand U2693 (N_2693,N_1737,N_1240);
nor U2694 (N_2694,N_1058,N_1554);
and U2695 (N_2695,N_1148,N_1773);
and U2696 (N_2696,N_1101,N_1956);
and U2697 (N_2697,N_1209,N_1099);
nand U2698 (N_2698,N_1358,N_1307);
or U2699 (N_2699,N_1529,N_1110);
nor U2700 (N_2700,N_1408,N_1415);
and U2701 (N_2701,N_1428,N_1820);
or U2702 (N_2702,N_1532,N_1450);
or U2703 (N_2703,N_1925,N_1461);
xor U2704 (N_2704,N_1926,N_1806);
or U2705 (N_2705,N_1418,N_1870);
nor U2706 (N_2706,N_1273,N_1391);
nand U2707 (N_2707,N_1566,N_1490);
and U2708 (N_2708,N_1559,N_1520);
or U2709 (N_2709,N_1552,N_1748);
and U2710 (N_2710,N_1976,N_1994);
or U2711 (N_2711,N_1927,N_1347);
nor U2712 (N_2712,N_1872,N_1679);
nor U2713 (N_2713,N_1389,N_1658);
nand U2714 (N_2714,N_1403,N_1263);
and U2715 (N_2715,N_1775,N_1912);
nand U2716 (N_2716,N_1239,N_1174);
nor U2717 (N_2717,N_1807,N_1699);
nand U2718 (N_2718,N_1326,N_1377);
and U2719 (N_2719,N_1173,N_1207);
or U2720 (N_2720,N_1723,N_1755);
xor U2721 (N_2721,N_1641,N_1108);
and U2722 (N_2722,N_1904,N_1205);
nor U2723 (N_2723,N_1314,N_1840);
and U2724 (N_2724,N_1454,N_1163);
nor U2725 (N_2725,N_1373,N_1304);
and U2726 (N_2726,N_1062,N_1609);
nor U2727 (N_2727,N_1797,N_1538);
or U2728 (N_2728,N_1529,N_1062);
nor U2729 (N_2729,N_1980,N_1537);
or U2730 (N_2730,N_1649,N_1945);
or U2731 (N_2731,N_1167,N_1921);
nand U2732 (N_2732,N_1506,N_1829);
and U2733 (N_2733,N_1677,N_1290);
or U2734 (N_2734,N_1744,N_1252);
or U2735 (N_2735,N_1603,N_1573);
or U2736 (N_2736,N_1391,N_1657);
or U2737 (N_2737,N_1736,N_1939);
nand U2738 (N_2738,N_1557,N_1300);
nand U2739 (N_2739,N_1661,N_1488);
nand U2740 (N_2740,N_1981,N_1860);
nand U2741 (N_2741,N_1844,N_1611);
nor U2742 (N_2742,N_1891,N_1907);
nand U2743 (N_2743,N_1363,N_1717);
nor U2744 (N_2744,N_1331,N_1315);
or U2745 (N_2745,N_1984,N_1257);
nand U2746 (N_2746,N_1326,N_1712);
or U2747 (N_2747,N_1116,N_1487);
nor U2748 (N_2748,N_1480,N_1574);
nand U2749 (N_2749,N_1482,N_1818);
and U2750 (N_2750,N_1404,N_1332);
or U2751 (N_2751,N_1163,N_1267);
xnor U2752 (N_2752,N_1593,N_1190);
and U2753 (N_2753,N_1852,N_1858);
or U2754 (N_2754,N_1297,N_1377);
or U2755 (N_2755,N_1652,N_1242);
nor U2756 (N_2756,N_1331,N_1027);
nor U2757 (N_2757,N_1509,N_1815);
nor U2758 (N_2758,N_1281,N_1968);
nand U2759 (N_2759,N_1322,N_1770);
and U2760 (N_2760,N_1598,N_1061);
xnor U2761 (N_2761,N_1203,N_1897);
and U2762 (N_2762,N_1325,N_1828);
nor U2763 (N_2763,N_1056,N_1646);
nor U2764 (N_2764,N_1366,N_1267);
nand U2765 (N_2765,N_1282,N_1808);
nor U2766 (N_2766,N_1159,N_1176);
or U2767 (N_2767,N_1138,N_1123);
nand U2768 (N_2768,N_1469,N_1918);
or U2769 (N_2769,N_1449,N_1048);
nand U2770 (N_2770,N_1197,N_1232);
nor U2771 (N_2771,N_1873,N_1216);
nor U2772 (N_2772,N_1373,N_1905);
or U2773 (N_2773,N_1615,N_1627);
or U2774 (N_2774,N_1957,N_1177);
nand U2775 (N_2775,N_1016,N_1739);
nand U2776 (N_2776,N_1460,N_1110);
and U2777 (N_2777,N_1151,N_1330);
and U2778 (N_2778,N_1414,N_1359);
and U2779 (N_2779,N_1158,N_1064);
or U2780 (N_2780,N_1469,N_1607);
or U2781 (N_2781,N_1788,N_1969);
nand U2782 (N_2782,N_1032,N_1060);
nor U2783 (N_2783,N_1620,N_1100);
nand U2784 (N_2784,N_1687,N_1391);
nand U2785 (N_2785,N_1938,N_1716);
nand U2786 (N_2786,N_1937,N_1944);
nor U2787 (N_2787,N_1335,N_1809);
and U2788 (N_2788,N_1985,N_1807);
or U2789 (N_2789,N_1056,N_1001);
nand U2790 (N_2790,N_1417,N_1552);
nand U2791 (N_2791,N_1353,N_1208);
or U2792 (N_2792,N_1513,N_1256);
nand U2793 (N_2793,N_1236,N_1978);
or U2794 (N_2794,N_1063,N_1243);
and U2795 (N_2795,N_1876,N_1572);
nor U2796 (N_2796,N_1862,N_1668);
nor U2797 (N_2797,N_1222,N_1589);
nand U2798 (N_2798,N_1272,N_1701);
or U2799 (N_2799,N_1135,N_1717);
or U2800 (N_2800,N_1232,N_1392);
or U2801 (N_2801,N_1329,N_1445);
nand U2802 (N_2802,N_1212,N_1287);
nor U2803 (N_2803,N_1819,N_1098);
nor U2804 (N_2804,N_1867,N_1178);
nand U2805 (N_2805,N_1501,N_1953);
or U2806 (N_2806,N_1910,N_1881);
nand U2807 (N_2807,N_1471,N_1656);
nor U2808 (N_2808,N_1945,N_1812);
nand U2809 (N_2809,N_1322,N_1592);
nand U2810 (N_2810,N_1874,N_1509);
or U2811 (N_2811,N_1101,N_1587);
nor U2812 (N_2812,N_1471,N_1812);
nor U2813 (N_2813,N_1365,N_1298);
nor U2814 (N_2814,N_1377,N_1237);
or U2815 (N_2815,N_1429,N_1716);
nand U2816 (N_2816,N_1744,N_1756);
or U2817 (N_2817,N_1152,N_1645);
or U2818 (N_2818,N_1018,N_1463);
nor U2819 (N_2819,N_1689,N_1076);
nor U2820 (N_2820,N_1250,N_1013);
nor U2821 (N_2821,N_1882,N_1072);
nor U2822 (N_2822,N_1397,N_1336);
and U2823 (N_2823,N_1560,N_1732);
nand U2824 (N_2824,N_1994,N_1526);
and U2825 (N_2825,N_1138,N_1878);
xor U2826 (N_2826,N_1599,N_1591);
nand U2827 (N_2827,N_1170,N_1816);
and U2828 (N_2828,N_1648,N_1694);
and U2829 (N_2829,N_1573,N_1060);
nor U2830 (N_2830,N_1714,N_1429);
nor U2831 (N_2831,N_1137,N_1448);
and U2832 (N_2832,N_1924,N_1666);
nor U2833 (N_2833,N_1927,N_1813);
or U2834 (N_2834,N_1180,N_1946);
or U2835 (N_2835,N_1317,N_1395);
or U2836 (N_2836,N_1792,N_1811);
and U2837 (N_2837,N_1250,N_1918);
nor U2838 (N_2838,N_1466,N_1635);
and U2839 (N_2839,N_1237,N_1636);
and U2840 (N_2840,N_1283,N_1102);
nor U2841 (N_2841,N_1255,N_1206);
nor U2842 (N_2842,N_1368,N_1865);
nand U2843 (N_2843,N_1082,N_1255);
nor U2844 (N_2844,N_1603,N_1671);
or U2845 (N_2845,N_1563,N_1241);
and U2846 (N_2846,N_1876,N_1901);
nand U2847 (N_2847,N_1335,N_1717);
and U2848 (N_2848,N_1359,N_1607);
nor U2849 (N_2849,N_1541,N_1044);
or U2850 (N_2850,N_1190,N_1188);
nand U2851 (N_2851,N_1815,N_1785);
nor U2852 (N_2852,N_1681,N_1617);
or U2853 (N_2853,N_1618,N_1678);
or U2854 (N_2854,N_1141,N_1462);
nand U2855 (N_2855,N_1521,N_1247);
nand U2856 (N_2856,N_1278,N_1560);
or U2857 (N_2857,N_1458,N_1833);
and U2858 (N_2858,N_1654,N_1786);
and U2859 (N_2859,N_1676,N_1786);
nor U2860 (N_2860,N_1707,N_1246);
nand U2861 (N_2861,N_1300,N_1043);
and U2862 (N_2862,N_1116,N_1753);
and U2863 (N_2863,N_1490,N_1485);
and U2864 (N_2864,N_1630,N_1307);
or U2865 (N_2865,N_1871,N_1512);
or U2866 (N_2866,N_1333,N_1763);
and U2867 (N_2867,N_1670,N_1308);
and U2868 (N_2868,N_1122,N_1306);
nand U2869 (N_2869,N_1181,N_1324);
or U2870 (N_2870,N_1471,N_1168);
and U2871 (N_2871,N_1948,N_1205);
nor U2872 (N_2872,N_1963,N_1030);
or U2873 (N_2873,N_1821,N_1372);
nand U2874 (N_2874,N_1507,N_1242);
nor U2875 (N_2875,N_1794,N_1474);
and U2876 (N_2876,N_1428,N_1474);
nand U2877 (N_2877,N_1573,N_1955);
and U2878 (N_2878,N_1320,N_1069);
and U2879 (N_2879,N_1122,N_1765);
nor U2880 (N_2880,N_1950,N_1964);
and U2881 (N_2881,N_1406,N_1811);
and U2882 (N_2882,N_1631,N_1353);
and U2883 (N_2883,N_1303,N_1933);
nand U2884 (N_2884,N_1525,N_1313);
nand U2885 (N_2885,N_1763,N_1575);
nor U2886 (N_2886,N_1031,N_1200);
and U2887 (N_2887,N_1941,N_1311);
and U2888 (N_2888,N_1882,N_1489);
nor U2889 (N_2889,N_1656,N_1031);
or U2890 (N_2890,N_1929,N_1553);
nand U2891 (N_2891,N_1519,N_1855);
nand U2892 (N_2892,N_1519,N_1719);
or U2893 (N_2893,N_1343,N_1727);
nor U2894 (N_2894,N_1812,N_1583);
nand U2895 (N_2895,N_1484,N_1002);
and U2896 (N_2896,N_1646,N_1926);
nor U2897 (N_2897,N_1471,N_1703);
and U2898 (N_2898,N_1047,N_1255);
or U2899 (N_2899,N_1575,N_1637);
and U2900 (N_2900,N_1949,N_1198);
nand U2901 (N_2901,N_1723,N_1722);
nand U2902 (N_2902,N_1293,N_1046);
or U2903 (N_2903,N_1376,N_1200);
nand U2904 (N_2904,N_1795,N_1193);
or U2905 (N_2905,N_1437,N_1639);
nand U2906 (N_2906,N_1986,N_1700);
or U2907 (N_2907,N_1238,N_1098);
nor U2908 (N_2908,N_1667,N_1748);
nand U2909 (N_2909,N_1033,N_1282);
or U2910 (N_2910,N_1641,N_1782);
nor U2911 (N_2911,N_1743,N_1427);
and U2912 (N_2912,N_1343,N_1840);
xor U2913 (N_2913,N_1939,N_1013);
nor U2914 (N_2914,N_1144,N_1735);
and U2915 (N_2915,N_1074,N_1539);
nand U2916 (N_2916,N_1828,N_1580);
nor U2917 (N_2917,N_1689,N_1578);
nor U2918 (N_2918,N_1215,N_1239);
and U2919 (N_2919,N_1011,N_1815);
or U2920 (N_2920,N_1200,N_1577);
and U2921 (N_2921,N_1329,N_1210);
and U2922 (N_2922,N_1071,N_1810);
and U2923 (N_2923,N_1435,N_1172);
and U2924 (N_2924,N_1081,N_1974);
nand U2925 (N_2925,N_1033,N_1960);
and U2926 (N_2926,N_1501,N_1697);
and U2927 (N_2927,N_1809,N_1123);
and U2928 (N_2928,N_1026,N_1822);
or U2929 (N_2929,N_1570,N_1612);
and U2930 (N_2930,N_1852,N_1819);
and U2931 (N_2931,N_1900,N_1926);
or U2932 (N_2932,N_1299,N_1586);
and U2933 (N_2933,N_1025,N_1275);
or U2934 (N_2934,N_1697,N_1522);
nor U2935 (N_2935,N_1225,N_1506);
nor U2936 (N_2936,N_1707,N_1489);
nand U2937 (N_2937,N_1424,N_1225);
and U2938 (N_2938,N_1403,N_1343);
or U2939 (N_2939,N_1908,N_1867);
nand U2940 (N_2940,N_1916,N_1357);
nand U2941 (N_2941,N_1046,N_1267);
nor U2942 (N_2942,N_1272,N_1582);
nor U2943 (N_2943,N_1024,N_1632);
nor U2944 (N_2944,N_1859,N_1809);
or U2945 (N_2945,N_1664,N_1709);
or U2946 (N_2946,N_1330,N_1123);
and U2947 (N_2947,N_1212,N_1843);
nor U2948 (N_2948,N_1003,N_1924);
nand U2949 (N_2949,N_1877,N_1766);
nor U2950 (N_2950,N_1883,N_1355);
and U2951 (N_2951,N_1437,N_1933);
or U2952 (N_2952,N_1557,N_1690);
nor U2953 (N_2953,N_1089,N_1363);
nand U2954 (N_2954,N_1700,N_1140);
and U2955 (N_2955,N_1110,N_1721);
or U2956 (N_2956,N_1272,N_1663);
nand U2957 (N_2957,N_1096,N_1338);
nand U2958 (N_2958,N_1765,N_1228);
or U2959 (N_2959,N_1884,N_1934);
nand U2960 (N_2960,N_1470,N_1512);
and U2961 (N_2961,N_1754,N_1536);
nor U2962 (N_2962,N_1418,N_1826);
nand U2963 (N_2963,N_1186,N_1146);
nor U2964 (N_2964,N_1769,N_1929);
nand U2965 (N_2965,N_1322,N_1562);
nand U2966 (N_2966,N_1167,N_1056);
nand U2967 (N_2967,N_1550,N_1720);
or U2968 (N_2968,N_1360,N_1961);
and U2969 (N_2969,N_1653,N_1181);
nor U2970 (N_2970,N_1921,N_1203);
or U2971 (N_2971,N_1514,N_1398);
nor U2972 (N_2972,N_1024,N_1022);
nand U2973 (N_2973,N_1243,N_1062);
xnor U2974 (N_2974,N_1869,N_1572);
nor U2975 (N_2975,N_1113,N_1282);
nor U2976 (N_2976,N_1526,N_1684);
or U2977 (N_2977,N_1075,N_1514);
or U2978 (N_2978,N_1092,N_1013);
xnor U2979 (N_2979,N_1138,N_1187);
or U2980 (N_2980,N_1447,N_1451);
nand U2981 (N_2981,N_1036,N_1327);
nor U2982 (N_2982,N_1056,N_1608);
or U2983 (N_2983,N_1577,N_1419);
and U2984 (N_2984,N_1505,N_1933);
nand U2985 (N_2985,N_1188,N_1573);
nor U2986 (N_2986,N_1153,N_1767);
nor U2987 (N_2987,N_1354,N_1411);
nand U2988 (N_2988,N_1736,N_1244);
nor U2989 (N_2989,N_1971,N_1186);
nor U2990 (N_2990,N_1231,N_1968);
or U2991 (N_2991,N_1397,N_1987);
nor U2992 (N_2992,N_1563,N_1870);
nor U2993 (N_2993,N_1209,N_1376);
nand U2994 (N_2994,N_1152,N_1515);
nor U2995 (N_2995,N_1193,N_1776);
and U2996 (N_2996,N_1827,N_1931);
nand U2997 (N_2997,N_1254,N_1426);
nand U2998 (N_2998,N_1462,N_1426);
or U2999 (N_2999,N_1279,N_1496);
nor U3000 (N_3000,N_2084,N_2904);
or U3001 (N_3001,N_2080,N_2970);
nand U3002 (N_3002,N_2065,N_2640);
or U3003 (N_3003,N_2418,N_2400);
nor U3004 (N_3004,N_2206,N_2965);
nor U3005 (N_3005,N_2258,N_2911);
nand U3006 (N_3006,N_2380,N_2518);
or U3007 (N_3007,N_2072,N_2044);
and U3008 (N_3008,N_2053,N_2057);
and U3009 (N_3009,N_2256,N_2980);
or U3010 (N_3010,N_2552,N_2601);
nor U3011 (N_3011,N_2990,N_2560);
or U3012 (N_3012,N_2326,N_2690);
nor U3013 (N_3013,N_2104,N_2567);
and U3014 (N_3014,N_2996,N_2986);
nand U3015 (N_3015,N_2482,N_2320);
nand U3016 (N_3016,N_2011,N_2271);
nand U3017 (N_3017,N_2670,N_2770);
or U3018 (N_3018,N_2162,N_2479);
or U3019 (N_3019,N_2116,N_2173);
nor U3020 (N_3020,N_2260,N_2696);
nand U3021 (N_3021,N_2950,N_2976);
or U3022 (N_3022,N_2780,N_2901);
nor U3023 (N_3023,N_2179,N_2798);
xor U3024 (N_3024,N_2815,N_2637);
and U3025 (N_3025,N_2630,N_2753);
xnor U3026 (N_3026,N_2559,N_2773);
nand U3027 (N_3027,N_2813,N_2296);
or U3028 (N_3028,N_2376,N_2136);
nand U3029 (N_3029,N_2349,N_2477);
nand U3030 (N_3030,N_2193,N_2681);
and U3031 (N_3031,N_2277,N_2828);
and U3032 (N_3032,N_2489,N_2473);
or U3033 (N_3033,N_2615,N_2997);
or U3034 (N_3034,N_2314,N_2267);
or U3035 (N_3035,N_2792,N_2283);
and U3036 (N_3036,N_2833,N_2379);
nor U3037 (N_3037,N_2840,N_2947);
xnor U3038 (N_3038,N_2705,N_2194);
and U3039 (N_3039,N_2437,N_2507);
nor U3040 (N_3040,N_2703,N_2159);
or U3041 (N_3041,N_2654,N_2971);
nor U3042 (N_3042,N_2881,N_2536);
nand U3043 (N_3043,N_2854,N_2834);
and U3044 (N_3044,N_2181,N_2363);
or U3045 (N_3045,N_2618,N_2768);
nor U3046 (N_3046,N_2960,N_2616);
or U3047 (N_3047,N_2564,N_2627);
and U3048 (N_3048,N_2750,N_2642);
nand U3049 (N_3049,N_2034,N_2701);
nor U3050 (N_3050,N_2577,N_2176);
or U3051 (N_3051,N_2808,N_2286);
or U3052 (N_3052,N_2839,N_2796);
and U3053 (N_3053,N_2078,N_2337);
nor U3054 (N_3054,N_2964,N_2748);
or U3055 (N_3055,N_2462,N_2830);
nand U3056 (N_3056,N_2280,N_2979);
nand U3057 (N_3057,N_2920,N_2663);
or U3058 (N_3058,N_2978,N_2086);
and U3059 (N_3059,N_2098,N_2413);
xnor U3060 (N_3060,N_2200,N_2935);
and U3061 (N_3061,N_2297,N_2861);
nand U3062 (N_3062,N_2146,N_2744);
and U3063 (N_3063,N_2617,N_2017);
nand U3064 (N_3064,N_2218,N_2747);
nand U3065 (N_3065,N_2102,N_2999);
or U3066 (N_3066,N_2248,N_2253);
nand U3067 (N_3067,N_2532,N_2421);
nor U3068 (N_3068,N_2668,N_2866);
and U3069 (N_3069,N_2524,N_2474);
or U3070 (N_3070,N_2676,N_2806);
nand U3071 (N_3071,N_2045,N_2801);
nand U3072 (N_3072,N_2344,N_2124);
nor U3073 (N_3073,N_2323,N_2902);
nor U3074 (N_3074,N_2390,N_2064);
and U3075 (N_3075,N_2936,N_2783);
or U3076 (N_3076,N_2984,N_2171);
or U3077 (N_3077,N_2804,N_2373);
nor U3078 (N_3078,N_2449,N_2991);
and U3079 (N_3079,N_2145,N_2397);
nor U3080 (N_3080,N_2679,N_2652);
or U3081 (N_3081,N_2180,N_2549);
nor U3082 (N_3082,N_2848,N_2907);
and U3083 (N_3083,N_2068,N_2809);
or U3084 (N_3084,N_2401,N_2417);
or U3085 (N_3085,N_2704,N_2915);
and U3086 (N_3086,N_2026,N_2740);
nor U3087 (N_3087,N_2844,N_2502);
nand U3088 (N_3088,N_2263,N_2148);
and U3089 (N_3089,N_2589,N_2369);
or U3090 (N_3090,N_2666,N_2528);
nand U3091 (N_3091,N_2096,N_2347);
nor U3092 (N_3092,N_2826,N_2092);
and U3093 (N_3093,N_2538,N_2227);
nor U3094 (N_3094,N_2435,N_2514);
or U3095 (N_3095,N_2731,N_2242);
nor U3096 (N_3096,N_2396,N_2223);
or U3097 (N_3097,N_2054,N_2983);
nor U3098 (N_3098,N_2623,N_2949);
nor U3099 (N_3099,N_2038,N_2995);
and U3100 (N_3100,N_2074,N_2232);
and U3101 (N_3101,N_2908,N_2251);
nor U3102 (N_3102,N_2154,N_2516);
nor U3103 (N_3103,N_2603,N_2183);
nor U3104 (N_3104,N_2358,N_2926);
nor U3105 (N_3105,N_2921,N_2459);
nand U3106 (N_3106,N_2655,N_2606);
and U3107 (N_3107,N_2877,N_2653);
nand U3108 (N_3108,N_2178,N_2952);
nor U3109 (N_3109,N_2662,N_2426);
xor U3110 (N_3110,N_2446,N_2879);
nor U3111 (N_3111,N_2475,N_2754);
nor U3112 (N_3112,N_2442,N_2752);
nand U3113 (N_3113,N_2931,N_2354);
and U3114 (N_3114,N_2718,N_2023);
nor U3115 (N_3115,N_2381,N_2091);
and U3116 (N_3116,N_2476,N_2678);
and U3117 (N_3117,N_2272,N_2082);
and U3118 (N_3118,N_2827,N_2024);
nand U3119 (N_3119,N_2634,N_2664);
nand U3120 (N_3120,N_2243,N_2450);
nand U3121 (N_3121,N_2781,N_2592);
and U3122 (N_3122,N_2455,N_2779);
nor U3123 (N_3123,N_2231,N_2147);
nor U3124 (N_3124,N_2706,N_2605);
nand U3125 (N_3125,N_2981,N_2939);
nand U3126 (N_3126,N_2556,N_2265);
or U3127 (N_3127,N_2742,N_2451);
nand U3128 (N_3128,N_2945,N_2070);
nor U3129 (N_3129,N_2644,N_2383);
and U3130 (N_3130,N_2353,N_2574);
and U3131 (N_3131,N_2805,N_2711);
and U3132 (N_3132,N_2942,N_2340);
or U3133 (N_3133,N_2168,N_2785);
and U3134 (N_3134,N_2444,N_2416);
and U3135 (N_3135,N_2571,N_2859);
and U3136 (N_3136,N_2389,N_2963);
nand U3137 (N_3137,N_2955,N_2115);
nand U3138 (N_3138,N_2727,N_2403);
nor U3139 (N_3139,N_2941,N_2725);
and U3140 (N_3140,N_2152,N_2262);
or U3141 (N_3141,N_2486,N_2002);
and U3142 (N_3142,N_2443,N_2432);
and U3143 (N_3143,N_2405,N_2423);
xor U3144 (N_3144,N_2910,N_2687);
nor U3145 (N_3145,N_2794,N_2710);
and U3146 (N_3146,N_2332,N_2348);
and U3147 (N_3147,N_2270,N_2582);
nand U3148 (N_3148,N_2281,N_2889);
and U3149 (N_3149,N_2000,N_2094);
xor U3150 (N_3150,N_2010,N_2599);
nor U3151 (N_3151,N_2867,N_2224);
nand U3152 (N_3152,N_2370,N_2018);
nand U3153 (N_3153,N_2974,N_2119);
or U3154 (N_3154,N_2728,N_2215);
nand U3155 (N_3155,N_2699,N_2487);
or U3156 (N_3156,N_2492,N_2305);
and U3157 (N_3157,N_2361,N_2628);
nand U3158 (N_3158,N_2133,N_2880);
or U3159 (N_3159,N_2745,N_2067);
and U3160 (N_3160,N_2483,N_2414);
and U3161 (N_3161,N_2987,N_2968);
nor U3162 (N_3162,N_2684,N_2519);
nor U3163 (N_3163,N_2743,N_2680);
or U3164 (N_3164,N_2334,N_2185);
and U3165 (N_3165,N_2555,N_2543);
or U3166 (N_3166,N_2860,N_2776);
or U3167 (N_3167,N_2558,N_2940);
and U3168 (N_3168,N_2204,N_2873);
and U3169 (N_3169,N_2106,N_2667);
nand U3170 (N_3170,N_2255,N_2249);
or U3171 (N_3171,N_2598,N_2408);
nand U3172 (N_3172,N_2737,N_2723);
nand U3173 (N_3173,N_2732,N_2112);
and U3174 (N_3174,N_2563,N_2686);
or U3175 (N_3175,N_2371,N_2130);
or U3176 (N_3176,N_2189,N_2391);
and U3177 (N_3177,N_2328,N_2862);
nor U3178 (N_3178,N_2876,N_2016);
or U3179 (N_3179,N_2409,N_2448);
or U3180 (N_3180,N_2188,N_2500);
and U3181 (N_3181,N_2778,N_2454);
or U3182 (N_3182,N_2504,N_2512);
or U3183 (N_3183,N_2647,N_2774);
nor U3184 (N_3184,N_2887,N_2759);
nand U3185 (N_3185,N_2914,N_2738);
nand U3186 (N_3186,N_2138,N_2338);
nand U3187 (N_3187,N_2894,N_2650);
nor U3188 (N_3188,N_2439,N_2175);
or U3189 (N_3189,N_2659,N_2665);
nor U3190 (N_3190,N_2816,N_2506);
nor U3191 (N_3191,N_2714,N_2143);
nor U3192 (N_3192,N_2734,N_2669);
nand U3193 (N_3193,N_2445,N_2021);
nor U3194 (N_3194,N_2318,N_2007);
or U3195 (N_3195,N_2386,N_2166);
nor U3196 (N_3196,N_2724,N_2051);
nor U3197 (N_3197,N_2544,N_2875);
and U3198 (N_3198,N_2932,N_2966);
and U3199 (N_3199,N_2890,N_2625);
nor U3200 (N_3200,N_2321,N_2037);
nor U3201 (N_3201,N_2292,N_2013);
nor U3202 (N_3202,N_2566,N_2675);
nand U3203 (N_3203,N_2851,N_2325);
and U3204 (N_3204,N_2682,N_2720);
or U3205 (N_3205,N_2129,N_2683);
nand U3206 (N_3206,N_2029,N_2847);
xor U3207 (N_3207,N_2685,N_2028);
nand U3208 (N_3208,N_2818,N_2893);
nor U3209 (N_3209,N_2523,N_2111);
nand U3210 (N_3210,N_2278,N_2244);
and U3211 (N_3211,N_2288,N_2144);
nand U3212 (N_3212,N_2638,N_2590);
or U3213 (N_3213,N_2060,N_2922);
nand U3214 (N_3214,N_2871,N_2375);
or U3215 (N_3215,N_2797,N_2327);
nand U3216 (N_3216,N_2641,N_2019);
nand U3217 (N_3217,N_2733,N_2020);
and U3218 (N_3218,N_2367,N_2619);
nor U3219 (N_3219,N_2657,N_2097);
nand U3220 (N_3220,N_2937,N_2122);
nand U3221 (N_3221,N_2858,N_2201);
nor U3222 (N_3222,N_2793,N_2174);
nor U3223 (N_3223,N_2190,N_2302);
and U3224 (N_3224,N_2431,N_2885);
and U3225 (N_3225,N_2043,N_2394);
nand U3226 (N_3226,N_2674,N_2635);
nor U3227 (N_3227,N_2460,N_2163);
or U3228 (N_3228,N_2125,N_2535);
nor U3229 (N_3229,N_2520,N_2509);
nand U3230 (N_3230,N_2656,N_2735);
and U3231 (N_3231,N_2303,N_2191);
or U3232 (N_3232,N_2259,N_2812);
nor U3233 (N_3233,N_2027,N_2469);
and U3234 (N_3234,N_2427,N_2071);
and U3235 (N_3235,N_2929,N_2632);
nand U3236 (N_3236,N_2578,N_2865);
and U3237 (N_3237,N_2093,N_2210);
nand U3238 (N_3238,N_2031,N_2357);
and U3239 (N_3239,N_2131,N_2447);
or U3240 (N_3240,N_2461,N_2081);
or U3241 (N_3241,N_2372,N_2114);
and U3242 (N_3242,N_2433,N_2550);
and U3243 (N_3243,N_2787,N_2693);
nand U3244 (N_3244,N_2220,N_2588);
nor U3245 (N_3245,N_2407,N_2843);
and U3246 (N_3246,N_2385,N_2241);
or U3247 (N_3247,N_2600,N_2203);
and U3248 (N_3248,N_2746,N_2722);
nor U3249 (N_3249,N_2436,N_2496);
or U3250 (N_3250,N_2891,N_2525);
nand U3251 (N_3251,N_2101,N_2756);
and U3252 (N_3252,N_2946,N_2398);
or U3253 (N_3253,N_2717,N_2782);
xor U3254 (N_3254,N_2150,N_2786);
or U3255 (N_3255,N_2584,N_2330);
nand U3256 (N_3256,N_2917,N_2766);
nor U3257 (N_3257,N_2410,N_2973);
nand U3258 (N_3258,N_2602,N_2003);
or U3259 (N_3259,N_2624,N_2471);
nand U3260 (N_3260,N_2790,N_2015);
xnor U3261 (N_3261,N_2621,N_2257);
nor U3262 (N_3262,N_2962,N_2298);
nand U3263 (N_3263,N_2040,N_2324);
or U3264 (N_3264,N_2004,N_2009);
nor U3265 (N_3265,N_2153,N_2059);
and U3266 (N_3266,N_2333,N_2882);
or U3267 (N_3267,N_2553,N_2485);
or U3268 (N_3268,N_2279,N_2594);
nand U3269 (N_3269,N_2368,N_2715);
nor U3270 (N_3270,N_2463,N_2359);
nand U3271 (N_3271,N_2484,N_2149);
nand U3272 (N_3272,N_2121,N_2835);
or U3273 (N_3273,N_2365,N_2763);
or U3274 (N_3274,N_2226,N_2415);
nor U3275 (N_3275,N_2275,N_2789);
nand U3276 (N_3276,N_2264,N_2749);
or U3277 (N_3277,N_2108,N_2692);
and U3278 (N_3278,N_2184,N_2633);
nor U3279 (N_3279,N_2042,N_2465);
and U3280 (N_3280,N_2276,N_2237);
and U3281 (N_3281,N_2364,N_2384);
nand U3282 (N_3282,N_2470,N_2478);
and U3283 (N_3283,N_2205,N_2360);
nor U3284 (N_3284,N_2382,N_2545);
nand U3285 (N_3285,N_2196,N_2105);
and U3286 (N_3286,N_2961,N_2075);
and U3287 (N_3287,N_2229,N_2551);
nand U3288 (N_3288,N_2689,N_2956);
nand U3289 (N_3289,N_2006,N_2845);
nor U3290 (N_3290,N_2800,N_2503);
nor U3291 (N_3291,N_2362,N_2140);
nand U3292 (N_3292,N_2565,N_2273);
or U3293 (N_3293,N_2355,N_2221);
or U3294 (N_3294,N_2139,N_2458);
and U3295 (N_3295,N_2036,N_2948);
or U3296 (N_3296,N_2586,N_2900);
xor U3297 (N_3297,N_2700,N_2857);
and U3298 (N_3298,N_2233,N_2831);
nor U3299 (N_3299,N_2729,N_2596);
nor U3300 (N_3300,N_2958,N_2245);
and U3301 (N_3301,N_2928,N_2671);
or U3302 (N_3302,N_2493,N_2807);
nor U3303 (N_3303,N_2411,N_2870);
nor U3304 (N_3304,N_2741,N_2972);
or U3305 (N_3305,N_2311,N_2772);
or U3306 (N_3306,N_2622,N_2169);
or U3307 (N_3307,N_2608,N_2425);
or U3308 (N_3308,N_2309,N_2250);
nand U3309 (N_3309,N_2698,N_2645);
nor U3310 (N_3310,N_2050,N_2195);
nor U3311 (N_3311,N_2951,N_2395);
nor U3312 (N_3312,N_2856,N_2762);
nor U3313 (N_3313,N_2672,N_2317);
and U3314 (N_3314,N_2366,N_2810);
nand U3315 (N_3315,N_2457,N_2300);
or U3316 (N_3316,N_2331,N_2755);
nor U3317 (N_3317,N_2083,N_2849);
and U3318 (N_3318,N_2261,N_2969);
or U3319 (N_3319,N_2982,N_2240);
and U3320 (N_3320,N_2490,N_2378);
nand U3321 (N_3321,N_2222,N_2899);
or U3322 (N_3322,N_2198,N_2607);
or U3323 (N_3323,N_2287,N_2883);
and U3324 (N_3324,N_2646,N_2295);
or U3325 (N_3325,N_2141,N_2924);
or U3326 (N_3326,N_2841,N_2660);
or U3327 (N_3327,N_2959,N_2906);
nand U3328 (N_3328,N_2252,N_2977);
or U3329 (N_3329,N_2468,N_2170);
and U3330 (N_3330,N_2167,N_2576);
or U3331 (N_3331,N_2869,N_2441);
or U3332 (N_3332,N_2160,N_2909);
or U3333 (N_3333,N_2118,N_2587);
and U3334 (N_3334,N_2117,N_2452);
nor U3335 (N_3335,N_2927,N_2923);
nor U3336 (N_3336,N_2254,N_2517);
and U3337 (N_3337,N_2505,N_2897);
nand U3338 (N_3338,N_2177,N_2895);
nand U3339 (N_3339,N_2246,N_2049);
or U3340 (N_3340,N_2719,N_2216);
nand U3341 (N_3341,N_2012,N_2537);
or U3342 (N_3342,N_2219,N_2819);
nand U3343 (N_3343,N_2100,N_2661);
nand U3344 (N_3344,N_2047,N_2211);
or U3345 (N_3345,N_2651,N_2716);
or U3346 (N_3346,N_2199,N_2878);
nand U3347 (N_3347,N_2356,N_2572);
or U3348 (N_3348,N_2613,N_2062);
nand U3349 (N_3349,N_2501,N_2868);
nor U3350 (N_3350,N_2850,N_2299);
nand U3351 (N_3351,N_2329,N_2322);
nor U3352 (N_3352,N_2202,N_2548);
or U3353 (N_3353,N_2898,N_2151);
nand U3354 (N_3354,N_2239,N_2351);
and U3355 (N_3355,N_2132,N_2301);
or U3356 (N_3356,N_2412,N_2648);
nand U3357 (N_3357,N_2495,N_2802);
xor U3358 (N_3358,N_2157,N_2316);
nand U3359 (N_3359,N_2041,N_2336);
nor U3360 (N_3360,N_2957,N_2533);
nand U3361 (N_3361,N_2268,N_2137);
nand U3362 (N_3362,N_2467,N_2998);
nor U3363 (N_3363,N_2025,N_2580);
and U3364 (N_3364,N_2821,N_2604);
nor U3365 (N_3365,N_2345,N_2304);
nand U3366 (N_3366,N_2499,N_2583);
nand U3367 (N_3367,N_2777,N_2341);
and U3368 (N_3368,N_2422,N_2597);
nor U3369 (N_3369,N_2730,N_2420);
nand U3370 (N_3370,N_2511,N_2829);
xor U3371 (N_3371,N_2079,N_2649);
xor U3372 (N_3372,N_2526,N_2691);
nand U3373 (N_3373,N_2063,N_2156);
or U3374 (N_3374,N_2836,N_2213);
and U3375 (N_3375,N_2274,N_2187);
or U3376 (N_3376,N_2530,N_2825);
xor U3377 (N_3377,N_2912,N_2110);
nor U3378 (N_3378,N_2842,N_2751);
or U3379 (N_3379,N_2557,N_2925);
or U3380 (N_3380,N_2757,N_2289);
nand U3381 (N_3381,N_2788,N_2142);
and U3382 (N_3382,N_2726,N_2943);
or U3383 (N_3383,N_2313,N_2784);
nor U3384 (N_3384,N_2282,N_2620);
nor U3385 (N_3385,N_2234,N_2614);
nand U3386 (N_3386,N_2208,N_2708);
and U3387 (N_3387,N_2335,N_2235);
or U3388 (N_3388,N_2838,N_2306);
nand U3389 (N_3389,N_2155,N_2569);
nand U3390 (N_3390,N_2498,N_2712);
nand U3391 (N_3391,N_2575,N_2822);
xnor U3392 (N_3392,N_2069,N_2769);
nand U3393 (N_3393,N_2527,N_2291);
nor U3394 (N_3394,N_2022,N_2612);
nor U3395 (N_3395,N_2758,N_2217);
nand U3396 (N_3396,N_2392,N_2032);
nand U3397 (N_3397,N_2052,N_2186);
nor U3398 (N_3398,N_2343,N_2985);
or U3399 (N_3399,N_2035,N_2944);
nor U3400 (N_3400,N_2214,N_2308);
or U3401 (N_3401,N_2872,N_2033);
and U3402 (N_3402,N_2429,N_2702);
nand U3403 (N_3403,N_2088,N_2992);
nor U3404 (N_3404,N_2374,N_2095);
nand U3405 (N_3405,N_2803,N_2058);
or U3406 (N_3406,N_2934,N_2158);
or U3407 (N_3407,N_2404,N_2387);
nor U3408 (N_3408,N_2464,N_2611);
nand U3409 (N_3409,N_2585,N_2434);
nand U3410 (N_3410,N_2077,N_2339);
nand U3411 (N_3411,N_2212,N_2192);
and U3412 (N_3412,N_2874,N_2795);
or U3413 (N_3413,N_2919,N_2497);
and U3414 (N_3414,N_2103,N_2440);
and U3415 (N_3415,N_2113,N_2342);
nor U3416 (N_3416,N_2739,N_2307);
and U3417 (N_3417,N_2547,N_2888);
and U3418 (N_3418,N_2595,N_2636);
nand U3419 (N_3419,N_2541,N_2938);
or U3420 (N_3420,N_2903,N_2135);
or U3421 (N_3421,N_2513,N_2430);
or U3422 (N_3422,N_2207,N_2066);
nand U3423 (N_3423,N_2428,N_2399);
and U3424 (N_3424,N_2388,N_2697);
or U3425 (N_3425,N_2561,N_2761);
nor U3426 (N_3426,N_2673,N_2820);
or U3427 (N_3427,N_2480,N_2542);
nand U3428 (N_3428,N_2481,N_2593);
or U3429 (N_3429,N_2852,N_2529);
or U3430 (N_3430,N_2126,N_2579);
and U3431 (N_3431,N_2515,N_2164);
and U3432 (N_3432,N_2377,N_2127);
nand U3433 (N_3433,N_2030,N_2087);
nand U3434 (N_3434,N_2466,N_2610);
and U3435 (N_3435,N_2546,N_2713);
or U3436 (N_3436,N_2236,N_2061);
or U3437 (N_3437,N_2228,N_2531);
nand U3438 (N_3438,N_2048,N_2993);
nand U3439 (N_3439,N_2290,N_2918);
nand U3440 (N_3440,N_2694,N_2832);
and U3441 (N_3441,N_2767,N_2319);
nor U3442 (N_3442,N_2472,N_2039);
or U3443 (N_3443,N_2197,N_2055);
and U3444 (N_3444,N_2350,N_2916);
nor U3445 (N_3445,N_2014,N_2312);
or U3446 (N_3446,N_2508,N_2609);
nand U3447 (N_3447,N_2269,N_2161);
and U3448 (N_3448,N_2953,N_2539);
nand U3449 (N_3449,N_2824,N_2721);
nand U3450 (N_3450,N_2853,N_2284);
nor U3451 (N_3451,N_2107,N_2811);
xor U3452 (N_3452,N_2456,N_2085);
nor U3453 (N_3453,N_2182,N_2230);
and U3454 (N_3454,N_2056,N_2709);
and U3455 (N_3455,N_2393,N_2238);
and U3456 (N_3456,N_2760,N_2315);
or U3457 (N_3457,N_2658,N_2090);
and U3458 (N_3458,N_2967,N_2954);
and U3459 (N_3459,N_2008,N_2905);
or U3460 (N_3460,N_2522,N_2294);
nand U3461 (N_3461,N_2688,N_2494);
or U3462 (N_3462,N_2293,N_2453);
or U3463 (N_3463,N_2099,N_2846);
nor U3464 (N_3464,N_2864,N_2406);
and U3465 (N_3465,N_2994,N_2165);
and U3466 (N_3466,N_2123,N_2591);
nand U3467 (N_3467,N_2975,N_2568);
and U3468 (N_3468,N_2562,N_2573);
and U3469 (N_3469,N_2172,N_2310);
nand U3470 (N_3470,N_2554,N_2643);
and U3471 (N_3471,N_2814,N_2247);
nand U3472 (N_3472,N_2765,N_2933);
or U3473 (N_3473,N_2346,N_2209);
and U3474 (N_3474,N_2855,N_2631);
nand U3475 (N_3475,N_2988,N_2823);
or U3476 (N_3476,N_2837,N_2352);
xnor U3477 (N_3477,N_2109,N_2073);
or U3478 (N_3478,N_2695,N_2491);
nand U3479 (N_3479,N_2225,N_2285);
nand U3480 (N_3480,N_2424,N_2913);
and U3481 (N_3481,N_2764,N_2266);
nor U3482 (N_3482,N_2677,N_2892);
nand U3483 (N_3483,N_2736,N_2771);
nor U3484 (N_3484,N_2639,N_2817);
or U3485 (N_3485,N_2626,N_2886);
or U3486 (N_3486,N_2076,N_2419);
nor U3487 (N_3487,N_2581,N_2402);
nor U3488 (N_3488,N_2775,N_2488);
nor U3489 (N_3489,N_2930,N_2863);
nor U3490 (N_3490,N_2540,N_2120);
or U3491 (N_3491,N_2989,N_2001);
nor U3492 (N_3492,N_2128,N_2005);
nor U3493 (N_3493,N_2896,N_2629);
nor U3494 (N_3494,N_2707,N_2521);
nand U3495 (N_3495,N_2884,N_2438);
and U3496 (N_3496,N_2134,N_2791);
nor U3497 (N_3497,N_2799,N_2046);
or U3498 (N_3498,N_2510,N_2570);
and U3499 (N_3499,N_2089,N_2534);
nand U3500 (N_3500,N_2020,N_2969);
nand U3501 (N_3501,N_2241,N_2295);
or U3502 (N_3502,N_2399,N_2994);
nor U3503 (N_3503,N_2966,N_2447);
nor U3504 (N_3504,N_2990,N_2574);
nor U3505 (N_3505,N_2628,N_2134);
and U3506 (N_3506,N_2936,N_2692);
nor U3507 (N_3507,N_2274,N_2851);
nand U3508 (N_3508,N_2511,N_2844);
and U3509 (N_3509,N_2647,N_2797);
nand U3510 (N_3510,N_2177,N_2455);
nor U3511 (N_3511,N_2508,N_2592);
or U3512 (N_3512,N_2019,N_2341);
nor U3513 (N_3513,N_2630,N_2167);
or U3514 (N_3514,N_2326,N_2644);
nor U3515 (N_3515,N_2205,N_2456);
nand U3516 (N_3516,N_2121,N_2994);
and U3517 (N_3517,N_2795,N_2102);
nor U3518 (N_3518,N_2110,N_2157);
nand U3519 (N_3519,N_2571,N_2504);
and U3520 (N_3520,N_2133,N_2181);
nor U3521 (N_3521,N_2554,N_2766);
nand U3522 (N_3522,N_2731,N_2780);
nor U3523 (N_3523,N_2550,N_2181);
nand U3524 (N_3524,N_2792,N_2856);
xor U3525 (N_3525,N_2581,N_2244);
xnor U3526 (N_3526,N_2946,N_2848);
or U3527 (N_3527,N_2452,N_2203);
nand U3528 (N_3528,N_2813,N_2646);
or U3529 (N_3529,N_2541,N_2902);
xor U3530 (N_3530,N_2869,N_2502);
or U3531 (N_3531,N_2381,N_2163);
and U3532 (N_3532,N_2214,N_2182);
nand U3533 (N_3533,N_2897,N_2884);
nor U3534 (N_3534,N_2005,N_2702);
and U3535 (N_3535,N_2937,N_2101);
nand U3536 (N_3536,N_2971,N_2422);
nor U3537 (N_3537,N_2578,N_2745);
and U3538 (N_3538,N_2564,N_2467);
or U3539 (N_3539,N_2717,N_2562);
nor U3540 (N_3540,N_2671,N_2969);
or U3541 (N_3541,N_2051,N_2082);
and U3542 (N_3542,N_2174,N_2949);
and U3543 (N_3543,N_2681,N_2302);
or U3544 (N_3544,N_2676,N_2334);
nand U3545 (N_3545,N_2730,N_2560);
nor U3546 (N_3546,N_2687,N_2547);
nor U3547 (N_3547,N_2138,N_2032);
or U3548 (N_3548,N_2176,N_2296);
nand U3549 (N_3549,N_2056,N_2041);
nor U3550 (N_3550,N_2187,N_2803);
or U3551 (N_3551,N_2054,N_2014);
nand U3552 (N_3552,N_2579,N_2789);
nand U3553 (N_3553,N_2786,N_2873);
nand U3554 (N_3554,N_2436,N_2831);
nor U3555 (N_3555,N_2613,N_2180);
nor U3556 (N_3556,N_2539,N_2662);
nor U3557 (N_3557,N_2655,N_2391);
nor U3558 (N_3558,N_2043,N_2565);
nor U3559 (N_3559,N_2215,N_2370);
nor U3560 (N_3560,N_2236,N_2258);
and U3561 (N_3561,N_2275,N_2256);
or U3562 (N_3562,N_2855,N_2514);
nand U3563 (N_3563,N_2156,N_2300);
nor U3564 (N_3564,N_2138,N_2523);
and U3565 (N_3565,N_2821,N_2716);
or U3566 (N_3566,N_2213,N_2705);
nand U3567 (N_3567,N_2892,N_2354);
nor U3568 (N_3568,N_2233,N_2604);
nor U3569 (N_3569,N_2998,N_2628);
xor U3570 (N_3570,N_2258,N_2461);
nor U3571 (N_3571,N_2358,N_2599);
and U3572 (N_3572,N_2307,N_2229);
and U3573 (N_3573,N_2160,N_2138);
nand U3574 (N_3574,N_2299,N_2630);
and U3575 (N_3575,N_2834,N_2264);
xor U3576 (N_3576,N_2834,N_2586);
or U3577 (N_3577,N_2221,N_2431);
nand U3578 (N_3578,N_2636,N_2123);
nor U3579 (N_3579,N_2393,N_2969);
and U3580 (N_3580,N_2364,N_2905);
nor U3581 (N_3581,N_2884,N_2877);
nand U3582 (N_3582,N_2016,N_2607);
or U3583 (N_3583,N_2853,N_2610);
nand U3584 (N_3584,N_2512,N_2726);
or U3585 (N_3585,N_2319,N_2802);
nand U3586 (N_3586,N_2684,N_2860);
nor U3587 (N_3587,N_2057,N_2931);
or U3588 (N_3588,N_2007,N_2486);
nand U3589 (N_3589,N_2911,N_2059);
or U3590 (N_3590,N_2636,N_2943);
or U3591 (N_3591,N_2295,N_2603);
and U3592 (N_3592,N_2177,N_2116);
or U3593 (N_3593,N_2240,N_2101);
and U3594 (N_3594,N_2442,N_2257);
xnor U3595 (N_3595,N_2296,N_2523);
or U3596 (N_3596,N_2741,N_2462);
nor U3597 (N_3597,N_2282,N_2833);
nand U3598 (N_3598,N_2232,N_2739);
and U3599 (N_3599,N_2815,N_2483);
and U3600 (N_3600,N_2270,N_2603);
and U3601 (N_3601,N_2981,N_2872);
nor U3602 (N_3602,N_2338,N_2323);
nor U3603 (N_3603,N_2443,N_2096);
and U3604 (N_3604,N_2366,N_2270);
and U3605 (N_3605,N_2037,N_2641);
nand U3606 (N_3606,N_2099,N_2608);
xnor U3607 (N_3607,N_2305,N_2851);
or U3608 (N_3608,N_2241,N_2200);
xor U3609 (N_3609,N_2239,N_2078);
or U3610 (N_3610,N_2668,N_2030);
nand U3611 (N_3611,N_2568,N_2812);
nand U3612 (N_3612,N_2394,N_2391);
and U3613 (N_3613,N_2355,N_2094);
nor U3614 (N_3614,N_2740,N_2705);
xnor U3615 (N_3615,N_2419,N_2694);
nor U3616 (N_3616,N_2706,N_2820);
or U3617 (N_3617,N_2391,N_2046);
or U3618 (N_3618,N_2157,N_2788);
or U3619 (N_3619,N_2970,N_2515);
nand U3620 (N_3620,N_2984,N_2799);
or U3621 (N_3621,N_2185,N_2660);
nand U3622 (N_3622,N_2201,N_2129);
nor U3623 (N_3623,N_2586,N_2805);
and U3624 (N_3624,N_2958,N_2960);
nand U3625 (N_3625,N_2982,N_2496);
xnor U3626 (N_3626,N_2067,N_2530);
and U3627 (N_3627,N_2157,N_2005);
and U3628 (N_3628,N_2167,N_2055);
nor U3629 (N_3629,N_2720,N_2502);
nor U3630 (N_3630,N_2704,N_2153);
nand U3631 (N_3631,N_2932,N_2917);
and U3632 (N_3632,N_2501,N_2149);
and U3633 (N_3633,N_2520,N_2826);
nand U3634 (N_3634,N_2670,N_2945);
nand U3635 (N_3635,N_2831,N_2657);
nor U3636 (N_3636,N_2635,N_2601);
nor U3637 (N_3637,N_2226,N_2938);
nand U3638 (N_3638,N_2156,N_2534);
nand U3639 (N_3639,N_2887,N_2543);
and U3640 (N_3640,N_2836,N_2553);
nand U3641 (N_3641,N_2203,N_2733);
nand U3642 (N_3642,N_2846,N_2685);
nor U3643 (N_3643,N_2157,N_2862);
nand U3644 (N_3644,N_2874,N_2180);
and U3645 (N_3645,N_2588,N_2961);
nor U3646 (N_3646,N_2054,N_2674);
or U3647 (N_3647,N_2770,N_2819);
or U3648 (N_3648,N_2137,N_2958);
nand U3649 (N_3649,N_2772,N_2723);
nor U3650 (N_3650,N_2519,N_2457);
nor U3651 (N_3651,N_2403,N_2899);
or U3652 (N_3652,N_2919,N_2408);
and U3653 (N_3653,N_2184,N_2722);
or U3654 (N_3654,N_2912,N_2687);
nor U3655 (N_3655,N_2279,N_2630);
nor U3656 (N_3656,N_2525,N_2822);
nor U3657 (N_3657,N_2434,N_2157);
or U3658 (N_3658,N_2233,N_2781);
nand U3659 (N_3659,N_2718,N_2737);
nand U3660 (N_3660,N_2931,N_2504);
nand U3661 (N_3661,N_2086,N_2403);
or U3662 (N_3662,N_2593,N_2108);
and U3663 (N_3663,N_2691,N_2716);
or U3664 (N_3664,N_2346,N_2268);
or U3665 (N_3665,N_2816,N_2118);
nand U3666 (N_3666,N_2035,N_2251);
or U3667 (N_3667,N_2011,N_2293);
nand U3668 (N_3668,N_2996,N_2204);
nor U3669 (N_3669,N_2681,N_2513);
or U3670 (N_3670,N_2710,N_2354);
nand U3671 (N_3671,N_2312,N_2385);
or U3672 (N_3672,N_2829,N_2124);
nand U3673 (N_3673,N_2605,N_2295);
nand U3674 (N_3674,N_2058,N_2856);
or U3675 (N_3675,N_2483,N_2991);
and U3676 (N_3676,N_2320,N_2155);
or U3677 (N_3677,N_2475,N_2173);
or U3678 (N_3678,N_2541,N_2993);
and U3679 (N_3679,N_2150,N_2599);
nand U3680 (N_3680,N_2082,N_2142);
or U3681 (N_3681,N_2193,N_2002);
or U3682 (N_3682,N_2430,N_2294);
or U3683 (N_3683,N_2910,N_2981);
xor U3684 (N_3684,N_2922,N_2475);
and U3685 (N_3685,N_2144,N_2757);
nor U3686 (N_3686,N_2583,N_2792);
nand U3687 (N_3687,N_2109,N_2152);
or U3688 (N_3688,N_2513,N_2939);
and U3689 (N_3689,N_2080,N_2821);
nor U3690 (N_3690,N_2307,N_2273);
or U3691 (N_3691,N_2678,N_2643);
nor U3692 (N_3692,N_2192,N_2945);
nand U3693 (N_3693,N_2669,N_2283);
or U3694 (N_3694,N_2631,N_2194);
or U3695 (N_3695,N_2530,N_2186);
nor U3696 (N_3696,N_2304,N_2287);
or U3697 (N_3697,N_2128,N_2460);
nor U3698 (N_3698,N_2800,N_2303);
and U3699 (N_3699,N_2884,N_2987);
xor U3700 (N_3700,N_2381,N_2546);
or U3701 (N_3701,N_2311,N_2871);
nor U3702 (N_3702,N_2673,N_2664);
nand U3703 (N_3703,N_2003,N_2236);
nor U3704 (N_3704,N_2022,N_2993);
and U3705 (N_3705,N_2441,N_2890);
nor U3706 (N_3706,N_2894,N_2668);
nand U3707 (N_3707,N_2550,N_2210);
or U3708 (N_3708,N_2173,N_2464);
nor U3709 (N_3709,N_2988,N_2381);
nand U3710 (N_3710,N_2185,N_2012);
nand U3711 (N_3711,N_2928,N_2846);
or U3712 (N_3712,N_2834,N_2742);
or U3713 (N_3713,N_2905,N_2360);
nand U3714 (N_3714,N_2231,N_2748);
or U3715 (N_3715,N_2321,N_2087);
nor U3716 (N_3716,N_2125,N_2394);
nor U3717 (N_3717,N_2852,N_2498);
or U3718 (N_3718,N_2651,N_2504);
nand U3719 (N_3719,N_2842,N_2350);
xnor U3720 (N_3720,N_2967,N_2873);
nor U3721 (N_3721,N_2373,N_2347);
nor U3722 (N_3722,N_2439,N_2952);
or U3723 (N_3723,N_2273,N_2713);
or U3724 (N_3724,N_2031,N_2794);
nand U3725 (N_3725,N_2437,N_2255);
nand U3726 (N_3726,N_2191,N_2097);
nand U3727 (N_3727,N_2355,N_2347);
or U3728 (N_3728,N_2117,N_2767);
nand U3729 (N_3729,N_2070,N_2508);
or U3730 (N_3730,N_2314,N_2053);
and U3731 (N_3731,N_2374,N_2926);
nand U3732 (N_3732,N_2662,N_2133);
and U3733 (N_3733,N_2518,N_2343);
and U3734 (N_3734,N_2307,N_2211);
xnor U3735 (N_3735,N_2296,N_2602);
nor U3736 (N_3736,N_2679,N_2593);
nor U3737 (N_3737,N_2402,N_2957);
nor U3738 (N_3738,N_2226,N_2746);
nand U3739 (N_3739,N_2002,N_2399);
nor U3740 (N_3740,N_2264,N_2590);
nand U3741 (N_3741,N_2460,N_2207);
and U3742 (N_3742,N_2991,N_2148);
nand U3743 (N_3743,N_2373,N_2357);
and U3744 (N_3744,N_2486,N_2412);
nor U3745 (N_3745,N_2389,N_2090);
and U3746 (N_3746,N_2214,N_2916);
nand U3747 (N_3747,N_2369,N_2749);
and U3748 (N_3748,N_2926,N_2475);
nand U3749 (N_3749,N_2018,N_2949);
nor U3750 (N_3750,N_2075,N_2668);
or U3751 (N_3751,N_2158,N_2905);
or U3752 (N_3752,N_2250,N_2383);
or U3753 (N_3753,N_2060,N_2565);
or U3754 (N_3754,N_2639,N_2169);
or U3755 (N_3755,N_2379,N_2903);
and U3756 (N_3756,N_2860,N_2441);
and U3757 (N_3757,N_2428,N_2367);
nor U3758 (N_3758,N_2671,N_2756);
and U3759 (N_3759,N_2746,N_2189);
and U3760 (N_3760,N_2372,N_2671);
nand U3761 (N_3761,N_2779,N_2378);
and U3762 (N_3762,N_2200,N_2845);
nor U3763 (N_3763,N_2341,N_2115);
nand U3764 (N_3764,N_2143,N_2881);
and U3765 (N_3765,N_2124,N_2319);
and U3766 (N_3766,N_2819,N_2991);
or U3767 (N_3767,N_2143,N_2952);
or U3768 (N_3768,N_2905,N_2622);
or U3769 (N_3769,N_2745,N_2166);
nand U3770 (N_3770,N_2887,N_2905);
or U3771 (N_3771,N_2117,N_2406);
or U3772 (N_3772,N_2524,N_2008);
and U3773 (N_3773,N_2261,N_2912);
nor U3774 (N_3774,N_2263,N_2586);
and U3775 (N_3775,N_2255,N_2328);
nand U3776 (N_3776,N_2527,N_2390);
nand U3777 (N_3777,N_2636,N_2864);
nand U3778 (N_3778,N_2024,N_2263);
nand U3779 (N_3779,N_2057,N_2745);
and U3780 (N_3780,N_2097,N_2892);
nor U3781 (N_3781,N_2770,N_2368);
and U3782 (N_3782,N_2701,N_2816);
or U3783 (N_3783,N_2927,N_2409);
nand U3784 (N_3784,N_2551,N_2215);
nor U3785 (N_3785,N_2947,N_2410);
or U3786 (N_3786,N_2232,N_2043);
or U3787 (N_3787,N_2805,N_2673);
and U3788 (N_3788,N_2550,N_2223);
nand U3789 (N_3789,N_2937,N_2179);
xnor U3790 (N_3790,N_2131,N_2897);
and U3791 (N_3791,N_2724,N_2156);
nor U3792 (N_3792,N_2342,N_2005);
and U3793 (N_3793,N_2115,N_2375);
nand U3794 (N_3794,N_2111,N_2956);
or U3795 (N_3795,N_2840,N_2059);
nand U3796 (N_3796,N_2731,N_2403);
nand U3797 (N_3797,N_2032,N_2960);
and U3798 (N_3798,N_2581,N_2693);
nor U3799 (N_3799,N_2302,N_2114);
and U3800 (N_3800,N_2125,N_2346);
nand U3801 (N_3801,N_2429,N_2930);
nand U3802 (N_3802,N_2596,N_2296);
or U3803 (N_3803,N_2653,N_2554);
nand U3804 (N_3804,N_2388,N_2738);
and U3805 (N_3805,N_2441,N_2562);
nand U3806 (N_3806,N_2924,N_2809);
or U3807 (N_3807,N_2789,N_2764);
or U3808 (N_3808,N_2011,N_2096);
and U3809 (N_3809,N_2313,N_2840);
or U3810 (N_3810,N_2636,N_2132);
and U3811 (N_3811,N_2635,N_2503);
and U3812 (N_3812,N_2045,N_2663);
or U3813 (N_3813,N_2068,N_2821);
nand U3814 (N_3814,N_2881,N_2111);
or U3815 (N_3815,N_2944,N_2101);
nand U3816 (N_3816,N_2114,N_2162);
nand U3817 (N_3817,N_2898,N_2747);
or U3818 (N_3818,N_2488,N_2320);
nand U3819 (N_3819,N_2493,N_2842);
or U3820 (N_3820,N_2616,N_2615);
or U3821 (N_3821,N_2950,N_2486);
nor U3822 (N_3822,N_2226,N_2003);
or U3823 (N_3823,N_2787,N_2035);
and U3824 (N_3824,N_2249,N_2044);
and U3825 (N_3825,N_2483,N_2325);
nand U3826 (N_3826,N_2149,N_2475);
and U3827 (N_3827,N_2831,N_2177);
nor U3828 (N_3828,N_2089,N_2726);
and U3829 (N_3829,N_2122,N_2394);
or U3830 (N_3830,N_2093,N_2006);
nor U3831 (N_3831,N_2018,N_2249);
nand U3832 (N_3832,N_2228,N_2155);
and U3833 (N_3833,N_2438,N_2146);
and U3834 (N_3834,N_2544,N_2506);
and U3835 (N_3835,N_2900,N_2365);
nor U3836 (N_3836,N_2328,N_2508);
nand U3837 (N_3837,N_2608,N_2376);
or U3838 (N_3838,N_2346,N_2280);
and U3839 (N_3839,N_2848,N_2258);
nor U3840 (N_3840,N_2968,N_2109);
nor U3841 (N_3841,N_2330,N_2336);
nand U3842 (N_3842,N_2493,N_2797);
xor U3843 (N_3843,N_2466,N_2391);
and U3844 (N_3844,N_2947,N_2920);
and U3845 (N_3845,N_2159,N_2865);
and U3846 (N_3846,N_2010,N_2700);
xnor U3847 (N_3847,N_2171,N_2802);
and U3848 (N_3848,N_2608,N_2098);
nand U3849 (N_3849,N_2473,N_2705);
and U3850 (N_3850,N_2126,N_2838);
nor U3851 (N_3851,N_2460,N_2812);
and U3852 (N_3852,N_2936,N_2898);
or U3853 (N_3853,N_2248,N_2147);
or U3854 (N_3854,N_2863,N_2877);
or U3855 (N_3855,N_2341,N_2358);
and U3856 (N_3856,N_2874,N_2634);
nand U3857 (N_3857,N_2186,N_2843);
and U3858 (N_3858,N_2413,N_2438);
and U3859 (N_3859,N_2437,N_2470);
and U3860 (N_3860,N_2962,N_2625);
nor U3861 (N_3861,N_2217,N_2126);
and U3862 (N_3862,N_2864,N_2882);
or U3863 (N_3863,N_2060,N_2427);
and U3864 (N_3864,N_2496,N_2023);
or U3865 (N_3865,N_2273,N_2324);
and U3866 (N_3866,N_2160,N_2039);
and U3867 (N_3867,N_2063,N_2027);
nor U3868 (N_3868,N_2685,N_2784);
or U3869 (N_3869,N_2126,N_2440);
nand U3870 (N_3870,N_2710,N_2924);
nand U3871 (N_3871,N_2345,N_2104);
nor U3872 (N_3872,N_2385,N_2395);
nand U3873 (N_3873,N_2047,N_2369);
and U3874 (N_3874,N_2634,N_2801);
nor U3875 (N_3875,N_2136,N_2859);
or U3876 (N_3876,N_2228,N_2738);
and U3877 (N_3877,N_2408,N_2014);
nor U3878 (N_3878,N_2220,N_2325);
nand U3879 (N_3879,N_2259,N_2763);
and U3880 (N_3880,N_2946,N_2197);
nor U3881 (N_3881,N_2301,N_2859);
nor U3882 (N_3882,N_2321,N_2655);
nor U3883 (N_3883,N_2023,N_2451);
xnor U3884 (N_3884,N_2995,N_2236);
nor U3885 (N_3885,N_2733,N_2971);
and U3886 (N_3886,N_2743,N_2079);
nand U3887 (N_3887,N_2350,N_2349);
nand U3888 (N_3888,N_2392,N_2932);
nor U3889 (N_3889,N_2736,N_2152);
xnor U3890 (N_3890,N_2901,N_2884);
and U3891 (N_3891,N_2410,N_2280);
or U3892 (N_3892,N_2680,N_2791);
or U3893 (N_3893,N_2496,N_2097);
and U3894 (N_3894,N_2673,N_2912);
nor U3895 (N_3895,N_2785,N_2897);
nor U3896 (N_3896,N_2342,N_2355);
nor U3897 (N_3897,N_2161,N_2976);
xor U3898 (N_3898,N_2422,N_2698);
or U3899 (N_3899,N_2625,N_2494);
nand U3900 (N_3900,N_2310,N_2526);
or U3901 (N_3901,N_2829,N_2500);
nand U3902 (N_3902,N_2103,N_2144);
nand U3903 (N_3903,N_2225,N_2737);
or U3904 (N_3904,N_2178,N_2865);
or U3905 (N_3905,N_2929,N_2504);
nand U3906 (N_3906,N_2828,N_2598);
and U3907 (N_3907,N_2828,N_2043);
nand U3908 (N_3908,N_2338,N_2466);
or U3909 (N_3909,N_2613,N_2671);
nand U3910 (N_3910,N_2523,N_2192);
nand U3911 (N_3911,N_2663,N_2282);
nand U3912 (N_3912,N_2390,N_2984);
nor U3913 (N_3913,N_2740,N_2571);
nor U3914 (N_3914,N_2650,N_2445);
nor U3915 (N_3915,N_2767,N_2476);
and U3916 (N_3916,N_2475,N_2429);
nand U3917 (N_3917,N_2647,N_2993);
nand U3918 (N_3918,N_2560,N_2625);
nand U3919 (N_3919,N_2581,N_2081);
and U3920 (N_3920,N_2943,N_2372);
nand U3921 (N_3921,N_2082,N_2030);
xor U3922 (N_3922,N_2926,N_2940);
and U3923 (N_3923,N_2457,N_2964);
and U3924 (N_3924,N_2533,N_2990);
and U3925 (N_3925,N_2501,N_2158);
or U3926 (N_3926,N_2983,N_2679);
and U3927 (N_3927,N_2101,N_2974);
nor U3928 (N_3928,N_2740,N_2800);
nand U3929 (N_3929,N_2861,N_2419);
and U3930 (N_3930,N_2293,N_2953);
or U3931 (N_3931,N_2119,N_2430);
nand U3932 (N_3932,N_2748,N_2615);
nand U3933 (N_3933,N_2400,N_2485);
nor U3934 (N_3934,N_2156,N_2743);
or U3935 (N_3935,N_2612,N_2909);
xnor U3936 (N_3936,N_2367,N_2578);
and U3937 (N_3937,N_2898,N_2109);
or U3938 (N_3938,N_2063,N_2870);
or U3939 (N_3939,N_2057,N_2509);
nand U3940 (N_3940,N_2850,N_2403);
and U3941 (N_3941,N_2312,N_2345);
or U3942 (N_3942,N_2006,N_2014);
nor U3943 (N_3943,N_2271,N_2995);
nand U3944 (N_3944,N_2606,N_2531);
and U3945 (N_3945,N_2178,N_2053);
or U3946 (N_3946,N_2060,N_2179);
or U3947 (N_3947,N_2657,N_2209);
and U3948 (N_3948,N_2364,N_2230);
or U3949 (N_3949,N_2393,N_2242);
and U3950 (N_3950,N_2033,N_2840);
xor U3951 (N_3951,N_2333,N_2629);
xor U3952 (N_3952,N_2049,N_2034);
and U3953 (N_3953,N_2374,N_2849);
nand U3954 (N_3954,N_2236,N_2539);
nor U3955 (N_3955,N_2489,N_2343);
nand U3956 (N_3956,N_2564,N_2881);
nor U3957 (N_3957,N_2768,N_2580);
nand U3958 (N_3958,N_2362,N_2135);
or U3959 (N_3959,N_2447,N_2667);
nor U3960 (N_3960,N_2777,N_2467);
nand U3961 (N_3961,N_2176,N_2522);
and U3962 (N_3962,N_2970,N_2630);
and U3963 (N_3963,N_2803,N_2287);
nand U3964 (N_3964,N_2819,N_2721);
and U3965 (N_3965,N_2750,N_2425);
nand U3966 (N_3966,N_2859,N_2691);
or U3967 (N_3967,N_2577,N_2985);
and U3968 (N_3968,N_2625,N_2333);
nor U3969 (N_3969,N_2298,N_2574);
nand U3970 (N_3970,N_2343,N_2910);
nor U3971 (N_3971,N_2763,N_2044);
nand U3972 (N_3972,N_2789,N_2044);
and U3973 (N_3973,N_2258,N_2101);
nand U3974 (N_3974,N_2916,N_2316);
xnor U3975 (N_3975,N_2043,N_2273);
or U3976 (N_3976,N_2573,N_2011);
or U3977 (N_3977,N_2240,N_2001);
and U3978 (N_3978,N_2533,N_2410);
or U3979 (N_3979,N_2565,N_2038);
nand U3980 (N_3980,N_2586,N_2944);
and U3981 (N_3981,N_2645,N_2585);
and U3982 (N_3982,N_2719,N_2695);
and U3983 (N_3983,N_2016,N_2030);
nand U3984 (N_3984,N_2763,N_2500);
nand U3985 (N_3985,N_2437,N_2245);
nor U3986 (N_3986,N_2449,N_2916);
and U3987 (N_3987,N_2637,N_2034);
nor U3988 (N_3988,N_2244,N_2435);
nand U3989 (N_3989,N_2965,N_2132);
nor U3990 (N_3990,N_2724,N_2025);
or U3991 (N_3991,N_2772,N_2652);
and U3992 (N_3992,N_2436,N_2936);
nor U3993 (N_3993,N_2564,N_2328);
and U3994 (N_3994,N_2391,N_2530);
and U3995 (N_3995,N_2299,N_2341);
or U3996 (N_3996,N_2904,N_2519);
nand U3997 (N_3997,N_2946,N_2543);
nand U3998 (N_3998,N_2120,N_2187);
or U3999 (N_3999,N_2936,N_2265);
or U4000 (N_4000,N_3978,N_3068);
nor U4001 (N_4001,N_3278,N_3173);
and U4002 (N_4002,N_3960,N_3267);
nor U4003 (N_4003,N_3134,N_3511);
nand U4004 (N_4004,N_3977,N_3467);
or U4005 (N_4005,N_3259,N_3917);
or U4006 (N_4006,N_3196,N_3652);
or U4007 (N_4007,N_3400,N_3739);
and U4008 (N_4008,N_3337,N_3265);
nand U4009 (N_4009,N_3148,N_3966);
nor U4010 (N_4010,N_3786,N_3307);
and U4011 (N_4011,N_3928,N_3813);
and U4012 (N_4012,N_3790,N_3581);
or U4013 (N_4013,N_3685,N_3546);
or U4014 (N_4014,N_3779,N_3998);
and U4015 (N_4015,N_3007,N_3863);
or U4016 (N_4016,N_3820,N_3482);
and U4017 (N_4017,N_3504,N_3205);
nor U4018 (N_4018,N_3553,N_3302);
and U4019 (N_4019,N_3980,N_3802);
or U4020 (N_4020,N_3251,N_3964);
nand U4021 (N_4021,N_3021,N_3164);
and U4022 (N_4022,N_3909,N_3975);
nand U4023 (N_4023,N_3049,N_3574);
nand U4024 (N_4024,N_3147,N_3984);
or U4025 (N_4025,N_3865,N_3279);
nand U4026 (N_4026,N_3835,N_3053);
and U4027 (N_4027,N_3392,N_3016);
nand U4028 (N_4028,N_3590,N_3605);
nand U4029 (N_4029,N_3564,N_3850);
or U4030 (N_4030,N_3014,N_3029);
and U4031 (N_4031,N_3247,N_3208);
and U4032 (N_4032,N_3241,N_3296);
and U4033 (N_4033,N_3602,N_3289);
nor U4034 (N_4034,N_3465,N_3498);
or U4035 (N_4035,N_3985,N_3712);
and U4036 (N_4036,N_3828,N_3249);
or U4037 (N_4037,N_3868,N_3988);
and U4038 (N_4038,N_3946,N_3209);
and U4039 (N_4039,N_3869,N_3027);
nand U4040 (N_4040,N_3615,N_3531);
nor U4041 (N_4041,N_3992,N_3806);
or U4042 (N_4042,N_3372,N_3993);
nor U4043 (N_4043,N_3672,N_3052);
nand U4044 (N_4044,N_3105,N_3922);
or U4045 (N_4045,N_3233,N_3000);
nor U4046 (N_4046,N_3810,N_3036);
and U4047 (N_4047,N_3461,N_3996);
or U4048 (N_4048,N_3074,N_3425);
or U4049 (N_4049,N_3862,N_3217);
or U4050 (N_4050,N_3558,N_3051);
and U4051 (N_4051,N_3312,N_3604);
xnor U4052 (N_4052,N_3211,N_3622);
or U4053 (N_4053,N_3124,N_3410);
and U4054 (N_4054,N_3837,N_3629);
nand U4055 (N_4055,N_3583,N_3385);
and U4056 (N_4056,N_3971,N_3152);
nand U4057 (N_4057,N_3018,N_3095);
nand U4058 (N_4058,N_3393,N_3576);
and U4059 (N_4059,N_3801,N_3623);
or U4060 (N_4060,N_3479,N_3765);
nor U4061 (N_4061,N_3065,N_3664);
or U4062 (N_4062,N_3642,N_3807);
or U4063 (N_4063,N_3663,N_3930);
xnor U4064 (N_4064,N_3509,N_3203);
and U4065 (N_4065,N_3476,N_3532);
or U4066 (N_4066,N_3376,N_3526);
or U4067 (N_4067,N_3387,N_3728);
xor U4068 (N_4068,N_3338,N_3167);
nand U4069 (N_4069,N_3731,N_3350);
nand U4070 (N_4070,N_3009,N_3874);
nand U4071 (N_4071,N_3543,N_3836);
nor U4072 (N_4072,N_3882,N_3236);
nand U4073 (N_4073,N_3643,N_3502);
and U4074 (N_4074,N_3774,N_3457);
xnor U4075 (N_4075,N_3035,N_3443);
nand U4076 (N_4076,N_3218,N_3128);
and U4077 (N_4077,N_3660,N_3157);
nor U4078 (N_4078,N_3573,N_3031);
nor U4079 (N_4079,N_3304,N_3495);
and U4080 (N_4080,N_3305,N_3441);
nor U4081 (N_4081,N_3488,N_3953);
or U4082 (N_4082,N_3618,N_3407);
or U4083 (N_4083,N_3194,N_3046);
nand U4084 (N_4084,N_3153,N_3800);
and U4085 (N_4085,N_3748,N_3055);
and U4086 (N_4086,N_3648,N_3355);
and U4087 (N_4087,N_3405,N_3780);
or U4088 (N_4088,N_3146,N_3037);
nor U4089 (N_4089,N_3131,N_3898);
nor U4090 (N_4090,N_3170,N_3635);
xor U4091 (N_4091,N_3151,N_3071);
or U4092 (N_4092,N_3261,N_3506);
nand U4093 (N_4093,N_3380,N_3881);
and U4094 (N_4094,N_3200,N_3115);
nand U4095 (N_4095,N_3655,N_3654);
or U4096 (N_4096,N_3831,N_3540);
nand U4097 (N_4097,N_3963,N_3178);
or U4098 (N_4098,N_3159,N_3453);
nand U4099 (N_4099,N_3704,N_3059);
nor U4100 (N_4100,N_3460,N_3693);
nor U4101 (N_4101,N_3340,N_3682);
xor U4102 (N_4102,N_3345,N_3673);
or U4103 (N_4103,N_3133,N_3891);
and U4104 (N_4104,N_3957,N_3593);
and U4105 (N_4105,N_3787,N_3058);
and U4106 (N_4106,N_3762,N_3269);
nor U4107 (N_4107,N_3137,N_3947);
nand U4108 (N_4108,N_3500,N_3149);
nor U4109 (N_4109,N_3421,N_3713);
xnor U4110 (N_4110,N_3944,N_3268);
or U4111 (N_4111,N_3180,N_3119);
nor U4112 (N_4112,N_3375,N_3794);
and U4113 (N_4113,N_3243,N_3462);
nor U4114 (N_4114,N_3478,N_3619);
nor U4115 (N_4115,N_3138,N_3219);
or U4116 (N_4116,N_3845,N_3078);
or U4117 (N_4117,N_3689,N_3044);
and U4118 (N_4118,N_3979,N_3444);
nor U4119 (N_4119,N_3588,N_3156);
or U4120 (N_4120,N_3606,N_3005);
or U4121 (N_4121,N_3033,N_3492);
or U4122 (N_4122,N_3601,N_3877);
or U4123 (N_4123,N_3950,N_3515);
nand U4124 (N_4124,N_3879,N_3730);
nor U4125 (N_4125,N_3120,N_3781);
or U4126 (N_4126,N_3347,N_3282);
nand U4127 (N_4127,N_3698,N_3143);
and U4128 (N_4128,N_3223,N_3633);
nand U4129 (N_4129,N_3314,N_3429);
nor U4130 (N_4130,N_3675,N_3534);
nand U4131 (N_4131,N_3079,N_3100);
nor U4132 (N_4132,N_3290,N_3199);
nor U4133 (N_4133,N_3113,N_3353);
and U4134 (N_4134,N_3741,N_3690);
nand U4135 (N_4135,N_3175,N_3808);
and U4136 (N_4136,N_3489,N_3589);
or U4137 (N_4137,N_3292,N_3439);
nand U4138 (N_4138,N_3545,N_3274);
nand U4139 (N_4139,N_3871,N_3132);
or U4140 (N_4140,N_3640,N_3067);
and U4141 (N_4141,N_3077,N_3649);
nor U4142 (N_4142,N_3603,N_3924);
or U4143 (N_4143,N_3771,N_3686);
and U4144 (N_4144,N_3291,N_3399);
nor U4145 (N_4145,N_3166,N_3123);
and U4146 (N_4146,N_3086,N_3396);
and U4147 (N_4147,N_3485,N_3112);
nand U4148 (N_4148,N_3644,N_3861);
nand U4149 (N_4149,N_3473,N_3755);
nor U4150 (N_4150,N_3165,N_3714);
or U4151 (N_4151,N_3093,N_3285);
nand U4152 (N_4152,N_3142,N_3263);
and U4153 (N_4153,N_3552,N_3094);
and U4154 (N_4154,N_3680,N_3880);
or U4155 (N_4155,N_3433,N_3384);
nor U4156 (N_4156,N_3325,N_3281);
nand U4157 (N_4157,N_3878,N_3008);
and U4158 (N_4158,N_3169,N_3856);
or U4159 (N_4159,N_3927,N_3620);
and U4160 (N_4160,N_3804,N_3459);
nor U4161 (N_4161,N_3313,N_3420);
and U4162 (N_4162,N_3791,N_3997);
nand U4163 (N_4163,N_3745,N_3542);
nand U4164 (N_4164,N_3404,N_3002);
and U4165 (N_4165,N_3426,N_3715);
or U4166 (N_4166,N_3413,N_3256);
and U4167 (N_4167,N_3557,N_3471);
nand U4168 (N_4168,N_3057,N_3162);
nor U4169 (N_4169,N_3773,N_3315);
and U4170 (N_4170,N_3104,N_3611);
and U4171 (N_4171,N_3674,N_3887);
and U4172 (N_4172,N_3150,N_3772);
or U4173 (N_4173,N_3554,N_3510);
and U4174 (N_4174,N_3535,N_3990);
nor U4175 (N_4175,N_3582,N_3419);
nand U4176 (N_4176,N_3976,N_3248);
nand U4177 (N_4177,N_3533,N_3207);
and U4178 (N_4178,N_3575,N_3215);
nand U4179 (N_4179,N_3254,N_3322);
nand U4180 (N_4180,N_3757,N_3161);
or U4181 (N_4181,N_3427,N_3452);
or U4182 (N_4182,N_3614,N_3587);
and U4183 (N_4183,N_3264,N_3799);
nand U4184 (N_4184,N_3702,N_3253);
and U4185 (N_4185,N_3965,N_3556);
xnor U4186 (N_4186,N_3190,N_3968);
or U4187 (N_4187,N_3592,N_3798);
or U4188 (N_4188,N_3395,N_3777);
nand U4189 (N_4189,N_3334,N_3516);
or U4190 (N_4190,N_3344,N_3567);
and U4191 (N_4191,N_3145,N_3232);
nand U4192 (N_4192,N_3273,N_3358);
nor U4193 (N_4193,N_3122,N_3106);
and U4194 (N_4194,N_3753,N_3885);
or U4195 (N_4195,N_3571,N_3902);
nand U4196 (N_4196,N_3328,N_3684);
and U4197 (N_4197,N_3499,N_3045);
or U4198 (N_4198,N_3701,N_3497);
and U4199 (N_4199,N_3906,N_3722);
nand U4200 (N_4200,N_3886,N_3659);
and U4201 (N_4201,N_3839,N_3933);
or U4202 (N_4202,N_3910,N_3025);
and U4203 (N_4203,N_3108,N_3570);
and U4204 (N_4204,N_3756,N_3843);
nor U4205 (N_4205,N_3359,N_3514);
and U4206 (N_4206,N_3080,N_3597);
nor U4207 (N_4207,N_3967,N_3691);
or U4208 (N_4208,N_3316,N_3809);
or U4209 (N_4209,N_3414,N_3003);
or U4210 (N_4210,N_3782,N_3637);
or U4211 (N_4211,N_3817,N_3069);
and U4212 (N_4212,N_3010,N_3555);
nor U4213 (N_4213,N_3607,N_3651);
and U4214 (N_4214,N_3948,N_3508);
nor U4215 (N_4215,N_3599,N_3107);
nand U4216 (N_4216,N_3921,N_3841);
nor U4217 (N_4217,N_3517,N_3415);
nor U4218 (N_4218,N_3747,N_3484);
nor U4219 (N_4219,N_3796,N_3284);
and U4220 (N_4220,N_3513,N_3280);
and U4221 (N_4221,N_3231,N_3222);
or U4222 (N_4222,N_3695,N_3671);
nand U4223 (N_4223,N_3491,N_3464);
nor U4224 (N_4224,N_3391,N_3901);
nor U4225 (N_4225,N_3923,N_3379);
and U4226 (N_4226,N_3524,N_3472);
nor U4227 (N_4227,N_3851,N_3198);
nor U4228 (N_4228,N_3110,N_3487);
nand U4229 (N_4229,N_3918,N_3463);
and U4230 (N_4230,N_3066,N_3125);
or U4231 (N_4231,N_3970,N_3949);
and U4232 (N_4232,N_3703,N_3854);
or U4233 (N_4233,N_3668,N_3445);
nor U4234 (N_4234,N_3667,N_3172);
nand U4235 (N_4235,N_3560,N_3934);
or U4236 (N_4236,N_3390,N_3617);
or U4237 (N_4237,N_3154,N_3317);
and U4238 (N_4238,N_3102,N_3039);
and U4239 (N_4239,N_3319,N_3048);
or U4240 (N_4240,N_3042,N_3099);
nor U4241 (N_4241,N_3306,N_3763);
and U4242 (N_4242,N_3266,N_3294);
or U4243 (N_4243,N_3189,N_3111);
nor U4244 (N_4244,N_3857,N_3889);
nand U4245 (N_4245,N_3406,N_3129);
xor U4246 (N_4246,N_3229,N_3665);
nor U4247 (N_4247,N_3752,N_3719);
and U4248 (N_4248,N_3028,N_3303);
nor U4249 (N_4249,N_3503,N_3174);
nor U4250 (N_4250,N_3913,N_3873);
nand U4251 (N_4251,N_3117,N_3367);
nand U4252 (N_4252,N_3494,N_3788);
and U4253 (N_4253,N_3864,N_3330);
nor U4254 (N_4254,N_3144,N_3805);
or U4255 (N_4255,N_3844,N_3013);
or U4256 (N_4256,N_3374,N_3234);
nand U4257 (N_4257,N_3213,N_3937);
nor U4258 (N_4258,N_3793,N_3116);
nand U4259 (N_4259,N_3182,N_3435);
and U4260 (N_4260,N_3432,N_3332);
and U4261 (N_4261,N_3724,N_3518);
or U4262 (N_4262,N_3521,N_3299);
nand U4263 (N_4263,N_3188,N_3608);
and U4264 (N_4264,N_3214,N_3321);
nand U4265 (N_4265,N_3226,N_3775);
nand U4266 (N_4266,N_3838,N_3335);
nor U4267 (N_4267,N_3795,N_3679);
xnor U4268 (N_4268,N_3666,N_3904);
nand U4269 (N_4269,N_3624,N_3210);
nor U4270 (N_4270,N_3382,N_3295);
or U4271 (N_4271,N_3015,N_3160);
nand U4272 (N_4272,N_3559,N_3610);
nor U4273 (N_4273,N_3830,N_3520);
or U4274 (N_4274,N_3056,N_3087);
nand U4275 (N_4275,N_3733,N_3536);
nand U4276 (N_4276,N_3181,N_3825);
or U4277 (N_4277,N_3446,N_3370);
or U4278 (N_4278,N_3754,N_3158);
and U4279 (N_4279,N_3721,N_3206);
and U4280 (N_4280,N_3797,N_3848);
and U4281 (N_4281,N_3434,N_3860);
and U4282 (N_4282,N_3293,N_3972);
or U4283 (N_4283,N_3938,N_3855);
nand U4284 (N_4284,N_3185,N_3186);
or U4285 (N_4285,N_3348,N_3600);
nor U4286 (N_4286,N_3477,N_3994);
and U4287 (N_4287,N_3041,N_3858);
and U4288 (N_4288,N_3054,N_3981);
nand U4289 (N_4289,N_3061,N_3101);
xor U4290 (N_4290,N_3237,N_3549);
nor U4291 (N_4291,N_3982,N_3778);
or U4292 (N_4292,N_3255,N_3512);
xnor U4293 (N_4293,N_3301,N_3076);
nand U4294 (N_4294,N_3935,N_3919);
and U4295 (N_4295,N_3431,N_3475);
nor U4296 (N_4296,N_3598,N_3866);
and U4297 (N_4297,N_3227,N_3287);
nor U4298 (N_4298,N_3230,N_3442);
nand U4299 (N_4299,N_3331,N_3789);
nand U4300 (N_4300,N_3566,N_3377);
nand U4301 (N_4301,N_3900,N_3720);
and U4302 (N_4302,N_3191,N_3951);
and U4303 (N_4303,N_3092,N_3272);
or U4304 (N_4304,N_3072,N_3677);
nor U4305 (N_4305,N_3939,N_3916);
nand U4306 (N_4306,N_3235,N_3995);
nand U4307 (N_4307,N_3818,N_3288);
and U4308 (N_4308,N_3245,N_3238);
and U4309 (N_4309,N_3271,N_3746);
or U4310 (N_4310,N_3723,N_3550);
or U4311 (N_4311,N_3811,N_3351);
xnor U4312 (N_4312,N_3883,N_3646);
or U4313 (N_4313,N_3539,N_3221);
xnor U4314 (N_4314,N_3662,N_3895);
xnor U4315 (N_4315,N_3631,N_3945);
nand U4316 (N_4316,N_3907,N_3091);
nand U4317 (N_4317,N_3070,N_3440);
and U4318 (N_4318,N_3941,N_3705);
and U4319 (N_4319,N_3023,N_3627);
xnor U4320 (N_4320,N_3171,N_3397);
or U4321 (N_4321,N_3929,N_3501);
nor U4322 (N_4322,N_3356,N_3011);
or U4323 (N_4323,N_3827,N_3639);
nor U4324 (N_4324,N_3468,N_3699);
nand U4325 (N_4325,N_3544,N_3636);
nor U4326 (N_4326,N_3676,N_3527);
and U4327 (N_4327,N_3139,N_3192);
and U4328 (N_4328,N_3661,N_3417);
nor U4329 (N_4329,N_3595,N_3656);
nor U4330 (N_4330,N_3034,N_3201);
nand U4331 (N_4331,N_3202,N_3803);
or U4332 (N_4332,N_3591,N_3038);
nor U4333 (N_4333,N_3381,N_3239);
nor U4334 (N_4334,N_3983,N_3456);
nor U4335 (N_4335,N_3650,N_3632);
and U4336 (N_4336,N_3451,N_3737);
or U4337 (N_4337,N_3899,N_3378);
nor U4338 (N_4338,N_3333,N_3759);
nand U4339 (N_4339,N_3454,N_3130);
or U4340 (N_4340,N_3709,N_3126);
nor U4341 (N_4341,N_3986,N_3341);
nor U4342 (N_4342,N_3075,N_3398);
and U4343 (N_4343,N_3692,N_3892);
or U4344 (N_4344,N_3228,N_3252);
nand U4345 (N_4345,N_3250,N_3257);
and U4346 (N_4346,N_3155,N_3389);
or U4347 (N_4347,N_3047,N_3565);
and U4348 (N_4348,N_3354,N_3784);
nand U4349 (N_4349,N_3954,N_3908);
nor U4350 (N_4350,N_3847,N_3840);
or U4351 (N_4351,N_3298,N_3019);
nor U4352 (N_4352,N_3750,N_3725);
nor U4353 (N_4353,N_3024,N_3541);
nor U4354 (N_4354,N_3323,N_3792);
and U4355 (N_4355,N_3177,N_3176);
or U4356 (N_4356,N_3824,N_3768);
or U4357 (N_4357,N_3262,N_3318);
nand U4358 (N_4358,N_3064,N_3483);
or U4359 (N_4359,N_3135,N_3926);
xnor U4360 (N_4360,N_3735,N_3326);
nand U4361 (N_4361,N_3140,N_3240);
nor U4362 (N_4362,N_3408,N_3630);
and U4363 (N_4363,N_3613,N_3537);
nand U4364 (N_4364,N_3829,N_3386);
or U4365 (N_4365,N_3700,N_3594);
nor U4366 (N_4366,N_3955,N_3320);
and U4367 (N_4367,N_3141,N_3530);
or U4368 (N_4368,N_3336,N_3876);
nand U4369 (N_4369,N_3849,N_3121);
xor U4370 (N_4370,N_3694,N_3548);
and U4371 (N_4371,N_3043,N_3991);
and U4372 (N_4372,N_3940,N_3342);
nand U4373 (N_4373,N_3022,N_3697);
and U4374 (N_4374,N_3767,N_3474);
and U4375 (N_4375,N_3496,N_3197);
nand U4376 (N_4376,N_3083,N_3727);
nor U4377 (N_4377,N_3311,N_3905);
and U4378 (N_4378,N_3505,N_3572);
and U4379 (N_4379,N_3961,N_3447);
nor U4380 (N_4380,N_3369,N_3383);
or U4381 (N_4381,N_3127,N_3696);
nand U4382 (N_4382,N_3062,N_3469);
nor U4383 (N_4383,N_3740,N_3578);
nor U4384 (N_4384,N_3932,N_3821);
nand U4385 (N_4385,N_3893,N_3989);
nor U4386 (N_4386,N_3846,N_3764);
or U4387 (N_4387,N_3678,N_3562);
or U4388 (N_4388,N_3276,N_3187);
and U4389 (N_4389,N_3911,N_3082);
nand U4390 (N_4390,N_3852,N_3450);
xnor U4391 (N_4391,N_3814,N_3084);
nand U4392 (N_4392,N_3621,N_3090);
and U4393 (N_4393,N_3364,N_3580);
nand U4394 (N_4394,N_3363,N_3738);
nor U4395 (N_4395,N_3073,N_3626);
or U4396 (N_4396,N_3920,N_3669);
nand U4397 (N_4397,N_3872,N_3834);
and U4398 (N_4398,N_3819,N_3822);
nand U4399 (N_4399,N_3523,N_3050);
nor U4400 (N_4400,N_3430,N_3212);
or U4401 (N_4401,N_3586,N_3455);
nand U4402 (N_4402,N_3815,N_3493);
and U4403 (N_4403,N_3224,N_3422);
and U4404 (N_4404,N_3958,N_3258);
nor U4405 (N_4405,N_3270,N_3758);
and U4406 (N_4406,N_3085,N_3402);
and U4407 (N_4407,N_3529,N_3436);
or U4408 (N_4408,N_3458,N_3179);
or U4409 (N_4409,N_3411,N_3569);
nor U4410 (N_4410,N_3718,N_3225);
or U4411 (N_4411,N_3522,N_3349);
and U4412 (N_4412,N_3744,N_3346);
nand U4413 (N_4413,N_3423,N_3641);
or U4414 (N_4414,N_3163,N_3418);
or U4415 (N_4415,N_3897,N_3109);
nand U4416 (N_4416,N_3388,N_3776);
and U4417 (N_4417,N_3030,N_3096);
or U4418 (N_4418,N_3769,N_3657);
xnor U4419 (N_4419,N_3711,N_3438);
or U4420 (N_4420,N_3726,N_3943);
nand U4421 (N_4421,N_3184,N_3625);
or U4422 (N_4422,N_3204,N_3584);
and U4423 (N_4423,N_3394,N_3097);
and U4424 (N_4424,N_3277,N_3244);
or U4425 (N_4425,N_3563,N_3357);
and U4426 (N_4426,N_3103,N_3300);
and U4427 (N_4427,N_3060,N_3361);
xnor U4428 (N_4428,N_3343,N_3373);
and U4429 (N_4429,N_3081,N_3216);
or U4430 (N_4430,N_3653,N_3716);
or U4431 (N_4431,N_3017,N_3729);
nand U4432 (N_4432,N_3596,N_3183);
nand U4433 (N_4433,N_3812,N_3412);
nor U4434 (N_4434,N_3551,N_3896);
or U4435 (N_4435,N_3638,N_3428);
or U4436 (N_4436,N_3365,N_3816);
and U4437 (N_4437,N_3761,N_3973);
or U4438 (N_4438,N_3890,N_3352);
nor U4439 (N_4439,N_3999,N_3339);
nand U4440 (N_4440,N_3195,N_3770);
nor U4441 (N_4441,N_3040,N_3360);
nor U4442 (N_4442,N_3751,N_3371);
nor U4443 (N_4443,N_3942,N_3853);
or U4444 (N_4444,N_3470,N_3585);
or U4445 (N_4445,N_3089,N_3118);
nor U4446 (N_4446,N_3708,N_3448);
nor U4447 (N_4447,N_3168,N_3688);
and U4448 (N_4448,N_3327,N_3063);
or U4449 (N_4449,N_3449,N_3760);
or U4450 (N_4450,N_3020,N_3275);
nand U4451 (N_4451,N_3310,N_3647);
and U4452 (N_4452,N_3974,N_3681);
and U4453 (N_4453,N_3088,N_3903);
nor U4454 (N_4454,N_3616,N_3519);
or U4455 (N_4455,N_3785,N_3006);
nor U4456 (N_4456,N_3687,N_3670);
or U4457 (N_4457,N_3736,N_3001);
or U4458 (N_4458,N_3579,N_3538);
or U4459 (N_4459,N_3634,N_3884);
or U4460 (N_4460,N_3561,N_3480);
nand U4461 (N_4461,N_3012,N_3888);
nand U4462 (N_4462,N_3658,N_3952);
or U4463 (N_4463,N_3547,N_3308);
xor U4464 (N_4464,N_3743,N_3842);
nor U4465 (N_4465,N_3416,N_3525);
or U4466 (N_4466,N_3568,N_3136);
xnor U4467 (N_4467,N_3914,N_3915);
nand U4468 (N_4468,N_3403,N_3437);
and U4469 (N_4469,N_3193,N_3286);
nor U4470 (N_4470,N_3706,N_3732);
nor U4471 (N_4471,N_3987,N_3242);
and U4472 (N_4472,N_3612,N_3826);
nor U4473 (N_4473,N_3833,N_3867);
or U4474 (N_4474,N_3098,N_3297);
and U4475 (N_4475,N_3324,N_3832);
and U4476 (N_4476,N_3894,N_3645);
nor U4477 (N_4477,N_3577,N_3875);
or U4478 (N_4478,N_3424,N_3368);
nor U4479 (N_4479,N_3742,N_3925);
nand U4480 (N_4480,N_3283,N_3956);
nor U4481 (N_4481,N_3628,N_3246);
and U4482 (N_4482,N_3366,N_3931);
and U4483 (N_4483,N_3466,N_3609);
or U4484 (N_4484,N_3962,N_3766);
and U4485 (N_4485,N_3329,N_3783);
and U4486 (N_4486,N_3912,N_3409);
or U4487 (N_4487,N_3490,N_3823);
nor U4488 (N_4488,N_3260,N_3528);
or U4489 (N_4489,N_3683,N_3401);
or U4490 (N_4490,N_3710,N_3707);
nor U4491 (N_4491,N_3507,N_3870);
and U4492 (N_4492,N_3734,N_3717);
or U4493 (N_4493,N_3481,N_3026);
and U4494 (N_4494,N_3004,N_3959);
nand U4495 (N_4495,N_3749,N_3362);
or U4496 (N_4496,N_3309,N_3114);
nor U4497 (N_4497,N_3859,N_3969);
and U4498 (N_4498,N_3936,N_3486);
or U4499 (N_4499,N_3220,N_3032);
nor U4500 (N_4500,N_3845,N_3320);
or U4501 (N_4501,N_3205,N_3858);
and U4502 (N_4502,N_3259,N_3124);
or U4503 (N_4503,N_3779,N_3365);
nand U4504 (N_4504,N_3429,N_3757);
and U4505 (N_4505,N_3422,N_3310);
nand U4506 (N_4506,N_3324,N_3480);
nor U4507 (N_4507,N_3219,N_3894);
or U4508 (N_4508,N_3692,N_3922);
nand U4509 (N_4509,N_3557,N_3829);
nor U4510 (N_4510,N_3783,N_3641);
and U4511 (N_4511,N_3342,N_3984);
or U4512 (N_4512,N_3801,N_3697);
or U4513 (N_4513,N_3323,N_3509);
nand U4514 (N_4514,N_3283,N_3450);
and U4515 (N_4515,N_3576,N_3676);
and U4516 (N_4516,N_3307,N_3973);
and U4517 (N_4517,N_3014,N_3239);
and U4518 (N_4518,N_3917,N_3271);
nor U4519 (N_4519,N_3519,N_3247);
or U4520 (N_4520,N_3371,N_3277);
nand U4521 (N_4521,N_3456,N_3590);
nand U4522 (N_4522,N_3220,N_3494);
nand U4523 (N_4523,N_3570,N_3381);
nand U4524 (N_4524,N_3356,N_3470);
and U4525 (N_4525,N_3355,N_3854);
nand U4526 (N_4526,N_3353,N_3164);
or U4527 (N_4527,N_3346,N_3675);
and U4528 (N_4528,N_3060,N_3495);
nor U4529 (N_4529,N_3233,N_3882);
nand U4530 (N_4530,N_3991,N_3681);
and U4531 (N_4531,N_3608,N_3527);
and U4532 (N_4532,N_3277,N_3416);
nand U4533 (N_4533,N_3664,N_3095);
nor U4534 (N_4534,N_3931,N_3482);
and U4535 (N_4535,N_3301,N_3079);
or U4536 (N_4536,N_3249,N_3573);
nor U4537 (N_4537,N_3464,N_3186);
and U4538 (N_4538,N_3443,N_3501);
and U4539 (N_4539,N_3811,N_3664);
or U4540 (N_4540,N_3262,N_3447);
nor U4541 (N_4541,N_3375,N_3712);
nor U4542 (N_4542,N_3517,N_3719);
nor U4543 (N_4543,N_3241,N_3601);
nand U4544 (N_4544,N_3752,N_3154);
and U4545 (N_4545,N_3430,N_3280);
nand U4546 (N_4546,N_3912,N_3133);
nor U4547 (N_4547,N_3632,N_3939);
nor U4548 (N_4548,N_3959,N_3113);
and U4549 (N_4549,N_3090,N_3989);
xnor U4550 (N_4550,N_3444,N_3219);
nor U4551 (N_4551,N_3385,N_3211);
and U4552 (N_4552,N_3825,N_3867);
nand U4553 (N_4553,N_3375,N_3457);
nand U4554 (N_4554,N_3702,N_3013);
nand U4555 (N_4555,N_3157,N_3748);
and U4556 (N_4556,N_3628,N_3910);
and U4557 (N_4557,N_3208,N_3348);
nor U4558 (N_4558,N_3947,N_3060);
and U4559 (N_4559,N_3679,N_3890);
nand U4560 (N_4560,N_3098,N_3114);
or U4561 (N_4561,N_3314,N_3014);
nand U4562 (N_4562,N_3009,N_3004);
and U4563 (N_4563,N_3067,N_3441);
or U4564 (N_4564,N_3285,N_3937);
nand U4565 (N_4565,N_3589,N_3990);
and U4566 (N_4566,N_3062,N_3929);
nand U4567 (N_4567,N_3188,N_3212);
nor U4568 (N_4568,N_3237,N_3217);
and U4569 (N_4569,N_3297,N_3624);
and U4570 (N_4570,N_3487,N_3398);
nor U4571 (N_4571,N_3966,N_3605);
nand U4572 (N_4572,N_3343,N_3803);
nor U4573 (N_4573,N_3317,N_3519);
or U4574 (N_4574,N_3717,N_3818);
and U4575 (N_4575,N_3258,N_3429);
and U4576 (N_4576,N_3178,N_3440);
nor U4577 (N_4577,N_3560,N_3495);
nand U4578 (N_4578,N_3076,N_3381);
nand U4579 (N_4579,N_3519,N_3981);
and U4580 (N_4580,N_3798,N_3691);
and U4581 (N_4581,N_3107,N_3019);
or U4582 (N_4582,N_3400,N_3013);
and U4583 (N_4583,N_3383,N_3802);
nor U4584 (N_4584,N_3699,N_3138);
nor U4585 (N_4585,N_3589,N_3437);
and U4586 (N_4586,N_3017,N_3905);
and U4587 (N_4587,N_3082,N_3558);
or U4588 (N_4588,N_3048,N_3538);
nand U4589 (N_4589,N_3224,N_3469);
nand U4590 (N_4590,N_3742,N_3816);
nand U4591 (N_4591,N_3947,N_3841);
or U4592 (N_4592,N_3740,N_3855);
and U4593 (N_4593,N_3423,N_3206);
nor U4594 (N_4594,N_3702,N_3257);
and U4595 (N_4595,N_3369,N_3612);
nor U4596 (N_4596,N_3784,N_3794);
and U4597 (N_4597,N_3718,N_3087);
and U4598 (N_4598,N_3602,N_3082);
or U4599 (N_4599,N_3235,N_3479);
nand U4600 (N_4600,N_3669,N_3150);
and U4601 (N_4601,N_3890,N_3699);
nand U4602 (N_4602,N_3078,N_3066);
and U4603 (N_4603,N_3252,N_3660);
or U4604 (N_4604,N_3607,N_3079);
and U4605 (N_4605,N_3946,N_3709);
and U4606 (N_4606,N_3291,N_3154);
nand U4607 (N_4607,N_3108,N_3758);
and U4608 (N_4608,N_3106,N_3955);
nand U4609 (N_4609,N_3395,N_3444);
and U4610 (N_4610,N_3058,N_3265);
nand U4611 (N_4611,N_3864,N_3174);
or U4612 (N_4612,N_3202,N_3634);
nand U4613 (N_4613,N_3039,N_3155);
and U4614 (N_4614,N_3338,N_3896);
nand U4615 (N_4615,N_3180,N_3177);
nand U4616 (N_4616,N_3268,N_3803);
nor U4617 (N_4617,N_3006,N_3529);
or U4618 (N_4618,N_3175,N_3104);
nand U4619 (N_4619,N_3164,N_3659);
and U4620 (N_4620,N_3064,N_3718);
nand U4621 (N_4621,N_3324,N_3175);
nor U4622 (N_4622,N_3969,N_3498);
or U4623 (N_4623,N_3106,N_3099);
nand U4624 (N_4624,N_3985,N_3066);
or U4625 (N_4625,N_3664,N_3497);
nor U4626 (N_4626,N_3477,N_3499);
nor U4627 (N_4627,N_3560,N_3384);
nand U4628 (N_4628,N_3559,N_3867);
nor U4629 (N_4629,N_3136,N_3786);
and U4630 (N_4630,N_3015,N_3411);
nand U4631 (N_4631,N_3622,N_3162);
nor U4632 (N_4632,N_3407,N_3173);
and U4633 (N_4633,N_3373,N_3694);
nor U4634 (N_4634,N_3251,N_3517);
and U4635 (N_4635,N_3843,N_3596);
nor U4636 (N_4636,N_3482,N_3034);
nor U4637 (N_4637,N_3069,N_3207);
nand U4638 (N_4638,N_3139,N_3150);
or U4639 (N_4639,N_3447,N_3328);
nand U4640 (N_4640,N_3645,N_3285);
nand U4641 (N_4641,N_3448,N_3668);
or U4642 (N_4642,N_3801,N_3165);
nand U4643 (N_4643,N_3822,N_3241);
nand U4644 (N_4644,N_3728,N_3623);
or U4645 (N_4645,N_3651,N_3041);
nand U4646 (N_4646,N_3283,N_3454);
and U4647 (N_4647,N_3576,N_3114);
nand U4648 (N_4648,N_3365,N_3374);
and U4649 (N_4649,N_3928,N_3882);
or U4650 (N_4650,N_3802,N_3170);
nand U4651 (N_4651,N_3152,N_3948);
and U4652 (N_4652,N_3047,N_3322);
nor U4653 (N_4653,N_3654,N_3565);
nand U4654 (N_4654,N_3715,N_3795);
or U4655 (N_4655,N_3009,N_3111);
nand U4656 (N_4656,N_3856,N_3295);
nor U4657 (N_4657,N_3519,N_3309);
and U4658 (N_4658,N_3347,N_3893);
and U4659 (N_4659,N_3120,N_3666);
or U4660 (N_4660,N_3992,N_3595);
nand U4661 (N_4661,N_3815,N_3128);
nor U4662 (N_4662,N_3933,N_3964);
or U4663 (N_4663,N_3127,N_3977);
nand U4664 (N_4664,N_3399,N_3213);
nand U4665 (N_4665,N_3457,N_3136);
nor U4666 (N_4666,N_3994,N_3387);
nor U4667 (N_4667,N_3581,N_3475);
nor U4668 (N_4668,N_3985,N_3182);
or U4669 (N_4669,N_3795,N_3942);
and U4670 (N_4670,N_3402,N_3462);
and U4671 (N_4671,N_3153,N_3313);
or U4672 (N_4672,N_3453,N_3510);
nor U4673 (N_4673,N_3359,N_3262);
nand U4674 (N_4674,N_3431,N_3692);
and U4675 (N_4675,N_3760,N_3095);
nand U4676 (N_4676,N_3705,N_3734);
and U4677 (N_4677,N_3734,N_3366);
nand U4678 (N_4678,N_3641,N_3995);
or U4679 (N_4679,N_3489,N_3864);
or U4680 (N_4680,N_3194,N_3058);
xor U4681 (N_4681,N_3768,N_3003);
nor U4682 (N_4682,N_3508,N_3048);
nor U4683 (N_4683,N_3700,N_3338);
xor U4684 (N_4684,N_3777,N_3480);
nand U4685 (N_4685,N_3803,N_3878);
or U4686 (N_4686,N_3996,N_3745);
nand U4687 (N_4687,N_3600,N_3924);
nand U4688 (N_4688,N_3241,N_3061);
or U4689 (N_4689,N_3080,N_3847);
or U4690 (N_4690,N_3050,N_3152);
and U4691 (N_4691,N_3663,N_3118);
and U4692 (N_4692,N_3825,N_3166);
nor U4693 (N_4693,N_3430,N_3249);
and U4694 (N_4694,N_3556,N_3058);
or U4695 (N_4695,N_3918,N_3735);
nand U4696 (N_4696,N_3099,N_3024);
and U4697 (N_4697,N_3574,N_3894);
or U4698 (N_4698,N_3763,N_3468);
or U4699 (N_4699,N_3323,N_3544);
and U4700 (N_4700,N_3848,N_3324);
nor U4701 (N_4701,N_3764,N_3503);
nor U4702 (N_4702,N_3732,N_3637);
nor U4703 (N_4703,N_3499,N_3934);
nor U4704 (N_4704,N_3425,N_3956);
and U4705 (N_4705,N_3580,N_3991);
and U4706 (N_4706,N_3166,N_3813);
and U4707 (N_4707,N_3027,N_3451);
and U4708 (N_4708,N_3791,N_3034);
nand U4709 (N_4709,N_3443,N_3214);
or U4710 (N_4710,N_3480,N_3812);
nor U4711 (N_4711,N_3501,N_3905);
nor U4712 (N_4712,N_3830,N_3070);
nand U4713 (N_4713,N_3655,N_3307);
nor U4714 (N_4714,N_3491,N_3765);
nand U4715 (N_4715,N_3653,N_3793);
nand U4716 (N_4716,N_3956,N_3973);
or U4717 (N_4717,N_3967,N_3225);
and U4718 (N_4718,N_3840,N_3012);
and U4719 (N_4719,N_3161,N_3239);
and U4720 (N_4720,N_3990,N_3393);
nand U4721 (N_4721,N_3195,N_3977);
nand U4722 (N_4722,N_3026,N_3437);
nand U4723 (N_4723,N_3063,N_3428);
and U4724 (N_4724,N_3734,N_3626);
nor U4725 (N_4725,N_3341,N_3581);
and U4726 (N_4726,N_3599,N_3344);
and U4727 (N_4727,N_3389,N_3074);
nand U4728 (N_4728,N_3218,N_3436);
or U4729 (N_4729,N_3114,N_3205);
nand U4730 (N_4730,N_3612,N_3463);
nand U4731 (N_4731,N_3523,N_3470);
nand U4732 (N_4732,N_3182,N_3444);
nor U4733 (N_4733,N_3405,N_3962);
or U4734 (N_4734,N_3572,N_3795);
nand U4735 (N_4735,N_3873,N_3059);
nand U4736 (N_4736,N_3518,N_3209);
nand U4737 (N_4737,N_3580,N_3980);
or U4738 (N_4738,N_3145,N_3138);
nand U4739 (N_4739,N_3333,N_3201);
nand U4740 (N_4740,N_3963,N_3360);
and U4741 (N_4741,N_3089,N_3202);
or U4742 (N_4742,N_3707,N_3296);
or U4743 (N_4743,N_3478,N_3631);
nand U4744 (N_4744,N_3147,N_3957);
or U4745 (N_4745,N_3689,N_3448);
nor U4746 (N_4746,N_3663,N_3673);
nand U4747 (N_4747,N_3362,N_3479);
nand U4748 (N_4748,N_3242,N_3063);
or U4749 (N_4749,N_3160,N_3351);
or U4750 (N_4750,N_3050,N_3681);
nand U4751 (N_4751,N_3428,N_3821);
nor U4752 (N_4752,N_3140,N_3552);
xor U4753 (N_4753,N_3827,N_3573);
and U4754 (N_4754,N_3108,N_3880);
nor U4755 (N_4755,N_3255,N_3679);
and U4756 (N_4756,N_3681,N_3035);
or U4757 (N_4757,N_3278,N_3172);
nand U4758 (N_4758,N_3567,N_3256);
or U4759 (N_4759,N_3290,N_3552);
or U4760 (N_4760,N_3339,N_3239);
nand U4761 (N_4761,N_3871,N_3656);
nand U4762 (N_4762,N_3175,N_3380);
nand U4763 (N_4763,N_3602,N_3849);
or U4764 (N_4764,N_3033,N_3598);
nor U4765 (N_4765,N_3380,N_3980);
and U4766 (N_4766,N_3100,N_3733);
xnor U4767 (N_4767,N_3159,N_3284);
nand U4768 (N_4768,N_3195,N_3221);
and U4769 (N_4769,N_3109,N_3633);
and U4770 (N_4770,N_3664,N_3843);
nor U4771 (N_4771,N_3268,N_3685);
or U4772 (N_4772,N_3472,N_3315);
or U4773 (N_4773,N_3905,N_3006);
nand U4774 (N_4774,N_3556,N_3375);
and U4775 (N_4775,N_3593,N_3733);
or U4776 (N_4776,N_3183,N_3109);
nor U4777 (N_4777,N_3244,N_3282);
or U4778 (N_4778,N_3458,N_3065);
and U4779 (N_4779,N_3205,N_3287);
or U4780 (N_4780,N_3556,N_3916);
and U4781 (N_4781,N_3506,N_3428);
and U4782 (N_4782,N_3724,N_3516);
nor U4783 (N_4783,N_3427,N_3056);
or U4784 (N_4784,N_3410,N_3626);
or U4785 (N_4785,N_3047,N_3636);
nor U4786 (N_4786,N_3241,N_3529);
and U4787 (N_4787,N_3644,N_3739);
nor U4788 (N_4788,N_3103,N_3097);
or U4789 (N_4789,N_3067,N_3304);
nand U4790 (N_4790,N_3944,N_3509);
xor U4791 (N_4791,N_3748,N_3242);
nor U4792 (N_4792,N_3342,N_3907);
nor U4793 (N_4793,N_3906,N_3736);
and U4794 (N_4794,N_3266,N_3082);
nor U4795 (N_4795,N_3755,N_3080);
nor U4796 (N_4796,N_3091,N_3737);
and U4797 (N_4797,N_3787,N_3347);
nand U4798 (N_4798,N_3865,N_3458);
nor U4799 (N_4799,N_3699,N_3776);
or U4800 (N_4800,N_3300,N_3571);
xnor U4801 (N_4801,N_3300,N_3604);
nand U4802 (N_4802,N_3733,N_3391);
xnor U4803 (N_4803,N_3063,N_3423);
nand U4804 (N_4804,N_3150,N_3831);
nand U4805 (N_4805,N_3349,N_3633);
and U4806 (N_4806,N_3397,N_3720);
nand U4807 (N_4807,N_3800,N_3986);
xnor U4808 (N_4808,N_3628,N_3270);
or U4809 (N_4809,N_3991,N_3217);
and U4810 (N_4810,N_3767,N_3585);
nand U4811 (N_4811,N_3387,N_3094);
and U4812 (N_4812,N_3199,N_3299);
nor U4813 (N_4813,N_3236,N_3592);
nand U4814 (N_4814,N_3782,N_3951);
and U4815 (N_4815,N_3869,N_3106);
nand U4816 (N_4816,N_3358,N_3458);
or U4817 (N_4817,N_3307,N_3244);
or U4818 (N_4818,N_3303,N_3352);
nand U4819 (N_4819,N_3955,N_3316);
or U4820 (N_4820,N_3683,N_3715);
or U4821 (N_4821,N_3845,N_3018);
nand U4822 (N_4822,N_3686,N_3187);
nand U4823 (N_4823,N_3747,N_3763);
nand U4824 (N_4824,N_3349,N_3230);
xnor U4825 (N_4825,N_3951,N_3899);
nor U4826 (N_4826,N_3332,N_3339);
and U4827 (N_4827,N_3211,N_3499);
or U4828 (N_4828,N_3154,N_3708);
or U4829 (N_4829,N_3981,N_3455);
nor U4830 (N_4830,N_3522,N_3664);
nor U4831 (N_4831,N_3879,N_3966);
nand U4832 (N_4832,N_3905,N_3853);
or U4833 (N_4833,N_3371,N_3085);
nor U4834 (N_4834,N_3169,N_3518);
and U4835 (N_4835,N_3075,N_3773);
nand U4836 (N_4836,N_3421,N_3664);
nor U4837 (N_4837,N_3159,N_3554);
and U4838 (N_4838,N_3501,N_3084);
nand U4839 (N_4839,N_3573,N_3911);
and U4840 (N_4840,N_3366,N_3995);
nor U4841 (N_4841,N_3529,N_3703);
nand U4842 (N_4842,N_3299,N_3707);
nand U4843 (N_4843,N_3257,N_3452);
and U4844 (N_4844,N_3186,N_3247);
nor U4845 (N_4845,N_3874,N_3625);
and U4846 (N_4846,N_3197,N_3698);
and U4847 (N_4847,N_3930,N_3305);
or U4848 (N_4848,N_3855,N_3749);
nand U4849 (N_4849,N_3319,N_3458);
nor U4850 (N_4850,N_3503,N_3574);
and U4851 (N_4851,N_3211,N_3836);
nand U4852 (N_4852,N_3798,N_3031);
nor U4853 (N_4853,N_3757,N_3365);
nor U4854 (N_4854,N_3435,N_3051);
nand U4855 (N_4855,N_3295,N_3770);
and U4856 (N_4856,N_3368,N_3993);
and U4857 (N_4857,N_3458,N_3800);
nand U4858 (N_4858,N_3581,N_3180);
or U4859 (N_4859,N_3345,N_3680);
nand U4860 (N_4860,N_3781,N_3088);
and U4861 (N_4861,N_3880,N_3417);
nor U4862 (N_4862,N_3169,N_3685);
nand U4863 (N_4863,N_3569,N_3161);
nand U4864 (N_4864,N_3650,N_3855);
nor U4865 (N_4865,N_3763,N_3429);
and U4866 (N_4866,N_3635,N_3150);
and U4867 (N_4867,N_3501,N_3026);
nor U4868 (N_4868,N_3191,N_3835);
nand U4869 (N_4869,N_3761,N_3790);
nand U4870 (N_4870,N_3335,N_3752);
nand U4871 (N_4871,N_3748,N_3151);
and U4872 (N_4872,N_3707,N_3291);
and U4873 (N_4873,N_3367,N_3827);
nand U4874 (N_4874,N_3868,N_3257);
and U4875 (N_4875,N_3298,N_3020);
or U4876 (N_4876,N_3462,N_3765);
or U4877 (N_4877,N_3605,N_3624);
or U4878 (N_4878,N_3249,N_3989);
or U4879 (N_4879,N_3189,N_3294);
nand U4880 (N_4880,N_3206,N_3809);
or U4881 (N_4881,N_3952,N_3670);
and U4882 (N_4882,N_3491,N_3023);
and U4883 (N_4883,N_3026,N_3209);
nand U4884 (N_4884,N_3215,N_3893);
and U4885 (N_4885,N_3348,N_3173);
and U4886 (N_4886,N_3689,N_3556);
and U4887 (N_4887,N_3970,N_3128);
nand U4888 (N_4888,N_3465,N_3405);
nor U4889 (N_4889,N_3875,N_3499);
nand U4890 (N_4890,N_3651,N_3246);
or U4891 (N_4891,N_3517,N_3615);
and U4892 (N_4892,N_3735,N_3675);
nor U4893 (N_4893,N_3552,N_3979);
nand U4894 (N_4894,N_3168,N_3028);
and U4895 (N_4895,N_3996,N_3843);
nor U4896 (N_4896,N_3883,N_3568);
nor U4897 (N_4897,N_3518,N_3184);
and U4898 (N_4898,N_3296,N_3885);
nor U4899 (N_4899,N_3368,N_3862);
nand U4900 (N_4900,N_3513,N_3289);
and U4901 (N_4901,N_3173,N_3413);
and U4902 (N_4902,N_3872,N_3223);
and U4903 (N_4903,N_3366,N_3294);
and U4904 (N_4904,N_3153,N_3705);
and U4905 (N_4905,N_3902,N_3097);
or U4906 (N_4906,N_3806,N_3345);
nand U4907 (N_4907,N_3518,N_3780);
nor U4908 (N_4908,N_3469,N_3561);
and U4909 (N_4909,N_3393,N_3881);
nand U4910 (N_4910,N_3198,N_3641);
nand U4911 (N_4911,N_3576,N_3610);
xor U4912 (N_4912,N_3075,N_3533);
and U4913 (N_4913,N_3575,N_3436);
nand U4914 (N_4914,N_3922,N_3032);
nand U4915 (N_4915,N_3606,N_3073);
nor U4916 (N_4916,N_3047,N_3095);
or U4917 (N_4917,N_3510,N_3428);
and U4918 (N_4918,N_3393,N_3953);
nand U4919 (N_4919,N_3008,N_3581);
and U4920 (N_4920,N_3020,N_3611);
nand U4921 (N_4921,N_3276,N_3562);
nand U4922 (N_4922,N_3178,N_3964);
and U4923 (N_4923,N_3267,N_3347);
nand U4924 (N_4924,N_3353,N_3250);
nor U4925 (N_4925,N_3069,N_3567);
nor U4926 (N_4926,N_3649,N_3789);
and U4927 (N_4927,N_3836,N_3006);
nor U4928 (N_4928,N_3186,N_3705);
or U4929 (N_4929,N_3156,N_3927);
nand U4930 (N_4930,N_3727,N_3255);
nand U4931 (N_4931,N_3494,N_3723);
nand U4932 (N_4932,N_3934,N_3645);
nor U4933 (N_4933,N_3619,N_3560);
nor U4934 (N_4934,N_3158,N_3742);
nor U4935 (N_4935,N_3984,N_3893);
nand U4936 (N_4936,N_3625,N_3041);
or U4937 (N_4937,N_3793,N_3977);
nand U4938 (N_4938,N_3253,N_3024);
and U4939 (N_4939,N_3573,N_3477);
and U4940 (N_4940,N_3103,N_3203);
nor U4941 (N_4941,N_3425,N_3318);
and U4942 (N_4942,N_3222,N_3445);
nor U4943 (N_4943,N_3977,N_3874);
nor U4944 (N_4944,N_3116,N_3086);
nor U4945 (N_4945,N_3246,N_3563);
or U4946 (N_4946,N_3880,N_3302);
or U4947 (N_4947,N_3797,N_3117);
or U4948 (N_4948,N_3225,N_3834);
xnor U4949 (N_4949,N_3169,N_3830);
and U4950 (N_4950,N_3495,N_3105);
nand U4951 (N_4951,N_3349,N_3739);
and U4952 (N_4952,N_3437,N_3343);
nand U4953 (N_4953,N_3207,N_3812);
or U4954 (N_4954,N_3703,N_3425);
nand U4955 (N_4955,N_3809,N_3662);
or U4956 (N_4956,N_3061,N_3696);
nor U4957 (N_4957,N_3978,N_3419);
or U4958 (N_4958,N_3325,N_3796);
nand U4959 (N_4959,N_3326,N_3495);
or U4960 (N_4960,N_3339,N_3592);
nor U4961 (N_4961,N_3797,N_3447);
and U4962 (N_4962,N_3941,N_3041);
nor U4963 (N_4963,N_3547,N_3839);
or U4964 (N_4964,N_3230,N_3196);
and U4965 (N_4965,N_3291,N_3715);
nand U4966 (N_4966,N_3498,N_3160);
and U4967 (N_4967,N_3972,N_3040);
and U4968 (N_4968,N_3080,N_3575);
nand U4969 (N_4969,N_3487,N_3925);
or U4970 (N_4970,N_3624,N_3572);
and U4971 (N_4971,N_3235,N_3015);
and U4972 (N_4972,N_3890,N_3715);
nor U4973 (N_4973,N_3067,N_3390);
or U4974 (N_4974,N_3780,N_3753);
nor U4975 (N_4975,N_3186,N_3765);
or U4976 (N_4976,N_3304,N_3895);
nor U4977 (N_4977,N_3692,N_3005);
or U4978 (N_4978,N_3942,N_3698);
and U4979 (N_4979,N_3596,N_3061);
nand U4980 (N_4980,N_3088,N_3562);
or U4981 (N_4981,N_3918,N_3851);
and U4982 (N_4982,N_3953,N_3699);
nor U4983 (N_4983,N_3461,N_3165);
nand U4984 (N_4984,N_3860,N_3487);
nand U4985 (N_4985,N_3040,N_3019);
xor U4986 (N_4986,N_3744,N_3300);
xnor U4987 (N_4987,N_3243,N_3451);
nand U4988 (N_4988,N_3231,N_3861);
nand U4989 (N_4989,N_3464,N_3656);
and U4990 (N_4990,N_3919,N_3541);
nand U4991 (N_4991,N_3656,N_3541);
or U4992 (N_4992,N_3076,N_3942);
and U4993 (N_4993,N_3666,N_3925);
nand U4994 (N_4994,N_3139,N_3582);
nand U4995 (N_4995,N_3105,N_3426);
xnor U4996 (N_4996,N_3094,N_3160);
and U4997 (N_4997,N_3882,N_3711);
and U4998 (N_4998,N_3537,N_3324);
nand U4999 (N_4999,N_3332,N_3996);
and UO_0 (O_0,N_4942,N_4578);
nor UO_1 (O_1,N_4298,N_4699);
or UO_2 (O_2,N_4005,N_4713);
or UO_3 (O_3,N_4488,N_4585);
nand UO_4 (O_4,N_4231,N_4099);
and UO_5 (O_5,N_4160,N_4893);
nand UO_6 (O_6,N_4588,N_4110);
and UO_7 (O_7,N_4093,N_4692);
nor UO_8 (O_8,N_4233,N_4626);
nor UO_9 (O_9,N_4218,N_4153);
and UO_10 (O_10,N_4994,N_4470);
and UO_11 (O_11,N_4234,N_4752);
nor UO_12 (O_12,N_4696,N_4781);
nor UO_13 (O_13,N_4611,N_4187);
nand UO_14 (O_14,N_4712,N_4569);
nor UO_15 (O_15,N_4982,N_4675);
and UO_16 (O_16,N_4481,N_4587);
nand UO_17 (O_17,N_4865,N_4209);
nand UO_18 (O_18,N_4782,N_4991);
nand UO_19 (O_19,N_4715,N_4315);
and UO_20 (O_20,N_4274,N_4076);
nand UO_21 (O_21,N_4156,N_4592);
nand UO_22 (O_22,N_4235,N_4911);
or UO_23 (O_23,N_4284,N_4571);
nand UO_24 (O_24,N_4908,N_4624);
or UO_25 (O_25,N_4538,N_4902);
or UO_26 (O_26,N_4743,N_4053);
or UO_27 (O_27,N_4772,N_4402);
nor UO_28 (O_28,N_4331,N_4679);
and UO_29 (O_29,N_4472,N_4547);
and UO_30 (O_30,N_4030,N_4293);
nor UO_31 (O_31,N_4381,N_4338);
and UO_32 (O_32,N_4168,N_4410);
nor UO_33 (O_33,N_4997,N_4213);
nor UO_34 (O_34,N_4098,N_4129);
and UO_35 (O_35,N_4403,N_4535);
or UO_36 (O_36,N_4738,N_4707);
xor UO_37 (O_37,N_4385,N_4066);
or UO_38 (O_38,N_4482,N_4075);
nand UO_39 (O_39,N_4924,N_4716);
nor UO_40 (O_40,N_4255,N_4515);
nor UO_41 (O_41,N_4246,N_4122);
nand UO_42 (O_42,N_4673,N_4605);
nand UO_43 (O_43,N_4217,N_4828);
nand UO_44 (O_44,N_4623,N_4064);
and UO_45 (O_45,N_4121,N_4379);
nor UO_46 (O_46,N_4377,N_4662);
nand UO_47 (O_47,N_4471,N_4559);
nor UO_48 (O_48,N_4469,N_4017);
and UO_49 (O_49,N_4989,N_4349);
nand UO_50 (O_50,N_4111,N_4748);
and UO_51 (O_51,N_4775,N_4404);
and UO_52 (O_52,N_4874,N_4895);
and UO_53 (O_53,N_4764,N_4549);
nor UO_54 (O_54,N_4340,N_4645);
nor UO_55 (O_55,N_4706,N_4632);
or UO_56 (O_56,N_4583,N_4146);
nor UO_57 (O_57,N_4079,N_4357);
and UO_58 (O_58,N_4910,N_4984);
and UO_59 (O_59,N_4789,N_4013);
nor UO_60 (O_60,N_4746,N_4964);
nor UO_61 (O_61,N_4452,N_4334);
or UO_62 (O_62,N_4616,N_4307);
nor UO_63 (O_63,N_4540,N_4629);
or UO_64 (O_64,N_4508,N_4926);
xnor UO_65 (O_65,N_4963,N_4424);
and UO_66 (O_66,N_4308,N_4837);
nand UO_67 (O_67,N_4207,N_4344);
and UO_68 (O_68,N_4798,N_4072);
or UO_69 (O_69,N_4316,N_4799);
xor UO_70 (O_70,N_4220,N_4126);
or UO_71 (O_71,N_4631,N_4788);
or UO_72 (O_72,N_4769,N_4498);
nand UO_73 (O_73,N_4822,N_4787);
nor UO_74 (O_74,N_4790,N_4195);
nor UO_75 (O_75,N_4130,N_4722);
nand UO_76 (O_76,N_4408,N_4271);
nor UO_77 (O_77,N_4650,N_4318);
nor UO_78 (O_78,N_4557,N_4927);
nand UO_79 (O_79,N_4528,N_4827);
nand UO_80 (O_80,N_4674,N_4177);
nand UO_81 (O_81,N_4336,N_4805);
nand UO_82 (O_82,N_4959,N_4918);
nand UO_83 (O_83,N_4561,N_4347);
and UO_84 (O_84,N_4023,N_4586);
and UO_85 (O_85,N_4247,N_4916);
nand UO_86 (O_86,N_4158,N_4059);
nor UO_87 (O_87,N_4229,N_4485);
or UO_88 (O_88,N_4483,N_4152);
and UO_89 (O_89,N_4800,N_4427);
nor UO_90 (O_90,N_4905,N_4061);
nor UO_91 (O_91,N_4714,N_4128);
nor UO_92 (O_92,N_4568,N_4060);
nand UO_93 (O_93,N_4590,N_4765);
or UO_94 (O_94,N_4957,N_4845);
nor UO_95 (O_95,N_4572,N_4194);
and UO_96 (O_96,N_4411,N_4056);
or UO_97 (O_97,N_4296,N_4660);
or UO_98 (O_98,N_4543,N_4007);
or UO_99 (O_99,N_4425,N_4178);
or UO_100 (O_100,N_4197,N_4343);
nor UO_101 (O_101,N_4371,N_4439);
nand UO_102 (O_102,N_4795,N_4533);
nand UO_103 (O_103,N_4232,N_4812);
and UO_104 (O_104,N_4850,N_4420);
nand UO_105 (O_105,N_4655,N_4857);
xnor UO_106 (O_106,N_4548,N_4763);
or UO_107 (O_107,N_4758,N_4906);
or UO_108 (O_108,N_4323,N_4433);
xor UO_109 (O_109,N_4211,N_4725);
and UO_110 (O_110,N_4443,N_4943);
or UO_111 (O_111,N_4651,N_4843);
nor UO_112 (O_112,N_4269,N_4816);
or UO_113 (O_113,N_4573,N_4328);
nand UO_114 (O_114,N_4505,N_4929);
or UO_115 (O_115,N_4976,N_4859);
nor UO_116 (O_116,N_4406,N_4276);
and UO_117 (O_117,N_4380,N_4742);
or UO_118 (O_118,N_4025,N_4045);
nand UO_119 (O_119,N_4301,N_4095);
and UO_120 (O_120,N_4806,N_4001);
nor UO_121 (O_121,N_4495,N_4200);
or UO_122 (O_122,N_4346,N_4360);
or UO_123 (O_123,N_4051,N_4074);
nand UO_124 (O_124,N_4201,N_4821);
nand UO_125 (O_125,N_4777,N_4219);
nor UO_126 (O_126,N_4412,N_4484);
or UO_127 (O_127,N_4441,N_4419);
and UO_128 (O_128,N_4574,N_4283);
nor UO_129 (O_129,N_4449,N_4981);
nor UO_130 (O_130,N_4191,N_4394);
and UO_131 (O_131,N_4919,N_4034);
and UO_132 (O_132,N_4831,N_4182);
nand UO_133 (O_133,N_4672,N_4398);
and UO_134 (O_134,N_4496,N_4175);
nand UO_135 (O_135,N_4597,N_4966);
nand UO_136 (O_136,N_4652,N_4909);
nor UO_137 (O_137,N_4251,N_4181);
or UO_138 (O_138,N_4387,N_4912);
and UO_139 (O_139,N_4878,N_4575);
or UO_140 (O_140,N_4526,N_4008);
or UO_141 (O_141,N_4148,N_4949);
nor UO_142 (O_142,N_4103,N_4451);
and UO_143 (O_143,N_4024,N_4581);
and UO_144 (O_144,N_4286,N_4537);
nor UO_145 (O_145,N_4029,N_4305);
or UO_146 (O_146,N_4500,N_4407);
or UO_147 (O_147,N_4796,N_4507);
and UO_148 (O_148,N_4084,N_4241);
or UO_149 (O_149,N_4872,N_4206);
nor UO_150 (O_150,N_4198,N_4820);
xor UO_151 (O_151,N_4304,N_4825);
or UO_152 (O_152,N_4445,N_4599);
and UO_153 (O_153,N_4958,N_4396);
nand UO_154 (O_154,N_4009,N_4999);
nor UO_155 (O_155,N_4657,N_4116);
and UO_156 (O_156,N_4117,N_4313);
and UO_157 (O_157,N_4506,N_4889);
and UO_158 (O_158,N_4460,N_4524);
nand UO_159 (O_159,N_4087,N_4238);
nand UO_160 (O_160,N_4532,N_4311);
and UO_161 (O_161,N_4431,N_4159);
or UO_162 (O_162,N_4339,N_4973);
and UO_163 (O_163,N_4539,N_4466);
nor UO_164 (O_164,N_4409,N_4327);
or UO_165 (O_165,N_4974,N_4118);
and UO_166 (O_166,N_4421,N_4904);
nand UO_167 (O_167,N_4648,N_4570);
and UO_168 (O_168,N_4179,N_4998);
or UO_169 (O_169,N_4925,N_4915);
and UO_170 (O_170,N_4279,N_4886);
xnor UO_171 (O_171,N_4668,N_4511);
and UO_172 (O_172,N_4851,N_4979);
nand UO_173 (O_173,N_4711,N_4267);
xnor UO_174 (O_174,N_4747,N_4726);
or UO_175 (O_175,N_4069,N_4317);
nor UO_176 (O_176,N_4996,N_4047);
nand UO_177 (O_177,N_4840,N_4803);
and UO_178 (O_178,N_4914,N_4202);
nor UO_179 (O_179,N_4666,N_4686);
nand UO_180 (O_180,N_4643,N_4947);
nand UO_181 (O_181,N_4576,N_4667);
nor UO_182 (O_182,N_4205,N_4480);
or UO_183 (O_183,N_4169,N_4444);
and UO_184 (O_184,N_4326,N_4355);
nor UO_185 (O_185,N_4625,N_4123);
nor UO_186 (O_186,N_4642,N_4085);
nand UO_187 (O_187,N_4373,N_4395);
or UO_188 (O_188,N_4939,N_4455);
or UO_189 (O_189,N_4767,N_4804);
nand UO_190 (O_190,N_4456,N_4734);
nor UO_191 (O_191,N_4504,N_4598);
or UO_192 (O_192,N_4223,N_4518);
or UO_193 (O_193,N_4855,N_4290);
and UO_194 (O_194,N_4002,N_4617);
nor UO_195 (O_195,N_4553,N_4832);
and UO_196 (O_196,N_4577,N_4397);
xnor UO_197 (O_197,N_4312,N_4501);
nand UO_198 (O_198,N_4432,N_4216);
and UO_199 (O_199,N_4704,N_4468);
or UO_200 (O_200,N_4491,N_4695);
or UO_201 (O_201,N_4558,N_4006);
nand UO_202 (O_202,N_4759,N_4188);
nor UO_203 (O_203,N_4353,N_4813);
and UO_204 (O_204,N_4442,N_4913);
or UO_205 (O_205,N_4644,N_4771);
nor UO_206 (O_206,N_4817,N_4281);
nand UO_207 (O_207,N_4094,N_4386);
nand UO_208 (O_208,N_4603,N_4310);
or UO_209 (O_209,N_4661,N_4363);
nand UO_210 (O_210,N_4658,N_4049);
and UO_211 (O_211,N_4426,N_4883);
and UO_212 (O_212,N_4950,N_4114);
nor UO_213 (O_213,N_4151,N_4749);
and UO_214 (O_214,N_4278,N_4641);
and UO_215 (O_215,N_4448,N_4729);
and UO_216 (O_216,N_4751,N_4523);
and UO_217 (O_217,N_4978,N_4091);
and UO_218 (O_218,N_4709,N_4776);
nor UO_219 (O_219,N_4719,N_4727);
and UO_220 (O_220,N_4541,N_4280);
nor UO_221 (O_221,N_4635,N_4299);
or UO_222 (O_222,N_4522,N_4415);
and UO_223 (O_223,N_4436,N_4842);
or UO_224 (O_224,N_4378,N_4778);
nor UO_225 (O_225,N_4733,N_4294);
nand UO_226 (O_226,N_4760,N_4637);
nand UO_227 (O_227,N_4627,N_4591);
nand UO_228 (O_228,N_4113,N_4794);
nand UO_229 (O_229,N_4184,N_4208);
and UO_230 (O_230,N_4614,N_4766);
and UO_231 (O_231,N_4730,N_4423);
nand UO_232 (O_232,N_4613,N_4601);
nand UO_233 (O_233,N_4262,N_4602);
nor UO_234 (O_234,N_4042,N_4365);
or UO_235 (O_235,N_4435,N_4221);
xor UO_236 (O_236,N_4993,N_4291);
nor UO_237 (O_237,N_4065,N_4165);
and UO_238 (O_238,N_4161,N_4604);
nor UO_239 (O_239,N_4309,N_4544);
or UO_240 (O_240,N_4853,N_4043);
nor UO_241 (O_241,N_4885,N_4285);
nor UO_242 (O_242,N_4057,N_4362);
nor UO_243 (O_243,N_4653,N_4938);
and UO_244 (O_244,N_4254,N_4955);
or UO_245 (O_245,N_4761,N_4698);
nand UO_246 (O_246,N_4757,N_4936);
nand UO_247 (O_247,N_4384,N_4849);
and UO_248 (O_248,N_4887,N_4756);
and UO_249 (O_249,N_4054,N_4870);
nand UO_250 (O_250,N_4487,N_4639);
or UO_251 (O_251,N_4401,N_4854);
and UO_252 (O_252,N_4622,N_4345);
or UO_253 (O_253,N_4277,N_4050);
nor UO_254 (O_254,N_4860,N_4871);
and UO_255 (O_255,N_4325,N_4021);
and UO_256 (O_256,N_4941,N_4606);
and UO_257 (O_257,N_4131,N_4154);
nor UO_258 (O_258,N_4633,N_4615);
nand UO_259 (O_259,N_4582,N_4295);
or UO_260 (O_260,N_4830,N_4257);
or UO_261 (O_261,N_4492,N_4961);
and UO_262 (O_262,N_4237,N_4392);
or UO_263 (O_263,N_4768,N_4770);
and UO_264 (O_264,N_4917,N_4732);
or UO_265 (O_265,N_4684,N_4628);
and UO_266 (O_266,N_4434,N_4741);
nor UO_267 (O_267,N_4861,N_4186);
nand UO_268 (O_268,N_4493,N_4882);
or UO_269 (O_269,N_4928,N_4092);
and UO_270 (O_270,N_4027,N_4429);
nor UO_271 (O_271,N_4676,N_4096);
nor UO_272 (O_272,N_4980,N_4088);
nand UO_273 (O_273,N_4951,N_4896);
nand UO_274 (O_274,N_4171,N_4516);
or UO_275 (O_275,N_4070,N_4841);
xor UO_276 (O_276,N_4203,N_4888);
or UO_277 (O_277,N_4105,N_4473);
nand UO_278 (O_278,N_4869,N_4400);
and UO_279 (O_279,N_4721,N_4527);
nor UO_280 (O_280,N_4014,N_4608);
or UO_281 (O_281,N_4133,N_4596);
or UO_282 (O_282,N_4440,N_4962);
xor UO_283 (O_283,N_4785,N_4900);
nor UO_284 (O_284,N_4971,N_4112);
or UO_285 (O_285,N_4986,N_4724);
or UO_286 (O_286,N_4248,N_4697);
and UO_287 (O_287,N_4731,N_4335);
or UO_288 (O_288,N_4370,N_4367);
or UO_289 (O_289,N_4879,N_4529);
and UO_290 (O_290,N_4120,N_4214);
or UO_291 (O_291,N_4352,N_4249);
or UO_292 (O_292,N_4953,N_4282);
and UO_293 (O_293,N_4867,N_4819);
and UO_294 (O_294,N_4933,N_4322);
nor UO_295 (O_295,N_4856,N_4797);
nand UO_296 (O_296,N_4791,N_4227);
and UO_297 (O_297,N_4802,N_4801);
xnor UO_298 (O_298,N_4382,N_4478);
or UO_299 (O_299,N_4147,N_4058);
and UO_300 (O_300,N_4173,N_4985);
xor UO_301 (O_301,N_4166,N_4204);
and UO_302 (O_302,N_4369,N_4467);
nor UO_303 (O_303,N_4388,N_4881);
and UO_304 (O_304,N_4390,N_4636);
or UO_305 (O_305,N_4475,N_4236);
or UO_306 (O_306,N_4612,N_4620);
or UO_307 (O_307,N_4640,N_4517);
nor UO_308 (O_308,N_4509,N_4052);
nand UO_309 (O_309,N_4580,N_4836);
nor UO_310 (O_310,N_4261,N_4245);
or UO_311 (O_311,N_4454,N_4786);
nand UO_312 (O_312,N_4755,N_4863);
and UO_313 (O_313,N_4563,N_4302);
xor UO_314 (O_314,N_4946,N_4036);
nor UO_315 (O_315,N_4844,N_4144);
nand UO_316 (O_316,N_4319,N_4225);
or UO_317 (O_317,N_4081,N_4497);
xor UO_318 (O_318,N_4474,N_4512);
nor UO_319 (O_319,N_4710,N_4104);
or UO_320 (O_320,N_4273,N_4534);
and UO_321 (O_321,N_4864,N_4383);
nor UO_322 (O_322,N_4372,N_4807);
nand UO_323 (O_323,N_4551,N_4546);
nand UO_324 (O_324,N_4438,N_4391);
nor UO_325 (O_325,N_4735,N_4359);
nand UO_326 (O_326,N_4048,N_4647);
or UO_327 (O_327,N_4969,N_4368);
nand UO_328 (O_328,N_4150,N_4170);
nand UO_329 (O_329,N_4965,N_4135);
nand UO_330 (O_330,N_4422,N_4514);
xor UO_331 (O_331,N_4073,N_4450);
nand UO_332 (O_332,N_4649,N_4185);
or UO_333 (O_333,N_4068,N_4823);
or UO_334 (O_334,N_4162,N_4172);
and UO_335 (O_335,N_4341,N_4808);
nor UO_336 (O_336,N_4366,N_4477);
nand UO_337 (O_337,N_4677,N_4320);
and UO_338 (O_338,N_4619,N_4654);
and UO_339 (O_339,N_4693,N_4288);
and UO_340 (O_340,N_4503,N_4463);
or UO_341 (O_341,N_4780,N_4189);
xnor UO_342 (O_342,N_4810,N_4015);
and UO_343 (O_343,N_4809,N_4826);
or UO_344 (O_344,N_4884,N_4321);
or UO_345 (O_345,N_4228,N_4145);
nor UO_346 (O_346,N_4708,N_4554);
or UO_347 (O_347,N_4545,N_4664);
nand UO_348 (O_348,N_4824,N_4499);
nand UO_349 (O_349,N_4656,N_4934);
nand UO_350 (O_350,N_4164,N_4155);
xnor UO_351 (O_351,N_4931,N_4089);
nor UO_352 (O_352,N_4354,N_4174);
or UO_353 (O_353,N_4740,N_4289);
nor UO_354 (O_354,N_4055,N_4106);
and UO_355 (O_355,N_4681,N_4413);
nor UO_356 (O_356,N_4020,N_4897);
or UO_357 (O_357,N_4678,N_4705);
nor UO_358 (O_358,N_4258,N_4292);
or UO_359 (O_359,N_4125,N_4838);
nand UO_360 (O_360,N_4811,N_4264);
nor UO_361 (O_361,N_4944,N_4519);
or UO_362 (O_362,N_4250,N_4542);
and UO_363 (O_363,N_4035,N_4784);
nand UO_364 (O_364,N_4031,N_4244);
or UO_365 (O_365,N_4132,N_4903);
nor UO_366 (O_366,N_4920,N_4670);
nand UO_367 (O_367,N_4930,N_4361);
nor UO_368 (O_368,N_4364,N_4521);
or UO_369 (O_369,N_4907,N_4922);
nand UO_370 (O_370,N_4399,N_4453);
or UO_371 (O_371,N_4960,N_4242);
nor UO_372 (O_372,N_4314,N_4037);
or UO_373 (O_373,N_4138,N_4531);
nor UO_374 (O_374,N_4038,N_4935);
and UO_375 (O_375,N_4040,N_4489);
and UO_376 (O_376,N_4252,N_4659);
or UO_377 (O_377,N_4945,N_4003);
and UO_378 (O_378,N_4536,N_4987);
or UO_379 (O_379,N_4875,N_4691);
or UO_380 (O_380,N_4330,N_4193);
nand UO_381 (O_381,N_4479,N_4595);
or UO_382 (O_382,N_4418,N_4028);
or UO_383 (O_383,N_4215,N_4033);
nor UO_384 (O_384,N_4899,N_4921);
or UO_385 (O_385,N_4901,N_4848);
or UO_386 (O_386,N_4892,N_4101);
or UO_387 (O_387,N_4259,N_4891);
nand UO_388 (O_388,N_4090,N_4968);
and UO_389 (O_389,N_4461,N_4967);
and UO_390 (O_390,N_4011,N_4833);
nor UO_391 (O_391,N_4665,N_4119);
and UO_392 (O_392,N_4745,N_4952);
and UO_393 (O_393,N_4815,N_4376);
and UO_394 (O_394,N_4513,N_4067);
xor UO_395 (O_395,N_4062,N_4701);
nand UO_396 (O_396,N_4127,N_4846);
or UO_397 (O_397,N_4723,N_4877);
nor UO_398 (O_398,N_4039,N_4222);
or UO_399 (O_399,N_4995,N_4212);
nor UO_400 (O_400,N_4753,N_4555);
and UO_401 (O_401,N_4682,N_4004);
nor UO_402 (O_402,N_4032,N_4703);
or UO_403 (O_403,N_4898,N_4562);
and UO_404 (O_404,N_4638,N_4275);
nor UO_405 (O_405,N_4022,N_4263);
nand UO_406 (O_406,N_4356,N_4970);
and UO_407 (O_407,N_4063,N_4272);
and UO_408 (O_408,N_4688,N_4773);
nor UO_409 (O_409,N_4685,N_4683);
or UO_410 (O_410,N_4550,N_4476);
nand UO_411 (O_411,N_4016,N_4520);
nor UO_412 (O_412,N_4983,N_4071);
nand UO_413 (O_413,N_4607,N_4502);
nand UO_414 (O_414,N_4754,N_4097);
or UO_415 (O_415,N_4894,N_4876);
nand UO_416 (O_416,N_4630,N_4142);
and UO_417 (O_417,N_4634,N_4306);
nor UO_418 (O_418,N_4702,N_4600);
and UO_419 (O_419,N_4124,N_4010);
nor UO_420 (O_420,N_4115,N_4416);
nor UO_421 (O_421,N_4937,N_4814);
nand UO_422 (O_422,N_4457,N_4462);
nor UO_423 (O_423,N_4584,N_4694);
or UO_424 (O_424,N_4265,N_4866);
and UO_425 (O_425,N_4774,N_4744);
nor UO_426 (O_426,N_4083,N_4680);
or UO_427 (O_427,N_4486,N_4720);
or UO_428 (O_428,N_4890,N_4226);
nand UO_429 (O_429,N_4190,N_4167);
nand UO_430 (O_430,N_4082,N_4210);
and UO_431 (O_431,N_4552,N_4972);
nor UO_432 (O_432,N_4077,N_4134);
and UO_433 (O_433,N_4332,N_4078);
nand UO_434 (O_434,N_4337,N_4046);
or UO_435 (O_435,N_4779,N_4464);
nor UO_436 (O_436,N_4988,N_4000);
or UO_437 (O_437,N_4762,N_4593);
or UO_438 (O_438,N_4646,N_4405);
nor UO_439 (O_439,N_4829,N_4287);
xor UO_440 (O_440,N_4447,N_4621);
or UO_441 (O_441,N_4932,N_4260);
nor UO_442 (O_442,N_4862,N_4792);
nor UO_443 (O_443,N_4737,N_4333);
nand UO_444 (O_444,N_4375,N_4510);
and UO_445 (O_445,N_4589,N_4149);
nand UO_446 (O_446,N_4736,N_4564);
nand UO_447 (O_447,N_4728,N_4618);
or UO_448 (O_448,N_4414,N_4012);
or UO_449 (O_449,N_4300,N_4610);
or UO_450 (O_450,N_4256,N_4358);
nand UO_451 (O_451,N_4530,N_4137);
nand UO_452 (O_452,N_4109,N_4609);
nand UO_453 (O_453,N_4954,N_4858);
nor UO_454 (O_454,N_4270,N_4818);
nand UO_455 (O_455,N_4793,N_4224);
and UO_456 (O_456,N_4690,N_4977);
nand UO_457 (O_457,N_4240,N_4107);
and UO_458 (O_458,N_4835,N_4992);
and UO_459 (O_459,N_4556,N_4230);
and UO_460 (O_460,N_4239,N_4393);
or UO_461 (O_461,N_4750,N_4594);
and UO_462 (O_462,N_4975,N_4689);
and UO_463 (O_463,N_4348,N_4739);
and UO_464 (O_464,N_4417,N_4044);
nor UO_465 (O_465,N_4140,N_4663);
or UO_466 (O_466,N_4566,N_4183);
or UO_467 (O_467,N_4100,N_4342);
nor UO_468 (O_468,N_4428,N_4266);
nor UO_469 (O_469,N_4446,N_4163);
or UO_470 (O_470,N_4847,N_4852);
or UO_471 (O_471,N_4437,N_4136);
or UO_472 (O_472,N_4687,N_4199);
and UO_473 (O_473,N_4303,N_4297);
nor UO_474 (O_474,N_4180,N_4565);
nor UO_475 (O_475,N_4880,N_4868);
or UO_476 (O_476,N_4459,N_4923);
nand UO_477 (O_477,N_4026,N_4329);
nor UO_478 (O_478,N_4157,N_4243);
xnor UO_479 (O_479,N_4041,N_4430);
or UO_480 (O_480,N_4494,N_4834);
nor UO_481 (O_481,N_4176,N_4490);
or UO_482 (O_482,N_4839,N_4192);
and UO_483 (O_483,N_4700,N_4948);
nor UO_484 (O_484,N_4669,N_4143);
nand UO_485 (O_485,N_4873,N_4956);
or UO_486 (O_486,N_4324,N_4018);
nand UO_487 (O_487,N_4374,N_4458);
and UO_488 (O_488,N_4351,N_4086);
nand UO_489 (O_489,N_4525,N_4389);
nor UO_490 (O_490,N_4567,N_4268);
or UO_491 (O_491,N_4465,N_4139);
nand UO_492 (O_492,N_4671,N_4102);
nand UO_493 (O_493,N_4990,N_4108);
and UO_494 (O_494,N_4579,N_4350);
or UO_495 (O_495,N_4560,N_4080);
nand UO_496 (O_496,N_4253,N_4940);
and UO_497 (O_497,N_4717,N_4718);
and UO_498 (O_498,N_4196,N_4141);
nor UO_499 (O_499,N_4783,N_4019);
nor UO_500 (O_500,N_4048,N_4966);
nand UO_501 (O_501,N_4036,N_4075);
nor UO_502 (O_502,N_4356,N_4416);
and UO_503 (O_503,N_4944,N_4404);
or UO_504 (O_504,N_4032,N_4493);
nand UO_505 (O_505,N_4144,N_4593);
or UO_506 (O_506,N_4737,N_4257);
or UO_507 (O_507,N_4201,N_4892);
and UO_508 (O_508,N_4122,N_4407);
nor UO_509 (O_509,N_4992,N_4659);
nand UO_510 (O_510,N_4898,N_4802);
and UO_511 (O_511,N_4349,N_4139);
and UO_512 (O_512,N_4179,N_4523);
and UO_513 (O_513,N_4923,N_4127);
nor UO_514 (O_514,N_4486,N_4866);
and UO_515 (O_515,N_4333,N_4235);
nand UO_516 (O_516,N_4403,N_4039);
and UO_517 (O_517,N_4542,N_4686);
or UO_518 (O_518,N_4026,N_4503);
nor UO_519 (O_519,N_4920,N_4402);
nor UO_520 (O_520,N_4756,N_4835);
and UO_521 (O_521,N_4602,N_4737);
nand UO_522 (O_522,N_4174,N_4357);
nand UO_523 (O_523,N_4070,N_4324);
and UO_524 (O_524,N_4460,N_4196);
or UO_525 (O_525,N_4659,N_4959);
nand UO_526 (O_526,N_4485,N_4805);
or UO_527 (O_527,N_4444,N_4975);
nor UO_528 (O_528,N_4901,N_4923);
nand UO_529 (O_529,N_4100,N_4666);
nand UO_530 (O_530,N_4316,N_4397);
nor UO_531 (O_531,N_4124,N_4601);
nor UO_532 (O_532,N_4844,N_4807);
nor UO_533 (O_533,N_4829,N_4922);
nor UO_534 (O_534,N_4944,N_4766);
or UO_535 (O_535,N_4058,N_4321);
or UO_536 (O_536,N_4965,N_4485);
nor UO_537 (O_537,N_4991,N_4896);
or UO_538 (O_538,N_4090,N_4333);
nand UO_539 (O_539,N_4351,N_4012);
and UO_540 (O_540,N_4187,N_4785);
and UO_541 (O_541,N_4999,N_4359);
and UO_542 (O_542,N_4916,N_4061);
and UO_543 (O_543,N_4767,N_4204);
or UO_544 (O_544,N_4372,N_4123);
nand UO_545 (O_545,N_4657,N_4395);
nand UO_546 (O_546,N_4660,N_4604);
nor UO_547 (O_547,N_4783,N_4184);
nor UO_548 (O_548,N_4234,N_4406);
nor UO_549 (O_549,N_4869,N_4842);
nor UO_550 (O_550,N_4690,N_4100);
and UO_551 (O_551,N_4681,N_4772);
and UO_552 (O_552,N_4580,N_4817);
xor UO_553 (O_553,N_4894,N_4955);
nand UO_554 (O_554,N_4736,N_4551);
and UO_555 (O_555,N_4410,N_4210);
nand UO_556 (O_556,N_4024,N_4773);
and UO_557 (O_557,N_4748,N_4817);
and UO_558 (O_558,N_4046,N_4596);
nor UO_559 (O_559,N_4417,N_4024);
and UO_560 (O_560,N_4552,N_4305);
nor UO_561 (O_561,N_4766,N_4680);
or UO_562 (O_562,N_4904,N_4519);
or UO_563 (O_563,N_4373,N_4448);
nand UO_564 (O_564,N_4378,N_4176);
nor UO_565 (O_565,N_4779,N_4062);
nor UO_566 (O_566,N_4720,N_4667);
xnor UO_567 (O_567,N_4036,N_4645);
nor UO_568 (O_568,N_4322,N_4638);
and UO_569 (O_569,N_4841,N_4541);
nand UO_570 (O_570,N_4003,N_4510);
nand UO_571 (O_571,N_4723,N_4020);
nand UO_572 (O_572,N_4748,N_4822);
and UO_573 (O_573,N_4691,N_4575);
xor UO_574 (O_574,N_4804,N_4102);
and UO_575 (O_575,N_4313,N_4444);
and UO_576 (O_576,N_4566,N_4119);
and UO_577 (O_577,N_4425,N_4727);
or UO_578 (O_578,N_4256,N_4395);
or UO_579 (O_579,N_4155,N_4350);
or UO_580 (O_580,N_4143,N_4850);
or UO_581 (O_581,N_4423,N_4024);
and UO_582 (O_582,N_4700,N_4915);
nor UO_583 (O_583,N_4603,N_4675);
and UO_584 (O_584,N_4347,N_4469);
or UO_585 (O_585,N_4428,N_4620);
nor UO_586 (O_586,N_4149,N_4632);
nand UO_587 (O_587,N_4632,N_4701);
or UO_588 (O_588,N_4632,N_4871);
and UO_589 (O_589,N_4532,N_4787);
and UO_590 (O_590,N_4708,N_4885);
and UO_591 (O_591,N_4652,N_4168);
nor UO_592 (O_592,N_4590,N_4598);
xnor UO_593 (O_593,N_4607,N_4093);
nand UO_594 (O_594,N_4638,N_4473);
or UO_595 (O_595,N_4489,N_4595);
or UO_596 (O_596,N_4183,N_4292);
or UO_597 (O_597,N_4976,N_4999);
nand UO_598 (O_598,N_4619,N_4932);
or UO_599 (O_599,N_4332,N_4482);
nor UO_600 (O_600,N_4309,N_4020);
nor UO_601 (O_601,N_4301,N_4590);
nand UO_602 (O_602,N_4885,N_4353);
and UO_603 (O_603,N_4386,N_4002);
and UO_604 (O_604,N_4842,N_4993);
and UO_605 (O_605,N_4275,N_4099);
or UO_606 (O_606,N_4082,N_4289);
nand UO_607 (O_607,N_4716,N_4881);
nor UO_608 (O_608,N_4657,N_4017);
or UO_609 (O_609,N_4191,N_4218);
or UO_610 (O_610,N_4550,N_4403);
nand UO_611 (O_611,N_4751,N_4163);
nor UO_612 (O_612,N_4873,N_4381);
xnor UO_613 (O_613,N_4774,N_4444);
or UO_614 (O_614,N_4561,N_4588);
and UO_615 (O_615,N_4149,N_4070);
and UO_616 (O_616,N_4358,N_4140);
or UO_617 (O_617,N_4469,N_4990);
or UO_618 (O_618,N_4091,N_4944);
nand UO_619 (O_619,N_4771,N_4797);
or UO_620 (O_620,N_4717,N_4037);
and UO_621 (O_621,N_4644,N_4121);
or UO_622 (O_622,N_4516,N_4925);
nor UO_623 (O_623,N_4100,N_4276);
and UO_624 (O_624,N_4345,N_4891);
and UO_625 (O_625,N_4362,N_4187);
or UO_626 (O_626,N_4585,N_4103);
or UO_627 (O_627,N_4495,N_4532);
or UO_628 (O_628,N_4545,N_4617);
or UO_629 (O_629,N_4663,N_4606);
and UO_630 (O_630,N_4296,N_4722);
nand UO_631 (O_631,N_4033,N_4533);
and UO_632 (O_632,N_4737,N_4474);
nor UO_633 (O_633,N_4037,N_4341);
or UO_634 (O_634,N_4614,N_4475);
or UO_635 (O_635,N_4071,N_4782);
and UO_636 (O_636,N_4478,N_4296);
nand UO_637 (O_637,N_4508,N_4626);
nor UO_638 (O_638,N_4119,N_4802);
or UO_639 (O_639,N_4719,N_4115);
nor UO_640 (O_640,N_4342,N_4045);
nand UO_641 (O_641,N_4114,N_4973);
nand UO_642 (O_642,N_4102,N_4741);
or UO_643 (O_643,N_4150,N_4132);
and UO_644 (O_644,N_4405,N_4924);
nand UO_645 (O_645,N_4377,N_4338);
nand UO_646 (O_646,N_4281,N_4816);
or UO_647 (O_647,N_4780,N_4521);
nand UO_648 (O_648,N_4368,N_4540);
or UO_649 (O_649,N_4920,N_4112);
nor UO_650 (O_650,N_4142,N_4937);
nor UO_651 (O_651,N_4500,N_4120);
and UO_652 (O_652,N_4019,N_4222);
and UO_653 (O_653,N_4441,N_4002);
or UO_654 (O_654,N_4591,N_4058);
nand UO_655 (O_655,N_4624,N_4431);
nand UO_656 (O_656,N_4801,N_4362);
nand UO_657 (O_657,N_4219,N_4567);
nor UO_658 (O_658,N_4342,N_4487);
nor UO_659 (O_659,N_4829,N_4608);
or UO_660 (O_660,N_4025,N_4001);
or UO_661 (O_661,N_4705,N_4005);
nand UO_662 (O_662,N_4242,N_4998);
nand UO_663 (O_663,N_4507,N_4859);
or UO_664 (O_664,N_4045,N_4621);
nor UO_665 (O_665,N_4257,N_4801);
nor UO_666 (O_666,N_4214,N_4949);
and UO_667 (O_667,N_4753,N_4981);
nand UO_668 (O_668,N_4260,N_4851);
and UO_669 (O_669,N_4514,N_4930);
nor UO_670 (O_670,N_4226,N_4802);
xor UO_671 (O_671,N_4878,N_4486);
or UO_672 (O_672,N_4453,N_4243);
nand UO_673 (O_673,N_4551,N_4785);
or UO_674 (O_674,N_4803,N_4462);
nor UO_675 (O_675,N_4229,N_4049);
nor UO_676 (O_676,N_4012,N_4977);
or UO_677 (O_677,N_4859,N_4891);
nand UO_678 (O_678,N_4706,N_4739);
and UO_679 (O_679,N_4295,N_4344);
or UO_680 (O_680,N_4274,N_4716);
and UO_681 (O_681,N_4135,N_4018);
or UO_682 (O_682,N_4660,N_4675);
nand UO_683 (O_683,N_4046,N_4147);
nor UO_684 (O_684,N_4783,N_4882);
nand UO_685 (O_685,N_4971,N_4901);
or UO_686 (O_686,N_4170,N_4482);
or UO_687 (O_687,N_4673,N_4424);
nand UO_688 (O_688,N_4637,N_4362);
and UO_689 (O_689,N_4148,N_4446);
or UO_690 (O_690,N_4513,N_4020);
and UO_691 (O_691,N_4386,N_4601);
or UO_692 (O_692,N_4014,N_4757);
nand UO_693 (O_693,N_4523,N_4403);
nor UO_694 (O_694,N_4187,N_4019);
or UO_695 (O_695,N_4540,N_4736);
nor UO_696 (O_696,N_4816,N_4335);
or UO_697 (O_697,N_4521,N_4808);
and UO_698 (O_698,N_4791,N_4573);
and UO_699 (O_699,N_4538,N_4870);
and UO_700 (O_700,N_4380,N_4610);
and UO_701 (O_701,N_4938,N_4983);
nand UO_702 (O_702,N_4393,N_4895);
or UO_703 (O_703,N_4348,N_4702);
and UO_704 (O_704,N_4277,N_4624);
and UO_705 (O_705,N_4228,N_4635);
nand UO_706 (O_706,N_4257,N_4000);
nor UO_707 (O_707,N_4148,N_4830);
or UO_708 (O_708,N_4266,N_4414);
nor UO_709 (O_709,N_4589,N_4180);
nand UO_710 (O_710,N_4512,N_4801);
nor UO_711 (O_711,N_4701,N_4666);
nand UO_712 (O_712,N_4266,N_4914);
and UO_713 (O_713,N_4411,N_4970);
and UO_714 (O_714,N_4765,N_4909);
or UO_715 (O_715,N_4876,N_4200);
nor UO_716 (O_716,N_4663,N_4935);
or UO_717 (O_717,N_4031,N_4785);
nor UO_718 (O_718,N_4576,N_4620);
and UO_719 (O_719,N_4861,N_4550);
nand UO_720 (O_720,N_4780,N_4681);
nor UO_721 (O_721,N_4369,N_4915);
nor UO_722 (O_722,N_4222,N_4321);
nor UO_723 (O_723,N_4880,N_4164);
and UO_724 (O_724,N_4165,N_4399);
or UO_725 (O_725,N_4742,N_4329);
or UO_726 (O_726,N_4107,N_4641);
or UO_727 (O_727,N_4767,N_4496);
and UO_728 (O_728,N_4971,N_4401);
nand UO_729 (O_729,N_4103,N_4108);
nand UO_730 (O_730,N_4387,N_4492);
or UO_731 (O_731,N_4959,N_4720);
or UO_732 (O_732,N_4554,N_4535);
nor UO_733 (O_733,N_4862,N_4809);
nor UO_734 (O_734,N_4297,N_4432);
or UO_735 (O_735,N_4263,N_4541);
nor UO_736 (O_736,N_4977,N_4669);
nor UO_737 (O_737,N_4219,N_4994);
nor UO_738 (O_738,N_4987,N_4171);
nor UO_739 (O_739,N_4703,N_4870);
or UO_740 (O_740,N_4514,N_4745);
or UO_741 (O_741,N_4284,N_4566);
nor UO_742 (O_742,N_4649,N_4094);
nor UO_743 (O_743,N_4372,N_4183);
and UO_744 (O_744,N_4440,N_4975);
or UO_745 (O_745,N_4358,N_4580);
nor UO_746 (O_746,N_4061,N_4192);
and UO_747 (O_747,N_4064,N_4388);
or UO_748 (O_748,N_4038,N_4063);
nor UO_749 (O_749,N_4079,N_4595);
or UO_750 (O_750,N_4430,N_4366);
nand UO_751 (O_751,N_4135,N_4780);
or UO_752 (O_752,N_4401,N_4429);
nor UO_753 (O_753,N_4340,N_4067);
nor UO_754 (O_754,N_4266,N_4757);
nor UO_755 (O_755,N_4459,N_4651);
nor UO_756 (O_756,N_4634,N_4141);
or UO_757 (O_757,N_4808,N_4863);
nor UO_758 (O_758,N_4843,N_4780);
and UO_759 (O_759,N_4855,N_4300);
or UO_760 (O_760,N_4735,N_4596);
or UO_761 (O_761,N_4042,N_4630);
or UO_762 (O_762,N_4937,N_4434);
nor UO_763 (O_763,N_4768,N_4479);
or UO_764 (O_764,N_4129,N_4360);
xnor UO_765 (O_765,N_4636,N_4962);
nand UO_766 (O_766,N_4894,N_4073);
or UO_767 (O_767,N_4309,N_4825);
nor UO_768 (O_768,N_4035,N_4577);
or UO_769 (O_769,N_4502,N_4701);
and UO_770 (O_770,N_4877,N_4924);
xnor UO_771 (O_771,N_4794,N_4640);
or UO_772 (O_772,N_4916,N_4706);
nand UO_773 (O_773,N_4444,N_4802);
nor UO_774 (O_774,N_4691,N_4098);
nor UO_775 (O_775,N_4749,N_4861);
nand UO_776 (O_776,N_4251,N_4298);
nand UO_777 (O_777,N_4686,N_4191);
and UO_778 (O_778,N_4019,N_4623);
and UO_779 (O_779,N_4183,N_4993);
nand UO_780 (O_780,N_4156,N_4002);
nand UO_781 (O_781,N_4707,N_4941);
nand UO_782 (O_782,N_4195,N_4192);
and UO_783 (O_783,N_4877,N_4249);
nor UO_784 (O_784,N_4591,N_4401);
and UO_785 (O_785,N_4896,N_4561);
nand UO_786 (O_786,N_4465,N_4985);
and UO_787 (O_787,N_4347,N_4965);
nor UO_788 (O_788,N_4920,N_4033);
or UO_789 (O_789,N_4654,N_4006);
and UO_790 (O_790,N_4510,N_4423);
or UO_791 (O_791,N_4882,N_4963);
or UO_792 (O_792,N_4823,N_4536);
or UO_793 (O_793,N_4923,N_4764);
or UO_794 (O_794,N_4052,N_4122);
or UO_795 (O_795,N_4780,N_4887);
and UO_796 (O_796,N_4770,N_4891);
nand UO_797 (O_797,N_4263,N_4043);
nand UO_798 (O_798,N_4720,N_4786);
nor UO_799 (O_799,N_4710,N_4967);
or UO_800 (O_800,N_4577,N_4150);
nor UO_801 (O_801,N_4890,N_4164);
xnor UO_802 (O_802,N_4809,N_4056);
and UO_803 (O_803,N_4495,N_4620);
nor UO_804 (O_804,N_4251,N_4147);
and UO_805 (O_805,N_4652,N_4182);
nor UO_806 (O_806,N_4819,N_4901);
nand UO_807 (O_807,N_4890,N_4641);
and UO_808 (O_808,N_4767,N_4295);
nor UO_809 (O_809,N_4044,N_4975);
nand UO_810 (O_810,N_4720,N_4371);
or UO_811 (O_811,N_4540,N_4481);
nand UO_812 (O_812,N_4611,N_4237);
and UO_813 (O_813,N_4849,N_4606);
and UO_814 (O_814,N_4212,N_4320);
and UO_815 (O_815,N_4189,N_4158);
or UO_816 (O_816,N_4785,N_4983);
and UO_817 (O_817,N_4922,N_4450);
nand UO_818 (O_818,N_4805,N_4474);
nor UO_819 (O_819,N_4851,N_4685);
nand UO_820 (O_820,N_4970,N_4543);
or UO_821 (O_821,N_4081,N_4289);
and UO_822 (O_822,N_4567,N_4712);
nand UO_823 (O_823,N_4664,N_4558);
or UO_824 (O_824,N_4740,N_4891);
nor UO_825 (O_825,N_4253,N_4262);
or UO_826 (O_826,N_4827,N_4631);
nor UO_827 (O_827,N_4278,N_4064);
nor UO_828 (O_828,N_4933,N_4534);
or UO_829 (O_829,N_4186,N_4973);
nand UO_830 (O_830,N_4425,N_4639);
and UO_831 (O_831,N_4970,N_4599);
nand UO_832 (O_832,N_4782,N_4606);
nor UO_833 (O_833,N_4494,N_4660);
nor UO_834 (O_834,N_4010,N_4527);
or UO_835 (O_835,N_4489,N_4037);
nand UO_836 (O_836,N_4697,N_4972);
and UO_837 (O_837,N_4632,N_4867);
and UO_838 (O_838,N_4131,N_4100);
nor UO_839 (O_839,N_4909,N_4052);
nand UO_840 (O_840,N_4204,N_4419);
nand UO_841 (O_841,N_4027,N_4444);
nand UO_842 (O_842,N_4561,N_4357);
nand UO_843 (O_843,N_4429,N_4122);
nand UO_844 (O_844,N_4125,N_4408);
nand UO_845 (O_845,N_4181,N_4991);
and UO_846 (O_846,N_4327,N_4984);
or UO_847 (O_847,N_4645,N_4272);
nor UO_848 (O_848,N_4534,N_4425);
or UO_849 (O_849,N_4690,N_4598);
and UO_850 (O_850,N_4058,N_4872);
nand UO_851 (O_851,N_4980,N_4534);
and UO_852 (O_852,N_4520,N_4141);
or UO_853 (O_853,N_4582,N_4660);
or UO_854 (O_854,N_4828,N_4929);
or UO_855 (O_855,N_4789,N_4845);
nand UO_856 (O_856,N_4989,N_4653);
nand UO_857 (O_857,N_4078,N_4349);
nor UO_858 (O_858,N_4558,N_4144);
nand UO_859 (O_859,N_4651,N_4061);
and UO_860 (O_860,N_4883,N_4945);
nand UO_861 (O_861,N_4710,N_4046);
or UO_862 (O_862,N_4910,N_4961);
and UO_863 (O_863,N_4919,N_4816);
and UO_864 (O_864,N_4813,N_4704);
or UO_865 (O_865,N_4377,N_4335);
or UO_866 (O_866,N_4492,N_4059);
nor UO_867 (O_867,N_4874,N_4576);
nand UO_868 (O_868,N_4256,N_4837);
nor UO_869 (O_869,N_4885,N_4502);
and UO_870 (O_870,N_4786,N_4430);
nor UO_871 (O_871,N_4499,N_4758);
nand UO_872 (O_872,N_4269,N_4030);
nand UO_873 (O_873,N_4386,N_4496);
nand UO_874 (O_874,N_4898,N_4878);
nand UO_875 (O_875,N_4134,N_4376);
or UO_876 (O_876,N_4980,N_4102);
nand UO_877 (O_877,N_4586,N_4335);
and UO_878 (O_878,N_4187,N_4870);
nor UO_879 (O_879,N_4018,N_4108);
xnor UO_880 (O_880,N_4057,N_4363);
nor UO_881 (O_881,N_4783,N_4128);
or UO_882 (O_882,N_4938,N_4766);
nand UO_883 (O_883,N_4536,N_4112);
or UO_884 (O_884,N_4402,N_4308);
nand UO_885 (O_885,N_4109,N_4043);
and UO_886 (O_886,N_4465,N_4940);
or UO_887 (O_887,N_4698,N_4939);
or UO_888 (O_888,N_4246,N_4256);
or UO_889 (O_889,N_4389,N_4921);
and UO_890 (O_890,N_4631,N_4453);
or UO_891 (O_891,N_4527,N_4327);
and UO_892 (O_892,N_4978,N_4700);
nand UO_893 (O_893,N_4997,N_4275);
or UO_894 (O_894,N_4663,N_4328);
nor UO_895 (O_895,N_4510,N_4263);
and UO_896 (O_896,N_4052,N_4278);
or UO_897 (O_897,N_4210,N_4676);
nor UO_898 (O_898,N_4250,N_4120);
nand UO_899 (O_899,N_4264,N_4466);
and UO_900 (O_900,N_4354,N_4408);
nand UO_901 (O_901,N_4309,N_4074);
and UO_902 (O_902,N_4713,N_4061);
nor UO_903 (O_903,N_4920,N_4598);
and UO_904 (O_904,N_4198,N_4464);
nor UO_905 (O_905,N_4308,N_4628);
nand UO_906 (O_906,N_4235,N_4169);
nand UO_907 (O_907,N_4455,N_4781);
or UO_908 (O_908,N_4945,N_4299);
nor UO_909 (O_909,N_4856,N_4690);
and UO_910 (O_910,N_4295,N_4345);
nor UO_911 (O_911,N_4109,N_4463);
or UO_912 (O_912,N_4017,N_4957);
nor UO_913 (O_913,N_4901,N_4271);
nand UO_914 (O_914,N_4568,N_4109);
or UO_915 (O_915,N_4887,N_4640);
nand UO_916 (O_916,N_4901,N_4609);
nor UO_917 (O_917,N_4005,N_4220);
and UO_918 (O_918,N_4092,N_4519);
or UO_919 (O_919,N_4077,N_4430);
and UO_920 (O_920,N_4222,N_4562);
and UO_921 (O_921,N_4468,N_4437);
and UO_922 (O_922,N_4685,N_4024);
nor UO_923 (O_923,N_4346,N_4057);
nand UO_924 (O_924,N_4895,N_4594);
nor UO_925 (O_925,N_4680,N_4975);
and UO_926 (O_926,N_4849,N_4144);
nand UO_927 (O_927,N_4883,N_4644);
nor UO_928 (O_928,N_4657,N_4432);
xnor UO_929 (O_929,N_4573,N_4551);
nor UO_930 (O_930,N_4821,N_4786);
or UO_931 (O_931,N_4863,N_4588);
nor UO_932 (O_932,N_4076,N_4671);
and UO_933 (O_933,N_4330,N_4907);
nand UO_934 (O_934,N_4474,N_4753);
or UO_935 (O_935,N_4010,N_4496);
nor UO_936 (O_936,N_4612,N_4942);
or UO_937 (O_937,N_4007,N_4662);
and UO_938 (O_938,N_4636,N_4579);
xor UO_939 (O_939,N_4265,N_4770);
nand UO_940 (O_940,N_4735,N_4563);
nor UO_941 (O_941,N_4365,N_4545);
or UO_942 (O_942,N_4645,N_4552);
nand UO_943 (O_943,N_4624,N_4653);
and UO_944 (O_944,N_4300,N_4198);
or UO_945 (O_945,N_4889,N_4636);
nor UO_946 (O_946,N_4169,N_4916);
and UO_947 (O_947,N_4602,N_4717);
and UO_948 (O_948,N_4617,N_4079);
or UO_949 (O_949,N_4309,N_4808);
or UO_950 (O_950,N_4673,N_4572);
or UO_951 (O_951,N_4260,N_4426);
nand UO_952 (O_952,N_4044,N_4481);
or UO_953 (O_953,N_4584,N_4126);
nand UO_954 (O_954,N_4536,N_4491);
and UO_955 (O_955,N_4549,N_4939);
or UO_956 (O_956,N_4153,N_4532);
nand UO_957 (O_957,N_4844,N_4801);
or UO_958 (O_958,N_4779,N_4590);
nor UO_959 (O_959,N_4779,N_4899);
nand UO_960 (O_960,N_4553,N_4954);
nand UO_961 (O_961,N_4955,N_4129);
and UO_962 (O_962,N_4660,N_4769);
nand UO_963 (O_963,N_4818,N_4666);
or UO_964 (O_964,N_4267,N_4268);
and UO_965 (O_965,N_4381,N_4722);
and UO_966 (O_966,N_4228,N_4292);
or UO_967 (O_967,N_4930,N_4815);
and UO_968 (O_968,N_4520,N_4383);
nand UO_969 (O_969,N_4048,N_4628);
and UO_970 (O_970,N_4820,N_4670);
nand UO_971 (O_971,N_4080,N_4431);
and UO_972 (O_972,N_4980,N_4218);
or UO_973 (O_973,N_4869,N_4877);
nor UO_974 (O_974,N_4327,N_4499);
nand UO_975 (O_975,N_4229,N_4667);
or UO_976 (O_976,N_4656,N_4337);
nand UO_977 (O_977,N_4360,N_4676);
nand UO_978 (O_978,N_4721,N_4157);
nor UO_979 (O_979,N_4128,N_4625);
and UO_980 (O_980,N_4643,N_4927);
or UO_981 (O_981,N_4732,N_4065);
and UO_982 (O_982,N_4135,N_4128);
or UO_983 (O_983,N_4706,N_4789);
nor UO_984 (O_984,N_4488,N_4124);
nand UO_985 (O_985,N_4571,N_4700);
and UO_986 (O_986,N_4747,N_4078);
nand UO_987 (O_987,N_4816,N_4794);
nand UO_988 (O_988,N_4720,N_4896);
or UO_989 (O_989,N_4829,N_4672);
nand UO_990 (O_990,N_4499,N_4130);
nor UO_991 (O_991,N_4247,N_4788);
nor UO_992 (O_992,N_4048,N_4335);
nor UO_993 (O_993,N_4025,N_4826);
nor UO_994 (O_994,N_4816,N_4608);
and UO_995 (O_995,N_4873,N_4605);
and UO_996 (O_996,N_4851,N_4061);
or UO_997 (O_997,N_4237,N_4803);
nor UO_998 (O_998,N_4627,N_4852);
or UO_999 (O_999,N_4598,N_4719);
endmodule