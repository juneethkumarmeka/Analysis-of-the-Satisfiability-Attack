module basic_1000_10000_1500_4_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nor U0 (N_0,In_816,In_362);
nand U1 (N_1,In_46,In_41);
nor U2 (N_2,In_294,In_292);
or U3 (N_3,In_879,In_479);
nand U4 (N_4,In_425,In_762);
nand U5 (N_5,In_528,In_549);
nand U6 (N_6,In_763,In_713);
nor U7 (N_7,In_443,In_183);
xnor U8 (N_8,In_393,In_585);
nor U9 (N_9,In_53,In_306);
or U10 (N_10,In_553,In_165);
and U11 (N_11,In_188,In_583);
nor U12 (N_12,In_821,In_21);
nand U13 (N_13,In_92,In_18);
nor U14 (N_14,In_96,In_375);
or U15 (N_15,In_197,In_285);
nand U16 (N_16,In_400,In_575);
nand U17 (N_17,In_789,In_345);
and U18 (N_18,In_771,In_941);
nor U19 (N_19,In_129,In_220);
nand U20 (N_20,In_350,In_904);
and U21 (N_21,In_358,In_113);
or U22 (N_22,In_132,In_245);
or U23 (N_23,In_711,In_335);
or U24 (N_24,In_330,In_311);
or U25 (N_25,In_300,In_656);
or U26 (N_26,In_986,In_647);
or U27 (N_27,In_557,In_288);
and U28 (N_28,In_80,In_338);
or U29 (N_29,In_938,In_686);
and U30 (N_30,In_935,In_864);
and U31 (N_31,In_396,In_861);
or U32 (N_32,In_468,In_377);
nor U33 (N_33,In_937,In_360);
or U34 (N_34,In_95,In_546);
nand U35 (N_35,In_392,In_431);
or U36 (N_36,In_442,In_20);
nor U37 (N_37,In_613,In_106);
nor U38 (N_38,In_796,In_397);
or U39 (N_39,In_695,In_888);
or U40 (N_40,In_54,In_232);
nor U41 (N_41,In_819,In_156);
nor U42 (N_42,In_641,In_445);
and U43 (N_43,In_812,In_174);
and U44 (N_44,In_40,In_138);
nand U45 (N_45,In_411,In_94);
nand U46 (N_46,In_595,In_952);
nor U47 (N_47,In_227,In_144);
and U48 (N_48,In_880,In_122);
nand U49 (N_49,In_191,In_620);
and U50 (N_50,In_126,In_459);
nand U51 (N_51,In_295,In_597);
nand U52 (N_52,In_190,In_718);
and U53 (N_53,In_507,In_200);
nand U54 (N_54,In_694,In_483);
and U55 (N_55,In_680,In_676);
xnor U56 (N_56,In_302,In_591);
or U57 (N_57,In_82,In_916);
nand U58 (N_58,In_139,In_145);
nand U59 (N_59,In_761,In_867);
nor U60 (N_60,In_811,In_262);
and U61 (N_61,In_517,In_240);
or U62 (N_62,In_348,In_572);
or U63 (N_63,In_540,In_838);
or U64 (N_64,In_7,In_353);
nor U65 (N_65,In_65,In_673);
nor U66 (N_66,In_351,In_389);
or U67 (N_67,In_604,In_498);
and U68 (N_68,In_461,In_851);
nor U69 (N_69,In_989,In_570);
nor U70 (N_70,In_973,In_870);
nor U71 (N_71,In_757,In_238);
nand U72 (N_72,In_746,In_751);
nor U73 (N_73,In_102,In_782);
or U74 (N_74,In_529,In_2);
or U75 (N_75,In_203,In_605);
nor U76 (N_76,In_76,In_963);
and U77 (N_77,In_667,In_648);
or U78 (N_78,In_634,In_551);
nor U79 (N_79,In_753,In_772);
nor U80 (N_80,In_632,In_171);
nor U81 (N_81,In_176,In_31);
nor U82 (N_82,In_592,In_697);
nor U83 (N_83,In_428,In_886);
nand U84 (N_84,In_602,In_317);
and U85 (N_85,In_755,In_419);
nor U86 (N_86,In_421,In_845);
and U87 (N_87,In_246,In_170);
and U88 (N_88,In_775,In_258);
nor U89 (N_89,In_930,In_93);
or U90 (N_90,In_434,In_924);
nor U91 (N_91,In_534,In_730);
and U92 (N_92,In_312,In_29);
or U93 (N_93,In_465,In_496);
nand U94 (N_94,In_919,In_902);
nand U95 (N_95,In_674,In_788);
nand U96 (N_96,In_162,In_361);
and U97 (N_97,In_38,In_325);
nor U98 (N_98,In_614,In_889);
and U99 (N_99,In_289,In_341);
nor U100 (N_100,In_731,In_12);
and U101 (N_101,In_467,In_412);
nand U102 (N_102,In_582,In_298);
and U103 (N_103,In_765,In_961);
nand U104 (N_104,In_424,In_505);
or U105 (N_105,In_542,In_630);
nor U106 (N_106,In_268,In_290);
nor U107 (N_107,In_482,In_305);
or U108 (N_108,In_901,In_573);
and U109 (N_109,In_148,In_208);
or U110 (N_110,In_115,In_172);
and U111 (N_111,In_150,In_355);
or U112 (N_112,In_652,In_635);
nand U113 (N_113,In_970,In_808);
nand U114 (N_114,In_503,In_803);
or U115 (N_115,In_568,In_844);
or U116 (N_116,In_678,In_975);
or U117 (N_117,In_908,In_315);
and U118 (N_118,In_35,In_742);
or U119 (N_119,In_233,In_881);
nand U120 (N_120,In_756,In_26);
or U121 (N_121,In_4,In_267);
or U122 (N_122,In_147,In_622);
or U123 (N_123,In_22,In_616);
and U124 (N_124,In_259,In_644);
nor U125 (N_125,In_559,In_600);
nand U126 (N_126,In_100,In_328);
or U127 (N_127,In_842,In_199);
nor U128 (N_128,In_956,In_669);
nand U129 (N_129,In_764,In_88);
nor U130 (N_130,In_194,In_60);
and U131 (N_131,In_463,In_284);
and U132 (N_132,In_776,In_719);
nand U133 (N_133,In_447,In_184);
nor U134 (N_134,In_318,In_903);
and U135 (N_135,In_965,In_633);
nand U136 (N_136,In_795,In_688);
and U137 (N_137,In_860,In_181);
or U138 (N_138,In_670,In_706);
and U139 (N_139,In_319,In_168);
nand U140 (N_140,In_728,In_455);
or U141 (N_141,In_805,In_394);
and U142 (N_142,In_417,In_687);
or U143 (N_143,In_502,In_642);
nor U144 (N_144,In_804,In_407);
nor U145 (N_145,In_940,In_110);
and U146 (N_146,In_433,In_942);
or U147 (N_147,In_485,In_690);
nand U148 (N_148,In_67,In_13);
or U149 (N_149,In_552,In_809);
xor U150 (N_150,In_979,In_160);
or U151 (N_151,In_276,In_875);
nand U152 (N_152,In_254,In_63);
nand U153 (N_153,In_367,In_155);
nand U154 (N_154,In_863,In_987);
or U155 (N_155,In_539,In_173);
nand U156 (N_156,In_725,In_905);
and U157 (N_157,In_235,In_950);
and U158 (N_158,In_66,In_855);
and U159 (N_159,In_726,In_493);
or U160 (N_160,In_117,In_663);
and U161 (N_161,In_167,In_737);
nand U162 (N_162,In_609,In_536);
nand U163 (N_163,In_273,In_717);
nor U164 (N_164,In_133,In_899);
xor U165 (N_165,In_215,In_266);
or U166 (N_166,In_177,In_786);
or U167 (N_167,In_696,In_42);
or U168 (N_168,In_187,In_621);
nor U169 (N_169,In_229,In_379);
nor U170 (N_170,In_499,In_453);
nand U171 (N_171,In_449,In_236);
nor U172 (N_172,In_698,In_943);
and U173 (N_173,In_286,In_234);
and U174 (N_174,In_998,In_885);
or U175 (N_175,In_506,In_857);
and U176 (N_176,In_140,In_967);
and U177 (N_177,In_391,In_612);
nand U178 (N_178,In_323,In_107);
and U179 (N_179,In_274,In_858);
nand U180 (N_180,In_301,In_303);
or U181 (N_181,In_475,In_256);
nor U182 (N_182,In_541,In_149);
nand U183 (N_183,In_270,In_959);
nand U184 (N_184,In_251,In_560);
and U185 (N_185,In_5,In_606);
nand U186 (N_186,In_783,In_747);
or U187 (N_187,In_985,In_263);
nor U188 (N_188,In_374,In_118);
nor U189 (N_189,In_221,In_334);
and U190 (N_190,In_11,In_287);
or U191 (N_191,In_624,In_797);
and U192 (N_192,In_932,In_225);
nor U193 (N_193,In_313,In_955);
or U194 (N_194,In_340,In_33);
nand U195 (N_195,In_324,In_957);
nand U196 (N_196,In_689,In_915);
nand U197 (N_197,In_531,In_121);
or U198 (N_198,In_481,In_662);
nor U199 (N_199,In_429,In_617);
and U200 (N_200,In_964,In_52);
or U201 (N_201,In_997,In_241);
or U202 (N_202,In_824,In_734);
nand U203 (N_203,In_370,In_566);
nor U204 (N_204,In_159,In_427);
and U205 (N_205,In_623,In_55);
nand U206 (N_206,In_395,In_137);
and U207 (N_207,In_972,In_32);
and U208 (N_208,In_206,In_525);
or U209 (N_209,In_849,In_834);
nand U210 (N_210,In_169,In_210);
nor U211 (N_211,In_712,In_527);
or U212 (N_212,In_587,In_835);
nor U213 (N_213,In_703,In_408);
nor U214 (N_214,In_212,In_253);
and U215 (N_215,In_887,In_28);
and U216 (N_216,In_39,In_247);
or U217 (N_217,In_671,In_15);
nor U218 (N_218,In_666,In_822);
or U219 (N_219,In_339,In_913);
nand U220 (N_220,In_320,In_770);
nor U221 (N_221,In_495,In_982);
and U222 (N_222,In_474,In_296);
and U223 (N_223,In_404,In_640);
or U224 (N_224,In_872,In_814);
nand U225 (N_225,In_920,In_205);
or U226 (N_226,In_836,In_509);
nor U227 (N_227,In_874,In_104);
and U228 (N_228,In_741,In_840);
nand U229 (N_229,In_657,In_626);
or U230 (N_230,In_265,In_114);
and U231 (N_231,In_564,In_580);
nor U232 (N_232,In_843,In_371);
nand U233 (N_233,In_37,In_629);
and U234 (N_234,In_709,In_142);
nand U235 (N_235,In_643,In_84);
xor U236 (N_236,In_494,In_388);
nor U237 (N_237,In_349,In_346);
nand U238 (N_238,In_399,In_900);
nor U239 (N_239,In_24,In_157);
nand U240 (N_240,In_794,In_213);
nor U241 (N_241,In_17,In_243);
nand U242 (N_242,In_226,In_448);
or U243 (N_243,In_639,In_6);
nor U244 (N_244,In_248,In_991);
or U245 (N_245,In_675,In_175);
and U246 (N_246,In_710,In_721);
and U247 (N_247,In_739,In_596);
nand U248 (N_248,In_146,In_951);
nor U249 (N_249,In_769,In_23);
or U250 (N_250,In_555,In_239);
nand U251 (N_251,In_131,In_768);
nand U252 (N_252,In_856,In_774);
nand U253 (N_253,In_598,In_34);
and U254 (N_254,In_577,In_58);
or U255 (N_255,In_70,In_309);
or U256 (N_256,In_519,In_672);
or U257 (N_257,In_754,In_890);
nand U258 (N_258,In_354,In_544);
and U259 (N_259,In_108,In_430);
and U260 (N_260,In_610,In_865);
or U261 (N_261,In_790,In_185);
nor U262 (N_262,In_594,In_550);
and U263 (N_263,In_378,In_948);
or U264 (N_264,In_261,In_299);
nand U265 (N_265,In_112,In_871);
nor U266 (N_266,In_841,In_599);
nor U267 (N_267,In_877,In_569);
nor U268 (N_268,In_882,In_61);
xor U269 (N_269,In_833,In_196);
nor U270 (N_270,In_272,In_120);
nand U271 (N_271,In_222,In_242);
and U272 (N_272,In_14,In_79);
nor U273 (N_273,In_522,In_193);
nand U274 (N_274,In_44,In_255);
and U275 (N_275,In_618,In_538);
nand U276 (N_276,In_356,In_615);
and U277 (N_277,In_883,In_446);
or U278 (N_278,In_578,In_105);
and U279 (N_279,In_166,In_501);
and U280 (N_280,In_87,In_535);
and U281 (N_281,In_476,In_75);
and U282 (N_282,In_418,In_907);
nor U283 (N_283,In_99,In_336);
nor U284 (N_284,In_401,In_83);
nand U285 (N_285,In_700,In_343);
nor U286 (N_286,In_178,In_347);
nor U287 (N_287,In_97,In_231);
and U288 (N_288,In_625,In_477);
and U289 (N_289,In_500,In_368);
nand U290 (N_290,In_876,In_659);
or U291 (N_291,In_969,In_278);
nor U292 (N_292,In_911,In_798);
nor U293 (N_293,In_369,In_484);
xor U294 (N_294,In_530,In_124);
nor U295 (N_295,In_590,In_151);
nand U296 (N_296,In_854,In_909);
and U297 (N_297,In_154,In_866);
or U298 (N_298,In_116,In_123);
or U299 (N_299,In_413,In_217);
or U300 (N_300,In_999,In_827);
nand U301 (N_301,In_420,In_664);
nand U302 (N_302,In_735,In_16);
and U303 (N_303,In_894,In_727);
or U304 (N_304,In_91,In_898);
and U305 (N_305,In_912,In_636);
nand U306 (N_306,In_548,In_415);
and U307 (N_307,In_103,In_0);
nand U308 (N_308,In_588,In_800);
and U309 (N_309,In_581,In_884);
nor U310 (N_310,In_163,In_611);
nand U311 (N_311,In_8,In_750);
or U312 (N_312,In_745,In_683);
or U313 (N_313,In_631,In_489);
or U314 (N_314,In_817,In_71);
nor U315 (N_315,In_852,In_56);
nand U316 (N_316,In_649,In_677);
xnor U317 (N_317,In_944,In_398);
nand U318 (N_318,In_279,In_486);
or U319 (N_319,In_219,In_781);
nor U320 (N_320,In_971,In_974);
nand U321 (N_321,In_988,In_204);
nand U322 (N_322,In_910,In_466);
and U323 (N_323,In_593,In_409);
nand U324 (N_324,In_724,In_416);
nand U325 (N_325,In_653,In_962);
and U326 (N_326,In_682,In_561);
and U327 (N_327,In_304,In_947);
nor U328 (N_328,In_510,In_651);
and U329 (N_329,In_977,In_976);
and U330 (N_330,In_638,In_422);
nand U331 (N_331,In_440,In_490);
xor U332 (N_332,In_778,In_224);
nand U333 (N_333,In_939,In_934);
and U334 (N_334,In_143,In_508);
or U335 (N_335,In_321,In_584);
and U336 (N_336,In_722,In_471);
or U337 (N_337,In_359,In_277);
or U338 (N_338,In_458,In_460);
nor U339 (N_339,In_738,In_1);
nand U340 (N_340,In_869,In_926);
or U341 (N_341,In_562,In_996);
nor U342 (N_342,In_314,In_310);
nor U343 (N_343,In_381,In_946);
nand U344 (N_344,In_567,In_787);
or U345 (N_345,In_576,In_980);
or U346 (N_346,In_19,In_152);
or U347 (N_347,In_101,In_511);
or U348 (N_348,In_981,In_237);
nand U349 (N_349,In_504,In_917);
nand U350 (N_350,In_281,In_820);
nand U351 (N_351,In_376,In_766);
or U352 (N_352,In_715,In_563);
and U353 (N_353,In_111,In_815);
nand U354 (N_354,In_383,In_352);
nor U355 (N_355,In_784,In_818);
or U356 (N_356,In_136,In_269);
and U357 (N_357,In_720,In_36);
nand U358 (N_358,In_936,In_921);
or U359 (N_359,In_89,In_480);
nand U360 (N_360,In_810,In_405);
xnor U361 (N_361,In_556,In_896);
nand U362 (N_362,In_382,In_373);
nand U363 (N_363,In_760,In_627);
nand U364 (N_364,In_785,In_520);
or U365 (N_365,In_994,In_729);
and U366 (N_366,In_848,In_223);
nor U367 (N_367,In_966,In_73);
nor U368 (N_368,In_515,In_859);
or U369 (N_369,In_329,In_823);
or U370 (N_370,In_492,In_707);
nand U371 (N_371,In_589,In_316);
or U372 (N_372,In_749,In_64);
and U373 (N_373,In_62,In_574);
and U374 (N_374,In_68,In_57);
or U375 (N_375,In_554,In_161);
nor U376 (N_376,In_608,In_47);
nand U377 (N_377,In_752,In_692);
nand U378 (N_378,In_839,In_792);
nand U379 (N_379,In_780,In_513);
nor U380 (N_380,In_125,In_332);
nor U381 (N_381,In_410,In_828);
nand U382 (N_382,In_462,In_189);
nand U383 (N_383,In_77,In_601);
and U384 (N_384,In_327,In_958);
or U385 (N_385,In_406,In_195);
and U386 (N_386,In_514,In_532);
and U387 (N_387,In_214,In_968);
nand U388 (N_388,In_873,In_260);
or U389 (N_389,In_211,In_846);
or U390 (N_390,In_586,In_660);
and U391 (N_391,In_565,In_579);
or U392 (N_392,In_78,In_9);
and U393 (N_393,In_773,In_469);
xor U394 (N_394,In_699,In_470);
nand U395 (N_395,In_128,In_439);
nor U396 (N_396,In_931,In_69);
nand U397 (N_397,In_923,In_230);
nor U398 (N_398,In_668,In_135);
nor U399 (N_399,In_436,In_645);
nor U400 (N_400,In_925,In_333);
nand U401 (N_401,In_252,In_830);
nand U402 (N_402,In_198,In_127);
nand U403 (N_403,In_293,In_244);
nor U404 (N_404,In_228,In_403);
nor U405 (N_405,In_435,In_723);
and U406 (N_406,In_134,In_654);
nor U407 (N_407,In_813,In_646);
or U408 (N_408,In_922,In_344);
nand U409 (N_409,In_49,In_806);
and U410 (N_410,In_895,In_130);
or U411 (N_411,In_868,In_691);
nand U412 (N_412,In_478,In_650);
and U413 (N_413,In_322,In_831);
nand U414 (N_414,In_3,In_337);
nand U415 (N_415,In_291,In_74);
xnor U416 (N_416,In_779,In_109);
nand U417 (N_417,In_825,In_450);
or U418 (N_418,In_521,In_43);
or U419 (N_419,In_826,In_533);
nand U420 (N_420,In_464,In_364);
nand U421 (N_421,In_209,In_10);
nor U422 (N_422,In_523,In_441);
nand U423 (N_423,In_207,In_202);
nor U424 (N_424,In_153,In_990);
nand U425 (N_425,In_98,In_283);
nor U426 (N_426,In_363,In_81);
or U427 (N_427,In_897,In_603);
nor U428 (N_428,In_704,In_59);
nand U429 (N_429,In_384,In_331);
nor U430 (N_430,In_452,In_685);
and U431 (N_431,In_491,In_141);
nor U432 (N_432,In_380,In_182);
and U433 (N_433,In_216,In_414);
nor U434 (N_434,In_893,In_949);
and U435 (N_435,In_250,In_847);
and U436 (N_436,In_862,In_85);
nor U437 (N_437,In_432,In_801);
or U438 (N_438,In_472,In_402);
nor U439 (N_439,In_953,In_702);
nand U440 (N_440,In_516,In_748);
nor U441 (N_441,In_264,In_619);
nand U442 (N_442,In_426,In_802);
and U443 (N_443,In_733,In_928);
nor U444 (N_444,In_119,In_164);
nand U445 (N_445,In_637,In_984);
or U446 (N_446,In_777,In_473);
nand U447 (N_447,In_48,In_497);
or U448 (N_448,In_558,In_454);
or U449 (N_449,In_27,In_456);
xor U450 (N_450,In_488,In_978);
nand U451 (N_451,In_832,In_387);
nand U452 (N_452,In_807,In_767);
nor U453 (N_453,In_192,In_249);
and U454 (N_454,In_326,In_906);
nand U455 (N_455,In_282,In_693);
and U456 (N_456,In_201,In_993);
or U457 (N_457,In_51,In_385);
nor U458 (N_458,In_72,In_714);
nor U459 (N_459,In_512,In_524);
nor U460 (N_460,In_954,In_927);
or U461 (N_461,In_661,In_892);
or U462 (N_462,In_50,In_372);
and U463 (N_463,In_366,In_179);
and U464 (N_464,In_918,In_758);
or U465 (N_465,In_357,In_992);
nand U466 (N_466,In_90,In_732);
and U467 (N_467,In_850,In_297);
xor U468 (N_468,In_829,In_543);
nor U469 (N_469,In_186,In_853);
or U470 (N_470,In_744,In_607);
nor U471 (N_471,In_679,In_655);
and U472 (N_472,In_218,In_736);
and U473 (N_473,In_280,In_390);
and U474 (N_474,In_571,In_342);
or U475 (N_475,In_945,In_929);
nand U476 (N_476,In_708,In_995);
or U477 (N_477,In_30,In_878);
nor U478 (N_478,In_933,In_518);
nand U479 (N_479,In_437,In_716);
xor U480 (N_480,In_628,In_545);
nor U481 (N_481,In_271,In_793);
nor U482 (N_482,In_537,In_307);
nor U483 (N_483,In_960,In_444);
or U484 (N_484,In_451,In_45);
xnor U485 (N_485,In_158,In_438);
nand U486 (N_486,In_86,In_891);
and U487 (N_487,In_526,In_423);
nor U488 (N_488,In_308,In_681);
and U489 (N_489,In_791,In_386);
nor U490 (N_490,In_658,In_983);
and U491 (N_491,In_547,In_914);
nand U492 (N_492,In_743,In_701);
and U493 (N_493,In_257,In_684);
nand U494 (N_494,In_275,In_705);
or U495 (N_495,In_799,In_487);
or U496 (N_496,In_365,In_759);
nand U497 (N_497,In_180,In_665);
nor U498 (N_498,In_740,In_25);
and U499 (N_499,In_837,In_457);
nand U500 (N_500,In_492,In_111);
nor U501 (N_501,In_278,In_233);
nand U502 (N_502,In_75,In_94);
or U503 (N_503,In_812,In_618);
nor U504 (N_504,In_631,In_140);
nor U505 (N_505,In_250,In_497);
nor U506 (N_506,In_981,In_962);
and U507 (N_507,In_678,In_827);
and U508 (N_508,In_996,In_420);
or U509 (N_509,In_868,In_54);
nor U510 (N_510,In_725,In_599);
or U511 (N_511,In_285,In_395);
nor U512 (N_512,In_558,In_368);
or U513 (N_513,In_462,In_855);
nand U514 (N_514,In_56,In_543);
nor U515 (N_515,In_314,In_692);
nand U516 (N_516,In_71,In_99);
and U517 (N_517,In_739,In_815);
nand U518 (N_518,In_589,In_122);
nand U519 (N_519,In_741,In_419);
nand U520 (N_520,In_169,In_845);
nand U521 (N_521,In_54,In_221);
nand U522 (N_522,In_262,In_768);
nand U523 (N_523,In_13,In_887);
nor U524 (N_524,In_987,In_160);
xnor U525 (N_525,In_678,In_123);
and U526 (N_526,In_289,In_462);
and U527 (N_527,In_383,In_388);
nand U528 (N_528,In_480,In_419);
nand U529 (N_529,In_51,In_228);
or U530 (N_530,In_490,In_608);
and U531 (N_531,In_453,In_379);
nor U532 (N_532,In_648,In_780);
xnor U533 (N_533,In_941,In_570);
or U534 (N_534,In_716,In_873);
nand U535 (N_535,In_865,In_695);
nand U536 (N_536,In_599,In_30);
or U537 (N_537,In_433,In_558);
nand U538 (N_538,In_704,In_755);
nand U539 (N_539,In_800,In_675);
or U540 (N_540,In_592,In_777);
nand U541 (N_541,In_442,In_969);
or U542 (N_542,In_686,In_512);
or U543 (N_543,In_445,In_140);
nor U544 (N_544,In_14,In_656);
and U545 (N_545,In_740,In_743);
nor U546 (N_546,In_795,In_709);
or U547 (N_547,In_336,In_449);
or U548 (N_548,In_451,In_686);
nand U549 (N_549,In_478,In_601);
or U550 (N_550,In_183,In_680);
or U551 (N_551,In_557,In_418);
or U552 (N_552,In_18,In_420);
nor U553 (N_553,In_286,In_827);
nor U554 (N_554,In_379,In_602);
and U555 (N_555,In_185,In_727);
or U556 (N_556,In_57,In_104);
or U557 (N_557,In_112,In_474);
and U558 (N_558,In_884,In_61);
or U559 (N_559,In_212,In_273);
and U560 (N_560,In_397,In_491);
or U561 (N_561,In_922,In_924);
nand U562 (N_562,In_578,In_690);
and U563 (N_563,In_242,In_990);
and U564 (N_564,In_768,In_484);
or U565 (N_565,In_894,In_381);
nand U566 (N_566,In_90,In_867);
nand U567 (N_567,In_19,In_735);
or U568 (N_568,In_587,In_701);
and U569 (N_569,In_930,In_397);
or U570 (N_570,In_246,In_134);
nand U571 (N_571,In_466,In_403);
nand U572 (N_572,In_968,In_836);
or U573 (N_573,In_692,In_185);
nor U574 (N_574,In_643,In_928);
nor U575 (N_575,In_609,In_358);
or U576 (N_576,In_632,In_307);
and U577 (N_577,In_799,In_834);
and U578 (N_578,In_994,In_378);
or U579 (N_579,In_955,In_929);
xor U580 (N_580,In_782,In_118);
nand U581 (N_581,In_974,In_213);
and U582 (N_582,In_93,In_807);
or U583 (N_583,In_613,In_159);
or U584 (N_584,In_104,In_924);
or U585 (N_585,In_439,In_123);
nor U586 (N_586,In_529,In_742);
nor U587 (N_587,In_176,In_800);
nor U588 (N_588,In_512,In_971);
nand U589 (N_589,In_953,In_839);
or U590 (N_590,In_338,In_952);
nor U591 (N_591,In_268,In_942);
nor U592 (N_592,In_836,In_60);
nand U593 (N_593,In_943,In_208);
nor U594 (N_594,In_215,In_906);
xnor U595 (N_595,In_261,In_650);
and U596 (N_596,In_951,In_401);
or U597 (N_597,In_524,In_43);
and U598 (N_598,In_808,In_709);
nand U599 (N_599,In_474,In_567);
nor U600 (N_600,In_429,In_272);
and U601 (N_601,In_779,In_728);
or U602 (N_602,In_495,In_805);
and U603 (N_603,In_257,In_844);
nor U604 (N_604,In_113,In_357);
and U605 (N_605,In_441,In_835);
nor U606 (N_606,In_361,In_549);
and U607 (N_607,In_981,In_145);
xor U608 (N_608,In_467,In_61);
or U609 (N_609,In_806,In_341);
nand U610 (N_610,In_1,In_470);
nor U611 (N_611,In_313,In_403);
nand U612 (N_612,In_593,In_75);
or U613 (N_613,In_91,In_732);
nor U614 (N_614,In_792,In_139);
nor U615 (N_615,In_979,In_79);
nor U616 (N_616,In_934,In_182);
nor U617 (N_617,In_766,In_66);
or U618 (N_618,In_301,In_804);
or U619 (N_619,In_451,In_59);
nor U620 (N_620,In_580,In_117);
or U621 (N_621,In_332,In_650);
nor U622 (N_622,In_366,In_986);
and U623 (N_623,In_140,In_44);
nor U624 (N_624,In_770,In_806);
and U625 (N_625,In_989,In_233);
nand U626 (N_626,In_178,In_401);
or U627 (N_627,In_145,In_488);
nor U628 (N_628,In_794,In_560);
nand U629 (N_629,In_28,In_503);
or U630 (N_630,In_570,In_223);
nand U631 (N_631,In_869,In_450);
and U632 (N_632,In_199,In_836);
xor U633 (N_633,In_844,In_333);
or U634 (N_634,In_351,In_421);
nand U635 (N_635,In_237,In_648);
nand U636 (N_636,In_234,In_65);
and U637 (N_637,In_577,In_944);
nor U638 (N_638,In_747,In_127);
and U639 (N_639,In_840,In_926);
and U640 (N_640,In_660,In_847);
or U641 (N_641,In_148,In_308);
nand U642 (N_642,In_492,In_42);
and U643 (N_643,In_445,In_474);
or U644 (N_644,In_116,In_217);
nor U645 (N_645,In_932,In_447);
nand U646 (N_646,In_553,In_698);
nand U647 (N_647,In_509,In_350);
or U648 (N_648,In_157,In_569);
nand U649 (N_649,In_948,In_276);
nor U650 (N_650,In_665,In_720);
nand U651 (N_651,In_571,In_594);
nand U652 (N_652,In_564,In_893);
nor U653 (N_653,In_822,In_782);
and U654 (N_654,In_719,In_601);
nand U655 (N_655,In_769,In_922);
nand U656 (N_656,In_611,In_251);
or U657 (N_657,In_571,In_297);
nand U658 (N_658,In_366,In_645);
nor U659 (N_659,In_170,In_440);
and U660 (N_660,In_759,In_813);
nor U661 (N_661,In_182,In_399);
nor U662 (N_662,In_761,In_59);
or U663 (N_663,In_240,In_934);
nor U664 (N_664,In_898,In_173);
or U665 (N_665,In_507,In_251);
nand U666 (N_666,In_250,In_586);
or U667 (N_667,In_129,In_295);
nor U668 (N_668,In_169,In_745);
nor U669 (N_669,In_386,In_604);
nand U670 (N_670,In_339,In_174);
or U671 (N_671,In_296,In_677);
or U672 (N_672,In_300,In_985);
or U673 (N_673,In_969,In_270);
nor U674 (N_674,In_521,In_722);
xnor U675 (N_675,In_643,In_65);
and U676 (N_676,In_909,In_87);
or U677 (N_677,In_584,In_482);
and U678 (N_678,In_167,In_611);
or U679 (N_679,In_568,In_894);
or U680 (N_680,In_590,In_267);
and U681 (N_681,In_81,In_87);
nand U682 (N_682,In_661,In_244);
nor U683 (N_683,In_342,In_270);
nor U684 (N_684,In_402,In_639);
nand U685 (N_685,In_851,In_214);
or U686 (N_686,In_492,In_355);
nor U687 (N_687,In_75,In_830);
nand U688 (N_688,In_312,In_181);
nand U689 (N_689,In_589,In_467);
and U690 (N_690,In_818,In_73);
nor U691 (N_691,In_410,In_758);
or U692 (N_692,In_561,In_776);
nor U693 (N_693,In_211,In_149);
and U694 (N_694,In_673,In_590);
nor U695 (N_695,In_806,In_255);
nand U696 (N_696,In_862,In_560);
nand U697 (N_697,In_16,In_451);
nand U698 (N_698,In_862,In_857);
and U699 (N_699,In_490,In_384);
xor U700 (N_700,In_125,In_217);
and U701 (N_701,In_579,In_404);
nand U702 (N_702,In_64,In_554);
and U703 (N_703,In_299,In_157);
or U704 (N_704,In_439,In_756);
nor U705 (N_705,In_774,In_136);
and U706 (N_706,In_350,In_405);
or U707 (N_707,In_229,In_661);
nor U708 (N_708,In_354,In_698);
nor U709 (N_709,In_254,In_556);
nor U710 (N_710,In_991,In_480);
and U711 (N_711,In_878,In_231);
nor U712 (N_712,In_814,In_659);
nand U713 (N_713,In_959,In_206);
nor U714 (N_714,In_129,In_502);
or U715 (N_715,In_25,In_641);
or U716 (N_716,In_674,In_250);
and U717 (N_717,In_495,In_666);
nor U718 (N_718,In_337,In_235);
or U719 (N_719,In_125,In_199);
nor U720 (N_720,In_339,In_695);
and U721 (N_721,In_250,In_190);
or U722 (N_722,In_988,In_68);
or U723 (N_723,In_858,In_605);
or U724 (N_724,In_45,In_317);
and U725 (N_725,In_336,In_499);
and U726 (N_726,In_200,In_642);
nor U727 (N_727,In_345,In_67);
xnor U728 (N_728,In_953,In_511);
and U729 (N_729,In_120,In_942);
or U730 (N_730,In_34,In_537);
nor U731 (N_731,In_970,In_966);
nand U732 (N_732,In_427,In_933);
nor U733 (N_733,In_379,In_60);
nor U734 (N_734,In_481,In_262);
or U735 (N_735,In_468,In_95);
nand U736 (N_736,In_112,In_684);
and U737 (N_737,In_631,In_346);
nand U738 (N_738,In_230,In_254);
nor U739 (N_739,In_389,In_777);
nor U740 (N_740,In_808,In_208);
and U741 (N_741,In_561,In_942);
and U742 (N_742,In_81,In_751);
nor U743 (N_743,In_640,In_985);
nand U744 (N_744,In_432,In_272);
nand U745 (N_745,In_608,In_149);
and U746 (N_746,In_469,In_422);
or U747 (N_747,In_870,In_281);
nor U748 (N_748,In_352,In_382);
or U749 (N_749,In_462,In_191);
and U750 (N_750,In_595,In_766);
nand U751 (N_751,In_643,In_123);
and U752 (N_752,In_290,In_881);
nor U753 (N_753,In_970,In_712);
and U754 (N_754,In_716,In_923);
and U755 (N_755,In_56,In_941);
nor U756 (N_756,In_617,In_455);
or U757 (N_757,In_995,In_216);
nor U758 (N_758,In_813,In_604);
nand U759 (N_759,In_218,In_572);
nor U760 (N_760,In_435,In_913);
nor U761 (N_761,In_549,In_251);
nand U762 (N_762,In_722,In_612);
and U763 (N_763,In_319,In_256);
and U764 (N_764,In_466,In_315);
nand U765 (N_765,In_35,In_711);
and U766 (N_766,In_708,In_23);
and U767 (N_767,In_157,In_670);
and U768 (N_768,In_356,In_693);
and U769 (N_769,In_984,In_433);
nor U770 (N_770,In_292,In_876);
nor U771 (N_771,In_642,In_62);
or U772 (N_772,In_576,In_133);
nand U773 (N_773,In_295,In_771);
nor U774 (N_774,In_14,In_415);
nor U775 (N_775,In_347,In_160);
nand U776 (N_776,In_48,In_174);
or U777 (N_777,In_254,In_710);
nand U778 (N_778,In_137,In_125);
and U779 (N_779,In_347,In_269);
or U780 (N_780,In_856,In_226);
nand U781 (N_781,In_850,In_34);
and U782 (N_782,In_700,In_15);
and U783 (N_783,In_982,In_569);
nor U784 (N_784,In_632,In_394);
nor U785 (N_785,In_265,In_529);
nand U786 (N_786,In_447,In_340);
and U787 (N_787,In_629,In_655);
nor U788 (N_788,In_744,In_515);
or U789 (N_789,In_101,In_724);
nand U790 (N_790,In_50,In_843);
or U791 (N_791,In_130,In_41);
nand U792 (N_792,In_733,In_790);
and U793 (N_793,In_124,In_184);
or U794 (N_794,In_594,In_427);
or U795 (N_795,In_26,In_680);
nand U796 (N_796,In_447,In_403);
or U797 (N_797,In_589,In_305);
nor U798 (N_798,In_121,In_455);
and U799 (N_799,In_401,In_664);
nand U800 (N_800,In_738,In_731);
or U801 (N_801,In_643,In_680);
or U802 (N_802,In_577,In_379);
or U803 (N_803,In_883,In_473);
and U804 (N_804,In_700,In_16);
or U805 (N_805,In_266,In_842);
nand U806 (N_806,In_252,In_833);
and U807 (N_807,In_808,In_143);
and U808 (N_808,In_144,In_143);
and U809 (N_809,In_931,In_55);
nor U810 (N_810,In_953,In_499);
or U811 (N_811,In_268,In_164);
and U812 (N_812,In_434,In_997);
nand U813 (N_813,In_945,In_888);
nor U814 (N_814,In_687,In_85);
and U815 (N_815,In_282,In_457);
nand U816 (N_816,In_887,In_757);
or U817 (N_817,In_996,In_858);
nand U818 (N_818,In_853,In_365);
nor U819 (N_819,In_792,In_545);
or U820 (N_820,In_582,In_588);
or U821 (N_821,In_478,In_71);
or U822 (N_822,In_576,In_750);
or U823 (N_823,In_247,In_353);
nand U824 (N_824,In_993,In_424);
and U825 (N_825,In_378,In_187);
nand U826 (N_826,In_330,In_5);
and U827 (N_827,In_987,In_946);
or U828 (N_828,In_843,In_299);
or U829 (N_829,In_239,In_657);
nand U830 (N_830,In_910,In_358);
nor U831 (N_831,In_33,In_280);
or U832 (N_832,In_714,In_556);
or U833 (N_833,In_216,In_354);
nor U834 (N_834,In_466,In_418);
nand U835 (N_835,In_556,In_25);
or U836 (N_836,In_756,In_599);
nand U837 (N_837,In_21,In_957);
nand U838 (N_838,In_270,In_163);
and U839 (N_839,In_782,In_357);
nor U840 (N_840,In_275,In_179);
nand U841 (N_841,In_282,In_221);
or U842 (N_842,In_539,In_79);
or U843 (N_843,In_729,In_460);
nor U844 (N_844,In_463,In_879);
xor U845 (N_845,In_34,In_545);
and U846 (N_846,In_647,In_248);
and U847 (N_847,In_211,In_867);
and U848 (N_848,In_812,In_358);
xnor U849 (N_849,In_892,In_555);
nand U850 (N_850,In_634,In_681);
and U851 (N_851,In_805,In_44);
nand U852 (N_852,In_565,In_346);
nor U853 (N_853,In_428,In_942);
or U854 (N_854,In_694,In_696);
nand U855 (N_855,In_460,In_546);
or U856 (N_856,In_260,In_880);
or U857 (N_857,In_394,In_335);
nand U858 (N_858,In_263,In_579);
nor U859 (N_859,In_541,In_186);
and U860 (N_860,In_816,In_196);
and U861 (N_861,In_153,In_28);
or U862 (N_862,In_739,In_841);
or U863 (N_863,In_210,In_781);
and U864 (N_864,In_677,In_247);
and U865 (N_865,In_373,In_214);
nor U866 (N_866,In_877,In_260);
nor U867 (N_867,In_573,In_527);
nand U868 (N_868,In_195,In_943);
or U869 (N_869,In_400,In_180);
or U870 (N_870,In_230,In_391);
nor U871 (N_871,In_546,In_891);
nand U872 (N_872,In_407,In_124);
or U873 (N_873,In_850,In_823);
nand U874 (N_874,In_967,In_899);
nand U875 (N_875,In_488,In_289);
or U876 (N_876,In_410,In_504);
or U877 (N_877,In_307,In_945);
or U878 (N_878,In_850,In_809);
nor U879 (N_879,In_760,In_403);
and U880 (N_880,In_468,In_576);
nor U881 (N_881,In_43,In_634);
nor U882 (N_882,In_405,In_508);
nand U883 (N_883,In_878,In_532);
and U884 (N_884,In_734,In_720);
nand U885 (N_885,In_804,In_217);
and U886 (N_886,In_30,In_704);
or U887 (N_887,In_745,In_794);
nand U888 (N_888,In_524,In_247);
or U889 (N_889,In_889,In_337);
or U890 (N_890,In_242,In_995);
xnor U891 (N_891,In_963,In_124);
and U892 (N_892,In_890,In_320);
or U893 (N_893,In_47,In_978);
nor U894 (N_894,In_168,In_958);
nand U895 (N_895,In_38,In_110);
or U896 (N_896,In_408,In_355);
nand U897 (N_897,In_944,In_964);
nand U898 (N_898,In_117,In_567);
or U899 (N_899,In_837,In_651);
and U900 (N_900,In_944,In_966);
and U901 (N_901,In_283,In_251);
and U902 (N_902,In_665,In_386);
or U903 (N_903,In_758,In_358);
nor U904 (N_904,In_898,In_193);
and U905 (N_905,In_906,In_7);
or U906 (N_906,In_504,In_521);
nand U907 (N_907,In_341,In_527);
nor U908 (N_908,In_62,In_559);
nand U909 (N_909,In_270,In_645);
or U910 (N_910,In_174,In_806);
nor U911 (N_911,In_389,In_781);
and U912 (N_912,In_317,In_840);
nor U913 (N_913,In_469,In_389);
nor U914 (N_914,In_89,In_381);
nand U915 (N_915,In_885,In_104);
nand U916 (N_916,In_351,In_641);
and U917 (N_917,In_117,In_672);
and U918 (N_918,In_134,In_239);
nand U919 (N_919,In_706,In_735);
or U920 (N_920,In_311,In_556);
or U921 (N_921,In_472,In_202);
nor U922 (N_922,In_573,In_754);
and U923 (N_923,In_134,In_253);
nand U924 (N_924,In_292,In_305);
and U925 (N_925,In_142,In_969);
and U926 (N_926,In_474,In_321);
nor U927 (N_927,In_245,In_282);
nor U928 (N_928,In_485,In_375);
and U929 (N_929,In_641,In_100);
nand U930 (N_930,In_781,In_273);
and U931 (N_931,In_356,In_450);
nand U932 (N_932,In_340,In_838);
and U933 (N_933,In_169,In_896);
nand U934 (N_934,In_442,In_355);
nand U935 (N_935,In_351,In_247);
nand U936 (N_936,In_49,In_594);
nor U937 (N_937,In_481,In_515);
or U938 (N_938,In_941,In_953);
and U939 (N_939,In_357,In_713);
nand U940 (N_940,In_828,In_237);
and U941 (N_941,In_326,In_596);
or U942 (N_942,In_816,In_571);
and U943 (N_943,In_979,In_95);
nor U944 (N_944,In_348,In_63);
and U945 (N_945,In_271,In_912);
and U946 (N_946,In_262,In_893);
or U947 (N_947,In_590,In_822);
nand U948 (N_948,In_793,In_578);
nand U949 (N_949,In_860,In_105);
and U950 (N_950,In_701,In_680);
nor U951 (N_951,In_555,In_519);
and U952 (N_952,In_762,In_234);
or U953 (N_953,In_291,In_655);
or U954 (N_954,In_819,In_332);
nand U955 (N_955,In_57,In_590);
nor U956 (N_956,In_459,In_43);
or U957 (N_957,In_1,In_135);
nor U958 (N_958,In_973,In_676);
or U959 (N_959,In_187,In_245);
nand U960 (N_960,In_11,In_725);
nor U961 (N_961,In_267,In_283);
nor U962 (N_962,In_144,In_231);
nand U963 (N_963,In_407,In_396);
or U964 (N_964,In_877,In_997);
nand U965 (N_965,In_548,In_236);
and U966 (N_966,In_477,In_78);
and U967 (N_967,In_16,In_160);
and U968 (N_968,In_428,In_657);
or U969 (N_969,In_861,In_578);
or U970 (N_970,In_666,In_921);
and U971 (N_971,In_535,In_814);
nor U972 (N_972,In_311,In_882);
and U973 (N_973,In_758,In_664);
nand U974 (N_974,In_887,In_211);
or U975 (N_975,In_161,In_432);
or U976 (N_976,In_268,In_119);
or U977 (N_977,In_677,In_138);
nor U978 (N_978,In_46,In_140);
nand U979 (N_979,In_87,In_388);
and U980 (N_980,In_414,In_656);
nor U981 (N_981,In_185,In_482);
nand U982 (N_982,In_839,In_364);
nor U983 (N_983,In_792,In_809);
nor U984 (N_984,In_732,In_729);
or U985 (N_985,In_342,In_907);
nand U986 (N_986,In_566,In_12);
or U987 (N_987,In_216,In_589);
nor U988 (N_988,In_703,In_167);
and U989 (N_989,In_668,In_751);
nor U990 (N_990,In_615,In_873);
nand U991 (N_991,In_788,In_136);
and U992 (N_992,In_791,In_467);
and U993 (N_993,In_823,In_582);
nand U994 (N_994,In_274,In_376);
or U995 (N_995,In_236,In_64);
and U996 (N_996,In_183,In_304);
or U997 (N_997,In_288,In_281);
and U998 (N_998,In_246,In_490);
or U999 (N_999,In_848,In_171);
nand U1000 (N_1000,In_689,In_205);
and U1001 (N_1001,In_971,In_399);
nor U1002 (N_1002,In_423,In_124);
and U1003 (N_1003,In_820,In_421);
and U1004 (N_1004,In_318,In_75);
nand U1005 (N_1005,In_247,In_841);
nand U1006 (N_1006,In_845,In_117);
nand U1007 (N_1007,In_63,In_925);
or U1008 (N_1008,In_694,In_628);
and U1009 (N_1009,In_320,In_270);
or U1010 (N_1010,In_621,In_127);
or U1011 (N_1011,In_637,In_810);
and U1012 (N_1012,In_840,In_214);
and U1013 (N_1013,In_124,In_383);
and U1014 (N_1014,In_377,In_154);
nand U1015 (N_1015,In_378,In_333);
nor U1016 (N_1016,In_784,In_143);
and U1017 (N_1017,In_690,In_201);
nand U1018 (N_1018,In_850,In_750);
nor U1019 (N_1019,In_684,In_80);
or U1020 (N_1020,In_712,In_536);
and U1021 (N_1021,In_46,In_961);
nand U1022 (N_1022,In_694,In_21);
or U1023 (N_1023,In_373,In_844);
nor U1024 (N_1024,In_793,In_394);
nand U1025 (N_1025,In_84,In_79);
nand U1026 (N_1026,In_219,In_379);
nand U1027 (N_1027,In_401,In_631);
nand U1028 (N_1028,In_438,In_141);
nand U1029 (N_1029,In_662,In_343);
nand U1030 (N_1030,In_691,In_631);
and U1031 (N_1031,In_116,In_10);
or U1032 (N_1032,In_793,In_693);
and U1033 (N_1033,In_791,In_430);
or U1034 (N_1034,In_625,In_782);
nor U1035 (N_1035,In_793,In_505);
nor U1036 (N_1036,In_525,In_945);
and U1037 (N_1037,In_944,In_458);
nor U1038 (N_1038,In_252,In_50);
nor U1039 (N_1039,In_428,In_623);
and U1040 (N_1040,In_466,In_67);
nand U1041 (N_1041,In_92,In_858);
nor U1042 (N_1042,In_257,In_479);
and U1043 (N_1043,In_404,In_882);
or U1044 (N_1044,In_862,In_484);
or U1045 (N_1045,In_534,In_224);
or U1046 (N_1046,In_851,In_20);
or U1047 (N_1047,In_447,In_569);
nand U1048 (N_1048,In_882,In_933);
nor U1049 (N_1049,In_1,In_846);
nor U1050 (N_1050,In_135,In_187);
nor U1051 (N_1051,In_774,In_561);
nor U1052 (N_1052,In_553,In_615);
nor U1053 (N_1053,In_712,In_241);
xor U1054 (N_1054,In_330,In_383);
nand U1055 (N_1055,In_595,In_753);
and U1056 (N_1056,In_400,In_706);
xor U1057 (N_1057,In_201,In_361);
or U1058 (N_1058,In_294,In_692);
nor U1059 (N_1059,In_162,In_869);
nor U1060 (N_1060,In_869,In_376);
nor U1061 (N_1061,In_45,In_828);
and U1062 (N_1062,In_901,In_515);
or U1063 (N_1063,In_573,In_966);
and U1064 (N_1064,In_786,In_784);
and U1065 (N_1065,In_642,In_627);
nand U1066 (N_1066,In_228,In_445);
and U1067 (N_1067,In_786,In_951);
and U1068 (N_1068,In_23,In_856);
and U1069 (N_1069,In_753,In_625);
nand U1070 (N_1070,In_878,In_400);
nand U1071 (N_1071,In_790,In_544);
nand U1072 (N_1072,In_349,In_4);
or U1073 (N_1073,In_990,In_19);
nand U1074 (N_1074,In_863,In_12);
nor U1075 (N_1075,In_775,In_508);
and U1076 (N_1076,In_860,In_781);
or U1077 (N_1077,In_575,In_510);
and U1078 (N_1078,In_823,In_997);
nor U1079 (N_1079,In_628,In_67);
and U1080 (N_1080,In_620,In_627);
and U1081 (N_1081,In_465,In_21);
nor U1082 (N_1082,In_620,In_30);
or U1083 (N_1083,In_891,In_361);
nand U1084 (N_1084,In_988,In_760);
or U1085 (N_1085,In_724,In_344);
or U1086 (N_1086,In_230,In_382);
and U1087 (N_1087,In_589,In_417);
nand U1088 (N_1088,In_866,In_366);
or U1089 (N_1089,In_951,In_481);
and U1090 (N_1090,In_456,In_269);
and U1091 (N_1091,In_733,In_165);
or U1092 (N_1092,In_512,In_275);
and U1093 (N_1093,In_602,In_32);
nor U1094 (N_1094,In_545,In_239);
nand U1095 (N_1095,In_273,In_52);
and U1096 (N_1096,In_852,In_163);
and U1097 (N_1097,In_582,In_244);
nand U1098 (N_1098,In_376,In_120);
nor U1099 (N_1099,In_292,In_911);
or U1100 (N_1100,In_817,In_285);
or U1101 (N_1101,In_353,In_352);
nand U1102 (N_1102,In_950,In_595);
and U1103 (N_1103,In_592,In_11);
and U1104 (N_1104,In_947,In_527);
or U1105 (N_1105,In_717,In_176);
nor U1106 (N_1106,In_32,In_702);
nand U1107 (N_1107,In_385,In_981);
and U1108 (N_1108,In_357,In_402);
or U1109 (N_1109,In_530,In_281);
or U1110 (N_1110,In_396,In_752);
or U1111 (N_1111,In_142,In_504);
or U1112 (N_1112,In_621,In_550);
nand U1113 (N_1113,In_437,In_850);
nor U1114 (N_1114,In_679,In_736);
and U1115 (N_1115,In_709,In_504);
nand U1116 (N_1116,In_161,In_807);
nor U1117 (N_1117,In_394,In_747);
or U1118 (N_1118,In_609,In_249);
or U1119 (N_1119,In_968,In_183);
nand U1120 (N_1120,In_656,In_451);
and U1121 (N_1121,In_362,In_272);
nor U1122 (N_1122,In_706,In_144);
and U1123 (N_1123,In_576,In_995);
nand U1124 (N_1124,In_967,In_674);
or U1125 (N_1125,In_799,In_592);
or U1126 (N_1126,In_954,In_307);
nand U1127 (N_1127,In_135,In_163);
nand U1128 (N_1128,In_846,In_395);
nand U1129 (N_1129,In_567,In_496);
nor U1130 (N_1130,In_550,In_510);
or U1131 (N_1131,In_590,In_391);
and U1132 (N_1132,In_508,In_421);
and U1133 (N_1133,In_566,In_485);
nor U1134 (N_1134,In_856,In_575);
or U1135 (N_1135,In_821,In_866);
nand U1136 (N_1136,In_225,In_380);
nor U1137 (N_1137,In_869,In_175);
nand U1138 (N_1138,In_866,In_944);
and U1139 (N_1139,In_549,In_55);
nand U1140 (N_1140,In_113,In_459);
or U1141 (N_1141,In_191,In_155);
nand U1142 (N_1142,In_70,In_460);
and U1143 (N_1143,In_968,In_218);
nor U1144 (N_1144,In_677,In_985);
nor U1145 (N_1145,In_428,In_21);
nand U1146 (N_1146,In_674,In_918);
or U1147 (N_1147,In_508,In_265);
nand U1148 (N_1148,In_821,In_176);
nor U1149 (N_1149,In_439,In_702);
nor U1150 (N_1150,In_926,In_2);
or U1151 (N_1151,In_131,In_217);
and U1152 (N_1152,In_340,In_98);
nand U1153 (N_1153,In_888,In_857);
nor U1154 (N_1154,In_112,In_507);
or U1155 (N_1155,In_352,In_455);
or U1156 (N_1156,In_706,In_861);
nor U1157 (N_1157,In_241,In_90);
xnor U1158 (N_1158,In_836,In_636);
and U1159 (N_1159,In_925,In_605);
and U1160 (N_1160,In_411,In_998);
nand U1161 (N_1161,In_112,In_423);
or U1162 (N_1162,In_879,In_586);
nor U1163 (N_1163,In_285,In_993);
or U1164 (N_1164,In_358,In_325);
nand U1165 (N_1165,In_745,In_936);
or U1166 (N_1166,In_54,In_327);
or U1167 (N_1167,In_455,In_276);
nor U1168 (N_1168,In_990,In_731);
nor U1169 (N_1169,In_867,In_302);
nor U1170 (N_1170,In_631,In_461);
nand U1171 (N_1171,In_643,In_21);
or U1172 (N_1172,In_264,In_379);
nor U1173 (N_1173,In_45,In_786);
nor U1174 (N_1174,In_899,In_839);
or U1175 (N_1175,In_186,In_105);
nand U1176 (N_1176,In_223,In_460);
nand U1177 (N_1177,In_710,In_401);
nor U1178 (N_1178,In_324,In_429);
nor U1179 (N_1179,In_342,In_47);
nor U1180 (N_1180,In_390,In_464);
or U1181 (N_1181,In_515,In_650);
nand U1182 (N_1182,In_698,In_965);
nand U1183 (N_1183,In_874,In_535);
and U1184 (N_1184,In_268,In_361);
and U1185 (N_1185,In_481,In_511);
nand U1186 (N_1186,In_788,In_536);
nor U1187 (N_1187,In_370,In_594);
nand U1188 (N_1188,In_289,In_267);
nor U1189 (N_1189,In_889,In_859);
nor U1190 (N_1190,In_14,In_577);
nor U1191 (N_1191,In_483,In_902);
nand U1192 (N_1192,In_251,In_762);
nor U1193 (N_1193,In_374,In_442);
nand U1194 (N_1194,In_685,In_307);
and U1195 (N_1195,In_204,In_546);
and U1196 (N_1196,In_351,In_83);
nor U1197 (N_1197,In_351,In_891);
or U1198 (N_1198,In_692,In_143);
and U1199 (N_1199,In_197,In_191);
nor U1200 (N_1200,In_977,In_876);
nor U1201 (N_1201,In_320,In_695);
nor U1202 (N_1202,In_321,In_325);
and U1203 (N_1203,In_713,In_312);
nor U1204 (N_1204,In_610,In_589);
nand U1205 (N_1205,In_272,In_17);
or U1206 (N_1206,In_227,In_551);
or U1207 (N_1207,In_330,In_474);
nand U1208 (N_1208,In_646,In_436);
nand U1209 (N_1209,In_368,In_106);
xnor U1210 (N_1210,In_728,In_93);
nand U1211 (N_1211,In_301,In_954);
nor U1212 (N_1212,In_478,In_83);
nor U1213 (N_1213,In_176,In_505);
nor U1214 (N_1214,In_697,In_247);
and U1215 (N_1215,In_224,In_853);
nand U1216 (N_1216,In_433,In_332);
or U1217 (N_1217,In_127,In_135);
and U1218 (N_1218,In_130,In_20);
and U1219 (N_1219,In_977,In_375);
nor U1220 (N_1220,In_943,In_12);
nand U1221 (N_1221,In_807,In_125);
or U1222 (N_1222,In_76,In_257);
or U1223 (N_1223,In_875,In_25);
or U1224 (N_1224,In_252,In_391);
nand U1225 (N_1225,In_886,In_772);
nand U1226 (N_1226,In_422,In_983);
and U1227 (N_1227,In_694,In_33);
nand U1228 (N_1228,In_992,In_902);
and U1229 (N_1229,In_525,In_291);
nand U1230 (N_1230,In_45,In_193);
or U1231 (N_1231,In_120,In_784);
nor U1232 (N_1232,In_715,In_74);
or U1233 (N_1233,In_306,In_63);
or U1234 (N_1234,In_697,In_46);
or U1235 (N_1235,In_393,In_939);
and U1236 (N_1236,In_203,In_844);
nand U1237 (N_1237,In_831,In_355);
nor U1238 (N_1238,In_420,In_211);
nor U1239 (N_1239,In_760,In_124);
and U1240 (N_1240,In_211,In_192);
nor U1241 (N_1241,In_209,In_673);
nand U1242 (N_1242,In_754,In_957);
and U1243 (N_1243,In_747,In_734);
nor U1244 (N_1244,In_138,In_455);
nor U1245 (N_1245,In_213,In_698);
nand U1246 (N_1246,In_150,In_179);
nor U1247 (N_1247,In_960,In_478);
nand U1248 (N_1248,In_647,In_352);
nand U1249 (N_1249,In_374,In_971);
or U1250 (N_1250,In_426,In_567);
or U1251 (N_1251,In_124,In_192);
nor U1252 (N_1252,In_628,In_940);
and U1253 (N_1253,In_488,In_466);
or U1254 (N_1254,In_305,In_805);
nand U1255 (N_1255,In_822,In_137);
and U1256 (N_1256,In_200,In_790);
nor U1257 (N_1257,In_542,In_184);
nand U1258 (N_1258,In_847,In_679);
or U1259 (N_1259,In_177,In_863);
nand U1260 (N_1260,In_335,In_200);
and U1261 (N_1261,In_755,In_626);
nor U1262 (N_1262,In_587,In_216);
or U1263 (N_1263,In_15,In_212);
or U1264 (N_1264,In_865,In_254);
nor U1265 (N_1265,In_526,In_82);
nand U1266 (N_1266,In_401,In_332);
nand U1267 (N_1267,In_848,In_444);
nand U1268 (N_1268,In_696,In_100);
nor U1269 (N_1269,In_714,In_876);
and U1270 (N_1270,In_235,In_851);
nand U1271 (N_1271,In_425,In_299);
nand U1272 (N_1272,In_329,In_504);
or U1273 (N_1273,In_59,In_349);
nand U1274 (N_1274,In_914,In_897);
nor U1275 (N_1275,In_311,In_395);
and U1276 (N_1276,In_587,In_853);
nor U1277 (N_1277,In_112,In_935);
xor U1278 (N_1278,In_880,In_502);
or U1279 (N_1279,In_698,In_620);
nand U1280 (N_1280,In_945,In_277);
nor U1281 (N_1281,In_780,In_956);
nand U1282 (N_1282,In_627,In_796);
nor U1283 (N_1283,In_162,In_740);
and U1284 (N_1284,In_786,In_399);
or U1285 (N_1285,In_556,In_963);
or U1286 (N_1286,In_837,In_327);
and U1287 (N_1287,In_743,In_118);
nand U1288 (N_1288,In_536,In_211);
nand U1289 (N_1289,In_687,In_812);
or U1290 (N_1290,In_762,In_465);
nand U1291 (N_1291,In_576,In_588);
or U1292 (N_1292,In_630,In_990);
nor U1293 (N_1293,In_970,In_795);
nor U1294 (N_1294,In_495,In_812);
nor U1295 (N_1295,In_17,In_561);
nor U1296 (N_1296,In_355,In_663);
nor U1297 (N_1297,In_899,In_527);
nand U1298 (N_1298,In_612,In_839);
and U1299 (N_1299,In_849,In_265);
nor U1300 (N_1300,In_777,In_444);
nor U1301 (N_1301,In_9,In_240);
and U1302 (N_1302,In_728,In_50);
nand U1303 (N_1303,In_593,In_9);
and U1304 (N_1304,In_411,In_573);
nor U1305 (N_1305,In_136,In_839);
and U1306 (N_1306,In_871,In_73);
nor U1307 (N_1307,In_346,In_348);
or U1308 (N_1308,In_581,In_715);
nor U1309 (N_1309,In_575,In_205);
nor U1310 (N_1310,In_840,In_691);
and U1311 (N_1311,In_540,In_969);
nor U1312 (N_1312,In_915,In_56);
and U1313 (N_1313,In_964,In_837);
nor U1314 (N_1314,In_93,In_468);
nand U1315 (N_1315,In_544,In_130);
and U1316 (N_1316,In_965,In_558);
nor U1317 (N_1317,In_729,In_601);
nand U1318 (N_1318,In_575,In_976);
nor U1319 (N_1319,In_548,In_721);
nor U1320 (N_1320,In_445,In_261);
nand U1321 (N_1321,In_580,In_591);
nor U1322 (N_1322,In_981,In_191);
or U1323 (N_1323,In_605,In_525);
nand U1324 (N_1324,In_119,In_257);
and U1325 (N_1325,In_425,In_142);
and U1326 (N_1326,In_639,In_124);
nor U1327 (N_1327,In_957,In_328);
nand U1328 (N_1328,In_131,In_226);
nor U1329 (N_1329,In_676,In_331);
or U1330 (N_1330,In_494,In_533);
nand U1331 (N_1331,In_733,In_789);
or U1332 (N_1332,In_752,In_912);
or U1333 (N_1333,In_820,In_22);
or U1334 (N_1334,In_458,In_608);
nor U1335 (N_1335,In_88,In_116);
nand U1336 (N_1336,In_76,In_109);
nor U1337 (N_1337,In_80,In_391);
and U1338 (N_1338,In_66,In_94);
nor U1339 (N_1339,In_626,In_282);
nand U1340 (N_1340,In_189,In_707);
nand U1341 (N_1341,In_298,In_53);
or U1342 (N_1342,In_374,In_262);
nor U1343 (N_1343,In_612,In_675);
nor U1344 (N_1344,In_555,In_316);
nand U1345 (N_1345,In_598,In_503);
nor U1346 (N_1346,In_624,In_509);
or U1347 (N_1347,In_22,In_827);
nor U1348 (N_1348,In_865,In_447);
or U1349 (N_1349,In_917,In_104);
and U1350 (N_1350,In_922,In_22);
and U1351 (N_1351,In_330,In_239);
nor U1352 (N_1352,In_189,In_413);
or U1353 (N_1353,In_251,In_616);
or U1354 (N_1354,In_44,In_455);
or U1355 (N_1355,In_976,In_802);
or U1356 (N_1356,In_236,In_505);
or U1357 (N_1357,In_113,In_808);
nand U1358 (N_1358,In_159,In_269);
and U1359 (N_1359,In_803,In_724);
nand U1360 (N_1360,In_32,In_170);
nor U1361 (N_1361,In_1,In_727);
and U1362 (N_1362,In_354,In_507);
nor U1363 (N_1363,In_516,In_433);
nand U1364 (N_1364,In_444,In_976);
nor U1365 (N_1365,In_342,In_681);
nor U1366 (N_1366,In_263,In_371);
or U1367 (N_1367,In_811,In_319);
or U1368 (N_1368,In_723,In_541);
or U1369 (N_1369,In_244,In_420);
and U1370 (N_1370,In_646,In_146);
nand U1371 (N_1371,In_957,In_489);
and U1372 (N_1372,In_313,In_856);
and U1373 (N_1373,In_319,In_885);
and U1374 (N_1374,In_989,In_663);
or U1375 (N_1375,In_896,In_809);
or U1376 (N_1376,In_386,In_728);
nor U1377 (N_1377,In_664,In_501);
nor U1378 (N_1378,In_301,In_982);
or U1379 (N_1379,In_416,In_115);
nand U1380 (N_1380,In_283,In_659);
nand U1381 (N_1381,In_100,In_84);
or U1382 (N_1382,In_377,In_700);
nor U1383 (N_1383,In_758,In_283);
nand U1384 (N_1384,In_192,In_970);
and U1385 (N_1385,In_689,In_4);
and U1386 (N_1386,In_446,In_491);
nor U1387 (N_1387,In_641,In_230);
nand U1388 (N_1388,In_754,In_698);
nand U1389 (N_1389,In_434,In_477);
nor U1390 (N_1390,In_274,In_36);
nand U1391 (N_1391,In_21,In_761);
nor U1392 (N_1392,In_377,In_362);
and U1393 (N_1393,In_649,In_31);
or U1394 (N_1394,In_502,In_666);
nand U1395 (N_1395,In_977,In_248);
and U1396 (N_1396,In_162,In_178);
nor U1397 (N_1397,In_213,In_404);
or U1398 (N_1398,In_319,In_522);
or U1399 (N_1399,In_212,In_632);
nor U1400 (N_1400,In_572,In_538);
and U1401 (N_1401,In_25,In_396);
or U1402 (N_1402,In_447,In_698);
nand U1403 (N_1403,In_835,In_377);
nand U1404 (N_1404,In_406,In_837);
or U1405 (N_1405,In_228,In_46);
nor U1406 (N_1406,In_495,In_250);
nor U1407 (N_1407,In_792,In_538);
nor U1408 (N_1408,In_82,In_260);
or U1409 (N_1409,In_539,In_756);
and U1410 (N_1410,In_789,In_211);
nand U1411 (N_1411,In_66,In_501);
nand U1412 (N_1412,In_339,In_807);
nor U1413 (N_1413,In_185,In_675);
and U1414 (N_1414,In_90,In_177);
nand U1415 (N_1415,In_473,In_735);
or U1416 (N_1416,In_734,In_984);
and U1417 (N_1417,In_557,In_875);
and U1418 (N_1418,In_361,In_635);
nand U1419 (N_1419,In_316,In_852);
and U1420 (N_1420,In_89,In_386);
nor U1421 (N_1421,In_164,In_736);
nand U1422 (N_1422,In_863,In_791);
nor U1423 (N_1423,In_815,In_666);
or U1424 (N_1424,In_779,In_73);
or U1425 (N_1425,In_956,In_568);
and U1426 (N_1426,In_665,In_641);
nor U1427 (N_1427,In_435,In_757);
and U1428 (N_1428,In_248,In_892);
nand U1429 (N_1429,In_892,In_340);
nand U1430 (N_1430,In_986,In_273);
nand U1431 (N_1431,In_353,In_159);
and U1432 (N_1432,In_953,In_139);
nand U1433 (N_1433,In_232,In_975);
nand U1434 (N_1434,In_286,In_327);
nor U1435 (N_1435,In_482,In_862);
and U1436 (N_1436,In_32,In_993);
nand U1437 (N_1437,In_767,In_20);
and U1438 (N_1438,In_651,In_450);
nand U1439 (N_1439,In_173,In_963);
nand U1440 (N_1440,In_196,In_622);
nor U1441 (N_1441,In_82,In_913);
or U1442 (N_1442,In_50,In_890);
nor U1443 (N_1443,In_895,In_741);
nand U1444 (N_1444,In_346,In_308);
xnor U1445 (N_1445,In_840,In_714);
and U1446 (N_1446,In_853,In_507);
or U1447 (N_1447,In_334,In_339);
nor U1448 (N_1448,In_768,In_783);
nor U1449 (N_1449,In_806,In_183);
nor U1450 (N_1450,In_220,In_783);
nand U1451 (N_1451,In_727,In_204);
nand U1452 (N_1452,In_454,In_383);
and U1453 (N_1453,In_447,In_517);
and U1454 (N_1454,In_184,In_335);
nand U1455 (N_1455,In_788,In_575);
nor U1456 (N_1456,In_662,In_768);
or U1457 (N_1457,In_697,In_410);
xnor U1458 (N_1458,In_333,In_56);
or U1459 (N_1459,In_799,In_16);
nor U1460 (N_1460,In_64,In_243);
nor U1461 (N_1461,In_687,In_509);
or U1462 (N_1462,In_375,In_234);
nor U1463 (N_1463,In_859,In_427);
nor U1464 (N_1464,In_967,In_969);
or U1465 (N_1465,In_960,In_941);
or U1466 (N_1466,In_453,In_422);
nor U1467 (N_1467,In_686,In_42);
nor U1468 (N_1468,In_40,In_108);
nand U1469 (N_1469,In_547,In_348);
nand U1470 (N_1470,In_675,In_863);
or U1471 (N_1471,In_619,In_918);
and U1472 (N_1472,In_400,In_213);
and U1473 (N_1473,In_424,In_808);
or U1474 (N_1474,In_243,In_400);
nand U1475 (N_1475,In_228,In_751);
nor U1476 (N_1476,In_496,In_356);
nor U1477 (N_1477,In_231,In_671);
nand U1478 (N_1478,In_155,In_254);
and U1479 (N_1479,In_915,In_519);
and U1480 (N_1480,In_163,In_513);
or U1481 (N_1481,In_87,In_720);
or U1482 (N_1482,In_746,In_224);
or U1483 (N_1483,In_533,In_633);
or U1484 (N_1484,In_741,In_861);
nor U1485 (N_1485,In_918,In_660);
nor U1486 (N_1486,In_248,In_72);
nand U1487 (N_1487,In_730,In_360);
or U1488 (N_1488,In_173,In_265);
and U1489 (N_1489,In_773,In_191);
nor U1490 (N_1490,In_625,In_370);
and U1491 (N_1491,In_510,In_500);
and U1492 (N_1492,In_250,In_582);
nor U1493 (N_1493,In_635,In_788);
and U1494 (N_1494,In_444,In_857);
or U1495 (N_1495,In_122,In_634);
or U1496 (N_1496,In_693,In_420);
or U1497 (N_1497,In_709,In_353);
nor U1498 (N_1498,In_383,In_647);
and U1499 (N_1499,In_451,In_746);
nand U1500 (N_1500,In_348,In_998);
nor U1501 (N_1501,In_675,In_832);
nand U1502 (N_1502,In_160,In_736);
nor U1503 (N_1503,In_511,In_864);
or U1504 (N_1504,In_176,In_963);
nand U1505 (N_1505,In_578,In_245);
nand U1506 (N_1506,In_939,In_501);
and U1507 (N_1507,In_427,In_739);
nand U1508 (N_1508,In_273,In_979);
or U1509 (N_1509,In_493,In_508);
and U1510 (N_1510,In_695,In_765);
nor U1511 (N_1511,In_849,In_15);
or U1512 (N_1512,In_382,In_762);
nor U1513 (N_1513,In_598,In_954);
nand U1514 (N_1514,In_190,In_107);
nor U1515 (N_1515,In_276,In_513);
or U1516 (N_1516,In_45,In_430);
or U1517 (N_1517,In_954,In_304);
and U1518 (N_1518,In_788,In_205);
nand U1519 (N_1519,In_979,In_523);
nor U1520 (N_1520,In_847,In_605);
and U1521 (N_1521,In_264,In_826);
nor U1522 (N_1522,In_856,In_587);
nor U1523 (N_1523,In_123,In_940);
or U1524 (N_1524,In_783,In_398);
and U1525 (N_1525,In_564,In_520);
or U1526 (N_1526,In_464,In_868);
nand U1527 (N_1527,In_909,In_290);
and U1528 (N_1528,In_222,In_670);
and U1529 (N_1529,In_278,In_946);
nor U1530 (N_1530,In_12,In_959);
and U1531 (N_1531,In_185,In_83);
and U1532 (N_1532,In_814,In_545);
nand U1533 (N_1533,In_355,In_296);
nand U1534 (N_1534,In_307,In_525);
nor U1535 (N_1535,In_988,In_457);
nor U1536 (N_1536,In_978,In_138);
and U1537 (N_1537,In_528,In_983);
or U1538 (N_1538,In_162,In_439);
nor U1539 (N_1539,In_734,In_188);
nor U1540 (N_1540,In_909,In_735);
and U1541 (N_1541,In_544,In_974);
or U1542 (N_1542,In_840,In_584);
or U1543 (N_1543,In_208,In_580);
nor U1544 (N_1544,In_575,In_844);
and U1545 (N_1545,In_716,In_393);
or U1546 (N_1546,In_798,In_374);
nor U1547 (N_1547,In_957,In_110);
and U1548 (N_1548,In_980,In_824);
nand U1549 (N_1549,In_81,In_127);
nor U1550 (N_1550,In_186,In_425);
nor U1551 (N_1551,In_159,In_225);
and U1552 (N_1552,In_853,In_848);
and U1553 (N_1553,In_235,In_266);
and U1554 (N_1554,In_309,In_781);
and U1555 (N_1555,In_701,In_793);
nor U1556 (N_1556,In_906,In_745);
nand U1557 (N_1557,In_104,In_977);
and U1558 (N_1558,In_73,In_655);
nand U1559 (N_1559,In_207,In_867);
and U1560 (N_1560,In_364,In_262);
and U1561 (N_1561,In_111,In_260);
nand U1562 (N_1562,In_866,In_457);
and U1563 (N_1563,In_188,In_95);
or U1564 (N_1564,In_333,In_35);
and U1565 (N_1565,In_888,In_971);
nor U1566 (N_1566,In_77,In_566);
nor U1567 (N_1567,In_248,In_349);
nor U1568 (N_1568,In_856,In_571);
or U1569 (N_1569,In_932,In_459);
and U1570 (N_1570,In_936,In_625);
nand U1571 (N_1571,In_196,In_152);
nand U1572 (N_1572,In_99,In_93);
nor U1573 (N_1573,In_124,In_756);
nor U1574 (N_1574,In_677,In_686);
nor U1575 (N_1575,In_283,In_382);
nor U1576 (N_1576,In_867,In_744);
nand U1577 (N_1577,In_493,In_762);
or U1578 (N_1578,In_326,In_745);
nand U1579 (N_1579,In_355,In_545);
and U1580 (N_1580,In_110,In_152);
nor U1581 (N_1581,In_835,In_26);
and U1582 (N_1582,In_115,In_901);
nand U1583 (N_1583,In_503,In_481);
or U1584 (N_1584,In_764,In_849);
nand U1585 (N_1585,In_79,In_532);
nand U1586 (N_1586,In_657,In_933);
nor U1587 (N_1587,In_300,In_634);
and U1588 (N_1588,In_886,In_132);
nand U1589 (N_1589,In_823,In_133);
nand U1590 (N_1590,In_313,In_42);
or U1591 (N_1591,In_586,In_359);
nand U1592 (N_1592,In_447,In_233);
nor U1593 (N_1593,In_100,In_39);
nor U1594 (N_1594,In_903,In_811);
or U1595 (N_1595,In_31,In_220);
nor U1596 (N_1596,In_118,In_827);
and U1597 (N_1597,In_519,In_122);
or U1598 (N_1598,In_294,In_686);
nand U1599 (N_1599,In_445,In_763);
xnor U1600 (N_1600,In_485,In_584);
or U1601 (N_1601,In_692,In_559);
and U1602 (N_1602,In_413,In_665);
and U1603 (N_1603,In_670,In_107);
nand U1604 (N_1604,In_339,In_176);
nand U1605 (N_1605,In_171,In_653);
nor U1606 (N_1606,In_824,In_260);
and U1607 (N_1607,In_913,In_974);
nor U1608 (N_1608,In_791,In_20);
and U1609 (N_1609,In_37,In_435);
nand U1610 (N_1610,In_975,In_847);
and U1611 (N_1611,In_503,In_190);
nor U1612 (N_1612,In_731,In_736);
nand U1613 (N_1613,In_652,In_48);
nor U1614 (N_1614,In_590,In_302);
nor U1615 (N_1615,In_939,In_311);
nand U1616 (N_1616,In_124,In_628);
nand U1617 (N_1617,In_393,In_381);
nor U1618 (N_1618,In_606,In_612);
nand U1619 (N_1619,In_879,In_487);
and U1620 (N_1620,In_749,In_980);
and U1621 (N_1621,In_729,In_167);
or U1622 (N_1622,In_186,In_872);
or U1623 (N_1623,In_567,In_705);
and U1624 (N_1624,In_63,In_418);
or U1625 (N_1625,In_455,In_490);
nor U1626 (N_1626,In_533,In_9);
and U1627 (N_1627,In_496,In_925);
and U1628 (N_1628,In_829,In_873);
nor U1629 (N_1629,In_235,In_170);
nand U1630 (N_1630,In_847,In_55);
or U1631 (N_1631,In_73,In_386);
or U1632 (N_1632,In_344,In_422);
or U1633 (N_1633,In_244,In_306);
nor U1634 (N_1634,In_307,In_578);
xor U1635 (N_1635,In_767,In_264);
and U1636 (N_1636,In_328,In_400);
or U1637 (N_1637,In_99,In_770);
or U1638 (N_1638,In_657,In_189);
and U1639 (N_1639,In_473,In_611);
nor U1640 (N_1640,In_632,In_890);
nor U1641 (N_1641,In_872,In_199);
nand U1642 (N_1642,In_925,In_986);
nor U1643 (N_1643,In_269,In_718);
and U1644 (N_1644,In_500,In_730);
or U1645 (N_1645,In_819,In_802);
nand U1646 (N_1646,In_628,In_959);
and U1647 (N_1647,In_576,In_298);
or U1648 (N_1648,In_305,In_120);
and U1649 (N_1649,In_55,In_114);
and U1650 (N_1650,In_669,In_412);
or U1651 (N_1651,In_59,In_519);
xor U1652 (N_1652,In_254,In_41);
and U1653 (N_1653,In_35,In_970);
nand U1654 (N_1654,In_631,In_780);
and U1655 (N_1655,In_163,In_998);
and U1656 (N_1656,In_407,In_693);
nor U1657 (N_1657,In_857,In_11);
nand U1658 (N_1658,In_354,In_518);
or U1659 (N_1659,In_608,In_625);
nand U1660 (N_1660,In_942,In_808);
nand U1661 (N_1661,In_588,In_918);
nor U1662 (N_1662,In_121,In_47);
and U1663 (N_1663,In_379,In_944);
or U1664 (N_1664,In_453,In_312);
nand U1665 (N_1665,In_751,In_814);
or U1666 (N_1666,In_215,In_76);
or U1667 (N_1667,In_112,In_473);
nor U1668 (N_1668,In_62,In_199);
nor U1669 (N_1669,In_869,In_599);
and U1670 (N_1670,In_114,In_750);
and U1671 (N_1671,In_682,In_666);
or U1672 (N_1672,In_503,In_882);
and U1673 (N_1673,In_879,In_126);
or U1674 (N_1674,In_166,In_811);
or U1675 (N_1675,In_188,In_748);
nor U1676 (N_1676,In_885,In_838);
nor U1677 (N_1677,In_407,In_339);
nor U1678 (N_1678,In_914,In_278);
and U1679 (N_1679,In_163,In_725);
nor U1680 (N_1680,In_724,In_12);
and U1681 (N_1681,In_771,In_852);
or U1682 (N_1682,In_740,In_710);
nor U1683 (N_1683,In_878,In_529);
or U1684 (N_1684,In_879,In_124);
or U1685 (N_1685,In_652,In_833);
nor U1686 (N_1686,In_611,In_521);
nand U1687 (N_1687,In_645,In_176);
nor U1688 (N_1688,In_141,In_980);
nor U1689 (N_1689,In_85,In_9);
or U1690 (N_1690,In_601,In_57);
and U1691 (N_1691,In_374,In_294);
nand U1692 (N_1692,In_789,In_177);
and U1693 (N_1693,In_291,In_951);
nand U1694 (N_1694,In_734,In_290);
nand U1695 (N_1695,In_624,In_8);
and U1696 (N_1696,In_916,In_911);
nor U1697 (N_1697,In_33,In_599);
nand U1698 (N_1698,In_726,In_849);
and U1699 (N_1699,In_750,In_507);
and U1700 (N_1700,In_916,In_467);
or U1701 (N_1701,In_751,In_349);
nor U1702 (N_1702,In_810,In_864);
nand U1703 (N_1703,In_882,In_427);
nor U1704 (N_1704,In_289,In_41);
and U1705 (N_1705,In_623,In_75);
nor U1706 (N_1706,In_427,In_515);
nor U1707 (N_1707,In_568,In_864);
nand U1708 (N_1708,In_164,In_640);
and U1709 (N_1709,In_242,In_504);
and U1710 (N_1710,In_469,In_683);
and U1711 (N_1711,In_728,In_378);
and U1712 (N_1712,In_499,In_660);
or U1713 (N_1713,In_466,In_772);
nand U1714 (N_1714,In_549,In_597);
nand U1715 (N_1715,In_982,In_18);
nand U1716 (N_1716,In_112,In_969);
and U1717 (N_1717,In_177,In_1);
or U1718 (N_1718,In_182,In_47);
and U1719 (N_1719,In_101,In_148);
nor U1720 (N_1720,In_261,In_557);
nor U1721 (N_1721,In_662,In_264);
and U1722 (N_1722,In_55,In_421);
or U1723 (N_1723,In_999,In_59);
nor U1724 (N_1724,In_732,In_43);
nor U1725 (N_1725,In_993,In_749);
nor U1726 (N_1726,In_368,In_619);
nor U1727 (N_1727,In_746,In_993);
nor U1728 (N_1728,In_850,In_245);
nand U1729 (N_1729,In_877,In_767);
nor U1730 (N_1730,In_188,In_801);
or U1731 (N_1731,In_870,In_771);
or U1732 (N_1732,In_828,In_883);
or U1733 (N_1733,In_122,In_147);
nor U1734 (N_1734,In_967,In_35);
or U1735 (N_1735,In_660,In_484);
or U1736 (N_1736,In_898,In_585);
nand U1737 (N_1737,In_845,In_932);
nand U1738 (N_1738,In_719,In_998);
nand U1739 (N_1739,In_647,In_307);
nor U1740 (N_1740,In_103,In_472);
and U1741 (N_1741,In_447,In_798);
nand U1742 (N_1742,In_670,In_927);
and U1743 (N_1743,In_554,In_225);
and U1744 (N_1744,In_696,In_974);
nand U1745 (N_1745,In_435,In_321);
or U1746 (N_1746,In_805,In_758);
or U1747 (N_1747,In_225,In_165);
nor U1748 (N_1748,In_770,In_445);
nand U1749 (N_1749,In_653,In_177);
and U1750 (N_1750,In_512,In_877);
nand U1751 (N_1751,In_829,In_833);
nand U1752 (N_1752,In_544,In_91);
xor U1753 (N_1753,In_94,In_184);
and U1754 (N_1754,In_404,In_610);
nor U1755 (N_1755,In_687,In_972);
nor U1756 (N_1756,In_168,In_367);
or U1757 (N_1757,In_958,In_559);
or U1758 (N_1758,In_641,In_289);
or U1759 (N_1759,In_304,In_407);
nand U1760 (N_1760,In_916,In_353);
and U1761 (N_1761,In_913,In_629);
nand U1762 (N_1762,In_530,In_217);
or U1763 (N_1763,In_679,In_986);
or U1764 (N_1764,In_274,In_111);
nand U1765 (N_1765,In_713,In_17);
and U1766 (N_1766,In_463,In_875);
and U1767 (N_1767,In_6,In_521);
and U1768 (N_1768,In_848,In_643);
or U1769 (N_1769,In_963,In_238);
and U1770 (N_1770,In_326,In_634);
nor U1771 (N_1771,In_593,In_774);
and U1772 (N_1772,In_622,In_401);
and U1773 (N_1773,In_541,In_307);
or U1774 (N_1774,In_375,In_373);
or U1775 (N_1775,In_513,In_310);
nor U1776 (N_1776,In_43,In_223);
nor U1777 (N_1777,In_218,In_737);
nor U1778 (N_1778,In_377,In_754);
nand U1779 (N_1779,In_806,In_583);
nor U1780 (N_1780,In_710,In_539);
or U1781 (N_1781,In_899,In_237);
nor U1782 (N_1782,In_197,In_697);
nand U1783 (N_1783,In_886,In_700);
nor U1784 (N_1784,In_766,In_904);
nor U1785 (N_1785,In_366,In_199);
or U1786 (N_1786,In_326,In_163);
or U1787 (N_1787,In_975,In_697);
nand U1788 (N_1788,In_827,In_662);
nand U1789 (N_1789,In_196,In_494);
xor U1790 (N_1790,In_140,In_998);
and U1791 (N_1791,In_120,In_629);
and U1792 (N_1792,In_282,In_658);
nand U1793 (N_1793,In_105,In_557);
nand U1794 (N_1794,In_104,In_422);
and U1795 (N_1795,In_757,In_545);
nand U1796 (N_1796,In_858,In_278);
and U1797 (N_1797,In_262,In_871);
and U1798 (N_1798,In_950,In_144);
or U1799 (N_1799,In_523,In_267);
nor U1800 (N_1800,In_725,In_657);
and U1801 (N_1801,In_602,In_855);
nand U1802 (N_1802,In_54,In_794);
or U1803 (N_1803,In_183,In_94);
nand U1804 (N_1804,In_62,In_285);
or U1805 (N_1805,In_816,In_19);
nand U1806 (N_1806,In_139,In_444);
or U1807 (N_1807,In_833,In_987);
nand U1808 (N_1808,In_425,In_200);
nand U1809 (N_1809,In_14,In_375);
nand U1810 (N_1810,In_438,In_50);
nor U1811 (N_1811,In_231,In_326);
nor U1812 (N_1812,In_322,In_780);
nand U1813 (N_1813,In_89,In_436);
nor U1814 (N_1814,In_885,In_123);
or U1815 (N_1815,In_444,In_248);
or U1816 (N_1816,In_901,In_329);
or U1817 (N_1817,In_845,In_913);
or U1818 (N_1818,In_82,In_614);
and U1819 (N_1819,In_480,In_338);
nor U1820 (N_1820,In_48,In_419);
nor U1821 (N_1821,In_786,In_681);
and U1822 (N_1822,In_798,In_99);
or U1823 (N_1823,In_643,In_420);
nor U1824 (N_1824,In_723,In_439);
or U1825 (N_1825,In_640,In_680);
nor U1826 (N_1826,In_511,In_63);
or U1827 (N_1827,In_208,In_65);
nand U1828 (N_1828,In_898,In_179);
or U1829 (N_1829,In_489,In_551);
or U1830 (N_1830,In_722,In_21);
or U1831 (N_1831,In_381,In_792);
nor U1832 (N_1832,In_914,In_665);
or U1833 (N_1833,In_44,In_513);
and U1834 (N_1834,In_475,In_790);
and U1835 (N_1835,In_700,In_79);
or U1836 (N_1836,In_419,In_373);
or U1837 (N_1837,In_984,In_372);
nand U1838 (N_1838,In_898,In_527);
nor U1839 (N_1839,In_469,In_492);
nor U1840 (N_1840,In_706,In_49);
nand U1841 (N_1841,In_108,In_95);
nand U1842 (N_1842,In_602,In_164);
and U1843 (N_1843,In_90,In_41);
and U1844 (N_1844,In_555,In_105);
nor U1845 (N_1845,In_194,In_354);
nor U1846 (N_1846,In_643,In_100);
nand U1847 (N_1847,In_737,In_54);
or U1848 (N_1848,In_71,In_321);
nand U1849 (N_1849,In_705,In_521);
nor U1850 (N_1850,In_346,In_2);
and U1851 (N_1851,In_837,In_65);
nand U1852 (N_1852,In_781,In_908);
and U1853 (N_1853,In_236,In_739);
and U1854 (N_1854,In_983,In_843);
or U1855 (N_1855,In_633,In_162);
and U1856 (N_1856,In_338,In_687);
and U1857 (N_1857,In_207,In_213);
nor U1858 (N_1858,In_330,In_722);
and U1859 (N_1859,In_140,In_640);
nor U1860 (N_1860,In_222,In_116);
nand U1861 (N_1861,In_682,In_192);
or U1862 (N_1862,In_402,In_687);
or U1863 (N_1863,In_396,In_162);
nand U1864 (N_1864,In_548,In_297);
nand U1865 (N_1865,In_988,In_372);
or U1866 (N_1866,In_179,In_691);
nand U1867 (N_1867,In_80,In_884);
nand U1868 (N_1868,In_133,In_740);
nand U1869 (N_1869,In_925,In_834);
nor U1870 (N_1870,In_387,In_363);
and U1871 (N_1871,In_718,In_641);
nand U1872 (N_1872,In_587,In_766);
or U1873 (N_1873,In_475,In_807);
and U1874 (N_1874,In_285,In_556);
nor U1875 (N_1875,In_692,In_280);
and U1876 (N_1876,In_603,In_787);
or U1877 (N_1877,In_421,In_573);
or U1878 (N_1878,In_445,In_904);
nor U1879 (N_1879,In_499,In_84);
nand U1880 (N_1880,In_717,In_26);
and U1881 (N_1881,In_883,In_341);
nor U1882 (N_1882,In_869,In_24);
or U1883 (N_1883,In_607,In_652);
or U1884 (N_1884,In_366,In_884);
nor U1885 (N_1885,In_743,In_95);
and U1886 (N_1886,In_560,In_694);
nor U1887 (N_1887,In_892,In_616);
nand U1888 (N_1888,In_837,In_169);
or U1889 (N_1889,In_715,In_860);
nor U1890 (N_1890,In_756,In_23);
or U1891 (N_1891,In_603,In_191);
nor U1892 (N_1892,In_244,In_936);
nor U1893 (N_1893,In_788,In_150);
and U1894 (N_1894,In_485,In_998);
nor U1895 (N_1895,In_84,In_395);
nor U1896 (N_1896,In_390,In_558);
or U1897 (N_1897,In_454,In_582);
nor U1898 (N_1898,In_295,In_757);
and U1899 (N_1899,In_701,In_133);
nor U1900 (N_1900,In_687,In_232);
and U1901 (N_1901,In_37,In_676);
nor U1902 (N_1902,In_336,In_26);
and U1903 (N_1903,In_125,In_760);
or U1904 (N_1904,In_92,In_212);
xnor U1905 (N_1905,In_295,In_635);
nand U1906 (N_1906,In_987,In_759);
nand U1907 (N_1907,In_644,In_490);
and U1908 (N_1908,In_166,In_136);
nand U1909 (N_1909,In_865,In_520);
nor U1910 (N_1910,In_113,In_884);
nor U1911 (N_1911,In_106,In_977);
and U1912 (N_1912,In_291,In_638);
or U1913 (N_1913,In_432,In_238);
and U1914 (N_1914,In_77,In_355);
nand U1915 (N_1915,In_855,In_491);
nor U1916 (N_1916,In_475,In_735);
nor U1917 (N_1917,In_522,In_750);
or U1918 (N_1918,In_998,In_331);
or U1919 (N_1919,In_29,In_984);
or U1920 (N_1920,In_604,In_942);
nor U1921 (N_1921,In_421,In_558);
or U1922 (N_1922,In_916,In_594);
nor U1923 (N_1923,In_33,In_321);
nor U1924 (N_1924,In_998,In_441);
nor U1925 (N_1925,In_843,In_242);
nand U1926 (N_1926,In_612,In_771);
and U1927 (N_1927,In_963,In_42);
nand U1928 (N_1928,In_494,In_66);
nor U1929 (N_1929,In_762,In_867);
nand U1930 (N_1930,In_196,In_614);
nor U1931 (N_1931,In_45,In_645);
and U1932 (N_1932,In_809,In_844);
nor U1933 (N_1933,In_444,In_629);
nor U1934 (N_1934,In_53,In_926);
and U1935 (N_1935,In_66,In_178);
and U1936 (N_1936,In_329,In_643);
and U1937 (N_1937,In_901,In_324);
nand U1938 (N_1938,In_230,In_643);
nor U1939 (N_1939,In_563,In_517);
nor U1940 (N_1940,In_636,In_200);
nor U1941 (N_1941,In_213,In_75);
nor U1942 (N_1942,In_232,In_772);
nand U1943 (N_1943,In_696,In_620);
and U1944 (N_1944,In_691,In_138);
and U1945 (N_1945,In_643,In_247);
nor U1946 (N_1946,In_379,In_419);
nand U1947 (N_1947,In_886,In_694);
and U1948 (N_1948,In_638,In_535);
nand U1949 (N_1949,In_437,In_827);
nand U1950 (N_1950,In_458,In_765);
or U1951 (N_1951,In_516,In_745);
and U1952 (N_1952,In_257,In_937);
nor U1953 (N_1953,In_741,In_199);
nand U1954 (N_1954,In_456,In_628);
or U1955 (N_1955,In_850,In_828);
or U1956 (N_1956,In_323,In_377);
and U1957 (N_1957,In_693,In_553);
nand U1958 (N_1958,In_355,In_145);
or U1959 (N_1959,In_80,In_81);
nor U1960 (N_1960,In_776,In_62);
or U1961 (N_1961,In_24,In_2);
nor U1962 (N_1962,In_182,In_815);
and U1963 (N_1963,In_960,In_94);
nand U1964 (N_1964,In_324,In_129);
xnor U1965 (N_1965,In_117,In_515);
and U1966 (N_1966,In_769,In_834);
nor U1967 (N_1967,In_559,In_860);
or U1968 (N_1968,In_640,In_637);
nand U1969 (N_1969,In_504,In_431);
nand U1970 (N_1970,In_648,In_879);
nand U1971 (N_1971,In_299,In_251);
nand U1972 (N_1972,In_39,In_328);
or U1973 (N_1973,In_405,In_816);
nor U1974 (N_1974,In_379,In_583);
nand U1975 (N_1975,In_462,In_900);
nor U1976 (N_1976,In_615,In_325);
nand U1977 (N_1977,In_477,In_482);
or U1978 (N_1978,In_696,In_482);
nor U1979 (N_1979,In_106,In_966);
or U1980 (N_1980,In_173,In_255);
nor U1981 (N_1981,In_44,In_366);
nor U1982 (N_1982,In_326,In_971);
or U1983 (N_1983,In_346,In_691);
or U1984 (N_1984,In_212,In_946);
nor U1985 (N_1985,In_4,In_508);
nand U1986 (N_1986,In_410,In_164);
or U1987 (N_1987,In_429,In_793);
and U1988 (N_1988,In_871,In_604);
and U1989 (N_1989,In_576,In_530);
nor U1990 (N_1990,In_612,In_451);
and U1991 (N_1991,In_880,In_541);
and U1992 (N_1992,In_124,In_38);
nor U1993 (N_1993,In_254,In_603);
xor U1994 (N_1994,In_423,In_687);
and U1995 (N_1995,In_743,In_247);
nor U1996 (N_1996,In_380,In_621);
and U1997 (N_1997,In_990,In_113);
nand U1998 (N_1998,In_800,In_343);
nor U1999 (N_1999,In_129,In_13);
nand U2000 (N_2000,In_979,In_88);
nor U2001 (N_2001,In_279,In_784);
or U2002 (N_2002,In_325,In_425);
nor U2003 (N_2003,In_86,In_797);
and U2004 (N_2004,In_528,In_98);
nand U2005 (N_2005,In_146,In_730);
and U2006 (N_2006,In_326,In_678);
and U2007 (N_2007,In_618,In_617);
and U2008 (N_2008,In_533,In_851);
or U2009 (N_2009,In_176,In_264);
and U2010 (N_2010,In_320,In_99);
nor U2011 (N_2011,In_515,In_780);
or U2012 (N_2012,In_782,In_43);
and U2013 (N_2013,In_440,In_89);
or U2014 (N_2014,In_547,In_719);
nor U2015 (N_2015,In_455,In_384);
nor U2016 (N_2016,In_137,In_88);
nor U2017 (N_2017,In_209,In_152);
nor U2018 (N_2018,In_988,In_940);
xnor U2019 (N_2019,In_124,In_548);
nor U2020 (N_2020,In_884,In_254);
and U2021 (N_2021,In_842,In_279);
and U2022 (N_2022,In_19,In_956);
or U2023 (N_2023,In_722,In_662);
nor U2024 (N_2024,In_880,In_134);
xor U2025 (N_2025,In_641,In_656);
nor U2026 (N_2026,In_566,In_903);
or U2027 (N_2027,In_307,In_606);
nor U2028 (N_2028,In_595,In_117);
nand U2029 (N_2029,In_619,In_538);
and U2030 (N_2030,In_95,In_78);
or U2031 (N_2031,In_947,In_604);
nand U2032 (N_2032,In_879,In_455);
nand U2033 (N_2033,In_47,In_225);
nor U2034 (N_2034,In_348,In_994);
and U2035 (N_2035,In_918,In_921);
nand U2036 (N_2036,In_838,In_250);
or U2037 (N_2037,In_377,In_533);
and U2038 (N_2038,In_500,In_578);
nor U2039 (N_2039,In_955,In_258);
and U2040 (N_2040,In_590,In_693);
nand U2041 (N_2041,In_131,In_510);
or U2042 (N_2042,In_639,In_874);
or U2043 (N_2043,In_410,In_818);
nand U2044 (N_2044,In_49,In_542);
nand U2045 (N_2045,In_69,In_890);
or U2046 (N_2046,In_558,In_203);
or U2047 (N_2047,In_409,In_289);
or U2048 (N_2048,In_590,In_730);
nand U2049 (N_2049,In_618,In_675);
nand U2050 (N_2050,In_943,In_185);
nor U2051 (N_2051,In_562,In_834);
or U2052 (N_2052,In_474,In_500);
or U2053 (N_2053,In_341,In_835);
nor U2054 (N_2054,In_768,In_397);
nand U2055 (N_2055,In_180,In_315);
or U2056 (N_2056,In_495,In_48);
nand U2057 (N_2057,In_597,In_440);
or U2058 (N_2058,In_310,In_890);
nand U2059 (N_2059,In_263,In_871);
or U2060 (N_2060,In_683,In_829);
and U2061 (N_2061,In_714,In_934);
nand U2062 (N_2062,In_762,In_282);
nand U2063 (N_2063,In_770,In_199);
nor U2064 (N_2064,In_25,In_44);
nor U2065 (N_2065,In_464,In_354);
and U2066 (N_2066,In_55,In_692);
nand U2067 (N_2067,In_44,In_143);
and U2068 (N_2068,In_152,In_651);
nor U2069 (N_2069,In_74,In_333);
nand U2070 (N_2070,In_54,In_678);
or U2071 (N_2071,In_468,In_109);
nand U2072 (N_2072,In_543,In_927);
and U2073 (N_2073,In_318,In_535);
and U2074 (N_2074,In_503,In_835);
nand U2075 (N_2075,In_345,In_693);
or U2076 (N_2076,In_29,In_666);
or U2077 (N_2077,In_14,In_260);
or U2078 (N_2078,In_867,In_279);
or U2079 (N_2079,In_542,In_158);
or U2080 (N_2080,In_48,In_761);
nand U2081 (N_2081,In_410,In_524);
or U2082 (N_2082,In_734,In_399);
or U2083 (N_2083,In_149,In_961);
or U2084 (N_2084,In_916,In_243);
or U2085 (N_2085,In_141,In_837);
and U2086 (N_2086,In_340,In_862);
and U2087 (N_2087,In_386,In_164);
nand U2088 (N_2088,In_357,In_701);
and U2089 (N_2089,In_335,In_130);
nand U2090 (N_2090,In_881,In_388);
nand U2091 (N_2091,In_878,In_592);
nor U2092 (N_2092,In_246,In_468);
nor U2093 (N_2093,In_551,In_185);
or U2094 (N_2094,In_870,In_167);
or U2095 (N_2095,In_691,In_425);
nand U2096 (N_2096,In_311,In_216);
and U2097 (N_2097,In_413,In_742);
and U2098 (N_2098,In_802,In_36);
nand U2099 (N_2099,In_297,In_172);
nand U2100 (N_2100,In_98,In_618);
nor U2101 (N_2101,In_191,In_291);
nor U2102 (N_2102,In_86,In_753);
nor U2103 (N_2103,In_40,In_842);
and U2104 (N_2104,In_191,In_690);
or U2105 (N_2105,In_853,In_171);
nor U2106 (N_2106,In_398,In_721);
and U2107 (N_2107,In_321,In_92);
or U2108 (N_2108,In_627,In_389);
and U2109 (N_2109,In_408,In_144);
nand U2110 (N_2110,In_559,In_818);
or U2111 (N_2111,In_198,In_766);
or U2112 (N_2112,In_324,In_188);
nor U2113 (N_2113,In_601,In_327);
or U2114 (N_2114,In_692,In_119);
and U2115 (N_2115,In_282,In_673);
and U2116 (N_2116,In_662,In_185);
nor U2117 (N_2117,In_350,In_759);
nand U2118 (N_2118,In_925,In_480);
nor U2119 (N_2119,In_812,In_614);
nor U2120 (N_2120,In_610,In_651);
nor U2121 (N_2121,In_370,In_520);
and U2122 (N_2122,In_811,In_803);
nor U2123 (N_2123,In_712,In_800);
and U2124 (N_2124,In_492,In_310);
and U2125 (N_2125,In_227,In_934);
nor U2126 (N_2126,In_133,In_231);
nand U2127 (N_2127,In_891,In_459);
or U2128 (N_2128,In_435,In_33);
nor U2129 (N_2129,In_587,In_133);
and U2130 (N_2130,In_864,In_573);
nor U2131 (N_2131,In_372,In_382);
nand U2132 (N_2132,In_385,In_690);
nor U2133 (N_2133,In_553,In_900);
and U2134 (N_2134,In_275,In_142);
and U2135 (N_2135,In_775,In_945);
or U2136 (N_2136,In_221,In_590);
nor U2137 (N_2137,In_624,In_908);
and U2138 (N_2138,In_334,In_367);
or U2139 (N_2139,In_193,In_377);
nor U2140 (N_2140,In_764,In_863);
or U2141 (N_2141,In_572,In_176);
and U2142 (N_2142,In_313,In_567);
nor U2143 (N_2143,In_896,In_469);
or U2144 (N_2144,In_671,In_821);
nand U2145 (N_2145,In_539,In_489);
nor U2146 (N_2146,In_235,In_254);
nand U2147 (N_2147,In_165,In_298);
nor U2148 (N_2148,In_7,In_247);
nand U2149 (N_2149,In_322,In_169);
and U2150 (N_2150,In_184,In_556);
and U2151 (N_2151,In_941,In_15);
and U2152 (N_2152,In_592,In_810);
and U2153 (N_2153,In_753,In_396);
nor U2154 (N_2154,In_121,In_45);
or U2155 (N_2155,In_896,In_806);
nand U2156 (N_2156,In_91,In_175);
nand U2157 (N_2157,In_651,In_740);
nand U2158 (N_2158,In_509,In_303);
nand U2159 (N_2159,In_568,In_31);
and U2160 (N_2160,In_598,In_274);
or U2161 (N_2161,In_330,In_131);
nand U2162 (N_2162,In_833,In_415);
and U2163 (N_2163,In_783,In_885);
nor U2164 (N_2164,In_124,In_60);
or U2165 (N_2165,In_214,In_229);
or U2166 (N_2166,In_743,In_940);
nand U2167 (N_2167,In_415,In_654);
or U2168 (N_2168,In_31,In_533);
or U2169 (N_2169,In_668,In_733);
nand U2170 (N_2170,In_628,In_699);
nor U2171 (N_2171,In_686,In_19);
nand U2172 (N_2172,In_762,In_223);
and U2173 (N_2173,In_4,In_743);
or U2174 (N_2174,In_408,In_927);
nor U2175 (N_2175,In_586,In_873);
nor U2176 (N_2176,In_679,In_821);
or U2177 (N_2177,In_291,In_98);
nand U2178 (N_2178,In_909,In_63);
nor U2179 (N_2179,In_130,In_219);
or U2180 (N_2180,In_39,In_9);
or U2181 (N_2181,In_52,In_262);
nand U2182 (N_2182,In_268,In_400);
nor U2183 (N_2183,In_88,In_529);
nor U2184 (N_2184,In_662,In_15);
nor U2185 (N_2185,In_770,In_205);
nand U2186 (N_2186,In_10,In_161);
or U2187 (N_2187,In_817,In_635);
or U2188 (N_2188,In_978,In_768);
nor U2189 (N_2189,In_206,In_828);
and U2190 (N_2190,In_73,In_540);
or U2191 (N_2191,In_597,In_866);
and U2192 (N_2192,In_140,In_353);
and U2193 (N_2193,In_54,In_699);
nor U2194 (N_2194,In_307,In_120);
and U2195 (N_2195,In_267,In_617);
or U2196 (N_2196,In_921,In_752);
and U2197 (N_2197,In_617,In_242);
xor U2198 (N_2198,In_230,In_512);
nand U2199 (N_2199,In_324,In_305);
or U2200 (N_2200,In_953,In_918);
or U2201 (N_2201,In_726,In_170);
xor U2202 (N_2202,In_413,In_685);
and U2203 (N_2203,In_828,In_55);
nand U2204 (N_2204,In_97,In_703);
and U2205 (N_2205,In_196,In_736);
nor U2206 (N_2206,In_876,In_444);
and U2207 (N_2207,In_858,In_699);
nand U2208 (N_2208,In_657,In_507);
nor U2209 (N_2209,In_111,In_778);
and U2210 (N_2210,In_387,In_508);
nor U2211 (N_2211,In_393,In_441);
and U2212 (N_2212,In_787,In_432);
and U2213 (N_2213,In_613,In_247);
nand U2214 (N_2214,In_803,In_901);
nor U2215 (N_2215,In_179,In_919);
nand U2216 (N_2216,In_110,In_21);
nand U2217 (N_2217,In_240,In_184);
and U2218 (N_2218,In_216,In_850);
or U2219 (N_2219,In_365,In_168);
or U2220 (N_2220,In_346,In_127);
or U2221 (N_2221,In_815,In_805);
nand U2222 (N_2222,In_342,In_720);
and U2223 (N_2223,In_913,In_91);
or U2224 (N_2224,In_628,In_777);
nor U2225 (N_2225,In_882,In_32);
nand U2226 (N_2226,In_992,In_866);
or U2227 (N_2227,In_565,In_480);
nor U2228 (N_2228,In_658,In_637);
nand U2229 (N_2229,In_156,In_656);
or U2230 (N_2230,In_856,In_432);
or U2231 (N_2231,In_899,In_792);
nor U2232 (N_2232,In_911,In_15);
and U2233 (N_2233,In_375,In_158);
and U2234 (N_2234,In_521,In_745);
nand U2235 (N_2235,In_973,In_439);
and U2236 (N_2236,In_130,In_996);
nor U2237 (N_2237,In_966,In_805);
nand U2238 (N_2238,In_638,In_996);
or U2239 (N_2239,In_365,In_69);
nor U2240 (N_2240,In_58,In_507);
nor U2241 (N_2241,In_14,In_480);
nand U2242 (N_2242,In_938,In_558);
xnor U2243 (N_2243,In_853,In_142);
or U2244 (N_2244,In_829,In_201);
nand U2245 (N_2245,In_257,In_401);
nand U2246 (N_2246,In_837,In_631);
and U2247 (N_2247,In_305,In_428);
nor U2248 (N_2248,In_373,In_984);
nor U2249 (N_2249,In_417,In_797);
and U2250 (N_2250,In_113,In_851);
and U2251 (N_2251,In_754,In_848);
and U2252 (N_2252,In_992,In_7);
nand U2253 (N_2253,In_552,In_285);
or U2254 (N_2254,In_199,In_560);
or U2255 (N_2255,In_23,In_305);
nor U2256 (N_2256,In_535,In_465);
and U2257 (N_2257,In_103,In_362);
or U2258 (N_2258,In_257,In_682);
or U2259 (N_2259,In_609,In_954);
nand U2260 (N_2260,In_870,In_754);
and U2261 (N_2261,In_873,In_79);
nor U2262 (N_2262,In_265,In_667);
nand U2263 (N_2263,In_824,In_764);
or U2264 (N_2264,In_919,In_202);
nand U2265 (N_2265,In_963,In_824);
or U2266 (N_2266,In_975,In_695);
nand U2267 (N_2267,In_933,In_410);
and U2268 (N_2268,In_912,In_208);
nand U2269 (N_2269,In_952,In_332);
nor U2270 (N_2270,In_670,In_161);
or U2271 (N_2271,In_127,In_408);
and U2272 (N_2272,In_206,In_436);
or U2273 (N_2273,In_768,In_520);
or U2274 (N_2274,In_473,In_476);
nor U2275 (N_2275,In_512,In_753);
nor U2276 (N_2276,In_454,In_847);
nor U2277 (N_2277,In_5,In_908);
nand U2278 (N_2278,In_354,In_212);
nand U2279 (N_2279,In_217,In_320);
and U2280 (N_2280,In_983,In_859);
and U2281 (N_2281,In_429,In_203);
and U2282 (N_2282,In_777,In_179);
nand U2283 (N_2283,In_963,In_822);
nor U2284 (N_2284,In_675,In_280);
or U2285 (N_2285,In_56,In_316);
nand U2286 (N_2286,In_318,In_927);
nor U2287 (N_2287,In_56,In_995);
or U2288 (N_2288,In_669,In_79);
or U2289 (N_2289,In_409,In_664);
and U2290 (N_2290,In_710,In_768);
nand U2291 (N_2291,In_952,In_689);
nor U2292 (N_2292,In_950,In_515);
and U2293 (N_2293,In_724,In_822);
or U2294 (N_2294,In_604,In_433);
or U2295 (N_2295,In_88,In_537);
or U2296 (N_2296,In_965,In_384);
nand U2297 (N_2297,In_766,In_787);
or U2298 (N_2298,In_141,In_214);
or U2299 (N_2299,In_886,In_162);
nand U2300 (N_2300,In_281,In_858);
nand U2301 (N_2301,In_271,In_159);
or U2302 (N_2302,In_108,In_794);
xor U2303 (N_2303,In_653,In_419);
and U2304 (N_2304,In_608,In_577);
and U2305 (N_2305,In_745,In_71);
or U2306 (N_2306,In_377,In_359);
nand U2307 (N_2307,In_762,In_351);
nor U2308 (N_2308,In_823,In_324);
or U2309 (N_2309,In_396,In_246);
nor U2310 (N_2310,In_541,In_630);
and U2311 (N_2311,In_547,In_863);
or U2312 (N_2312,In_801,In_811);
nor U2313 (N_2313,In_97,In_777);
and U2314 (N_2314,In_337,In_851);
nand U2315 (N_2315,In_628,In_454);
and U2316 (N_2316,In_977,In_51);
nor U2317 (N_2317,In_565,In_36);
and U2318 (N_2318,In_235,In_893);
or U2319 (N_2319,In_179,In_866);
or U2320 (N_2320,In_300,In_91);
or U2321 (N_2321,In_450,In_568);
or U2322 (N_2322,In_166,In_80);
nor U2323 (N_2323,In_92,In_80);
nand U2324 (N_2324,In_140,In_911);
and U2325 (N_2325,In_777,In_14);
or U2326 (N_2326,In_214,In_696);
or U2327 (N_2327,In_342,In_768);
or U2328 (N_2328,In_994,In_901);
nor U2329 (N_2329,In_164,In_561);
or U2330 (N_2330,In_400,In_847);
nand U2331 (N_2331,In_325,In_123);
or U2332 (N_2332,In_944,In_146);
and U2333 (N_2333,In_311,In_924);
or U2334 (N_2334,In_623,In_777);
nand U2335 (N_2335,In_546,In_556);
nor U2336 (N_2336,In_218,In_377);
nand U2337 (N_2337,In_38,In_327);
or U2338 (N_2338,In_724,In_825);
nand U2339 (N_2339,In_588,In_695);
nor U2340 (N_2340,In_293,In_908);
and U2341 (N_2341,In_174,In_982);
nor U2342 (N_2342,In_404,In_688);
or U2343 (N_2343,In_386,In_879);
nor U2344 (N_2344,In_194,In_25);
nand U2345 (N_2345,In_416,In_167);
nand U2346 (N_2346,In_561,In_400);
and U2347 (N_2347,In_885,In_447);
or U2348 (N_2348,In_773,In_481);
xnor U2349 (N_2349,In_102,In_248);
xnor U2350 (N_2350,In_306,In_881);
nand U2351 (N_2351,In_38,In_677);
or U2352 (N_2352,In_932,In_989);
or U2353 (N_2353,In_142,In_270);
or U2354 (N_2354,In_339,In_287);
and U2355 (N_2355,In_105,In_994);
or U2356 (N_2356,In_569,In_297);
nand U2357 (N_2357,In_613,In_673);
and U2358 (N_2358,In_46,In_706);
or U2359 (N_2359,In_557,In_884);
nor U2360 (N_2360,In_518,In_385);
and U2361 (N_2361,In_322,In_630);
nor U2362 (N_2362,In_539,In_346);
nor U2363 (N_2363,In_961,In_181);
or U2364 (N_2364,In_949,In_645);
nand U2365 (N_2365,In_776,In_977);
nor U2366 (N_2366,In_331,In_607);
nor U2367 (N_2367,In_229,In_856);
or U2368 (N_2368,In_524,In_461);
nor U2369 (N_2369,In_477,In_523);
and U2370 (N_2370,In_346,In_61);
or U2371 (N_2371,In_425,In_907);
nor U2372 (N_2372,In_249,In_115);
xor U2373 (N_2373,In_499,In_701);
nor U2374 (N_2374,In_403,In_22);
nor U2375 (N_2375,In_216,In_548);
nand U2376 (N_2376,In_495,In_649);
nor U2377 (N_2377,In_365,In_692);
nand U2378 (N_2378,In_28,In_630);
or U2379 (N_2379,In_590,In_60);
nand U2380 (N_2380,In_635,In_988);
nand U2381 (N_2381,In_688,In_806);
and U2382 (N_2382,In_58,In_20);
and U2383 (N_2383,In_938,In_2);
and U2384 (N_2384,In_899,In_188);
nand U2385 (N_2385,In_48,In_774);
nor U2386 (N_2386,In_868,In_972);
nand U2387 (N_2387,In_784,In_238);
and U2388 (N_2388,In_6,In_90);
nand U2389 (N_2389,In_614,In_5);
nor U2390 (N_2390,In_774,In_857);
nor U2391 (N_2391,In_976,In_423);
or U2392 (N_2392,In_71,In_111);
and U2393 (N_2393,In_306,In_748);
nand U2394 (N_2394,In_850,In_303);
or U2395 (N_2395,In_720,In_335);
and U2396 (N_2396,In_107,In_474);
or U2397 (N_2397,In_215,In_571);
nor U2398 (N_2398,In_643,In_413);
or U2399 (N_2399,In_989,In_917);
nor U2400 (N_2400,In_165,In_122);
nand U2401 (N_2401,In_93,In_622);
nand U2402 (N_2402,In_705,In_644);
nor U2403 (N_2403,In_942,In_612);
and U2404 (N_2404,In_742,In_500);
or U2405 (N_2405,In_10,In_704);
nor U2406 (N_2406,In_958,In_379);
or U2407 (N_2407,In_38,In_918);
xor U2408 (N_2408,In_592,In_709);
nor U2409 (N_2409,In_969,In_710);
and U2410 (N_2410,In_640,In_337);
nor U2411 (N_2411,In_657,In_132);
and U2412 (N_2412,In_620,In_63);
or U2413 (N_2413,In_430,In_451);
and U2414 (N_2414,In_857,In_973);
or U2415 (N_2415,In_925,In_882);
nand U2416 (N_2416,In_715,In_258);
and U2417 (N_2417,In_505,In_328);
nor U2418 (N_2418,In_661,In_420);
or U2419 (N_2419,In_924,In_816);
nand U2420 (N_2420,In_628,In_675);
and U2421 (N_2421,In_180,In_917);
nor U2422 (N_2422,In_629,In_178);
and U2423 (N_2423,In_386,In_468);
and U2424 (N_2424,In_382,In_124);
nor U2425 (N_2425,In_105,In_282);
nand U2426 (N_2426,In_948,In_265);
nor U2427 (N_2427,In_811,In_37);
and U2428 (N_2428,In_19,In_623);
or U2429 (N_2429,In_750,In_573);
nor U2430 (N_2430,In_883,In_694);
or U2431 (N_2431,In_590,In_318);
and U2432 (N_2432,In_887,In_807);
and U2433 (N_2433,In_766,In_269);
and U2434 (N_2434,In_972,In_281);
nand U2435 (N_2435,In_725,In_560);
nand U2436 (N_2436,In_423,In_854);
and U2437 (N_2437,In_604,In_635);
nor U2438 (N_2438,In_82,In_317);
nor U2439 (N_2439,In_614,In_845);
and U2440 (N_2440,In_469,In_372);
or U2441 (N_2441,In_312,In_631);
nand U2442 (N_2442,In_549,In_629);
nor U2443 (N_2443,In_557,In_395);
nor U2444 (N_2444,In_546,In_660);
or U2445 (N_2445,In_945,In_635);
nand U2446 (N_2446,In_755,In_701);
and U2447 (N_2447,In_385,In_382);
or U2448 (N_2448,In_300,In_995);
and U2449 (N_2449,In_619,In_753);
or U2450 (N_2450,In_409,In_900);
or U2451 (N_2451,In_578,In_494);
or U2452 (N_2452,In_69,In_550);
and U2453 (N_2453,In_738,In_482);
nor U2454 (N_2454,In_938,In_193);
or U2455 (N_2455,In_255,In_845);
nand U2456 (N_2456,In_839,In_950);
nor U2457 (N_2457,In_989,In_438);
nand U2458 (N_2458,In_213,In_598);
nand U2459 (N_2459,In_520,In_837);
nand U2460 (N_2460,In_282,In_88);
nand U2461 (N_2461,In_717,In_506);
nor U2462 (N_2462,In_581,In_988);
nand U2463 (N_2463,In_67,In_531);
and U2464 (N_2464,In_417,In_769);
nand U2465 (N_2465,In_945,In_69);
and U2466 (N_2466,In_240,In_347);
nand U2467 (N_2467,In_74,In_969);
and U2468 (N_2468,In_888,In_116);
nand U2469 (N_2469,In_322,In_377);
or U2470 (N_2470,In_597,In_296);
and U2471 (N_2471,In_247,In_250);
and U2472 (N_2472,In_250,In_499);
and U2473 (N_2473,In_149,In_902);
and U2474 (N_2474,In_432,In_45);
and U2475 (N_2475,In_690,In_650);
nand U2476 (N_2476,In_974,In_722);
or U2477 (N_2477,In_810,In_518);
or U2478 (N_2478,In_140,In_459);
and U2479 (N_2479,In_998,In_841);
nor U2480 (N_2480,In_356,In_39);
nand U2481 (N_2481,In_429,In_728);
nand U2482 (N_2482,In_191,In_651);
or U2483 (N_2483,In_100,In_665);
nand U2484 (N_2484,In_188,In_25);
and U2485 (N_2485,In_351,In_57);
nor U2486 (N_2486,In_443,In_757);
or U2487 (N_2487,In_16,In_990);
and U2488 (N_2488,In_417,In_715);
nand U2489 (N_2489,In_768,In_521);
and U2490 (N_2490,In_529,In_557);
nand U2491 (N_2491,In_945,In_401);
and U2492 (N_2492,In_978,In_879);
or U2493 (N_2493,In_192,In_237);
nand U2494 (N_2494,In_80,In_472);
and U2495 (N_2495,In_201,In_151);
or U2496 (N_2496,In_149,In_523);
or U2497 (N_2497,In_597,In_537);
nand U2498 (N_2498,In_690,In_401);
and U2499 (N_2499,In_739,In_185);
and U2500 (N_2500,N_244,N_1142);
nor U2501 (N_2501,N_666,N_147);
nor U2502 (N_2502,N_1067,N_1671);
nand U2503 (N_2503,N_1410,N_1688);
nand U2504 (N_2504,N_980,N_2298);
nor U2505 (N_2505,N_2354,N_1642);
nor U2506 (N_2506,N_1480,N_1794);
or U2507 (N_2507,N_1973,N_10);
and U2508 (N_2508,N_2369,N_1710);
and U2509 (N_2509,N_146,N_2119);
nand U2510 (N_2510,N_261,N_1938);
nor U2511 (N_2511,N_644,N_1173);
nand U2512 (N_2512,N_1300,N_1704);
and U2513 (N_2513,N_1074,N_1780);
nor U2514 (N_2514,N_1620,N_1983);
or U2515 (N_2515,N_1931,N_1213);
and U2516 (N_2516,N_1148,N_583);
or U2517 (N_2517,N_654,N_1701);
nor U2518 (N_2518,N_458,N_2042);
nand U2519 (N_2519,N_1644,N_1250);
and U2520 (N_2520,N_167,N_1376);
or U2521 (N_2521,N_813,N_158);
and U2522 (N_2522,N_2426,N_1234);
or U2523 (N_2523,N_1838,N_214);
nand U2524 (N_2524,N_1334,N_700);
nor U2525 (N_2525,N_625,N_997);
nor U2526 (N_2526,N_889,N_199);
nand U2527 (N_2527,N_2289,N_1050);
nor U2528 (N_2528,N_2445,N_2222);
nand U2529 (N_2529,N_807,N_2013);
and U2530 (N_2530,N_2319,N_1637);
nor U2531 (N_2531,N_2323,N_400);
nor U2532 (N_2532,N_80,N_1869);
and U2533 (N_2533,N_1842,N_641);
nor U2534 (N_2534,N_1221,N_114);
and U2535 (N_2535,N_2364,N_760);
nor U2536 (N_2536,N_1757,N_2328);
and U2537 (N_2537,N_2460,N_2341);
nor U2538 (N_2538,N_1291,N_2370);
and U2539 (N_2539,N_1564,N_1925);
nor U2540 (N_2540,N_1723,N_172);
nor U2541 (N_2541,N_2416,N_2009);
or U2542 (N_2542,N_821,N_313);
or U2543 (N_2543,N_349,N_990);
or U2544 (N_2544,N_98,N_1242);
nand U2545 (N_2545,N_32,N_1206);
nand U2546 (N_2546,N_374,N_1280);
and U2547 (N_2547,N_1229,N_229);
nand U2548 (N_2548,N_470,N_2349);
or U2549 (N_2549,N_1285,N_717);
xor U2550 (N_2550,N_1429,N_1005);
nand U2551 (N_2551,N_1498,N_2188);
nor U2552 (N_2552,N_651,N_1354);
or U2553 (N_2553,N_88,N_2083);
nand U2554 (N_2554,N_2483,N_691);
nor U2555 (N_2555,N_44,N_1699);
nand U2556 (N_2556,N_2431,N_2037);
nand U2557 (N_2557,N_1478,N_1967);
or U2558 (N_2558,N_1651,N_1488);
xnor U2559 (N_2559,N_148,N_2297);
nor U2560 (N_2560,N_433,N_956);
nor U2561 (N_2561,N_58,N_733);
and U2562 (N_2562,N_1135,N_833);
nand U2563 (N_2563,N_436,N_2146);
and U2564 (N_2564,N_2060,N_588);
or U2565 (N_2565,N_1076,N_828);
nor U2566 (N_2566,N_1158,N_271);
nor U2567 (N_2567,N_2288,N_2311);
nor U2568 (N_2568,N_438,N_2064);
or U2569 (N_2569,N_1874,N_1260);
nor U2570 (N_2570,N_1835,N_1729);
and U2571 (N_2571,N_721,N_1871);
or U2572 (N_2572,N_239,N_1433);
nand U2573 (N_2573,N_942,N_1787);
nor U2574 (N_2574,N_2330,N_316);
nor U2575 (N_2575,N_1316,N_1408);
nand U2576 (N_2576,N_1361,N_521);
nor U2577 (N_2577,N_1774,N_97);
and U2578 (N_2578,N_1094,N_623);
nor U2579 (N_2579,N_617,N_318);
and U2580 (N_2580,N_1960,N_2317);
nand U2581 (N_2581,N_480,N_2129);
or U2582 (N_2582,N_1303,N_1176);
or U2583 (N_2583,N_1430,N_96);
nand U2584 (N_2584,N_2286,N_2007);
nand U2585 (N_2585,N_993,N_2342);
nand U2586 (N_2586,N_1544,N_16);
nand U2587 (N_2587,N_402,N_2466);
and U2588 (N_2588,N_327,N_151);
nand U2589 (N_2589,N_501,N_379);
or U2590 (N_2590,N_1330,N_2137);
and U2591 (N_2591,N_1855,N_1385);
nand U2592 (N_2592,N_2246,N_134);
and U2593 (N_2593,N_742,N_1395);
and U2594 (N_2594,N_2391,N_2467);
and U2595 (N_2595,N_1128,N_2320);
or U2596 (N_2596,N_1188,N_1006);
and U2597 (N_2597,N_1437,N_636);
and U2598 (N_2598,N_1026,N_1039);
and U2599 (N_2599,N_876,N_26);
nand U2600 (N_2600,N_863,N_1347);
or U2601 (N_2601,N_163,N_2266);
and U2602 (N_2602,N_1661,N_1321);
and U2603 (N_2603,N_2475,N_99);
nor U2604 (N_2604,N_2403,N_1272);
or U2605 (N_2605,N_325,N_355);
or U2606 (N_2606,N_2187,N_631);
nor U2607 (N_2607,N_1692,N_1216);
and U2608 (N_2608,N_2443,N_484);
nor U2609 (N_2609,N_1129,N_1824);
or U2610 (N_2610,N_973,N_1293);
nand U2611 (N_2611,N_818,N_1634);
nor U2612 (N_2612,N_1359,N_345);
nor U2613 (N_2613,N_2059,N_1177);
nor U2614 (N_2614,N_684,N_1986);
xnor U2615 (N_2615,N_1784,N_2294);
nor U2616 (N_2616,N_2281,N_1271);
and U2617 (N_2617,N_2014,N_1868);
nor U2618 (N_2618,N_1734,N_444);
or U2619 (N_2619,N_1058,N_587);
or U2620 (N_2620,N_423,N_1220);
and U2621 (N_2621,N_523,N_429);
or U2622 (N_2622,N_1218,N_1970);
and U2623 (N_2623,N_220,N_2499);
and U2624 (N_2624,N_991,N_2025);
xor U2625 (N_2625,N_1889,N_552);
nor U2626 (N_2626,N_560,N_2149);
nand U2627 (N_2627,N_2293,N_912);
or U2628 (N_2628,N_2240,N_1989);
nor U2629 (N_2629,N_1759,N_1618);
nor U2630 (N_2630,N_1298,N_2295);
nand U2631 (N_2631,N_2350,N_1265);
and U2632 (N_2632,N_1543,N_779);
and U2633 (N_2633,N_1880,N_15);
nor U2634 (N_2634,N_756,N_49);
nand U2635 (N_2635,N_1594,N_2331);
nor U2636 (N_2636,N_1565,N_213);
or U2637 (N_2637,N_279,N_1217);
or U2638 (N_2638,N_683,N_1553);
nand U2639 (N_2639,N_2248,N_1537);
and U2640 (N_2640,N_1524,N_500);
nand U2641 (N_2641,N_1600,N_795);
nor U2642 (N_2642,N_573,N_887);
and U2643 (N_2643,N_1647,N_2136);
nor U2644 (N_2644,N_2357,N_1288);
nand U2645 (N_2645,N_2262,N_2408);
and U2646 (N_2646,N_1903,N_2169);
and U2647 (N_2647,N_1223,N_1004);
and U2648 (N_2648,N_2175,N_600);
nand U2649 (N_2649,N_2128,N_1735);
nand U2650 (N_2650,N_1578,N_1980);
and U2651 (N_2651,N_1664,N_2429);
nand U2652 (N_2652,N_1130,N_826);
or U2653 (N_2653,N_2232,N_531);
nor U2654 (N_2654,N_720,N_1782);
nand U2655 (N_2655,N_19,N_357);
and U2656 (N_2656,N_710,N_2425);
and U2657 (N_2657,N_1160,N_320);
or U2658 (N_2658,N_2110,N_1152);
nor U2659 (N_2659,N_2315,N_1904);
nor U2660 (N_2660,N_1629,N_321);
or U2661 (N_2661,N_926,N_2300);
and U2662 (N_2662,N_515,N_2045);
or U2663 (N_2663,N_1415,N_1314);
or U2664 (N_2664,N_2305,N_2296);
or U2665 (N_2665,N_2327,N_1523);
nand U2666 (N_2666,N_1231,N_743);
nand U2667 (N_2667,N_1048,N_1845);
or U2668 (N_2668,N_95,N_2356);
or U2669 (N_2669,N_1161,N_2435);
and U2670 (N_2670,N_1682,N_2145);
nor U2671 (N_2671,N_106,N_2267);
and U2672 (N_2672,N_2276,N_1091);
or U2673 (N_2673,N_609,N_1950);
or U2674 (N_2674,N_4,N_1261);
or U2675 (N_2675,N_897,N_2155);
nand U2676 (N_2676,N_2264,N_690);
nand U2677 (N_2677,N_1089,N_1088);
or U2678 (N_2678,N_109,N_1133);
nand U2679 (N_2679,N_1412,N_285);
and U2680 (N_2680,N_100,N_2474);
or U2681 (N_2681,N_249,N_2338);
nand U2682 (N_2682,N_1294,N_2143);
nor U2683 (N_2683,N_935,N_2035);
xnor U2684 (N_2684,N_270,N_326);
nor U2685 (N_2685,N_1849,N_749);
nor U2686 (N_2686,N_1696,N_1055);
nor U2687 (N_2687,N_1910,N_1905);
nand U2688 (N_2688,N_79,N_800);
nand U2689 (N_2689,N_1317,N_1561);
or U2690 (N_2690,N_2157,N_1653);
nor U2691 (N_2691,N_464,N_102);
or U2692 (N_2692,N_554,N_2046);
and U2693 (N_2693,N_525,N_1222);
or U2694 (N_2694,N_2406,N_2131);
and U2695 (N_2695,N_1147,N_1918);
and U2696 (N_2696,N_442,N_362);
nand U2697 (N_2697,N_1105,N_2352);
nor U2698 (N_2698,N_919,N_472);
or U2699 (N_2699,N_203,N_723);
or U2700 (N_2700,N_759,N_984);
nor U2701 (N_2701,N_2167,N_370);
or U2702 (N_2702,N_1820,N_2388);
and U2703 (N_2703,N_70,N_1636);
or U2704 (N_2704,N_881,N_2049);
nand U2705 (N_2705,N_1964,N_473);
nand U2706 (N_2706,N_844,N_810);
nor U2707 (N_2707,N_2290,N_1859);
nand U2708 (N_2708,N_1597,N_200);
or U2709 (N_2709,N_698,N_2337);
nor U2710 (N_2710,N_1659,N_1801);
nand U2711 (N_2711,N_1396,N_1358);
or U2712 (N_2712,N_596,N_2029);
nand U2713 (N_2713,N_788,N_1718);
and U2714 (N_2714,N_1079,N_384);
or U2715 (N_2715,N_622,N_86);
nand U2716 (N_2716,N_1436,N_864);
and U2717 (N_2717,N_1401,N_1350);
nand U2718 (N_2718,N_1806,N_1063);
and U2719 (N_2719,N_555,N_2132);
nor U2720 (N_2720,N_1694,N_794);
and U2721 (N_2721,N_1848,N_767);
nand U2722 (N_2722,N_1592,N_1827);
and U2723 (N_2723,N_1149,N_453);
and U2724 (N_2724,N_2056,N_708);
or U2725 (N_2725,N_2068,N_1154);
or U2726 (N_2726,N_862,N_2359);
or U2727 (N_2727,N_1752,N_116);
nand U2728 (N_2728,N_1164,N_2306);
or U2729 (N_2729,N_787,N_849);
nand U2730 (N_2730,N_286,N_761);
or U2731 (N_2731,N_1695,N_1425);
and U2732 (N_2732,N_837,N_404);
and U2733 (N_2733,N_724,N_675);
or U2734 (N_2734,N_1573,N_288);
nor U2735 (N_2735,N_455,N_1822);
nand U2736 (N_2736,N_1252,N_1962);
nor U2737 (N_2737,N_1484,N_1096);
or U2738 (N_2738,N_1598,N_1035);
nor U2739 (N_2739,N_1958,N_2393);
nand U2740 (N_2740,N_605,N_242);
and U2741 (N_2741,N_1036,N_1018);
nor U2742 (N_2742,N_2008,N_45);
nor U2743 (N_2743,N_69,N_972);
nor U2744 (N_2744,N_226,N_1021);
and U2745 (N_2745,N_1595,N_445);
or U2746 (N_2746,N_1509,N_1447);
or U2747 (N_2747,N_2252,N_888);
or U2748 (N_2748,N_373,N_1828);
and U2749 (N_2749,N_882,N_2072);
or U2750 (N_2750,N_1900,N_2186);
nand U2751 (N_2751,N_34,N_1405);
and U2752 (N_2752,N_1716,N_171);
and U2753 (N_2753,N_1325,N_629);
and U2754 (N_2754,N_1483,N_2441);
nor U2755 (N_2755,N_447,N_2150);
nand U2756 (N_2756,N_2057,N_2253);
and U2757 (N_2757,N_1807,N_806);
or U2758 (N_2758,N_2032,N_76);
nand U2759 (N_2759,N_1529,N_1273);
or U2760 (N_2760,N_1712,N_1001);
nand U2761 (N_2761,N_1468,N_390);
or U2762 (N_2762,N_1506,N_1626);
nor U2763 (N_2763,N_730,N_2115);
nor U2764 (N_2764,N_1451,N_75);
or U2765 (N_2765,N_1539,N_1377);
nor U2766 (N_2766,N_1715,N_187);
xnor U2767 (N_2767,N_2422,N_1496);
nor U2768 (N_2768,N_677,N_931);
and U2769 (N_2769,N_1745,N_274);
nor U2770 (N_2770,N_2133,N_928);
nor U2771 (N_2771,N_1031,N_1282);
and U2772 (N_2772,N_948,N_1374);
nand U2773 (N_2773,N_1215,N_658);
and U2774 (N_2774,N_1525,N_1403);
and U2775 (N_2775,N_777,N_1940);
nand U2776 (N_2776,N_2274,N_1398);
and U2777 (N_2777,N_1665,N_1179);
and U2778 (N_2778,N_1894,N_299);
nor U2779 (N_2779,N_856,N_101);
and U2780 (N_2780,N_1858,N_1440);
nor U2781 (N_2781,N_1053,N_178);
and U2782 (N_2782,N_2480,N_1028);
nor U2783 (N_2783,N_1623,N_1362);
nand U2784 (N_2784,N_389,N_2263);
and U2785 (N_2785,N_1107,N_2421);
and U2786 (N_2786,N_1514,N_1235);
or U2787 (N_2787,N_2279,N_2148);
nor U2788 (N_2788,N_1382,N_2023);
nand U2789 (N_2789,N_1934,N_1134);
nand U2790 (N_2790,N_1344,N_1587);
and U2791 (N_2791,N_1011,N_2490);
and U2792 (N_2792,N_2401,N_869);
and U2793 (N_2793,N_1556,N_1302);
and U2794 (N_2794,N_1205,N_2449);
or U2795 (N_2795,N_2050,N_342);
nand U2796 (N_2796,N_1741,N_2268);
nor U2797 (N_2797,N_1500,N_1551);
or U2798 (N_2798,N_2107,N_2478);
and U2799 (N_2799,N_1789,N_660);
nand U2800 (N_2800,N_2385,N_1475);
nand U2801 (N_2801,N_115,N_1755);
nand U2802 (N_2802,N_944,N_1615);
and U2803 (N_2803,N_386,N_584);
nand U2804 (N_2804,N_55,N_2250);
nand U2805 (N_2805,N_1356,N_1126);
xor U2806 (N_2806,N_1109,N_1424);
or U2807 (N_2807,N_2247,N_2255);
or U2808 (N_2808,N_1375,N_574);
and U2809 (N_2809,N_1571,N_1240);
nand U2810 (N_2810,N_1608,N_2473);
nor U2811 (N_2811,N_385,N_1228);
nor U2812 (N_2812,N_1337,N_238);
nand U2813 (N_2813,N_865,N_1178);
nor U2814 (N_2814,N_145,N_1137);
and U2815 (N_2815,N_434,N_780);
or U2816 (N_2816,N_283,N_2417);
nor U2817 (N_2817,N_1071,N_2114);
and U2818 (N_2818,N_2447,N_808);
nand U2819 (N_2819,N_111,N_469);
and U2820 (N_2820,N_1531,N_1559);
or U2821 (N_2821,N_466,N_1990);
nand U2822 (N_2822,N_2402,N_2204);
or U2823 (N_2823,N_2237,N_517);
and U2824 (N_2824,N_785,N_1702);
nor U2825 (N_2825,N_563,N_2171);
or U2826 (N_2826,N_485,N_2095);
and U2827 (N_2827,N_1837,N_567);
nand U2828 (N_2828,N_1323,N_893);
nor U2829 (N_2829,N_565,N_890);
nand U2830 (N_2830,N_996,N_1454);
or U2831 (N_2831,N_1917,N_872);
and U2832 (N_2832,N_1909,N_918);
nor U2833 (N_2833,N_399,N_1856);
and U2834 (N_2834,N_2205,N_1125);
and U2835 (N_2835,N_1369,N_2384);
nand U2836 (N_2836,N_2244,N_2440);
and U2837 (N_2837,N_1533,N_1567);
nand U2838 (N_2838,N_62,N_278);
nand U2839 (N_2839,N_257,N_248);
nand U2840 (N_2840,N_830,N_2081);
nor U2841 (N_2841,N_1679,N_923);
or U2842 (N_2842,N_1033,N_2005);
and U2843 (N_2843,N_1777,N_222);
or U2844 (N_2844,N_728,N_191);
nand U2845 (N_2845,N_1054,N_713);
and U2846 (N_2846,N_2021,N_1459);
and U2847 (N_2847,N_394,N_1965);
nor U2848 (N_2848,N_435,N_443);
or U2849 (N_2849,N_614,N_1144);
nand U2850 (N_2850,N_1681,N_152);
and U2851 (N_2851,N_1996,N_2127);
and U2852 (N_2852,N_1799,N_144);
or U2853 (N_2853,N_1274,N_611);
or U2854 (N_2854,N_689,N_1439);
nand U2855 (N_2855,N_1087,N_981);
or U2856 (N_2856,N_1913,N_359);
and U2857 (N_2857,N_843,N_1230);
or U2858 (N_2858,N_2074,N_263);
nor U2859 (N_2859,N_1810,N_1490);
and U2860 (N_2860,N_2452,N_1009);
nand U2861 (N_2861,N_2418,N_2217);
and U2862 (N_2862,N_2363,N_514);
and U2863 (N_2863,N_121,N_858);
or U2864 (N_2864,N_906,N_2271);
nor U2865 (N_2865,N_256,N_1227);
nand U2866 (N_2866,N_946,N_1530);
nor U2867 (N_2867,N_934,N_1499);
and U2868 (N_2868,N_857,N_140);
nor U2869 (N_2869,N_2041,N_254);
or U2870 (N_2870,N_1301,N_1654);
and U2871 (N_2871,N_352,N_1332);
nor U2872 (N_2872,N_2113,N_1435);
and U2873 (N_2873,N_620,N_2075);
nand U2874 (N_2874,N_1093,N_2302);
and U2875 (N_2875,N_1819,N_608);
or U2876 (N_2876,N_2026,N_712);
or U2877 (N_2877,N_1897,N_2151);
nor U2878 (N_2878,N_1120,N_1491);
or U2879 (N_2879,N_678,N_1550);
and U2880 (N_2880,N_543,N_1645);
nor U2881 (N_2881,N_1946,N_1628);
or U2882 (N_2882,N_426,N_347);
and U2883 (N_2883,N_1972,N_259);
nor U2884 (N_2884,N_2206,N_2170);
and U2885 (N_2885,N_796,N_2096);
and U2886 (N_2886,N_1110,N_2079);
or U2887 (N_2887,N_2344,N_1180);
nor U2888 (N_2888,N_2482,N_1977);
nand U2889 (N_2889,N_282,N_1527);
nor U2890 (N_2890,N_1951,N_153);
or U2891 (N_2891,N_1102,N_561);
and U2892 (N_2892,N_334,N_1870);
and U2893 (N_2893,N_1373,N_477);
nand U2894 (N_2894,N_1731,N_2138);
nor U2895 (N_2895,N_1511,N_1726);
and U2896 (N_2896,N_456,N_894);
nand U2897 (N_2897,N_2099,N_489);
and U2898 (N_2898,N_1943,N_1577);
nand U2899 (N_2899,N_1995,N_917);
or U2900 (N_2900,N_1453,N_361);
nand U2901 (N_2901,N_2378,N_1119);
or U2902 (N_2902,N_2278,N_2396);
or U2903 (N_2903,N_1208,N_706);
or U2904 (N_2904,N_1025,N_1997);
or U2905 (N_2905,N_1601,N_524);
and U2906 (N_2906,N_1365,N_372);
nor U2907 (N_2907,N_1762,N_245);
nor U2908 (N_2908,N_2351,N_2454);
nand U2909 (N_2909,N_982,N_964);
and U2910 (N_2910,N_1669,N_1812);
nor U2911 (N_2911,N_1413,N_309);
or U2912 (N_2912,N_2367,N_891);
nand U2913 (N_2913,N_2314,N_1896);
nor U2914 (N_2914,N_1319,N_971);
and U2915 (N_2915,N_48,N_1717);
or U2916 (N_2916,N_1010,N_548);
nand U2917 (N_2917,N_91,N_1570);
or U2918 (N_2918,N_838,N_1211);
nor U2919 (N_2919,N_1985,N_495);
nor U2920 (N_2920,N_781,N_1020);
nand U2921 (N_2921,N_417,N_527);
xor U2922 (N_2922,N_750,N_542);
xor U2923 (N_2923,N_1497,N_23);
nand U2924 (N_2924,N_36,N_989);
or U2925 (N_2925,N_1778,N_1426);
nand U2926 (N_2926,N_1086,N_5);
and U2927 (N_2927,N_2208,N_1748);
nor U2928 (N_2928,N_992,N_746);
and U2929 (N_2929,N_896,N_606);
or U2930 (N_2930,N_1493,N_507);
or U2931 (N_2931,N_262,N_2090);
and U2932 (N_2932,N_705,N_1814);
and U2933 (N_2933,N_1185,N_1522);
nand U2934 (N_2934,N_1516,N_1742);
nor U2935 (N_2935,N_1893,N_1753);
nand U2936 (N_2936,N_2193,N_142);
or U2937 (N_2937,N_2180,N_2471);
or U2938 (N_2938,N_680,N_1312);
nor U2939 (N_2939,N_2409,N_860);
nand U2940 (N_2940,N_873,N_255);
or U2941 (N_2941,N_1649,N_1928);
nand U2942 (N_2942,N_770,N_2434);
xnor U2943 (N_2943,N_156,N_1568);
or U2944 (N_2944,N_1790,N_1061);
nand U2945 (N_2945,N_1434,N_1472);
nor U2946 (N_2946,N_2310,N_1226);
nor U2947 (N_2947,N_2335,N_2088);
nor U2948 (N_2948,N_1077,N_2481);
and U2949 (N_2949,N_532,N_1898);
and U2950 (N_2950,N_1428,N_2343);
nor U2951 (N_2951,N_1821,N_353);
and U2952 (N_2952,N_1486,N_490);
nor U2953 (N_2953,N_1341,N_1090);
nor U2954 (N_2954,N_1467,N_886);
nor U2955 (N_2955,N_2018,N_1037);
nand U2956 (N_2956,N_162,N_2368);
nor U2957 (N_2957,N_269,N_1507);
or U2958 (N_2958,N_1246,N_2275);
nand U2959 (N_2959,N_635,N_1324);
nor U2960 (N_2960,N_1582,N_594);
or U2961 (N_2961,N_1342,N_1363);
nor U2962 (N_2962,N_804,N_241);
nor U2963 (N_2963,N_637,N_303);
nand U2964 (N_2964,N_314,N_820);
or U2965 (N_2965,N_251,N_2174);
nor U2966 (N_2966,N_441,N_2185);
and U2967 (N_2967,N_2439,N_2413);
or U2968 (N_2968,N_578,N_1232);
or U2969 (N_2969,N_1966,N_722);
or U2970 (N_2970,N_1936,N_401);
nand U2971 (N_2971,N_415,N_2106);
nor U2972 (N_2972,N_29,N_1825);
nand U2973 (N_2973,N_2055,N_2325);
nor U2974 (N_2974,N_2197,N_411);
nor U2975 (N_2975,N_2303,N_1040);
or U2976 (N_2976,N_762,N_1992);
and U2977 (N_2977,N_440,N_166);
nor U2978 (N_2978,N_468,N_396);
and U2979 (N_2979,N_487,N_1318);
or U2980 (N_2980,N_28,N_1933);
or U2981 (N_2981,N_1993,N_701);
nor U2982 (N_2982,N_2027,N_2153);
xnor U2983 (N_2983,N_2446,N_1007);
nand U2984 (N_2984,N_2433,N_1915);
and U2985 (N_2985,N_12,N_1542);
and U2986 (N_2986,N_758,N_481);
and U2987 (N_2987,N_1032,N_929);
nor U2988 (N_2988,N_180,N_598);
or U2989 (N_2989,N_930,N_2010);
or U2990 (N_2990,N_2047,N_413);
and U2991 (N_2991,N_1655,N_2051);
nor U2992 (N_2992,N_575,N_694);
nor U2993 (N_2993,N_1823,N_1326);
or U2994 (N_2994,N_1482,N_789);
nor U2995 (N_2995,N_518,N_1195);
and U2996 (N_2996,N_296,N_1008);
or U2997 (N_2997,N_300,N_510);
xor U2998 (N_2998,N_378,N_911);
or U2999 (N_2999,N_38,N_768);
nor U3000 (N_3000,N_845,N_2191);
nand U3001 (N_3001,N_1059,N_1954);
or U3002 (N_3002,N_2100,N_949);
nor U3003 (N_3003,N_1257,N_1526);
nor U3004 (N_3004,N_1612,N_1355);
nand U3005 (N_3005,N_1225,N_1908);
and U3006 (N_3006,N_735,N_71);
nor U3007 (N_3007,N_317,N_2484);
nor U3008 (N_3008,N_1576,N_363);
or U3009 (N_3009,N_848,N_1092);
or U3010 (N_3010,N_1698,N_1172);
and U3011 (N_3011,N_1877,N_2233);
nor U3012 (N_3012,N_711,N_1987);
and U3013 (N_3013,N_1023,N_586);
nand U3014 (N_3014,N_2124,N_963);
or U3015 (N_3015,N_1719,N_2380);
and U3016 (N_3016,N_1157,N_1586);
nor U3017 (N_3017,N_987,N_1448);
xor U3018 (N_3018,N_1192,N_1268);
and U3019 (N_3019,N_2016,N_1183);
nand U3020 (N_3020,N_1998,N_59);
nor U3021 (N_3021,N_737,N_1277);
or U3022 (N_3022,N_1236,N_1163);
and U3023 (N_3023,N_1101,N_580);
or U3024 (N_3024,N_859,N_2097);
or U3025 (N_3025,N_1443,N_2238);
or U3026 (N_3026,N_757,N_853);
nor U3027 (N_3027,N_1540,N_2235);
nand U3028 (N_3028,N_615,N_2257);
and U3029 (N_3029,N_1818,N_265);
and U3030 (N_3030,N_1667,N_452);
nor U3031 (N_3031,N_842,N_2236);
or U3032 (N_3032,N_1627,N_1836);
nor U3033 (N_3033,N_1839,N_335);
nor U3034 (N_3034,N_1560,N_2472);
nor U3035 (N_3035,N_1136,N_1060);
or U3036 (N_3036,N_966,N_939);
nor U3037 (N_3037,N_538,N_1418);
nand U3038 (N_3038,N_427,N_2147);
and U3039 (N_3039,N_792,N_2242);
and U3040 (N_3040,N_1924,N_688);
nand U3041 (N_3041,N_1674,N_2160);
nand U3042 (N_3042,N_2491,N_1492);
nand U3043 (N_3043,N_1432,N_405);
and U3044 (N_3044,N_2166,N_2375);
and U3045 (N_3045,N_2182,N_1269);
and U3046 (N_3046,N_2420,N_1833);
nand U3047 (N_3047,N_1150,N_1760);
and U3048 (N_3048,N_1469,N_1563);
nor U3049 (N_3049,N_2033,N_1788);
nand U3050 (N_3050,N_1515,N_1815);
nor U3051 (N_3051,N_183,N_324);
or U3052 (N_3052,N_909,N_607);
nor U3053 (N_3053,N_1663,N_476);
or U3054 (N_3054,N_1714,N_1263);
or U3055 (N_3055,N_940,N_2273);
nand U3056 (N_3056,N_383,N_281);
nand U3057 (N_3057,N_1746,N_1322);
nand U3058 (N_3058,N_37,N_976);
and U3059 (N_3059,N_297,N_1999);
or U3060 (N_3060,N_1168,N_0);
nand U3061 (N_3061,N_2102,N_1387);
and U3062 (N_3062,N_1166,N_1327);
nand U3063 (N_3063,N_280,N_40);
nor U3064 (N_3064,N_582,N_2152);
nor U3065 (N_3065,N_1034,N_1638);
or U3066 (N_3066,N_901,N_670);
nor U3067 (N_3067,N_1536,N_1445);
or U3068 (N_3068,N_2230,N_137);
and U3069 (N_3069,N_2105,N_253);
nor U3070 (N_3070,N_1895,N_686);
or U3071 (N_3071,N_1854,N_1400);
nand U3072 (N_3072,N_572,N_2123);
nor U3073 (N_3073,N_2339,N_1886);
nand U3074 (N_3074,N_1155,N_977);
nor U3075 (N_3075,N_2428,N_633);
nor U3076 (N_3076,N_1141,N_503);
and U3077 (N_3077,N_290,N_343);
nand U3078 (N_3078,N_1057,N_593);
and U3079 (N_3079,N_1182,N_1923);
nor U3080 (N_3080,N_9,N_1552);
nor U3081 (N_3081,N_1545,N_168);
nor U3082 (N_3082,N_576,N_805);
nor U3083 (N_3083,N_1393,N_1975);
and U3084 (N_3084,N_1963,N_437);
and U3085 (N_3085,N_1541,N_1419);
nor U3086 (N_3086,N_1941,N_425);
or U3087 (N_3087,N_1899,N_1463);
nand U3088 (N_3088,N_454,N_884);
nand U3089 (N_3089,N_2073,N_551);
nand U3090 (N_3090,N_112,N_663);
or U3091 (N_3091,N_138,N_2098);
nand U3092 (N_3092,N_1705,N_1124);
or U3093 (N_3093,N_1795,N_2358);
nor U3094 (N_3094,N_105,N_161);
and U3095 (N_3095,N_451,N_2168);
or U3096 (N_3096,N_1214,N_589);
nor U3097 (N_3097,N_159,N_1611);
nor U3098 (N_3098,N_2398,N_1779);
or U3099 (N_3099,N_2414,N_772);
and U3100 (N_3100,N_937,N_1184);
nand U3101 (N_3101,N_165,N_1722);
or U3102 (N_3102,N_2340,N_1733);
and U3103 (N_3103,N_613,N_1115);
and U3104 (N_3104,N_1557,N_1861);
or U3105 (N_3105,N_1357,N_155);
or U3106 (N_3106,N_653,N_907);
nand U3107 (N_3107,N_1813,N_1707);
nand U3108 (N_3108,N_504,N_85);
or U3109 (N_3109,N_1680,N_1198);
or U3110 (N_3110,N_356,N_1850);
xnor U3111 (N_3111,N_1012,N_1749);
or U3112 (N_3112,N_260,N_1811);
nor U3113 (N_3113,N_764,N_2468);
and U3114 (N_3114,N_1015,N_1421);
nor U3115 (N_3115,N_1736,N_185);
and U3116 (N_3116,N_467,N_2334);
nor U3117 (N_3117,N_366,N_1508);
nor U3118 (N_3118,N_17,N_1069);
nor U3119 (N_3119,N_2223,N_1817);
or U3120 (N_3120,N_817,N_53);
nor U3121 (N_3121,N_408,N_2112);
or U3122 (N_3122,N_2430,N_73);
nor U3123 (N_3123,N_988,N_1391);
or U3124 (N_3124,N_2094,N_1340);
nor U3125 (N_3125,N_2091,N_656);
or U3126 (N_3126,N_983,N_1932);
nor U3127 (N_3127,N_1386,N_39);
nor U3128 (N_3128,N_2400,N_1098);
nor U3129 (N_3129,N_2386,N_292);
and U3130 (N_3130,N_83,N_516);
and U3131 (N_3131,N_209,N_2231);
or U3132 (N_3132,N_1689,N_92);
nand U3133 (N_3133,N_2292,N_1911);
nor U3134 (N_3134,N_1381,N_773);
nand U3135 (N_3135,N_782,N_266);
or U3136 (N_3136,N_212,N_1417);
or U3137 (N_3137,N_2432,N_2063);
and U3138 (N_3138,N_1593,N_1153);
nand U3139 (N_3139,N_1279,N_695);
nand U3140 (N_3140,N_1535,N_1367);
or U3141 (N_3141,N_1307,N_1464);
and U3142 (N_3142,N_246,N_422);
or U3143 (N_3143,N_2371,N_2054);
or U3144 (N_3144,N_537,N_585);
and U3145 (N_3145,N_306,N_741);
nor U3146 (N_3146,N_420,N_2141);
nand U3147 (N_3147,N_1081,N_682);
nand U3148 (N_3148,N_2347,N_130);
or U3149 (N_3149,N_752,N_1914);
and U3150 (N_3150,N_522,N_344);
and U3151 (N_3151,N_903,N_1580);
nand U3152 (N_3152,N_2280,N_1056);
and U3153 (N_3153,N_432,N_358);
and U3154 (N_3154,N_1579,N_2002);
and U3155 (N_3155,N_228,N_225);
nand U3156 (N_3156,N_298,N_638);
or U3157 (N_3157,N_1264,N_947);
nand U3158 (N_3158,N_179,N_751);
nand U3159 (N_3159,N_2165,N_90);
nand U3160 (N_3160,N_969,N_645);
and U3161 (N_3161,N_1520,N_305);
nand U3162 (N_3162,N_1331,N_42);
or U3163 (N_3163,N_1052,N_509);
nand U3164 (N_3164,N_1585,N_914);
nand U3165 (N_3165,N_380,N_1668);
or U3166 (N_3166,N_1423,N_267);
nand U3167 (N_3167,N_136,N_2058);
and U3168 (N_3168,N_1534,N_2203);
or U3169 (N_3169,N_646,N_719);
and U3170 (N_3170,N_545,N_2179);
nand U3171 (N_3171,N_135,N_2229);
and U3172 (N_3172,N_395,N_1030);
nor U3173 (N_3173,N_954,N_1721);
nand U3174 (N_3174,N_2399,N_703);
or U3175 (N_3175,N_661,N_368);
nor U3176 (N_3176,N_1479,N_1662);
and U3177 (N_3177,N_128,N_1043);
nor U3178 (N_3178,N_1832,N_1919);
nor U3179 (N_3179,N_1384,N_1796);
xor U3180 (N_3180,N_1194,N_1657);
and U3181 (N_3181,N_1792,N_1175);
nor U3182 (N_3182,N_175,N_104);
or U3183 (N_3183,N_2156,N_1766);
nand U3184 (N_3184,N_925,N_775);
nand U3185 (N_3185,N_3,N_1872);
and U3186 (N_3186,N_1083,N_2486);
nand U3187 (N_3187,N_197,N_1343);
or U3188 (N_3188,N_2234,N_1633);
nand U3189 (N_3189,N_1554,N_346);
nand U3190 (N_3190,N_331,N_2423);
or U3191 (N_3191,N_2022,N_718);
or U3192 (N_3192,N_1860,N_194);
and U3193 (N_3193,N_177,N_1968);
or U3194 (N_3194,N_508,N_129);
nor U3195 (N_3195,N_1471,N_340);
or U3196 (N_3196,N_1084,N_2366);
nand U3197 (N_3197,N_2382,N_193);
nand U3198 (N_3198,N_2043,N_618);
nand U3199 (N_3199,N_94,N_642);
or U3200 (N_3200,N_943,N_1513);
and U3201 (N_3201,N_1394,N_1569);
and U3202 (N_3202,N_736,N_1191);
and U3203 (N_3203,N_916,N_1407);
and U3204 (N_3204,N_93,N_1785);
or U3205 (N_3205,N_459,N_1399);
and U3206 (N_3206,N_189,N_132);
or U3207 (N_3207,N_1197,N_2078);
and U3208 (N_3208,N_921,N_2077);
xnor U3209 (N_3209,N_716,N_2154);
nand U3210 (N_3210,N_412,N_2318);
or U3211 (N_3211,N_1641,N_1504);
nor U3212 (N_3212,N_1202,N_558);
nor U3213 (N_3213,N_382,N_562);
and U3214 (N_3214,N_1632,N_13);
xor U3215 (N_3215,N_2158,N_293);
and U3216 (N_3216,N_230,N_416);
xnor U3217 (N_3217,N_900,N_702);
or U3218 (N_3218,N_765,N_41);
and U3219 (N_3219,N_2039,N_46);
or U3220 (N_3220,N_1487,N_2020);
or U3221 (N_3221,N_421,N_1402);
nand U3222 (N_3222,N_559,N_2412);
and U3223 (N_3223,N_1863,N_2116);
or U3224 (N_3224,N_364,N_235);
and U3225 (N_3225,N_494,N_1121);
or U3226 (N_3226,N_1921,N_2254);
nand U3227 (N_3227,N_1851,N_878);
nor U3228 (N_3228,N_1174,N_1131);
nor U3229 (N_3229,N_2092,N_850);
and U3230 (N_3230,N_1427,N_1614);
nor U3231 (N_3231,N_1306,N_1099);
nor U3232 (N_3232,N_2256,N_709);
or U3233 (N_3233,N_323,N_840);
and U3234 (N_3234,N_2415,N_2065);
nor U3235 (N_3235,N_1047,N_1768);
or U3236 (N_3236,N_1605,N_1609);
nor U3237 (N_3237,N_2450,N_2361);
and U3238 (N_3238,N_513,N_938);
nor U3239 (N_3239,N_1847,N_206);
and U3240 (N_3240,N_2488,N_1866);
nor U3241 (N_3241,N_1684,N_164);
nand U3242 (N_3242,N_955,N_502);
nor U3243 (N_3243,N_1151,N_289);
or U3244 (N_3244,N_2457,N_2397);
or U3245 (N_3245,N_143,N_192);
and U3246 (N_3246,N_2161,N_124);
nand U3247 (N_3247,N_1349,N_2269);
and U3248 (N_3248,N_2453,N_814);
nor U3249 (N_3249,N_650,N_1621);
or U3250 (N_3250,N_2285,N_1957);
and U3251 (N_3251,N_1650,N_1404);
and U3252 (N_3252,N_2071,N_1117);
nor U3253 (N_3253,N_1624,N_1431);
or U3254 (N_3254,N_2392,N_2086);
and U3255 (N_3255,N_2213,N_1831);
nand U3256 (N_3256,N_2178,N_1687);
and U3257 (N_3257,N_196,N_904);
and U3258 (N_3258,N_2066,N_1920);
and U3259 (N_3259,N_968,N_1466);
nand U3260 (N_3260,N_273,N_846);
nand U3261 (N_3261,N_439,N_122);
or U3262 (N_3262,N_1283,N_920);
and U3263 (N_3263,N_117,N_67);
or U3264 (N_3264,N_498,N_839);
nand U3265 (N_3265,N_2463,N_1596);
nor U3266 (N_3266,N_2465,N_2444);
or U3267 (N_3267,N_729,N_1769);
nor U3268 (N_3268,N_360,N_7);
nand U3269 (N_3269,N_1458,N_113);
and U3270 (N_3270,N_1844,N_874);
and U3271 (N_3271,N_291,N_198);
and U3272 (N_3272,N_2067,N_2);
nand U3273 (N_3273,N_1019,N_665);
nand U3274 (N_3274,N_1652,N_210);
or U3275 (N_3275,N_1474,N_915);
or U3276 (N_3276,N_1262,N_2436);
or U3277 (N_3277,N_186,N_2108);
or U3278 (N_3278,N_726,N_1690);
nand U3279 (N_3279,N_1064,N_236);
nor U3280 (N_3280,N_1730,N_381);
nand U3281 (N_3281,N_960,N_831);
nor U3282 (N_3282,N_995,N_414);
and U3283 (N_3283,N_205,N_1495);
nor U3284 (N_3284,N_1276,N_2118);
and U3285 (N_3285,N_824,N_1104);
and U3286 (N_3286,N_2216,N_528);
and U3287 (N_3287,N_2215,N_376);
nand U3288 (N_3288,N_482,N_2282);
nor U3289 (N_3289,N_530,N_57);
nand U3290 (N_3290,N_329,N_579);
or U3291 (N_3291,N_2004,N_672);
or U3292 (N_3292,N_870,N_961);
or U3293 (N_3293,N_219,N_471);
or U3294 (N_3294,N_243,N_696);
nand U3295 (N_3295,N_24,N_2456);
or U3296 (N_3296,N_1809,N_2498);
nor U3297 (N_3297,N_630,N_1132);
and U3298 (N_3298,N_1066,N_1336);
nand U3299 (N_3299,N_1333,N_2405);
nand U3300 (N_3300,N_2006,N_237);
and U3301 (N_3301,N_1713,N_371);
nand U3302 (N_3302,N_892,N_1485);
and U3303 (N_3303,N_1572,N_341);
and U3304 (N_3304,N_284,N_871);
nand U3305 (N_3305,N_2117,N_2390);
nand U3306 (N_3306,N_1635,N_1313);
or U3307 (N_3307,N_2219,N_188);
nor U3308 (N_3308,N_1082,N_1978);
nand U3309 (N_3309,N_2496,N_799);
nand U3310 (N_3310,N_1670,N_365);
and U3311 (N_3311,N_1438,N_591);
and U3312 (N_3312,N_1840,N_173);
and U3313 (N_3313,N_208,N_1248);
and U3314 (N_3314,N_2087,N_1170);
nor U3315 (N_3315,N_1673,N_201);
and U3316 (N_3316,N_1613,N_740);
and U3317 (N_3317,N_1584,N_2309);
or U3318 (N_3318,N_1097,N_1517);
nor U3319 (N_3319,N_1465,N_1209);
and U3320 (N_3320,N_2410,N_2053);
nand U3321 (N_3321,N_1024,N_258);
nor U3322 (N_3322,N_577,N_406);
nand U3323 (N_3323,N_6,N_330);
or U3324 (N_3324,N_965,N_81);
nand U3325 (N_3325,N_2373,N_350);
nor U3326 (N_3326,N_885,N_1826);
and U3327 (N_3327,N_307,N_2336);
or U3328 (N_3328,N_571,N_511);
and U3329 (N_3329,N_478,N_174);
nor U3330 (N_3330,N_994,N_2459);
and U3331 (N_3331,N_1841,N_1862);
nand U3332 (N_3332,N_1189,N_2200);
nor U3333 (N_3333,N_127,N_21);
and U3334 (N_3334,N_1219,N_2048);
nand U3335 (N_3335,N_1470,N_1446);
nor U3336 (N_3336,N_217,N_1955);
nor U3337 (N_3337,N_1187,N_1027);
nand U3338 (N_3338,N_311,N_1378);
and U3339 (N_3339,N_2135,N_2209);
nor U3340 (N_3340,N_1442,N_861);
or U3341 (N_3341,N_535,N_1816);
nand U3342 (N_3342,N_2015,N_1732);
nand U3343 (N_3343,N_1292,N_1138);
nor U3344 (N_3344,N_479,N_836);
and U3345 (N_3345,N_1555,N_149);
nand U3346 (N_3346,N_847,N_2265);
or U3347 (N_3347,N_2299,N_1390);
and U3348 (N_3348,N_1971,N_2031);
nor U3349 (N_3349,N_1589,N_1473);
and U3350 (N_3350,N_2227,N_35);
nor U3351 (N_3351,N_655,N_2194);
or U3352 (N_3352,N_108,N_1666);
nor U3353 (N_3353,N_211,N_1095);
and U3354 (N_3354,N_549,N_332);
nor U3355 (N_3355,N_2424,N_2212);
or U3356 (N_3356,N_1961,N_2304);
nor U3357 (N_3357,N_546,N_950);
nand U3358 (N_3358,N_1740,N_601);
nor U3359 (N_3359,N_154,N_986);
nor U3360 (N_3360,N_2495,N_951);
nand U3361 (N_3361,N_669,N_1146);
nor U3362 (N_3362,N_391,N_1887);
nand U3363 (N_3363,N_766,N_1460);
and U3364 (N_3364,N_68,N_2052);
or U3365 (N_3365,N_1750,N_1267);
or U3366 (N_3366,N_56,N_1397);
nand U3367 (N_3367,N_1979,N_2181);
nand U3368 (N_3368,N_2301,N_449);
nor U3369 (N_3369,N_1640,N_63);
nor U3370 (N_3370,N_1830,N_2419);
nor U3371 (N_3371,N_2261,N_553);
nand U3372 (N_3372,N_1159,N_1338);
nand U3373 (N_3373,N_339,N_1754);
and U3374 (N_3374,N_160,N_1708);
and U3375 (N_3375,N_754,N_2455);
nor U3376 (N_3376,N_1364,N_1366);
nor U3377 (N_3377,N_2040,N_51);
nand U3378 (N_3378,N_461,N_1720);
nor U3379 (N_3379,N_1075,N_1602);
and U3380 (N_3380,N_139,N_457);
nor U3381 (N_3381,N_979,N_310);
nor U3382 (N_3382,N_2485,N_2379);
or U3383 (N_3383,N_998,N_2355);
and U3384 (N_3384,N_1875,N_1883);
nand U3385 (N_3385,N_727,N_927);
nand U3386 (N_3386,N_1287,N_223);
nand U3387 (N_3387,N_14,N_1616);
or U3388 (N_3388,N_1703,N_1379);
and U3389 (N_3389,N_2464,N_2122);
or U3390 (N_3390,N_277,N_627);
and U3391 (N_3391,N_1683,N_2258);
or U3392 (N_3392,N_1685,N_1884);
nand U3393 (N_3393,N_2394,N_1575);
nand U3394 (N_3394,N_739,N_506);
nand U3395 (N_3395,N_556,N_784);
and U3396 (N_3396,N_657,N_215);
or U3397 (N_3397,N_1372,N_1286);
or U3398 (N_3398,N_33,N_1902);
nand U3399 (N_3399,N_2283,N_2196);
or U3400 (N_3400,N_107,N_922);
nand U3401 (N_3401,N_2469,N_1013);
and U3402 (N_3402,N_119,N_1255);
or U3403 (N_3403,N_899,N_1113);
nor U3404 (N_3404,N_1411,N_1199);
nand U3405 (N_3405,N_2192,N_564);
and U3406 (N_3406,N_491,N_2163);
and U3407 (N_3407,N_1581,N_626);
nor U3408 (N_3408,N_2427,N_1000);
or U3409 (N_3409,N_1253,N_1743);
nor U3410 (N_3410,N_962,N_933);
and U3411 (N_3411,N_2225,N_483);
nor U3412 (N_3412,N_1706,N_875);
nand U3413 (N_3413,N_970,N_74);
and U3414 (N_3414,N_1237,N_774);
nand U3415 (N_3415,N_744,N_1353);
or U3416 (N_3416,N_308,N_866);
nor U3417 (N_3417,N_150,N_2082);
nor U3418 (N_3418,N_1737,N_1348);
nand U3419 (N_3419,N_715,N_793);
nand U3420 (N_3420,N_2489,N_1041);
nor U3421 (N_3421,N_233,N_2322);
nand U3422 (N_3422,N_1622,N_936);
nand U3423 (N_3423,N_1853,N_707);
nand U3424 (N_3424,N_1532,N_448);
nor U3425 (N_3425,N_1370,N_1462);
nand U3426 (N_3426,N_1646,N_1901);
nand U3427 (N_3427,N_27,N_1519);
and U3428 (N_3428,N_1619,N_1797);
or U3429 (N_3429,N_82,N_66);
or U3430 (N_3430,N_1045,N_338);
or U3431 (N_3431,N_2076,N_1203);
nand U3432 (N_3432,N_1643,N_811);
nor U3433 (N_3433,N_624,N_1888);
nor U3434 (N_3434,N_1106,N_570);
nand U3435 (N_3435,N_2458,N_822);
and U3436 (N_3436,N_692,N_1781);
nor U3437 (N_3437,N_714,N_190);
or U3438 (N_3438,N_648,N_1078);
and U3439 (N_3439,N_2214,N_232);
and U3440 (N_3440,N_2228,N_2411);
and U3441 (N_3441,N_763,N_1724);
nor U3442 (N_3442,N_131,N_1776);
or U3443 (N_3443,N_1243,N_797);
nor U3444 (N_3444,N_393,N_1744);
nand U3445 (N_3445,N_647,N_72);
nor U3446 (N_3446,N_2172,N_388);
nor U3447 (N_3447,N_1912,N_1538);
nand U3448 (N_3448,N_852,N_409);
nand U3449 (N_3449,N_1922,N_1389);
and U3450 (N_3450,N_1281,N_103);
nor U3451 (N_3451,N_170,N_958);
or U3452 (N_3452,N_2316,N_43);
or U3453 (N_3453,N_2176,N_1648);
nand U3454 (N_3454,N_1739,N_1956);
nor U3455 (N_3455,N_2395,N_499);
xnor U3456 (N_3456,N_2332,N_2017);
and U3457 (N_3457,N_1546,N_2345);
nor U3458 (N_3458,N_1112,N_2476);
nand U3459 (N_3459,N_1444,N_568);
or U3460 (N_3460,N_1658,N_1065);
nand U3461 (N_3461,N_1254,N_2284);
nor U3462 (N_3462,N_659,N_2120);
and U3463 (N_3463,N_550,N_825);
nand U3464 (N_3464,N_1140,N_815);
nor U3465 (N_3465,N_2070,N_880);
and U3466 (N_3466,N_2348,N_60);
nor U3467 (N_3467,N_2492,N_216);
and U3468 (N_3468,N_985,N_2251);
and U3469 (N_3469,N_1583,N_2470);
or U3470 (N_3470,N_2211,N_1420);
and U3471 (N_3471,N_240,N_547);
or U3472 (N_3472,N_687,N_616);
nor U3473 (N_3473,N_1204,N_533);
nor U3474 (N_3474,N_2226,N_1793);
nor U3475 (N_3475,N_1873,N_419);
nand U3476 (N_3476,N_526,N_1016);
or U3477 (N_3477,N_184,N_539);
or U3478 (N_3478,N_1042,N_430);
nor U3479 (N_3479,N_47,N_854);
and U3480 (N_3480,N_460,N_957);
and U3481 (N_3481,N_520,N_1879);
xnor U3482 (N_3482,N_2201,N_628);
or U3483 (N_3483,N_2000,N_2177);
and U3484 (N_3484,N_639,N_1625);
nor U3485 (N_3485,N_1284,N_333);
and U3486 (N_3486,N_446,N_247);
or U3487 (N_3487,N_776,N_664);
and U3488 (N_3488,N_1617,N_118);
and U3489 (N_3489,N_2277,N_1456);
nor U3490 (N_3490,N_84,N_908);
and U3491 (N_3491,N_2487,N_1360);
xnor U3492 (N_3492,N_369,N_769);
and U3493 (N_3493,N_1022,N_941);
and U3494 (N_3494,N_581,N_1103);
nor U3495 (N_3495,N_276,N_1867);
and U3496 (N_3496,N_1123,N_1630);
nor U3497 (N_3497,N_20,N_1259);
and U3498 (N_3498,N_1604,N_604);
nor U3499 (N_3499,N_2093,N_557);
and U3500 (N_3500,N_2308,N_428);
or U3501 (N_3501,N_1335,N_867);
nor U3502 (N_3502,N_1165,N_2069);
nor U3503 (N_3503,N_1270,N_463);
or U3504 (N_3504,N_2190,N_2360);
nor U3505 (N_3505,N_877,N_632);
nand U3506 (N_3506,N_2243,N_778);
or U3507 (N_3507,N_8,N_1275);
or U3508 (N_3508,N_924,N_397);
or U3509 (N_3509,N_78,N_275);
and U3510 (N_3510,N_204,N_337);
nand U3511 (N_3511,N_1761,N_169);
nand U3512 (N_3512,N_704,N_1196);
or U3513 (N_3513,N_2291,N_2313);
nand U3514 (N_3514,N_1116,N_1994);
xor U3515 (N_3515,N_1518,N_685);
nand U3516 (N_3516,N_1046,N_431);
nand U3517 (N_3517,N_1878,N_1786);
nand U3518 (N_3518,N_1603,N_133);
nand U3519 (N_3519,N_2407,N_2321);
xor U3520 (N_3520,N_667,N_1072);
nor U3521 (N_3521,N_1297,N_302);
or U3522 (N_3522,N_599,N_250);
or U3523 (N_3523,N_2272,N_1711);
and U3524 (N_3524,N_1591,N_1239);
and U3525 (N_3525,N_2210,N_1145);
nand U3526 (N_3526,N_227,N_2239);
nand U3527 (N_3527,N_182,N_2494);
and U3528 (N_3528,N_2084,N_2144);
and U3529 (N_3529,N_264,N_1891);
and U3530 (N_3530,N_2270,N_1773);
or U3531 (N_3531,N_392,N_2245);
or U3532 (N_3532,N_1441,N_218);
nor U3533 (N_3533,N_2030,N_348);
nand U3534 (N_3534,N_1080,N_2365);
nand U3535 (N_3535,N_2044,N_1590);
or U3536 (N_3536,N_1241,N_1907);
or U3537 (N_3537,N_1315,N_1111);
and U3538 (N_3538,N_1309,N_534);
or U3539 (N_3539,N_328,N_2477);
nor U3540 (N_3540,N_1143,N_895);
nand U3541 (N_3541,N_2381,N_1489);
nand U3542 (N_3542,N_2061,N_1974);
nand U3543 (N_3543,N_676,N_829);
or U3544 (N_3544,N_231,N_2383);
nand U3545 (N_3545,N_1422,N_1368);
and U3546 (N_3546,N_1660,N_207);
and U3547 (N_3547,N_673,N_1455);
or U3548 (N_3548,N_734,N_540);
or U3549 (N_3549,N_1803,N_1038);
and U3550 (N_3550,N_351,N_410);
nor U3551 (N_3551,N_2036,N_1070);
nor U3552 (N_3552,N_512,N_791);
nand U3553 (N_3553,N_1890,N_1311);
nor U3554 (N_3554,N_1114,N_294);
or U3555 (N_3555,N_1481,N_832);
or U3556 (N_3556,N_827,N_272);
and U3557 (N_3557,N_2329,N_2438);
nor U3558 (N_3558,N_1388,N_1798);
nand U3559 (N_3559,N_1201,N_745);
and U3560 (N_3560,N_1599,N_1953);
or U3561 (N_3561,N_1003,N_1127);
nand U3562 (N_3562,N_1212,N_322);
or U3563 (N_3563,N_1639,N_544);
or U3564 (N_3564,N_1501,N_1002);
nand U3565 (N_3565,N_1139,N_1186);
nor U3566 (N_3566,N_1606,N_1245);
and U3567 (N_3567,N_2287,N_755);
nor U3568 (N_3568,N_1521,N_1547);
or U3569 (N_3569,N_375,N_1512);
and U3570 (N_3570,N_1258,N_1200);
or U3571 (N_3571,N_819,N_1686);
and U3572 (N_3572,N_975,N_1503);
nor U3573 (N_3573,N_2101,N_1691);
or U3574 (N_3574,N_835,N_1251);
nor U3575 (N_3575,N_731,N_2333);
and U3576 (N_3576,N_902,N_398);
nor U3577 (N_3577,N_1278,N_2479);
nor U3578 (N_3578,N_1457,N_2462);
nand U3579 (N_3579,N_126,N_1927);
or U3580 (N_3580,N_974,N_2140);
nand U3581 (N_3581,N_1371,N_354);
or U3582 (N_3582,N_519,N_1767);
or U3583 (N_3583,N_1725,N_2448);
nor U3584 (N_3584,N_1224,N_748);
nor U3585 (N_3585,N_2134,N_1476);
and U3586 (N_3586,N_674,N_693);
nor U3587 (N_3587,N_798,N_2326);
nor U3588 (N_3588,N_2139,N_1945);
nand U3589 (N_3589,N_649,N_54);
nand U3590 (N_3590,N_1939,N_1329);
and U3591 (N_3591,N_1193,N_1935);
or U3592 (N_3592,N_541,N_125);
xor U3593 (N_3593,N_418,N_1804);
and U3594 (N_3594,N_2387,N_1049);
or U3595 (N_3595,N_2404,N_387);
and U3596 (N_3596,N_224,N_952);
nand U3597 (N_3597,N_790,N_1295);
nor U3598 (N_3598,N_295,N_967);
and U3599 (N_3599,N_377,N_643);
or U3600 (N_3600,N_1693,N_2121);
and U3601 (N_3601,N_2224,N_1770);
nand U3602 (N_3602,N_1947,N_1328);
or U3603 (N_3603,N_1763,N_2437);
or U3604 (N_3604,N_1029,N_1510);
and U3605 (N_3605,N_1452,N_1607);
nor U3606 (N_3606,N_1944,N_2024);
and U3607 (N_3607,N_2198,N_681);
and U3608 (N_3608,N_1352,N_1865);
and U3609 (N_3609,N_1014,N_898);
nor U3610 (N_3610,N_855,N_1167);
and U3611 (N_3611,N_87,N_2011);
or U3612 (N_3612,N_1709,N_403);
or U3613 (N_3613,N_803,N_475);
nor U3614 (N_3614,N_841,N_1450);
or U3615 (N_3615,N_1771,N_1162);
nor U3616 (N_3616,N_181,N_932);
nand U3617 (N_3617,N_2034,N_913);
nor U3618 (N_3618,N_2080,N_1406);
and U3619 (N_3619,N_597,N_31);
nor U3620 (N_3620,N_1846,N_1308);
nand U3621 (N_3621,N_2346,N_2104);
or U3622 (N_3622,N_1558,N_783);
and U3623 (N_3623,N_1305,N_621);
or U3624 (N_3624,N_1892,N_1296);
nand U3625 (N_3625,N_1528,N_64);
or U3626 (N_3626,N_268,N_978);
nand U3627 (N_3627,N_61,N_753);
nor U3628 (N_3628,N_1805,N_1548);
and U3629 (N_3629,N_679,N_492);
nand U3630 (N_3630,N_1449,N_18);
and U3631 (N_3631,N_1677,N_1764);
and U3632 (N_3632,N_1244,N_1416);
nor U3633 (N_3633,N_1588,N_603);
and U3634 (N_3634,N_1549,N_2038);
nor U3635 (N_3635,N_652,N_1233);
nor U3636 (N_3636,N_2389,N_1085);
or U3637 (N_3637,N_1738,N_304);
nor U3638 (N_3638,N_2377,N_474);
or U3639 (N_3639,N_315,N_1929);
nand U3640 (N_3640,N_640,N_1);
or U3641 (N_3641,N_1290,N_488);
or U3642 (N_3642,N_1249,N_883);
and U3643 (N_3643,N_1256,N_1461);
and U3644 (N_3644,N_1808,N_1952);
and U3645 (N_3645,N_771,N_1477);
nand U3646 (N_3646,N_1247,N_1697);
xnor U3647 (N_3647,N_834,N_202);
nor U3648 (N_3648,N_1320,N_497);
nor U3649 (N_3649,N_619,N_2442);
and U3650 (N_3650,N_1857,N_945);
nand U3651 (N_3651,N_1834,N_407);
or U3652 (N_3652,N_2260,N_1976);
or U3653 (N_3653,N_2461,N_2374);
nor U3654 (N_3654,N_1345,N_2085);
or U3655 (N_3655,N_89,N_1392);
nand U3656 (N_3656,N_953,N_2376);
or U3657 (N_3657,N_1843,N_634);
or U3658 (N_3658,N_2130,N_2164);
or U3659 (N_3659,N_1068,N_2162);
or U3660 (N_3660,N_2451,N_566);
nand U3661 (N_3661,N_2353,N_1991);
xnor U3662 (N_3662,N_496,N_486);
and U3663 (N_3663,N_2195,N_287);
nor U3664 (N_3664,N_2372,N_612);
nor U3665 (N_3665,N_1728,N_1266);
nor U3666 (N_3666,N_1409,N_1675);
and U3667 (N_3667,N_1969,N_157);
or U3668 (N_3668,N_1505,N_802);
or U3669 (N_3669,N_738,N_2202);
and U3670 (N_3670,N_1747,N_595);
nand U3671 (N_3671,N_1210,N_2028);
nand U3672 (N_3672,N_2062,N_319);
nor U3673 (N_3673,N_699,N_1289);
nand U3674 (N_3674,N_1981,N_879);
nor U3675 (N_3675,N_301,N_1238);
and U3676 (N_3676,N_823,N_336);
nand U3677 (N_3677,N_1906,N_1414);
and U3678 (N_3678,N_1864,N_801);
nor U3679 (N_3679,N_1383,N_2001);
and U3680 (N_3680,N_2497,N_25);
and U3681 (N_3681,N_465,N_1171);
and U3682 (N_3682,N_1800,N_662);
nor U3683 (N_3683,N_1656,N_529);
and U3684 (N_3684,N_1756,N_1751);
and U3685 (N_3685,N_2173,N_1017);
or U3686 (N_3686,N_1876,N_2183);
nand U3687 (N_3687,N_732,N_1930);
nor U3688 (N_3688,N_2126,N_312);
nor U3689 (N_3689,N_602,N_536);
nand U3690 (N_3690,N_1304,N_1926);
and U3691 (N_3691,N_1181,N_2199);
nand U3692 (N_3692,N_1339,N_1882);
nor U3693 (N_3693,N_1044,N_999);
and U3694 (N_3694,N_1916,N_1988);
nand U3695 (N_3695,N_1676,N_1775);
nor U3696 (N_3696,N_65,N_1959);
or U3697 (N_3697,N_1169,N_2259);
nand U3698 (N_3698,N_2249,N_2493);
nand U3699 (N_3699,N_1299,N_2324);
or U3700 (N_3700,N_816,N_50);
nand U3701 (N_3701,N_1062,N_505);
nor U3702 (N_3702,N_77,N_1852);
or U3703 (N_3703,N_2307,N_450);
or U3704 (N_3704,N_30,N_1984);
and U3705 (N_3705,N_493,N_1678);
and U3706 (N_3706,N_1672,N_195);
nor U3707 (N_3707,N_905,N_2012);
nor U3708 (N_3708,N_910,N_1346);
or U3709 (N_3709,N_1982,N_1829);
nor U3710 (N_3710,N_1631,N_747);
nor U3711 (N_3711,N_1118,N_1051);
nor U3712 (N_3712,N_725,N_590);
nor U3713 (N_3713,N_1156,N_2241);
nor U3714 (N_3714,N_2125,N_592);
nand U3715 (N_3715,N_1100,N_1562);
nor U3716 (N_3716,N_1783,N_610);
or U3717 (N_3717,N_1073,N_812);
and U3718 (N_3718,N_11,N_671);
and U3719 (N_3719,N_424,N_1122);
and U3720 (N_3720,N_1772,N_2111);
or U3721 (N_3721,N_367,N_2218);
nor U3722 (N_3722,N_959,N_2103);
or U3723 (N_3723,N_809,N_2019);
nand U3724 (N_3724,N_1937,N_221);
nand U3725 (N_3725,N_2089,N_1700);
or U3726 (N_3726,N_1190,N_1727);
nor U3727 (N_3727,N_462,N_1574);
or U3728 (N_3728,N_22,N_697);
nor U3729 (N_3729,N_123,N_1791);
and U3730 (N_3730,N_1351,N_786);
nand U3731 (N_3731,N_2189,N_1494);
nand U3732 (N_3732,N_1610,N_2159);
and U3733 (N_3733,N_1310,N_1765);
nand U3734 (N_3734,N_868,N_1380);
nand U3735 (N_3735,N_2312,N_1942);
nand U3736 (N_3736,N_2142,N_141);
nand U3737 (N_3737,N_1881,N_234);
or U3738 (N_3738,N_110,N_2362);
or U3739 (N_3739,N_52,N_2109);
nor U3740 (N_3740,N_2220,N_2003);
xnor U3741 (N_3741,N_1885,N_2184);
nand U3742 (N_3742,N_176,N_1502);
nor U3743 (N_3743,N_1949,N_569);
or U3744 (N_3744,N_1802,N_1758);
nor U3745 (N_3745,N_668,N_1566);
and U3746 (N_3746,N_120,N_1948);
nand U3747 (N_3747,N_1207,N_2221);
and U3748 (N_3748,N_2207,N_1108);
nand U3749 (N_3749,N_252,N_851);
and U3750 (N_3750,N_235,N_1560);
nand U3751 (N_3751,N_2258,N_720);
nor U3752 (N_3752,N_1541,N_1769);
nand U3753 (N_3753,N_2255,N_265);
or U3754 (N_3754,N_1727,N_1025);
nand U3755 (N_3755,N_2361,N_1460);
nor U3756 (N_3756,N_759,N_1993);
and U3757 (N_3757,N_2006,N_625);
nor U3758 (N_3758,N_1886,N_2024);
or U3759 (N_3759,N_352,N_995);
nor U3760 (N_3760,N_660,N_2108);
or U3761 (N_3761,N_1360,N_704);
nand U3762 (N_3762,N_1030,N_2391);
nand U3763 (N_3763,N_2296,N_1585);
or U3764 (N_3764,N_2085,N_40);
or U3765 (N_3765,N_2117,N_1128);
nor U3766 (N_3766,N_1518,N_2128);
and U3767 (N_3767,N_882,N_2475);
nand U3768 (N_3768,N_1346,N_894);
nor U3769 (N_3769,N_1727,N_217);
nand U3770 (N_3770,N_1945,N_1964);
nand U3771 (N_3771,N_802,N_969);
nand U3772 (N_3772,N_400,N_1893);
and U3773 (N_3773,N_1779,N_640);
nand U3774 (N_3774,N_598,N_1112);
or U3775 (N_3775,N_247,N_725);
nor U3776 (N_3776,N_735,N_2248);
nor U3777 (N_3777,N_950,N_2176);
and U3778 (N_3778,N_1687,N_1043);
and U3779 (N_3779,N_314,N_28);
nand U3780 (N_3780,N_2298,N_2183);
and U3781 (N_3781,N_1191,N_420);
or U3782 (N_3782,N_904,N_2148);
and U3783 (N_3783,N_189,N_817);
nor U3784 (N_3784,N_988,N_1699);
or U3785 (N_3785,N_561,N_904);
nor U3786 (N_3786,N_1368,N_804);
and U3787 (N_3787,N_1441,N_1866);
nor U3788 (N_3788,N_266,N_1464);
and U3789 (N_3789,N_2271,N_180);
or U3790 (N_3790,N_760,N_411);
and U3791 (N_3791,N_878,N_174);
nand U3792 (N_3792,N_1213,N_544);
nor U3793 (N_3793,N_128,N_1941);
and U3794 (N_3794,N_1583,N_433);
nand U3795 (N_3795,N_530,N_2293);
or U3796 (N_3796,N_949,N_2432);
nor U3797 (N_3797,N_797,N_2093);
and U3798 (N_3798,N_1815,N_2048);
and U3799 (N_3799,N_2195,N_948);
or U3800 (N_3800,N_339,N_362);
or U3801 (N_3801,N_1508,N_1937);
and U3802 (N_3802,N_1391,N_2463);
nor U3803 (N_3803,N_2185,N_1595);
or U3804 (N_3804,N_2312,N_138);
or U3805 (N_3805,N_66,N_456);
nand U3806 (N_3806,N_2430,N_129);
nor U3807 (N_3807,N_1628,N_1922);
or U3808 (N_3808,N_1936,N_1475);
or U3809 (N_3809,N_278,N_486);
nand U3810 (N_3810,N_2289,N_1915);
nand U3811 (N_3811,N_109,N_976);
nand U3812 (N_3812,N_693,N_1801);
nor U3813 (N_3813,N_953,N_1707);
or U3814 (N_3814,N_365,N_368);
nand U3815 (N_3815,N_348,N_1432);
or U3816 (N_3816,N_219,N_1202);
or U3817 (N_3817,N_49,N_178);
nand U3818 (N_3818,N_1000,N_2039);
or U3819 (N_3819,N_1051,N_1669);
nand U3820 (N_3820,N_526,N_1769);
nand U3821 (N_3821,N_1648,N_1151);
and U3822 (N_3822,N_1210,N_577);
and U3823 (N_3823,N_845,N_148);
nand U3824 (N_3824,N_2403,N_1759);
or U3825 (N_3825,N_586,N_2378);
or U3826 (N_3826,N_879,N_1889);
or U3827 (N_3827,N_1875,N_424);
and U3828 (N_3828,N_528,N_981);
or U3829 (N_3829,N_573,N_499);
and U3830 (N_3830,N_310,N_1151);
nand U3831 (N_3831,N_1501,N_1631);
and U3832 (N_3832,N_291,N_1155);
and U3833 (N_3833,N_1370,N_294);
or U3834 (N_3834,N_2013,N_429);
xor U3835 (N_3835,N_2324,N_2348);
nor U3836 (N_3836,N_2430,N_1569);
and U3837 (N_3837,N_414,N_790);
nand U3838 (N_3838,N_1423,N_2164);
nand U3839 (N_3839,N_2411,N_691);
and U3840 (N_3840,N_2359,N_1936);
nor U3841 (N_3841,N_1028,N_1074);
and U3842 (N_3842,N_816,N_1131);
nand U3843 (N_3843,N_1004,N_2490);
nand U3844 (N_3844,N_1517,N_861);
nand U3845 (N_3845,N_1063,N_2095);
or U3846 (N_3846,N_2303,N_1339);
nand U3847 (N_3847,N_1953,N_2220);
nand U3848 (N_3848,N_179,N_1923);
nor U3849 (N_3849,N_370,N_256);
and U3850 (N_3850,N_1570,N_714);
or U3851 (N_3851,N_692,N_931);
or U3852 (N_3852,N_2346,N_959);
and U3853 (N_3853,N_686,N_1393);
nand U3854 (N_3854,N_638,N_1386);
and U3855 (N_3855,N_1805,N_1574);
nor U3856 (N_3856,N_379,N_185);
nand U3857 (N_3857,N_1642,N_563);
and U3858 (N_3858,N_1575,N_2253);
and U3859 (N_3859,N_596,N_1618);
and U3860 (N_3860,N_580,N_2045);
nand U3861 (N_3861,N_1843,N_461);
or U3862 (N_3862,N_9,N_1892);
nor U3863 (N_3863,N_2083,N_489);
and U3864 (N_3864,N_685,N_1188);
and U3865 (N_3865,N_1401,N_2453);
nor U3866 (N_3866,N_430,N_2273);
and U3867 (N_3867,N_1458,N_145);
and U3868 (N_3868,N_1245,N_120);
nor U3869 (N_3869,N_1072,N_1975);
nand U3870 (N_3870,N_410,N_2277);
and U3871 (N_3871,N_565,N_705);
and U3872 (N_3872,N_398,N_2207);
nand U3873 (N_3873,N_1518,N_605);
and U3874 (N_3874,N_771,N_1274);
nand U3875 (N_3875,N_443,N_545);
xnor U3876 (N_3876,N_1131,N_207);
and U3877 (N_3877,N_1293,N_1362);
nand U3878 (N_3878,N_1644,N_189);
nand U3879 (N_3879,N_2498,N_2092);
nand U3880 (N_3880,N_2433,N_2248);
and U3881 (N_3881,N_1164,N_2185);
and U3882 (N_3882,N_458,N_938);
or U3883 (N_3883,N_1497,N_783);
and U3884 (N_3884,N_1285,N_56);
and U3885 (N_3885,N_1185,N_2484);
nor U3886 (N_3886,N_2085,N_1256);
nor U3887 (N_3887,N_1374,N_895);
or U3888 (N_3888,N_791,N_1126);
nor U3889 (N_3889,N_2099,N_1806);
nor U3890 (N_3890,N_533,N_1049);
or U3891 (N_3891,N_258,N_2217);
or U3892 (N_3892,N_2081,N_1524);
nor U3893 (N_3893,N_1916,N_1895);
nand U3894 (N_3894,N_811,N_1608);
nand U3895 (N_3895,N_1444,N_1723);
nor U3896 (N_3896,N_2012,N_186);
nor U3897 (N_3897,N_371,N_1733);
or U3898 (N_3898,N_1094,N_1236);
and U3899 (N_3899,N_2398,N_868);
nor U3900 (N_3900,N_390,N_1687);
nor U3901 (N_3901,N_1748,N_1724);
nor U3902 (N_3902,N_599,N_1477);
nor U3903 (N_3903,N_1651,N_1598);
nand U3904 (N_3904,N_2403,N_2012);
and U3905 (N_3905,N_19,N_2006);
nand U3906 (N_3906,N_298,N_903);
nand U3907 (N_3907,N_604,N_965);
or U3908 (N_3908,N_1660,N_290);
or U3909 (N_3909,N_898,N_303);
or U3910 (N_3910,N_1809,N_328);
nand U3911 (N_3911,N_615,N_227);
or U3912 (N_3912,N_614,N_387);
or U3913 (N_3913,N_416,N_2025);
or U3914 (N_3914,N_1151,N_499);
and U3915 (N_3915,N_1379,N_119);
or U3916 (N_3916,N_599,N_2287);
xor U3917 (N_3917,N_86,N_1435);
and U3918 (N_3918,N_449,N_871);
or U3919 (N_3919,N_1639,N_1123);
nand U3920 (N_3920,N_931,N_1438);
nand U3921 (N_3921,N_1267,N_59);
and U3922 (N_3922,N_1005,N_733);
nor U3923 (N_3923,N_1433,N_1711);
and U3924 (N_3924,N_2222,N_1292);
or U3925 (N_3925,N_1259,N_920);
nand U3926 (N_3926,N_2310,N_1006);
and U3927 (N_3927,N_560,N_339);
and U3928 (N_3928,N_163,N_288);
nand U3929 (N_3929,N_141,N_913);
or U3930 (N_3930,N_508,N_1052);
or U3931 (N_3931,N_1430,N_1697);
nand U3932 (N_3932,N_1247,N_1774);
or U3933 (N_3933,N_428,N_629);
nor U3934 (N_3934,N_731,N_450);
or U3935 (N_3935,N_752,N_1531);
nor U3936 (N_3936,N_186,N_314);
nand U3937 (N_3937,N_2000,N_1860);
nand U3938 (N_3938,N_348,N_651);
nor U3939 (N_3939,N_1562,N_2042);
and U3940 (N_3940,N_1412,N_1661);
or U3941 (N_3941,N_897,N_159);
nand U3942 (N_3942,N_671,N_1545);
and U3943 (N_3943,N_184,N_945);
or U3944 (N_3944,N_2470,N_1191);
or U3945 (N_3945,N_1183,N_1317);
nand U3946 (N_3946,N_419,N_203);
nor U3947 (N_3947,N_88,N_1367);
nand U3948 (N_3948,N_2390,N_1205);
nor U3949 (N_3949,N_1646,N_1670);
or U3950 (N_3950,N_1633,N_2356);
and U3951 (N_3951,N_1467,N_69);
and U3952 (N_3952,N_1476,N_1116);
nor U3953 (N_3953,N_557,N_975);
xor U3954 (N_3954,N_1256,N_1815);
or U3955 (N_3955,N_1730,N_574);
nor U3956 (N_3956,N_2098,N_1566);
nand U3957 (N_3957,N_735,N_1999);
or U3958 (N_3958,N_2018,N_1223);
nand U3959 (N_3959,N_2199,N_477);
nand U3960 (N_3960,N_491,N_816);
nor U3961 (N_3961,N_2461,N_670);
nor U3962 (N_3962,N_844,N_594);
nor U3963 (N_3963,N_1147,N_831);
or U3964 (N_3964,N_654,N_1816);
nand U3965 (N_3965,N_1367,N_521);
and U3966 (N_3966,N_2159,N_497);
nand U3967 (N_3967,N_1928,N_250);
nand U3968 (N_3968,N_476,N_414);
and U3969 (N_3969,N_1513,N_816);
or U3970 (N_3970,N_1912,N_164);
nor U3971 (N_3971,N_1812,N_594);
or U3972 (N_3972,N_879,N_1178);
or U3973 (N_3973,N_768,N_2316);
or U3974 (N_3974,N_469,N_698);
and U3975 (N_3975,N_780,N_770);
nand U3976 (N_3976,N_772,N_2);
and U3977 (N_3977,N_2450,N_2309);
and U3978 (N_3978,N_572,N_268);
and U3979 (N_3979,N_1427,N_319);
or U3980 (N_3980,N_2454,N_701);
nor U3981 (N_3981,N_895,N_2194);
nand U3982 (N_3982,N_698,N_2402);
and U3983 (N_3983,N_432,N_231);
nand U3984 (N_3984,N_548,N_1047);
or U3985 (N_3985,N_938,N_754);
nand U3986 (N_3986,N_2072,N_104);
nand U3987 (N_3987,N_984,N_333);
or U3988 (N_3988,N_1771,N_2495);
nand U3989 (N_3989,N_926,N_2290);
nor U3990 (N_3990,N_1789,N_2471);
nor U3991 (N_3991,N_1986,N_2486);
or U3992 (N_3992,N_803,N_2402);
or U3993 (N_3993,N_2185,N_1348);
and U3994 (N_3994,N_1744,N_1455);
and U3995 (N_3995,N_1658,N_345);
nor U3996 (N_3996,N_930,N_2193);
and U3997 (N_3997,N_2241,N_2105);
nand U3998 (N_3998,N_2475,N_1139);
xnor U3999 (N_3999,N_1358,N_1729);
nand U4000 (N_4000,N_1147,N_1152);
nand U4001 (N_4001,N_1763,N_1275);
and U4002 (N_4002,N_260,N_527);
nand U4003 (N_4003,N_1036,N_1952);
and U4004 (N_4004,N_1903,N_1322);
and U4005 (N_4005,N_2410,N_998);
or U4006 (N_4006,N_2389,N_1678);
nor U4007 (N_4007,N_260,N_2041);
and U4008 (N_4008,N_1148,N_581);
nor U4009 (N_4009,N_493,N_859);
or U4010 (N_4010,N_986,N_1661);
or U4011 (N_4011,N_505,N_929);
nand U4012 (N_4012,N_33,N_2110);
nand U4013 (N_4013,N_458,N_510);
or U4014 (N_4014,N_2453,N_698);
or U4015 (N_4015,N_1010,N_1036);
nand U4016 (N_4016,N_1539,N_146);
nand U4017 (N_4017,N_2397,N_346);
and U4018 (N_4018,N_1669,N_788);
nand U4019 (N_4019,N_1380,N_1054);
nor U4020 (N_4020,N_468,N_2361);
nand U4021 (N_4021,N_1932,N_366);
nor U4022 (N_4022,N_2142,N_1246);
nor U4023 (N_4023,N_1844,N_2240);
and U4024 (N_4024,N_128,N_105);
nor U4025 (N_4025,N_211,N_1059);
nor U4026 (N_4026,N_1352,N_1057);
nand U4027 (N_4027,N_1170,N_634);
nor U4028 (N_4028,N_369,N_2215);
and U4029 (N_4029,N_134,N_497);
nor U4030 (N_4030,N_2388,N_2167);
nor U4031 (N_4031,N_1033,N_428);
nand U4032 (N_4032,N_777,N_1633);
or U4033 (N_4033,N_1497,N_707);
or U4034 (N_4034,N_1587,N_800);
nor U4035 (N_4035,N_2251,N_1258);
nand U4036 (N_4036,N_1600,N_1286);
nand U4037 (N_4037,N_926,N_2043);
and U4038 (N_4038,N_674,N_39);
nor U4039 (N_4039,N_2109,N_707);
or U4040 (N_4040,N_353,N_1596);
and U4041 (N_4041,N_1110,N_746);
nand U4042 (N_4042,N_190,N_1473);
nor U4043 (N_4043,N_1476,N_2438);
nor U4044 (N_4044,N_676,N_960);
nand U4045 (N_4045,N_157,N_2061);
nor U4046 (N_4046,N_1815,N_1230);
nor U4047 (N_4047,N_2229,N_825);
or U4048 (N_4048,N_1448,N_2236);
nor U4049 (N_4049,N_488,N_1367);
nor U4050 (N_4050,N_1125,N_1538);
nand U4051 (N_4051,N_1124,N_114);
nand U4052 (N_4052,N_512,N_1219);
nand U4053 (N_4053,N_1211,N_1485);
nand U4054 (N_4054,N_187,N_114);
nand U4055 (N_4055,N_57,N_1954);
and U4056 (N_4056,N_2083,N_966);
nor U4057 (N_4057,N_1265,N_1071);
nor U4058 (N_4058,N_1102,N_1112);
nor U4059 (N_4059,N_1704,N_163);
or U4060 (N_4060,N_906,N_1063);
nor U4061 (N_4061,N_879,N_773);
and U4062 (N_4062,N_1281,N_1440);
nor U4063 (N_4063,N_2471,N_390);
nor U4064 (N_4064,N_1406,N_1848);
and U4065 (N_4065,N_1758,N_888);
nor U4066 (N_4066,N_821,N_2376);
and U4067 (N_4067,N_488,N_298);
nand U4068 (N_4068,N_1539,N_991);
or U4069 (N_4069,N_766,N_135);
or U4070 (N_4070,N_527,N_2225);
nand U4071 (N_4071,N_428,N_1809);
and U4072 (N_4072,N_63,N_861);
nand U4073 (N_4073,N_82,N_1793);
nand U4074 (N_4074,N_2240,N_2204);
nor U4075 (N_4075,N_2138,N_2189);
and U4076 (N_4076,N_1760,N_1241);
and U4077 (N_4077,N_611,N_1595);
nand U4078 (N_4078,N_2040,N_903);
nand U4079 (N_4079,N_735,N_443);
nand U4080 (N_4080,N_204,N_744);
or U4081 (N_4081,N_368,N_1122);
or U4082 (N_4082,N_1114,N_1678);
nor U4083 (N_4083,N_288,N_511);
nand U4084 (N_4084,N_1942,N_13);
nand U4085 (N_4085,N_2104,N_703);
nand U4086 (N_4086,N_2403,N_2395);
nor U4087 (N_4087,N_243,N_564);
and U4088 (N_4088,N_2146,N_1932);
and U4089 (N_4089,N_1797,N_45);
nand U4090 (N_4090,N_341,N_1806);
or U4091 (N_4091,N_1810,N_2334);
nor U4092 (N_4092,N_1624,N_19);
nand U4093 (N_4093,N_1702,N_1365);
nand U4094 (N_4094,N_515,N_864);
or U4095 (N_4095,N_156,N_1768);
nor U4096 (N_4096,N_2467,N_933);
and U4097 (N_4097,N_1255,N_1665);
and U4098 (N_4098,N_1560,N_688);
nor U4099 (N_4099,N_2283,N_302);
or U4100 (N_4100,N_417,N_953);
nor U4101 (N_4101,N_1307,N_1892);
and U4102 (N_4102,N_269,N_734);
or U4103 (N_4103,N_74,N_1290);
or U4104 (N_4104,N_82,N_1534);
and U4105 (N_4105,N_2265,N_933);
or U4106 (N_4106,N_889,N_485);
and U4107 (N_4107,N_661,N_2457);
nor U4108 (N_4108,N_1126,N_164);
nor U4109 (N_4109,N_2211,N_704);
and U4110 (N_4110,N_1567,N_453);
nand U4111 (N_4111,N_2003,N_1774);
nor U4112 (N_4112,N_1043,N_1306);
nor U4113 (N_4113,N_980,N_1177);
nand U4114 (N_4114,N_1760,N_1849);
nand U4115 (N_4115,N_1166,N_1886);
nand U4116 (N_4116,N_263,N_1142);
nand U4117 (N_4117,N_1014,N_1124);
or U4118 (N_4118,N_1246,N_859);
or U4119 (N_4119,N_1045,N_1770);
nand U4120 (N_4120,N_1285,N_1861);
and U4121 (N_4121,N_753,N_965);
nand U4122 (N_4122,N_401,N_1188);
and U4123 (N_4123,N_500,N_620);
and U4124 (N_4124,N_1089,N_1756);
or U4125 (N_4125,N_57,N_1239);
or U4126 (N_4126,N_2379,N_1998);
nand U4127 (N_4127,N_838,N_831);
nand U4128 (N_4128,N_1755,N_24);
and U4129 (N_4129,N_1148,N_2111);
nor U4130 (N_4130,N_1659,N_297);
nor U4131 (N_4131,N_652,N_1469);
nor U4132 (N_4132,N_205,N_1370);
and U4133 (N_4133,N_1907,N_1801);
or U4134 (N_4134,N_2124,N_903);
nand U4135 (N_4135,N_891,N_185);
nand U4136 (N_4136,N_2095,N_1333);
nor U4137 (N_4137,N_1222,N_1410);
nor U4138 (N_4138,N_2383,N_1685);
and U4139 (N_4139,N_1352,N_586);
or U4140 (N_4140,N_307,N_441);
and U4141 (N_4141,N_2131,N_888);
and U4142 (N_4142,N_2380,N_2067);
or U4143 (N_4143,N_1175,N_1138);
nand U4144 (N_4144,N_620,N_2144);
or U4145 (N_4145,N_26,N_1520);
nor U4146 (N_4146,N_523,N_1807);
or U4147 (N_4147,N_675,N_1584);
nor U4148 (N_4148,N_1927,N_253);
and U4149 (N_4149,N_1993,N_1888);
nor U4150 (N_4150,N_295,N_691);
nand U4151 (N_4151,N_1227,N_2128);
nor U4152 (N_4152,N_523,N_403);
nor U4153 (N_4153,N_1723,N_2188);
nor U4154 (N_4154,N_2144,N_1785);
and U4155 (N_4155,N_1086,N_2122);
nor U4156 (N_4156,N_264,N_1628);
xor U4157 (N_4157,N_202,N_1153);
or U4158 (N_4158,N_1417,N_108);
nor U4159 (N_4159,N_1101,N_251);
and U4160 (N_4160,N_1903,N_1231);
or U4161 (N_4161,N_2493,N_1207);
or U4162 (N_4162,N_540,N_1855);
and U4163 (N_4163,N_1340,N_1165);
nand U4164 (N_4164,N_1199,N_363);
or U4165 (N_4165,N_2004,N_1631);
and U4166 (N_4166,N_133,N_1290);
nand U4167 (N_4167,N_1050,N_1981);
and U4168 (N_4168,N_610,N_117);
and U4169 (N_4169,N_1538,N_1492);
nor U4170 (N_4170,N_1759,N_1745);
or U4171 (N_4171,N_1930,N_1191);
nand U4172 (N_4172,N_1247,N_621);
nor U4173 (N_4173,N_1330,N_2365);
or U4174 (N_4174,N_2000,N_760);
or U4175 (N_4175,N_261,N_1068);
nor U4176 (N_4176,N_662,N_1211);
nor U4177 (N_4177,N_769,N_218);
nor U4178 (N_4178,N_1950,N_859);
or U4179 (N_4179,N_1626,N_999);
and U4180 (N_4180,N_916,N_2443);
and U4181 (N_4181,N_118,N_911);
and U4182 (N_4182,N_1152,N_1309);
nand U4183 (N_4183,N_134,N_2100);
nor U4184 (N_4184,N_1108,N_210);
nor U4185 (N_4185,N_2349,N_1255);
nand U4186 (N_4186,N_1689,N_1067);
nor U4187 (N_4187,N_2070,N_205);
nor U4188 (N_4188,N_1294,N_1897);
nor U4189 (N_4189,N_2458,N_288);
or U4190 (N_4190,N_2343,N_2361);
and U4191 (N_4191,N_1376,N_2083);
nor U4192 (N_4192,N_2037,N_1468);
nand U4193 (N_4193,N_269,N_1749);
xor U4194 (N_4194,N_974,N_1765);
and U4195 (N_4195,N_1549,N_1967);
and U4196 (N_4196,N_672,N_1544);
and U4197 (N_4197,N_1545,N_666);
or U4198 (N_4198,N_1595,N_1193);
and U4199 (N_4199,N_1711,N_1039);
nor U4200 (N_4200,N_17,N_1591);
and U4201 (N_4201,N_2417,N_2261);
nor U4202 (N_4202,N_1372,N_489);
nor U4203 (N_4203,N_2244,N_398);
or U4204 (N_4204,N_1411,N_200);
nand U4205 (N_4205,N_135,N_1773);
or U4206 (N_4206,N_2229,N_5);
xor U4207 (N_4207,N_1148,N_1180);
nor U4208 (N_4208,N_538,N_1851);
or U4209 (N_4209,N_26,N_1498);
nand U4210 (N_4210,N_1657,N_4);
or U4211 (N_4211,N_79,N_63);
and U4212 (N_4212,N_2392,N_49);
nand U4213 (N_4213,N_2376,N_2289);
and U4214 (N_4214,N_1637,N_570);
nor U4215 (N_4215,N_569,N_2247);
and U4216 (N_4216,N_2458,N_316);
nor U4217 (N_4217,N_350,N_1548);
nor U4218 (N_4218,N_759,N_2337);
and U4219 (N_4219,N_296,N_1933);
nand U4220 (N_4220,N_850,N_2167);
nor U4221 (N_4221,N_1458,N_2237);
and U4222 (N_4222,N_1928,N_981);
nand U4223 (N_4223,N_42,N_1027);
nor U4224 (N_4224,N_1051,N_1896);
and U4225 (N_4225,N_1261,N_1100);
or U4226 (N_4226,N_913,N_1033);
nor U4227 (N_4227,N_2092,N_925);
nor U4228 (N_4228,N_679,N_489);
nor U4229 (N_4229,N_136,N_366);
and U4230 (N_4230,N_1162,N_275);
nor U4231 (N_4231,N_30,N_385);
nor U4232 (N_4232,N_2402,N_13);
nor U4233 (N_4233,N_426,N_253);
nor U4234 (N_4234,N_1622,N_2131);
nand U4235 (N_4235,N_1519,N_860);
or U4236 (N_4236,N_2099,N_1704);
nand U4237 (N_4237,N_907,N_1447);
and U4238 (N_4238,N_1229,N_1963);
and U4239 (N_4239,N_2482,N_2463);
and U4240 (N_4240,N_1061,N_1226);
and U4241 (N_4241,N_2417,N_217);
nand U4242 (N_4242,N_2491,N_1009);
nand U4243 (N_4243,N_1065,N_1254);
nand U4244 (N_4244,N_1742,N_369);
and U4245 (N_4245,N_1617,N_1576);
nor U4246 (N_4246,N_1643,N_1453);
nand U4247 (N_4247,N_479,N_1228);
or U4248 (N_4248,N_557,N_957);
nor U4249 (N_4249,N_1276,N_2224);
or U4250 (N_4250,N_1150,N_1613);
nand U4251 (N_4251,N_2256,N_964);
or U4252 (N_4252,N_2042,N_1009);
or U4253 (N_4253,N_1676,N_961);
nor U4254 (N_4254,N_1190,N_25);
or U4255 (N_4255,N_388,N_1965);
and U4256 (N_4256,N_621,N_944);
or U4257 (N_4257,N_557,N_140);
nor U4258 (N_4258,N_2371,N_744);
nor U4259 (N_4259,N_1900,N_2331);
and U4260 (N_4260,N_1591,N_1819);
and U4261 (N_4261,N_2278,N_1901);
nor U4262 (N_4262,N_1312,N_446);
and U4263 (N_4263,N_1231,N_1102);
nor U4264 (N_4264,N_1386,N_63);
nor U4265 (N_4265,N_33,N_1612);
nand U4266 (N_4266,N_2218,N_90);
nor U4267 (N_4267,N_2339,N_880);
and U4268 (N_4268,N_2232,N_1244);
and U4269 (N_4269,N_2331,N_1086);
or U4270 (N_4270,N_418,N_1121);
nor U4271 (N_4271,N_2195,N_1871);
or U4272 (N_4272,N_1505,N_2141);
or U4273 (N_4273,N_2180,N_532);
and U4274 (N_4274,N_1212,N_1537);
or U4275 (N_4275,N_1631,N_2143);
xor U4276 (N_4276,N_2387,N_815);
and U4277 (N_4277,N_230,N_332);
nor U4278 (N_4278,N_2355,N_878);
and U4279 (N_4279,N_43,N_1225);
nand U4280 (N_4280,N_1273,N_1411);
and U4281 (N_4281,N_981,N_857);
and U4282 (N_4282,N_130,N_2424);
nand U4283 (N_4283,N_963,N_2229);
or U4284 (N_4284,N_1509,N_522);
nor U4285 (N_4285,N_2039,N_2091);
and U4286 (N_4286,N_58,N_2005);
nor U4287 (N_4287,N_1026,N_2067);
nand U4288 (N_4288,N_2087,N_229);
nor U4289 (N_4289,N_2283,N_777);
nor U4290 (N_4290,N_1946,N_921);
nor U4291 (N_4291,N_45,N_1163);
nand U4292 (N_4292,N_1034,N_2396);
nand U4293 (N_4293,N_553,N_1693);
and U4294 (N_4294,N_1803,N_884);
nor U4295 (N_4295,N_1766,N_290);
nor U4296 (N_4296,N_955,N_876);
and U4297 (N_4297,N_1539,N_72);
or U4298 (N_4298,N_965,N_433);
nor U4299 (N_4299,N_611,N_1024);
nor U4300 (N_4300,N_376,N_541);
nand U4301 (N_4301,N_1090,N_1473);
and U4302 (N_4302,N_365,N_2242);
or U4303 (N_4303,N_844,N_1573);
nor U4304 (N_4304,N_1081,N_2432);
nor U4305 (N_4305,N_388,N_897);
and U4306 (N_4306,N_2351,N_1578);
nand U4307 (N_4307,N_857,N_361);
and U4308 (N_4308,N_492,N_1703);
nand U4309 (N_4309,N_2145,N_1149);
nand U4310 (N_4310,N_1538,N_1950);
and U4311 (N_4311,N_2394,N_818);
nand U4312 (N_4312,N_1382,N_2270);
or U4313 (N_4313,N_2222,N_1077);
or U4314 (N_4314,N_525,N_560);
nor U4315 (N_4315,N_1118,N_582);
nand U4316 (N_4316,N_70,N_2331);
nand U4317 (N_4317,N_1274,N_478);
nand U4318 (N_4318,N_1663,N_1615);
nand U4319 (N_4319,N_1879,N_2421);
and U4320 (N_4320,N_977,N_1768);
or U4321 (N_4321,N_171,N_923);
nor U4322 (N_4322,N_218,N_89);
and U4323 (N_4323,N_2486,N_1399);
or U4324 (N_4324,N_695,N_2374);
nand U4325 (N_4325,N_645,N_2402);
or U4326 (N_4326,N_758,N_2390);
and U4327 (N_4327,N_1748,N_2377);
nor U4328 (N_4328,N_211,N_871);
and U4329 (N_4329,N_1041,N_685);
or U4330 (N_4330,N_363,N_852);
or U4331 (N_4331,N_1750,N_611);
nand U4332 (N_4332,N_1709,N_2003);
and U4333 (N_4333,N_100,N_1839);
or U4334 (N_4334,N_1300,N_819);
and U4335 (N_4335,N_2367,N_313);
nor U4336 (N_4336,N_350,N_1132);
or U4337 (N_4337,N_1453,N_451);
nor U4338 (N_4338,N_1495,N_1019);
and U4339 (N_4339,N_1034,N_1041);
or U4340 (N_4340,N_515,N_1581);
or U4341 (N_4341,N_1562,N_2114);
nand U4342 (N_4342,N_1233,N_2412);
nand U4343 (N_4343,N_150,N_2285);
nor U4344 (N_4344,N_1683,N_1448);
nand U4345 (N_4345,N_1397,N_565);
xor U4346 (N_4346,N_1899,N_1167);
and U4347 (N_4347,N_2281,N_2000);
nand U4348 (N_4348,N_1261,N_1305);
or U4349 (N_4349,N_2317,N_99);
or U4350 (N_4350,N_498,N_2334);
or U4351 (N_4351,N_1021,N_852);
and U4352 (N_4352,N_278,N_1743);
nor U4353 (N_4353,N_223,N_1029);
nor U4354 (N_4354,N_1106,N_2293);
or U4355 (N_4355,N_680,N_675);
and U4356 (N_4356,N_97,N_1483);
nor U4357 (N_4357,N_2062,N_1739);
and U4358 (N_4358,N_2205,N_2083);
nor U4359 (N_4359,N_143,N_1613);
nor U4360 (N_4360,N_478,N_1915);
nor U4361 (N_4361,N_1046,N_893);
nand U4362 (N_4362,N_692,N_152);
nand U4363 (N_4363,N_1855,N_1884);
nand U4364 (N_4364,N_2082,N_1518);
nand U4365 (N_4365,N_1070,N_721);
and U4366 (N_4366,N_2158,N_2047);
nor U4367 (N_4367,N_2074,N_2086);
or U4368 (N_4368,N_220,N_1952);
nand U4369 (N_4369,N_2311,N_951);
nand U4370 (N_4370,N_1063,N_200);
and U4371 (N_4371,N_54,N_2251);
or U4372 (N_4372,N_331,N_2184);
nor U4373 (N_4373,N_1616,N_1615);
and U4374 (N_4374,N_1304,N_60);
or U4375 (N_4375,N_196,N_625);
or U4376 (N_4376,N_2294,N_514);
nor U4377 (N_4377,N_1744,N_1888);
and U4378 (N_4378,N_2271,N_2247);
and U4379 (N_4379,N_491,N_1271);
or U4380 (N_4380,N_2250,N_2200);
and U4381 (N_4381,N_2281,N_1462);
nor U4382 (N_4382,N_1512,N_472);
or U4383 (N_4383,N_1562,N_351);
nor U4384 (N_4384,N_737,N_65);
nor U4385 (N_4385,N_523,N_584);
or U4386 (N_4386,N_1384,N_590);
nor U4387 (N_4387,N_1124,N_1560);
nand U4388 (N_4388,N_2492,N_1246);
or U4389 (N_4389,N_334,N_996);
or U4390 (N_4390,N_693,N_1630);
and U4391 (N_4391,N_489,N_1084);
nand U4392 (N_4392,N_2433,N_1384);
and U4393 (N_4393,N_64,N_906);
nand U4394 (N_4394,N_620,N_1845);
and U4395 (N_4395,N_1447,N_1984);
or U4396 (N_4396,N_1163,N_77);
nor U4397 (N_4397,N_2053,N_1722);
nand U4398 (N_4398,N_1743,N_2366);
or U4399 (N_4399,N_1747,N_1547);
nor U4400 (N_4400,N_2320,N_1465);
nor U4401 (N_4401,N_401,N_1593);
nand U4402 (N_4402,N_1919,N_199);
nor U4403 (N_4403,N_1107,N_62);
nand U4404 (N_4404,N_97,N_1295);
or U4405 (N_4405,N_1510,N_1592);
or U4406 (N_4406,N_136,N_209);
nand U4407 (N_4407,N_2385,N_1625);
nand U4408 (N_4408,N_2277,N_1893);
and U4409 (N_4409,N_444,N_2276);
nor U4410 (N_4410,N_659,N_1891);
and U4411 (N_4411,N_1796,N_303);
nor U4412 (N_4412,N_844,N_981);
nand U4413 (N_4413,N_2338,N_1773);
nand U4414 (N_4414,N_2302,N_1111);
or U4415 (N_4415,N_2219,N_447);
or U4416 (N_4416,N_1424,N_564);
nand U4417 (N_4417,N_1042,N_112);
nand U4418 (N_4418,N_316,N_890);
nand U4419 (N_4419,N_1189,N_2469);
or U4420 (N_4420,N_1058,N_892);
or U4421 (N_4421,N_76,N_730);
nand U4422 (N_4422,N_1816,N_1519);
or U4423 (N_4423,N_2162,N_992);
nor U4424 (N_4424,N_2473,N_397);
or U4425 (N_4425,N_2419,N_814);
and U4426 (N_4426,N_931,N_319);
or U4427 (N_4427,N_258,N_278);
nand U4428 (N_4428,N_189,N_503);
nand U4429 (N_4429,N_747,N_861);
nand U4430 (N_4430,N_511,N_113);
nand U4431 (N_4431,N_1046,N_1223);
nand U4432 (N_4432,N_363,N_431);
or U4433 (N_4433,N_1441,N_2314);
or U4434 (N_4434,N_549,N_142);
nand U4435 (N_4435,N_1889,N_2395);
nand U4436 (N_4436,N_2399,N_487);
nand U4437 (N_4437,N_1692,N_429);
nand U4438 (N_4438,N_727,N_743);
and U4439 (N_4439,N_1139,N_1836);
or U4440 (N_4440,N_894,N_2418);
or U4441 (N_4441,N_1718,N_814);
xor U4442 (N_4442,N_894,N_1267);
and U4443 (N_4443,N_727,N_472);
and U4444 (N_4444,N_66,N_886);
nand U4445 (N_4445,N_1017,N_2277);
nor U4446 (N_4446,N_806,N_1131);
or U4447 (N_4447,N_1724,N_1338);
and U4448 (N_4448,N_1015,N_20);
nand U4449 (N_4449,N_1445,N_312);
nand U4450 (N_4450,N_1582,N_1571);
or U4451 (N_4451,N_1324,N_1372);
nand U4452 (N_4452,N_31,N_632);
nand U4453 (N_4453,N_1523,N_689);
nor U4454 (N_4454,N_972,N_1463);
and U4455 (N_4455,N_129,N_559);
or U4456 (N_4456,N_2099,N_491);
or U4457 (N_4457,N_1443,N_1782);
nand U4458 (N_4458,N_1177,N_1058);
xnor U4459 (N_4459,N_512,N_1357);
nor U4460 (N_4460,N_1901,N_1572);
nor U4461 (N_4461,N_1464,N_2055);
or U4462 (N_4462,N_831,N_2063);
or U4463 (N_4463,N_913,N_979);
nor U4464 (N_4464,N_666,N_2000);
and U4465 (N_4465,N_856,N_2250);
nor U4466 (N_4466,N_1117,N_319);
nand U4467 (N_4467,N_244,N_1603);
or U4468 (N_4468,N_2252,N_1758);
nor U4469 (N_4469,N_648,N_714);
or U4470 (N_4470,N_426,N_1995);
nand U4471 (N_4471,N_2211,N_1757);
nor U4472 (N_4472,N_1340,N_232);
nand U4473 (N_4473,N_1845,N_616);
or U4474 (N_4474,N_1930,N_1184);
nor U4475 (N_4475,N_1547,N_2401);
or U4476 (N_4476,N_2119,N_1820);
and U4477 (N_4477,N_1640,N_2303);
nor U4478 (N_4478,N_920,N_86);
nand U4479 (N_4479,N_2306,N_163);
or U4480 (N_4480,N_2280,N_1008);
nor U4481 (N_4481,N_1266,N_571);
nand U4482 (N_4482,N_935,N_667);
or U4483 (N_4483,N_336,N_1957);
or U4484 (N_4484,N_2158,N_1944);
or U4485 (N_4485,N_2078,N_2261);
nand U4486 (N_4486,N_832,N_2476);
nand U4487 (N_4487,N_2172,N_2262);
and U4488 (N_4488,N_2087,N_1587);
and U4489 (N_4489,N_1028,N_2471);
nor U4490 (N_4490,N_910,N_829);
or U4491 (N_4491,N_300,N_611);
nand U4492 (N_4492,N_407,N_1823);
nand U4493 (N_4493,N_216,N_204);
nand U4494 (N_4494,N_2405,N_791);
nand U4495 (N_4495,N_880,N_1162);
nand U4496 (N_4496,N_234,N_1675);
nor U4497 (N_4497,N_549,N_297);
nor U4498 (N_4498,N_86,N_1416);
nor U4499 (N_4499,N_2346,N_1606);
and U4500 (N_4500,N_286,N_2427);
and U4501 (N_4501,N_1432,N_340);
or U4502 (N_4502,N_924,N_2278);
and U4503 (N_4503,N_1101,N_22);
and U4504 (N_4504,N_917,N_684);
or U4505 (N_4505,N_1989,N_746);
nand U4506 (N_4506,N_541,N_854);
nor U4507 (N_4507,N_1471,N_2058);
and U4508 (N_4508,N_180,N_2288);
or U4509 (N_4509,N_2430,N_404);
or U4510 (N_4510,N_1280,N_1853);
and U4511 (N_4511,N_841,N_1351);
or U4512 (N_4512,N_1548,N_617);
nand U4513 (N_4513,N_1195,N_1711);
nor U4514 (N_4514,N_612,N_926);
nand U4515 (N_4515,N_2038,N_1541);
nand U4516 (N_4516,N_394,N_1879);
nor U4517 (N_4517,N_2363,N_1180);
nand U4518 (N_4518,N_418,N_724);
nor U4519 (N_4519,N_1709,N_311);
or U4520 (N_4520,N_482,N_410);
or U4521 (N_4521,N_1253,N_1357);
and U4522 (N_4522,N_1189,N_928);
and U4523 (N_4523,N_1821,N_606);
or U4524 (N_4524,N_630,N_475);
nand U4525 (N_4525,N_2275,N_937);
nand U4526 (N_4526,N_791,N_1945);
nor U4527 (N_4527,N_1096,N_1209);
and U4528 (N_4528,N_1670,N_2268);
and U4529 (N_4529,N_1987,N_2410);
nor U4530 (N_4530,N_662,N_2417);
nand U4531 (N_4531,N_1272,N_2344);
nand U4532 (N_4532,N_1961,N_2264);
and U4533 (N_4533,N_245,N_798);
nor U4534 (N_4534,N_1025,N_511);
nor U4535 (N_4535,N_10,N_950);
nand U4536 (N_4536,N_868,N_407);
and U4537 (N_4537,N_2478,N_729);
or U4538 (N_4538,N_1681,N_2162);
or U4539 (N_4539,N_2173,N_2102);
or U4540 (N_4540,N_578,N_1166);
nand U4541 (N_4541,N_375,N_2358);
nor U4542 (N_4542,N_239,N_1089);
or U4543 (N_4543,N_1674,N_30);
nand U4544 (N_4544,N_1877,N_2404);
and U4545 (N_4545,N_508,N_162);
or U4546 (N_4546,N_2078,N_1955);
or U4547 (N_4547,N_750,N_104);
or U4548 (N_4548,N_76,N_731);
and U4549 (N_4549,N_1887,N_2085);
and U4550 (N_4550,N_1801,N_2280);
or U4551 (N_4551,N_607,N_319);
or U4552 (N_4552,N_368,N_1680);
nor U4553 (N_4553,N_1606,N_454);
nor U4554 (N_4554,N_2338,N_1817);
nand U4555 (N_4555,N_1665,N_471);
and U4556 (N_4556,N_711,N_1874);
or U4557 (N_4557,N_2312,N_2223);
nor U4558 (N_4558,N_2316,N_955);
and U4559 (N_4559,N_2238,N_666);
nor U4560 (N_4560,N_1181,N_1362);
nor U4561 (N_4561,N_775,N_877);
and U4562 (N_4562,N_1761,N_1051);
nor U4563 (N_4563,N_959,N_1083);
nor U4564 (N_4564,N_1358,N_1911);
and U4565 (N_4565,N_271,N_907);
nor U4566 (N_4566,N_2440,N_524);
nor U4567 (N_4567,N_1732,N_2291);
or U4568 (N_4568,N_905,N_1455);
and U4569 (N_4569,N_949,N_535);
nor U4570 (N_4570,N_683,N_2304);
nor U4571 (N_4571,N_405,N_998);
or U4572 (N_4572,N_2218,N_1179);
nor U4573 (N_4573,N_2212,N_738);
xor U4574 (N_4574,N_402,N_2396);
and U4575 (N_4575,N_1385,N_2276);
and U4576 (N_4576,N_2000,N_1773);
and U4577 (N_4577,N_338,N_1669);
and U4578 (N_4578,N_1645,N_953);
nand U4579 (N_4579,N_669,N_1734);
or U4580 (N_4580,N_1177,N_2011);
nor U4581 (N_4581,N_1445,N_400);
or U4582 (N_4582,N_2066,N_1295);
nand U4583 (N_4583,N_2182,N_1256);
nor U4584 (N_4584,N_2294,N_792);
or U4585 (N_4585,N_694,N_1896);
nor U4586 (N_4586,N_2308,N_1999);
and U4587 (N_4587,N_431,N_471);
and U4588 (N_4588,N_1016,N_714);
nor U4589 (N_4589,N_1313,N_2237);
and U4590 (N_4590,N_166,N_880);
or U4591 (N_4591,N_776,N_2322);
or U4592 (N_4592,N_2122,N_339);
or U4593 (N_4593,N_1545,N_478);
nor U4594 (N_4594,N_1280,N_1730);
nor U4595 (N_4595,N_359,N_2434);
or U4596 (N_4596,N_2331,N_1523);
or U4597 (N_4597,N_1828,N_1162);
or U4598 (N_4598,N_885,N_279);
nor U4599 (N_4599,N_2399,N_2142);
nand U4600 (N_4600,N_193,N_43);
nor U4601 (N_4601,N_1214,N_2412);
and U4602 (N_4602,N_1377,N_181);
nor U4603 (N_4603,N_387,N_773);
nand U4604 (N_4604,N_1728,N_1732);
nor U4605 (N_4605,N_48,N_1064);
nand U4606 (N_4606,N_353,N_924);
nand U4607 (N_4607,N_2236,N_2088);
nor U4608 (N_4608,N_1709,N_1348);
nand U4609 (N_4609,N_1690,N_2366);
or U4610 (N_4610,N_385,N_2107);
nand U4611 (N_4611,N_1251,N_2153);
or U4612 (N_4612,N_1711,N_898);
and U4613 (N_4613,N_2137,N_2077);
nand U4614 (N_4614,N_1192,N_1601);
or U4615 (N_4615,N_264,N_535);
nand U4616 (N_4616,N_1776,N_1232);
and U4617 (N_4617,N_462,N_93);
nor U4618 (N_4618,N_73,N_1169);
nand U4619 (N_4619,N_1706,N_318);
nand U4620 (N_4620,N_1772,N_88);
nand U4621 (N_4621,N_2005,N_1418);
or U4622 (N_4622,N_1342,N_397);
and U4623 (N_4623,N_843,N_531);
and U4624 (N_4624,N_2195,N_1011);
or U4625 (N_4625,N_483,N_1452);
and U4626 (N_4626,N_578,N_596);
or U4627 (N_4627,N_867,N_2294);
nor U4628 (N_4628,N_1167,N_1783);
nor U4629 (N_4629,N_691,N_1835);
or U4630 (N_4630,N_693,N_1708);
nor U4631 (N_4631,N_1439,N_1714);
nand U4632 (N_4632,N_2403,N_1405);
nand U4633 (N_4633,N_1601,N_822);
nand U4634 (N_4634,N_1993,N_238);
nor U4635 (N_4635,N_3,N_277);
nor U4636 (N_4636,N_1466,N_2361);
nor U4637 (N_4637,N_222,N_278);
xnor U4638 (N_4638,N_881,N_2062);
or U4639 (N_4639,N_998,N_2487);
nor U4640 (N_4640,N_1482,N_474);
nand U4641 (N_4641,N_2360,N_1320);
or U4642 (N_4642,N_2199,N_2142);
nand U4643 (N_4643,N_1656,N_744);
nor U4644 (N_4644,N_857,N_511);
or U4645 (N_4645,N_1534,N_1870);
and U4646 (N_4646,N_1020,N_144);
and U4647 (N_4647,N_410,N_1110);
nand U4648 (N_4648,N_1766,N_344);
nand U4649 (N_4649,N_1310,N_1);
and U4650 (N_4650,N_1744,N_197);
and U4651 (N_4651,N_1506,N_1122);
nand U4652 (N_4652,N_736,N_795);
nand U4653 (N_4653,N_790,N_2052);
or U4654 (N_4654,N_2463,N_1703);
or U4655 (N_4655,N_2130,N_1053);
nor U4656 (N_4656,N_1162,N_1168);
nor U4657 (N_4657,N_662,N_737);
nor U4658 (N_4658,N_1152,N_954);
nor U4659 (N_4659,N_1043,N_284);
and U4660 (N_4660,N_2209,N_2241);
and U4661 (N_4661,N_1204,N_1008);
nand U4662 (N_4662,N_2105,N_2063);
and U4663 (N_4663,N_971,N_1839);
or U4664 (N_4664,N_1178,N_2421);
and U4665 (N_4665,N_1976,N_765);
nand U4666 (N_4666,N_1955,N_2026);
nand U4667 (N_4667,N_631,N_843);
nor U4668 (N_4668,N_1761,N_1604);
nor U4669 (N_4669,N_1067,N_527);
or U4670 (N_4670,N_117,N_2418);
or U4671 (N_4671,N_1478,N_1231);
or U4672 (N_4672,N_1652,N_2038);
nand U4673 (N_4673,N_1689,N_1075);
nand U4674 (N_4674,N_462,N_1230);
and U4675 (N_4675,N_2333,N_625);
nand U4676 (N_4676,N_973,N_526);
nand U4677 (N_4677,N_187,N_2167);
and U4678 (N_4678,N_950,N_2395);
or U4679 (N_4679,N_144,N_2490);
and U4680 (N_4680,N_841,N_2445);
or U4681 (N_4681,N_1011,N_1694);
nand U4682 (N_4682,N_1776,N_663);
or U4683 (N_4683,N_2404,N_463);
nor U4684 (N_4684,N_939,N_1847);
nor U4685 (N_4685,N_489,N_966);
nand U4686 (N_4686,N_393,N_2);
nand U4687 (N_4687,N_1135,N_2285);
and U4688 (N_4688,N_2128,N_1622);
nor U4689 (N_4689,N_2113,N_1343);
and U4690 (N_4690,N_1257,N_1311);
or U4691 (N_4691,N_495,N_1820);
nor U4692 (N_4692,N_268,N_1289);
or U4693 (N_4693,N_2486,N_1143);
nor U4694 (N_4694,N_1330,N_1731);
nor U4695 (N_4695,N_2208,N_2225);
or U4696 (N_4696,N_642,N_534);
nor U4697 (N_4697,N_1719,N_477);
nor U4698 (N_4698,N_2293,N_1840);
nand U4699 (N_4699,N_2313,N_2288);
nand U4700 (N_4700,N_2477,N_1043);
or U4701 (N_4701,N_182,N_1502);
nor U4702 (N_4702,N_333,N_51);
or U4703 (N_4703,N_1372,N_1185);
nand U4704 (N_4704,N_327,N_1442);
nand U4705 (N_4705,N_1538,N_1056);
or U4706 (N_4706,N_2160,N_2087);
or U4707 (N_4707,N_2233,N_1523);
nor U4708 (N_4708,N_1578,N_2447);
nand U4709 (N_4709,N_1446,N_1052);
or U4710 (N_4710,N_2171,N_2002);
nand U4711 (N_4711,N_2115,N_1950);
or U4712 (N_4712,N_359,N_663);
or U4713 (N_4713,N_1664,N_60);
nor U4714 (N_4714,N_752,N_1403);
or U4715 (N_4715,N_1351,N_2469);
nor U4716 (N_4716,N_1768,N_1092);
nand U4717 (N_4717,N_1747,N_1137);
or U4718 (N_4718,N_1999,N_1371);
nand U4719 (N_4719,N_659,N_1583);
and U4720 (N_4720,N_515,N_2258);
nor U4721 (N_4721,N_2327,N_2017);
nand U4722 (N_4722,N_25,N_582);
or U4723 (N_4723,N_2445,N_881);
and U4724 (N_4724,N_1928,N_2073);
or U4725 (N_4725,N_1953,N_1450);
xor U4726 (N_4726,N_1480,N_889);
and U4727 (N_4727,N_802,N_1214);
and U4728 (N_4728,N_322,N_1708);
and U4729 (N_4729,N_1476,N_171);
nor U4730 (N_4730,N_2281,N_23);
nand U4731 (N_4731,N_1483,N_2005);
nand U4732 (N_4732,N_864,N_2297);
or U4733 (N_4733,N_926,N_963);
nor U4734 (N_4734,N_1530,N_1645);
or U4735 (N_4735,N_1275,N_2092);
or U4736 (N_4736,N_1849,N_1645);
nand U4737 (N_4737,N_398,N_104);
or U4738 (N_4738,N_847,N_327);
nand U4739 (N_4739,N_364,N_1399);
nor U4740 (N_4740,N_2262,N_933);
and U4741 (N_4741,N_909,N_1220);
xnor U4742 (N_4742,N_149,N_856);
or U4743 (N_4743,N_1432,N_2120);
and U4744 (N_4744,N_2276,N_1546);
nand U4745 (N_4745,N_325,N_1569);
and U4746 (N_4746,N_2218,N_1131);
nand U4747 (N_4747,N_2183,N_652);
or U4748 (N_4748,N_1977,N_1303);
nor U4749 (N_4749,N_436,N_2418);
nor U4750 (N_4750,N_2051,N_2236);
and U4751 (N_4751,N_1235,N_1773);
or U4752 (N_4752,N_1285,N_299);
or U4753 (N_4753,N_357,N_1063);
or U4754 (N_4754,N_46,N_51);
nor U4755 (N_4755,N_1857,N_1542);
nand U4756 (N_4756,N_1078,N_1200);
and U4757 (N_4757,N_1447,N_1411);
nor U4758 (N_4758,N_936,N_1763);
or U4759 (N_4759,N_1569,N_907);
nand U4760 (N_4760,N_2218,N_1156);
nand U4761 (N_4761,N_1415,N_1375);
and U4762 (N_4762,N_1390,N_346);
and U4763 (N_4763,N_2343,N_1231);
or U4764 (N_4764,N_1934,N_1122);
nand U4765 (N_4765,N_2080,N_928);
nand U4766 (N_4766,N_2388,N_2223);
or U4767 (N_4767,N_254,N_529);
or U4768 (N_4768,N_602,N_904);
nor U4769 (N_4769,N_1537,N_1939);
and U4770 (N_4770,N_1517,N_1289);
nand U4771 (N_4771,N_2336,N_2389);
or U4772 (N_4772,N_484,N_2305);
or U4773 (N_4773,N_383,N_489);
or U4774 (N_4774,N_922,N_1174);
nor U4775 (N_4775,N_1237,N_1935);
nand U4776 (N_4776,N_1218,N_1517);
nor U4777 (N_4777,N_2278,N_1029);
and U4778 (N_4778,N_2401,N_1191);
nor U4779 (N_4779,N_327,N_611);
nand U4780 (N_4780,N_958,N_928);
or U4781 (N_4781,N_1504,N_1611);
nand U4782 (N_4782,N_1979,N_1413);
nand U4783 (N_4783,N_836,N_581);
nand U4784 (N_4784,N_1028,N_727);
nor U4785 (N_4785,N_2189,N_943);
or U4786 (N_4786,N_199,N_1399);
nand U4787 (N_4787,N_1967,N_356);
and U4788 (N_4788,N_1317,N_844);
nor U4789 (N_4789,N_1723,N_1900);
or U4790 (N_4790,N_447,N_4);
nor U4791 (N_4791,N_2420,N_939);
nand U4792 (N_4792,N_1159,N_425);
or U4793 (N_4793,N_1955,N_710);
or U4794 (N_4794,N_15,N_2038);
and U4795 (N_4795,N_2428,N_321);
nand U4796 (N_4796,N_2067,N_2245);
and U4797 (N_4797,N_175,N_227);
and U4798 (N_4798,N_1372,N_1976);
or U4799 (N_4799,N_248,N_2168);
nor U4800 (N_4800,N_1283,N_2491);
nand U4801 (N_4801,N_1809,N_1778);
nor U4802 (N_4802,N_1724,N_1401);
nor U4803 (N_4803,N_1039,N_390);
nor U4804 (N_4804,N_1403,N_2289);
or U4805 (N_4805,N_473,N_2140);
or U4806 (N_4806,N_131,N_305);
nor U4807 (N_4807,N_1106,N_250);
or U4808 (N_4808,N_524,N_187);
and U4809 (N_4809,N_1055,N_1007);
xor U4810 (N_4810,N_1584,N_1423);
and U4811 (N_4811,N_1815,N_925);
nand U4812 (N_4812,N_543,N_689);
and U4813 (N_4813,N_223,N_60);
nand U4814 (N_4814,N_260,N_2115);
or U4815 (N_4815,N_503,N_228);
nand U4816 (N_4816,N_45,N_1590);
nand U4817 (N_4817,N_2412,N_651);
nor U4818 (N_4818,N_277,N_216);
nor U4819 (N_4819,N_1420,N_2361);
nand U4820 (N_4820,N_739,N_929);
nor U4821 (N_4821,N_738,N_2492);
nand U4822 (N_4822,N_2442,N_1981);
nor U4823 (N_4823,N_1406,N_941);
or U4824 (N_4824,N_1297,N_251);
nand U4825 (N_4825,N_2222,N_2004);
and U4826 (N_4826,N_2094,N_933);
nand U4827 (N_4827,N_2260,N_1516);
or U4828 (N_4828,N_464,N_1044);
and U4829 (N_4829,N_205,N_1768);
nand U4830 (N_4830,N_2192,N_523);
nand U4831 (N_4831,N_2124,N_2152);
nor U4832 (N_4832,N_843,N_1037);
and U4833 (N_4833,N_2238,N_840);
nand U4834 (N_4834,N_1669,N_916);
nor U4835 (N_4835,N_144,N_1313);
nand U4836 (N_4836,N_1651,N_751);
or U4837 (N_4837,N_141,N_272);
or U4838 (N_4838,N_1054,N_2067);
or U4839 (N_4839,N_2201,N_955);
and U4840 (N_4840,N_1543,N_2150);
and U4841 (N_4841,N_1455,N_1460);
or U4842 (N_4842,N_353,N_259);
xor U4843 (N_4843,N_672,N_2444);
and U4844 (N_4844,N_1527,N_1338);
nand U4845 (N_4845,N_2403,N_276);
nand U4846 (N_4846,N_2312,N_7);
and U4847 (N_4847,N_128,N_1133);
or U4848 (N_4848,N_796,N_1050);
nand U4849 (N_4849,N_1007,N_1401);
and U4850 (N_4850,N_1522,N_573);
nand U4851 (N_4851,N_2020,N_967);
nor U4852 (N_4852,N_937,N_1111);
nor U4853 (N_4853,N_1490,N_1270);
nand U4854 (N_4854,N_1519,N_697);
or U4855 (N_4855,N_84,N_1520);
and U4856 (N_4856,N_1866,N_907);
nor U4857 (N_4857,N_1881,N_2256);
and U4858 (N_4858,N_1102,N_432);
or U4859 (N_4859,N_2177,N_39);
nor U4860 (N_4860,N_1583,N_1790);
nand U4861 (N_4861,N_1192,N_1574);
nand U4862 (N_4862,N_791,N_1485);
and U4863 (N_4863,N_211,N_1923);
or U4864 (N_4864,N_562,N_1376);
nor U4865 (N_4865,N_680,N_562);
nand U4866 (N_4866,N_1175,N_2193);
or U4867 (N_4867,N_2222,N_1222);
or U4868 (N_4868,N_1323,N_1495);
nand U4869 (N_4869,N_722,N_1533);
and U4870 (N_4870,N_665,N_172);
nor U4871 (N_4871,N_1818,N_2322);
or U4872 (N_4872,N_2094,N_311);
and U4873 (N_4873,N_1005,N_852);
nor U4874 (N_4874,N_1039,N_2379);
nand U4875 (N_4875,N_1216,N_1258);
and U4876 (N_4876,N_307,N_434);
or U4877 (N_4877,N_476,N_428);
nand U4878 (N_4878,N_691,N_55);
or U4879 (N_4879,N_1210,N_1959);
nand U4880 (N_4880,N_615,N_2316);
nor U4881 (N_4881,N_648,N_515);
nand U4882 (N_4882,N_2145,N_1361);
nand U4883 (N_4883,N_2229,N_2255);
nand U4884 (N_4884,N_433,N_1381);
or U4885 (N_4885,N_1335,N_767);
and U4886 (N_4886,N_174,N_597);
nand U4887 (N_4887,N_1717,N_1310);
and U4888 (N_4888,N_1050,N_176);
nor U4889 (N_4889,N_280,N_1481);
nor U4890 (N_4890,N_1527,N_1655);
or U4891 (N_4891,N_835,N_335);
nand U4892 (N_4892,N_723,N_960);
and U4893 (N_4893,N_436,N_861);
nor U4894 (N_4894,N_1916,N_1591);
or U4895 (N_4895,N_2080,N_716);
and U4896 (N_4896,N_4,N_1266);
nor U4897 (N_4897,N_2117,N_1451);
or U4898 (N_4898,N_889,N_2413);
or U4899 (N_4899,N_1617,N_1282);
and U4900 (N_4900,N_813,N_1608);
and U4901 (N_4901,N_99,N_832);
and U4902 (N_4902,N_419,N_1811);
nor U4903 (N_4903,N_1402,N_1291);
and U4904 (N_4904,N_1173,N_1053);
and U4905 (N_4905,N_741,N_2295);
nand U4906 (N_4906,N_1620,N_727);
nand U4907 (N_4907,N_2098,N_677);
nand U4908 (N_4908,N_1004,N_619);
nand U4909 (N_4909,N_1237,N_2103);
or U4910 (N_4910,N_241,N_1779);
nor U4911 (N_4911,N_1328,N_747);
or U4912 (N_4912,N_1095,N_428);
or U4913 (N_4913,N_161,N_501);
or U4914 (N_4914,N_224,N_487);
nor U4915 (N_4915,N_72,N_1157);
nand U4916 (N_4916,N_558,N_1652);
or U4917 (N_4917,N_1106,N_323);
and U4918 (N_4918,N_1889,N_1199);
or U4919 (N_4919,N_1772,N_1269);
or U4920 (N_4920,N_1422,N_1483);
and U4921 (N_4921,N_1013,N_857);
nor U4922 (N_4922,N_485,N_1615);
nand U4923 (N_4923,N_1122,N_1601);
nor U4924 (N_4924,N_1940,N_1192);
nand U4925 (N_4925,N_1852,N_1757);
and U4926 (N_4926,N_485,N_628);
nor U4927 (N_4927,N_1954,N_2455);
nor U4928 (N_4928,N_847,N_1668);
nor U4929 (N_4929,N_223,N_272);
nor U4930 (N_4930,N_2434,N_252);
nor U4931 (N_4931,N_1883,N_1621);
nor U4932 (N_4932,N_137,N_97);
or U4933 (N_4933,N_263,N_122);
and U4934 (N_4934,N_1490,N_493);
or U4935 (N_4935,N_271,N_962);
nor U4936 (N_4936,N_1040,N_1382);
and U4937 (N_4937,N_858,N_2024);
and U4938 (N_4938,N_1988,N_39);
and U4939 (N_4939,N_2009,N_2398);
or U4940 (N_4940,N_184,N_1668);
and U4941 (N_4941,N_690,N_1659);
and U4942 (N_4942,N_1605,N_1241);
nand U4943 (N_4943,N_2041,N_1234);
nor U4944 (N_4944,N_1010,N_1719);
and U4945 (N_4945,N_1292,N_14);
nor U4946 (N_4946,N_1706,N_2092);
and U4947 (N_4947,N_832,N_2455);
nor U4948 (N_4948,N_668,N_465);
nand U4949 (N_4949,N_2362,N_906);
nand U4950 (N_4950,N_1468,N_2330);
and U4951 (N_4951,N_264,N_837);
or U4952 (N_4952,N_2389,N_1193);
nor U4953 (N_4953,N_714,N_220);
nand U4954 (N_4954,N_1575,N_2289);
nor U4955 (N_4955,N_1166,N_200);
nor U4956 (N_4956,N_1895,N_777);
or U4957 (N_4957,N_240,N_1105);
and U4958 (N_4958,N_1079,N_25);
and U4959 (N_4959,N_1034,N_1814);
nor U4960 (N_4960,N_606,N_1816);
or U4961 (N_4961,N_272,N_2156);
nand U4962 (N_4962,N_812,N_1837);
nand U4963 (N_4963,N_1619,N_2387);
nand U4964 (N_4964,N_2392,N_1802);
or U4965 (N_4965,N_2438,N_594);
or U4966 (N_4966,N_1265,N_1751);
or U4967 (N_4967,N_2274,N_1255);
and U4968 (N_4968,N_1039,N_1531);
nand U4969 (N_4969,N_1114,N_15);
or U4970 (N_4970,N_2036,N_1185);
or U4971 (N_4971,N_2034,N_1446);
nor U4972 (N_4972,N_1086,N_1548);
nand U4973 (N_4973,N_2023,N_1799);
nor U4974 (N_4974,N_1658,N_2492);
or U4975 (N_4975,N_1341,N_669);
nand U4976 (N_4976,N_1813,N_1292);
or U4977 (N_4977,N_1249,N_209);
nor U4978 (N_4978,N_929,N_1112);
or U4979 (N_4979,N_95,N_2476);
nor U4980 (N_4980,N_653,N_2428);
nor U4981 (N_4981,N_426,N_1311);
nand U4982 (N_4982,N_1624,N_689);
nor U4983 (N_4983,N_1233,N_2305);
nand U4984 (N_4984,N_853,N_1175);
or U4985 (N_4985,N_1161,N_1070);
and U4986 (N_4986,N_1396,N_1408);
and U4987 (N_4987,N_224,N_1651);
and U4988 (N_4988,N_606,N_1023);
or U4989 (N_4989,N_2442,N_1750);
nor U4990 (N_4990,N_2231,N_216);
xnor U4991 (N_4991,N_672,N_1486);
nand U4992 (N_4992,N_1465,N_491);
or U4993 (N_4993,N_1811,N_451);
or U4994 (N_4994,N_537,N_487);
or U4995 (N_4995,N_1636,N_2290);
or U4996 (N_4996,N_2463,N_1931);
nand U4997 (N_4997,N_1941,N_1693);
and U4998 (N_4998,N_2200,N_2065);
and U4999 (N_4999,N_2033,N_622);
nor U5000 (N_5000,N_3331,N_4278);
or U5001 (N_5001,N_3802,N_2695);
nor U5002 (N_5002,N_4191,N_4035);
nand U5003 (N_5003,N_3966,N_4720);
or U5004 (N_5004,N_4598,N_2805);
nand U5005 (N_5005,N_4784,N_3516);
nor U5006 (N_5006,N_2691,N_2553);
or U5007 (N_5007,N_2956,N_4241);
or U5008 (N_5008,N_4971,N_3911);
or U5009 (N_5009,N_2779,N_2617);
or U5010 (N_5010,N_3017,N_4815);
and U5011 (N_5011,N_2751,N_3361);
nor U5012 (N_5012,N_4381,N_2801);
and U5013 (N_5013,N_4669,N_4458);
or U5014 (N_5014,N_4510,N_2628);
nor U5015 (N_5015,N_3836,N_4385);
and U5016 (N_5016,N_4781,N_4681);
nor U5017 (N_5017,N_3565,N_3750);
nor U5018 (N_5018,N_4963,N_3968);
or U5019 (N_5019,N_3106,N_3265);
and U5020 (N_5020,N_4700,N_4026);
nand U5021 (N_5021,N_4183,N_4780);
nor U5022 (N_5022,N_4198,N_2931);
or U5023 (N_5023,N_3125,N_3528);
or U5024 (N_5024,N_3792,N_3041);
xnor U5025 (N_5025,N_4133,N_3057);
and U5026 (N_5026,N_3897,N_4264);
or U5027 (N_5027,N_3891,N_4379);
or U5028 (N_5028,N_4178,N_3138);
and U5029 (N_5029,N_4674,N_4365);
nor U5030 (N_5030,N_3373,N_3590);
and U5031 (N_5031,N_4748,N_3163);
and U5032 (N_5032,N_3408,N_4473);
and U5033 (N_5033,N_4616,N_3292);
and U5034 (N_5034,N_2888,N_3922);
nand U5035 (N_5035,N_3886,N_4369);
and U5036 (N_5036,N_3845,N_2596);
and U5037 (N_5037,N_2775,N_3183);
or U5038 (N_5038,N_4668,N_2761);
nand U5039 (N_5039,N_3915,N_4362);
nand U5040 (N_5040,N_3664,N_3986);
nor U5041 (N_5041,N_3320,N_3753);
nand U5042 (N_5042,N_4307,N_3152);
or U5043 (N_5043,N_4130,N_3964);
or U5044 (N_5044,N_3522,N_2788);
or U5045 (N_5045,N_4829,N_4097);
nand U5046 (N_5046,N_2750,N_3839);
or U5047 (N_5047,N_2627,N_3310);
nor U5048 (N_5048,N_2629,N_2702);
or U5049 (N_5049,N_3427,N_2744);
nor U5050 (N_5050,N_4931,N_4934);
nand U5051 (N_5051,N_2656,N_2684);
xor U5052 (N_5052,N_4438,N_2624);
or U5053 (N_5053,N_4476,N_3712);
or U5054 (N_5054,N_3296,N_3413);
nand U5055 (N_5055,N_4922,N_4747);
nand U5056 (N_5056,N_3527,N_3114);
nand U5057 (N_5057,N_3141,N_3688);
xor U5058 (N_5058,N_4749,N_4865);
nand U5059 (N_5059,N_3757,N_4965);
nor U5060 (N_5060,N_4347,N_4452);
nand U5061 (N_5061,N_2698,N_3488);
xnor U5062 (N_5062,N_3953,N_3875);
or U5063 (N_5063,N_3404,N_4111);
nor U5064 (N_5064,N_4515,N_3094);
or U5065 (N_5065,N_2918,N_2559);
nand U5066 (N_5066,N_4550,N_3020);
and U5067 (N_5067,N_4481,N_3500);
or U5068 (N_5068,N_4858,N_3949);
nand U5069 (N_5069,N_3301,N_2982);
nand U5070 (N_5070,N_4479,N_4275);
nor U5071 (N_5071,N_4165,N_2643);
nor U5072 (N_5072,N_4132,N_2570);
and U5073 (N_5073,N_3594,N_4454);
and U5074 (N_5074,N_4055,N_4078);
or U5075 (N_5075,N_4779,N_4057);
or U5076 (N_5076,N_3402,N_3199);
and U5077 (N_5077,N_3606,N_3666);
nand U5078 (N_5078,N_4228,N_4527);
nand U5079 (N_5079,N_3696,N_3126);
nand U5080 (N_5080,N_4041,N_4734);
and U5081 (N_5081,N_3015,N_2590);
or U5082 (N_5082,N_4764,N_4936);
nand U5083 (N_5083,N_3720,N_3066);
nor U5084 (N_5084,N_4214,N_4786);
or U5085 (N_5085,N_3054,N_2675);
or U5086 (N_5086,N_4575,N_3476);
nand U5087 (N_5087,N_4290,N_2708);
or U5088 (N_5088,N_3730,N_3214);
nor U5089 (N_5089,N_3190,N_4870);
nor U5090 (N_5090,N_4868,N_4951);
nor U5091 (N_5091,N_4488,N_3904);
and U5092 (N_5092,N_4155,N_4617);
nor U5093 (N_5093,N_2520,N_2631);
and U5094 (N_5094,N_3863,N_4195);
nand U5095 (N_5095,N_4088,N_4698);
and U5096 (N_5096,N_4895,N_4845);
nand U5097 (N_5097,N_4728,N_2842);
nand U5098 (N_5098,N_4832,N_4590);
or U5099 (N_5099,N_4554,N_2641);
and U5100 (N_5100,N_4975,N_3317);
or U5101 (N_5101,N_4619,N_4478);
nand U5102 (N_5102,N_4382,N_4083);
nor U5103 (N_5103,N_4713,N_3458);
nor U5104 (N_5104,N_3139,N_4240);
nand U5105 (N_5105,N_3110,N_4467);
and U5106 (N_5106,N_3959,N_3080);
nand U5107 (N_5107,N_4830,N_2604);
nand U5108 (N_5108,N_2839,N_2968);
or U5109 (N_5109,N_4653,N_3780);
and U5110 (N_5110,N_3625,N_4059);
nand U5111 (N_5111,N_4937,N_4269);
and U5112 (N_5112,N_2734,N_4646);
nor U5113 (N_5113,N_2940,N_2996);
or U5114 (N_5114,N_3702,N_4735);
nor U5115 (N_5115,N_3943,N_4732);
and U5116 (N_5116,N_3001,N_4631);
nor U5117 (N_5117,N_4533,N_3853);
or U5118 (N_5118,N_2546,N_4042);
nor U5119 (N_5119,N_3651,N_4577);
nand U5120 (N_5120,N_3832,N_4933);
or U5121 (N_5121,N_4945,N_3890);
nand U5122 (N_5122,N_4657,N_2738);
or U5123 (N_5123,N_4346,N_3652);
nor U5124 (N_5124,N_3266,N_4153);
and U5125 (N_5125,N_4691,N_4246);
nor U5126 (N_5126,N_3771,N_4265);
and U5127 (N_5127,N_3867,N_4463);
and U5128 (N_5128,N_4798,N_3555);
nand U5129 (N_5129,N_2605,N_4303);
nor U5130 (N_5130,N_4816,N_3703);
or U5131 (N_5131,N_4163,N_3604);
nand U5132 (N_5132,N_3043,N_3831);
nand U5133 (N_5133,N_2938,N_4885);
nand U5134 (N_5134,N_3866,N_3270);
or U5135 (N_5135,N_4518,N_3396);
or U5136 (N_5136,N_3686,N_4243);
and U5137 (N_5137,N_4753,N_4604);
or U5138 (N_5138,N_3465,N_4536);
or U5139 (N_5139,N_3460,N_4161);
nand U5140 (N_5140,N_4245,N_4392);
and U5141 (N_5141,N_3036,N_4710);
and U5142 (N_5142,N_2509,N_3777);
and U5143 (N_5143,N_4609,N_4349);
and U5144 (N_5144,N_2531,N_2609);
and U5145 (N_5145,N_3477,N_4840);
nor U5146 (N_5146,N_4082,N_4677);
and U5147 (N_5147,N_4876,N_3807);
nor U5148 (N_5148,N_3992,N_3400);
or U5149 (N_5149,N_2522,N_4799);
nor U5150 (N_5150,N_4750,N_3096);
nand U5151 (N_5151,N_3805,N_4216);
nand U5152 (N_5152,N_2655,N_3000);
and U5153 (N_5153,N_3646,N_2715);
nor U5154 (N_5154,N_4549,N_4137);
nand U5155 (N_5155,N_4022,N_2584);
nor U5156 (N_5156,N_4139,N_4149);
or U5157 (N_5157,N_3142,N_4109);
and U5158 (N_5158,N_4135,N_3228);
and U5159 (N_5159,N_4557,N_4172);
and U5160 (N_5160,N_4623,N_3473);
nand U5161 (N_5161,N_2731,N_3305);
or U5162 (N_5162,N_4356,N_3491);
nor U5163 (N_5163,N_3165,N_3362);
and U5164 (N_5164,N_4642,N_3207);
nand U5165 (N_5165,N_4571,N_3583);
nand U5166 (N_5166,N_3678,N_4996);
and U5167 (N_5167,N_4225,N_3613);
and U5168 (N_5168,N_4875,N_4411);
nor U5169 (N_5169,N_3668,N_2828);
and U5170 (N_5170,N_3605,N_2713);
nor U5171 (N_5171,N_3737,N_4008);
and U5172 (N_5172,N_4974,N_4414);
nand U5173 (N_5173,N_3193,N_3562);
nor U5174 (N_5174,N_4923,N_3963);
nor U5175 (N_5175,N_4866,N_2814);
nor U5176 (N_5176,N_3916,N_2957);
or U5177 (N_5177,N_3436,N_3632);
and U5178 (N_5178,N_2662,N_3821);
nand U5179 (N_5179,N_4138,N_2625);
nor U5180 (N_5180,N_4917,N_3541);
and U5181 (N_5181,N_2985,N_2860);
and U5182 (N_5182,N_4304,N_4867);
nand U5183 (N_5183,N_4390,N_3761);
or U5184 (N_5184,N_3824,N_4158);
nor U5185 (N_5185,N_4104,N_2886);
nor U5186 (N_5186,N_4474,N_3573);
nand U5187 (N_5187,N_4625,N_4632);
and U5188 (N_5188,N_2883,N_2780);
nand U5189 (N_5189,N_4920,N_3869);
and U5190 (N_5190,N_2733,N_4806);
nand U5191 (N_5191,N_3425,N_4233);
nand U5192 (N_5192,N_3294,N_3468);
nor U5193 (N_5193,N_3628,N_4511);
or U5194 (N_5194,N_4256,N_4320);
or U5195 (N_5195,N_3826,N_2526);
and U5196 (N_5196,N_4864,N_3903);
or U5197 (N_5197,N_2567,N_3731);
or U5198 (N_5198,N_3439,N_4020);
or U5199 (N_5199,N_3850,N_3449);
and U5200 (N_5200,N_3407,N_3459);
nand U5201 (N_5201,N_4767,N_3336);
and U5202 (N_5202,N_4206,N_4108);
and U5203 (N_5203,N_4095,N_3797);
and U5204 (N_5204,N_3254,N_3622);
or U5205 (N_5205,N_4475,N_4589);
and U5206 (N_5206,N_4599,N_4812);
or U5207 (N_5207,N_4859,N_2554);
nor U5208 (N_5208,N_4721,N_2549);
and U5209 (N_5209,N_3976,N_2669);
xnor U5210 (N_5210,N_4074,N_4400);
xnor U5211 (N_5211,N_2992,N_4558);
nand U5212 (N_5212,N_2727,N_2569);
nor U5213 (N_5213,N_4449,N_3578);
and U5214 (N_5214,N_3470,N_3834);
or U5215 (N_5215,N_3290,N_3596);
nand U5216 (N_5216,N_3506,N_3258);
xnor U5217 (N_5217,N_3155,N_4730);
and U5218 (N_5218,N_3127,N_2634);
or U5219 (N_5219,N_4384,N_3655);
and U5220 (N_5220,N_4402,N_4368);
nor U5221 (N_5221,N_3377,N_3406);
and U5222 (N_5222,N_3929,N_3558);
xor U5223 (N_5223,N_4719,N_2545);
nand U5224 (N_5224,N_3372,N_3205);
and U5225 (N_5225,N_4424,N_4912);
nor U5226 (N_5226,N_2706,N_3711);
and U5227 (N_5227,N_2615,N_2626);
and U5228 (N_5228,N_3116,N_4938);
nand U5229 (N_5229,N_2762,N_3092);
or U5230 (N_5230,N_3724,N_4224);
nor U5231 (N_5231,N_4089,N_4982);
or U5232 (N_5232,N_4101,N_3859);
nor U5233 (N_5233,N_3243,N_4699);
and U5234 (N_5234,N_4763,N_4039);
and U5235 (N_5235,N_4027,N_2885);
nand U5236 (N_5236,N_3184,N_3539);
or U5237 (N_5237,N_4964,N_3932);
or U5238 (N_5238,N_4879,N_4497);
and U5239 (N_5239,N_4582,N_4021);
and U5240 (N_5240,N_3283,N_4373);
nand U5241 (N_5241,N_3739,N_4120);
nor U5242 (N_5242,N_3151,N_2867);
or U5243 (N_5243,N_4236,N_4501);
and U5244 (N_5244,N_2873,N_2671);
and U5245 (N_5245,N_4546,N_3879);
and U5246 (N_5246,N_4237,N_4493);
and U5247 (N_5247,N_2840,N_4523);
or U5248 (N_5248,N_4338,N_4796);
or U5249 (N_5249,N_3638,N_4890);
nor U5250 (N_5250,N_4555,N_3050);
nor U5251 (N_5251,N_3658,N_4926);
and U5252 (N_5252,N_3412,N_3671);
or U5253 (N_5253,N_2673,N_3872);
nor U5254 (N_5254,N_3769,N_4913);
or U5255 (N_5255,N_4628,N_4988);
or U5256 (N_5256,N_3849,N_4134);
nor U5257 (N_5257,N_4073,N_4976);
and U5258 (N_5258,N_4332,N_3572);
and U5259 (N_5259,N_3918,N_2682);
and U5260 (N_5260,N_4871,N_4387);
nand U5261 (N_5261,N_4239,N_2786);
and U5262 (N_5262,N_2862,N_2757);
or U5263 (N_5263,N_3004,N_3800);
and U5264 (N_5264,N_4408,N_2517);
and U5265 (N_5265,N_4655,N_4397);
and U5266 (N_5266,N_3942,N_4298);
nand U5267 (N_5267,N_3038,N_4521);
nor U5268 (N_5268,N_4308,N_3715);
and U5269 (N_5269,N_3551,N_3593);
nand U5270 (N_5270,N_4560,N_4086);
and U5271 (N_5271,N_4855,N_2991);
nand U5272 (N_5272,N_4319,N_4260);
and U5273 (N_5273,N_3157,N_3028);
and U5274 (N_5274,N_2848,N_3765);
or U5275 (N_5275,N_3740,N_3670);
or U5276 (N_5276,N_2776,N_4645);
or U5277 (N_5277,N_2793,N_3095);
xor U5278 (N_5278,N_4189,N_2932);
or U5279 (N_5279,N_2893,N_4990);
nor U5280 (N_5280,N_2622,N_4650);
and U5281 (N_5281,N_3383,N_3612);
and U5282 (N_5282,N_3549,N_4363);
and U5283 (N_5283,N_3014,N_3371);
and U5284 (N_5284,N_2723,N_3498);
and U5285 (N_5285,N_2610,N_2777);
and U5286 (N_5286,N_4266,N_2965);
nand U5287 (N_5287,N_4722,N_3816);
nor U5288 (N_5288,N_2937,N_2829);
nor U5289 (N_5289,N_3128,N_3033);
and U5290 (N_5290,N_3926,N_4181);
nand U5291 (N_5291,N_2753,N_3692);
and U5292 (N_5292,N_4462,N_4306);
or U5293 (N_5293,N_3502,N_3431);
nor U5294 (N_5294,N_3405,N_2635);
or U5295 (N_5295,N_3923,N_4099);
nor U5296 (N_5296,N_3277,N_2581);
and U5297 (N_5297,N_4383,N_3817);
or U5298 (N_5298,N_4957,N_2688);
or U5299 (N_5299,N_3636,N_3617);
nor U5300 (N_5300,N_2623,N_3677);
nand U5301 (N_5301,N_3087,N_2606);
and U5302 (N_5302,N_4037,N_4643);
nor U5303 (N_5303,N_3230,N_3443);
or U5304 (N_5304,N_3961,N_3812);
nand U5305 (N_5305,N_3211,N_3830);
and U5306 (N_5306,N_2863,N_3643);
and U5307 (N_5307,N_2905,N_4826);
or U5308 (N_5308,N_4828,N_4354);
or U5309 (N_5309,N_4440,N_4552);
nor U5310 (N_5310,N_3453,N_3563);
nor U5311 (N_5311,N_4234,N_3418);
xnor U5312 (N_5312,N_3735,N_4076);
or U5313 (N_5313,N_4238,N_2974);
nand U5314 (N_5314,N_4118,N_4066);
or U5315 (N_5315,N_2525,N_4192);
nand U5316 (N_5316,N_4268,N_2571);
and U5317 (N_5317,N_3888,N_4831);
nor U5318 (N_5318,N_3180,N_3415);
and U5319 (N_5319,N_4051,N_2815);
or U5320 (N_5320,N_3798,N_2797);
or U5321 (N_5321,N_2592,N_3181);
nor U5322 (N_5322,N_4814,N_4640);
nand U5323 (N_5323,N_4935,N_2557);
or U5324 (N_5324,N_3838,N_3168);
nor U5325 (N_5325,N_3073,N_3469);
nand U5326 (N_5326,N_3284,N_3633);
and U5327 (N_5327,N_2972,N_3329);
and U5328 (N_5328,N_2701,N_3321);
and U5329 (N_5329,N_3068,N_2999);
and U5330 (N_5330,N_3945,N_4348);
xnor U5331 (N_5331,N_3389,N_4091);
nand U5332 (N_5332,N_4407,N_3162);
nand U5333 (N_5333,N_3238,N_4904);
or U5334 (N_5334,N_3602,N_3006);
nor U5335 (N_5335,N_4992,N_3393);
or U5336 (N_5336,N_3382,N_4084);
nand U5337 (N_5337,N_3704,N_2506);
or U5338 (N_5338,N_2948,N_3881);
xnor U5339 (N_5339,N_4248,N_4952);
and U5340 (N_5340,N_4342,N_3182);
and U5341 (N_5341,N_4803,N_3280);
nor U5342 (N_5342,N_4393,N_2687);
and U5343 (N_5343,N_2789,N_3454);
nand U5344 (N_5344,N_3889,N_2954);
nor U5345 (N_5345,N_4100,N_3176);
nand U5346 (N_5346,N_4466,N_4991);
and U5347 (N_5347,N_4092,N_3084);
nor U5348 (N_5348,N_3525,N_4105);
or U5349 (N_5349,N_2952,N_4662);
or U5350 (N_5350,N_3360,N_3591);
nor U5351 (N_5351,N_3755,N_4649);
or U5352 (N_5352,N_4607,N_3718);
and U5353 (N_5353,N_3260,N_2650);
or U5354 (N_5354,N_4002,N_4514);
nor U5355 (N_5355,N_3510,N_4726);
nand U5356 (N_5356,N_4124,N_3137);
nor U5357 (N_5357,N_2544,N_4615);
and U5358 (N_5358,N_3356,N_3131);
and U5359 (N_5359,N_4883,N_4334);
and U5360 (N_5360,N_4359,N_4053);
nor U5361 (N_5361,N_3399,N_4289);
nand U5362 (N_5362,N_2647,N_2690);
nand U5363 (N_5363,N_3917,N_4716);
and U5364 (N_5364,N_2737,N_4014);
nor U5365 (N_5365,N_3883,N_3973);
and U5366 (N_5366,N_3642,N_2804);
or U5367 (N_5367,N_4046,N_4597);
and U5368 (N_5368,N_3363,N_3354);
xor U5369 (N_5369,N_3895,N_4506);
and U5370 (N_5370,N_2812,N_2568);
or U5371 (N_5371,N_3056,N_2927);
nor U5372 (N_5372,N_3269,N_3315);
nor U5373 (N_5373,N_3093,N_2836);
nand U5374 (N_5374,N_4672,N_3010);
nor U5375 (N_5375,N_2746,N_4503);
and U5376 (N_5376,N_4851,N_3620);
nand U5377 (N_5377,N_4955,N_2660);
nor U5378 (N_5378,N_3936,N_2740);
and U5379 (N_5379,N_4353,N_2664);
nor U5380 (N_5380,N_2551,N_3191);
nand U5381 (N_5381,N_3312,N_4223);
nand U5382 (N_5382,N_2646,N_4603);
nor U5383 (N_5383,N_3723,N_3451);
nor U5384 (N_5384,N_3219,N_4659);
or U5385 (N_5385,N_4184,N_4508);
nor U5386 (N_5386,N_3414,N_4509);
nand U5387 (N_5387,N_2849,N_2979);
or U5388 (N_5388,N_3592,N_4333);
nand U5389 (N_5389,N_3115,N_3774);
or U5390 (N_5390,N_3878,N_2649);
nor U5391 (N_5391,N_3263,N_3101);
nor U5392 (N_5392,N_4556,N_4929);
nand U5393 (N_5393,N_3107,N_3367);
and U5394 (N_5394,N_4434,N_4707);
and U5395 (N_5395,N_3421,N_4244);
nor U5396 (N_5396,N_4112,N_3385);
and U5397 (N_5397,N_2847,N_3055);
nand U5398 (N_5398,N_2816,N_3603);
nand U5399 (N_5399,N_3504,N_2935);
nor U5400 (N_5400,N_3120,N_3744);
nand U5401 (N_5401,N_3540,N_3351);
nand U5402 (N_5402,N_4056,N_3983);
or U5403 (N_5403,N_3278,N_3341);
or U5404 (N_5404,N_4924,N_4459);
nor U5405 (N_5405,N_3687,N_4778);
nor U5406 (N_5406,N_3854,N_3577);
or U5407 (N_5407,N_4854,N_3833);
nor U5408 (N_5408,N_3585,N_3919);
and U5409 (N_5409,N_4811,N_2644);
or U5410 (N_5410,N_3870,N_4512);
nor U5411 (N_5411,N_4441,N_4877);
and U5412 (N_5412,N_2966,N_2859);
nor U5413 (N_5413,N_2897,N_3040);
and U5414 (N_5414,N_4154,N_3884);
or U5415 (N_5415,N_3322,N_2722);
xnor U5416 (N_5416,N_4760,N_2721);
and U5417 (N_5417,N_3194,N_3700);
nand U5418 (N_5418,N_3795,N_3218);
and U5419 (N_5419,N_4094,N_3524);
nand U5420 (N_5420,N_4921,N_2855);
nand U5421 (N_5421,N_4959,N_4067);
nor U5422 (N_5422,N_3898,N_3318);
nand U5423 (N_5423,N_4121,N_4071);
nor U5424 (N_5424,N_3342,N_2679);
or U5425 (N_5425,N_4351,N_4213);
and U5426 (N_5426,N_4993,N_3829);
nor U5427 (N_5427,N_4998,N_2705);
nor U5428 (N_5428,N_3257,N_4916);
nor U5429 (N_5429,N_3991,N_3693);
and U5430 (N_5430,N_3289,N_3996);
or U5431 (N_5431,N_4257,N_3815);
nor U5432 (N_5432,N_2958,N_3995);
or U5433 (N_5433,N_2959,N_2826);
nand U5434 (N_5434,N_3464,N_3801);
and U5435 (N_5435,N_3308,N_2600);
xnor U5436 (N_5436,N_3698,N_2668);
and U5437 (N_5437,N_3426,N_4423);
and U5438 (N_5438,N_3158,N_3071);
nor U5439 (N_5439,N_2739,N_2764);
or U5440 (N_5440,N_3235,N_3272);
nand U5441 (N_5441,N_3287,N_3104);
nor U5442 (N_5442,N_2730,N_2541);
nor U5443 (N_5443,N_4682,N_3791);
or U5444 (N_5444,N_3175,N_3103);
nor U5445 (N_5445,N_2798,N_3143);
nand U5446 (N_5446,N_3375,N_3988);
nand U5447 (N_5447,N_4480,N_3249);
and U5448 (N_5448,N_2936,N_4773);
nand U5449 (N_5449,N_3660,N_3629);
nand U5450 (N_5450,N_4939,N_4807);
or U5451 (N_5451,N_4667,N_3031);
nor U5452 (N_5452,N_4435,N_3734);
nand U5453 (N_5453,N_3448,N_3124);
nand U5454 (N_5454,N_3999,N_4167);
and U5455 (N_5455,N_4850,N_4302);
nor U5456 (N_5456,N_3980,N_2983);
nand U5457 (N_5457,N_2903,N_3144);
and U5458 (N_5458,N_4507,N_3259);
or U5459 (N_5459,N_2939,N_3417);
and U5460 (N_5460,N_2768,N_3848);
and U5461 (N_5461,N_4502,N_3647);
nor U5462 (N_5462,N_2852,N_2736);
or U5463 (N_5463,N_3164,N_4562);
or U5464 (N_5464,N_3857,N_2790);
nand U5465 (N_5465,N_3754,N_4277);
nand U5466 (N_5466,N_4455,N_2833);
or U5467 (N_5467,N_4862,N_2864);
and U5468 (N_5468,N_3552,N_3669);
and U5469 (N_5469,N_2621,N_4419);
nor U5470 (N_5470,N_3275,N_4412);
or U5471 (N_5471,N_4326,N_3948);
nor U5472 (N_5472,N_3333,N_4622);
nor U5473 (N_5473,N_3167,N_4430);
or U5474 (N_5474,N_3865,N_4910);
nor U5475 (N_5475,N_3195,N_4606);
nor U5476 (N_5476,N_3352,N_2533);
or U5477 (N_5477,N_3083,N_2562);
nor U5478 (N_5478,N_2585,N_3580);
nor U5479 (N_5479,N_3546,N_4313);
or U5480 (N_5480,N_4340,N_4420);
and U5481 (N_5481,N_4309,N_4752);
nor U5482 (N_5482,N_3529,N_3295);
or U5483 (N_5483,N_2763,N_3298);
or U5484 (N_5484,N_3847,N_3098);
or U5485 (N_5485,N_4162,N_4633);
or U5486 (N_5486,N_4834,N_3785);
xnor U5487 (N_5487,N_3672,N_2795);
nor U5488 (N_5488,N_4274,N_2637);
nor U5489 (N_5489,N_3256,N_4563);
nand U5490 (N_5490,N_4495,N_4499);
nor U5491 (N_5491,N_2575,N_3334);
nor U5492 (N_5492,N_4583,N_2534);
and U5493 (N_5493,N_3044,N_2854);
nor U5494 (N_5494,N_3571,N_3570);
and U5495 (N_5495,N_3481,N_4925);
nor U5496 (N_5496,N_3483,N_3062);
nor U5497 (N_5497,N_3099,N_4946);
nand U5498 (N_5498,N_4572,N_3749);
or U5499 (N_5499,N_3457,N_3022);
xnor U5500 (N_5500,N_3485,N_4001);
nand U5501 (N_5501,N_4727,N_3683);
or U5502 (N_5502,N_4352,N_3088);
or U5503 (N_5503,N_4838,N_3746);
nand U5504 (N_5504,N_3011,N_4000);
nand U5505 (N_5505,N_3077,N_3349);
or U5506 (N_5506,N_3306,N_2603);
or U5507 (N_5507,N_3021,N_2718);
nand U5508 (N_5508,N_4788,N_3751);
nor U5509 (N_5509,N_4003,N_4742);
nor U5510 (N_5510,N_3689,N_3132);
nor U5511 (N_5511,N_3216,N_4894);
xnor U5512 (N_5512,N_2941,N_2728);
and U5513 (N_5513,N_2891,N_2765);
nand U5514 (N_5514,N_3912,N_3150);
nor U5515 (N_5515,N_4882,N_4310);
and U5516 (N_5516,N_2875,N_4596);
nand U5517 (N_5517,N_4335,N_4187);
or U5518 (N_5518,N_4697,N_4884);
and U5519 (N_5519,N_4398,N_3928);
and U5520 (N_5520,N_3496,N_4116);
or U5521 (N_5521,N_3337,N_3039);
nor U5522 (N_5522,N_3741,N_4947);
or U5523 (N_5523,N_3113,N_2537);
nand U5524 (N_5524,N_4034,N_3224);
nand U5525 (N_5525,N_3378,N_3907);
and U5526 (N_5526,N_3058,N_3111);
and U5527 (N_5527,N_3433,N_2880);
nor U5528 (N_5528,N_4415,N_3047);
nor U5529 (N_5529,N_3819,N_3611);
nand U5530 (N_5530,N_3411,N_4341);
or U5531 (N_5531,N_4418,N_2505);
and U5532 (N_5532,N_2946,N_3630);
nor U5533 (N_5533,N_3745,N_4860);
nor U5534 (N_5534,N_4427,N_3474);
and U5535 (N_5535,N_4566,N_4374);
and U5536 (N_5536,N_2699,N_4775);
or U5537 (N_5537,N_3575,N_2747);
and U5538 (N_5538,N_2619,N_3758);
nand U5539 (N_5539,N_4712,N_3925);
and U5540 (N_5540,N_4787,N_2703);
and U5541 (N_5541,N_2792,N_3582);
nand U5542 (N_5542,N_3856,N_4209);
nor U5543 (N_5543,N_3533,N_4644);
nor U5544 (N_5544,N_4956,N_4725);
or U5545 (N_5545,N_2672,N_4821);
nor U5546 (N_5546,N_4594,N_4872);
and U5547 (N_5547,N_3763,N_4437);
nor U5548 (N_5548,N_3067,N_2841);
nand U5549 (N_5549,N_4123,N_3788);
and U5550 (N_5550,N_3186,N_3121);
and U5551 (N_5551,N_4018,N_3429);
nor U5552 (N_5552,N_2856,N_2922);
nand U5553 (N_5553,N_4090,N_4177);
and U5554 (N_5554,N_3392,N_4805);
or U5555 (N_5555,N_4680,N_2561);
or U5556 (N_5556,N_3676,N_4410);
or U5557 (N_5557,N_3369,N_4880);
nand U5558 (N_5558,N_3521,N_2716);
nor U5559 (N_5559,N_4809,N_4220);
and U5560 (N_5560,N_2962,N_4630);
or U5561 (N_5561,N_3534,N_4626);
nor U5562 (N_5562,N_3989,N_2872);
nand U5563 (N_5563,N_2785,N_4063);
and U5564 (N_5564,N_4291,N_2555);
nand U5565 (N_5565,N_2923,N_4272);
and U5566 (N_5566,N_4629,N_3675);
nand U5567 (N_5567,N_4673,N_3007);
or U5568 (N_5568,N_2831,N_4023);
nand U5569 (N_5569,N_4869,N_4496);
nor U5570 (N_5570,N_4079,N_3727);
nor U5571 (N_5571,N_2611,N_2942);
and U5572 (N_5572,N_3924,N_2945);
nor U5573 (N_5573,N_3424,N_3049);
nand U5574 (N_5574,N_4769,N_3387);
or U5575 (N_5575,N_4180,N_4025);
nand U5576 (N_5576,N_3665,N_4144);
or U5577 (N_5577,N_4588,N_3530);
or U5578 (N_5578,N_4820,N_4881);
and U5579 (N_5579,N_2658,N_3231);
nor U5580 (N_5580,N_2512,N_4126);
nand U5581 (N_5581,N_4136,N_4399);
and U5582 (N_5582,N_4911,N_2539);
and U5583 (N_5583,N_3673,N_3659);
or U5584 (N_5584,N_3053,N_3507);
or U5585 (N_5585,N_4469,N_4045);
and U5586 (N_5586,N_4848,N_2724);
or U5587 (N_5587,N_4833,N_4689);
or U5588 (N_5588,N_2822,N_2726);
nand U5589 (N_5589,N_3222,N_3958);
or U5590 (N_5590,N_4110,N_2565);
or U5591 (N_5591,N_4958,N_2970);
nand U5592 (N_5592,N_4358,N_4321);
and U5593 (N_5593,N_2830,N_3212);
and U5594 (N_5594,N_2916,N_4818);
or U5595 (N_5595,N_2642,N_4186);
nand U5596 (N_5596,N_3595,N_4694);
or U5597 (N_5597,N_3173,N_4075);
and U5598 (N_5598,N_4054,N_3538);
nand U5599 (N_5599,N_3579,N_3302);
nand U5600 (N_5600,N_2528,N_2951);
nand U5601 (N_5601,N_2953,N_3844);
and U5602 (N_5602,N_4205,N_2986);
or U5603 (N_5603,N_3100,N_3624);
nor U5604 (N_5604,N_4896,N_4733);
or U5605 (N_5605,N_3971,N_4717);
or U5606 (N_5606,N_4842,N_3246);
nand U5607 (N_5607,N_2574,N_3944);
nand U5608 (N_5608,N_4064,N_4665);
nor U5609 (N_5609,N_3281,N_4768);
or U5610 (N_5610,N_3217,N_4620);
or U5611 (N_5611,N_4490,N_3707);
nor U5612 (N_5612,N_4361,N_3543);
nand U5613 (N_5613,N_4230,N_3215);
and U5614 (N_5614,N_4685,N_4979);
and U5615 (N_5615,N_4724,N_3019);
and U5616 (N_5616,N_4280,N_3026);
and U5617 (N_5617,N_4741,N_2906);
and U5618 (N_5618,N_4601,N_3052);
or U5619 (N_5619,N_4252,N_3240);
or U5620 (N_5620,N_4007,N_4758);
nand U5621 (N_5621,N_4038,N_4808);
nand U5622 (N_5622,N_4201,N_3348);
and U5623 (N_5623,N_2502,N_4581);
nand U5624 (N_5624,N_4729,N_3775);
or U5625 (N_5625,N_4432,N_2787);
or U5626 (N_5626,N_4893,N_3203);
nand U5627 (N_5627,N_4157,N_4261);
and U5628 (N_5628,N_3467,N_3174);
nor U5629 (N_5629,N_2694,N_3846);
nand U5630 (N_5630,N_3455,N_2799);
nand U5631 (N_5631,N_3828,N_3234);
or U5632 (N_5632,N_4004,N_3370);
and U5633 (N_5633,N_4574,N_2990);
or U5634 (N_5634,N_3887,N_2573);
and U5635 (N_5635,N_4903,N_3514);
and U5636 (N_5636,N_4901,N_3435);
nand U5637 (N_5637,N_3398,N_2593);
nand U5638 (N_5638,N_4541,N_4849);
and U5639 (N_5639,N_4914,N_3639);
and U5640 (N_5640,N_3499,N_4547);
and U5641 (N_5641,N_2889,N_3109);
nand U5642 (N_5642,N_3742,N_4428);
nand U5643 (N_5643,N_2920,N_3082);
and U5644 (N_5644,N_4448,N_3442);
and U5645 (N_5645,N_3220,N_3154);
nor U5646 (N_5646,N_4185,N_2997);
or U5647 (N_5647,N_4179,N_3350);
nor U5648 (N_5648,N_3877,N_4442);
nor U5649 (N_5649,N_3025,N_2511);
nor U5650 (N_5650,N_2515,N_2781);
and U5651 (N_5651,N_3061,N_4857);
or U5652 (N_5652,N_2563,N_4336);
and U5653 (N_5653,N_3192,N_4844);
and U5654 (N_5654,N_3786,N_3880);
or U5655 (N_5655,N_4843,N_4287);
and U5656 (N_5656,N_4776,N_4047);
nor U5657 (N_5657,N_4032,N_4520);
and U5658 (N_5658,N_4426,N_3759);
or U5659 (N_5659,N_4810,N_4666);
and U5660 (N_5660,N_3598,N_4380);
nor U5661 (N_5661,N_2552,N_4370);
or U5662 (N_5662,N_2608,N_4036);
nand U5663 (N_5663,N_2527,N_4141);
and U5664 (N_5664,N_4790,N_4927);
nor U5665 (N_5665,N_2898,N_3987);
xor U5666 (N_5666,N_3489,N_4487);
or U5667 (N_5667,N_3233,N_2774);
nand U5668 (N_5668,N_4431,N_3209);
or U5669 (N_5669,N_2714,N_2910);
nor U5670 (N_5670,N_4174,N_3119);
nor U5671 (N_5671,N_3471,N_2674);
nor U5672 (N_5672,N_4247,N_4970);
or U5673 (N_5673,N_4695,N_3781);
nor U5674 (N_5674,N_4900,N_3939);
and U5675 (N_5675,N_3286,N_4602);
nand U5676 (N_5676,N_2930,N_4551);
nor U5677 (N_5677,N_4033,N_4460);
nand U5678 (N_5678,N_3146,N_3279);
xor U5679 (N_5679,N_3714,N_4115);
nor U5680 (N_5680,N_2741,N_2835);
nor U5681 (N_5681,N_3536,N_3013);
or U5682 (N_5682,N_2800,N_2524);
and U5683 (N_5683,N_3475,N_3909);
nor U5684 (N_5684,N_3564,N_4986);
or U5685 (N_5685,N_3934,N_4098);
or U5686 (N_5686,N_4439,N_3931);
or U5687 (N_5687,N_4981,N_4175);
or U5688 (N_5688,N_2978,N_4706);
nor U5689 (N_5689,N_2601,N_3804);
or U5690 (N_5690,N_4143,N_3268);
nand U5691 (N_5691,N_4006,N_2712);
and U5692 (N_5692,N_4482,N_3079);
or U5693 (N_5693,N_3862,N_4658);
or U5694 (N_5694,N_2929,N_3914);
nor U5695 (N_5695,N_4166,N_3364);
nand U5696 (N_5696,N_3045,N_4156);
or U5697 (N_5697,N_2663,N_3790);
nand U5698 (N_5698,N_4394,N_4058);
or U5699 (N_5699,N_3705,N_3905);
nand U5700 (N_5700,N_3225,N_3063);
xor U5701 (N_5701,N_4548,N_3484);
nand U5702 (N_5702,N_4255,N_4827);
or U5703 (N_5703,N_3251,N_4663);
or U5704 (N_5704,N_4202,N_3239);
or U5705 (N_5705,N_4738,N_2630);
nand U5706 (N_5706,N_3076,N_4543);
nor U5707 (N_5707,N_3479,N_4836);
nand U5708 (N_5708,N_4229,N_2548);
and U5709 (N_5709,N_4251,N_3641);
nand U5710 (N_5710,N_3353,N_2784);
nand U5711 (N_5711,N_3782,N_3316);
nand U5712 (N_5712,N_4436,N_3237);
or U5713 (N_5713,N_4802,N_3051);
nor U5714 (N_5714,N_4909,N_4614);
or U5715 (N_5715,N_4751,N_3072);
nand U5716 (N_5716,N_4538,N_3937);
or U5717 (N_5717,N_3616,N_3503);
nand U5718 (N_5718,N_4966,N_4823);
nand U5719 (N_5719,N_3713,N_3979);
and U5720 (N_5720,N_4621,N_4977);
nand U5721 (N_5721,N_2519,N_2857);
nand U5722 (N_5722,N_3472,N_4030);
nor U5723 (N_5723,N_3255,N_4997);
nor U5724 (N_5724,N_2899,N_3309);
nor U5725 (N_5725,N_2975,N_2667);
nor U5726 (N_5726,N_3208,N_4425);
or U5727 (N_5727,N_4950,N_4331);
or U5728 (N_5728,N_3323,N_3338);
nor U5729 (N_5729,N_4417,N_4453);
nor U5730 (N_5730,N_2607,N_3016);
or U5731 (N_5731,N_2823,N_3610);
nand U5732 (N_5732,N_3008,N_2813);
nor U5733 (N_5733,N_2904,N_4081);
nand U5734 (N_5734,N_4887,N_2870);
nand U5735 (N_5735,N_3589,N_3747);
and U5736 (N_5736,N_4276,N_4969);
nor U5737 (N_5737,N_4196,N_2586);
nor U5738 (N_5738,N_3947,N_4576);
or U5739 (N_5739,N_4782,N_2588);
and U5740 (N_5740,N_3920,N_2681);
nor U5741 (N_5741,N_3147,N_3981);
nor U5742 (N_5742,N_2558,N_2907);
or U5743 (N_5743,N_4285,N_4793);
and U5744 (N_5744,N_3701,N_4584);
nor U5745 (N_5745,N_4888,N_3456);
nand U5746 (N_5746,N_3030,N_3009);
nand U5747 (N_5747,N_3328,N_4061);
and U5748 (N_5748,N_3314,N_3631);
and U5749 (N_5749,N_4841,N_3085);
nand U5750 (N_5750,N_2894,N_3447);
nand U5751 (N_5751,N_3397,N_3493);
or U5752 (N_5752,N_4405,N_4686);
nor U5753 (N_5753,N_3046,N_4279);
or U5754 (N_5754,N_4822,N_2811);
nor U5755 (N_5755,N_3674,N_3307);
nor U5756 (N_5756,N_4500,N_4323);
nand U5757 (N_5757,N_2973,N_3873);
and U5758 (N_5758,N_4113,N_4314);
nand U5759 (N_5759,N_3122,N_2530);
and U5760 (N_5760,N_4565,N_3561);
nand U5761 (N_5761,N_3975,N_4915);
or U5762 (N_5762,N_4783,N_3105);
or U5763 (N_5763,N_2693,N_4570);
nand U5764 (N_5764,N_4015,N_4176);
nor U5765 (N_5765,N_4972,N_4147);
and U5766 (N_5766,N_4164,N_3434);
or U5767 (N_5767,N_3438,N_2676);
nor U5768 (N_5768,N_3490,N_3166);
or U5769 (N_5769,N_2652,N_3822);
and U5770 (N_5770,N_3576,N_4660);
nor U5771 (N_5771,N_2579,N_4254);
or U5772 (N_5772,N_3118,N_2861);
nand U5773 (N_5773,N_2874,N_3882);
and U5774 (N_5774,N_2824,N_4794);
or U5775 (N_5775,N_3970,N_4774);
or U5776 (N_5776,N_4366,N_4978);
nand U5777 (N_5777,N_3492,N_4789);
nor U5778 (N_5778,N_2881,N_4498);
nand U5779 (N_5779,N_2538,N_2955);
or U5780 (N_5780,N_3160,N_4009);
or U5781 (N_5781,N_4005,N_3102);
and U5782 (N_5782,N_4173,N_3149);
nor U5783 (N_5783,N_4817,N_3568);
and U5784 (N_5784,N_3764,N_3330);
xnor U5785 (N_5785,N_3654,N_4017);
or U5786 (N_5786,N_4117,N_4070);
or U5787 (N_5787,N_4861,N_3627);
nor U5788 (N_5788,N_2640,N_4847);
nand U5789 (N_5789,N_4564,N_3515);
or U5790 (N_5790,N_3027,N_4941);
and U5791 (N_5791,N_4486,N_4253);
and U5792 (N_5792,N_3960,N_4270);
nand U5793 (N_5793,N_4627,N_3940);
and U5794 (N_5794,N_4701,N_3808);
nand U5795 (N_5795,N_4388,N_2843);
and U5796 (N_5796,N_4207,N_2745);
and U5797 (N_5797,N_3691,N_3684);
or U5798 (N_5798,N_4226,N_3423);
and U5799 (N_5799,N_3767,N_4612);
nor U5800 (N_5800,N_3197,N_3708);
or U5801 (N_5801,N_2846,N_4675);
nand U5802 (N_5802,N_3480,N_3559);
nand U5803 (N_5803,N_4391,N_2577);
nand U5804 (N_5804,N_3452,N_4114);
nor U5805 (N_5805,N_3874,N_3282);
nand U5806 (N_5806,N_4754,N_4960);
nand U5807 (N_5807,N_4522,N_4403);
nor U5808 (N_5808,N_4928,N_3840);
nand U5809 (N_5809,N_4445,N_4282);
nor U5810 (N_5810,N_3140,N_2677);
nor U5811 (N_5811,N_2670,N_4740);
or U5812 (N_5812,N_3324,N_3608);
nor U5813 (N_5813,N_4446,N_3221);
and U5814 (N_5814,N_3716,N_4169);
nor U5815 (N_5815,N_3913,N_4048);
nand U5816 (N_5816,N_4210,N_2648);
nor U5817 (N_5817,N_2773,N_4647);
or U5818 (N_5818,N_4283,N_3967);
or U5819 (N_5819,N_4918,N_3326);
nand U5820 (N_5820,N_3793,N_4122);
nor U5821 (N_5821,N_2535,N_3778);
nor U5822 (N_5822,N_4553,N_4561);
nor U5823 (N_5823,N_4127,N_4654);
and U5824 (N_5824,N_3933,N_4693);
nand U5825 (N_5825,N_4204,N_3512);
or U5826 (N_5826,N_4919,N_4839);
or U5827 (N_5827,N_2877,N_3178);
nand U5828 (N_5828,N_4968,N_4406);
nand U5829 (N_5829,N_4389,N_3390);
or U5830 (N_5830,N_3366,N_2981);
or U5831 (N_5831,N_3172,N_4182);
and U5832 (N_5832,N_4148,N_4468);
nor U5833 (N_5833,N_4690,N_4595);
and U5834 (N_5834,N_2556,N_4043);
or U5835 (N_5835,N_3129,N_4532);
or U5836 (N_5836,N_4517,N_4142);
nor U5837 (N_5837,N_4168,N_3261);
or U5838 (N_5838,N_3615,N_3064);
and U5839 (N_5839,N_3069,N_4610);
nand U5840 (N_5840,N_4343,N_3841);
or U5841 (N_5841,N_3645,N_2532);
nor U5842 (N_5842,N_4696,N_3444);
nand U5843 (N_5843,N_4364,N_4222);
nand U5844 (N_5844,N_4618,N_3601);
and U5845 (N_5845,N_4286,N_3902);
nand U5846 (N_5846,N_4932,N_3206);
or U5847 (N_5847,N_2513,N_4757);
nand U5848 (N_5848,N_3679,N_2987);
nor U5849 (N_5849,N_2969,N_3784);
and U5850 (N_5850,N_4267,N_4451);
nand U5851 (N_5851,N_4077,N_4150);
nor U5852 (N_5852,N_2500,N_3956);
nor U5853 (N_5853,N_4835,N_2845);
or U5854 (N_5854,N_4159,N_4489);
nor U5855 (N_5855,N_2882,N_2767);
nor U5856 (N_5856,N_3059,N_3358);
nor U5857 (N_5857,N_3388,N_3074);
nand U5858 (N_5858,N_4249,N_3621);
nor U5859 (N_5859,N_4852,N_4305);
nand U5860 (N_5860,N_4160,N_3232);
or U5861 (N_5861,N_2709,N_4470);
nor U5862 (N_5862,N_4227,N_2572);
and U5863 (N_5863,N_3274,N_3285);
nor U5864 (N_5864,N_4258,N_2659);
xor U5865 (N_5865,N_3505,N_3520);
or U5866 (N_5866,N_3461,N_3227);
nand U5867 (N_5867,N_4146,N_3938);
nand U5868 (N_5868,N_3951,N_3722);
or U5869 (N_5869,N_3544,N_3843);
nand U5870 (N_5870,N_3796,N_3721);
and U5871 (N_5871,N_4197,N_4028);
and U5872 (N_5872,N_4944,N_3532);
nor U5873 (N_5873,N_3210,N_3303);
nand U5874 (N_5874,N_2547,N_4422);
nand U5875 (N_5875,N_3123,N_4300);
nor U5876 (N_5876,N_2866,N_4648);
nand U5877 (N_5877,N_4372,N_4898);
nor U5878 (N_5878,N_2853,N_4050);
or U5879 (N_5879,N_3680,N_2583);
and U5880 (N_5880,N_4943,N_4524);
nor U5881 (N_5881,N_4819,N_3990);
and U5882 (N_5882,N_2892,N_2998);
nor U5883 (N_5883,N_3820,N_3169);
nand U5884 (N_5884,N_3410,N_3299);
and U5885 (N_5885,N_2766,N_3213);
nand U5886 (N_5886,N_4967,N_4367);
or U5887 (N_5887,N_2633,N_3374);
and U5888 (N_5888,N_3478,N_3494);
nand U5889 (N_5889,N_3732,N_4190);
or U5890 (N_5890,N_3710,N_2977);
or U5891 (N_5891,N_4519,N_3264);
and U5892 (N_5892,N_2919,N_2685);
nand U5893 (N_5893,N_4980,N_4770);
nand U5894 (N_5894,N_3993,N_3823);
or U5895 (N_5895,N_2501,N_2944);
and U5896 (N_5896,N_3760,N_2665);
and U5897 (N_5897,N_4709,N_3896);
nor U5898 (N_5898,N_3738,N_3226);
or U5899 (N_5899,N_2602,N_2661);
nor U5900 (N_5900,N_4906,N_4294);
or U5901 (N_5901,N_3644,N_3656);
nor U5902 (N_5902,N_2808,N_4284);
nand U5903 (N_5903,N_3548,N_2791);
nor U5904 (N_5904,N_2890,N_4128);
or U5905 (N_5905,N_4813,N_4777);
or U5906 (N_5906,N_4443,N_3519);
nand U5907 (N_5907,N_4327,N_2666);
and U5908 (N_5908,N_2858,N_2884);
nand U5909 (N_5909,N_3189,N_3930);
nand U5910 (N_5910,N_2717,N_4611);
nand U5911 (N_5911,N_2802,N_4995);
or U5912 (N_5912,N_2810,N_4355);
or U5913 (N_5913,N_2503,N_3466);
or U5914 (N_5914,N_3482,N_4542);
nand U5915 (N_5915,N_2510,N_2995);
nor U5916 (N_5916,N_4371,N_2819);
and U5917 (N_5917,N_4386,N_3892);
nor U5918 (N_5918,N_3252,N_3395);
nand U5919 (N_5919,N_4477,N_3024);
nor U5920 (N_5920,N_3267,N_4444);
or U5921 (N_5921,N_2578,N_4069);
nor U5922 (N_5922,N_4737,N_3587);
and U5923 (N_5923,N_4908,N_4396);
or U5924 (N_5924,N_4940,N_4404);
nand U5925 (N_5925,N_4200,N_4591);
or U5926 (N_5926,N_4525,N_3648);
or U5927 (N_5927,N_4962,N_4170);
nor U5928 (N_5928,N_4472,N_2851);
or U5929 (N_5929,N_3635,N_4624);
nand U5930 (N_5930,N_4344,N_3695);
or U5931 (N_5931,N_2818,N_3609);
or U5932 (N_5932,N_2536,N_3409);
or U5933 (N_5933,N_4746,N_4723);
nor U5934 (N_5934,N_4714,N_3368);
and U5935 (N_5935,N_3032,N_3667);
and U5936 (N_5936,N_3495,N_4878);
nand U5937 (N_5937,N_4221,N_4483);
and U5938 (N_5938,N_3177,N_2756);
nor U5939 (N_5939,N_2934,N_3972);
nand U5940 (N_5940,N_4401,N_3954);
or U5941 (N_5941,N_3547,N_4540);
nand U5942 (N_5942,N_2752,N_3553);
and U5943 (N_5943,N_3835,N_3657);
or U5944 (N_5944,N_4825,N_2869);
or U5945 (N_5945,N_3313,N_4052);
and U5946 (N_5946,N_3242,N_2504);
or U5947 (N_5947,N_2963,N_4587);
and U5948 (N_5948,N_3946,N_4635);
nor U5949 (N_5949,N_3523,N_4580);
nand U5950 (N_5950,N_4062,N_2614);
nor U5951 (N_5951,N_3344,N_2950);
nand U5952 (N_5952,N_2529,N_3799);
nand U5953 (N_5953,N_4954,N_4421);
nor U5954 (N_5954,N_3825,N_3921);
nor U5955 (N_5955,N_2921,N_3416);
or U5956 (N_5956,N_2725,N_4856);
nor U5957 (N_5957,N_4211,N_3952);
and U5958 (N_5958,N_4605,N_2803);
xnor U5959 (N_5959,N_3245,N_3600);
nand U5960 (N_5960,N_3187,N_3463);
nand U5961 (N_5961,N_3871,N_2878);
nand U5962 (N_5962,N_3597,N_2589);
nand U5963 (N_5963,N_4044,N_4705);
nor U5964 (N_5964,N_2964,N_4494);
or U5965 (N_5965,N_4378,N_3153);
nand U5966 (N_5966,N_4683,N_3327);
or U5967 (N_5967,N_4317,N_2580);
and U5968 (N_5968,N_3276,N_2678);
or U5969 (N_5969,N_3002,N_3376);
nor U5970 (N_5970,N_4271,N_2778);
and U5971 (N_5971,N_2516,N_4465);
nor U5972 (N_5972,N_4457,N_2782);
or U5973 (N_5973,N_2928,N_3381);
nor U5974 (N_5974,N_2587,N_3201);
nand U5975 (N_5975,N_4040,N_3005);
nor U5976 (N_5976,N_2560,N_3300);
or U5977 (N_5977,N_3697,N_2926);
or U5978 (N_5978,N_3347,N_2707);
xnor U5979 (N_5979,N_2993,N_2599);
or U5980 (N_5980,N_3814,N_3650);
nor U5981 (N_5981,N_3229,N_4377);
nand U5982 (N_5982,N_3661,N_3725);
nor U5983 (N_5983,N_4450,N_4330);
or U5984 (N_5984,N_2967,N_2924);
nand U5985 (N_5985,N_4592,N_3860);
nor U5986 (N_5986,N_4636,N_2711);
nor U5987 (N_5987,N_3196,N_4085);
and U5988 (N_5988,N_3086,N_4119);
nand U5989 (N_5989,N_2850,N_4199);
nand U5990 (N_5990,N_4639,N_3772);
or U5991 (N_5991,N_2865,N_3566);
or U5992 (N_5992,N_4049,N_3486);
nand U5993 (N_5993,N_4687,N_2769);
nor U5994 (N_5994,N_2988,N_3462);
nand U5995 (N_5995,N_4152,N_3885);
nand U5996 (N_5996,N_2523,N_4529);
nand U5997 (N_5997,N_3599,N_3690);
or U5998 (N_5998,N_3060,N_2618);
and U5999 (N_5999,N_4013,N_3649);
nand U6000 (N_6000,N_3728,N_2732);
nor U6001 (N_6001,N_3401,N_3581);
and U6002 (N_6002,N_2755,N_3908);
nand U6003 (N_6003,N_4983,N_3623);
nand U6004 (N_6004,N_4664,N_2913);
nor U6005 (N_6005,N_4263,N_4375);
or U6006 (N_6006,N_2749,N_4218);
nor U6007 (N_6007,N_3012,N_4907);
nand U6008 (N_6008,N_3900,N_2912);
or U6009 (N_6009,N_2832,N_2735);
nor U6010 (N_6010,N_4785,N_4953);
and U6011 (N_6011,N_2632,N_4103);
and U6012 (N_6012,N_3699,N_3223);
and U6013 (N_6013,N_3241,N_4315);
nand U6014 (N_6014,N_3332,N_4107);
nor U6015 (N_6015,N_2697,N_4296);
nor U6016 (N_6016,N_2582,N_3380);
or U6017 (N_6017,N_3185,N_3584);
nor U6018 (N_6018,N_4311,N_3818);
nor U6019 (N_6019,N_2868,N_3813);
nor U6020 (N_6020,N_3974,N_3156);
and U6021 (N_6021,N_4010,N_3508);
and U6022 (N_6022,N_3985,N_2844);
nor U6023 (N_6023,N_4129,N_3766);
nand U6024 (N_6024,N_2759,N_4545);
nand U6025 (N_6025,N_4301,N_2827);
or U6026 (N_6026,N_4765,N_4350);
or U6027 (N_6027,N_4060,N_3288);
and U6028 (N_6028,N_4745,N_3253);
nor U6029 (N_6029,N_2909,N_2994);
nand U6030 (N_6030,N_2540,N_2820);
and U6031 (N_6031,N_4212,N_3962);
nand U6032 (N_6032,N_3037,N_3343);
nor U6033 (N_6033,N_4188,N_2902);
and U6034 (N_6034,N_4711,N_4989);
nand U6035 (N_6035,N_3248,N_2900);
and U6036 (N_6036,N_2613,N_4600);
and U6037 (N_6037,N_3545,N_3384);
or U6038 (N_6038,N_2908,N_4949);
or U6039 (N_6039,N_3023,N_3770);
nor U6040 (N_6040,N_4208,N_3517);
nor U6041 (N_6041,N_3065,N_2770);
and U6042 (N_6042,N_4131,N_4325);
nor U6043 (N_6043,N_4637,N_3810);
and U6044 (N_6044,N_2976,N_4526);
and U6045 (N_6045,N_3335,N_4948);
nand U6046 (N_6046,N_3779,N_4031);
and U6047 (N_6047,N_4930,N_3273);
or U6048 (N_6048,N_4259,N_2943);
or U6049 (N_6049,N_4568,N_3861);
nand U6050 (N_6050,N_4012,N_4608);
nor U6051 (N_6051,N_3391,N_4891);
or U6052 (N_6052,N_4801,N_3430);
and U6053 (N_6053,N_2760,N_4539);
nor U6054 (N_6054,N_2657,N_2692);
or U6055 (N_6055,N_2809,N_3634);
and U6056 (N_6056,N_4634,N_3135);
nor U6057 (N_6057,N_2543,N_4535);
or U6058 (N_6058,N_4708,N_2911);
and U6059 (N_6059,N_4569,N_2783);
or U6060 (N_6060,N_3899,N_3204);
nand U6061 (N_6061,N_3717,N_2729);
nor U6062 (N_6062,N_4318,N_4638);
and U6063 (N_6063,N_3179,N_3081);
nor U6064 (N_6064,N_3607,N_4102);
nor U6065 (N_6065,N_3682,N_2507);
or U6066 (N_6066,N_4072,N_2689);
nand U6067 (N_6067,N_4718,N_2825);
xor U6068 (N_6068,N_3588,N_4019);
nand U6069 (N_6069,N_4987,N_2704);
or U6070 (N_6070,N_3941,N_3837);
or U6071 (N_6071,N_3554,N_4316);
and U6072 (N_6072,N_3526,N_4151);
or U6073 (N_6073,N_3864,N_4395);
nor U6074 (N_6074,N_4339,N_2542);
or U6075 (N_6075,N_3783,N_3346);
nor U6076 (N_6076,N_3511,N_3048);
nand U6077 (N_6077,N_2651,N_4961);
nand U6078 (N_6078,N_2653,N_2639);
nor U6079 (N_6079,N_3509,N_4766);
nor U6080 (N_6080,N_4641,N_3756);
or U6081 (N_6081,N_3787,N_4288);
nand U6082 (N_6082,N_2598,N_3748);
nor U6083 (N_6083,N_2742,N_4899);
or U6084 (N_6084,N_3662,N_4759);
nor U6085 (N_6085,N_3876,N_4837);
or U6086 (N_6086,N_2960,N_3733);
or U6087 (N_6087,N_4093,N_2595);
or U6088 (N_6088,N_2597,N_3736);
or U6089 (N_6089,N_4702,N_2796);
nor U6090 (N_6090,N_2806,N_4905);
or U6091 (N_6091,N_3097,N_4744);
and U6092 (N_6092,N_3136,N_4889);
nand U6093 (N_6093,N_4846,N_3977);
or U6094 (N_6094,N_2683,N_4329);
or U6095 (N_6095,N_3319,N_4409);
or U6096 (N_6096,N_4242,N_4863);
and U6097 (N_6097,N_4544,N_4065);
xor U6098 (N_6098,N_3171,N_4232);
or U6099 (N_6099,N_4016,N_4292);
nor U6100 (N_6100,N_4772,N_4531);
or U6101 (N_6101,N_4736,N_3957);
and U6102 (N_6102,N_3161,N_3803);
or U6103 (N_6103,N_4337,N_4250);
nor U6104 (N_6104,N_2901,N_4125);
nand U6105 (N_6105,N_4231,N_4219);
or U6106 (N_6106,N_4771,N_3906);
nand U6107 (N_6107,N_4293,N_3078);
or U6108 (N_6108,N_4537,N_3513);
and U6109 (N_6109,N_4235,N_4999);
and U6110 (N_6110,N_3497,N_4613);
nor U6111 (N_6111,N_3794,N_2771);
or U6112 (N_6112,N_3441,N_2654);
or U6113 (N_6113,N_4973,N_3557);
or U6114 (N_6114,N_3719,N_3729);
and U6115 (N_6115,N_4985,N_3018);
and U6116 (N_6116,N_3950,N_2961);
nand U6117 (N_6117,N_3450,N_4873);
or U6118 (N_6118,N_3969,N_4886);
nand U6119 (N_6119,N_3112,N_2838);
nor U6120 (N_6120,N_3145,N_2754);
nor U6121 (N_6121,N_3029,N_3556);
nand U6122 (N_6122,N_2564,N_4492);
nand U6123 (N_6123,N_2638,N_2720);
nor U6124 (N_6124,N_4762,N_4559);
or U6125 (N_6125,N_4273,N_2917);
or U6126 (N_6126,N_2591,N_3542);
or U6127 (N_6127,N_3198,N_4688);
nor U6128 (N_6128,N_4464,N_3537);
or U6129 (N_6129,N_3518,N_4743);
nand U6130 (N_6130,N_2896,N_4106);
or U6131 (N_6131,N_2645,N_2895);
and U6132 (N_6132,N_3340,N_3117);
nand U6133 (N_6133,N_2576,N_2837);
and U6134 (N_6134,N_3379,N_3901);
nand U6135 (N_6135,N_4262,N_2933);
and U6136 (N_6136,N_2748,N_4902);
nand U6137 (N_6137,N_3202,N_3709);
or U6138 (N_6138,N_3236,N_3440);
or U6139 (N_6139,N_4676,N_4534);
and U6140 (N_6140,N_2636,N_2620);
or U6141 (N_6141,N_4656,N_4360);
nor U6142 (N_6142,N_4471,N_3535);
nor U6143 (N_6143,N_4892,N_2834);
nand U6144 (N_6144,N_2719,N_4461);
and U6145 (N_6145,N_2566,N_3003);
and U6146 (N_6146,N_3851,N_2989);
nor U6147 (N_6147,N_2879,N_3560);
or U6148 (N_6148,N_3910,N_3994);
and U6149 (N_6149,N_3619,N_3042);
or U6150 (N_6150,N_4080,N_4322);
nand U6151 (N_6151,N_2817,N_3743);
nand U6152 (N_6152,N_3428,N_3681);
or U6153 (N_6153,N_4715,N_4096);
and U6154 (N_6154,N_3359,N_2514);
and U6155 (N_6155,N_4874,N_3927);
nor U6156 (N_6156,N_3271,N_3984);
and U6157 (N_6157,N_3247,N_2696);
nor U6158 (N_6158,N_3614,N_3200);
and U6159 (N_6159,N_2949,N_3569);
or U6160 (N_6160,N_4447,N_3365);
or U6161 (N_6161,N_3035,N_4024);
or U6162 (N_6162,N_3419,N_3386);
or U6163 (N_6163,N_3355,N_2710);
nand U6164 (N_6164,N_3752,N_3893);
nor U6165 (N_6165,N_4791,N_3297);
nand U6166 (N_6166,N_3806,N_3574);
or U6167 (N_6167,N_4804,N_3637);
and U6168 (N_6168,N_3982,N_4345);
xor U6169 (N_6169,N_2521,N_2925);
nand U6170 (N_6170,N_3852,N_3776);
nand U6171 (N_6171,N_3244,N_4678);
nor U6172 (N_6172,N_4217,N_4679);
nor U6173 (N_6173,N_4853,N_3394);
and U6174 (N_6174,N_4193,N_3090);
nand U6175 (N_6175,N_4145,N_4579);
nor U6176 (N_6176,N_3773,N_3653);
nor U6177 (N_6177,N_3894,N_4897);
nor U6178 (N_6178,N_3706,N_3550);
or U6179 (N_6179,N_4994,N_4651);
xor U6180 (N_6180,N_3445,N_4140);
nor U6181 (N_6181,N_3311,N_4456);
nand U6182 (N_6182,N_4797,N_3789);
and U6183 (N_6183,N_3997,N_3487);
nor U6184 (N_6184,N_3858,N_2971);
nand U6185 (N_6185,N_4573,N_3304);
or U6186 (N_6186,N_4670,N_3586);
nor U6187 (N_6187,N_3357,N_4756);
nand U6188 (N_6188,N_4376,N_3075);
and U6189 (N_6189,N_2887,N_2594);
or U6190 (N_6190,N_3446,N_3663);
and U6191 (N_6191,N_3955,N_3626);
nor U6192 (N_6192,N_3148,N_4593);
nand U6193 (N_6193,N_3089,N_4416);
or U6194 (N_6194,N_3768,N_3437);
or U6195 (N_6195,N_2743,N_2915);
and U6196 (N_6196,N_3501,N_3935);
nor U6197 (N_6197,N_4011,N_3827);
or U6198 (N_6198,N_3809,N_3070);
nand U6199 (N_6199,N_3108,N_2980);
nand U6200 (N_6200,N_4297,N_4530);
nor U6201 (N_6201,N_2871,N_4215);
and U6202 (N_6202,N_4578,N_3842);
and U6203 (N_6203,N_4792,N_4513);
and U6204 (N_6204,N_4528,N_4692);
nor U6205 (N_6205,N_2772,N_4328);
and U6206 (N_6206,N_4585,N_3325);
nand U6207 (N_6207,N_2550,N_4413);
and U6208 (N_6208,N_2914,N_4761);
nor U6209 (N_6209,N_3262,N_3868);
nor U6210 (N_6210,N_4357,N_4491);
nand U6211 (N_6211,N_2700,N_4312);
nor U6212 (N_6212,N_3170,N_3685);
nor U6213 (N_6213,N_4433,N_3291);
and U6214 (N_6214,N_3640,N_2984);
nand U6215 (N_6215,N_4739,N_3531);
nor U6216 (N_6216,N_4942,N_3694);
or U6217 (N_6217,N_2758,N_3339);
and U6218 (N_6218,N_4795,N_2518);
nand U6219 (N_6219,N_4299,N_3130);
and U6220 (N_6220,N_4516,N_4661);
nor U6221 (N_6221,N_3293,N_4485);
or U6222 (N_6222,N_3567,N_4203);
nor U6223 (N_6223,N_4194,N_4429);
nand U6224 (N_6224,N_4671,N_3998);
xnor U6225 (N_6225,N_4704,N_4586);
xnor U6226 (N_6226,N_4505,N_4171);
nand U6227 (N_6227,N_4755,N_3811);
and U6228 (N_6228,N_2947,N_3134);
and U6229 (N_6229,N_4824,N_3432);
nor U6230 (N_6230,N_3965,N_2612);
or U6231 (N_6231,N_4029,N_4567);
or U6232 (N_6232,N_4087,N_2508);
nand U6233 (N_6233,N_3133,N_3855);
nand U6234 (N_6234,N_4295,N_3978);
nand U6235 (N_6235,N_2680,N_4504);
and U6236 (N_6236,N_3726,N_2686);
nand U6237 (N_6237,N_3618,N_3159);
nor U6238 (N_6238,N_2807,N_4703);
or U6239 (N_6239,N_3762,N_4800);
and U6240 (N_6240,N_3422,N_2616);
and U6241 (N_6241,N_4652,N_4684);
and U6242 (N_6242,N_3034,N_4068);
nand U6243 (N_6243,N_4281,N_3420);
or U6244 (N_6244,N_3091,N_3188);
and U6245 (N_6245,N_2821,N_4731);
and U6246 (N_6246,N_4984,N_3345);
nand U6247 (N_6247,N_4324,N_2876);
nor U6248 (N_6248,N_3403,N_3250);
nand U6249 (N_6249,N_4484,N_2794);
nor U6250 (N_6250,N_2823,N_3453);
or U6251 (N_6251,N_3762,N_3822);
nor U6252 (N_6252,N_3733,N_2696);
nor U6253 (N_6253,N_3637,N_2510);
nand U6254 (N_6254,N_2503,N_4904);
and U6255 (N_6255,N_4398,N_4325);
xnor U6256 (N_6256,N_2678,N_4382);
or U6257 (N_6257,N_3189,N_3136);
nand U6258 (N_6258,N_2757,N_3751);
or U6259 (N_6259,N_3373,N_2905);
nor U6260 (N_6260,N_3344,N_4845);
nand U6261 (N_6261,N_4830,N_3267);
and U6262 (N_6262,N_3125,N_4941);
nor U6263 (N_6263,N_4300,N_3691);
nor U6264 (N_6264,N_4360,N_4975);
nand U6265 (N_6265,N_4095,N_3469);
nor U6266 (N_6266,N_3378,N_4568);
and U6267 (N_6267,N_4271,N_4905);
nand U6268 (N_6268,N_4096,N_3340);
or U6269 (N_6269,N_3449,N_3122);
and U6270 (N_6270,N_3857,N_2717);
or U6271 (N_6271,N_4200,N_4148);
or U6272 (N_6272,N_3364,N_3509);
nand U6273 (N_6273,N_3479,N_4892);
nor U6274 (N_6274,N_3679,N_3144);
nand U6275 (N_6275,N_4691,N_4470);
or U6276 (N_6276,N_3552,N_2835);
nor U6277 (N_6277,N_4699,N_4526);
and U6278 (N_6278,N_4470,N_3919);
nand U6279 (N_6279,N_4153,N_4093);
and U6280 (N_6280,N_4883,N_3612);
nand U6281 (N_6281,N_4832,N_4139);
nor U6282 (N_6282,N_3455,N_3093);
or U6283 (N_6283,N_2559,N_2755);
and U6284 (N_6284,N_3682,N_3835);
nor U6285 (N_6285,N_4875,N_3755);
nor U6286 (N_6286,N_3875,N_3381);
and U6287 (N_6287,N_4300,N_2656);
nand U6288 (N_6288,N_2612,N_4752);
nor U6289 (N_6289,N_3801,N_2544);
nor U6290 (N_6290,N_4402,N_2556);
xor U6291 (N_6291,N_4613,N_3347);
nand U6292 (N_6292,N_3827,N_2966);
nor U6293 (N_6293,N_4688,N_3533);
nor U6294 (N_6294,N_3715,N_2560);
or U6295 (N_6295,N_4439,N_4791);
or U6296 (N_6296,N_4161,N_3113);
nor U6297 (N_6297,N_3306,N_3247);
nand U6298 (N_6298,N_4538,N_2907);
nor U6299 (N_6299,N_2879,N_2987);
nand U6300 (N_6300,N_3400,N_4458);
nor U6301 (N_6301,N_3225,N_2870);
and U6302 (N_6302,N_2949,N_3486);
and U6303 (N_6303,N_2796,N_3137);
and U6304 (N_6304,N_4981,N_4852);
nor U6305 (N_6305,N_4766,N_3440);
and U6306 (N_6306,N_2666,N_3501);
nand U6307 (N_6307,N_4542,N_4016);
nand U6308 (N_6308,N_2760,N_3321);
nor U6309 (N_6309,N_3794,N_3105);
nor U6310 (N_6310,N_3917,N_3178);
nor U6311 (N_6311,N_3767,N_3486);
nand U6312 (N_6312,N_3081,N_3923);
nand U6313 (N_6313,N_4571,N_4269);
nor U6314 (N_6314,N_2699,N_2731);
and U6315 (N_6315,N_2561,N_4036);
or U6316 (N_6316,N_3415,N_3434);
and U6317 (N_6317,N_4828,N_2651);
xor U6318 (N_6318,N_3773,N_4822);
and U6319 (N_6319,N_4510,N_4651);
nor U6320 (N_6320,N_4123,N_3384);
or U6321 (N_6321,N_3495,N_4963);
and U6322 (N_6322,N_3740,N_4736);
xnor U6323 (N_6323,N_3656,N_2513);
or U6324 (N_6324,N_4783,N_3577);
nand U6325 (N_6325,N_3576,N_3537);
and U6326 (N_6326,N_4572,N_4405);
nor U6327 (N_6327,N_4330,N_4638);
or U6328 (N_6328,N_2673,N_2725);
and U6329 (N_6329,N_3971,N_4621);
or U6330 (N_6330,N_3845,N_3181);
or U6331 (N_6331,N_4256,N_2626);
and U6332 (N_6332,N_3744,N_4078);
xnor U6333 (N_6333,N_4592,N_4087);
nor U6334 (N_6334,N_4974,N_4457);
and U6335 (N_6335,N_3105,N_3883);
or U6336 (N_6336,N_4223,N_3840);
and U6337 (N_6337,N_4667,N_4089);
or U6338 (N_6338,N_2818,N_2770);
nand U6339 (N_6339,N_3637,N_3369);
nand U6340 (N_6340,N_3003,N_2640);
nor U6341 (N_6341,N_3082,N_3884);
nand U6342 (N_6342,N_3889,N_2552);
nor U6343 (N_6343,N_3769,N_3069);
or U6344 (N_6344,N_3676,N_4467);
or U6345 (N_6345,N_3947,N_3154);
or U6346 (N_6346,N_4503,N_3740);
nand U6347 (N_6347,N_4014,N_4695);
and U6348 (N_6348,N_4359,N_2691);
nand U6349 (N_6349,N_2947,N_3811);
or U6350 (N_6350,N_4245,N_3543);
nand U6351 (N_6351,N_4348,N_2860);
and U6352 (N_6352,N_4482,N_4048);
or U6353 (N_6353,N_2769,N_2925);
nand U6354 (N_6354,N_4790,N_3581);
and U6355 (N_6355,N_2943,N_3794);
or U6356 (N_6356,N_2572,N_2703);
or U6357 (N_6357,N_4513,N_3960);
or U6358 (N_6358,N_3295,N_3930);
nand U6359 (N_6359,N_3693,N_4312);
or U6360 (N_6360,N_4800,N_3619);
or U6361 (N_6361,N_4391,N_3156);
nand U6362 (N_6362,N_4878,N_4302);
or U6363 (N_6363,N_3797,N_4001);
nand U6364 (N_6364,N_2861,N_3015);
nand U6365 (N_6365,N_4122,N_3539);
nand U6366 (N_6366,N_4868,N_4227);
nor U6367 (N_6367,N_3266,N_4148);
nor U6368 (N_6368,N_4914,N_3708);
nor U6369 (N_6369,N_2798,N_4767);
and U6370 (N_6370,N_4889,N_2648);
and U6371 (N_6371,N_3388,N_4615);
nand U6372 (N_6372,N_4656,N_2529);
nor U6373 (N_6373,N_3320,N_3485);
nor U6374 (N_6374,N_4245,N_3734);
or U6375 (N_6375,N_2515,N_2640);
or U6376 (N_6376,N_4494,N_3240);
nor U6377 (N_6377,N_3616,N_4463);
or U6378 (N_6378,N_3766,N_3095);
or U6379 (N_6379,N_2700,N_3614);
nor U6380 (N_6380,N_2528,N_3348);
and U6381 (N_6381,N_2856,N_3194);
and U6382 (N_6382,N_3205,N_3043);
and U6383 (N_6383,N_3884,N_3966);
or U6384 (N_6384,N_4875,N_3667);
or U6385 (N_6385,N_3975,N_4318);
or U6386 (N_6386,N_3278,N_4645);
and U6387 (N_6387,N_2602,N_3420);
nand U6388 (N_6388,N_3802,N_3008);
nand U6389 (N_6389,N_3947,N_3740);
nand U6390 (N_6390,N_3657,N_3820);
or U6391 (N_6391,N_3754,N_4544);
and U6392 (N_6392,N_3062,N_2699);
and U6393 (N_6393,N_3486,N_3150);
or U6394 (N_6394,N_3629,N_4396);
nor U6395 (N_6395,N_3028,N_3576);
or U6396 (N_6396,N_3279,N_3147);
and U6397 (N_6397,N_2632,N_3790);
or U6398 (N_6398,N_3679,N_3281);
or U6399 (N_6399,N_2953,N_4843);
nor U6400 (N_6400,N_2587,N_3102);
nor U6401 (N_6401,N_4053,N_3938);
nand U6402 (N_6402,N_3674,N_4283);
nand U6403 (N_6403,N_4824,N_4574);
and U6404 (N_6404,N_4453,N_4699);
or U6405 (N_6405,N_3106,N_4144);
nor U6406 (N_6406,N_3640,N_4602);
and U6407 (N_6407,N_3557,N_3191);
nor U6408 (N_6408,N_3238,N_4852);
and U6409 (N_6409,N_2610,N_3746);
or U6410 (N_6410,N_4502,N_4528);
nor U6411 (N_6411,N_3632,N_3143);
nand U6412 (N_6412,N_4130,N_3903);
or U6413 (N_6413,N_2647,N_4060);
or U6414 (N_6414,N_3007,N_3536);
or U6415 (N_6415,N_4966,N_2664);
nand U6416 (N_6416,N_3597,N_3922);
and U6417 (N_6417,N_2907,N_3226);
nor U6418 (N_6418,N_4463,N_4065);
nor U6419 (N_6419,N_3878,N_3513);
nor U6420 (N_6420,N_3496,N_4015);
and U6421 (N_6421,N_2583,N_3094);
or U6422 (N_6422,N_3159,N_4073);
and U6423 (N_6423,N_4758,N_2717);
nand U6424 (N_6424,N_3285,N_3102);
or U6425 (N_6425,N_2581,N_2869);
and U6426 (N_6426,N_2853,N_3782);
nor U6427 (N_6427,N_3999,N_2801);
and U6428 (N_6428,N_3733,N_4930);
or U6429 (N_6429,N_3084,N_4795);
nand U6430 (N_6430,N_4735,N_3526);
or U6431 (N_6431,N_3952,N_3895);
nor U6432 (N_6432,N_2886,N_3101);
nor U6433 (N_6433,N_2526,N_2714);
nor U6434 (N_6434,N_3344,N_4444);
or U6435 (N_6435,N_3814,N_4979);
and U6436 (N_6436,N_4009,N_4438);
nor U6437 (N_6437,N_3126,N_4847);
or U6438 (N_6438,N_3873,N_4111);
nor U6439 (N_6439,N_3455,N_4291);
and U6440 (N_6440,N_3441,N_3853);
and U6441 (N_6441,N_3294,N_3684);
and U6442 (N_6442,N_2738,N_4890);
or U6443 (N_6443,N_3325,N_4748);
and U6444 (N_6444,N_4319,N_3287);
and U6445 (N_6445,N_2736,N_4492);
and U6446 (N_6446,N_4457,N_3022);
and U6447 (N_6447,N_4143,N_4231);
nor U6448 (N_6448,N_3306,N_3499);
xor U6449 (N_6449,N_4342,N_2753);
nand U6450 (N_6450,N_4771,N_2906);
and U6451 (N_6451,N_3504,N_3830);
nor U6452 (N_6452,N_4433,N_3661);
or U6453 (N_6453,N_4488,N_2679);
or U6454 (N_6454,N_3958,N_4560);
and U6455 (N_6455,N_4729,N_3851);
nand U6456 (N_6456,N_2851,N_3582);
and U6457 (N_6457,N_3568,N_3944);
nor U6458 (N_6458,N_3423,N_2931);
or U6459 (N_6459,N_4631,N_3268);
nor U6460 (N_6460,N_3741,N_3669);
and U6461 (N_6461,N_4777,N_2811);
nand U6462 (N_6462,N_3522,N_4503);
and U6463 (N_6463,N_2710,N_3835);
nor U6464 (N_6464,N_3095,N_4598);
and U6465 (N_6465,N_2824,N_3394);
and U6466 (N_6466,N_3623,N_4417);
or U6467 (N_6467,N_2624,N_2637);
nand U6468 (N_6468,N_4424,N_3113);
nor U6469 (N_6469,N_2804,N_4930);
nor U6470 (N_6470,N_3611,N_2783);
or U6471 (N_6471,N_3473,N_4884);
and U6472 (N_6472,N_2910,N_4999);
nand U6473 (N_6473,N_2771,N_4347);
or U6474 (N_6474,N_3937,N_3851);
and U6475 (N_6475,N_3189,N_4116);
nand U6476 (N_6476,N_3531,N_3744);
or U6477 (N_6477,N_2639,N_3284);
nor U6478 (N_6478,N_3044,N_4754);
nor U6479 (N_6479,N_3344,N_4203);
or U6480 (N_6480,N_3657,N_4143);
or U6481 (N_6481,N_3433,N_4514);
nand U6482 (N_6482,N_4545,N_3131);
nand U6483 (N_6483,N_3777,N_4848);
nand U6484 (N_6484,N_3654,N_3326);
or U6485 (N_6485,N_4934,N_4761);
nor U6486 (N_6486,N_3304,N_3315);
and U6487 (N_6487,N_4164,N_2941);
nor U6488 (N_6488,N_3736,N_3893);
and U6489 (N_6489,N_3932,N_3168);
nor U6490 (N_6490,N_3829,N_3601);
or U6491 (N_6491,N_3042,N_3782);
and U6492 (N_6492,N_4253,N_2879);
nor U6493 (N_6493,N_2841,N_3389);
or U6494 (N_6494,N_2863,N_3276);
or U6495 (N_6495,N_2955,N_3386);
nand U6496 (N_6496,N_2930,N_3684);
nor U6497 (N_6497,N_2924,N_4544);
or U6498 (N_6498,N_4527,N_3659);
nor U6499 (N_6499,N_4071,N_3553);
xor U6500 (N_6500,N_4564,N_2517);
nand U6501 (N_6501,N_3762,N_4312);
and U6502 (N_6502,N_3900,N_4951);
nor U6503 (N_6503,N_2616,N_2827);
nand U6504 (N_6504,N_3494,N_4527);
nor U6505 (N_6505,N_3737,N_4521);
nand U6506 (N_6506,N_3007,N_4616);
and U6507 (N_6507,N_4521,N_3609);
nand U6508 (N_6508,N_4210,N_3235);
and U6509 (N_6509,N_4632,N_4901);
and U6510 (N_6510,N_2644,N_2727);
or U6511 (N_6511,N_3788,N_4738);
and U6512 (N_6512,N_3883,N_4542);
and U6513 (N_6513,N_2692,N_4227);
nand U6514 (N_6514,N_4465,N_2623);
nand U6515 (N_6515,N_3777,N_4807);
nor U6516 (N_6516,N_4458,N_3584);
nand U6517 (N_6517,N_3490,N_3411);
nor U6518 (N_6518,N_4733,N_4272);
nor U6519 (N_6519,N_4329,N_3607);
and U6520 (N_6520,N_3572,N_4287);
nor U6521 (N_6521,N_3454,N_4200);
nor U6522 (N_6522,N_2625,N_4905);
and U6523 (N_6523,N_4840,N_2650);
nand U6524 (N_6524,N_2729,N_3189);
or U6525 (N_6525,N_3998,N_3479);
nand U6526 (N_6526,N_4503,N_2799);
nand U6527 (N_6527,N_4159,N_4958);
or U6528 (N_6528,N_2762,N_3033);
or U6529 (N_6529,N_4521,N_2603);
nor U6530 (N_6530,N_3426,N_4406);
or U6531 (N_6531,N_4806,N_3345);
or U6532 (N_6532,N_3574,N_3345);
or U6533 (N_6533,N_4010,N_3720);
and U6534 (N_6534,N_3862,N_3345);
nor U6535 (N_6535,N_3971,N_4113);
nand U6536 (N_6536,N_4986,N_2907);
nor U6537 (N_6537,N_4606,N_4859);
and U6538 (N_6538,N_3110,N_4297);
nor U6539 (N_6539,N_3750,N_4624);
nor U6540 (N_6540,N_4552,N_4707);
nor U6541 (N_6541,N_3513,N_3465);
nand U6542 (N_6542,N_4973,N_2822);
or U6543 (N_6543,N_3566,N_4244);
nor U6544 (N_6544,N_2812,N_3998);
nand U6545 (N_6545,N_4401,N_4478);
or U6546 (N_6546,N_3336,N_4658);
and U6547 (N_6547,N_3889,N_4633);
or U6548 (N_6548,N_4130,N_3518);
nand U6549 (N_6549,N_3869,N_3922);
and U6550 (N_6550,N_3445,N_4282);
nand U6551 (N_6551,N_3087,N_3062);
or U6552 (N_6552,N_4783,N_4079);
nor U6553 (N_6553,N_4909,N_4125);
nand U6554 (N_6554,N_4937,N_3411);
or U6555 (N_6555,N_4893,N_2780);
and U6556 (N_6556,N_3217,N_4363);
and U6557 (N_6557,N_3568,N_3241);
nor U6558 (N_6558,N_4896,N_2996);
and U6559 (N_6559,N_4253,N_4829);
nor U6560 (N_6560,N_2915,N_3989);
nand U6561 (N_6561,N_4137,N_4502);
nor U6562 (N_6562,N_4635,N_3196);
nand U6563 (N_6563,N_2573,N_4249);
or U6564 (N_6564,N_4951,N_3238);
or U6565 (N_6565,N_3829,N_3891);
nor U6566 (N_6566,N_4523,N_4776);
or U6567 (N_6567,N_2972,N_4935);
or U6568 (N_6568,N_3592,N_4895);
nand U6569 (N_6569,N_4926,N_3007);
or U6570 (N_6570,N_4179,N_3330);
nand U6571 (N_6571,N_3967,N_4020);
nand U6572 (N_6572,N_2630,N_2799);
or U6573 (N_6573,N_4668,N_3411);
or U6574 (N_6574,N_3085,N_4107);
nand U6575 (N_6575,N_2953,N_4089);
or U6576 (N_6576,N_4726,N_4722);
nor U6577 (N_6577,N_2937,N_4177);
and U6578 (N_6578,N_4041,N_4204);
nor U6579 (N_6579,N_2845,N_4152);
and U6580 (N_6580,N_4470,N_4751);
nand U6581 (N_6581,N_4841,N_3488);
nor U6582 (N_6582,N_2619,N_4365);
and U6583 (N_6583,N_4220,N_3106);
nor U6584 (N_6584,N_4947,N_3519);
nand U6585 (N_6585,N_3119,N_4823);
nand U6586 (N_6586,N_4100,N_4694);
and U6587 (N_6587,N_4724,N_4156);
or U6588 (N_6588,N_4125,N_2947);
and U6589 (N_6589,N_3262,N_4404);
nor U6590 (N_6590,N_3700,N_4065);
and U6591 (N_6591,N_2961,N_4724);
or U6592 (N_6592,N_4333,N_3208);
nor U6593 (N_6593,N_4288,N_4447);
nor U6594 (N_6594,N_4875,N_3119);
nor U6595 (N_6595,N_4760,N_3051);
nor U6596 (N_6596,N_3314,N_2958);
nor U6597 (N_6597,N_4900,N_2500);
nand U6598 (N_6598,N_3794,N_3225);
or U6599 (N_6599,N_3091,N_4075);
nand U6600 (N_6600,N_4831,N_4593);
and U6601 (N_6601,N_3861,N_3745);
nor U6602 (N_6602,N_2654,N_2945);
and U6603 (N_6603,N_3548,N_4220);
nor U6604 (N_6604,N_4552,N_4699);
nand U6605 (N_6605,N_3827,N_2898);
nand U6606 (N_6606,N_4071,N_3698);
nand U6607 (N_6607,N_4283,N_2669);
nand U6608 (N_6608,N_2948,N_3228);
nor U6609 (N_6609,N_3031,N_3938);
and U6610 (N_6610,N_3197,N_3263);
or U6611 (N_6611,N_2560,N_4144);
and U6612 (N_6612,N_3130,N_2721);
and U6613 (N_6613,N_4684,N_2657);
xor U6614 (N_6614,N_2719,N_4934);
or U6615 (N_6615,N_4841,N_4388);
xor U6616 (N_6616,N_3296,N_2633);
or U6617 (N_6617,N_2880,N_4992);
nor U6618 (N_6618,N_2507,N_2661);
or U6619 (N_6619,N_4759,N_4899);
nand U6620 (N_6620,N_2684,N_4976);
or U6621 (N_6621,N_3539,N_4914);
or U6622 (N_6622,N_3282,N_3979);
and U6623 (N_6623,N_4464,N_2530);
nor U6624 (N_6624,N_3416,N_4692);
and U6625 (N_6625,N_2870,N_3734);
and U6626 (N_6626,N_4353,N_3387);
or U6627 (N_6627,N_2629,N_3500);
and U6628 (N_6628,N_2869,N_3955);
or U6629 (N_6629,N_3097,N_3197);
nor U6630 (N_6630,N_4414,N_4310);
xnor U6631 (N_6631,N_2950,N_3529);
or U6632 (N_6632,N_3235,N_2526);
or U6633 (N_6633,N_3092,N_2726);
or U6634 (N_6634,N_3956,N_4301);
and U6635 (N_6635,N_3739,N_3372);
and U6636 (N_6636,N_2998,N_4457);
and U6637 (N_6637,N_4249,N_2870);
nor U6638 (N_6638,N_4754,N_3628);
nor U6639 (N_6639,N_4169,N_3566);
nor U6640 (N_6640,N_4558,N_3451);
nand U6641 (N_6641,N_3617,N_4563);
nand U6642 (N_6642,N_4976,N_2996);
and U6643 (N_6643,N_4569,N_3353);
nand U6644 (N_6644,N_2927,N_3542);
and U6645 (N_6645,N_4103,N_2861);
or U6646 (N_6646,N_3411,N_4514);
nor U6647 (N_6647,N_2922,N_2758);
and U6648 (N_6648,N_2904,N_2750);
nand U6649 (N_6649,N_2650,N_4787);
and U6650 (N_6650,N_2544,N_3113);
and U6651 (N_6651,N_2749,N_4896);
nand U6652 (N_6652,N_2518,N_4234);
nor U6653 (N_6653,N_4447,N_4179);
or U6654 (N_6654,N_4798,N_2659);
nand U6655 (N_6655,N_3302,N_4710);
nor U6656 (N_6656,N_4203,N_3257);
and U6657 (N_6657,N_2576,N_3470);
xnor U6658 (N_6658,N_2665,N_3443);
nor U6659 (N_6659,N_3036,N_3563);
nor U6660 (N_6660,N_2716,N_3001);
and U6661 (N_6661,N_4750,N_3920);
or U6662 (N_6662,N_2502,N_3173);
and U6663 (N_6663,N_4461,N_3430);
nor U6664 (N_6664,N_4191,N_3142);
nor U6665 (N_6665,N_3109,N_2929);
or U6666 (N_6666,N_3667,N_4267);
and U6667 (N_6667,N_4726,N_3269);
or U6668 (N_6668,N_2723,N_4058);
nor U6669 (N_6669,N_4050,N_2737);
nand U6670 (N_6670,N_2825,N_2945);
nor U6671 (N_6671,N_4226,N_3000);
or U6672 (N_6672,N_2978,N_2608);
nand U6673 (N_6673,N_2825,N_4854);
xor U6674 (N_6674,N_3138,N_2832);
and U6675 (N_6675,N_3684,N_4273);
nand U6676 (N_6676,N_3571,N_2628);
and U6677 (N_6677,N_4415,N_4257);
or U6678 (N_6678,N_3383,N_3275);
nor U6679 (N_6679,N_4162,N_3325);
or U6680 (N_6680,N_2568,N_3312);
nor U6681 (N_6681,N_4475,N_4400);
nor U6682 (N_6682,N_3172,N_2714);
nand U6683 (N_6683,N_4966,N_3757);
nor U6684 (N_6684,N_4994,N_3637);
nand U6685 (N_6685,N_3742,N_4445);
nor U6686 (N_6686,N_3709,N_2943);
nand U6687 (N_6687,N_4733,N_3836);
xor U6688 (N_6688,N_4901,N_4441);
nor U6689 (N_6689,N_4883,N_4467);
and U6690 (N_6690,N_4816,N_3524);
nor U6691 (N_6691,N_3332,N_3679);
or U6692 (N_6692,N_3623,N_4194);
nor U6693 (N_6693,N_3381,N_2560);
nor U6694 (N_6694,N_3802,N_4332);
nand U6695 (N_6695,N_3112,N_3107);
nor U6696 (N_6696,N_3093,N_3111);
nor U6697 (N_6697,N_4468,N_3571);
nor U6698 (N_6698,N_4141,N_3997);
nor U6699 (N_6699,N_4867,N_3768);
and U6700 (N_6700,N_4620,N_4701);
and U6701 (N_6701,N_4726,N_4497);
nor U6702 (N_6702,N_3851,N_3648);
nor U6703 (N_6703,N_2624,N_4833);
nor U6704 (N_6704,N_3955,N_4204);
nand U6705 (N_6705,N_4145,N_2649);
nor U6706 (N_6706,N_4566,N_2770);
nor U6707 (N_6707,N_3232,N_4950);
nand U6708 (N_6708,N_2710,N_3350);
nand U6709 (N_6709,N_3974,N_3031);
or U6710 (N_6710,N_4187,N_4348);
nor U6711 (N_6711,N_4974,N_4581);
nand U6712 (N_6712,N_3963,N_3598);
or U6713 (N_6713,N_2699,N_4221);
nand U6714 (N_6714,N_2601,N_3320);
or U6715 (N_6715,N_4771,N_4778);
nor U6716 (N_6716,N_3981,N_3810);
or U6717 (N_6717,N_4990,N_3776);
nand U6718 (N_6718,N_3050,N_3140);
nand U6719 (N_6719,N_3115,N_3369);
and U6720 (N_6720,N_4586,N_4416);
nand U6721 (N_6721,N_4469,N_3529);
and U6722 (N_6722,N_4969,N_3893);
and U6723 (N_6723,N_3856,N_3293);
or U6724 (N_6724,N_4397,N_3176);
and U6725 (N_6725,N_4968,N_2792);
and U6726 (N_6726,N_4524,N_3973);
or U6727 (N_6727,N_3818,N_2667);
nor U6728 (N_6728,N_2521,N_3343);
and U6729 (N_6729,N_4473,N_3750);
and U6730 (N_6730,N_2985,N_2839);
nor U6731 (N_6731,N_3778,N_3780);
nor U6732 (N_6732,N_3357,N_4997);
nor U6733 (N_6733,N_4564,N_2819);
and U6734 (N_6734,N_4506,N_3013);
or U6735 (N_6735,N_4380,N_2515);
nand U6736 (N_6736,N_3552,N_4551);
and U6737 (N_6737,N_4920,N_4127);
or U6738 (N_6738,N_4102,N_3009);
nor U6739 (N_6739,N_3202,N_3688);
nor U6740 (N_6740,N_4235,N_2519);
or U6741 (N_6741,N_3533,N_2856);
or U6742 (N_6742,N_3641,N_2837);
and U6743 (N_6743,N_3574,N_3984);
nor U6744 (N_6744,N_4354,N_4877);
nor U6745 (N_6745,N_3331,N_3901);
and U6746 (N_6746,N_3869,N_3757);
and U6747 (N_6747,N_2833,N_3676);
nand U6748 (N_6748,N_2679,N_3699);
nor U6749 (N_6749,N_3506,N_4992);
or U6750 (N_6750,N_3240,N_3871);
nor U6751 (N_6751,N_3206,N_3603);
nor U6752 (N_6752,N_3541,N_4906);
nor U6753 (N_6753,N_2806,N_4550);
nand U6754 (N_6754,N_3904,N_3044);
or U6755 (N_6755,N_3409,N_2626);
nor U6756 (N_6756,N_3448,N_2741);
nor U6757 (N_6757,N_3276,N_4931);
or U6758 (N_6758,N_4293,N_2931);
nor U6759 (N_6759,N_3021,N_4565);
or U6760 (N_6760,N_3648,N_4061);
xor U6761 (N_6761,N_4840,N_4820);
nand U6762 (N_6762,N_3961,N_4950);
nand U6763 (N_6763,N_2765,N_3379);
nand U6764 (N_6764,N_4148,N_3153);
or U6765 (N_6765,N_4210,N_3686);
nand U6766 (N_6766,N_2515,N_3207);
and U6767 (N_6767,N_4982,N_3257);
and U6768 (N_6768,N_3270,N_4792);
or U6769 (N_6769,N_3845,N_2550);
nor U6770 (N_6770,N_3319,N_3503);
nand U6771 (N_6771,N_2513,N_3883);
nor U6772 (N_6772,N_4029,N_4836);
nand U6773 (N_6773,N_3088,N_4761);
nor U6774 (N_6774,N_4179,N_2994);
and U6775 (N_6775,N_4517,N_3418);
and U6776 (N_6776,N_2795,N_3501);
nor U6777 (N_6777,N_2641,N_3487);
and U6778 (N_6778,N_3411,N_4161);
nand U6779 (N_6779,N_2984,N_2911);
or U6780 (N_6780,N_4112,N_4234);
nor U6781 (N_6781,N_3685,N_4521);
and U6782 (N_6782,N_4345,N_4848);
nor U6783 (N_6783,N_3665,N_4493);
nor U6784 (N_6784,N_4215,N_3510);
nor U6785 (N_6785,N_4447,N_3502);
and U6786 (N_6786,N_2667,N_2781);
nor U6787 (N_6787,N_4476,N_3113);
or U6788 (N_6788,N_4831,N_2601);
nor U6789 (N_6789,N_2979,N_4641);
nor U6790 (N_6790,N_4816,N_4906);
nand U6791 (N_6791,N_4958,N_2748);
nor U6792 (N_6792,N_2533,N_3382);
nand U6793 (N_6793,N_3100,N_2985);
nand U6794 (N_6794,N_4523,N_4721);
nor U6795 (N_6795,N_3497,N_4175);
nand U6796 (N_6796,N_4101,N_3333);
nand U6797 (N_6797,N_3887,N_2533);
nand U6798 (N_6798,N_3831,N_3402);
nand U6799 (N_6799,N_4845,N_4013);
nand U6800 (N_6800,N_4901,N_4363);
nand U6801 (N_6801,N_4805,N_3474);
nand U6802 (N_6802,N_2555,N_4627);
or U6803 (N_6803,N_2978,N_3834);
and U6804 (N_6804,N_4119,N_2715);
or U6805 (N_6805,N_3121,N_3314);
nor U6806 (N_6806,N_4539,N_2811);
nand U6807 (N_6807,N_4311,N_4966);
nand U6808 (N_6808,N_3650,N_4209);
nand U6809 (N_6809,N_3513,N_3201);
and U6810 (N_6810,N_4636,N_4279);
nor U6811 (N_6811,N_2548,N_4129);
nand U6812 (N_6812,N_4580,N_3385);
and U6813 (N_6813,N_3677,N_3722);
nor U6814 (N_6814,N_4455,N_3685);
and U6815 (N_6815,N_4257,N_3572);
nor U6816 (N_6816,N_3483,N_2745);
nor U6817 (N_6817,N_4722,N_4227);
and U6818 (N_6818,N_4162,N_4341);
and U6819 (N_6819,N_2906,N_3590);
or U6820 (N_6820,N_2577,N_4013);
nand U6821 (N_6821,N_4680,N_4461);
or U6822 (N_6822,N_4094,N_4636);
and U6823 (N_6823,N_2806,N_3398);
nand U6824 (N_6824,N_3715,N_4236);
nor U6825 (N_6825,N_2745,N_3745);
nor U6826 (N_6826,N_3100,N_2945);
and U6827 (N_6827,N_3862,N_3022);
and U6828 (N_6828,N_4781,N_3021);
nand U6829 (N_6829,N_3767,N_3699);
nor U6830 (N_6830,N_4607,N_3381);
xor U6831 (N_6831,N_4695,N_3954);
nor U6832 (N_6832,N_4679,N_2694);
nor U6833 (N_6833,N_2656,N_4891);
nand U6834 (N_6834,N_3656,N_4794);
nand U6835 (N_6835,N_2567,N_4205);
nand U6836 (N_6836,N_3297,N_4655);
and U6837 (N_6837,N_3800,N_4762);
nand U6838 (N_6838,N_4781,N_3525);
and U6839 (N_6839,N_4339,N_4464);
or U6840 (N_6840,N_3045,N_4259);
and U6841 (N_6841,N_4578,N_4275);
and U6842 (N_6842,N_2849,N_4786);
nand U6843 (N_6843,N_3557,N_4852);
nor U6844 (N_6844,N_4790,N_3452);
or U6845 (N_6845,N_3217,N_2666);
nor U6846 (N_6846,N_2807,N_2654);
nand U6847 (N_6847,N_4510,N_4241);
nor U6848 (N_6848,N_3389,N_2797);
nor U6849 (N_6849,N_2596,N_3597);
and U6850 (N_6850,N_2886,N_3244);
or U6851 (N_6851,N_4165,N_3649);
nand U6852 (N_6852,N_2826,N_4456);
nor U6853 (N_6853,N_3496,N_4266);
or U6854 (N_6854,N_3211,N_3186);
nor U6855 (N_6855,N_4336,N_2790);
and U6856 (N_6856,N_4387,N_2994);
nand U6857 (N_6857,N_3636,N_2907);
nor U6858 (N_6858,N_3308,N_3998);
or U6859 (N_6859,N_3659,N_3921);
and U6860 (N_6860,N_2752,N_4238);
nor U6861 (N_6861,N_3305,N_3688);
or U6862 (N_6862,N_4336,N_4125);
nor U6863 (N_6863,N_4648,N_2694);
xor U6864 (N_6864,N_4193,N_4390);
nand U6865 (N_6865,N_4486,N_4384);
nor U6866 (N_6866,N_4463,N_4331);
nand U6867 (N_6867,N_3651,N_4041);
and U6868 (N_6868,N_3528,N_2787);
nor U6869 (N_6869,N_3221,N_4585);
nor U6870 (N_6870,N_4476,N_3213);
nor U6871 (N_6871,N_3082,N_2567);
nand U6872 (N_6872,N_4342,N_3178);
xnor U6873 (N_6873,N_3470,N_4137);
and U6874 (N_6874,N_4203,N_4053);
or U6875 (N_6875,N_3452,N_4352);
nor U6876 (N_6876,N_4145,N_3786);
or U6877 (N_6877,N_3827,N_3580);
nor U6878 (N_6878,N_4956,N_3979);
nand U6879 (N_6879,N_4209,N_3904);
nand U6880 (N_6880,N_3905,N_4738);
nand U6881 (N_6881,N_4014,N_3178);
and U6882 (N_6882,N_3498,N_4529);
and U6883 (N_6883,N_3920,N_4353);
and U6884 (N_6884,N_3135,N_4276);
or U6885 (N_6885,N_3508,N_4698);
and U6886 (N_6886,N_4976,N_4189);
or U6887 (N_6887,N_2892,N_4866);
nor U6888 (N_6888,N_4855,N_4696);
nor U6889 (N_6889,N_3598,N_4883);
nor U6890 (N_6890,N_4383,N_3828);
or U6891 (N_6891,N_2872,N_2821);
nor U6892 (N_6892,N_4848,N_3398);
nor U6893 (N_6893,N_2932,N_3382);
and U6894 (N_6894,N_4742,N_4720);
nand U6895 (N_6895,N_2947,N_3102);
and U6896 (N_6896,N_2983,N_3068);
and U6897 (N_6897,N_2887,N_3484);
and U6898 (N_6898,N_2698,N_4109);
nor U6899 (N_6899,N_3055,N_3653);
nor U6900 (N_6900,N_3143,N_3152);
and U6901 (N_6901,N_4929,N_3160);
nand U6902 (N_6902,N_4579,N_4243);
nand U6903 (N_6903,N_4916,N_3083);
and U6904 (N_6904,N_2975,N_2864);
nand U6905 (N_6905,N_4814,N_2955);
nand U6906 (N_6906,N_3963,N_2677);
nand U6907 (N_6907,N_3394,N_2615);
and U6908 (N_6908,N_4603,N_4997);
and U6909 (N_6909,N_4169,N_2773);
nand U6910 (N_6910,N_3509,N_3070);
and U6911 (N_6911,N_4608,N_3152);
or U6912 (N_6912,N_3136,N_4340);
and U6913 (N_6913,N_4512,N_3712);
nor U6914 (N_6914,N_2749,N_3731);
or U6915 (N_6915,N_3913,N_3410);
nand U6916 (N_6916,N_4427,N_4981);
nor U6917 (N_6917,N_3724,N_2995);
and U6918 (N_6918,N_2515,N_4796);
or U6919 (N_6919,N_3330,N_2518);
or U6920 (N_6920,N_3923,N_3540);
nand U6921 (N_6921,N_3311,N_4374);
and U6922 (N_6922,N_3209,N_3066);
nor U6923 (N_6923,N_4565,N_4570);
nor U6924 (N_6924,N_2663,N_4017);
or U6925 (N_6925,N_3414,N_2620);
nor U6926 (N_6926,N_4348,N_2610);
nor U6927 (N_6927,N_3303,N_4484);
nor U6928 (N_6928,N_3566,N_3658);
nor U6929 (N_6929,N_3058,N_3567);
or U6930 (N_6930,N_4175,N_3047);
nor U6931 (N_6931,N_4217,N_3563);
and U6932 (N_6932,N_3834,N_4326);
and U6933 (N_6933,N_2989,N_4371);
nor U6934 (N_6934,N_2516,N_2858);
or U6935 (N_6935,N_3275,N_3191);
or U6936 (N_6936,N_3761,N_4104);
and U6937 (N_6937,N_4417,N_3219);
nand U6938 (N_6938,N_3116,N_4475);
or U6939 (N_6939,N_3339,N_3858);
or U6940 (N_6940,N_4172,N_3452);
and U6941 (N_6941,N_3253,N_2937);
nor U6942 (N_6942,N_2795,N_3925);
or U6943 (N_6943,N_4258,N_3911);
and U6944 (N_6944,N_3716,N_4594);
nor U6945 (N_6945,N_4567,N_4611);
nor U6946 (N_6946,N_4882,N_3063);
or U6947 (N_6947,N_3960,N_4264);
or U6948 (N_6948,N_3831,N_3239);
and U6949 (N_6949,N_3171,N_3493);
and U6950 (N_6950,N_4941,N_2641);
or U6951 (N_6951,N_2569,N_3958);
nand U6952 (N_6952,N_2560,N_2772);
and U6953 (N_6953,N_3853,N_3742);
and U6954 (N_6954,N_4349,N_2956);
and U6955 (N_6955,N_4673,N_3716);
nand U6956 (N_6956,N_2964,N_3216);
nor U6957 (N_6957,N_3183,N_4471);
or U6958 (N_6958,N_3149,N_3305);
nand U6959 (N_6959,N_4680,N_2862);
or U6960 (N_6960,N_3396,N_4148);
or U6961 (N_6961,N_4881,N_3100);
nor U6962 (N_6962,N_3609,N_3029);
and U6963 (N_6963,N_4219,N_2535);
xor U6964 (N_6964,N_3945,N_3542);
and U6965 (N_6965,N_3800,N_4826);
or U6966 (N_6966,N_3007,N_3934);
nand U6967 (N_6967,N_4951,N_3575);
and U6968 (N_6968,N_2569,N_3289);
and U6969 (N_6969,N_3811,N_4216);
or U6970 (N_6970,N_4603,N_4007);
and U6971 (N_6971,N_3695,N_3686);
nor U6972 (N_6972,N_2940,N_4992);
or U6973 (N_6973,N_4868,N_4585);
or U6974 (N_6974,N_3177,N_3633);
nand U6975 (N_6975,N_4239,N_4042);
and U6976 (N_6976,N_3999,N_3119);
and U6977 (N_6977,N_4813,N_3276);
nor U6978 (N_6978,N_4502,N_4654);
nand U6979 (N_6979,N_4382,N_4302);
and U6980 (N_6980,N_3424,N_4955);
nor U6981 (N_6981,N_3976,N_4861);
nand U6982 (N_6982,N_2617,N_4679);
nand U6983 (N_6983,N_3007,N_4796);
nand U6984 (N_6984,N_3493,N_3475);
or U6985 (N_6985,N_2519,N_4171);
nand U6986 (N_6986,N_4486,N_3096);
nor U6987 (N_6987,N_3042,N_3763);
and U6988 (N_6988,N_3658,N_3219);
nand U6989 (N_6989,N_2867,N_3275);
nor U6990 (N_6990,N_4699,N_4338);
and U6991 (N_6991,N_3072,N_2693);
and U6992 (N_6992,N_4270,N_3153);
nor U6993 (N_6993,N_3366,N_4388);
nand U6994 (N_6994,N_3293,N_2851);
nand U6995 (N_6995,N_3609,N_3186);
nand U6996 (N_6996,N_3985,N_3898);
nor U6997 (N_6997,N_3605,N_3508);
nand U6998 (N_6998,N_4629,N_2974);
nand U6999 (N_6999,N_4683,N_2751);
and U7000 (N_7000,N_3484,N_2719);
xnor U7001 (N_7001,N_3910,N_3434);
nor U7002 (N_7002,N_2931,N_2807);
or U7003 (N_7003,N_3891,N_4803);
and U7004 (N_7004,N_3360,N_2813);
or U7005 (N_7005,N_4534,N_4444);
and U7006 (N_7006,N_3326,N_4058);
or U7007 (N_7007,N_2867,N_4723);
and U7008 (N_7008,N_2989,N_3229);
nor U7009 (N_7009,N_2628,N_2595);
or U7010 (N_7010,N_2837,N_3686);
xor U7011 (N_7011,N_3209,N_3241);
nand U7012 (N_7012,N_3985,N_2823);
and U7013 (N_7013,N_2943,N_4988);
and U7014 (N_7014,N_2689,N_4892);
nor U7015 (N_7015,N_3615,N_3415);
nand U7016 (N_7016,N_4634,N_3447);
nand U7017 (N_7017,N_3900,N_4956);
or U7018 (N_7018,N_4976,N_2971);
nand U7019 (N_7019,N_3726,N_4935);
nand U7020 (N_7020,N_3479,N_4419);
and U7021 (N_7021,N_3599,N_4693);
and U7022 (N_7022,N_2895,N_2563);
nand U7023 (N_7023,N_3519,N_3860);
or U7024 (N_7024,N_3638,N_2881);
nand U7025 (N_7025,N_4358,N_3250);
nand U7026 (N_7026,N_4785,N_4440);
or U7027 (N_7027,N_2938,N_3063);
nand U7028 (N_7028,N_3651,N_4378);
or U7029 (N_7029,N_2678,N_3810);
or U7030 (N_7030,N_4815,N_4480);
nor U7031 (N_7031,N_2501,N_4353);
and U7032 (N_7032,N_2614,N_3202);
nand U7033 (N_7033,N_4785,N_2577);
and U7034 (N_7034,N_4367,N_4333);
nor U7035 (N_7035,N_3802,N_4245);
and U7036 (N_7036,N_3651,N_2819);
or U7037 (N_7037,N_4379,N_4338);
and U7038 (N_7038,N_4536,N_3257);
or U7039 (N_7039,N_3541,N_4423);
nand U7040 (N_7040,N_2947,N_3359);
nor U7041 (N_7041,N_3166,N_4411);
or U7042 (N_7042,N_3935,N_3970);
nor U7043 (N_7043,N_3443,N_4435);
nor U7044 (N_7044,N_3599,N_4390);
and U7045 (N_7045,N_4350,N_3698);
or U7046 (N_7046,N_4468,N_2692);
and U7047 (N_7047,N_3634,N_3868);
or U7048 (N_7048,N_3467,N_4260);
and U7049 (N_7049,N_2708,N_2844);
or U7050 (N_7050,N_2651,N_4417);
and U7051 (N_7051,N_2597,N_4293);
nor U7052 (N_7052,N_4338,N_4835);
nor U7053 (N_7053,N_3241,N_3337);
or U7054 (N_7054,N_4095,N_3397);
nand U7055 (N_7055,N_2601,N_3628);
or U7056 (N_7056,N_4282,N_4512);
and U7057 (N_7057,N_3195,N_4108);
nand U7058 (N_7058,N_3547,N_4225);
and U7059 (N_7059,N_3269,N_4605);
nand U7060 (N_7060,N_3285,N_2729);
nand U7061 (N_7061,N_3508,N_4767);
or U7062 (N_7062,N_3262,N_4472);
nor U7063 (N_7063,N_4910,N_3708);
nor U7064 (N_7064,N_3235,N_2687);
nor U7065 (N_7065,N_3797,N_4314);
nor U7066 (N_7066,N_3322,N_3214);
or U7067 (N_7067,N_4637,N_2593);
or U7068 (N_7068,N_4517,N_2636);
or U7069 (N_7069,N_4062,N_3063);
or U7070 (N_7070,N_4914,N_4949);
or U7071 (N_7071,N_3310,N_3577);
and U7072 (N_7072,N_4178,N_2921);
nor U7073 (N_7073,N_3229,N_3040);
and U7074 (N_7074,N_4380,N_4296);
or U7075 (N_7075,N_3867,N_4341);
nor U7076 (N_7076,N_3553,N_4860);
and U7077 (N_7077,N_4930,N_2905);
and U7078 (N_7078,N_2594,N_4514);
xor U7079 (N_7079,N_3865,N_3060);
nand U7080 (N_7080,N_3954,N_4849);
nand U7081 (N_7081,N_3527,N_4873);
nand U7082 (N_7082,N_2579,N_4785);
nor U7083 (N_7083,N_2745,N_2764);
nor U7084 (N_7084,N_4336,N_4294);
nor U7085 (N_7085,N_2544,N_3126);
nor U7086 (N_7086,N_3966,N_3973);
nor U7087 (N_7087,N_3224,N_4174);
xnor U7088 (N_7088,N_2840,N_3993);
nand U7089 (N_7089,N_3501,N_4152);
or U7090 (N_7090,N_4251,N_2865);
and U7091 (N_7091,N_4554,N_3896);
and U7092 (N_7092,N_3272,N_3048);
or U7093 (N_7093,N_3599,N_4863);
and U7094 (N_7094,N_3096,N_3959);
or U7095 (N_7095,N_3482,N_3563);
nor U7096 (N_7096,N_3253,N_2969);
nor U7097 (N_7097,N_2755,N_2663);
or U7098 (N_7098,N_4694,N_2830);
nand U7099 (N_7099,N_3570,N_3484);
nor U7100 (N_7100,N_3273,N_4579);
nor U7101 (N_7101,N_4444,N_4277);
nand U7102 (N_7102,N_4954,N_4107);
nor U7103 (N_7103,N_4394,N_2580);
and U7104 (N_7104,N_4839,N_2514);
xnor U7105 (N_7105,N_4678,N_4692);
or U7106 (N_7106,N_4560,N_3595);
and U7107 (N_7107,N_3499,N_3287);
and U7108 (N_7108,N_2748,N_2525);
or U7109 (N_7109,N_4189,N_3117);
and U7110 (N_7110,N_3964,N_4313);
and U7111 (N_7111,N_4840,N_3014);
or U7112 (N_7112,N_3855,N_4300);
nor U7113 (N_7113,N_4499,N_3375);
and U7114 (N_7114,N_4859,N_3424);
nor U7115 (N_7115,N_4605,N_2765);
nor U7116 (N_7116,N_4486,N_4044);
nand U7117 (N_7117,N_3688,N_4659);
and U7118 (N_7118,N_3937,N_3439);
or U7119 (N_7119,N_4691,N_3235);
nor U7120 (N_7120,N_3782,N_4233);
or U7121 (N_7121,N_4499,N_2804);
and U7122 (N_7122,N_3601,N_4057);
or U7123 (N_7123,N_3313,N_4074);
nand U7124 (N_7124,N_4306,N_3120);
nand U7125 (N_7125,N_4631,N_3634);
and U7126 (N_7126,N_3827,N_4407);
xnor U7127 (N_7127,N_3248,N_3882);
and U7128 (N_7128,N_4085,N_4196);
and U7129 (N_7129,N_2554,N_4780);
nand U7130 (N_7130,N_2808,N_4018);
and U7131 (N_7131,N_4792,N_2690);
nand U7132 (N_7132,N_4865,N_4839);
and U7133 (N_7133,N_3939,N_4457);
nor U7134 (N_7134,N_2533,N_3577);
and U7135 (N_7135,N_3784,N_2723);
nor U7136 (N_7136,N_4953,N_4179);
nor U7137 (N_7137,N_4719,N_3757);
nand U7138 (N_7138,N_4380,N_4334);
nor U7139 (N_7139,N_3416,N_2836);
and U7140 (N_7140,N_2766,N_3385);
nor U7141 (N_7141,N_2762,N_4290);
or U7142 (N_7142,N_3352,N_3935);
or U7143 (N_7143,N_4486,N_4707);
nor U7144 (N_7144,N_4157,N_2546);
and U7145 (N_7145,N_4385,N_2821);
and U7146 (N_7146,N_4485,N_4527);
xnor U7147 (N_7147,N_2822,N_3355);
or U7148 (N_7148,N_2794,N_2677);
nor U7149 (N_7149,N_3253,N_3221);
or U7150 (N_7150,N_4144,N_4774);
or U7151 (N_7151,N_3363,N_4688);
nand U7152 (N_7152,N_4193,N_3240);
or U7153 (N_7153,N_4269,N_3865);
nand U7154 (N_7154,N_4898,N_3760);
and U7155 (N_7155,N_2887,N_4949);
nand U7156 (N_7156,N_4203,N_3019);
and U7157 (N_7157,N_2902,N_4667);
and U7158 (N_7158,N_2590,N_3393);
nand U7159 (N_7159,N_4921,N_4823);
nor U7160 (N_7160,N_4392,N_4773);
or U7161 (N_7161,N_4198,N_2962);
nor U7162 (N_7162,N_4726,N_3243);
nand U7163 (N_7163,N_2739,N_4768);
or U7164 (N_7164,N_2721,N_4249);
nand U7165 (N_7165,N_4185,N_3710);
nand U7166 (N_7166,N_2514,N_3436);
and U7167 (N_7167,N_2532,N_2615);
or U7168 (N_7168,N_4669,N_3380);
and U7169 (N_7169,N_3939,N_3421);
or U7170 (N_7170,N_2846,N_4220);
or U7171 (N_7171,N_3344,N_2847);
or U7172 (N_7172,N_3947,N_3419);
and U7173 (N_7173,N_4368,N_2606);
nor U7174 (N_7174,N_4169,N_4699);
nand U7175 (N_7175,N_3854,N_3700);
and U7176 (N_7176,N_4358,N_2608);
or U7177 (N_7177,N_3321,N_2837);
and U7178 (N_7178,N_4757,N_3984);
nand U7179 (N_7179,N_3238,N_4026);
nand U7180 (N_7180,N_2652,N_2526);
nor U7181 (N_7181,N_4820,N_4699);
or U7182 (N_7182,N_2518,N_4605);
nor U7183 (N_7183,N_3489,N_2801);
nor U7184 (N_7184,N_4911,N_2770);
nand U7185 (N_7185,N_3265,N_4589);
or U7186 (N_7186,N_4864,N_4079);
nor U7187 (N_7187,N_3311,N_3753);
or U7188 (N_7188,N_4264,N_3384);
nor U7189 (N_7189,N_3809,N_4000);
and U7190 (N_7190,N_4582,N_4417);
and U7191 (N_7191,N_3912,N_4158);
or U7192 (N_7192,N_3241,N_3307);
or U7193 (N_7193,N_4331,N_4468);
nand U7194 (N_7194,N_3646,N_2615);
and U7195 (N_7195,N_2635,N_4652);
and U7196 (N_7196,N_4819,N_3296);
nor U7197 (N_7197,N_4287,N_3653);
nand U7198 (N_7198,N_3612,N_2555);
or U7199 (N_7199,N_3162,N_3259);
nor U7200 (N_7200,N_4047,N_3677);
and U7201 (N_7201,N_3857,N_4452);
nand U7202 (N_7202,N_3963,N_3951);
nand U7203 (N_7203,N_3600,N_4560);
nor U7204 (N_7204,N_3774,N_2783);
nand U7205 (N_7205,N_3128,N_4379);
and U7206 (N_7206,N_2797,N_4624);
nand U7207 (N_7207,N_3888,N_4003);
nand U7208 (N_7208,N_3823,N_3918);
nor U7209 (N_7209,N_4497,N_3011);
or U7210 (N_7210,N_3873,N_4524);
nor U7211 (N_7211,N_3884,N_4653);
or U7212 (N_7212,N_3101,N_3301);
and U7213 (N_7213,N_4478,N_2657);
and U7214 (N_7214,N_2529,N_4331);
nand U7215 (N_7215,N_3050,N_2516);
nand U7216 (N_7216,N_3992,N_3284);
nor U7217 (N_7217,N_3796,N_3910);
and U7218 (N_7218,N_4340,N_4632);
or U7219 (N_7219,N_2767,N_2944);
or U7220 (N_7220,N_2811,N_3481);
or U7221 (N_7221,N_2758,N_4305);
or U7222 (N_7222,N_4159,N_4609);
and U7223 (N_7223,N_4668,N_3143);
and U7224 (N_7224,N_3284,N_3121);
nor U7225 (N_7225,N_3968,N_3617);
nand U7226 (N_7226,N_2590,N_4065);
or U7227 (N_7227,N_3145,N_3567);
nand U7228 (N_7228,N_2585,N_4225);
or U7229 (N_7229,N_4061,N_3959);
nor U7230 (N_7230,N_4311,N_3921);
and U7231 (N_7231,N_3474,N_4772);
and U7232 (N_7232,N_4294,N_3541);
nand U7233 (N_7233,N_2573,N_3381);
nor U7234 (N_7234,N_4188,N_4321);
or U7235 (N_7235,N_3788,N_4448);
nor U7236 (N_7236,N_4126,N_3324);
nor U7237 (N_7237,N_3541,N_3781);
or U7238 (N_7238,N_4960,N_4073);
and U7239 (N_7239,N_2538,N_3951);
and U7240 (N_7240,N_4978,N_3873);
or U7241 (N_7241,N_3135,N_3750);
or U7242 (N_7242,N_3896,N_3511);
or U7243 (N_7243,N_4368,N_4056);
nor U7244 (N_7244,N_3015,N_4272);
nand U7245 (N_7245,N_4526,N_3404);
nand U7246 (N_7246,N_3050,N_3083);
nor U7247 (N_7247,N_3122,N_3370);
or U7248 (N_7248,N_2939,N_4817);
nor U7249 (N_7249,N_4451,N_4278);
nand U7250 (N_7250,N_2775,N_4641);
xor U7251 (N_7251,N_4785,N_4095);
or U7252 (N_7252,N_3130,N_3873);
or U7253 (N_7253,N_3724,N_3780);
nand U7254 (N_7254,N_4049,N_4323);
or U7255 (N_7255,N_2785,N_4383);
and U7256 (N_7256,N_2758,N_2581);
and U7257 (N_7257,N_3019,N_3686);
nand U7258 (N_7258,N_4669,N_3759);
or U7259 (N_7259,N_3457,N_4708);
and U7260 (N_7260,N_3139,N_3069);
and U7261 (N_7261,N_3613,N_4570);
nand U7262 (N_7262,N_3669,N_2874);
and U7263 (N_7263,N_2740,N_4541);
and U7264 (N_7264,N_4169,N_3907);
nand U7265 (N_7265,N_2674,N_4419);
nand U7266 (N_7266,N_4714,N_2965);
or U7267 (N_7267,N_4919,N_2561);
nand U7268 (N_7268,N_3103,N_2630);
and U7269 (N_7269,N_2837,N_4591);
nand U7270 (N_7270,N_4837,N_4482);
or U7271 (N_7271,N_3767,N_3240);
nand U7272 (N_7272,N_2767,N_2550);
nand U7273 (N_7273,N_3913,N_2640);
nand U7274 (N_7274,N_4847,N_3676);
nor U7275 (N_7275,N_4277,N_3118);
and U7276 (N_7276,N_4686,N_3789);
and U7277 (N_7277,N_4693,N_3848);
nor U7278 (N_7278,N_3425,N_3973);
nor U7279 (N_7279,N_2563,N_4105);
and U7280 (N_7280,N_4596,N_4277);
or U7281 (N_7281,N_4335,N_4512);
and U7282 (N_7282,N_4196,N_3395);
and U7283 (N_7283,N_2654,N_4200);
nor U7284 (N_7284,N_3605,N_4593);
or U7285 (N_7285,N_4370,N_2707);
and U7286 (N_7286,N_4591,N_3932);
nand U7287 (N_7287,N_3733,N_3521);
nor U7288 (N_7288,N_3229,N_3162);
and U7289 (N_7289,N_3349,N_4842);
nand U7290 (N_7290,N_2602,N_4628);
nand U7291 (N_7291,N_3115,N_2682);
and U7292 (N_7292,N_4629,N_3395);
nor U7293 (N_7293,N_3907,N_3387);
or U7294 (N_7294,N_2506,N_2818);
and U7295 (N_7295,N_4643,N_3474);
and U7296 (N_7296,N_3357,N_3821);
or U7297 (N_7297,N_2561,N_4490);
and U7298 (N_7298,N_4782,N_2860);
or U7299 (N_7299,N_2813,N_4714);
and U7300 (N_7300,N_3032,N_4972);
or U7301 (N_7301,N_3615,N_4365);
and U7302 (N_7302,N_3260,N_4951);
nor U7303 (N_7303,N_4039,N_4502);
and U7304 (N_7304,N_2808,N_3182);
nor U7305 (N_7305,N_3805,N_4137);
and U7306 (N_7306,N_3581,N_2663);
or U7307 (N_7307,N_3099,N_4069);
nand U7308 (N_7308,N_3986,N_4683);
or U7309 (N_7309,N_3858,N_3922);
or U7310 (N_7310,N_4558,N_2733);
and U7311 (N_7311,N_2773,N_3200);
nor U7312 (N_7312,N_3394,N_4998);
nor U7313 (N_7313,N_4731,N_4621);
nor U7314 (N_7314,N_2546,N_2864);
nand U7315 (N_7315,N_3637,N_3892);
or U7316 (N_7316,N_2825,N_4572);
nor U7317 (N_7317,N_4268,N_3830);
nor U7318 (N_7318,N_2806,N_4998);
and U7319 (N_7319,N_2684,N_2906);
and U7320 (N_7320,N_3752,N_3561);
nor U7321 (N_7321,N_3511,N_4805);
nand U7322 (N_7322,N_3205,N_4644);
or U7323 (N_7323,N_3045,N_4171);
xnor U7324 (N_7324,N_2773,N_2618);
or U7325 (N_7325,N_4226,N_4146);
or U7326 (N_7326,N_3564,N_3145);
nand U7327 (N_7327,N_4773,N_3003);
nand U7328 (N_7328,N_4718,N_3028);
nand U7329 (N_7329,N_4253,N_2595);
nor U7330 (N_7330,N_3555,N_2933);
nand U7331 (N_7331,N_3690,N_3160);
nor U7332 (N_7332,N_4666,N_4026);
nand U7333 (N_7333,N_3013,N_4906);
nand U7334 (N_7334,N_3304,N_3990);
nand U7335 (N_7335,N_3013,N_3716);
or U7336 (N_7336,N_3706,N_3377);
nor U7337 (N_7337,N_2840,N_4932);
or U7338 (N_7338,N_3709,N_4545);
nand U7339 (N_7339,N_4784,N_4092);
or U7340 (N_7340,N_3705,N_4094);
nand U7341 (N_7341,N_2509,N_4732);
nor U7342 (N_7342,N_4705,N_4273);
nand U7343 (N_7343,N_3031,N_4805);
nand U7344 (N_7344,N_3551,N_3967);
nand U7345 (N_7345,N_2663,N_4141);
nor U7346 (N_7346,N_4664,N_3634);
nand U7347 (N_7347,N_4249,N_3106);
nor U7348 (N_7348,N_3708,N_4410);
nand U7349 (N_7349,N_4387,N_2842);
nand U7350 (N_7350,N_2626,N_4822);
nor U7351 (N_7351,N_3513,N_4157);
and U7352 (N_7352,N_3313,N_3489);
or U7353 (N_7353,N_2836,N_3523);
nor U7354 (N_7354,N_3793,N_2887);
nor U7355 (N_7355,N_3525,N_2551);
and U7356 (N_7356,N_4708,N_4206);
nor U7357 (N_7357,N_4418,N_4679);
nand U7358 (N_7358,N_4341,N_4355);
and U7359 (N_7359,N_2609,N_2934);
nand U7360 (N_7360,N_3518,N_2948);
nand U7361 (N_7361,N_4516,N_2882);
nand U7362 (N_7362,N_3494,N_3414);
or U7363 (N_7363,N_3936,N_4056);
nor U7364 (N_7364,N_3196,N_3160);
or U7365 (N_7365,N_4773,N_2986);
nor U7366 (N_7366,N_4406,N_4892);
nand U7367 (N_7367,N_2528,N_3408);
or U7368 (N_7368,N_2984,N_3721);
nand U7369 (N_7369,N_4199,N_2596);
or U7370 (N_7370,N_3311,N_4760);
and U7371 (N_7371,N_2792,N_4778);
and U7372 (N_7372,N_2601,N_3930);
and U7373 (N_7373,N_3449,N_4519);
nor U7374 (N_7374,N_2546,N_3115);
nor U7375 (N_7375,N_4320,N_2565);
nand U7376 (N_7376,N_3996,N_3056);
nand U7377 (N_7377,N_4162,N_4403);
nor U7378 (N_7378,N_2639,N_3815);
or U7379 (N_7379,N_2696,N_2729);
nor U7380 (N_7380,N_4037,N_4007);
nand U7381 (N_7381,N_4217,N_4278);
or U7382 (N_7382,N_4116,N_2581);
nor U7383 (N_7383,N_2574,N_4679);
and U7384 (N_7384,N_3311,N_4517);
and U7385 (N_7385,N_3275,N_2550);
or U7386 (N_7386,N_4659,N_4274);
nand U7387 (N_7387,N_2879,N_3053);
or U7388 (N_7388,N_2871,N_4882);
nand U7389 (N_7389,N_3208,N_3073);
nand U7390 (N_7390,N_4241,N_3572);
and U7391 (N_7391,N_2814,N_3764);
and U7392 (N_7392,N_3400,N_2593);
or U7393 (N_7393,N_4189,N_2936);
and U7394 (N_7394,N_3119,N_3091);
nor U7395 (N_7395,N_4575,N_3221);
or U7396 (N_7396,N_3097,N_3394);
nor U7397 (N_7397,N_4161,N_4677);
nand U7398 (N_7398,N_2768,N_3973);
and U7399 (N_7399,N_2593,N_2878);
nand U7400 (N_7400,N_4234,N_4249);
or U7401 (N_7401,N_4243,N_4003);
or U7402 (N_7402,N_4535,N_3281);
or U7403 (N_7403,N_4827,N_3255);
and U7404 (N_7404,N_3447,N_4573);
nor U7405 (N_7405,N_2597,N_2926);
and U7406 (N_7406,N_3987,N_3526);
or U7407 (N_7407,N_4256,N_3262);
nor U7408 (N_7408,N_2666,N_3443);
nor U7409 (N_7409,N_3392,N_3249);
nand U7410 (N_7410,N_4407,N_4351);
and U7411 (N_7411,N_3208,N_4095);
or U7412 (N_7412,N_2939,N_2691);
nand U7413 (N_7413,N_4241,N_3465);
nand U7414 (N_7414,N_2610,N_3941);
nand U7415 (N_7415,N_4308,N_3670);
and U7416 (N_7416,N_3698,N_4574);
nor U7417 (N_7417,N_3659,N_4154);
and U7418 (N_7418,N_3293,N_4190);
or U7419 (N_7419,N_3904,N_3401);
or U7420 (N_7420,N_4152,N_2733);
nor U7421 (N_7421,N_3437,N_4103);
nor U7422 (N_7422,N_4339,N_4946);
nand U7423 (N_7423,N_3655,N_3428);
nand U7424 (N_7424,N_3184,N_3210);
nand U7425 (N_7425,N_4719,N_2535);
or U7426 (N_7426,N_3433,N_2591);
nand U7427 (N_7427,N_3852,N_3215);
and U7428 (N_7428,N_2527,N_4673);
nor U7429 (N_7429,N_4629,N_4376);
and U7430 (N_7430,N_2690,N_3570);
nand U7431 (N_7431,N_4197,N_3825);
and U7432 (N_7432,N_4527,N_4417);
or U7433 (N_7433,N_4731,N_2991);
nor U7434 (N_7434,N_4324,N_2894);
or U7435 (N_7435,N_4769,N_3787);
or U7436 (N_7436,N_3662,N_4566);
and U7437 (N_7437,N_4559,N_2615);
and U7438 (N_7438,N_2591,N_2989);
or U7439 (N_7439,N_2532,N_3749);
and U7440 (N_7440,N_3264,N_4673);
or U7441 (N_7441,N_4386,N_2552);
and U7442 (N_7442,N_3654,N_3079);
nand U7443 (N_7443,N_4926,N_3687);
and U7444 (N_7444,N_2647,N_3124);
and U7445 (N_7445,N_3121,N_3187);
and U7446 (N_7446,N_4967,N_3984);
nand U7447 (N_7447,N_4387,N_2685);
and U7448 (N_7448,N_4167,N_4813);
and U7449 (N_7449,N_3958,N_4333);
nor U7450 (N_7450,N_2525,N_3378);
and U7451 (N_7451,N_4095,N_4832);
or U7452 (N_7452,N_4969,N_3874);
nand U7453 (N_7453,N_4249,N_3330);
nor U7454 (N_7454,N_2813,N_2532);
or U7455 (N_7455,N_4896,N_3218);
nand U7456 (N_7456,N_3243,N_4076);
and U7457 (N_7457,N_4661,N_2741);
or U7458 (N_7458,N_3770,N_3930);
nand U7459 (N_7459,N_4984,N_2904);
nor U7460 (N_7460,N_4146,N_4933);
nor U7461 (N_7461,N_4311,N_2600);
or U7462 (N_7462,N_4275,N_4599);
or U7463 (N_7463,N_4030,N_4745);
nand U7464 (N_7464,N_3886,N_4260);
and U7465 (N_7465,N_3600,N_4138);
and U7466 (N_7466,N_3762,N_3903);
or U7467 (N_7467,N_3262,N_3366);
or U7468 (N_7468,N_2550,N_4461);
nand U7469 (N_7469,N_3775,N_3502);
and U7470 (N_7470,N_2695,N_2917);
and U7471 (N_7471,N_4255,N_4181);
or U7472 (N_7472,N_2799,N_3429);
nor U7473 (N_7473,N_4907,N_3030);
and U7474 (N_7474,N_4641,N_4703);
or U7475 (N_7475,N_4407,N_4574);
or U7476 (N_7476,N_3055,N_4135);
and U7477 (N_7477,N_4591,N_2926);
nand U7478 (N_7478,N_3144,N_4148);
or U7479 (N_7479,N_3065,N_2987);
and U7480 (N_7480,N_2746,N_3329);
nand U7481 (N_7481,N_3302,N_2915);
nand U7482 (N_7482,N_4971,N_4998);
nor U7483 (N_7483,N_3385,N_4703);
or U7484 (N_7484,N_2706,N_4655);
and U7485 (N_7485,N_3258,N_4389);
and U7486 (N_7486,N_2827,N_2872);
or U7487 (N_7487,N_2885,N_3809);
or U7488 (N_7488,N_2587,N_2904);
xnor U7489 (N_7489,N_3893,N_4173);
or U7490 (N_7490,N_4226,N_3263);
nor U7491 (N_7491,N_3722,N_3752);
nand U7492 (N_7492,N_4621,N_2975);
nor U7493 (N_7493,N_2616,N_2972);
nand U7494 (N_7494,N_4984,N_4187);
nor U7495 (N_7495,N_4157,N_4026);
or U7496 (N_7496,N_3651,N_2911);
nor U7497 (N_7497,N_4433,N_4284);
and U7498 (N_7498,N_3326,N_2690);
xor U7499 (N_7499,N_2729,N_4681);
and U7500 (N_7500,N_5360,N_6888);
nand U7501 (N_7501,N_6188,N_5441);
and U7502 (N_7502,N_6919,N_6117);
or U7503 (N_7503,N_7015,N_5781);
and U7504 (N_7504,N_6741,N_7317);
nor U7505 (N_7505,N_5334,N_6957);
or U7506 (N_7506,N_6271,N_6149);
nor U7507 (N_7507,N_5969,N_5159);
or U7508 (N_7508,N_6799,N_6296);
nand U7509 (N_7509,N_6399,N_5089);
nand U7510 (N_7510,N_6776,N_6407);
or U7511 (N_7511,N_6406,N_5020);
nand U7512 (N_7512,N_6718,N_6381);
nand U7513 (N_7513,N_7463,N_5099);
and U7514 (N_7514,N_7452,N_6508);
and U7515 (N_7515,N_6654,N_5551);
or U7516 (N_7516,N_7343,N_7323);
nor U7517 (N_7517,N_5478,N_6600);
and U7518 (N_7518,N_5405,N_5784);
or U7519 (N_7519,N_7217,N_6275);
nand U7520 (N_7520,N_7035,N_6802);
nand U7521 (N_7521,N_5297,N_6861);
nor U7522 (N_7522,N_6205,N_6754);
or U7523 (N_7523,N_6092,N_6766);
or U7524 (N_7524,N_7387,N_5131);
xnor U7525 (N_7525,N_7451,N_6518);
or U7526 (N_7526,N_5510,N_6962);
nand U7527 (N_7527,N_7489,N_5892);
or U7528 (N_7528,N_6926,N_6783);
xnor U7529 (N_7529,N_7213,N_5101);
and U7530 (N_7530,N_5536,N_5746);
nor U7531 (N_7531,N_6862,N_6699);
or U7532 (N_7532,N_5030,N_6071);
and U7533 (N_7533,N_6915,N_5212);
nor U7534 (N_7534,N_7426,N_6476);
and U7535 (N_7535,N_6881,N_7047);
and U7536 (N_7536,N_7245,N_7469);
and U7537 (N_7537,N_5198,N_5028);
or U7538 (N_7538,N_6498,N_5715);
or U7539 (N_7539,N_5565,N_6527);
and U7540 (N_7540,N_5820,N_6429);
nor U7541 (N_7541,N_7432,N_6907);
nor U7542 (N_7542,N_7382,N_6686);
nor U7543 (N_7543,N_7383,N_5581);
and U7544 (N_7544,N_6025,N_6836);
nand U7545 (N_7545,N_6289,N_5435);
or U7546 (N_7546,N_5262,N_7362);
nor U7547 (N_7547,N_5883,N_7214);
nor U7548 (N_7548,N_7110,N_6528);
and U7549 (N_7549,N_7369,N_5514);
nand U7550 (N_7550,N_5224,N_6769);
and U7551 (N_7551,N_6450,N_7385);
nand U7552 (N_7552,N_7099,N_7365);
nor U7553 (N_7553,N_5677,N_6300);
or U7554 (N_7554,N_5366,N_5719);
or U7555 (N_7555,N_6930,N_7439);
and U7556 (N_7556,N_6049,N_6577);
nand U7557 (N_7557,N_5307,N_5049);
nor U7558 (N_7558,N_6259,N_6107);
and U7559 (N_7559,N_5091,N_6545);
nand U7560 (N_7560,N_6648,N_5445);
nand U7561 (N_7561,N_5525,N_5359);
nor U7562 (N_7562,N_5233,N_6257);
nor U7563 (N_7563,N_6212,N_5523);
xor U7564 (N_7564,N_5162,N_7078);
nor U7565 (N_7565,N_5472,N_5662);
nor U7566 (N_7566,N_5109,N_5838);
or U7567 (N_7567,N_5817,N_6288);
nor U7568 (N_7568,N_6520,N_7253);
nand U7569 (N_7569,N_5379,N_5696);
nor U7570 (N_7570,N_5807,N_5654);
nor U7571 (N_7571,N_6727,N_6878);
or U7572 (N_7572,N_7422,N_5544);
and U7573 (N_7573,N_5084,N_5929);
and U7574 (N_7574,N_6643,N_6671);
and U7575 (N_7575,N_5306,N_5195);
nor U7576 (N_7576,N_7325,N_5680);
nor U7577 (N_7577,N_6869,N_5736);
nand U7578 (N_7578,N_6100,N_6094);
or U7579 (N_7579,N_5163,N_5216);
nor U7580 (N_7580,N_5701,N_5246);
or U7581 (N_7581,N_7416,N_7410);
nor U7582 (N_7582,N_7315,N_5583);
and U7583 (N_7583,N_6142,N_5596);
nand U7584 (N_7584,N_6052,N_5710);
nand U7585 (N_7585,N_6831,N_5970);
and U7586 (N_7586,N_5376,N_5505);
nand U7587 (N_7587,N_6599,N_5175);
or U7588 (N_7588,N_7468,N_6183);
nand U7589 (N_7589,N_5661,N_6765);
nand U7590 (N_7590,N_6085,N_6088);
xor U7591 (N_7591,N_6101,N_6298);
or U7592 (N_7592,N_6646,N_6917);
nor U7593 (N_7593,N_6041,N_5403);
nand U7594 (N_7594,N_5646,N_6638);
nor U7595 (N_7595,N_5954,N_7311);
nand U7596 (N_7596,N_5862,N_5672);
or U7597 (N_7597,N_5380,N_7005);
and U7598 (N_7598,N_6375,N_5276);
and U7599 (N_7599,N_6361,N_6390);
and U7600 (N_7600,N_5322,N_6285);
nand U7601 (N_7601,N_5716,N_5941);
or U7602 (N_7602,N_5870,N_6369);
or U7603 (N_7603,N_6291,N_6224);
or U7604 (N_7604,N_7490,N_6204);
nor U7605 (N_7605,N_6416,N_6753);
nor U7606 (N_7606,N_6672,N_7273);
or U7607 (N_7607,N_6384,N_5595);
nor U7608 (N_7608,N_7310,N_6093);
nand U7609 (N_7609,N_5888,N_7073);
and U7610 (N_7610,N_6113,N_6689);
nor U7611 (N_7611,N_5465,N_6811);
and U7612 (N_7612,N_5760,N_5125);
nor U7613 (N_7613,N_6480,N_6504);
or U7614 (N_7614,N_5190,N_5401);
nand U7615 (N_7615,N_6095,N_5408);
nor U7616 (N_7616,N_7384,N_6295);
and U7617 (N_7617,N_7093,N_6303);
nand U7618 (N_7618,N_6922,N_6220);
nor U7619 (N_7619,N_6155,N_5873);
nand U7620 (N_7620,N_5563,N_7006);
nor U7621 (N_7621,N_5168,N_6346);
and U7622 (N_7622,N_6465,N_5913);
nor U7623 (N_7623,N_7037,N_6372);
and U7624 (N_7624,N_5210,N_6377);
nand U7625 (N_7625,N_6552,N_6758);
nand U7626 (N_7626,N_6780,N_5787);
and U7627 (N_7627,N_5147,N_6002);
or U7628 (N_7628,N_6939,N_5001);
and U7629 (N_7629,N_7464,N_6409);
and U7630 (N_7630,N_5768,N_5013);
nor U7631 (N_7631,N_6130,N_6510);
nor U7632 (N_7632,N_6236,N_5587);
and U7633 (N_7633,N_6421,N_6326);
nand U7634 (N_7634,N_7041,N_6162);
nor U7635 (N_7635,N_5777,N_7212);
nor U7636 (N_7636,N_5763,N_6873);
and U7637 (N_7637,N_6124,N_7004);
nor U7638 (N_7638,N_5464,N_6268);
nand U7639 (N_7639,N_5278,N_6311);
nor U7640 (N_7640,N_6830,N_5118);
nor U7641 (N_7641,N_5902,N_5676);
nor U7642 (N_7642,N_5610,N_6229);
nor U7643 (N_7643,N_5048,N_7431);
or U7644 (N_7644,N_6637,N_7318);
nor U7645 (N_7645,N_5113,N_6357);
nand U7646 (N_7646,N_5062,N_7061);
or U7647 (N_7647,N_6193,N_7351);
and U7648 (N_7648,N_6234,N_6437);
nand U7649 (N_7649,N_6609,N_6075);
nor U7650 (N_7650,N_7062,N_6458);
nand U7651 (N_7651,N_6854,N_5729);
or U7652 (N_7652,N_6573,N_6173);
nand U7653 (N_7653,N_6143,N_6323);
or U7654 (N_7654,N_6281,N_6354);
nor U7655 (N_7655,N_6422,N_6106);
nand U7656 (N_7656,N_5259,N_6099);
nor U7657 (N_7657,N_5429,N_7491);
nor U7658 (N_7658,N_5611,N_5200);
and U7659 (N_7659,N_5882,N_5880);
and U7660 (N_7660,N_6687,N_6876);
nor U7661 (N_7661,N_5766,N_5406);
and U7662 (N_7662,N_5957,N_6233);
or U7663 (N_7663,N_7207,N_5891);
nor U7664 (N_7664,N_5274,N_6807);
nand U7665 (N_7665,N_5151,N_6969);
nor U7666 (N_7666,N_6729,N_5364);
or U7667 (N_7667,N_6161,N_6994);
nand U7668 (N_7668,N_7172,N_6184);
and U7669 (N_7669,N_7086,N_5384);
nand U7670 (N_7670,N_6841,N_5998);
nand U7671 (N_7671,N_5456,N_6277);
nor U7672 (N_7672,N_7268,N_7444);
and U7673 (N_7673,N_5263,N_5064);
or U7674 (N_7674,N_6096,N_6808);
and U7675 (N_7675,N_7412,N_6440);
nand U7676 (N_7676,N_5327,N_6290);
nand U7677 (N_7677,N_6227,N_5112);
nor U7678 (N_7678,N_6519,N_5219);
or U7679 (N_7679,N_5675,N_7085);
nand U7680 (N_7680,N_6078,N_6514);
nor U7681 (N_7681,N_7329,N_6970);
nor U7682 (N_7682,N_6571,N_6984);
or U7683 (N_7683,N_5556,N_5493);
or U7684 (N_7684,N_6832,N_5819);
nor U7685 (N_7685,N_7406,N_6089);
and U7686 (N_7686,N_6287,N_5252);
nor U7687 (N_7687,N_5744,N_5180);
or U7688 (N_7688,N_7413,N_7151);
nor U7689 (N_7689,N_6985,N_5318);
and U7690 (N_7690,N_5721,N_6951);
nand U7691 (N_7691,N_7333,N_6713);
and U7692 (N_7692,N_5548,N_5197);
or U7693 (N_7693,N_6840,N_5336);
nand U7694 (N_7694,N_5330,N_6669);
or U7695 (N_7695,N_6091,N_5031);
and U7696 (N_7696,N_6180,N_7056);
or U7697 (N_7697,N_5560,N_5457);
or U7698 (N_7698,N_6859,N_6104);
or U7699 (N_7699,N_6006,N_5841);
and U7700 (N_7700,N_6252,N_5280);
and U7701 (N_7701,N_5698,N_7097);
and U7702 (N_7702,N_7033,N_5177);
nor U7703 (N_7703,N_7316,N_5966);
nand U7704 (N_7704,N_6114,N_7197);
or U7705 (N_7705,N_7157,N_7359);
nor U7706 (N_7706,N_5962,N_5215);
and U7707 (N_7707,N_5847,N_5628);
nor U7708 (N_7708,N_5973,N_7026);
nor U7709 (N_7709,N_5533,N_7155);
or U7710 (N_7710,N_5114,N_5461);
nor U7711 (N_7711,N_6209,N_6884);
and U7712 (N_7712,N_6568,N_6007);
nor U7713 (N_7713,N_7052,N_7448);
nor U7714 (N_7714,N_6054,N_5550);
and U7715 (N_7715,N_7427,N_6011);
or U7716 (N_7716,N_7358,N_7462);
or U7717 (N_7717,N_6339,N_5779);
nand U7718 (N_7718,N_6784,N_7152);
nand U7719 (N_7719,N_6431,N_7265);
or U7720 (N_7720,N_5639,N_5642);
nand U7721 (N_7721,N_6097,N_6855);
nand U7722 (N_7722,N_7081,N_5846);
and U7723 (N_7723,N_5050,N_6594);
or U7724 (N_7724,N_7119,N_6653);
nor U7725 (N_7725,N_5810,N_5019);
nor U7726 (N_7726,N_6292,N_6785);
and U7727 (N_7727,N_6256,N_6449);
nand U7728 (N_7728,N_5617,N_7044);
nand U7729 (N_7729,N_5221,N_7084);
nor U7730 (N_7730,N_5585,N_5124);
nor U7731 (N_7731,N_7092,N_6787);
or U7732 (N_7732,N_5358,N_5409);
and U7733 (N_7733,N_5727,N_5886);
nand U7734 (N_7734,N_5612,N_7189);
nor U7735 (N_7735,N_6214,N_5607);
and U7736 (N_7736,N_5992,N_5993);
and U7737 (N_7737,N_5723,N_6507);
nand U7738 (N_7738,N_7367,N_6650);
and U7739 (N_7739,N_6631,N_7190);
nor U7740 (N_7740,N_6613,N_5349);
nand U7741 (N_7741,N_7294,N_5265);
nand U7742 (N_7742,N_5598,N_6263);
and U7743 (N_7743,N_7372,N_6196);
nor U7744 (N_7744,N_6363,N_6283);
nor U7745 (N_7745,N_7461,N_7205);
nor U7746 (N_7746,N_5632,N_5561);
or U7747 (N_7747,N_6477,N_7336);
nor U7748 (N_7748,N_5440,N_6265);
nand U7749 (N_7749,N_5343,N_5641);
and U7750 (N_7750,N_5059,N_5378);
nand U7751 (N_7751,N_5622,N_6316);
and U7752 (N_7752,N_5910,N_6742);
nand U7753 (N_7753,N_5105,N_5389);
or U7754 (N_7754,N_7058,N_6387);
nor U7755 (N_7755,N_6417,N_5485);
nand U7756 (N_7756,N_6560,N_6066);
or U7757 (N_7757,N_5293,N_5712);
or U7758 (N_7758,N_6745,N_7171);
nand U7759 (N_7759,N_6062,N_6353);
or U7760 (N_7760,N_5039,N_7445);
or U7761 (N_7761,N_7378,N_5305);
nor U7762 (N_7762,N_5481,N_7342);
nand U7763 (N_7763,N_5931,N_6175);
or U7764 (N_7764,N_6222,N_6358);
or U7765 (N_7765,N_6176,N_6691);
and U7766 (N_7766,N_6058,N_6436);
nand U7767 (N_7767,N_6128,N_6735);
nand U7768 (N_7768,N_7292,N_5094);
and U7769 (N_7769,N_5422,N_5961);
and U7770 (N_7770,N_6160,N_6614);
and U7771 (N_7771,N_5313,N_6694);
nand U7772 (N_7772,N_7269,N_7348);
nand U7773 (N_7773,N_5885,N_6329);
nor U7774 (N_7774,N_7140,N_6837);
nand U7775 (N_7775,N_7039,N_6167);
and U7776 (N_7776,N_5771,N_5836);
or U7777 (N_7777,N_6129,N_5069);
or U7778 (N_7778,N_6842,N_7256);
nand U7779 (N_7779,N_6269,N_6338);
nor U7780 (N_7780,N_7174,N_5983);
nand U7781 (N_7781,N_5521,N_5024);
and U7782 (N_7782,N_6661,N_5936);
and U7783 (N_7783,N_5949,N_5415);
or U7784 (N_7784,N_6241,N_7442);
or U7785 (N_7785,N_6424,N_7218);
nor U7786 (N_7786,N_5428,N_6991);
and U7787 (N_7787,N_7364,N_7109);
or U7788 (N_7788,N_6068,N_6115);
nand U7789 (N_7789,N_6714,N_5522);
and U7790 (N_7790,N_5439,N_5673);
nand U7791 (N_7791,N_6971,N_6082);
nor U7792 (N_7792,N_6243,N_5156);
nor U7793 (N_7793,N_6730,N_5541);
or U7794 (N_7794,N_6634,N_6703);
nor U7795 (N_7795,N_6500,N_5803);
or U7796 (N_7796,N_6156,N_7079);
nand U7797 (N_7797,N_6366,N_6469);
or U7798 (N_7798,N_6966,N_5745);
or U7799 (N_7799,N_7178,N_6886);
and U7800 (N_7800,N_5713,N_6319);
nand U7801 (N_7801,N_6667,N_6817);
nand U7802 (N_7802,N_6000,N_7398);
or U7803 (N_7803,N_6544,N_5483);
and U7804 (N_7804,N_5773,N_6202);
nand U7805 (N_7805,N_6056,N_6997);
nor U7806 (N_7806,N_5799,N_5547);
nor U7807 (N_7807,N_6902,N_6911);
and U7808 (N_7808,N_6549,N_7159);
or U7809 (N_7809,N_7195,N_7186);
and U7810 (N_7810,N_6165,N_6451);
nand U7811 (N_7811,N_6564,N_5545);
or U7812 (N_7812,N_5291,N_7430);
nor U7813 (N_7813,N_6415,N_6427);
nand U7814 (N_7814,N_5738,N_5243);
nand U7815 (N_7815,N_6135,N_6644);
nor U7816 (N_7816,N_5669,N_7022);
nand U7817 (N_7817,N_6213,N_6809);
and U7818 (N_7818,N_6558,N_6944);
nand U7819 (N_7819,N_7117,N_7250);
nor U7820 (N_7820,N_5828,N_6928);
nor U7821 (N_7821,N_6487,N_5468);
or U7822 (N_7822,N_7390,N_6762);
nand U7823 (N_7823,N_5249,N_5145);
or U7824 (N_7824,N_7115,N_7350);
nand U7825 (N_7825,N_5255,N_5021);
nand U7826 (N_7826,N_7143,N_5597);
or U7827 (N_7827,N_7193,N_6286);
or U7828 (N_7828,N_7227,N_6812);
nor U7829 (N_7829,N_6628,N_5630);
nand U7830 (N_7830,N_5199,N_5423);
nand U7831 (N_7831,N_7482,N_6750);
and U7832 (N_7832,N_6029,N_5346);
and U7833 (N_7833,N_6702,N_6759);
and U7834 (N_7834,N_6551,N_7070);
and U7835 (N_7835,N_6466,N_7339);
and U7836 (N_7836,N_6174,N_5507);
and U7837 (N_7837,N_7446,N_7304);
nand U7838 (N_7838,N_6591,N_5267);
nand U7839 (N_7839,N_6941,N_6356);
or U7840 (N_7840,N_7279,N_5381);
nand U7841 (N_7841,N_5154,N_6617);
nand U7842 (N_7842,N_7302,N_6616);
and U7843 (N_7843,N_5692,N_6035);
and U7844 (N_7844,N_7419,N_5095);
or U7845 (N_7845,N_6582,N_7179);
or U7846 (N_7846,N_6748,N_7392);
or U7847 (N_7847,N_7375,N_7307);
nor U7848 (N_7848,N_5446,N_6526);
or U7849 (N_7849,N_5747,N_7170);
nand U7850 (N_7850,N_6736,N_7361);
nor U7851 (N_7851,N_7328,N_6197);
or U7852 (N_7852,N_6746,N_6335);
and U7853 (N_7853,N_6839,N_6502);
nand U7854 (N_7854,N_5244,N_5640);
nand U7855 (N_7855,N_6327,N_5849);
nor U7856 (N_7856,N_7135,N_6084);
or U7857 (N_7857,N_5593,N_6801);
or U7858 (N_7858,N_5275,N_5621);
or U7859 (N_7859,N_6219,N_7353);
nand U7860 (N_7860,N_7054,N_6833);
or U7861 (N_7861,N_6822,N_7286);
or U7862 (N_7862,N_7335,N_6144);
nor U7863 (N_7863,N_6909,N_5996);
nand U7864 (N_7864,N_5627,N_5239);
or U7865 (N_7865,N_7454,N_5288);
nand U7866 (N_7866,N_6586,N_5682);
nand U7867 (N_7867,N_6566,N_6074);
nor U7868 (N_7868,N_5842,N_7118);
xor U7869 (N_7869,N_6774,N_5916);
or U7870 (N_7870,N_6537,N_5577);
nor U7871 (N_7871,N_6182,N_6931);
and U7872 (N_7872,N_5955,N_6993);
nand U7873 (N_7873,N_5491,N_6444);
and U7874 (N_7874,N_5658,N_6344);
nand U7875 (N_7875,N_6565,N_6053);
or U7876 (N_7876,N_7133,N_6662);
and U7877 (N_7877,N_7421,N_5344);
and U7878 (N_7878,N_6652,N_6732);
and U7879 (N_7879,N_5899,N_5071);
and U7880 (N_7880,N_6225,N_6118);
nand U7881 (N_7881,N_6711,N_5111);
or U7882 (N_7882,N_5398,N_6136);
nor U7883 (N_7883,N_7238,N_6898);
nand U7884 (N_7884,N_7497,N_5009);
nor U7885 (N_7885,N_6413,N_5394);
nor U7886 (N_7886,N_5589,N_5826);
nor U7887 (N_7887,N_5853,N_6701);
and U7888 (N_7888,N_5207,N_7449);
nand U7889 (N_7889,N_6889,N_5315);
or U7890 (N_7890,N_7088,N_6756);
nand U7891 (N_7891,N_7113,N_5134);
nor U7892 (N_7892,N_5012,N_7418);
and U7893 (N_7893,N_6535,N_5976);
and U7894 (N_7894,N_6547,N_5535);
or U7895 (N_7895,N_7300,N_5374);
nand U7896 (N_7896,N_5129,N_5930);
and U7897 (N_7897,N_5363,N_7080);
nor U7898 (N_7898,N_6813,N_6455);
and U7899 (N_7899,N_6245,N_6150);
and U7900 (N_7900,N_6555,N_7262);
nor U7901 (N_7901,N_7074,N_7401);
or U7902 (N_7902,N_5908,N_5753);
nor U7903 (N_7903,N_6904,N_7209);
or U7904 (N_7904,N_5832,N_6244);
nor U7905 (N_7905,N_5476,N_6673);
nand U7906 (N_7906,N_6460,N_6590);
nand U7907 (N_7907,N_7065,N_6423);
nor U7908 (N_7908,N_5829,N_5005);
nor U7909 (N_7909,N_5856,N_5191);
nor U7910 (N_7910,N_5761,N_6629);
and U7911 (N_7911,N_5789,N_7082);
and U7912 (N_7912,N_6664,N_6470);
xor U7913 (N_7913,N_6747,N_6249);
or U7914 (N_7914,N_6359,N_7312);
or U7915 (N_7915,N_6647,N_6844);
nand U7916 (N_7916,N_6072,N_5504);
and U7917 (N_7917,N_5311,N_7319);
nand U7918 (N_7918,N_5643,N_5447);
nand U7919 (N_7919,N_7123,N_7409);
nand U7920 (N_7920,N_6843,N_6408);
or U7921 (N_7921,N_6967,N_6438);
or U7922 (N_7922,N_6601,N_7141);
and U7923 (N_7923,N_5868,N_6334);
nor U7924 (N_7924,N_5127,N_5732);
or U7925 (N_7925,N_6336,N_6632);
nand U7926 (N_7926,N_6952,N_6005);
nor U7927 (N_7927,N_5567,N_5117);
and U7928 (N_7928,N_6924,N_5958);
nor U7929 (N_7929,N_7103,N_6540);
nand U7930 (N_7930,N_6786,N_5116);
or U7931 (N_7931,N_5726,N_5448);
nor U7932 (N_7932,N_6262,N_5097);
nand U7933 (N_7933,N_6955,N_6598);
or U7934 (N_7934,N_7411,N_7349);
nor U7935 (N_7935,N_5798,N_5214);
or U7936 (N_7936,N_6719,N_6990);
nor U7937 (N_7937,N_7067,N_6867);
and U7938 (N_7938,N_6850,N_6294);
and U7939 (N_7939,N_7486,N_6501);
or U7940 (N_7940,N_7139,N_5659);
or U7941 (N_7941,N_5161,N_6032);
and U7942 (N_7942,N_7255,N_5792);
and U7943 (N_7943,N_7124,N_6761);
or U7944 (N_7944,N_5090,N_5011);
or U7945 (N_7945,N_5179,N_6973);
nand U7946 (N_7946,N_6119,N_6297);
nand U7947 (N_7947,N_5361,N_6059);
nand U7948 (N_7948,N_5733,N_5411);
and U7949 (N_7949,N_5731,N_5905);
or U7950 (N_7950,N_6561,N_6302);
nor U7951 (N_7951,N_7038,N_5484);
or U7952 (N_7952,N_6491,N_6668);
or U7953 (N_7953,N_6461,N_6933);
nor U7954 (N_7954,N_5815,N_6168);
nand U7955 (N_7955,N_6770,N_5325);
nor U7956 (N_7956,N_5755,N_5354);
and U7957 (N_7957,N_7308,N_5827);
or U7958 (N_7958,N_7018,N_6342);
nand U7959 (N_7959,N_6457,N_5876);
nand U7960 (N_7960,N_7147,N_7199);
nand U7961 (N_7961,N_6685,N_6620);
nand U7962 (N_7962,N_6821,N_7063);
nor U7963 (N_7963,N_5754,N_5903);
or U7964 (N_7964,N_6584,N_6309);
nand U7965 (N_7965,N_5473,N_5277);
and U7966 (N_7966,N_5946,N_6148);
nor U7967 (N_7967,N_5086,N_5321);
or U7968 (N_7968,N_5173,N_6001);
or U7969 (N_7969,N_6376,N_6557);
and U7970 (N_7970,N_5489,N_5811);
and U7971 (N_7971,N_7121,N_6726);
nor U7972 (N_7972,N_6704,N_6863);
nor U7973 (N_7973,N_6166,N_5750);
and U7974 (N_7974,N_5816,N_5390);
nor U7975 (N_7975,N_5000,N_7478);
and U7976 (N_7976,N_5248,N_7053);
or U7977 (N_7977,N_7211,N_5959);
nand U7978 (N_7978,N_6996,N_5512);
nor U7979 (N_7979,N_7183,N_5500);
or U7980 (N_7980,N_6879,N_5742);
nand U7981 (N_7981,N_5332,N_5704);
and U7982 (N_7982,N_5337,N_6827);
nand U7983 (N_7983,N_6988,N_5382);
and U7984 (N_7984,N_5901,N_5620);
and U7985 (N_7985,N_7066,N_6481);
and U7986 (N_7986,N_5629,N_6874);
nand U7987 (N_7987,N_7331,N_5287);
and U7988 (N_7988,N_5132,N_6237);
or U7989 (N_7989,N_5917,N_5201);
nor U7990 (N_7990,N_6773,N_5149);
and U7991 (N_7991,N_5036,N_6467);
nand U7992 (N_7992,N_5553,N_5558);
and U7993 (N_7993,N_7259,N_5889);
nor U7994 (N_7994,N_5531,N_5513);
or U7995 (N_7995,N_5418,N_6442);
nand U7996 (N_7996,N_5273,N_5532);
nor U7997 (N_7997,N_7188,N_7068);
or U7998 (N_7998,N_5060,N_7156);
nand U7999 (N_7999,N_6818,N_5320);
or U8000 (N_8000,N_7475,N_5982);
or U8001 (N_8001,N_6154,N_7233);
or U8002 (N_8002,N_5061,N_6987);
nor U8003 (N_8003,N_6706,N_5740);
and U8004 (N_8004,N_5580,N_5702);
or U8005 (N_8005,N_5671,N_6912);
and U8006 (N_8006,N_6989,N_6127);
and U8007 (N_8007,N_5352,N_5140);
xor U8008 (N_8008,N_7100,N_7034);
nand U8009 (N_8009,N_6927,N_6192);
and U8010 (N_8010,N_5927,N_5029);
or U8011 (N_8011,N_5187,N_7011);
nor U8012 (N_8012,N_5648,N_5534);
or U8013 (N_8013,N_6153,N_6386);
and U8014 (N_8014,N_7072,N_7281);
xnor U8015 (N_8015,N_5488,N_7404);
or U8016 (N_8016,N_5206,N_6098);
and U8017 (N_8017,N_7346,N_6828);
nand U8018 (N_8018,N_5764,N_6475);
nand U8019 (N_8019,N_7020,N_6883);
nand U8020 (N_8020,N_7050,N_7275);
or U8021 (N_8021,N_7280,N_7228);
nor U8022 (N_8022,N_5237,N_5143);
and U8023 (N_8023,N_5752,N_5404);
nand U8024 (N_8024,N_5647,N_6728);
nor U8025 (N_8025,N_7243,N_5636);
or U8026 (N_8026,N_5527,N_6314);
nor U8027 (N_8027,N_5718,N_5804);
and U8028 (N_8028,N_5092,N_6998);
nand U8029 (N_8029,N_5269,N_5139);
nand U8030 (N_8030,N_6208,N_6597);
nor U8031 (N_8031,N_6435,N_7499);
or U8032 (N_8032,N_5963,N_5106);
or U8033 (N_8033,N_6345,N_7158);
nor U8034 (N_8034,N_6251,N_7003);
and U8035 (N_8035,N_6892,N_7340);
or U8036 (N_8036,N_6943,N_5679);
and U8037 (N_8037,N_7208,N_5865);
nor U8038 (N_8038,N_5073,N_6246);
nor U8039 (N_8039,N_7376,N_7287);
nor U8040 (N_8040,N_6411,N_7232);
nor U8041 (N_8041,N_6145,N_5229);
and U8042 (N_8042,N_7059,N_7297);
nand U8043 (N_8043,N_6374,N_6315);
nand U8044 (N_8044,N_6958,N_7373);
nor U8045 (N_8045,N_6485,N_5100);
nand U8046 (N_8046,N_6028,N_7138);
or U8047 (N_8047,N_6509,N_6640);
or U8048 (N_8048,N_5586,N_5034);
or U8049 (N_8049,N_5054,N_6956);
or U8050 (N_8050,N_5751,N_5458);
nand U8051 (N_8051,N_6038,N_5271);
nor U8052 (N_8052,N_5425,N_5835);
and U8053 (N_8053,N_6757,N_6459);
nand U8054 (N_8054,N_5314,N_5881);
nand U8055 (N_8055,N_7386,N_6578);
and U8056 (N_8056,N_6462,N_5474);
or U8057 (N_8057,N_6624,N_6061);
nand U8058 (N_8058,N_7394,N_5309);
nor U8059 (N_8059,N_5797,N_6918);
nand U8060 (N_8060,N_5502,N_5470);
nor U8061 (N_8061,N_5205,N_7192);
nand U8062 (N_8062,N_5331,N_5096);
nand U8063 (N_8063,N_6936,N_7009);
nor U8064 (N_8064,N_6282,N_5290);
or U8065 (N_8065,N_7354,N_5482);
and U8066 (N_8066,N_6925,N_5171);
nor U8067 (N_8067,N_7222,N_5167);
nor U8068 (N_8068,N_5837,N_6965);
or U8069 (N_8069,N_6425,N_6897);
nor U8070 (N_8070,N_7105,N_5506);
nand U8071 (N_8071,N_7127,N_7370);
nor U8072 (N_8072,N_6362,N_5032);
nor U8073 (N_8073,N_6923,N_6447);
or U8074 (N_8074,N_6125,N_6221);
or U8075 (N_8075,N_5790,N_6806);
or U8076 (N_8076,N_6218,N_6781);
nor U8077 (N_8077,N_6299,N_5040);
nor U8078 (N_8078,N_6189,N_6798);
nor U8079 (N_8079,N_5391,N_5437);
nand U8080 (N_8080,N_7324,N_6017);
or U8081 (N_8081,N_6057,N_6569);
nand U8082 (N_8082,N_7322,N_6393);
nor U8083 (N_8083,N_5192,N_5935);
and U8084 (N_8084,N_6343,N_5426);
nor U8085 (N_8085,N_6529,N_7241);
or U8086 (N_8086,N_5912,N_5421);
nor U8087 (N_8087,N_5257,N_6382);
nor U8088 (N_8088,N_6397,N_7283);
nand U8089 (N_8089,N_6796,N_5555);
and U8090 (N_8090,N_6630,N_7476);
nand U8091 (N_8091,N_6838,N_6014);
or U8092 (N_8092,N_7104,N_5757);
nand U8093 (N_8093,N_6023,N_5339);
or U8094 (N_8094,N_6261,N_6804);
nor U8095 (N_8095,N_5578,N_7069);
and U8096 (N_8096,N_5072,N_7166);
or U8097 (N_8097,N_6013,N_6740);
nor U8098 (N_8098,N_5310,N_6080);
or U8099 (N_8099,N_5150,N_5264);
or U8100 (N_8100,N_6649,N_7176);
nor U8101 (N_8101,N_6723,N_6108);
nand U8102 (N_8102,N_7111,N_6553);
nor U8103 (N_8103,N_5025,N_5087);
or U8104 (N_8104,N_5254,N_6875);
or U8105 (N_8105,N_7374,N_6797);
and U8106 (N_8106,N_5759,N_7064);
nor U8107 (N_8107,N_5057,N_5743);
nand U8108 (N_8108,N_6083,N_6328);
or U8109 (N_8109,N_5076,N_6039);
and U8110 (N_8110,N_5463,N_6511);
nand U8111 (N_8111,N_6304,N_5449);
and U8112 (N_8112,N_6446,N_6716);
or U8113 (N_8113,N_6322,N_6999);
nor U8114 (N_8114,N_7291,N_6697);
or U8115 (N_8115,N_5281,N_7060);
nand U8116 (N_8116,N_7028,N_5933);
nor U8117 (N_8117,N_6133,N_6069);
and U8118 (N_8118,N_5487,N_6280);
or U8119 (N_8119,N_6050,N_6468);
or U8120 (N_8120,N_6385,N_7402);
and U8121 (N_8121,N_7023,N_5951);
nor U8122 (N_8122,N_6771,N_6793);
nor U8123 (N_8123,N_5778,N_6492);
nand U8124 (N_8124,N_5964,N_7443);
and U8125 (N_8125,N_5539,N_5135);
nand U8126 (N_8126,N_6030,N_6420);
and U8127 (N_8127,N_5519,N_5295);
nand U8128 (N_8128,N_6178,N_5774);
or U8129 (N_8129,N_6379,N_6258);
and U8130 (N_8130,N_6708,N_7242);
nor U8131 (N_8131,N_5802,N_6810);
nor U8132 (N_8132,N_5653,N_6554);
or U8133 (N_8133,N_7301,N_5345);
and U8134 (N_8134,N_6206,N_6496);
xnor U8135 (N_8135,N_7276,N_6720);
or U8136 (N_8136,N_6789,N_7008);
nand U8137 (N_8137,N_5107,N_5614);
nand U8138 (N_8138,N_6199,N_5362);
or U8139 (N_8139,N_6151,N_7397);
or U8140 (N_8140,N_7000,N_6659);
nand U8141 (N_8141,N_7168,N_6493);
nor U8142 (N_8142,N_5980,N_6276);
nand U8143 (N_8143,N_6274,N_5944);
and U8144 (N_8144,N_5542,N_5312);
nand U8145 (N_8145,N_6312,N_7032);
or U8146 (N_8146,N_7338,N_5368);
or U8147 (N_8147,N_5232,N_6090);
or U8148 (N_8148,N_7405,N_5213);
and U8149 (N_8149,N_6497,N_6725);
nor U8150 (N_8150,N_5635,N_5017);
nand U8151 (N_8151,N_7040,N_6618);
or U8152 (N_8152,N_6949,N_5296);
nor U8153 (N_8153,N_6087,N_6751);
or U8154 (N_8154,N_6835,N_6378);
or U8155 (N_8155,N_5416,N_5939);
or U8156 (N_8156,N_5645,N_6076);
and U8157 (N_8157,N_5388,N_6534);
nand U8158 (N_8158,N_6665,N_5496);
nor U8159 (N_8159,N_6147,N_7290);
nand U8160 (N_8160,N_5524,N_5342);
and U8161 (N_8161,N_5971,N_5896);
and U8162 (N_8162,N_5991,N_6306);
and U8163 (N_8163,N_5431,N_6688);
or U8164 (N_8164,N_5678,N_6682);
or U8165 (N_8165,N_5083,N_5999);
or U8166 (N_8166,N_5308,N_5579);
nand U8167 (N_8167,N_6367,N_6722);
and U8168 (N_8168,N_6383,N_7380);
and U8169 (N_8169,N_6216,N_7030);
nand U8170 (N_8170,N_5765,N_5226);
or U8171 (N_8171,N_6712,N_6541);
or U8172 (N_8172,N_5402,N_6004);
nor U8173 (N_8173,N_6605,N_5104);
nand U8174 (N_8174,N_6036,N_6775);
or U8175 (N_8175,N_5681,N_7252);
and U8176 (N_8176,N_5965,N_6279);
or U8177 (N_8177,N_7477,N_5022);
nor U8178 (N_8178,N_7479,N_7010);
and U8179 (N_8179,N_6250,N_6894);
or U8180 (N_8180,N_5795,N_5146);
nor U8181 (N_8181,N_5608,N_7379);
or U8182 (N_8182,N_5576,N_5786);
nor U8183 (N_8183,N_6595,N_5907);
or U8184 (N_8184,N_5538,N_5316);
or U8185 (N_8185,N_5302,N_5004);
nand U8186 (N_8186,N_6240,N_5157);
or U8187 (N_8187,N_6895,N_6942);
nor U8188 (N_8188,N_6042,N_5245);
nand U8189 (N_8189,N_6621,N_5469);
nand U8190 (N_8190,N_6333,N_6610);
or U8191 (N_8191,N_6163,N_6820);
nor U8192 (N_8192,N_6579,N_7146);
or U8193 (N_8193,N_7150,N_5093);
or U8194 (N_8194,N_5085,N_6583);
nor U8195 (N_8195,N_5748,N_5102);
and U8196 (N_8196,N_6045,N_6891);
and U8197 (N_8197,N_7237,N_6805);
and U8198 (N_8198,N_5656,N_5575);
or U8199 (N_8199,N_5686,N_7025);
and U8200 (N_8200,N_6611,N_5737);
nand U8201 (N_8201,N_7481,N_5347);
nand U8202 (N_8202,N_7389,N_7264);
or U8203 (N_8203,N_5844,N_7494);
or U8204 (N_8204,N_5338,N_5010);
and U8205 (N_8205,N_7142,N_6739);
nor U8206 (N_8206,N_5285,N_5420);
and U8207 (N_8207,N_5051,N_5279);
nor U8208 (N_8208,N_5367,N_6337);
and U8209 (N_8209,N_5014,N_6681);
nor U8210 (N_8210,N_5995,N_5395);
and U8211 (N_8211,N_5626,N_6903);
and U8212 (N_8212,N_5741,N_7017);
or U8213 (N_8213,N_5714,N_6570);
nor U8214 (N_8214,N_6506,N_6763);
nor U8215 (N_8215,N_5793,N_7347);
nor U8216 (N_8216,N_7029,N_7094);
nor U8217 (N_8217,N_6232,N_6683);
nand U8218 (N_8218,N_7224,N_6678);
nor U8219 (N_8219,N_7220,N_7055);
nor U8220 (N_8220,N_5631,N_5383);
nand U8221 (N_8221,N_5979,N_6473);
nor U8222 (N_8222,N_6823,N_5919);
and U8223 (N_8223,N_5918,N_6938);
and U8224 (N_8224,N_6619,N_6950);
xnor U8225 (N_8225,N_5088,N_7456);
nor U8226 (N_8226,N_7249,N_5924);
nand U8227 (N_8227,N_5015,N_5854);
nand U8228 (N_8228,N_6207,N_7087);
nand U8229 (N_8229,N_5372,N_5861);
or U8230 (N_8230,N_7203,N_7210);
nor U8231 (N_8231,N_6733,N_5840);
and U8232 (N_8232,N_5968,N_5341);
and U8233 (N_8233,N_6364,N_7447);
nand U8234 (N_8234,N_7298,N_5317);
nor U8235 (N_8235,N_5562,N_5898);
xnor U8236 (N_8236,N_6472,N_6679);
or U8237 (N_8237,N_6932,N_5365);
or U8238 (N_8238,N_5133,N_6482);
or U8239 (N_8239,N_5251,N_5894);
and U8240 (N_8240,N_5915,N_6021);
and U8241 (N_8241,N_7165,N_6680);
nand U8242 (N_8242,N_6351,N_5045);
or U8243 (N_8243,N_6081,N_6846);
nand U8244 (N_8244,N_5193,N_6441);
nand U8245 (N_8245,N_7305,N_6857);
nand U8246 (N_8246,N_6392,N_6159);
and U8247 (N_8247,N_6211,N_5451);
nor U8248 (N_8248,N_5185,N_5230);
nor U8249 (N_8249,N_6235,N_7438);
nand U8250 (N_8250,N_6051,N_6471);
nor U8251 (N_8251,N_5574,N_7167);
nand U8252 (N_8252,N_6645,N_5684);
nor U8253 (N_8253,N_5165,N_6456);
and U8254 (N_8254,N_5356,N_5294);
and U8255 (N_8255,N_5227,N_7460);
and U8256 (N_8256,N_5926,N_6137);
nand U8257 (N_8257,N_5734,N_5780);
nor U8258 (N_8258,N_6868,N_7363);
nand U8259 (N_8259,N_7089,N_7075);
or U8260 (N_8260,N_6588,N_6937);
xor U8261 (N_8261,N_5651,N_5668);
nor U8262 (N_8262,N_7164,N_7388);
nand U8263 (N_8263,N_5223,N_5475);
or U8264 (N_8264,N_5989,N_7435);
or U8265 (N_8265,N_5667,N_6490);
nand U8266 (N_8266,N_5335,N_5801);
nor U8267 (N_8267,N_6239,N_7048);
and U8268 (N_8268,N_5182,N_7019);
and U8269 (N_8269,N_5932,N_5911);
and U8270 (N_8270,N_5674,N_6738);
and U8271 (N_8271,N_6929,N_6737);
or U8272 (N_8272,N_5110,N_5594);
nor U8273 (N_8273,N_6960,N_6849);
nor U8274 (N_8274,N_6266,N_5503);
or U8275 (N_8275,N_7126,N_6320);
or U8276 (N_8276,N_5813,N_6479);
and U8277 (N_8277,N_7288,N_5900);
and U8278 (N_8278,N_7101,N_6201);
nor U8279 (N_8279,N_6870,N_5848);
nand U8280 (N_8280,N_5497,N_5130);
nor U8281 (N_8281,N_6331,N_6517);
nand U8282 (N_8282,N_5711,N_5490);
nor U8283 (N_8283,N_6651,N_5152);
nand U8284 (N_8284,N_5455,N_6305);
or U8285 (N_8285,N_7355,N_6433);
nor U8286 (N_8286,N_5566,N_5174);
nand U8287 (N_8287,N_5169,N_6330);
nor U8288 (N_8288,N_5529,N_7299);
and U8289 (N_8289,N_6253,N_6731);
nand U8290 (N_8290,N_7021,N_6077);
nand U8291 (N_8291,N_7272,N_5528);
or U8292 (N_8292,N_7057,N_6946);
nand U8293 (N_8293,N_7395,N_6405);
nand U8294 (N_8294,N_7225,N_7235);
nand U8295 (N_8295,N_6858,N_5075);
nand U8296 (N_8296,N_5058,N_6010);
nor U8297 (N_8297,N_5300,N_5978);
nand U8298 (N_8298,N_6428,N_6845);
nand U8299 (N_8299,N_5081,N_6660);
or U8300 (N_8300,N_5831,N_6454);
and U8301 (N_8301,N_5984,N_6948);
or U8302 (N_8302,N_7120,N_5685);
or U8303 (N_8303,N_6968,N_5272);
nand U8304 (N_8304,N_5082,N_5783);
nor U8305 (N_8305,N_6191,N_5897);
or U8306 (N_8306,N_6388,N_7096);
and U8307 (N_8307,N_5136,N_6102);
or U8308 (N_8308,N_7129,N_6574);
nor U8309 (N_8309,N_6576,N_5557);
or U8310 (N_8310,N_7196,N_7108);
or U8311 (N_8311,N_5063,N_7071);
or U8312 (N_8312,N_6860,N_5806);
nand U8313 (N_8313,N_5033,N_5690);
nand U8314 (N_8314,N_6141,N_7043);
or U8315 (N_8315,N_5950,N_6012);
or U8316 (N_8316,N_5370,N_7366);
and U8317 (N_8317,N_7270,N_6079);
nand U8318 (N_8318,N_6419,N_5800);
and U8319 (N_8319,N_5559,N_5253);
nor U8320 (N_8320,N_5633,N_6788);
nand U8321 (N_8321,N_7027,N_5833);
nor U8322 (N_8322,N_6418,N_6744);
or U8323 (N_8323,N_5466,N_6864);
nor U8324 (N_8324,N_6349,N_6819);
nand U8325 (N_8325,N_5144,N_5707);
or U8326 (N_8326,N_6921,N_6448);
or U8327 (N_8327,N_6825,N_7393);
and U8328 (N_8328,N_6489,N_7453);
and U8329 (N_8329,N_6360,N_5644);
nand U8330 (N_8330,N_5121,N_5720);
nand U8331 (N_8331,N_5805,N_5517);
and U8332 (N_8332,N_7295,N_5670);
or U8333 (N_8333,N_5920,N_7434);
or U8334 (N_8334,N_5235,N_6131);
nor U8335 (N_8335,N_6979,N_5666);
nand U8336 (N_8336,N_7145,N_6478);
nor U8337 (N_8337,N_6453,N_5739);
nand U8338 (N_8338,N_5289,N_5986);
and U8339 (N_8339,N_5689,N_7492);
nand U8340 (N_8340,N_7016,N_6543);
and U8341 (N_8341,N_7267,N_5814);
nand U8342 (N_8342,N_7360,N_7231);
or U8343 (N_8343,N_7429,N_6272);
nor U8344 (N_8344,N_7173,N_6116);
and U8345 (N_8345,N_6318,N_5728);
and U8346 (N_8346,N_5070,N_6139);
and U8347 (N_8347,N_5434,N_5947);
or U8348 (N_8348,N_7134,N_7031);
nand U8349 (N_8349,N_5238,N_6037);
and U8350 (N_8350,N_5397,N_5634);
or U8351 (N_8351,N_7472,N_6675);
or U8352 (N_8352,N_5649,N_5874);
nor U8353 (N_8353,N_6871,N_7153);
and U8354 (N_8354,N_5438,N_5537);
nor U8355 (N_8355,N_5665,N_5592);
or U8356 (N_8356,N_7136,N_6636);
nand U8357 (N_8357,N_6103,N_6715);
or U8358 (N_8358,N_7107,N_7001);
and U8359 (N_8359,N_5776,N_6550);
or U8360 (N_8360,N_7484,N_6978);
and U8361 (N_8361,N_7046,N_6105);
and U8362 (N_8362,N_6992,N_6426);
and U8363 (N_8363,N_7083,N_5921);
nor U8364 (N_8364,N_5377,N_6777);
nand U8365 (N_8365,N_6580,N_5960);
xnor U8366 (N_8366,N_5186,N_6572);
xor U8367 (N_8367,N_5462,N_6522);
nand U8368 (N_8368,N_6070,N_7013);
and U8369 (N_8369,N_6816,N_6852);
nor U8370 (N_8370,N_5467,N_5023);
and U8371 (N_8371,N_6710,N_5530);
nand U8372 (N_8372,N_7357,N_5914);
nor U8373 (N_8373,N_5074,N_5572);
or U8374 (N_8374,N_5956,N_5824);
and U8375 (N_8375,N_6210,N_5725);
nand U8376 (N_8376,N_7163,N_6513);
or U8377 (N_8377,N_5410,N_5808);
and U8378 (N_8378,N_5172,N_5823);
nor U8379 (N_8379,N_6794,N_6676);
or U8380 (N_8380,N_7391,N_5479);
nor U8381 (N_8381,N_5887,N_6575);
nand U8382 (N_8382,N_6947,N_7216);
nand U8383 (N_8383,N_7090,N_5211);
nor U8384 (N_8384,N_7122,N_6008);
nand U8385 (N_8385,N_5943,N_7403);
and U8386 (N_8386,N_6768,N_6365);
nand U8387 (N_8387,N_6608,N_7326);
and U8388 (N_8388,N_6186,N_6060);
nor U8389 (N_8389,N_5994,N_5722);
and U8390 (N_8390,N_5353,N_5584);
and U8391 (N_8391,N_7420,N_5859);
nor U8392 (N_8392,N_6604,N_7181);
nor U8393 (N_8393,N_6499,N_6721);
and U8394 (N_8394,N_7495,N_6340);
nor U8395 (N_8395,N_5357,N_5042);
or U8396 (N_8396,N_5228,N_5494);
nand U8397 (N_8397,N_6692,N_6533);
nor U8398 (N_8398,N_6179,N_6890);
and U8399 (N_8399,N_6185,N_6228);
or U8400 (N_8400,N_7128,N_7125);
nand U8401 (N_8401,N_6981,N_6693);
nand U8402 (N_8402,N_5564,N_5142);
nor U8403 (N_8403,N_5413,N_5373);
nand U8404 (N_8404,N_6935,N_7345);
nor U8405 (N_8405,N_6523,N_6521);
and U8406 (N_8406,N_5974,N_5967);
nor U8407 (N_8407,N_5664,N_7330);
nor U8408 (N_8408,N_5972,N_6684);
nand U8409 (N_8409,N_5925,N_7187);
nor U8410 (N_8410,N_7334,N_5098);
and U8411 (N_8411,N_5052,N_6494);
or U8412 (N_8412,N_6635,N_5303);
or U8413 (N_8413,N_6255,N_5044);
or U8414 (N_8414,N_7396,N_5498);
nor U8415 (N_8415,N_6194,N_5791);
nor U8416 (N_8416,N_5188,N_6132);
nor U8417 (N_8417,N_5735,N_7215);
nor U8418 (N_8418,N_5137,N_6432);
nor U8419 (N_8419,N_6690,N_6980);
nand U8420 (N_8420,N_5866,N_7441);
nor U8421 (N_8421,N_6800,N_6603);
and U8422 (N_8422,N_5509,N_5938);
nor U8423 (N_8423,N_5234,N_7465);
nor U8424 (N_8424,N_6626,N_5785);
nor U8425 (N_8425,N_5948,N_7185);
and U8426 (N_8426,N_5606,N_7198);
or U8427 (N_8427,N_7077,N_5518);
or U8428 (N_8428,N_7239,N_6190);
nor U8429 (N_8429,N_5203,N_6982);
and U8430 (N_8430,N_5250,N_5055);
nand U8431 (N_8431,N_5225,N_7049);
or U8432 (N_8432,N_7488,N_7313);
and U8433 (N_8433,N_6767,N_6772);
or U8434 (N_8434,N_5471,N_5700);
or U8435 (N_8435,N_5706,N_7175);
and U8436 (N_8436,N_5879,N_6677);
or U8437 (N_8437,N_6814,N_5196);
nand U8438 (N_8438,N_5003,N_6348);
or U8439 (N_8439,N_5480,N_6503);
nor U8440 (N_8440,N_6963,N_6301);
nand U8441 (N_8441,N_5623,N_7480);
nor U8442 (N_8442,N_5788,N_6164);
and U8443 (N_8443,N_5080,N_5266);
xor U8444 (N_8444,N_7160,N_6972);
or U8445 (N_8445,N_6495,N_6400);
nor U8446 (N_8446,N_7114,N_5450);
nand U8447 (N_8447,N_5202,N_5526);
and U8448 (N_8448,N_5292,N_6371);
and U8449 (N_8449,N_6589,N_6016);
nand U8450 (N_8450,N_7266,N_7191);
nand U8451 (N_8451,N_7470,N_5977);
nand U8452 (N_8452,N_6865,N_5189);
or U8453 (N_8453,N_5047,N_5657);
nand U8454 (N_8454,N_5018,N_6187);
and U8455 (N_8455,N_7036,N_5845);
and U8456 (N_8456,N_6581,N_7493);
nand U8457 (N_8457,N_6824,N_6934);
nand U8458 (N_8458,N_6264,N_7162);
nand U8459 (N_8459,N_5184,N_5066);
xnor U8460 (N_8460,N_7485,N_5940);
or U8461 (N_8461,N_7095,N_5922);
and U8462 (N_8462,N_5619,N_5906);
nand U8463 (N_8463,N_6152,N_5419);
and U8464 (N_8464,N_5283,N_6542);
and U8465 (N_8465,N_5770,N_7440);
or U8466 (N_8466,N_6906,N_6847);
nor U8467 (N_8467,N_6063,N_7332);
or U8468 (N_8468,N_6044,N_7285);
or U8469 (N_8469,N_6592,N_5895);
or U8470 (N_8470,N_7002,N_5459);
and U8471 (N_8471,N_7425,N_6247);
xor U8472 (N_8472,N_6404,N_5822);
and U8473 (N_8473,N_6200,N_5928);
nand U8474 (N_8474,N_6882,N_6217);
nor U8475 (N_8475,N_7467,N_6532);
or U8476 (N_8476,N_5724,N_6138);
or U8477 (N_8477,N_6959,N_7278);
and U8478 (N_8478,N_7161,N_6705);
nor U8479 (N_8479,N_6623,N_5120);
nand U8480 (N_8480,N_5242,N_6172);
nor U8481 (N_8481,N_7261,N_6905);
and U8482 (N_8482,N_7091,N_5348);
or U8483 (N_8483,N_7206,N_5222);
xnor U8484 (N_8484,N_5769,N_5399);
or U8485 (N_8485,N_7282,N_6398);
nor U8486 (N_8486,N_5477,N_6226);
or U8487 (N_8487,N_5717,N_6412);
nor U8488 (N_8488,N_7204,N_6880);
and U8489 (N_8489,N_5427,N_7230);
and U8490 (N_8490,N_6003,N_6238);
nor U8491 (N_8491,N_7303,N_5386);
nand U8492 (N_8492,N_5601,N_6964);
or U8493 (N_8493,N_5430,N_6696);
or U8494 (N_8494,N_5355,N_6146);
nor U8495 (N_8495,N_7024,N_5486);
nor U8496 (N_8496,N_6121,N_5351);
or U8497 (N_8497,N_5119,N_5282);
nor U8498 (N_8498,N_6655,N_7399);
nor U8499 (N_8499,N_5153,N_6403);
nand U8500 (N_8500,N_6803,N_5923);
and U8501 (N_8501,N_5260,N_6625);
nor U8502 (N_8502,N_7377,N_7473);
and U8503 (N_8503,N_7428,N_6065);
and U8504 (N_8504,N_6709,N_7012);
nand U8505 (N_8505,N_5843,N_5603);
nor U8506 (N_8506,N_5387,N_5687);
nand U8507 (N_8507,N_6607,N_5301);
nor U8508 (N_8508,N_7144,N_6396);
nor U8509 (N_8509,N_7116,N_5371);
and U8510 (N_8510,N_5625,N_7202);
nand U8511 (N_8511,N_5975,N_6040);
nand U8512 (N_8512,N_6486,N_5442);
nor U8513 (N_8513,N_6439,N_6606);
and U8514 (N_8514,N_5041,N_6866);
or U8515 (N_8515,N_6033,N_6452);
nand U8516 (N_8516,N_5181,N_6402);
and U8517 (N_8517,N_6347,N_5220);
or U8518 (N_8518,N_7424,N_6267);
nor U8519 (N_8519,N_7260,N_5767);
nor U8520 (N_8520,N_7051,N_5588);
and U8521 (N_8521,N_6596,N_7076);
and U8522 (N_8522,N_6464,N_7130);
nand U8523 (N_8523,N_5953,N_6764);
nor U8524 (N_8524,N_6556,N_5573);
nor U8525 (N_8525,N_6826,N_5851);
nand U8526 (N_8526,N_7352,N_7471);
nor U8527 (N_8527,N_5333,N_5329);
nor U8528 (N_8528,N_6018,N_7277);
nand U8529 (N_8529,N_7474,N_6027);
and U8530 (N_8530,N_7466,N_6530);
nor U8531 (N_8531,N_6639,N_5600);
or U8532 (N_8532,N_5053,N_6920);
xnor U8533 (N_8533,N_6977,N_7414);
or U8534 (N_8534,N_5065,N_6791);
nand U8535 (N_8535,N_5038,N_5869);
and U8536 (N_8536,N_6254,N_5217);
xnor U8537 (N_8537,N_5890,N_6110);
nor U8538 (N_8538,N_6734,N_6986);
nand U8539 (N_8539,N_6851,N_5762);
or U8540 (N_8540,N_5400,N_7344);
nor U8541 (N_8541,N_5158,N_5204);
nor U8542 (N_8542,N_5241,N_6707);
or U8543 (N_8543,N_5934,N_7455);
nor U8544 (N_8544,N_5141,N_6046);
nand U8545 (N_8545,N_7415,N_7483);
and U8546 (N_8546,N_6834,N_6009);
and U8547 (N_8547,N_6181,N_5615);
and U8548 (N_8548,N_6157,N_6559);
nand U8549 (N_8549,N_7423,N_5122);
and U8550 (N_8550,N_5543,N_5694);
or U8551 (N_8551,N_6562,N_7149);
and U8552 (N_8552,N_6284,N_7131);
nor U8553 (N_8553,N_6612,N_6749);
or U8554 (N_8554,N_6203,N_7271);
or U8555 (N_8555,N_6512,N_5270);
or U8556 (N_8556,N_7007,N_6048);
nor U8557 (N_8557,N_6853,N_5652);
and U8558 (N_8558,N_7106,N_5208);
or U8559 (N_8559,N_6067,N_6563);
nor U8560 (N_8560,N_5569,N_6782);
nor U8561 (N_8561,N_6389,N_7219);
nor U8562 (N_8562,N_7132,N_5319);
nand U8563 (N_8563,N_5350,N_5236);
nor U8564 (N_8564,N_5396,N_7223);
or U8565 (N_8565,N_6109,N_7337);
nand U8566 (N_8566,N_5508,N_7247);
nor U8567 (N_8567,N_5414,N_7498);
or U8568 (N_8568,N_5218,N_6230);
or U8569 (N_8569,N_5782,N_6242);
nand U8570 (N_8570,N_6717,N_6410);
and U8571 (N_8571,N_7368,N_5749);
nor U8572 (N_8572,N_7169,N_5703);
or U8573 (N_8573,N_6627,N_6815);
and U8574 (N_8574,N_5304,N_6674);
or U8575 (N_8575,N_7381,N_6434);
or U8576 (N_8576,N_5412,N_5990);
or U8577 (N_8577,N_5392,N_6198);
and U8578 (N_8578,N_5942,N_6901);
nor U8579 (N_8579,N_6899,N_5170);
or U8580 (N_8580,N_5148,N_5693);
nor U8581 (N_8581,N_6792,N_7045);
or U8582 (N_8582,N_5160,N_5176);
or U8583 (N_8583,N_7458,N_5591);
nand U8584 (N_8584,N_6463,N_5166);
nand U8585 (N_8585,N_6031,N_5650);
and U8586 (N_8586,N_7408,N_5126);
and U8587 (N_8587,N_5540,N_7284);
nand U8588 (N_8588,N_5436,N_5699);
nand U8589 (N_8589,N_6215,N_6352);
nand U8590 (N_8590,N_6278,N_5369);
nor U8591 (N_8591,N_5834,N_6086);
nor U8592 (N_8592,N_5909,N_6896);
and U8593 (N_8593,N_5209,N_6633);
nand U8594 (N_8594,N_5155,N_5756);
nor U8595 (N_8595,N_6177,N_7014);
and U8596 (N_8596,N_5663,N_5867);
and U8597 (N_8597,N_6380,N_5258);
and U8598 (N_8598,N_5552,N_7433);
or U8599 (N_8599,N_6195,N_5006);
nand U8600 (N_8600,N_6663,N_6401);
and U8601 (N_8601,N_6332,N_7263);
nand U8602 (N_8602,N_5812,N_5794);
nand U8603 (N_8603,N_5893,N_7221);
and U8604 (N_8604,N_5655,N_6593);
or U8605 (N_8605,N_6974,N_7177);
and U8606 (N_8606,N_6995,N_5945);
nand U8607 (N_8607,N_6525,N_6666);
and U8608 (N_8608,N_5618,N_6310);
or U8609 (N_8609,N_7437,N_6515);
nor U8610 (N_8610,N_7200,N_6020);
and U8611 (N_8611,N_5328,N_5952);
or U8612 (N_8612,N_5385,N_6585);
nor U8613 (N_8613,N_5850,N_6170);
or U8614 (N_8614,N_5284,N_6140);
or U8615 (N_8615,N_6325,N_5871);
nor U8616 (N_8616,N_7327,N_7293);
nand U8617 (N_8617,N_6724,N_6567);
nand U8618 (N_8618,N_6546,N_6313);
or U8619 (N_8619,N_6531,N_6856);
nand U8620 (N_8620,N_5417,N_7148);
or U8621 (N_8621,N_7251,N_6916);
or U8622 (N_8622,N_7240,N_5877);
and U8623 (N_8623,N_7236,N_6872);
nand U8624 (N_8624,N_5407,N_5231);
and U8625 (N_8625,N_5549,N_6961);
xor U8626 (N_8626,N_5590,N_6760);
nor U8627 (N_8627,N_5872,N_7112);
nor U8628 (N_8628,N_6112,N_6536);
and U8629 (N_8629,N_5444,N_6430);
or U8630 (N_8630,N_5582,N_5987);
and U8631 (N_8631,N_6047,N_5079);
or U8632 (N_8632,N_5904,N_7417);
nor U8633 (N_8633,N_6394,N_7487);
nor U8634 (N_8634,N_6538,N_5852);
and U8635 (N_8635,N_7459,N_7457);
and U8636 (N_8636,N_5599,N_7289);
or U8637 (N_8637,N_7234,N_5078);
nor U8638 (N_8638,N_5604,N_5697);
or U8639 (N_8639,N_7137,N_6910);
nor U8640 (N_8640,N_5299,N_6270);
or U8641 (N_8641,N_5638,N_7184);
and U8642 (N_8642,N_7254,N_5609);
and U8643 (N_8643,N_5256,N_6248);
and U8644 (N_8644,N_6122,N_6954);
nor U8645 (N_8645,N_6445,N_5007);
nand U8646 (N_8646,N_6223,N_6395);
or U8647 (N_8647,N_5863,N_5056);
or U8648 (N_8648,N_5884,N_6043);
or U8649 (N_8649,N_5605,N_5691);
and U8650 (N_8650,N_6945,N_6321);
nor U8651 (N_8651,N_6698,N_6656);
nor U8652 (N_8652,N_6877,N_6307);
or U8653 (N_8653,N_5830,N_7496);
or U8654 (N_8654,N_5068,N_5571);
nor U8655 (N_8655,N_7042,N_7257);
or U8656 (N_8656,N_6953,N_5695);
nor U8657 (N_8657,N_5460,N_6355);
nor U8658 (N_8658,N_6260,N_7246);
and U8659 (N_8659,N_7320,N_6908);
nor U8660 (N_8660,N_5138,N_6975);
and U8661 (N_8661,N_7229,N_5511);
nand U8662 (N_8662,N_6913,N_5520);
or U8663 (N_8663,N_7450,N_6350);
nand U8664 (N_8664,N_6615,N_6034);
or U8665 (N_8665,N_5178,N_5046);
and U8666 (N_8666,N_6829,N_6743);
nor U8667 (N_8667,N_6539,N_5077);
or U8668 (N_8668,N_6488,N_5708);
nor U8669 (N_8669,N_5103,N_7306);
nor U8670 (N_8670,N_7321,N_6976);
nor U8671 (N_8671,N_5016,N_5183);
and U8672 (N_8672,N_5997,N_6293);
or U8673 (N_8673,N_7154,N_5758);
nand U8674 (N_8674,N_6134,N_5286);
or U8675 (N_8675,N_6778,N_5037);
nor U8676 (N_8676,N_5008,N_6795);
and U8677 (N_8677,N_6273,N_6171);
nor U8678 (N_8678,N_5602,N_7201);
xor U8679 (N_8679,N_7098,N_6779);
nor U8680 (N_8680,N_5454,N_5002);
and U8681 (N_8681,N_6126,N_6169);
or U8682 (N_8682,N_6324,N_7309);
nor U8683 (N_8683,N_6026,N_6505);
or U8684 (N_8684,N_7258,N_6524);
nor U8685 (N_8685,N_5043,N_5613);
and U8686 (N_8686,N_6231,N_6370);
nand U8687 (N_8687,N_6790,N_6900);
and U8688 (N_8688,N_5115,N_5937);
nand U8689 (N_8689,N_6414,N_5128);
or U8690 (N_8690,N_5108,N_6695);
and U8691 (N_8691,N_7226,N_5857);
nor U8692 (N_8692,N_6019,N_5433);
and U8693 (N_8693,N_6641,N_5340);
nor U8694 (N_8694,N_6622,N_7371);
nor U8695 (N_8695,N_5035,N_5683);
nor U8696 (N_8696,N_6700,N_5268);
nand U8697 (N_8697,N_5546,N_6887);
nor U8698 (N_8698,N_7407,N_6373);
or U8699 (N_8699,N_5492,N_7102);
and U8700 (N_8700,N_5452,N_6983);
nor U8701 (N_8701,N_6885,N_5123);
xor U8702 (N_8702,N_6548,N_5261);
and U8703 (N_8703,N_7400,N_5809);
or U8704 (N_8704,N_6602,N_5554);
and U8705 (N_8705,N_6123,N_5424);
nor U8706 (N_8706,N_6341,N_5375);
and U8707 (N_8707,N_5501,N_5570);
xor U8708 (N_8708,N_5495,N_6484);
or U8709 (N_8709,N_6658,N_5067);
nand U8710 (N_8710,N_6024,N_5194);
nor U8711 (N_8711,N_5324,N_5616);
nand U8712 (N_8712,N_7314,N_5775);
and U8713 (N_8713,N_5709,N_5818);
nor U8714 (N_8714,N_6642,N_6015);
and U8715 (N_8715,N_5443,N_5298);
nand U8716 (N_8716,N_7182,N_5240);
nand U8717 (N_8717,N_6893,N_5860);
nand U8718 (N_8718,N_7436,N_5568);
and U8719 (N_8719,N_5026,N_5660);
and U8720 (N_8720,N_5624,N_7180);
nand U8721 (N_8721,N_7341,N_5772);
or U8722 (N_8722,N_6848,N_5247);
nor U8723 (N_8723,N_6914,N_6073);
and U8724 (N_8724,N_5516,N_5875);
and U8725 (N_8725,N_5164,N_6516);
nand U8726 (N_8726,N_6368,N_5864);
or U8727 (N_8727,N_5825,N_5988);
or U8728 (N_8728,N_5688,N_6308);
and U8729 (N_8729,N_5323,N_5858);
nand U8730 (N_8730,N_6391,N_6317);
nand U8731 (N_8731,N_7296,N_6443);
or U8732 (N_8732,N_5499,N_6670);
nor U8733 (N_8733,N_6940,N_6055);
nand U8734 (N_8734,N_6474,N_5326);
nor U8735 (N_8735,N_5839,N_7274);
nand U8736 (N_8736,N_5821,N_6752);
and U8737 (N_8737,N_5796,N_6483);
nand U8738 (N_8738,N_6587,N_6120);
or U8739 (N_8739,N_5515,N_5393);
nor U8740 (N_8740,N_5027,N_5432);
or U8741 (N_8741,N_6111,N_5981);
or U8742 (N_8742,N_6064,N_6755);
and U8743 (N_8743,N_6022,N_5453);
or U8744 (N_8744,N_5878,N_6657);
or U8745 (N_8745,N_6158,N_7356);
or U8746 (N_8746,N_7244,N_7194);
nor U8747 (N_8747,N_7248,N_5985);
nand U8748 (N_8748,N_5855,N_5637);
or U8749 (N_8749,N_5705,N_5730);
nand U8750 (N_8750,N_6124,N_6007);
nor U8751 (N_8751,N_7287,N_5221);
nor U8752 (N_8752,N_5761,N_5709);
or U8753 (N_8753,N_5087,N_7156);
nand U8754 (N_8754,N_5510,N_5920);
nand U8755 (N_8755,N_6951,N_6853);
and U8756 (N_8756,N_6160,N_6604);
and U8757 (N_8757,N_7252,N_7365);
nand U8758 (N_8758,N_5252,N_7318);
and U8759 (N_8759,N_6396,N_5303);
nand U8760 (N_8760,N_6242,N_6545);
or U8761 (N_8761,N_5140,N_6345);
nand U8762 (N_8762,N_5111,N_5208);
nand U8763 (N_8763,N_7364,N_5093);
or U8764 (N_8764,N_6833,N_7465);
nand U8765 (N_8765,N_5472,N_6023);
or U8766 (N_8766,N_5310,N_6518);
or U8767 (N_8767,N_6015,N_6713);
nor U8768 (N_8768,N_7056,N_7203);
or U8769 (N_8769,N_6476,N_7355);
and U8770 (N_8770,N_7165,N_6854);
and U8771 (N_8771,N_5633,N_5876);
and U8772 (N_8772,N_5788,N_5380);
nor U8773 (N_8773,N_5987,N_7263);
nand U8774 (N_8774,N_6649,N_5409);
nor U8775 (N_8775,N_5793,N_6014);
nor U8776 (N_8776,N_5008,N_7275);
nor U8777 (N_8777,N_5034,N_6951);
or U8778 (N_8778,N_5949,N_5584);
or U8779 (N_8779,N_6022,N_5369);
nand U8780 (N_8780,N_7393,N_7071);
and U8781 (N_8781,N_6956,N_5941);
nor U8782 (N_8782,N_5617,N_5476);
nor U8783 (N_8783,N_5942,N_6887);
or U8784 (N_8784,N_7262,N_6106);
or U8785 (N_8785,N_5516,N_5822);
nor U8786 (N_8786,N_5173,N_5426);
and U8787 (N_8787,N_6435,N_6113);
and U8788 (N_8788,N_7345,N_5562);
or U8789 (N_8789,N_5942,N_6111);
nor U8790 (N_8790,N_6518,N_5150);
and U8791 (N_8791,N_5766,N_5755);
and U8792 (N_8792,N_5711,N_5876);
or U8793 (N_8793,N_5201,N_5932);
nor U8794 (N_8794,N_6235,N_6488);
xnor U8795 (N_8795,N_7195,N_5911);
nor U8796 (N_8796,N_7290,N_5530);
and U8797 (N_8797,N_5616,N_6891);
nor U8798 (N_8798,N_5479,N_6574);
nand U8799 (N_8799,N_5481,N_6574);
or U8800 (N_8800,N_6772,N_5904);
or U8801 (N_8801,N_5789,N_6428);
nor U8802 (N_8802,N_5427,N_6117);
or U8803 (N_8803,N_6934,N_6384);
nand U8804 (N_8804,N_6482,N_6489);
nand U8805 (N_8805,N_5347,N_5085);
and U8806 (N_8806,N_7178,N_7176);
or U8807 (N_8807,N_5380,N_6753);
nor U8808 (N_8808,N_7380,N_5865);
or U8809 (N_8809,N_6504,N_5990);
and U8810 (N_8810,N_7152,N_5437);
and U8811 (N_8811,N_6934,N_7040);
nand U8812 (N_8812,N_5521,N_6337);
nor U8813 (N_8813,N_7359,N_5469);
xnor U8814 (N_8814,N_6070,N_5174);
nor U8815 (N_8815,N_6324,N_5651);
or U8816 (N_8816,N_5557,N_6459);
and U8817 (N_8817,N_7350,N_5262);
or U8818 (N_8818,N_5145,N_5571);
nor U8819 (N_8819,N_6789,N_7186);
or U8820 (N_8820,N_5010,N_7209);
nor U8821 (N_8821,N_5430,N_7068);
and U8822 (N_8822,N_6818,N_6688);
nand U8823 (N_8823,N_5080,N_5793);
nand U8824 (N_8824,N_7260,N_5678);
nand U8825 (N_8825,N_5757,N_5716);
nor U8826 (N_8826,N_5383,N_6048);
nor U8827 (N_8827,N_6873,N_6690);
or U8828 (N_8828,N_5708,N_6444);
nand U8829 (N_8829,N_6901,N_7493);
nand U8830 (N_8830,N_6346,N_5681);
and U8831 (N_8831,N_6299,N_7257);
or U8832 (N_8832,N_7104,N_6032);
nor U8833 (N_8833,N_5954,N_6174);
xnor U8834 (N_8834,N_5837,N_5827);
nand U8835 (N_8835,N_5682,N_5043);
nor U8836 (N_8836,N_6695,N_6521);
and U8837 (N_8837,N_5545,N_5019);
nor U8838 (N_8838,N_5375,N_6385);
or U8839 (N_8839,N_7420,N_5565);
and U8840 (N_8840,N_7214,N_6642);
nor U8841 (N_8841,N_5863,N_7243);
xnor U8842 (N_8842,N_6358,N_5579);
nand U8843 (N_8843,N_7486,N_5699);
nand U8844 (N_8844,N_6630,N_5664);
or U8845 (N_8845,N_5232,N_5245);
nor U8846 (N_8846,N_5063,N_7162);
nand U8847 (N_8847,N_6586,N_7350);
and U8848 (N_8848,N_5679,N_5113);
or U8849 (N_8849,N_5047,N_7210);
or U8850 (N_8850,N_7253,N_5706);
and U8851 (N_8851,N_5019,N_6124);
and U8852 (N_8852,N_5546,N_6838);
nor U8853 (N_8853,N_6057,N_6437);
and U8854 (N_8854,N_6947,N_5677);
nor U8855 (N_8855,N_6960,N_5740);
nand U8856 (N_8856,N_5467,N_6768);
nor U8857 (N_8857,N_6026,N_5215);
and U8858 (N_8858,N_5907,N_6936);
nand U8859 (N_8859,N_5059,N_6341);
nand U8860 (N_8860,N_5768,N_6482);
and U8861 (N_8861,N_6862,N_5694);
nor U8862 (N_8862,N_6163,N_6653);
nand U8863 (N_8863,N_6257,N_6754);
or U8864 (N_8864,N_5280,N_5315);
and U8865 (N_8865,N_5339,N_6641);
and U8866 (N_8866,N_5537,N_5916);
and U8867 (N_8867,N_6202,N_5598);
or U8868 (N_8868,N_6503,N_5504);
nor U8869 (N_8869,N_6578,N_5307);
and U8870 (N_8870,N_7133,N_7305);
or U8871 (N_8871,N_6791,N_5818);
or U8872 (N_8872,N_5047,N_5779);
nand U8873 (N_8873,N_7438,N_7298);
and U8874 (N_8874,N_5028,N_6489);
nor U8875 (N_8875,N_5614,N_6233);
or U8876 (N_8876,N_5403,N_7082);
or U8877 (N_8877,N_5764,N_5003);
or U8878 (N_8878,N_6107,N_5564);
or U8879 (N_8879,N_6810,N_5638);
nor U8880 (N_8880,N_6252,N_7459);
or U8881 (N_8881,N_5229,N_6305);
nor U8882 (N_8882,N_5835,N_6546);
nor U8883 (N_8883,N_6729,N_6417);
and U8884 (N_8884,N_7467,N_5266);
and U8885 (N_8885,N_6691,N_6991);
or U8886 (N_8886,N_5865,N_6389);
nor U8887 (N_8887,N_6048,N_7228);
nand U8888 (N_8888,N_5006,N_5665);
nand U8889 (N_8889,N_6019,N_6935);
or U8890 (N_8890,N_5579,N_7472);
nor U8891 (N_8891,N_7200,N_5112);
or U8892 (N_8892,N_5685,N_6362);
nor U8893 (N_8893,N_5400,N_6921);
nor U8894 (N_8894,N_7178,N_7405);
nand U8895 (N_8895,N_5884,N_5306);
and U8896 (N_8896,N_5025,N_5045);
or U8897 (N_8897,N_6011,N_5615);
and U8898 (N_8898,N_5214,N_6942);
nor U8899 (N_8899,N_5479,N_5937);
nor U8900 (N_8900,N_6135,N_6391);
or U8901 (N_8901,N_7349,N_5153);
or U8902 (N_8902,N_6446,N_6046);
nand U8903 (N_8903,N_6905,N_5742);
nand U8904 (N_8904,N_5378,N_7489);
nor U8905 (N_8905,N_6691,N_5236);
or U8906 (N_8906,N_6821,N_5720);
and U8907 (N_8907,N_5928,N_6028);
nor U8908 (N_8908,N_5084,N_5611);
nand U8909 (N_8909,N_6292,N_5024);
nor U8910 (N_8910,N_6940,N_6302);
or U8911 (N_8911,N_5756,N_6147);
and U8912 (N_8912,N_6419,N_6528);
or U8913 (N_8913,N_7187,N_5934);
and U8914 (N_8914,N_6033,N_5539);
nand U8915 (N_8915,N_7417,N_5305);
nand U8916 (N_8916,N_6172,N_5944);
or U8917 (N_8917,N_5530,N_5894);
or U8918 (N_8918,N_6180,N_5661);
nor U8919 (N_8919,N_5792,N_5353);
xor U8920 (N_8920,N_5117,N_5650);
nor U8921 (N_8921,N_6334,N_7006);
nand U8922 (N_8922,N_5269,N_5604);
and U8923 (N_8923,N_6005,N_5824);
nand U8924 (N_8924,N_7400,N_5890);
nand U8925 (N_8925,N_7416,N_5365);
nand U8926 (N_8926,N_7288,N_6683);
or U8927 (N_8927,N_5337,N_6807);
or U8928 (N_8928,N_7041,N_5726);
nor U8929 (N_8929,N_6923,N_5425);
and U8930 (N_8930,N_5692,N_7212);
or U8931 (N_8931,N_7486,N_5707);
nand U8932 (N_8932,N_5811,N_7276);
or U8933 (N_8933,N_6215,N_7138);
nor U8934 (N_8934,N_5630,N_6893);
nor U8935 (N_8935,N_6938,N_5917);
and U8936 (N_8936,N_7320,N_6256);
nand U8937 (N_8937,N_6521,N_6690);
nor U8938 (N_8938,N_6416,N_5057);
or U8939 (N_8939,N_5107,N_5189);
or U8940 (N_8940,N_5134,N_7277);
nor U8941 (N_8941,N_6019,N_7450);
or U8942 (N_8942,N_5896,N_5529);
or U8943 (N_8943,N_6206,N_5691);
nand U8944 (N_8944,N_6801,N_5025);
or U8945 (N_8945,N_5206,N_5575);
and U8946 (N_8946,N_7217,N_6070);
and U8947 (N_8947,N_5644,N_7400);
nand U8948 (N_8948,N_6280,N_6533);
nor U8949 (N_8949,N_6902,N_6025);
nor U8950 (N_8950,N_6768,N_6490);
and U8951 (N_8951,N_5447,N_6528);
or U8952 (N_8952,N_6740,N_5768);
nand U8953 (N_8953,N_7421,N_6707);
nand U8954 (N_8954,N_5716,N_7403);
or U8955 (N_8955,N_7096,N_6226);
nand U8956 (N_8956,N_6212,N_6249);
and U8957 (N_8957,N_7193,N_6336);
and U8958 (N_8958,N_6915,N_5648);
or U8959 (N_8959,N_7165,N_5779);
nand U8960 (N_8960,N_5349,N_5390);
nor U8961 (N_8961,N_6477,N_6706);
or U8962 (N_8962,N_6584,N_6347);
and U8963 (N_8963,N_5767,N_6972);
or U8964 (N_8964,N_6675,N_5630);
nand U8965 (N_8965,N_5312,N_6493);
and U8966 (N_8966,N_6273,N_7478);
or U8967 (N_8967,N_6235,N_7002);
and U8968 (N_8968,N_5139,N_7326);
nand U8969 (N_8969,N_5950,N_5929);
or U8970 (N_8970,N_5932,N_6101);
nand U8971 (N_8971,N_5471,N_5288);
or U8972 (N_8972,N_5584,N_6267);
or U8973 (N_8973,N_6168,N_6924);
nand U8974 (N_8974,N_5790,N_7082);
nand U8975 (N_8975,N_7111,N_7022);
nor U8976 (N_8976,N_5322,N_5456);
nand U8977 (N_8977,N_5405,N_5205);
nor U8978 (N_8978,N_7096,N_7143);
nor U8979 (N_8979,N_5075,N_5635);
nand U8980 (N_8980,N_6077,N_5477);
nor U8981 (N_8981,N_6064,N_6214);
or U8982 (N_8982,N_6153,N_6562);
xor U8983 (N_8983,N_6270,N_6129);
nand U8984 (N_8984,N_6001,N_5526);
and U8985 (N_8985,N_7276,N_7088);
nor U8986 (N_8986,N_6795,N_5474);
nand U8987 (N_8987,N_5004,N_5657);
or U8988 (N_8988,N_7444,N_5644);
nor U8989 (N_8989,N_6349,N_6256);
or U8990 (N_8990,N_5530,N_6657);
nor U8991 (N_8991,N_5042,N_5450);
nor U8992 (N_8992,N_6650,N_5611);
nor U8993 (N_8993,N_6292,N_6262);
and U8994 (N_8994,N_6910,N_5632);
and U8995 (N_8995,N_6508,N_6057);
and U8996 (N_8996,N_5435,N_6707);
or U8997 (N_8997,N_6202,N_5494);
or U8998 (N_8998,N_6948,N_5840);
nand U8999 (N_8999,N_5403,N_5716);
nor U9000 (N_9000,N_7040,N_6186);
and U9001 (N_9001,N_6084,N_5701);
nand U9002 (N_9002,N_5189,N_7293);
nor U9003 (N_9003,N_6172,N_6269);
and U9004 (N_9004,N_6624,N_7162);
nor U9005 (N_9005,N_5157,N_5682);
and U9006 (N_9006,N_7433,N_6541);
nand U9007 (N_9007,N_5070,N_6764);
and U9008 (N_9008,N_6088,N_6770);
or U9009 (N_9009,N_5155,N_5306);
nor U9010 (N_9010,N_5154,N_6421);
or U9011 (N_9011,N_5612,N_5423);
nand U9012 (N_9012,N_5079,N_7103);
nor U9013 (N_9013,N_7290,N_6339);
nor U9014 (N_9014,N_5803,N_6348);
or U9015 (N_9015,N_6111,N_7312);
or U9016 (N_9016,N_6184,N_5308);
and U9017 (N_9017,N_6691,N_5170);
nand U9018 (N_9018,N_5384,N_7080);
or U9019 (N_9019,N_6298,N_7064);
nand U9020 (N_9020,N_6176,N_5600);
and U9021 (N_9021,N_5860,N_5726);
nand U9022 (N_9022,N_5476,N_7368);
nor U9023 (N_9023,N_6012,N_5716);
and U9024 (N_9024,N_7171,N_6678);
nor U9025 (N_9025,N_5163,N_5966);
and U9026 (N_9026,N_7439,N_5124);
nand U9027 (N_9027,N_5684,N_5058);
nand U9028 (N_9028,N_6790,N_5138);
and U9029 (N_9029,N_6946,N_6998);
nand U9030 (N_9030,N_5463,N_6709);
nor U9031 (N_9031,N_5741,N_6254);
or U9032 (N_9032,N_7216,N_5948);
and U9033 (N_9033,N_5778,N_5600);
nor U9034 (N_9034,N_6335,N_6603);
or U9035 (N_9035,N_6262,N_6153);
and U9036 (N_9036,N_5322,N_6599);
nor U9037 (N_9037,N_6308,N_6465);
or U9038 (N_9038,N_7457,N_6207);
and U9039 (N_9039,N_6287,N_7398);
and U9040 (N_9040,N_6240,N_6494);
and U9041 (N_9041,N_5742,N_5739);
nand U9042 (N_9042,N_5613,N_5767);
and U9043 (N_9043,N_5116,N_5188);
nor U9044 (N_9044,N_7388,N_5564);
or U9045 (N_9045,N_6520,N_6774);
and U9046 (N_9046,N_5232,N_6117);
nand U9047 (N_9047,N_5854,N_7276);
nand U9048 (N_9048,N_6346,N_5357);
and U9049 (N_9049,N_6497,N_5383);
nand U9050 (N_9050,N_5611,N_7414);
or U9051 (N_9051,N_7154,N_5936);
nor U9052 (N_9052,N_7080,N_7356);
or U9053 (N_9053,N_6276,N_6999);
and U9054 (N_9054,N_6187,N_6161);
and U9055 (N_9055,N_6487,N_6524);
and U9056 (N_9056,N_5883,N_6689);
nand U9057 (N_9057,N_6069,N_6851);
or U9058 (N_9058,N_5361,N_5306);
or U9059 (N_9059,N_7169,N_5321);
and U9060 (N_9060,N_5910,N_7424);
and U9061 (N_9061,N_6515,N_6345);
or U9062 (N_9062,N_6943,N_6018);
and U9063 (N_9063,N_7272,N_6408);
nand U9064 (N_9064,N_7244,N_7321);
nand U9065 (N_9065,N_6908,N_5404);
and U9066 (N_9066,N_6551,N_6286);
nor U9067 (N_9067,N_5228,N_5292);
nor U9068 (N_9068,N_6196,N_6832);
and U9069 (N_9069,N_6902,N_5913);
and U9070 (N_9070,N_6576,N_6218);
nand U9071 (N_9071,N_7272,N_6551);
nor U9072 (N_9072,N_6779,N_6234);
and U9073 (N_9073,N_6122,N_7154);
nand U9074 (N_9074,N_5903,N_5657);
or U9075 (N_9075,N_5286,N_6976);
nor U9076 (N_9076,N_6642,N_6513);
and U9077 (N_9077,N_7105,N_6723);
or U9078 (N_9078,N_6248,N_5732);
or U9079 (N_9079,N_7276,N_6374);
and U9080 (N_9080,N_5274,N_6612);
nor U9081 (N_9081,N_5796,N_5510);
or U9082 (N_9082,N_5106,N_6356);
nand U9083 (N_9083,N_7237,N_7362);
nand U9084 (N_9084,N_7426,N_5899);
and U9085 (N_9085,N_7094,N_6229);
and U9086 (N_9086,N_5244,N_5778);
nor U9087 (N_9087,N_6398,N_5121);
nor U9088 (N_9088,N_5914,N_5660);
nor U9089 (N_9089,N_7191,N_5562);
nor U9090 (N_9090,N_5160,N_5570);
nand U9091 (N_9091,N_6447,N_6970);
and U9092 (N_9092,N_6644,N_6176);
nand U9093 (N_9093,N_6072,N_6876);
nand U9094 (N_9094,N_7468,N_6830);
nand U9095 (N_9095,N_6080,N_5518);
and U9096 (N_9096,N_6163,N_5715);
and U9097 (N_9097,N_6726,N_5500);
nand U9098 (N_9098,N_6505,N_7167);
nor U9099 (N_9099,N_7260,N_5137);
and U9100 (N_9100,N_5139,N_7498);
nand U9101 (N_9101,N_6350,N_5961);
and U9102 (N_9102,N_6993,N_5268);
and U9103 (N_9103,N_7080,N_5709);
or U9104 (N_9104,N_5101,N_7408);
nor U9105 (N_9105,N_6035,N_5662);
xnor U9106 (N_9106,N_6256,N_5027);
nor U9107 (N_9107,N_5388,N_7010);
and U9108 (N_9108,N_7093,N_5002);
or U9109 (N_9109,N_5928,N_5485);
nor U9110 (N_9110,N_5942,N_6526);
nor U9111 (N_9111,N_5666,N_5877);
or U9112 (N_9112,N_5987,N_5393);
and U9113 (N_9113,N_6835,N_6368);
or U9114 (N_9114,N_6334,N_7266);
and U9115 (N_9115,N_7044,N_5610);
and U9116 (N_9116,N_5564,N_6299);
xor U9117 (N_9117,N_6403,N_6785);
or U9118 (N_9118,N_5829,N_5671);
and U9119 (N_9119,N_6047,N_7077);
nand U9120 (N_9120,N_5702,N_5636);
nand U9121 (N_9121,N_5750,N_6596);
or U9122 (N_9122,N_5881,N_6984);
and U9123 (N_9123,N_6746,N_5903);
or U9124 (N_9124,N_6496,N_6730);
nor U9125 (N_9125,N_5682,N_5938);
and U9126 (N_9126,N_5013,N_6177);
and U9127 (N_9127,N_5819,N_6606);
or U9128 (N_9128,N_5441,N_6436);
or U9129 (N_9129,N_5087,N_6810);
nand U9130 (N_9130,N_5378,N_5825);
and U9131 (N_9131,N_6706,N_6308);
nand U9132 (N_9132,N_5136,N_5784);
nor U9133 (N_9133,N_5366,N_5604);
or U9134 (N_9134,N_6019,N_6073);
nor U9135 (N_9135,N_5349,N_5962);
or U9136 (N_9136,N_6805,N_5379);
or U9137 (N_9137,N_6579,N_5213);
nand U9138 (N_9138,N_7045,N_6415);
nor U9139 (N_9139,N_6799,N_5091);
and U9140 (N_9140,N_6096,N_6519);
and U9141 (N_9141,N_7133,N_5747);
nand U9142 (N_9142,N_7257,N_5893);
nor U9143 (N_9143,N_5851,N_6043);
and U9144 (N_9144,N_5159,N_7228);
and U9145 (N_9145,N_5777,N_5638);
and U9146 (N_9146,N_7123,N_6696);
nor U9147 (N_9147,N_6124,N_5286);
nor U9148 (N_9148,N_6022,N_6907);
nand U9149 (N_9149,N_6570,N_6554);
nor U9150 (N_9150,N_5046,N_6659);
or U9151 (N_9151,N_6715,N_5051);
and U9152 (N_9152,N_6657,N_7486);
or U9153 (N_9153,N_5490,N_6490);
nand U9154 (N_9154,N_5628,N_6452);
nand U9155 (N_9155,N_7025,N_7090);
nand U9156 (N_9156,N_6861,N_7141);
or U9157 (N_9157,N_5886,N_5234);
nand U9158 (N_9158,N_5143,N_5597);
and U9159 (N_9159,N_6958,N_7129);
nand U9160 (N_9160,N_6050,N_6226);
nor U9161 (N_9161,N_5285,N_6784);
and U9162 (N_9162,N_6235,N_7324);
or U9163 (N_9163,N_5153,N_5752);
or U9164 (N_9164,N_5357,N_5940);
nand U9165 (N_9165,N_6623,N_5636);
or U9166 (N_9166,N_7383,N_6221);
xor U9167 (N_9167,N_6885,N_5874);
nor U9168 (N_9168,N_5407,N_5133);
nand U9169 (N_9169,N_6817,N_6885);
and U9170 (N_9170,N_6418,N_6156);
nand U9171 (N_9171,N_6731,N_5043);
nand U9172 (N_9172,N_6576,N_5641);
nor U9173 (N_9173,N_7431,N_7104);
nand U9174 (N_9174,N_6257,N_5495);
or U9175 (N_9175,N_5505,N_5359);
and U9176 (N_9176,N_5318,N_5761);
or U9177 (N_9177,N_6041,N_6751);
or U9178 (N_9178,N_6510,N_7352);
and U9179 (N_9179,N_5369,N_5466);
nand U9180 (N_9180,N_5403,N_5287);
or U9181 (N_9181,N_6456,N_6935);
nor U9182 (N_9182,N_7471,N_6094);
or U9183 (N_9183,N_7421,N_7262);
nor U9184 (N_9184,N_6652,N_6526);
or U9185 (N_9185,N_7339,N_6198);
and U9186 (N_9186,N_5931,N_7368);
nor U9187 (N_9187,N_5388,N_6913);
nor U9188 (N_9188,N_5083,N_7180);
nor U9189 (N_9189,N_7435,N_5770);
and U9190 (N_9190,N_6454,N_6674);
or U9191 (N_9191,N_6702,N_6622);
nor U9192 (N_9192,N_5139,N_5142);
or U9193 (N_9193,N_6504,N_7150);
nand U9194 (N_9194,N_7090,N_7486);
and U9195 (N_9195,N_7036,N_6605);
or U9196 (N_9196,N_6345,N_6992);
nand U9197 (N_9197,N_7413,N_7334);
nor U9198 (N_9198,N_5740,N_5842);
and U9199 (N_9199,N_6707,N_6343);
nor U9200 (N_9200,N_6630,N_5534);
and U9201 (N_9201,N_5194,N_7014);
and U9202 (N_9202,N_7077,N_5827);
nor U9203 (N_9203,N_6049,N_5638);
or U9204 (N_9204,N_5922,N_6735);
nor U9205 (N_9205,N_6922,N_6915);
nand U9206 (N_9206,N_7308,N_5445);
and U9207 (N_9207,N_6046,N_6291);
and U9208 (N_9208,N_6629,N_7459);
nand U9209 (N_9209,N_6025,N_6648);
or U9210 (N_9210,N_6706,N_7409);
nor U9211 (N_9211,N_6287,N_7438);
and U9212 (N_9212,N_5301,N_6030);
or U9213 (N_9213,N_5674,N_7365);
nand U9214 (N_9214,N_5523,N_7464);
and U9215 (N_9215,N_5943,N_5061);
and U9216 (N_9216,N_7178,N_5436);
nor U9217 (N_9217,N_5565,N_7072);
xnor U9218 (N_9218,N_5007,N_5414);
nand U9219 (N_9219,N_6891,N_6220);
or U9220 (N_9220,N_7049,N_5190);
or U9221 (N_9221,N_7345,N_6365);
or U9222 (N_9222,N_7298,N_6060);
nand U9223 (N_9223,N_6602,N_7225);
nor U9224 (N_9224,N_6478,N_6721);
and U9225 (N_9225,N_6789,N_6715);
nor U9226 (N_9226,N_5862,N_5456);
or U9227 (N_9227,N_6672,N_6300);
and U9228 (N_9228,N_5728,N_6563);
xor U9229 (N_9229,N_6528,N_5226);
and U9230 (N_9230,N_6506,N_6464);
or U9231 (N_9231,N_7237,N_6606);
or U9232 (N_9232,N_5446,N_5616);
nand U9233 (N_9233,N_5701,N_7421);
and U9234 (N_9234,N_5524,N_5144);
nand U9235 (N_9235,N_5397,N_5277);
or U9236 (N_9236,N_5500,N_7323);
nor U9237 (N_9237,N_6359,N_6517);
nor U9238 (N_9238,N_5573,N_5980);
and U9239 (N_9239,N_7039,N_6766);
nand U9240 (N_9240,N_5140,N_7002);
xor U9241 (N_9241,N_7117,N_6853);
and U9242 (N_9242,N_6129,N_5896);
nand U9243 (N_9243,N_6821,N_5129);
and U9244 (N_9244,N_6840,N_5962);
nor U9245 (N_9245,N_6586,N_6712);
nor U9246 (N_9246,N_7018,N_6016);
nand U9247 (N_9247,N_7205,N_5911);
and U9248 (N_9248,N_5822,N_6098);
nand U9249 (N_9249,N_6484,N_7155);
or U9250 (N_9250,N_5759,N_5479);
nor U9251 (N_9251,N_5550,N_7330);
and U9252 (N_9252,N_5474,N_5655);
or U9253 (N_9253,N_7187,N_5290);
nor U9254 (N_9254,N_6223,N_5576);
and U9255 (N_9255,N_7124,N_7237);
nand U9256 (N_9256,N_7127,N_5347);
and U9257 (N_9257,N_5509,N_6960);
and U9258 (N_9258,N_5366,N_6275);
or U9259 (N_9259,N_5984,N_6069);
nor U9260 (N_9260,N_7330,N_6971);
or U9261 (N_9261,N_6805,N_6251);
nor U9262 (N_9262,N_6962,N_5626);
or U9263 (N_9263,N_7109,N_7456);
nor U9264 (N_9264,N_5610,N_6504);
and U9265 (N_9265,N_5276,N_6801);
or U9266 (N_9266,N_7080,N_6841);
nand U9267 (N_9267,N_7175,N_6944);
nand U9268 (N_9268,N_7336,N_6891);
or U9269 (N_9269,N_5935,N_7392);
nor U9270 (N_9270,N_6812,N_5957);
nand U9271 (N_9271,N_5844,N_6643);
nor U9272 (N_9272,N_7281,N_6891);
nand U9273 (N_9273,N_7332,N_5916);
or U9274 (N_9274,N_6404,N_6402);
nand U9275 (N_9275,N_6266,N_5066);
and U9276 (N_9276,N_6630,N_6655);
nand U9277 (N_9277,N_5274,N_6251);
or U9278 (N_9278,N_6757,N_6062);
nor U9279 (N_9279,N_5440,N_6260);
nand U9280 (N_9280,N_5922,N_7202);
or U9281 (N_9281,N_6646,N_5285);
and U9282 (N_9282,N_6173,N_6767);
and U9283 (N_9283,N_6686,N_7205);
and U9284 (N_9284,N_5644,N_5252);
nor U9285 (N_9285,N_6785,N_6316);
or U9286 (N_9286,N_6369,N_7430);
nand U9287 (N_9287,N_7390,N_6737);
or U9288 (N_9288,N_6829,N_5055);
and U9289 (N_9289,N_5489,N_6561);
nor U9290 (N_9290,N_6456,N_5056);
nand U9291 (N_9291,N_5675,N_6212);
nand U9292 (N_9292,N_5201,N_6049);
or U9293 (N_9293,N_5468,N_5647);
nor U9294 (N_9294,N_5003,N_5438);
or U9295 (N_9295,N_5825,N_7454);
or U9296 (N_9296,N_5168,N_6282);
nor U9297 (N_9297,N_6401,N_6055);
or U9298 (N_9298,N_5997,N_6418);
nand U9299 (N_9299,N_7294,N_5076);
nor U9300 (N_9300,N_6759,N_5620);
xnor U9301 (N_9301,N_7380,N_5387);
or U9302 (N_9302,N_7262,N_5951);
nand U9303 (N_9303,N_7206,N_6343);
and U9304 (N_9304,N_6289,N_6535);
nor U9305 (N_9305,N_6431,N_5455);
or U9306 (N_9306,N_6928,N_5075);
or U9307 (N_9307,N_7190,N_6085);
nor U9308 (N_9308,N_6372,N_5812);
or U9309 (N_9309,N_7167,N_6313);
or U9310 (N_9310,N_7457,N_5399);
nor U9311 (N_9311,N_5124,N_5245);
or U9312 (N_9312,N_7003,N_6759);
and U9313 (N_9313,N_6265,N_5188);
nor U9314 (N_9314,N_5899,N_5623);
nor U9315 (N_9315,N_5445,N_5714);
nand U9316 (N_9316,N_7319,N_5532);
and U9317 (N_9317,N_5777,N_7490);
and U9318 (N_9318,N_6054,N_7266);
nor U9319 (N_9319,N_5234,N_6839);
nand U9320 (N_9320,N_6605,N_6433);
and U9321 (N_9321,N_6064,N_5921);
and U9322 (N_9322,N_5831,N_6500);
nor U9323 (N_9323,N_5492,N_5471);
nor U9324 (N_9324,N_6695,N_6944);
nor U9325 (N_9325,N_6815,N_5426);
nand U9326 (N_9326,N_5870,N_6389);
nand U9327 (N_9327,N_7420,N_6539);
nand U9328 (N_9328,N_5142,N_6441);
nand U9329 (N_9329,N_6348,N_7284);
nand U9330 (N_9330,N_5806,N_7099);
and U9331 (N_9331,N_7444,N_6016);
nand U9332 (N_9332,N_6813,N_7251);
and U9333 (N_9333,N_6086,N_6950);
nor U9334 (N_9334,N_5672,N_5130);
or U9335 (N_9335,N_5081,N_5187);
nor U9336 (N_9336,N_7375,N_5299);
or U9337 (N_9337,N_6439,N_5819);
and U9338 (N_9338,N_7174,N_5471);
or U9339 (N_9339,N_7288,N_7345);
nor U9340 (N_9340,N_6240,N_6456);
nor U9341 (N_9341,N_5292,N_5304);
nor U9342 (N_9342,N_6013,N_5422);
nor U9343 (N_9343,N_6583,N_6358);
or U9344 (N_9344,N_5465,N_6585);
or U9345 (N_9345,N_7263,N_7014);
nor U9346 (N_9346,N_5131,N_6749);
nand U9347 (N_9347,N_5221,N_5230);
or U9348 (N_9348,N_6531,N_5588);
nand U9349 (N_9349,N_5846,N_5877);
nand U9350 (N_9350,N_6576,N_7159);
nor U9351 (N_9351,N_6349,N_6124);
nor U9352 (N_9352,N_6593,N_7274);
or U9353 (N_9353,N_5130,N_5746);
nor U9354 (N_9354,N_6634,N_5545);
nand U9355 (N_9355,N_5846,N_7015);
nand U9356 (N_9356,N_7262,N_6561);
or U9357 (N_9357,N_6435,N_6484);
xor U9358 (N_9358,N_5207,N_7248);
and U9359 (N_9359,N_7314,N_6504);
nor U9360 (N_9360,N_7140,N_7393);
and U9361 (N_9361,N_6507,N_5203);
nand U9362 (N_9362,N_5472,N_6747);
or U9363 (N_9363,N_6273,N_7365);
or U9364 (N_9364,N_5835,N_7016);
and U9365 (N_9365,N_6397,N_6931);
or U9366 (N_9366,N_7015,N_6319);
and U9367 (N_9367,N_6853,N_7360);
and U9368 (N_9368,N_5675,N_5857);
or U9369 (N_9369,N_6452,N_7428);
and U9370 (N_9370,N_6726,N_5172);
nor U9371 (N_9371,N_6939,N_7346);
or U9372 (N_9372,N_6068,N_7043);
nor U9373 (N_9373,N_5691,N_6768);
and U9374 (N_9374,N_7438,N_5380);
nor U9375 (N_9375,N_7137,N_7051);
and U9376 (N_9376,N_6784,N_5257);
or U9377 (N_9377,N_6341,N_6728);
or U9378 (N_9378,N_6605,N_7072);
xnor U9379 (N_9379,N_6142,N_6898);
or U9380 (N_9380,N_6890,N_5506);
nand U9381 (N_9381,N_7049,N_6685);
or U9382 (N_9382,N_5324,N_6825);
nor U9383 (N_9383,N_7183,N_5587);
and U9384 (N_9384,N_7164,N_5139);
nor U9385 (N_9385,N_7381,N_7300);
and U9386 (N_9386,N_6679,N_7387);
or U9387 (N_9387,N_6061,N_5043);
or U9388 (N_9388,N_5925,N_5843);
nand U9389 (N_9389,N_7221,N_6458);
and U9390 (N_9390,N_5074,N_6746);
nor U9391 (N_9391,N_7007,N_7407);
or U9392 (N_9392,N_6914,N_7437);
nor U9393 (N_9393,N_6269,N_7401);
and U9394 (N_9394,N_5534,N_6059);
and U9395 (N_9395,N_5177,N_5403);
nand U9396 (N_9396,N_5768,N_5187);
and U9397 (N_9397,N_5965,N_6499);
and U9398 (N_9398,N_5774,N_7379);
nand U9399 (N_9399,N_5412,N_6534);
and U9400 (N_9400,N_5832,N_5873);
nand U9401 (N_9401,N_6351,N_5644);
and U9402 (N_9402,N_5838,N_6328);
nand U9403 (N_9403,N_5594,N_5234);
nor U9404 (N_9404,N_6430,N_5137);
or U9405 (N_9405,N_5610,N_5776);
and U9406 (N_9406,N_5201,N_6534);
nor U9407 (N_9407,N_6065,N_5069);
nor U9408 (N_9408,N_7074,N_6999);
or U9409 (N_9409,N_6534,N_6516);
nor U9410 (N_9410,N_6435,N_7326);
and U9411 (N_9411,N_5781,N_7461);
and U9412 (N_9412,N_6074,N_6580);
nor U9413 (N_9413,N_7241,N_5387);
nor U9414 (N_9414,N_5345,N_6327);
nor U9415 (N_9415,N_5960,N_5799);
or U9416 (N_9416,N_6742,N_6789);
nor U9417 (N_9417,N_6405,N_5613);
nand U9418 (N_9418,N_6801,N_6052);
and U9419 (N_9419,N_5665,N_5325);
nand U9420 (N_9420,N_6374,N_6743);
nor U9421 (N_9421,N_6390,N_7484);
or U9422 (N_9422,N_7358,N_5105);
and U9423 (N_9423,N_5172,N_6509);
nand U9424 (N_9424,N_6251,N_6886);
or U9425 (N_9425,N_7064,N_5973);
nor U9426 (N_9426,N_5143,N_6052);
nand U9427 (N_9427,N_7173,N_6466);
and U9428 (N_9428,N_5875,N_6707);
or U9429 (N_9429,N_7498,N_5212);
or U9430 (N_9430,N_6939,N_6002);
nor U9431 (N_9431,N_6950,N_5762);
nor U9432 (N_9432,N_7124,N_7290);
nor U9433 (N_9433,N_7017,N_6695);
and U9434 (N_9434,N_6641,N_5890);
or U9435 (N_9435,N_5068,N_6971);
or U9436 (N_9436,N_6107,N_7221);
nor U9437 (N_9437,N_6306,N_5761);
nor U9438 (N_9438,N_5945,N_6672);
and U9439 (N_9439,N_6685,N_6985);
nor U9440 (N_9440,N_6910,N_6463);
nor U9441 (N_9441,N_7279,N_7137);
and U9442 (N_9442,N_5403,N_6491);
or U9443 (N_9443,N_5931,N_5626);
and U9444 (N_9444,N_7427,N_5467);
nand U9445 (N_9445,N_6549,N_6567);
nand U9446 (N_9446,N_7069,N_7187);
nand U9447 (N_9447,N_5173,N_6793);
nand U9448 (N_9448,N_6331,N_6072);
nand U9449 (N_9449,N_6314,N_6736);
nand U9450 (N_9450,N_5294,N_6970);
xnor U9451 (N_9451,N_7359,N_6001);
and U9452 (N_9452,N_7410,N_5509);
or U9453 (N_9453,N_6334,N_7260);
nand U9454 (N_9454,N_6333,N_7272);
and U9455 (N_9455,N_7028,N_6037);
nor U9456 (N_9456,N_6218,N_6984);
nand U9457 (N_9457,N_7406,N_5050);
or U9458 (N_9458,N_5076,N_6179);
or U9459 (N_9459,N_7397,N_6259);
nor U9460 (N_9460,N_7075,N_5149);
nand U9461 (N_9461,N_5326,N_6356);
nand U9462 (N_9462,N_7214,N_6415);
nor U9463 (N_9463,N_5723,N_6495);
nand U9464 (N_9464,N_6295,N_5194);
nand U9465 (N_9465,N_6703,N_6869);
nor U9466 (N_9466,N_6950,N_5616);
nor U9467 (N_9467,N_6380,N_7493);
and U9468 (N_9468,N_6287,N_7188);
nor U9469 (N_9469,N_5548,N_7105);
and U9470 (N_9470,N_7281,N_6696);
nand U9471 (N_9471,N_5455,N_6508);
and U9472 (N_9472,N_6068,N_6931);
and U9473 (N_9473,N_5297,N_6715);
nor U9474 (N_9474,N_7111,N_6357);
or U9475 (N_9475,N_5561,N_7414);
nand U9476 (N_9476,N_5477,N_7086);
nor U9477 (N_9477,N_6648,N_6533);
and U9478 (N_9478,N_5708,N_5626);
or U9479 (N_9479,N_6683,N_7166);
or U9480 (N_9480,N_6497,N_5807);
and U9481 (N_9481,N_6071,N_5423);
or U9482 (N_9482,N_5254,N_6165);
or U9483 (N_9483,N_5040,N_5931);
or U9484 (N_9484,N_5777,N_7046);
and U9485 (N_9485,N_5936,N_6949);
nand U9486 (N_9486,N_5408,N_5597);
nor U9487 (N_9487,N_7498,N_6005);
and U9488 (N_9488,N_5913,N_5995);
nand U9489 (N_9489,N_5364,N_5607);
and U9490 (N_9490,N_5446,N_6885);
nand U9491 (N_9491,N_6309,N_6081);
nor U9492 (N_9492,N_5470,N_7178);
nor U9493 (N_9493,N_6270,N_5014);
or U9494 (N_9494,N_5880,N_5846);
nand U9495 (N_9495,N_6955,N_5940);
nand U9496 (N_9496,N_6659,N_7391);
nand U9497 (N_9497,N_5434,N_5709);
nor U9498 (N_9498,N_5370,N_6344);
nor U9499 (N_9499,N_5050,N_6889);
nor U9500 (N_9500,N_6053,N_7257);
and U9501 (N_9501,N_5734,N_6525);
and U9502 (N_9502,N_6612,N_6717);
nor U9503 (N_9503,N_6508,N_7016);
and U9504 (N_9504,N_5316,N_5569);
nor U9505 (N_9505,N_5249,N_7197);
and U9506 (N_9506,N_7210,N_5910);
and U9507 (N_9507,N_5876,N_7473);
nand U9508 (N_9508,N_7326,N_5653);
and U9509 (N_9509,N_7169,N_6244);
or U9510 (N_9510,N_5062,N_7035);
and U9511 (N_9511,N_5850,N_5392);
and U9512 (N_9512,N_5799,N_6801);
nor U9513 (N_9513,N_6024,N_5431);
xnor U9514 (N_9514,N_5007,N_5995);
or U9515 (N_9515,N_5324,N_7052);
and U9516 (N_9516,N_5185,N_5691);
and U9517 (N_9517,N_7452,N_6550);
xor U9518 (N_9518,N_5585,N_6883);
or U9519 (N_9519,N_5389,N_6213);
nor U9520 (N_9520,N_7225,N_6469);
or U9521 (N_9521,N_5730,N_5081);
nand U9522 (N_9522,N_6313,N_6716);
nor U9523 (N_9523,N_7263,N_6210);
or U9524 (N_9524,N_6006,N_5886);
or U9525 (N_9525,N_7353,N_6740);
nor U9526 (N_9526,N_5285,N_6811);
nor U9527 (N_9527,N_5201,N_7073);
or U9528 (N_9528,N_6352,N_5261);
or U9529 (N_9529,N_5651,N_6171);
or U9530 (N_9530,N_6400,N_5850);
and U9531 (N_9531,N_5296,N_6756);
and U9532 (N_9532,N_5516,N_7176);
nand U9533 (N_9533,N_5177,N_5698);
nor U9534 (N_9534,N_6901,N_6724);
or U9535 (N_9535,N_5569,N_5468);
nand U9536 (N_9536,N_6690,N_5200);
nand U9537 (N_9537,N_5580,N_5780);
nand U9538 (N_9538,N_5963,N_6841);
and U9539 (N_9539,N_5703,N_7109);
and U9540 (N_9540,N_5707,N_6834);
or U9541 (N_9541,N_5640,N_7317);
nor U9542 (N_9542,N_5954,N_6628);
or U9543 (N_9543,N_7143,N_7429);
or U9544 (N_9544,N_5105,N_7102);
or U9545 (N_9545,N_5461,N_6963);
xnor U9546 (N_9546,N_5623,N_6274);
nand U9547 (N_9547,N_5547,N_6414);
nand U9548 (N_9548,N_6314,N_6582);
and U9549 (N_9549,N_6125,N_5214);
nor U9550 (N_9550,N_6536,N_5325);
or U9551 (N_9551,N_5258,N_5638);
nor U9552 (N_9552,N_5939,N_5319);
nand U9553 (N_9553,N_6605,N_7235);
or U9554 (N_9554,N_6519,N_7177);
or U9555 (N_9555,N_5623,N_6911);
nand U9556 (N_9556,N_7074,N_5226);
or U9557 (N_9557,N_5450,N_5949);
or U9558 (N_9558,N_6319,N_6131);
and U9559 (N_9559,N_6718,N_5952);
or U9560 (N_9560,N_6578,N_6550);
or U9561 (N_9561,N_6257,N_6807);
and U9562 (N_9562,N_7376,N_5728);
and U9563 (N_9563,N_7446,N_5198);
nand U9564 (N_9564,N_5515,N_7153);
nand U9565 (N_9565,N_6607,N_6012);
and U9566 (N_9566,N_6353,N_5894);
nor U9567 (N_9567,N_6226,N_6202);
xnor U9568 (N_9568,N_6937,N_6721);
nor U9569 (N_9569,N_5466,N_6354);
nand U9570 (N_9570,N_6940,N_6321);
nand U9571 (N_9571,N_7169,N_6569);
or U9572 (N_9572,N_5129,N_6018);
or U9573 (N_9573,N_5335,N_6131);
or U9574 (N_9574,N_5324,N_7377);
and U9575 (N_9575,N_6176,N_6823);
and U9576 (N_9576,N_7268,N_6200);
nand U9577 (N_9577,N_7058,N_5058);
or U9578 (N_9578,N_7104,N_6121);
and U9579 (N_9579,N_6757,N_5150);
nor U9580 (N_9580,N_5590,N_5305);
nor U9581 (N_9581,N_6680,N_6264);
or U9582 (N_9582,N_7077,N_6181);
nor U9583 (N_9583,N_5495,N_5822);
nor U9584 (N_9584,N_5835,N_6282);
and U9585 (N_9585,N_6399,N_6856);
or U9586 (N_9586,N_5964,N_7372);
and U9587 (N_9587,N_5543,N_6970);
nor U9588 (N_9588,N_6843,N_6831);
nand U9589 (N_9589,N_6542,N_6725);
and U9590 (N_9590,N_7068,N_7232);
nand U9591 (N_9591,N_7419,N_5847);
nor U9592 (N_9592,N_5017,N_6152);
or U9593 (N_9593,N_7110,N_7231);
nand U9594 (N_9594,N_6456,N_7019);
nor U9595 (N_9595,N_7001,N_5778);
and U9596 (N_9596,N_6459,N_5092);
nor U9597 (N_9597,N_5794,N_5232);
nor U9598 (N_9598,N_5849,N_6457);
nor U9599 (N_9599,N_7025,N_5351);
and U9600 (N_9600,N_7312,N_7315);
nor U9601 (N_9601,N_7141,N_5835);
and U9602 (N_9602,N_6848,N_7251);
or U9603 (N_9603,N_6066,N_6058);
and U9604 (N_9604,N_6367,N_7131);
and U9605 (N_9605,N_5599,N_5359);
nor U9606 (N_9606,N_6662,N_6830);
nor U9607 (N_9607,N_7477,N_5572);
and U9608 (N_9608,N_6784,N_5847);
nand U9609 (N_9609,N_7215,N_7285);
nand U9610 (N_9610,N_6151,N_6587);
and U9611 (N_9611,N_6710,N_5102);
nor U9612 (N_9612,N_6836,N_7435);
or U9613 (N_9613,N_6084,N_6423);
nor U9614 (N_9614,N_5816,N_6121);
and U9615 (N_9615,N_7122,N_6749);
nor U9616 (N_9616,N_5255,N_6554);
nand U9617 (N_9617,N_5916,N_6529);
and U9618 (N_9618,N_7165,N_6644);
nor U9619 (N_9619,N_5340,N_7122);
or U9620 (N_9620,N_5556,N_6155);
nand U9621 (N_9621,N_6859,N_5015);
and U9622 (N_9622,N_6333,N_6326);
nor U9623 (N_9623,N_5721,N_6729);
nand U9624 (N_9624,N_5878,N_6865);
or U9625 (N_9625,N_5547,N_7189);
and U9626 (N_9626,N_6828,N_5875);
or U9627 (N_9627,N_5202,N_5129);
or U9628 (N_9628,N_5542,N_5223);
nor U9629 (N_9629,N_6276,N_6030);
and U9630 (N_9630,N_7174,N_6897);
nand U9631 (N_9631,N_6837,N_5063);
nor U9632 (N_9632,N_5419,N_6378);
nor U9633 (N_9633,N_6710,N_6685);
nor U9634 (N_9634,N_6936,N_6076);
nand U9635 (N_9635,N_5743,N_7185);
or U9636 (N_9636,N_6007,N_5150);
nor U9637 (N_9637,N_5027,N_5152);
nor U9638 (N_9638,N_5610,N_6226);
nand U9639 (N_9639,N_6813,N_5717);
and U9640 (N_9640,N_6064,N_7226);
nand U9641 (N_9641,N_5863,N_5657);
nor U9642 (N_9642,N_7212,N_6256);
or U9643 (N_9643,N_6826,N_5892);
nand U9644 (N_9644,N_5315,N_7253);
and U9645 (N_9645,N_5694,N_6912);
or U9646 (N_9646,N_5217,N_5306);
nor U9647 (N_9647,N_7105,N_6555);
nand U9648 (N_9648,N_5753,N_5400);
or U9649 (N_9649,N_6609,N_5858);
nand U9650 (N_9650,N_6092,N_7345);
or U9651 (N_9651,N_5551,N_5206);
nor U9652 (N_9652,N_7346,N_6774);
or U9653 (N_9653,N_6063,N_5308);
nor U9654 (N_9654,N_5220,N_5351);
or U9655 (N_9655,N_5348,N_6824);
or U9656 (N_9656,N_6832,N_6730);
nand U9657 (N_9657,N_6154,N_6671);
nor U9658 (N_9658,N_6505,N_6971);
nor U9659 (N_9659,N_5728,N_6346);
nand U9660 (N_9660,N_7152,N_6063);
nand U9661 (N_9661,N_6933,N_5624);
nand U9662 (N_9662,N_5201,N_7362);
nand U9663 (N_9663,N_6809,N_6222);
nor U9664 (N_9664,N_5857,N_6965);
nand U9665 (N_9665,N_5308,N_6471);
nand U9666 (N_9666,N_5771,N_5849);
nand U9667 (N_9667,N_5914,N_5084);
xor U9668 (N_9668,N_7487,N_6874);
and U9669 (N_9669,N_6987,N_5106);
nor U9670 (N_9670,N_7457,N_5334);
and U9671 (N_9671,N_6521,N_5571);
or U9672 (N_9672,N_5173,N_6429);
and U9673 (N_9673,N_5091,N_5804);
nand U9674 (N_9674,N_5204,N_6225);
nor U9675 (N_9675,N_5255,N_5072);
xnor U9676 (N_9676,N_5675,N_6232);
and U9677 (N_9677,N_5277,N_6023);
nor U9678 (N_9678,N_6885,N_6041);
nand U9679 (N_9679,N_6476,N_6365);
nand U9680 (N_9680,N_7136,N_6155);
nor U9681 (N_9681,N_5833,N_5111);
or U9682 (N_9682,N_5341,N_7220);
nor U9683 (N_9683,N_6723,N_7256);
nor U9684 (N_9684,N_6232,N_5601);
nand U9685 (N_9685,N_6641,N_7027);
and U9686 (N_9686,N_7184,N_6709);
and U9687 (N_9687,N_6304,N_5016);
nand U9688 (N_9688,N_6122,N_5505);
and U9689 (N_9689,N_5712,N_6291);
or U9690 (N_9690,N_5104,N_5094);
or U9691 (N_9691,N_7494,N_5360);
nor U9692 (N_9692,N_7369,N_6979);
nand U9693 (N_9693,N_6555,N_6009);
and U9694 (N_9694,N_7153,N_6759);
and U9695 (N_9695,N_6305,N_5210);
nor U9696 (N_9696,N_7190,N_5467);
nor U9697 (N_9697,N_5637,N_5800);
nand U9698 (N_9698,N_6573,N_5284);
nor U9699 (N_9699,N_5268,N_5278);
and U9700 (N_9700,N_6432,N_5236);
nand U9701 (N_9701,N_6812,N_6356);
nor U9702 (N_9702,N_6117,N_6121);
or U9703 (N_9703,N_7116,N_6775);
or U9704 (N_9704,N_6717,N_6247);
or U9705 (N_9705,N_6328,N_7402);
or U9706 (N_9706,N_5315,N_6742);
nand U9707 (N_9707,N_5312,N_5097);
nor U9708 (N_9708,N_6130,N_5511);
and U9709 (N_9709,N_6962,N_5304);
nor U9710 (N_9710,N_6104,N_6678);
or U9711 (N_9711,N_5161,N_7340);
nand U9712 (N_9712,N_5058,N_5372);
nand U9713 (N_9713,N_6179,N_6608);
nand U9714 (N_9714,N_5746,N_6073);
nor U9715 (N_9715,N_5502,N_5962);
nand U9716 (N_9716,N_5227,N_7397);
nor U9717 (N_9717,N_6539,N_7057);
or U9718 (N_9718,N_6481,N_5877);
and U9719 (N_9719,N_5192,N_5895);
or U9720 (N_9720,N_6548,N_5469);
nor U9721 (N_9721,N_7495,N_5918);
nand U9722 (N_9722,N_6743,N_5335);
nand U9723 (N_9723,N_5743,N_5093);
nand U9724 (N_9724,N_5030,N_5610);
nor U9725 (N_9725,N_7455,N_5787);
and U9726 (N_9726,N_6584,N_5718);
and U9727 (N_9727,N_6038,N_6893);
or U9728 (N_9728,N_5766,N_7204);
and U9729 (N_9729,N_6302,N_6488);
and U9730 (N_9730,N_6573,N_5410);
nor U9731 (N_9731,N_5628,N_6696);
and U9732 (N_9732,N_5133,N_5870);
nor U9733 (N_9733,N_5702,N_6017);
and U9734 (N_9734,N_7076,N_7020);
nor U9735 (N_9735,N_6206,N_6777);
nand U9736 (N_9736,N_7142,N_5253);
or U9737 (N_9737,N_6535,N_5395);
or U9738 (N_9738,N_6642,N_6716);
nand U9739 (N_9739,N_7439,N_5949);
nor U9740 (N_9740,N_5537,N_6435);
or U9741 (N_9741,N_5356,N_7051);
nor U9742 (N_9742,N_5460,N_6305);
or U9743 (N_9743,N_5431,N_5327);
nand U9744 (N_9744,N_6420,N_6391);
or U9745 (N_9745,N_6904,N_7016);
or U9746 (N_9746,N_5765,N_6054);
or U9747 (N_9747,N_5172,N_7407);
nand U9748 (N_9748,N_7131,N_5438);
nor U9749 (N_9749,N_5256,N_6094);
or U9750 (N_9750,N_6147,N_6438);
and U9751 (N_9751,N_7187,N_5631);
nor U9752 (N_9752,N_5241,N_6359);
and U9753 (N_9753,N_5527,N_5966);
nor U9754 (N_9754,N_6019,N_6319);
or U9755 (N_9755,N_6116,N_5945);
nor U9756 (N_9756,N_7068,N_5403);
and U9757 (N_9757,N_5602,N_5220);
nor U9758 (N_9758,N_6676,N_5084);
nand U9759 (N_9759,N_5542,N_5682);
nand U9760 (N_9760,N_5529,N_6304);
nor U9761 (N_9761,N_5937,N_7265);
nor U9762 (N_9762,N_6772,N_5167);
and U9763 (N_9763,N_5106,N_6728);
or U9764 (N_9764,N_7401,N_6239);
and U9765 (N_9765,N_7153,N_5929);
nand U9766 (N_9766,N_6189,N_6506);
and U9767 (N_9767,N_6972,N_5097);
nor U9768 (N_9768,N_7273,N_6680);
nand U9769 (N_9769,N_6167,N_6217);
and U9770 (N_9770,N_7394,N_5473);
xor U9771 (N_9771,N_6788,N_6200);
nor U9772 (N_9772,N_6235,N_6687);
or U9773 (N_9773,N_6039,N_6015);
nand U9774 (N_9774,N_6452,N_5489);
or U9775 (N_9775,N_6570,N_6931);
and U9776 (N_9776,N_6875,N_7199);
and U9777 (N_9777,N_5207,N_6729);
and U9778 (N_9778,N_5232,N_6532);
and U9779 (N_9779,N_6040,N_6212);
and U9780 (N_9780,N_6115,N_5139);
nand U9781 (N_9781,N_6196,N_6241);
or U9782 (N_9782,N_5086,N_7054);
nor U9783 (N_9783,N_7244,N_6491);
or U9784 (N_9784,N_5694,N_5449);
nor U9785 (N_9785,N_6683,N_6565);
nand U9786 (N_9786,N_5727,N_6065);
nor U9787 (N_9787,N_5002,N_5077);
nand U9788 (N_9788,N_5245,N_6008);
nor U9789 (N_9789,N_5124,N_6898);
or U9790 (N_9790,N_6943,N_7179);
nand U9791 (N_9791,N_5930,N_6487);
nand U9792 (N_9792,N_6548,N_6442);
nor U9793 (N_9793,N_6807,N_5733);
or U9794 (N_9794,N_6777,N_7214);
nand U9795 (N_9795,N_6044,N_5154);
nor U9796 (N_9796,N_6426,N_5974);
and U9797 (N_9797,N_6427,N_6211);
and U9798 (N_9798,N_6545,N_6933);
or U9799 (N_9799,N_5272,N_6051);
nand U9800 (N_9800,N_6313,N_5017);
and U9801 (N_9801,N_6053,N_5548);
nor U9802 (N_9802,N_6724,N_6183);
or U9803 (N_9803,N_5066,N_7473);
nor U9804 (N_9804,N_6584,N_5807);
or U9805 (N_9805,N_5461,N_5055);
nor U9806 (N_9806,N_5854,N_5902);
and U9807 (N_9807,N_6893,N_7117);
nand U9808 (N_9808,N_5243,N_7144);
nor U9809 (N_9809,N_7196,N_7359);
nor U9810 (N_9810,N_5918,N_5040);
nor U9811 (N_9811,N_5339,N_5450);
nor U9812 (N_9812,N_6386,N_6735);
nand U9813 (N_9813,N_5474,N_7253);
nor U9814 (N_9814,N_6769,N_7129);
or U9815 (N_9815,N_6732,N_5400);
nand U9816 (N_9816,N_5384,N_5389);
nand U9817 (N_9817,N_6520,N_7276);
and U9818 (N_9818,N_7284,N_5829);
nand U9819 (N_9819,N_5247,N_5868);
nor U9820 (N_9820,N_6057,N_6843);
and U9821 (N_9821,N_5932,N_6699);
nor U9822 (N_9822,N_5656,N_6866);
and U9823 (N_9823,N_5897,N_6153);
and U9824 (N_9824,N_6600,N_6441);
or U9825 (N_9825,N_5502,N_6222);
nor U9826 (N_9826,N_6833,N_6677);
or U9827 (N_9827,N_6174,N_5084);
nand U9828 (N_9828,N_5074,N_6345);
or U9829 (N_9829,N_5691,N_5416);
or U9830 (N_9830,N_5307,N_5750);
nand U9831 (N_9831,N_5671,N_7114);
nor U9832 (N_9832,N_5262,N_6529);
nor U9833 (N_9833,N_6514,N_6308);
or U9834 (N_9834,N_6658,N_5405);
or U9835 (N_9835,N_7068,N_5195);
nand U9836 (N_9836,N_6962,N_5543);
and U9837 (N_9837,N_7215,N_6420);
or U9838 (N_9838,N_6075,N_6044);
nor U9839 (N_9839,N_5038,N_5261);
xor U9840 (N_9840,N_6634,N_5766);
nor U9841 (N_9841,N_6528,N_5594);
nand U9842 (N_9842,N_5130,N_6099);
and U9843 (N_9843,N_7191,N_6821);
nand U9844 (N_9844,N_7096,N_6327);
or U9845 (N_9845,N_5474,N_5771);
or U9846 (N_9846,N_7022,N_6622);
nor U9847 (N_9847,N_5986,N_5645);
and U9848 (N_9848,N_5119,N_5032);
and U9849 (N_9849,N_6824,N_6527);
nor U9850 (N_9850,N_5144,N_6801);
or U9851 (N_9851,N_7121,N_6040);
nand U9852 (N_9852,N_6717,N_7027);
nand U9853 (N_9853,N_6541,N_5155);
nor U9854 (N_9854,N_6313,N_6444);
nand U9855 (N_9855,N_6174,N_5771);
nand U9856 (N_9856,N_5766,N_5303);
and U9857 (N_9857,N_7319,N_5842);
and U9858 (N_9858,N_7182,N_5610);
nand U9859 (N_9859,N_5633,N_6120);
and U9860 (N_9860,N_7054,N_6558);
nor U9861 (N_9861,N_5366,N_5515);
xor U9862 (N_9862,N_6172,N_7238);
nand U9863 (N_9863,N_5203,N_5225);
nor U9864 (N_9864,N_5531,N_5044);
or U9865 (N_9865,N_5700,N_6981);
nand U9866 (N_9866,N_6731,N_6145);
nor U9867 (N_9867,N_5986,N_6453);
or U9868 (N_9868,N_6215,N_6056);
nor U9869 (N_9869,N_6334,N_6588);
and U9870 (N_9870,N_6842,N_6636);
nor U9871 (N_9871,N_5772,N_6280);
or U9872 (N_9872,N_5029,N_6294);
nand U9873 (N_9873,N_7407,N_7446);
or U9874 (N_9874,N_5378,N_6827);
and U9875 (N_9875,N_6143,N_7198);
nand U9876 (N_9876,N_6498,N_5404);
nor U9877 (N_9877,N_6139,N_6395);
or U9878 (N_9878,N_6657,N_6138);
nand U9879 (N_9879,N_6618,N_7169);
nand U9880 (N_9880,N_6166,N_6428);
xor U9881 (N_9881,N_6157,N_5323);
xnor U9882 (N_9882,N_6693,N_6896);
nor U9883 (N_9883,N_5685,N_5468);
xor U9884 (N_9884,N_6067,N_5131);
nor U9885 (N_9885,N_6774,N_5268);
or U9886 (N_9886,N_6553,N_5440);
nor U9887 (N_9887,N_5990,N_6804);
nand U9888 (N_9888,N_6018,N_6922);
nand U9889 (N_9889,N_7097,N_7180);
nand U9890 (N_9890,N_5413,N_5824);
or U9891 (N_9891,N_7312,N_5032);
nand U9892 (N_9892,N_5634,N_7374);
and U9893 (N_9893,N_7143,N_6843);
nor U9894 (N_9894,N_5906,N_5547);
nor U9895 (N_9895,N_5920,N_5828);
nand U9896 (N_9896,N_5733,N_6646);
and U9897 (N_9897,N_6821,N_6269);
and U9898 (N_9898,N_7106,N_5925);
or U9899 (N_9899,N_5179,N_6669);
or U9900 (N_9900,N_5821,N_6179);
and U9901 (N_9901,N_5997,N_5897);
nor U9902 (N_9902,N_7486,N_6877);
nand U9903 (N_9903,N_6797,N_6962);
or U9904 (N_9904,N_7245,N_6184);
nor U9905 (N_9905,N_7485,N_6363);
or U9906 (N_9906,N_6648,N_7401);
or U9907 (N_9907,N_6398,N_5091);
and U9908 (N_9908,N_5534,N_6944);
nand U9909 (N_9909,N_6996,N_5249);
or U9910 (N_9910,N_6072,N_7034);
nand U9911 (N_9911,N_5553,N_6078);
and U9912 (N_9912,N_5076,N_6185);
xor U9913 (N_9913,N_5092,N_6907);
or U9914 (N_9914,N_6345,N_5767);
nor U9915 (N_9915,N_5692,N_6173);
and U9916 (N_9916,N_7413,N_7314);
nand U9917 (N_9917,N_5640,N_6391);
or U9918 (N_9918,N_5805,N_6208);
nand U9919 (N_9919,N_7448,N_5371);
nor U9920 (N_9920,N_7354,N_5786);
xnor U9921 (N_9921,N_5400,N_5322);
and U9922 (N_9922,N_6428,N_6690);
or U9923 (N_9923,N_5446,N_5052);
or U9924 (N_9924,N_6408,N_7146);
or U9925 (N_9925,N_7368,N_7261);
or U9926 (N_9926,N_6730,N_5263);
nor U9927 (N_9927,N_6500,N_7313);
nand U9928 (N_9928,N_5506,N_5271);
nor U9929 (N_9929,N_5010,N_7135);
nor U9930 (N_9930,N_5828,N_5947);
and U9931 (N_9931,N_7112,N_7046);
nor U9932 (N_9932,N_5880,N_6079);
and U9933 (N_9933,N_6981,N_6099);
and U9934 (N_9934,N_6670,N_5921);
nor U9935 (N_9935,N_5420,N_5044);
and U9936 (N_9936,N_7421,N_5949);
nor U9937 (N_9937,N_6692,N_6935);
and U9938 (N_9938,N_6277,N_6219);
or U9939 (N_9939,N_7102,N_7175);
or U9940 (N_9940,N_6070,N_5690);
and U9941 (N_9941,N_5320,N_7060);
nand U9942 (N_9942,N_7348,N_5517);
and U9943 (N_9943,N_6205,N_6731);
nor U9944 (N_9944,N_5956,N_6930);
or U9945 (N_9945,N_5122,N_5569);
and U9946 (N_9946,N_5988,N_5671);
and U9947 (N_9947,N_5626,N_7435);
nand U9948 (N_9948,N_6768,N_6812);
nand U9949 (N_9949,N_5262,N_5525);
or U9950 (N_9950,N_5464,N_5630);
or U9951 (N_9951,N_7194,N_5094);
or U9952 (N_9952,N_5729,N_6476);
nand U9953 (N_9953,N_5511,N_5649);
nand U9954 (N_9954,N_6071,N_6443);
or U9955 (N_9955,N_7498,N_5453);
nor U9956 (N_9956,N_7437,N_6529);
and U9957 (N_9957,N_6828,N_6525);
nand U9958 (N_9958,N_5257,N_6060);
nand U9959 (N_9959,N_6204,N_6568);
or U9960 (N_9960,N_5732,N_5614);
nand U9961 (N_9961,N_5684,N_5571);
or U9962 (N_9962,N_5846,N_6074);
nor U9963 (N_9963,N_5200,N_7176);
or U9964 (N_9964,N_7215,N_5176);
nor U9965 (N_9965,N_6764,N_5905);
or U9966 (N_9966,N_6216,N_6671);
or U9967 (N_9967,N_5607,N_6871);
and U9968 (N_9968,N_5509,N_5918);
nor U9969 (N_9969,N_5348,N_5493);
nor U9970 (N_9970,N_6641,N_5616);
and U9971 (N_9971,N_6366,N_6651);
nand U9972 (N_9972,N_5118,N_6747);
and U9973 (N_9973,N_6577,N_5551);
xor U9974 (N_9974,N_7074,N_5327);
nand U9975 (N_9975,N_5901,N_7468);
and U9976 (N_9976,N_5537,N_5600);
nor U9977 (N_9977,N_5926,N_7227);
nand U9978 (N_9978,N_6474,N_6939);
nor U9979 (N_9979,N_6755,N_6390);
nor U9980 (N_9980,N_6658,N_5622);
nor U9981 (N_9981,N_5064,N_6721);
or U9982 (N_9982,N_6878,N_5287);
nand U9983 (N_9983,N_5086,N_7315);
or U9984 (N_9984,N_7493,N_5499);
nand U9985 (N_9985,N_6328,N_5003);
or U9986 (N_9986,N_5929,N_6901);
nand U9987 (N_9987,N_5810,N_6039);
nand U9988 (N_9988,N_5677,N_5292);
nor U9989 (N_9989,N_6253,N_6386);
nand U9990 (N_9990,N_5595,N_6584);
or U9991 (N_9991,N_6339,N_7431);
nand U9992 (N_9992,N_5186,N_6591);
and U9993 (N_9993,N_7372,N_6384);
nor U9994 (N_9994,N_6152,N_5872);
nand U9995 (N_9995,N_5030,N_5272);
or U9996 (N_9996,N_6499,N_5453);
nand U9997 (N_9997,N_5865,N_6983);
nor U9998 (N_9998,N_6610,N_5693);
nor U9999 (N_9999,N_5778,N_7485);
nand UO_0 (O_0,N_9602,N_8929);
nand UO_1 (O_1,N_8781,N_7508);
nor UO_2 (O_2,N_9142,N_7901);
and UO_3 (O_3,N_7516,N_9014);
nor UO_4 (O_4,N_7689,N_7861);
nor UO_5 (O_5,N_8985,N_9271);
or UO_6 (O_6,N_8420,N_9692);
nand UO_7 (O_7,N_8477,N_9789);
nand UO_8 (O_8,N_8837,N_9410);
nor UO_9 (O_9,N_7620,N_9729);
nand UO_10 (O_10,N_9574,N_7852);
nand UO_11 (O_11,N_8805,N_8979);
or UO_12 (O_12,N_9198,N_9021);
nor UO_13 (O_13,N_9000,N_8458);
nor UO_14 (O_14,N_9714,N_7552);
nor UO_15 (O_15,N_9205,N_8573);
nand UO_16 (O_16,N_8005,N_9066);
or UO_17 (O_17,N_7695,N_9258);
nand UO_18 (O_18,N_7616,N_8958);
or UO_19 (O_19,N_9759,N_9826);
nor UO_20 (O_20,N_9735,N_7835);
nor UO_21 (O_21,N_9501,N_7906);
nor UO_22 (O_22,N_9380,N_9564);
nor UO_23 (O_23,N_7859,N_9229);
nor UO_24 (O_24,N_8390,N_8565);
nor UO_25 (O_25,N_8762,N_8697);
nor UO_26 (O_26,N_8728,N_8620);
nor UO_27 (O_27,N_9458,N_8130);
nor UO_28 (O_28,N_9805,N_9466);
nand UO_29 (O_29,N_8609,N_8400);
nand UO_30 (O_30,N_9660,N_9561);
or UO_31 (O_31,N_8914,N_7992);
or UO_32 (O_32,N_8944,N_9024);
nand UO_33 (O_33,N_7868,N_8124);
and UO_34 (O_34,N_8838,N_8969);
and UO_35 (O_35,N_8933,N_9304);
or UO_36 (O_36,N_9423,N_9983);
nand UO_37 (O_37,N_8167,N_8798);
and UO_38 (O_38,N_9935,N_9573);
and UO_39 (O_39,N_7925,N_7533);
nor UO_40 (O_40,N_9074,N_7717);
nand UO_41 (O_41,N_9740,N_8426);
or UO_42 (O_42,N_9494,N_8419);
and UO_43 (O_43,N_7606,N_8309);
nor UO_44 (O_44,N_9543,N_7826);
nand UO_45 (O_45,N_9912,N_8399);
and UO_46 (O_46,N_8909,N_9474);
and UO_47 (O_47,N_8118,N_9617);
and UO_48 (O_48,N_9623,N_7625);
and UO_49 (O_49,N_7989,N_9227);
nor UO_50 (O_50,N_9450,N_8389);
and UO_51 (O_51,N_9545,N_8441);
nand UO_52 (O_52,N_8513,N_9815);
or UO_53 (O_53,N_8651,N_7786);
nand UO_54 (O_54,N_8931,N_9788);
or UO_55 (O_55,N_8563,N_9876);
nor UO_56 (O_56,N_9678,N_8025);
nand UO_57 (O_57,N_9129,N_7823);
nor UO_58 (O_58,N_9092,N_8231);
nand UO_59 (O_59,N_8382,N_9875);
and UO_60 (O_60,N_9784,N_7542);
nand UO_61 (O_61,N_8219,N_7936);
nand UO_62 (O_62,N_8073,N_9381);
nor UO_63 (O_63,N_8726,N_8258);
nand UO_64 (O_64,N_8230,N_8248);
nor UO_65 (O_65,N_8644,N_7774);
nand UO_66 (O_66,N_7768,N_8751);
and UO_67 (O_67,N_9916,N_9975);
nand UO_68 (O_68,N_7685,N_8997);
and UO_69 (O_69,N_9974,N_9313);
and UO_70 (O_70,N_9048,N_7720);
nor UO_71 (O_71,N_9001,N_9799);
nor UO_72 (O_72,N_9103,N_9322);
nor UO_73 (O_73,N_8558,N_8430);
or UO_74 (O_74,N_8113,N_8431);
nor UO_75 (O_75,N_8013,N_8171);
or UO_76 (O_76,N_9084,N_9584);
nand UO_77 (O_77,N_8666,N_9080);
or UO_78 (O_78,N_9200,N_8050);
nand UO_79 (O_79,N_7547,N_8746);
nor UO_80 (O_80,N_8294,N_8061);
nor UO_81 (O_81,N_9090,N_8404);
nor UO_82 (O_82,N_8634,N_9987);
nor UO_83 (O_83,N_9982,N_8191);
nand UO_84 (O_84,N_9694,N_9592);
or UO_85 (O_85,N_8024,N_9931);
and UO_86 (O_86,N_7876,N_9881);
and UO_87 (O_87,N_8069,N_8597);
nand UO_88 (O_88,N_7645,N_8974);
and UO_89 (O_89,N_9721,N_9144);
nand UO_90 (O_90,N_8981,N_8353);
and UO_91 (O_91,N_7964,N_9559);
nand UO_92 (O_92,N_8650,N_8999);
nor UO_93 (O_93,N_7562,N_9862);
or UO_94 (O_94,N_8352,N_7808);
or UO_95 (O_95,N_7512,N_8938);
nand UO_96 (O_96,N_8589,N_8684);
nand UO_97 (O_97,N_8495,N_8953);
and UO_98 (O_98,N_7810,N_7754);
or UO_99 (O_99,N_8412,N_8383);
nand UO_100 (O_100,N_7621,N_7913);
nand UO_101 (O_101,N_9757,N_7990);
and UO_102 (O_102,N_9715,N_7760);
nor UO_103 (O_103,N_9940,N_9747);
and UO_104 (O_104,N_8827,N_9513);
nand UO_105 (O_105,N_8306,N_7982);
or UO_106 (O_106,N_9107,N_9923);
or UO_107 (O_107,N_9634,N_9842);
nor UO_108 (O_108,N_9036,N_8525);
nor UO_109 (O_109,N_7713,N_8063);
and UO_110 (O_110,N_8244,N_7587);
or UO_111 (O_111,N_8311,N_8302);
and UO_112 (O_112,N_9065,N_8755);
nor UO_113 (O_113,N_8160,N_9254);
or UO_114 (O_114,N_9956,N_8022);
and UO_115 (O_115,N_8575,N_9595);
nor UO_116 (O_116,N_8688,N_9582);
or UO_117 (O_117,N_9417,N_7657);
or UO_118 (O_118,N_9087,N_8801);
and UO_119 (O_119,N_8267,N_7986);
and UO_120 (O_120,N_7895,N_8872);
nand UO_121 (O_121,N_8682,N_8698);
xor UO_122 (O_122,N_8741,N_8304);
or UO_123 (O_123,N_8036,N_7812);
nand UO_124 (O_124,N_9492,N_8894);
or UO_125 (O_125,N_8208,N_7513);
nand UO_126 (O_126,N_8445,N_8657);
and UO_127 (O_127,N_9658,N_8438);
nand UO_128 (O_128,N_9894,N_8694);
nand UO_129 (O_129,N_8181,N_7752);
nand UO_130 (O_130,N_7984,N_9125);
or UO_131 (O_131,N_8328,N_9857);
and UO_132 (O_132,N_8917,N_8580);
nor UO_133 (O_133,N_8183,N_9625);
and UO_134 (O_134,N_7762,N_9057);
and UO_135 (O_135,N_9877,N_8767);
nor UO_136 (O_136,N_8713,N_7784);
nand UO_137 (O_137,N_9929,N_8531);
or UO_138 (O_138,N_8515,N_9638);
nand UO_139 (O_139,N_8176,N_8239);
and UO_140 (O_140,N_8615,N_9452);
nand UO_141 (O_141,N_9155,N_7523);
nand UO_142 (O_142,N_8284,N_8295);
and UO_143 (O_143,N_8840,N_7694);
or UO_144 (O_144,N_9343,N_9674);
nand UO_145 (O_145,N_8507,N_8481);
or UO_146 (O_146,N_7904,N_9756);
nor UO_147 (O_147,N_8749,N_9893);
xnor UO_148 (O_148,N_9713,N_8004);
or UO_149 (O_149,N_8133,N_8395);
or UO_150 (O_150,N_8165,N_8137);
nand UO_151 (O_151,N_9994,N_8845);
nor UO_152 (O_152,N_8280,N_9320);
nand UO_153 (O_153,N_8885,N_8355);
or UO_154 (O_154,N_8829,N_9578);
nor UO_155 (O_155,N_9774,N_9978);
nand UO_156 (O_156,N_9791,N_7806);
or UO_157 (O_157,N_8897,N_8460);
nand UO_158 (O_158,N_9299,N_8660);
nand UO_159 (O_159,N_8444,N_8970);
and UO_160 (O_160,N_8119,N_8928);
nand UO_161 (O_161,N_7544,N_9314);
nor UO_162 (O_162,N_8792,N_8593);
and UO_163 (O_163,N_7951,N_7961);
or UO_164 (O_164,N_9897,N_8008);
nand UO_165 (O_165,N_7738,N_7858);
nand UO_166 (O_166,N_8966,N_9079);
nand UO_167 (O_167,N_7800,N_9888);
nor UO_168 (O_168,N_9253,N_8936);
nor UO_169 (O_169,N_8910,N_7672);
nor UO_170 (O_170,N_7912,N_9848);
nand UO_171 (O_171,N_8027,N_7734);
or UO_172 (O_172,N_8057,N_8707);
nor UO_173 (O_173,N_8806,N_7642);
nor UO_174 (O_174,N_8003,N_8105);
nand UO_175 (O_175,N_8822,N_9828);
nand UO_176 (O_176,N_9618,N_9403);
nand UO_177 (O_177,N_7837,N_9977);
nor UO_178 (O_178,N_7952,N_9095);
nand UO_179 (O_179,N_8791,N_8376);
and UO_180 (O_180,N_9123,N_9162);
or UO_181 (O_181,N_9588,N_8907);
or UO_182 (O_182,N_9363,N_9599);
nand UO_183 (O_183,N_8312,N_9546);
nor UO_184 (O_184,N_8059,N_9062);
nor UO_185 (O_185,N_8566,N_8711);
nor UO_186 (O_186,N_8942,N_7704);
or UO_187 (O_187,N_9244,N_9432);
nor UO_188 (O_188,N_8347,N_7598);
or UO_189 (O_189,N_8537,N_8740);
nor UO_190 (O_190,N_8807,N_8529);
and UO_191 (O_191,N_9840,N_9701);
and UO_192 (O_192,N_9918,N_8014);
nand UO_193 (O_193,N_8182,N_7789);
nor UO_194 (O_194,N_8315,N_9484);
or UO_195 (O_195,N_7770,N_7920);
and UO_196 (O_196,N_8492,N_9909);
and UO_197 (O_197,N_7622,N_9708);
or UO_198 (O_198,N_8152,N_7945);
nand UO_199 (O_199,N_8672,N_9239);
nand UO_200 (O_200,N_8645,N_9454);
nor UO_201 (O_201,N_7898,N_7613);
or UO_202 (O_202,N_9814,N_8342);
nor UO_203 (O_203,N_9976,N_9053);
nand UO_204 (O_204,N_7847,N_9807);
xnor UO_205 (O_205,N_9248,N_9712);
or UO_206 (O_206,N_7502,N_7710);
nor UO_207 (O_207,N_8300,N_8247);
and UO_208 (O_208,N_9158,N_8766);
nand UO_209 (O_209,N_9136,N_7579);
and UO_210 (O_210,N_8368,N_9115);
or UO_211 (O_211,N_9269,N_9211);
or UO_212 (O_212,N_9521,N_9113);
nand UO_213 (O_213,N_8269,N_7865);
nor UO_214 (O_214,N_9216,N_9839);
nand UO_215 (O_215,N_9769,N_9058);
and UO_216 (O_216,N_9621,N_9568);
or UO_217 (O_217,N_8864,N_8560);
and UO_218 (O_218,N_9161,N_9420);
nor UO_219 (O_219,N_7853,N_7571);
or UO_220 (O_220,N_7905,N_8384);
nand UO_221 (O_221,N_8019,N_7791);
nand UO_222 (O_222,N_7742,N_8147);
nand UO_223 (O_223,N_8877,N_9972);
or UO_224 (O_224,N_7527,N_8718);
or UO_225 (O_225,N_9265,N_8144);
nor UO_226 (O_226,N_9147,N_9849);
nand UO_227 (O_227,N_8629,N_9159);
and UO_228 (O_228,N_7630,N_9991);
or UO_229 (O_229,N_8636,N_8453);
nor UO_230 (O_230,N_9139,N_8029);
and UO_231 (O_231,N_8341,N_9440);
nor UO_232 (O_232,N_8918,N_8317);
nand UO_233 (O_233,N_9288,N_9699);
and UO_234 (O_234,N_8948,N_9823);
nand UO_235 (O_235,N_8185,N_9919);
and UO_236 (O_236,N_8452,N_8545);
nand UO_237 (O_237,N_7666,N_9117);
or UO_238 (O_238,N_7997,N_9263);
nor UO_239 (O_239,N_9743,N_8223);
nor UO_240 (O_240,N_7707,N_7922);
or UO_241 (O_241,N_8818,N_9270);
nor UO_242 (O_242,N_8415,N_8879);
or UO_243 (O_243,N_9750,N_9981);
nand UO_244 (O_244,N_8401,N_7712);
nand UO_245 (O_245,N_7680,N_9698);
nand UO_246 (O_246,N_9030,N_7797);
nand UO_247 (O_247,N_8546,N_8861);
nor UO_248 (O_248,N_8346,N_9984);
nor UO_249 (O_249,N_9645,N_9586);
or UO_250 (O_250,N_7545,N_9127);
or UO_251 (O_251,N_9996,N_9368);
nand UO_252 (O_252,N_8583,N_7883);
nor UO_253 (O_253,N_8963,N_9950);
nor UO_254 (O_254,N_8703,N_9089);
nor UO_255 (O_255,N_8808,N_9910);
and UO_256 (O_256,N_8964,N_9635);
or UO_257 (O_257,N_7652,N_9643);
and UO_258 (O_258,N_7924,N_8476);
or UO_259 (O_259,N_7677,N_7850);
nand UO_260 (O_260,N_8709,N_8344);
and UO_261 (O_261,N_8141,N_8018);
or UO_262 (O_262,N_9177,N_9203);
and UO_263 (O_263,N_9844,N_7698);
or UO_264 (O_264,N_8474,N_8721);
and UO_265 (O_265,N_7785,N_9583);
nor UO_266 (O_266,N_8220,N_8539);
and UO_267 (O_267,N_9359,N_9422);
nor UO_268 (O_268,N_8202,N_7880);
nand UO_269 (O_269,N_8282,N_7661);
or UO_270 (O_270,N_8483,N_9971);
and UO_271 (O_271,N_9151,N_7519);
nor UO_272 (O_272,N_8784,N_9291);
or UO_273 (O_273,N_7687,N_9310);
nand UO_274 (O_274,N_8442,N_8117);
nand UO_275 (O_275,N_8002,N_7975);
nor UO_276 (O_276,N_8139,N_9306);
or UO_277 (O_277,N_9519,N_9356);
or UO_278 (O_278,N_8333,N_7801);
nand UO_279 (O_279,N_7960,N_7888);
nor UO_280 (O_280,N_9329,N_7716);
nor UO_281 (O_281,N_9206,N_8544);
nor UO_282 (O_282,N_8257,N_9668);
nor UO_283 (O_283,N_8530,N_8890);
nor UO_284 (O_284,N_9182,N_8735);
nor UO_285 (O_285,N_8725,N_8285);
xnor UO_286 (O_286,N_9471,N_8564);
nand UO_287 (O_287,N_9413,N_8490);
and UO_288 (O_288,N_9847,N_7809);
or UO_289 (O_289,N_9609,N_8641);
nand UO_290 (O_290,N_9215,N_8816);
nor UO_291 (O_291,N_8243,N_7553);
nand UO_292 (O_292,N_8648,N_8043);
and UO_293 (O_293,N_8339,N_9226);
nor UO_294 (O_294,N_9869,N_7885);
and UO_295 (O_295,N_8823,N_7841);
nand UO_296 (O_296,N_8760,N_9949);
nor UO_297 (O_297,N_7813,N_9149);
nand UO_298 (O_298,N_9187,N_8463);
nand UO_299 (O_299,N_9914,N_8060);
nor UO_300 (O_300,N_7766,N_8567);
and UO_301 (O_301,N_9832,N_9398);
and UO_302 (O_302,N_9015,N_9575);
or UO_303 (O_303,N_9082,N_9855);
nor UO_304 (O_304,N_9455,N_8790);
nor UO_305 (O_305,N_9020,N_8689);
nor UO_306 (O_306,N_7977,N_9746);
and UO_307 (O_307,N_7627,N_9331);
or UO_308 (O_308,N_9696,N_8475);
and UO_309 (O_309,N_7996,N_7667);
or UO_310 (O_310,N_8775,N_8407);
and UO_311 (O_311,N_9489,N_7804);
and UO_312 (O_312,N_8461,N_9662);
or UO_313 (O_313,N_8209,N_8148);
nand UO_314 (O_314,N_9346,N_8950);
or UO_315 (O_315,N_8858,N_9580);
nor UO_316 (O_316,N_7546,N_9164);
nor UO_317 (O_317,N_7958,N_7656);
nor UO_318 (O_318,N_9146,N_7724);
nand UO_319 (O_319,N_9407,N_8913);
nor UO_320 (O_320,N_8486,N_8600);
nand UO_321 (O_321,N_9402,N_8848);
nor UO_322 (O_322,N_8523,N_8482);
nor UO_323 (O_323,N_8548,N_9899);
or UO_324 (O_324,N_7634,N_9763);
nor UO_325 (O_325,N_9041,N_8192);
or UO_326 (O_326,N_8750,N_9262);
nand UO_327 (O_327,N_9672,N_9439);
nand UO_328 (O_328,N_9605,N_7658);
nor UO_329 (O_329,N_8321,N_9811);
nand UO_330 (O_330,N_8677,N_9386);
nand UO_331 (O_331,N_8883,N_8072);
and UO_332 (O_332,N_7615,N_9808);
nand UO_333 (O_333,N_7691,N_8131);
or UO_334 (O_334,N_8594,N_7524);
xnor UO_335 (O_335,N_9340,N_9004);
nor UO_336 (O_336,N_9510,N_8626);
and UO_337 (O_337,N_9833,N_7970);
nor UO_338 (O_338,N_8758,N_8142);
nand UO_339 (O_339,N_7769,N_9207);
and UO_340 (O_340,N_8180,N_8394);
or UO_341 (O_341,N_7974,N_9507);
or UO_342 (O_342,N_8947,N_8042);
nor UO_343 (O_343,N_9154,N_9552);
and UO_344 (O_344,N_7911,N_9184);
or UO_345 (O_345,N_9770,N_8241);
nor UO_346 (O_346,N_8602,N_8109);
and UO_347 (O_347,N_9677,N_9333);
nor UO_348 (O_348,N_7592,N_8251);
nand UO_349 (O_349,N_9094,N_8210);
nand UO_350 (O_350,N_8363,N_9795);
nand UO_351 (O_351,N_7739,N_9453);
or UO_352 (O_352,N_8068,N_8814);
nand UO_353 (O_353,N_7973,N_7910);
nor UO_354 (O_354,N_9539,N_8994);
and UO_355 (O_355,N_9490,N_9554);
nand UO_356 (O_356,N_9383,N_8417);
nand UO_357 (O_357,N_8880,N_9597);
nand UO_358 (O_358,N_7543,N_8071);
nor UO_359 (O_359,N_9027,N_9734);
and UO_360 (O_360,N_8608,N_7675);
or UO_361 (O_361,N_9682,N_8824);
or UO_362 (O_362,N_7683,N_9045);
nand UO_363 (O_363,N_7648,N_8528);
nand UO_364 (O_364,N_8542,N_7708);
and UO_365 (O_365,N_9050,N_8015);
or UO_366 (O_366,N_9236,N_8654);
nor UO_367 (O_367,N_8291,N_9273);
or UO_368 (O_368,N_9649,N_9813);
nand UO_369 (O_369,N_8611,N_9793);
nor UO_370 (O_370,N_9557,N_7651);
or UO_371 (O_371,N_8278,N_8038);
and UO_372 (O_372,N_9934,N_9470);
nand UO_373 (O_373,N_9879,N_9056);
and UO_374 (O_374,N_9111,N_8723);
nor UO_375 (O_375,N_8314,N_8279);
nand UO_376 (O_376,N_8356,N_9110);
or UO_377 (O_377,N_7521,N_9531);
and UO_378 (O_378,N_9797,N_8813);
nand UO_379 (O_379,N_7511,N_8017);
or UO_380 (O_380,N_8048,N_8421);
and UO_381 (O_381,N_7879,N_9292);
and UO_382 (O_382,N_7640,N_9819);
or UO_383 (O_383,N_8954,N_9278);
nor UO_384 (O_384,N_9366,N_7732);
nand UO_385 (O_385,N_9870,N_9208);
nor UO_386 (O_386,N_8955,N_8561);
nor UO_387 (O_387,N_7686,N_8518);
or UO_388 (O_388,N_7749,N_9655);
and UO_389 (O_389,N_7583,N_8896);
nand UO_390 (O_390,N_7890,N_8586);
or UO_391 (O_391,N_9705,N_9874);
nor UO_392 (O_392,N_8331,N_8932);
and UO_393 (O_393,N_7550,N_7854);
nor UO_394 (O_394,N_7978,N_9347);
or UO_395 (O_395,N_9619,N_9775);
and UO_396 (O_396,N_7551,N_9687);
nor UO_397 (O_397,N_9391,N_9749);
nor UO_398 (O_398,N_8836,N_7926);
and UO_399 (O_399,N_9863,N_9165);
and UO_400 (O_400,N_7946,N_9859);
and UO_401 (O_401,N_8206,N_8323);
nor UO_402 (O_402,N_8570,N_8381);
or UO_403 (O_403,N_8770,N_8372);
nor UO_404 (O_404,N_8850,N_7827);
nor UO_405 (O_405,N_9424,N_9629);
nor UO_406 (O_406,N_9852,N_8487);
nand UO_407 (O_407,N_9902,N_9491);
nand UO_408 (O_408,N_7845,N_9630);
nor UO_409 (O_409,N_9824,N_8099);
and UO_410 (O_410,N_8313,N_8056);
nor UO_411 (O_411,N_7862,N_8519);
or UO_412 (O_412,N_9081,N_9318);
nor UO_413 (O_413,N_8887,N_8177);
and UO_414 (O_414,N_9010,N_7582);
nor UO_415 (O_415,N_8949,N_8406);
and UO_416 (O_416,N_9483,N_8326);
or UO_417 (O_417,N_8360,N_8268);
and UO_418 (O_418,N_9632,N_9719);
or UO_419 (O_419,N_7690,N_7709);
and UO_420 (O_420,N_9078,N_9370);
nor UO_421 (O_421,N_7908,N_9684);
nand UO_422 (O_422,N_9153,N_7846);
or UO_423 (O_423,N_9109,N_8283);
nand UO_424 (O_424,N_8794,N_8643);
or UO_425 (O_425,N_8164,N_8842);
nand UO_426 (O_426,N_9913,N_8538);
nand UO_427 (O_427,N_9915,N_9404);
nand UO_428 (O_428,N_9190,N_9102);
nor UO_429 (O_429,N_9120,N_8473);
nor UO_430 (O_430,N_9480,N_7601);
nor UO_431 (O_431,N_7585,N_8987);
and UO_432 (O_432,N_8865,N_7594);
nor UO_433 (O_433,N_9556,N_8912);
nor UO_434 (O_434,N_8380,N_8856);
and UO_435 (O_435,N_8178,N_8493);
nor UO_436 (O_436,N_7733,N_9419);
nand UO_437 (O_437,N_9406,N_7864);
nor UO_438 (O_438,N_7765,N_9388);
nor UO_439 (O_439,N_8026,N_9108);
nor UO_440 (O_440,N_8195,N_8470);
nor UO_441 (O_441,N_7570,N_8977);
or UO_442 (O_442,N_8745,N_9528);
nand UO_443 (O_443,N_9943,N_7772);
nand UO_444 (O_444,N_8965,N_7962);
nor UO_445 (O_445,N_9512,N_7662);
nand UO_446 (O_446,N_8956,N_9055);
or UO_447 (O_447,N_9099,N_8354);
nor UO_448 (O_448,N_9937,N_9339);
or UO_449 (O_449,N_8370,N_8536);
and UO_450 (O_450,N_8578,N_9114);
nand UO_451 (O_451,N_9890,N_9251);
and UO_452 (O_452,N_7919,N_8797);
nor UO_453 (O_453,N_8982,N_8098);
or UO_454 (O_454,N_9724,N_8995);
or UO_455 (O_455,N_9738,N_9904);
or UO_456 (O_456,N_8778,N_7897);
nor UO_457 (O_457,N_7877,N_9830);
and UO_458 (O_458,N_7856,N_8574);
and UO_459 (O_459,N_8768,N_9733);
and UO_460 (O_460,N_8081,N_9921);
nor UO_461 (O_461,N_9603,N_9547);
nor UO_462 (O_462,N_9332,N_7987);
nand UO_463 (O_463,N_8386,N_9898);
nand UO_464 (O_464,N_9871,N_8882);
nor UO_465 (O_465,N_8957,N_8708);
and UO_466 (O_466,N_8437,N_9858);
or UO_467 (O_467,N_9042,N_7700);
nor UO_468 (O_468,N_7777,N_7900);
nand UO_469 (O_469,N_8093,N_8676);
nor UO_470 (O_470,N_9666,N_8450);
nor UO_471 (O_471,N_9119,N_8802);
nand UO_472 (O_472,N_8815,N_9193);
and UO_473 (O_473,N_7814,N_8174);
or UO_474 (O_474,N_8673,N_9969);
nand UO_475 (O_475,N_8738,N_8335);
nand UO_476 (O_476,N_9148,N_8753);
or UO_477 (O_477,N_7927,N_8101);
and UO_478 (O_478,N_9341,N_9903);
and UO_479 (O_479,N_8522,N_8028);
and UO_480 (O_480,N_8110,N_9375);
and UO_481 (O_481,N_9171,N_9298);
or UO_482 (O_482,N_7819,N_8127);
or UO_483 (O_483,N_8780,N_9163);
or UO_484 (O_484,N_9502,N_7820);
nand UO_485 (O_485,N_8526,N_8855);
and UO_486 (O_486,N_8397,N_8275);
nor UO_487 (O_487,N_8973,N_8710);
and UO_488 (O_488,N_8378,N_8705);
and UO_489 (O_489,N_9328,N_8270);
or UO_490 (O_490,N_7572,N_8034);
nand UO_491 (O_491,N_9970,N_8961);
nor UO_492 (O_492,N_7863,N_9019);
nand UO_493 (O_493,N_8759,N_9167);
or UO_494 (O_494,N_8464,N_8764);
nand UO_495 (O_495,N_8429,N_9604);
or UO_496 (O_496,N_7914,N_8862);
nor UO_497 (O_497,N_7949,N_9275);
or UO_498 (O_498,N_7848,N_9003);
nand UO_499 (O_499,N_9071,N_8067);
nand UO_500 (O_500,N_7560,N_7539);
and UO_501 (O_501,N_8901,N_9002);
or UO_502 (O_502,N_7860,N_9284);
and UO_503 (O_503,N_9191,N_9717);
or UO_504 (O_504,N_8681,N_9435);
nand UO_505 (O_505,N_7849,N_9059);
nor UO_506 (O_506,N_8075,N_9237);
or UO_507 (O_507,N_8761,N_8662);
or UO_508 (O_508,N_7855,N_7617);
nand UO_509 (O_509,N_8729,N_9965);
or UO_510 (O_510,N_9628,N_7663);
or UO_511 (O_511,N_9214,N_7679);
and UO_512 (O_512,N_9234,N_7923);
nand UO_513 (O_513,N_7916,N_9296);
nand UO_514 (O_514,N_8106,N_9720);
nand UO_515 (O_515,N_7501,N_7815);
and UO_516 (O_516,N_9992,N_8252);
nor UO_517 (O_517,N_8996,N_8720);
nand UO_518 (O_518,N_8184,N_9463);
or UO_519 (O_519,N_7573,N_9371);
or UO_520 (O_520,N_9880,N_9782);
and UO_521 (O_521,N_8904,N_9009);
or UO_522 (O_522,N_9106,N_9377);
nand UO_523 (O_523,N_8607,N_8627);
nand UO_524 (O_524,N_7816,N_9952);
nor UO_525 (O_525,N_9924,N_9865);
and UO_526 (O_526,N_9755,N_9412);
nand UO_527 (O_527,N_8250,N_9098);
nor UO_528 (O_528,N_9787,N_7824);
nor UO_529 (O_529,N_8699,N_9500);
or UO_530 (O_530,N_8074,N_9933);
and UO_531 (O_531,N_8039,N_9196);
nand UO_532 (O_532,N_7595,N_8221);
nor UO_533 (O_533,N_7518,N_9083);
nand UO_534 (O_534,N_7699,N_9192);
and UO_535 (O_535,N_7736,N_7534);
and UO_536 (O_536,N_8085,N_9442);
nor UO_537 (O_537,N_9567,N_9425);
or UO_538 (O_538,N_9854,N_7610);
nor UO_539 (O_539,N_8655,N_9954);
nor UO_540 (O_540,N_9895,N_7793);
or UO_541 (O_541,N_8844,N_8554);
nand UO_542 (O_542,N_7894,N_8783);
nand UO_543 (O_543,N_8937,N_8217);
or UO_544 (O_544,N_9864,N_8079);
nor UO_545 (O_545,N_8757,N_9882);
and UO_546 (O_546,N_8047,N_8795);
nor UO_547 (O_547,N_7755,N_9540);
nor UO_548 (O_548,N_8508,N_9688);
nor UO_549 (O_549,N_7576,N_9063);
and UO_550 (O_550,N_8799,N_8524);
and UO_551 (O_551,N_8527,N_8290);
or UO_552 (O_552,N_9961,N_9948);
nand UO_553 (O_553,N_7776,N_9637);
and UO_554 (O_554,N_9511,N_8610);
or UO_555 (O_555,N_8310,N_8906);
or UO_556 (O_556,N_8488,N_9464);
nand UO_557 (O_557,N_9307,N_8103);
or UO_558 (O_558,N_9695,N_7728);
and UO_559 (O_559,N_8197,N_8227);
or UO_560 (O_560,N_7991,N_9487);
and UO_561 (O_561,N_7889,N_9212);
and UO_562 (O_562,N_7702,N_9731);
or UO_563 (O_563,N_9277,N_9364);
nor UO_564 (O_564,N_9768,N_8203);
nor UO_565 (O_565,N_8035,N_8878);
or UO_566 (O_566,N_7743,N_9017);
nor UO_567 (O_567,N_7748,N_9741);
nor UO_568 (O_568,N_9224,N_8604);
nor UO_569 (O_569,N_9018,N_8196);
nand UO_570 (O_570,N_7998,N_7943);
and UO_571 (O_571,N_9772,N_8534);
xor UO_572 (O_572,N_8277,N_8467);
nor UO_573 (O_573,N_8375,N_8521);
or UO_574 (O_574,N_7753,N_9105);
or UO_575 (O_575,N_9256,N_9220);
nor UO_576 (O_576,N_8946,N_8193);
nand UO_577 (O_577,N_9989,N_9186);
or UO_578 (O_578,N_8114,N_8112);
nor UO_579 (O_579,N_9944,N_9527);
nand UO_580 (O_580,N_9892,N_8145);
or UO_581 (O_581,N_8585,N_8841);
nand UO_582 (O_582,N_7969,N_8338);
nand UO_583 (O_583,N_8693,N_8543);
nand UO_584 (O_584,N_7780,N_9508);
nor UO_585 (O_585,N_8789,N_9397);
and UO_586 (O_586,N_9379,N_7623);
xor UO_587 (O_587,N_8296,N_7872);
nor UO_588 (O_588,N_8998,N_9067);
or UO_589 (O_589,N_8871,N_8516);
nand UO_590 (O_590,N_8991,N_8308);
or UO_591 (O_591,N_9047,N_8410);
or UO_592 (O_592,N_7715,N_8064);
nand UO_593 (O_593,N_9646,N_9429);
nor UO_594 (O_594,N_9960,N_9469);
xor UO_595 (O_595,N_8359,N_9607);
or UO_596 (O_596,N_8943,N_8930);
nand UO_597 (O_597,N_8188,N_7740);
or UO_598 (O_598,N_8062,N_8867);
nor UO_599 (O_599,N_8993,N_8215);
and UO_600 (O_600,N_7684,N_7701);
nor UO_601 (O_601,N_8447,N_8642);
and UO_602 (O_602,N_8934,N_8053);
and UO_603 (O_603,N_8754,N_7574);
or UO_604 (O_604,N_9408,N_9744);
or UO_605 (O_605,N_9088,N_7798);
nand UO_606 (O_606,N_8502,N_8409);
and UO_607 (O_607,N_9670,N_7878);
nand UO_608 (O_608,N_7631,N_9798);
nand UO_609 (O_609,N_8161,N_8379);
and UO_610 (O_610,N_7597,N_8175);
nand UO_611 (O_611,N_7559,N_9267);
nor UO_612 (O_612,N_9112,N_8983);
or UO_613 (O_613,N_8212,N_9663);
or UO_614 (O_614,N_8076,N_9315);
nor UO_615 (O_615,N_9286,N_9199);
nand UO_616 (O_616,N_9572,N_9690);
nor UO_617 (O_617,N_7871,N_9765);
and UO_618 (O_618,N_7761,N_8860);
nand UO_619 (O_619,N_8023,N_9927);
and UO_620 (O_620,N_9321,N_8007);
nand UO_621 (O_621,N_8416,N_9443);
nor UO_622 (O_622,N_9594,N_8935);
or UO_623 (O_623,N_8424,N_9570);
nand UO_624 (O_624,N_8941,N_9069);
nor UO_625 (O_625,N_9963,N_7950);
nor UO_626 (O_626,N_8922,N_7703);
nand UO_627 (O_627,N_7535,N_8224);
and UO_628 (O_628,N_9185,N_8211);
and UO_629 (O_629,N_9495,N_8719);
nor UO_630 (O_630,N_7857,N_8786);
nand UO_631 (O_631,N_8653,N_8329);
or UO_632 (O_632,N_9669,N_8205);
nand UO_633 (O_633,N_7884,N_9901);
nand UO_634 (O_634,N_9651,N_8125);
xnor UO_635 (O_635,N_7635,N_8540);
nor UO_636 (O_636,N_7504,N_8361);
and UO_637 (O_637,N_9073,N_8553);
and UO_638 (O_638,N_8318,N_9803);
and UO_639 (O_639,N_8456,N_9338);
nand UO_640 (O_640,N_8033,N_7722);
nor UO_641 (O_641,N_9168,N_8364);
and UO_642 (O_642,N_9433,N_8108);
or UO_643 (O_643,N_8612,N_9642);
and UO_644 (O_644,N_8687,N_9250);
and UO_645 (O_645,N_9702,N_8040);
nand UO_646 (O_646,N_8204,N_8266);
nor UO_647 (O_647,N_9143,N_9938);
nor UO_648 (O_648,N_8049,N_8533);
nor UO_649 (O_649,N_8501,N_9884);
nand UO_650 (O_650,N_8249,N_8520);
nor UO_651 (O_651,N_8595,N_9707);
and UO_652 (O_652,N_7718,N_8170);
nand UO_653 (O_653,N_8489,N_8869);
nor UO_654 (O_654,N_7891,N_9447);
nand UO_655 (O_655,N_9806,N_8925);
nand UO_656 (O_656,N_9885,N_9353);
or UO_657 (O_657,N_8235,N_8276);
and UO_658 (O_658,N_9344,N_9118);
or UO_659 (O_659,N_7638,N_8863);
or UO_660 (O_660,N_8664,N_8552);
and UO_661 (O_661,N_8569,N_9345);
nor UO_662 (O_662,N_9932,N_9966);
nand UO_663 (O_663,N_7719,N_7588);
nand UO_664 (O_664,N_9636,N_8685);
nor UO_665 (O_665,N_7935,N_8485);
or UO_666 (O_666,N_7730,N_7633);
nand UO_667 (O_667,N_8281,N_8596);
nand UO_668 (O_668,N_7938,N_9357);
nand UO_669 (O_669,N_7840,N_9405);
nor UO_670 (O_670,N_8398,N_8680);
or UO_671 (O_671,N_9418,N_9093);
and UO_672 (O_672,N_9276,N_8201);
and UO_673 (O_673,N_8480,N_8834);
or UO_674 (O_674,N_8451,N_7603);
nor UO_675 (O_675,N_9661,N_8572);
or UO_676 (O_676,N_9745,N_8393);
nor UO_677 (O_677,N_8151,N_7775);
nor UO_678 (O_678,N_9804,N_9247);
nor UO_679 (O_679,N_9778,N_8462);
nand UO_680 (O_680,N_7981,N_7520);
and UO_681 (O_681,N_9101,N_7942);
nor UO_682 (O_682,N_7972,N_9640);
or UO_683 (O_683,N_9786,N_8286);
nand UO_684 (O_684,N_8095,N_9485);
nor UO_685 (O_685,N_7612,N_9920);
and UO_686 (O_686,N_8509,N_8854);
nand UO_687 (O_687,N_9861,N_9967);
nor UO_688 (O_688,N_8976,N_7993);
and UO_689 (O_689,N_9926,N_9421);
and UO_690 (O_690,N_9174,N_9008);
or UO_691 (O_691,N_9121,N_9548);
and UO_692 (O_692,N_9964,N_8245);
or UO_693 (O_693,N_9323,N_8873);
nand UO_694 (O_694,N_9348,N_9550);
or UO_695 (O_695,N_9070,N_7832);
and UO_696 (O_696,N_9360,N_9133);
or UO_697 (O_697,N_9563,N_9846);
and UO_698 (O_698,N_8632,N_9681);
nand UO_699 (O_699,N_8639,N_8598);
and UO_700 (O_700,N_9558,N_8469);
nand UO_701 (O_701,N_9475,N_8091);
nand UO_702 (O_702,N_9426,N_8012);
nand UO_703 (O_703,N_8228,N_7725);
nand UO_704 (O_704,N_9183,N_8218);
nand UO_705 (O_705,N_9361,N_7829);
nand UO_706 (O_706,N_8340,N_8911);
nand UO_707 (O_707,N_9999,N_9626);
and UO_708 (O_708,N_8927,N_8606);
or UO_709 (O_709,N_7909,N_8123);
or UO_710 (O_710,N_7655,N_9238);
or UO_711 (O_711,N_8960,N_9627);
and UO_712 (O_712,N_7746,N_8817);
nor UO_713 (O_713,N_9657,N_8138);
nor UO_714 (O_714,N_7688,N_9016);
nand UO_715 (O_715,N_8769,N_8683);
nand UO_716 (O_716,N_9831,N_7506);
or UO_717 (O_717,N_9526,N_8273);
nor UO_718 (O_718,N_9822,N_9906);
or UO_719 (O_719,N_7794,N_7618);
or UO_720 (O_720,N_9029,N_8498);
or UO_721 (O_721,N_8616,N_8866);
nor UO_722 (O_722,N_9930,N_8097);
or UO_723 (O_723,N_9802,N_8692);
nor UO_724 (O_724,N_7792,N_8920);
or UO_725 (O_725,N_8288,N_8839);
nand UO_726 (O_726,N_8150,N_8679);
or UO_727 (O_727,N_7747,N_9727);
or UO_728 (O_728,N_8874,N_9362);
nor UO_729 (O_729,N_9156,N_8357);
or UO_730 (O_730,N_8793,N_8506);
nand UO_731 (O_731,N_9232,N_9596);
nor UO_732 (O_732,N_9436,N_8514);
and UO_733 (O_733,N_8293,N_8591);
nor UO_734 (O_734,N_8695,N_8070);
nand UO_735 (O_735,N_9478,N_7607);
nor UO_736 (O_736,N_8614,N_8274);
and UO_737 (O_737,N_8436,N_9585);
and UO_738 (O_738,N_8875,N_9941);
nand UO_739 (O_739,N_9068,N_9973);
nand UO_740 (O_740,N_8345,N_9243);
or UO_741 (O_741,N_9172,N_9317);
nand UO_742 (O_742,N_9665,N_8893);
and UO_743 (O_743,N_9441,N_9241);
nor UO_744 (O_744,N_7532,N_9958);
nor UO_745 (O_745,N_9128,N_8155);
nand UO_746 (O_746,N_8299,N_8365);
and UO_747 (O_747,N_9221,N_8849);
and UO_748 (O_748,N_8898,N_8562);
nand UO_749 (O_749,N_8661,N_8625);
and UO_750 (O_750,N_9838,N_9593);
nand UO_751 (O_751,N_7941,N_7896);
nor UO_752 (O_752,N_9820,N_9825);
or UO_753 (O_753,N_9231,N_8923);
and UO_754 (O_754,N_8638,N_9104);
or UO_755 (O_755,N_7971,N_7628);
and UO_756 (O_756,N_8128,N_8763);
or UO_757 (O_757,N_8358,N_9896);
nor UO_758 (O_758,N_8222,N_8603);
and UO_759 (O_759,N_8041,N_8468);
nand UO_760 (O_760,N_8439,N_7515);
nor UO_761 (O_761,N_7584,N_7994);
and UO_762 (O_762,N_7807,N_7526);
or UO_763 (O_763,N_8225,N_9038);
and UO_764 (O_764,N_7995,N_9551);
nor UO_765 (O_765,N_9279,N_9012);
nand UO_766 (O_766,N_8001,N_8392);
or UO_767 (O_767,N_9395,N_8571);
or UO_768 (O_768,N_9600,N_8289);
nand UO_769 (O_769,N_8058,N_7781);
nand UO_770 (O_770,N_9210,N_9033);
or UO_771 (O_771,N_9945,N_7930);
or UO_772 (O_772,N_9810,N_8497);
or UO_773 (O_773,N_8262,N_8717);
nor UO_774 (O_774,N_7756,N_9394);
or UO_775 (O_775,N_9130,N_9060);
nor UO_776 (O_776,N_8089,N_9085);
or UO_777 (O_777,N_9736,N_9986);
or UO_778 (O_778,N_9219,N_8556);
and UO_779 (O_779,N_7985,N_8232);
and UO_780 (O_780,N_7605,N_9261);
and UO_781 (O_781,N_9641,N_9444);
nand UO_782 (O_782,N_8146,N_9005);
and UO_783 (O_783,N_9536,N_8576);
and UO_784 (O_784,N_9166,N_9372);
or UO_785 (O_785,N_7744,N_7937);
and UO_786 (O_786,N_9257,N_9335);
nand UO_787 (O_787,N_7948,N_9202);
nor UO_788 (O_788,N_9225,N_9761);
nor UO_789 (O_789,N_9622,N_9639);
or UO_790 (O_790,N_9504,N_9122);
and UO_791 (O_791,N_9061,N_9387);
and UO_792 (O_792,N_7940,N_9922);
nor UO_793 (O_793,N_8427,N_9579);
nand UO_794 (O_794,N_8301,N_8715);
or UO_795 (O_795,N_7842,N_8088);
and UO_796 (O_796,N_7509,N_8986);
and UO_797 (O_797,N_7869,N_9462);
nand UO_798 (O_798,N_9096,N_8478);
or UO_799 (O_799,N_9473,N_9451);
and UO_800 (O_800,N_8859,N_7561);
nand UO_801 (O_801,N_8975,N_9389);
nor UO_802 (O_802,N_9282,N_8748);
nor UO_803 (O_803,N_8756,N_7902);
nor UO_804 (O_804,N_8157,N_7676);
nor UO_805 (O_805,N_9851,N_8830);
and UO_806 (O_806,N_8846,N_8387);
nor UO_807 (O_807,N_8812,N_8772);
and UO_808 (O_808,N_9608,N_9514);
nand UO_809 (O_809,N_7682,N_9845);
or UO_810 (O_810,N_8045,N_9650);
nor UO_811 (O_811,N_9549,N_8959);
nor UO_812 (O_812,N_9006,N_7650);
nor UO_813 (O_813,N_9285,N_8122);
and UO_814 (O_814,N_8242,N_8104);
or UO_815 (O_815,N_8156,N_8065);
nor UO_816 (O_816,N_9289,N_7822);
nand UO_817 (O_817,N_9040,N_8111);
and UO_818 (O_818,N_9648,N_9259);
or UO_819 (O_819,N_7873,N_9354);
nor UO_820 (O_820,N_9946,N_9091);
nor UO_821 (O_821,N_9754,N_9428);
nor UO_822 (O_822,N_8351,N_8143);
nor UO_823 (O_823,N_9457,N_8391);
nor UO_824 (O_824,N_9779,N_7538);
nand UO_825 (O_825,N_9327,N_8334);
nand UO_826 (O_826,N_7531,N_9242);
nor UO_827 (O_827,N_8199,N_7654);
nor UO_828 (O_828,N_9620,N_7731);
or UO_829 (O_829,N_9297,N_9290);
and UO_830 (O_830,N_9498,N_7788);
nor UO_831 (O_831,N_9951,N_7929);
nor UO_832 (O_832,N_7555,N_8316);
nor UO_833 (O_833,N_9295,N_7647);
or UO_834 (O_834,N_8126,N_8256);
nor UO_835 (O_835,N_9416,N_9785);
nor UO_836 (O_836,N_9124,N_9610);
or UO_837 (O_837,N_7763,N_9409);
and UO_838 (O_838,N_7578,N_8752);
and UO_839 (O_839,N_9499,N_9959);
nor UO_840 (O_840,N_7758,N_9330);
nor UO_841 (O_841,N_8853,N_7568);
nor UO_842 (O_842,N_9722,N_7874);
nor UO_843 (O_843,N_8163,N_9131);
and UO_844 (O_844,N_9201,N_9766);
nand UO_845 (O_845,N_7589,N_9553);
nor UO_846 (O_846,N_9301,N_7779);
and UO_847 (O_847,N_7664,N_7783);
nand UO_848 (O_848,N_8733,N_9886);
and UO_849 (O_849,N_8852,N_7575);
nand UO_850 (O_850,N_8226,N_9725);
or UO_851 (O_851,N_7659,N_7563);
nand UO_852 (O_852,N_8265,N_8646);
nand UO_853 (O_853,N_9393,N_7795);
nor UO_854 (O_854,N_9342,N_7503);
and UO_855 (O_855,N_7903,N_8200);
nor UO_856 (O_856,N_7678,N_9195);
and UO_857 (O_857,N_7567,N_7931);
and UO_858 (O_858,N_9497,N_9382);
nand UO_859 (O_859,N_8884,N_7529);
nor UO_860 (O_860,N_7821,N_8621);
nor UO_861 (O_861,N_8631,N_9995);
nand UO_862 (O_862,N_9860,N_7541);
nor UO_863 (O_863,N_8332,N_9565);
and UO_864 (O_864,N_9664,N_8630);
nand UO_865 (O_865,N_9367,N_8535);
nand UO_866 (O_866,N_9689,N_9525);
and UO_867 (O_867,N_9049,N_8908);
xnor UO_868 (O_868,N_8952,N_9523);
or UO_869 (O_869,N_7773,N_7836);
or UO_870 (O_870,N_7639,N_8272);
nand UO_871 (O_871,N_9868,N_9336);
or UO_872 (O_872,N_7851,N_7921);
and UO_873 (O_873,N_8411,N_9710);
or UO_874 (O_874,N_7886,N_7818);
nand UO_875 (O_875,N_9097,N_9032);
nand UO_876 (O_876,N_7549,N_8303);
or UO_877 (O_877,N_8663,N_9516);
nand UO_878 (O_878,N_8077,N_8804);
nor UO_879 (O_879,N_8238,N_8254);
nor UO_880 (O_880,N_7619,N_8819);
and UO_881 (O_881,N_9883,N_8702);
or UO_882 (O_882,N_8547,N_8833);
nand UO_883 (O_883,N_9493,N_9576);
or UO_884 (O_884,N_8154,N_9039);
or UO_885 (O_885,N_9654,N_8647);
nor UO_886 (O_886,N_8433,N_8945);
nand UO_887 (O_887,N_8229,N_9272);
xor UO_888 (O_888,N_8440,N_7830);
and UO_889 (O_889,N_8472,N_9503);
or UO_890 (O_890,N_9274,N_7918);
or UO_891 (O_891,N_7802,N_9482);
and UO_892 (O_892,N_7608,N_9169);
nor UO_893 (O_893,N_8577,N_8418);
nor UO_894 (O_894,N_9249,N_8924);
nor UO_895 (O_895,N_9866,N_9378);
and UO_896 (O_896,N_9350,N_9856);
and UO_897 (O_897,N_9223,N_9467);
and UO_898 (O_898,N_8588,N_9479);
nor UO_899 (O_899,N_8902,N_9587);
or UO_900 (O_900,N_9998,N_8322);
and UO_901 (O_901,N_9827,N_8635);
or UO_902 (O_902,N_7668,N_9522);
or UO_903 (O_903,N_7614,N_9534);
nor UO_904 (O_904,N_8510,N_8066);
nor UO_905 (O_905,N_9790,N_9283);
or UO_906 (O_906,N_7843,N_9997);
or UO_907 (O_907,N_9145,N_8237);
and UO_908 (O_908,N_8500,N_8905);
nand UO_909 (O_909,N_9302,N_9137);
and UO_910 (O_910,N_8253,N_8449);
nor UO_911 (O_911,N_9606,N_8327);
and UO_912 (O_912,N_8054,N_7649);
nand UO_913 (O_913,N_9415,N_9086);
xor UO_914 (O_914,N_8587,N_8216);
nor UO_915 (O_915,N_8967,N_9737);
nand UO_916 (O_916,N_9025,N_7644);
nand UO_917 (O_917,N_8402,N_9653);
and UO_918 (O_918,N_9373,N_9365);
nand UO_919 (O_919,N_8851,N_8712);
or UO_920 (O_920,N_8491,N_9152);
nor UO_921 (O_921,N_7745,N_7530);
nand UO_922 (O_922,N_9035,N_9656);
and UO_923 (O_923,N_9566,N_7590);
xnor UO_924 (O_924,N_8747,N_7510);
or UO_925 (O_925,N_8826,N_9776);
and UO_926 (O_926,N_8857,N_7825);
and UO_927 (O_927,N_8736,N_8408);
nand UO_928 (O_928,N_8055,N_7750);
nand UO_929 (O_929,N_7507,N_8009);
and UO_930 (O_930,N_8305,N_7629);
nor UO_931 (O_931,N_8876,N_9753);
or UO_932 (O_932,N_9515,N_8658);
nand UO_933 (O_933,N_8669,N_8366);
or UO_934 (O_934,N_9456,N_8706);
or UO_935 (O_935,N_8086,N_9676);
nor UO_936 (O_936,N_8457,N_7681);
nor UO_937 (O_937,N_7591,N_8984);
or UO_938 (O_938,N_9077,N_8581);
nor UO_939 (O_939,N_8350,N_8739);
and UO_940 (O_940,N_9197,N_8549);
or UO_941 (O_941,N_9217,N_8021);
nor UO_942 (O_942,N_9911,N_7522);
and UO_943 (O_943,N_7641,N_9703);
nor UO_944 (O_944,N_9872,N_9524);
or UO_945 (O_945,N_8559,N_9644);
or UO_946 (O_946,N_7669,N_8494);
or UO_947 (O_947,N_8136,N_8990);
or UO_948 (O_948,N_8168,N_9718);
nor UO_949 (O_949,N_7932,N_8972);
nand UO_950 (O_950,N_8371,N_9324);
nor UO_951 (O_951,N_8512,N_9517);
and UO_952 (O_952,N_9616,N_8617);
nor UO_953 (O_953,N_7505,N_8337);
and UO_954 (O_954,N_8623,N_9843);
and UO_955 (O_955,N_8190,N_8307);
nor UO_956 (O_956,N_8889,N_7956);
nor UO_957 (O_957,N_8096,N_7556);
nand UO_958 (O_958,N_7811,N_7887);
nand UO_959 (O_959,N_8691,N_7596);
nand UO_960 (O_960,N_9160,N_8434);
and UO_961 (O_961,N_8704,N_9541);
nand UO_962 (O_962,N_8135,N_8443);
and UO_963 (O_963,N_8169,N_8737);
nand UO_964 (O_964,N_9671,N_8233);
or UO_965 (O_965,N_8832,N_7670);
nand UO_966 (O_966,N_9836,N_8348);
or UO_967 (O_967,N_9817,N_8921);
nor UO_968 (O_968,N_8568,N_7692);
nand UO_969 (O_969,N_8771,N_7525);
nand UO_970 (O_970,N_9376,N_8324);
or UO_971 (O_971,N_7844,N_8555);
nor UO_972 (O_972,N_8377,N_8129);
nand UO_973 (O_973,N_9777,N_7711);
nor UO_974 (O_974,N_7751,N_9873);
nor UO_975 (O_975,N_9334,N_8140);
nor UO_976 (O_976,N_9264,N_9170);
nor UO_977 (O_977,N_7980,N_9246);
nor UO_978 (O_978,N_9569,N_8659);
or UO_979 (O_979,N_8649,N_8435);
nor UO_980 (O_980,N_8189,N_7564);
nand UO_981 (O_981,N_8744,N_8052);
nor UO_982 (O_982,N_9679,N_7833);
or UO_983 (O_983,N_8665,N_7599);
or UO_984 (O_984,N_8330,N_8601);
nand UO_985 (O_985,N_8788,N_8432);
nand UO_986 (O_986,N_7706,N_8425);
and UO_987 (O_987,N_7565,N_8207);
or UO_988 (O_988,N_8466,N_8084);
nor UO_989 (O_989,N_8159,N_8613);
nand UO_990 (O_990,N_9281,N_8263);
and UO_991 (O_991,N_9598,N_7965);
and UO_992 (O_992,N_7955,N_8696);
or UO_993 (O_993,N_7834,N_9673);
and UO_994 (O_994,N_8810,N_8448);
nor UO_995 (O_995,N_8459,N_8989);
and UO_996 (O_996,N_8100,N_8903);
nand UO_997 (O_997,N_9555,N_9046);
nand UO_998 (O_998,N_9374,N_9685);
and UO_999 (O_999,N_8083,N_9140);
nor UO_1000 (O_1000,N_9472,N_9538);
and UO_1001 (O_1001,N_9659,N_9581);
nand UO_1002 (O_1002,N_9562,N_7828);
nand UO_1003 (O_1003,N_7653,N_8796);
and UO_1004 (O_1004,N_8724,N_8782);
nand UO_1005 (O_1005,N_8809,N_9647);
nand UO_1006 (O_1006,N_9800,N_7705);
nor UO_1007 (O_1007,N_9905,N_8939);
nand UO_1008 (O_1008,N_9878,N_9173);
and UO_1009 (O_1009,N_9213,N_8132);
nor UO_1010 (O_1010,N_9783,N_8325);
or UO_1011 (O_1011,N_9691,N_8940);
nor UO_1012 (O_1012,N_7968,N_8484);
nand UO_1013 (O_1013,N_9764,N_8671);
nand UO_1014 (O_1014,N_8373,N_8951);
and UO_1015 (O_1015,N_8020,N_7723);
nor UO_1016 (O_1016,N_7870,N_7696);
xnor UO_1017 (O_1017,N_9533,N_8622);
or UO_1018 (O_1018,N_9506,N_8465);
or UO_1019 (O_1019,N_9181,N_9399);
nor UO_1020 (O_1020,N_9993,N_7536);
and UO_1021 (O_1021,N_8686,N_7593);
nor UO_1022 (O_1022,N_9175,N_8102);
nor UO_1023 (O_1023,N_7759,N_8803);
and UO_1024 (O_1024,N_9023,N_8881);
and UO_1025 (O_1025,N_9044,N_7566);
nor UO_1026 (O_1026,N_8246,N_9957);
nor UO_1027 (O_1027,N_9268,N_9532);
nand UO_1028 (O_1028,N_8640,N_8454);
or UO_1029 (O_1029,N_7899,N_7817);
nor UO_1030 (O_1030,N_9400,N_8980);
and UO_1031 (O_1031,N_7867,N_8892);
or UO_1032 (O_1032,N_9459,N_9985);
nand UO_1033 (O_1033,N_8116,N_8115);
or UO_1034 (O_1034,N_9007,N_8926);
nand UO_1035 (O_1035,N_7976,N_7764);
or UO_1036 (O_1036,N_8811,N_7939);
or UO_1037 (O_1037,N_9615,N_8773);
nand UO_1038 (O_1038,N_9385,N_9431);
and UO_1039 (O_1039,N_9686,N_9716);
nand UO_1040 (O_1040,N_9437,N_9188);
nand UO_1041 (O_1041,N_9990,N_9189);
or UO_1042 (O_1042,N_8271,N_7548);
nor UO_1043 (O_1043,N_8633,N_9723);
nand UO_1044 (O_1044,N_7966,N_9542);
and UO_1045 (O_1045,N_8446,N_7580);
nor UO_1046 (O_1046,N_7729,N_7983);
nand UO_1047 (O_1047,N_7632,N_7838);
and UO_1048 (O_1048,N_9652,N_8888);
nor UO_1049 (O_1049,N_9349,N_9809);
nor UO_1050 (O_1050,N_8800,N_9853);
or UO_1051 (O_1051,N_8413,N_9461);
nand UO_1052 (O_1052,N_8320,N_8517);
and UO_1053 (O_1053,N_9309,N_7767);
and UO_1054 (O_1054,N_9022,N_9028);
or UO_1055 (O_1055,N_9667,N_8011);
nor UO_1056 (O_1056,N_8504,N_7665);
nand UO_1057 (O_1057,N_9352,N_8779);
and UO_1058 (O_1058,N_8261,N_8700);
xnor UO_1059 (O_1059,N_8010,N_9031);
or UO_1060 (O_1060,N_9075,N_8891);
nand UO_1061 (O_1061,N_9138,N_9939);
and UO_1062 (O_1062,N_8618,N_9781);
nand UO_1063 (O_1063,N_8000,N_9700);
nor UO_1064 (O_1064,N_9414,N_9230);
and UO_1065 (O_1065,N_7637,N_7881);
or UO_1066 (O_1066,N_9390,N_8044);
or UO_1067 (O_1067,N_7609,N_9011);
or UO_1068 (O_1068,N_7626,N_9752);
nor UO_1069 (O_1069,N_8153,N_9446);
nor UO_1070 (O_1070,N_8785,N_8988);
nand UO_1071 (O_1071,N_8732,N_9358);
or UO_1072 (O_1072,N_9116,N_9233);
or UO_1073 (O_1073,N_9132,N_8158);
nand UO_1074 (O_1074,N_8670,N_9209);
nand UO_1075 (O_1075,N_8240,N_7933);
xnor UO_1076 (O_1076,N_7569,N_9255);
and UO_1077 (O_1077,N_7907,N_9591);
and UO_1078 (O_1078,N_8087,N_9518);
and UO_1079 (O_1079,N_9887,N_7928);
and UO_1080 (O_1080,N_7643,N_8722);
or UO_1081 (O_1081,N_8962,N_8628);
and UO_1082 (O_1082,N_7660,N_9955);
and UO_1083 (O_1083,N_8428,N_9293);
or UO_1084 (O_1084,N_7979,N_8557);
nor UO_1085 (O_1085,N_9305,N_7517);
and UO_1086 (O_1086,N_7602,N_8579);
nor UO_1087 (O_1087,N_8369,N_9325);
and UO_1088 (O_1088,N_9739,N_9796);
xnor UO_1089 (O_1089,N_8082,N_7787);
nor UO_1090 (O_1090,N_9013,N_8403);
nor UO_1091 (O_1091,N_9889,N_8541);
or UO_1092 (O_1092,N_8499,N_8186);
nor UO_1093 (O_1093,N_8843,N_8343);
nor UO_1094 (O_1094,N_8742,N_8765);
or UO_1095 (O_1095,N_9697,N_9834);
nand UO_1096 (O_1096,N_8590,N_9728);
nand UO_1097 (O_1097,N_9351,N_9204);
and UO_1098 (O_1098,N_8886,N_9613);
or UO_1099 (O_1099,N_7600,N_7959);
or UO_1100 (O_1100,N_7790,N_8847);
nand UO_1101 (O_1101,N_8187,N_8455);
nor UO_1102 (O_1102,N_7917,N_9837);
nand UO_1103 (O_1103,N_7799,N_9384);
or UO_1104 (O_1104,N_8776,N_8349);
xnor UO_1105 (O_1105,N_9821,N_9908);
nand UO_1106 (O_1106,N_9726,N_8652);
or UO_1107 (O_1107,N_9157,N_8422);
or UO_1108 (O_1108,N_8016,N_8166);
nor UO_1109 (O_1109,N_8992,N_9792);
nand UO_1110 (O_1110,N_9337,N_9280);
nor UO_1111 (O_1111,N_9732,N_8046);
nand UO_1112 (O_1112,N_8582,N_8374);
and UO_1113 (O_1113,N_8236,N_7586);
nand UO_1114 (O_1114,N_7944,N_8668);
or UO_1115 (O_1115,N_8532,N_9134);
and UO_1116 (O_1116,N_8505,N_9891);
and UO_1117 (O_1117,N_9026,N_9460);
nor UO_1118 (O_1118,N_9816,N_7882);
nand UO_1119 (O_1119,N_7557,N_8619);
and UO_1120 (O_1120,N_8213,N_9326);
nand UO_1121 (O_1121,N_8774,N_7674);
nor UO_1122 (O_1122,N_8624,N_7757);
and UO_1123 (O_1123,N_9486,N_8362);
nand UO_1124 (O_1124,N_9611,N_8870);
nand UO_1125 (O_1125,N_9245,N_9794);
nand UO_1126 (O_1126,N_9150,N_9812);
and UO_1127 (O_1127,N_8078,N_9801);
nor UO_1128 (O_1128,N_8255,N_9936);
nand UO_1129 (O_1129,N_8675,N_8092);
nand UO_1130 (O_1130,N_9590,N_7947);
nand UO_1131 (O_1131,N_7540,N_9537);
and UO_1132 (O_1132,N_8198,N_8423);
xor UO_1133 (O_1133,N_9612,N_8584);
nor UO_1134 (O_1134,N_7624,N_9680);
nor UO_1135 (O_1135,N_8405,N_9624);
and UO_1136 (O_1136,N_7727,N_8592);
nand UO_1137 (O_1137,N_9530,N_8667);
and UO_1138 (O_1138,N_8835,N_8388);
nor UO_1139 (O_1139,N_9907,N_8551);
nor UO_1140 (O_1140,N_9037,N_8821);
and UO_1141 (O_1141,N_8678,N_9294);
nand UO_1142 (O_1142,N_7735,N_9633);
or UO_1143 (O_1143,N_8298,N_8094);
or UO_1144 (O_1144,N_8259,N_9709);
or UO_1145 (O_1145,N_8260,N_9052);
or UO_1146 (O_1146,N_8599,N_8214);
or UO_1147 (O_1147,N_9544,N_9051);
nor UO_1148 (O_1148,N_8396,N_8971);
nand UO_1149 (O_1149,N_7697,N_8173);
and UO_1150 (O_1150,N_9228,N_9043);
or UO_1151 (O_1151,N_9303,N_8031);
nand UO_1152 (O_1152,N_7999,N_7726);
nor UO_1153 (O_1153,N_9218,N_8162);
nand UO_1154 (O_1154,N_9266,N_9135);
and UO_1155 (O_1155,N_9176,N_9704);
nor UO_1156 (O_1156,N_7671,N_9064);
and UO_1157 (O_1157,N_9505,N_9308);
and UO_1158 (O_1158,N_8264,N_8968);
or UO_1159 (O_1159,N_8367,N_8731);
and UO_1160 (O_1160,N_8820,N_8828);
nor UO_1161 (O_1161,N_7805,N_9683);
nor UO_1162 (O_1162,N_8037,N_9928);
nor UO_1163 (O_1163,N_9589,N_8550);
nor UO_1164 (O_1164,N_9535,N_9867);
nand UO_1165 (O_1165,N_9180,N_7558);
and UO_1166 (O_1166,N_7514,N_8656);
nand UO_1167 (O_1167,N_9742,N_9835);
nand UO_1168 (O_1168,N_7673,N_9947);
nand UO_1169 (O_1169,N_8496,N_8080);
nor UO_1170 (O_1170,N_8336,N_9773);
and UO_1171 (O_1171,N_9235,N_9434);
nand UO_1172 (O_1172,N_7528,N_9980);
nor UO_1173 (O_1173,N_8716,N_9829);
or UO_1174 (O_1174,N_7803,N_9316);
nor UO_1175 (O_1175,N_8734,N_7611);
nor UO_1176 (O_1176,N_9468,N_9841);
nor UO_1177 (O_1177,N_9369,N_9034);
and UO_1178 (O_1178,N_7714,N_9392);
and UO_1179 (O_1179,N_7988,N_7915);
nor UO_1180 (O_1180,N_9287,N_8120);
nor UO_1181 (O_1181,N_7953,N_9900);
nor UO_1182 (O_1182,N_8414,N_8234);
nor UO_1183 (O_1183,N_8030,N_7839);
nand UO_1184 (O_1184,N_8121,N_9675);
or UO_1185 (O_1185,N_9300,N_9942);
nor UO_1186 (O_1186,N_9222,N_7537);
nand UO_1187 (O_1187,N_8471,N_7796);
nand UO_1188 (O_1188,N_9601,N_7866);
and UO_1189 (O_1189,N_7693,N_8051);
or UO_1190 (O_1190,N_9762,N_9438);
nor UO_1191 (O_1191,N_8919,N_9751);
or UO_1192 (O_1192,N_8701,N_8714);
nand UO_1193 (O_1193,N_9126,N_9449);
nor UO_1194 (O_1194,N_9758,N_9076);
nand UO_1195 (O_1195,N_7893,N_9529);
nor UO_1196 (O_1196,N_7831,N_8978);
and UO_1197 (O_1197,N_9312,N_8297);
nand UO_1198 (O_1198,N_8179,N_8292);
nor UO_1199 (O_1199,N_8194,N_7782);
nand UO_1200 (O_1200,N_8503,N_9968);
nor UO_1201 (O_1201,N_9988,N_8743);
or UO_1202 (O_1202,N_9445,N_8149);
or UO_1203 (O_1203,N_9953,N_8032);
and UO_1204 (O_1204,N_9925,N_8787);
nor UO_1205 (O_1205,N_7577,N_9979);
or UO_1206 (O_1206,N_8727,N_8899);
nor UO_1207 (O_1207,N_7721,N_9917);
nand UO_1208 (O_1208,N_7963,N_8674);
nor UO_1209 (O_1209,N_8479,N_8900);
nor UO_1210 (O_1210,N_9730,N_9850);
nand UO_1211 (O_1211,N_8825,N_8287);
nand UO_1212 (O_1212,N_7892,N_7934);
or UO_1213 (O_1213,N_8831,N_9430);
and UO_1214 (O_1214,N_9818,N_9179);
and UO_1215 (O_1215,N_9396,N_8915);
nand UO_1216 (O_1216,N_7875,N_9072);
nor UO_1217 (O_1217,N_9355,N_9706);
nand UO_1218 (O_1218,N_8637,N_7636);
nor UO_1219 (O_1219,N_9319,N_9711);
and UO_1220 (O_1220,N_9476,N_8868);
nor UO_1221 (O_1221,N_7967,N_7604);
nand UO_1222 (O_1222,N_9260,N_8690);
nor UO_1223 (O_1223,N_9962,N_9748);
and UO_1224 (O_1224,N_9631,N_8385);
nor UO_1225 (O_1225,N_9178,N_9194);
nand UO_1226 (O_1226,N_9141,N_9780);
nor UO_1227 (O_1227,N_9577,N_7741);
or UO_1228 (O_1228,N_8895,N_8006);
and UO_1229 (O_1229,N_9401,N_9411);
nor UO_1230 (O_1230,N_9571,N_7957);
nor UO_1231 (O_1231,N_7646,N_9693);
and UO_1232 (O_1232,N_8107,N_9054);
and UO_1233 (O_1233,N_9488,N_9509);
nor UO_1234 (O_1234,N_9477,N_9760);
nand UO_1235 (O_1235,N_9767,N_8916);
nor UO_1236 (O_1236,N_9240,N_8777);
nor UO_1237 (O_1237,N_9520,N_9465);
or UO_1238 (O_1238,N_9448,N_8172);
nand UO_1239 (O_1239,N_8090,N_7778);
nand UO_1240 (O_1240,N_9481,N_7554);
and UO_1241 (O_1241,N_9100,N_8605);
nor UO_1242 (O_1242,N_9614,N_8319);
and UO_1243 (O_1243,N_7737,N_9496);
and UO_1244 (O_1244,N_8134,N_7954);
or UO_1245 (O_1245,N_9771,N_9560);
nand UO_1246 (O_1246,N_9252,N_7500);
and UO_1247 (O_1247,N_8511,N_7581);
or UO_1248 (O_1248,N_8730,N_9311);
nor UO_1249 (O_1249,N_7771,N_9427);
or UO_1250 (O_1250,N_9289,N_8752);
and UO_1251 (O_1251,N_8930,N_9615);
nor UO_1252 (O_1252,N_9601,N_9479);
or UO_1253 (O_1253,N_9623,N_8124);
or UO_1254 (O_1254,N_8566,N_8315);
and UO_1255 (O_1255,N_9451,N_9076);
and UO_1256 (O_1256,N_9105,N_9437);
and UO_1257 (O_1257,N_9904,N_7629);
nor UO_1258 (O_1258,N_9987,N_7570);
nand UO_1259 (O_1259,N_9057,N_9448);
and UO_1260 (O_1260,N_9158,N_8306);
and UO_1261 (O_1261,N_8625,N_9008);
nand UO_1262 (O_1262,N_9387,N_8342);
nor UO_1263 (O_1263,N_9079,N_8002);
and UO_1264 (O_1264,N_7904,N_8361);
nand UO_1265 (O_1265,N_8830,N_8932);
or UO_1266 (O_1266,N_9393,N_9162);
and UO_1267 (O_1267,N_7739,N_8510);
and UO_1268 (O_1268,N_8178,N_9144);
nand UO_1269 (O_1269,N_9718,N_8613);
or UO_1270 (O_1270,N_7873,N_8689);
nand UO_1271 (O_1271,N_9944,N_9028);
nor UO_1272 (O_1272,N_8804,N_8326);
nand UO_1273 (O_1273,N_8823,N_7819);
or UO_1274 (O_1274,N_8272,N_9709);
nand UO_1275 (O_1275,N_9768,N_7978);
and UO_1276 (O_1276,N_8054,N_9040);
or UO_1277 (O_1277,N_8225,N_8368);
nor UO_1278 (O_1278,N_9461,N_9459);
and UO_1279 (O_1279,N_9074,N_7916);
nor UO_1280 (O_1280,N_8442,N_8045);
or UO_1281 (O_1281,N_9933,N_8880);
and UO_1282 (O_1282,N_7649,N_7594);
nor UO_1283 (O_1283,N_7899,N_8891);
nor UO_1284 (O_1284,N_8916,N_8863);
or UO_1285 (O_1285,N_9237,N_8780);
and UO_1286 (O_1286,N_8554,N_8258);
and UO_1287 (O_1287,N_9630,N_8875);
and UO_1288 (O_1288,N_9113,N_9660);
nor UO_1289 (O_1289,N_9326,N_8479);
xor UO_1290 (O_1290,N_9536,N_9660);
and UO_1291 (O_1291,N_9696,N_8530);
nand UO_1292 (O_1292,N_8575,N_8090);
nand UO_1293 (O_1293,N_7685,N_7905);
nand UO_1294 (O_1294,N_8967,N_8920);
nor UO_1295 (O_1295,N_9433,N_9330);
nor UO_1296 (O_1296,N_8372,N_7961);
nand UO_1297 (O_1297,N_8835,N_7554);
nand UO_1298 (O_1298,N_8052,N_9473);
or UO_1299 (O_1299,N_9951,N_8863);
and UO_1300 (O_1300,N_8594,N_8673);
or UO_1301 (O_1301,N_8439,N_9832);
or UO_1302 (O_1302,N_8418,N_9642);
nand UO_1303 (O_1303,N_7626,N_8379);
nor UO_1304 (O_1304,N_9157,N_9333);
and UO_1305 (O_1305,N_8966,N_8776);
or UO_1306 (O_1306,N_9617,N_8544);
and UO_1307 (O_1307,N_8364,N_9475);
nand UO_1308 (O_1308,N_8615,N_7580);
nor UO_1309 (O_1309,N_9677,N_8665);
nand UO_1310 (O_1310,N_7723,N_9834);
or UO_1311 (O_1311,N_9408,N_9915);
nand UO_1312 (O_1312,N_8337,N_9877);
nand UO_1313 (O_1313,N_8406,N_9737);
and UO_1314 (O_1314,N_9662,N_9289);
nand UO_1315 (O_1315,N_8199,N_8471);
nand UO_1316 (O_1316,N_9646,N_9284);
nand UO_1317 (O_1317,N_9715,N_9746);
or UO_1318 (O_1318,N_8362,N_8941);
and UO_1319 (O_1319,N_8895,N_9238);
and UO_1320 (O_1320,N_7704,N_7633);
nand UO_1321 (O_1321,N_9775,N_8701);
nor UO_1322 (O_1322,N_8027,N_8702);
nor UO_1323 (O_1323,N_8131,N_9197);
nand UO_1324 (O_1324,N_9531,N_9159);
nand UO_1325 (O_1325,N_8779,N_9716);
and UO_1326 (O_1326,N_8456,N_9301);
and UO_1327 (O_1327,N_8730,N_8587);
or UO_1328 (O_1328,N_9250,N_8374);
and UO_1329 (O_1329,N_9344,N_9750);
or UO_1330 (O_1330,N_7592,N_8297);
and UO_1331 (O_1331,N_7722,N_9674);
or UO_1332 (O_1332,N_8918,N_7663);
and UO_1333 (O_1333,N_8841,N_9927);
or UO_1334 (O_1334,N_7652,N_9890);
or UO_1335 (O_1335,N_8561,N_8025);
nor UO_1336 (O_1336,N_8281,N_8813);
and UO_1337 (O_1337,N_8620,N_8573);
or UO_1338 (O_1338,N_7626,N_9696);
or UO_1339 (O_1339,N_9952,N_9161);
nor UO_1340 (O_1340,N_9250,N_8865);
nand UO_1341 (O_1341,N_8421,N_8827);
nor UO_1342 (O_1342,N_9881,N_9024);
nor UO_1343 (O_1343,N_9752,N_9256);
nor UO_1344 (O_1344,N_9678,N_8103);
nor UO_1345 (O_1345,N_8949,N_9194);
nor UO_1346 (O_1346,N_8741,N_8112);
and UO_1347 (O_1347,N_9481,N_8721);
nor UO_1348 (O_1348,N_9281,N_9491);
or UO_1349 (O_1349,N_8905,N_8068);
nor UO_1350 (O_1350,N_9109,N_9381);
nor UO_1351 (O_1351,N_9026,N_7958);
and UO_1352 (O_1352,N_8037,N_8201);
and UO_1353 (O_1353,N_8482,N_9070);
or UO_1354 (O_1354,N_7965,N_9587);
nor UO_1355 (O_1355,N_7763,N_9436);
nor UO_1356 (O_1356,N_8149,N_9080);
and UO_1357 (O_1357,N_9958,N_7663);
and UO_1358 (O_1358,N_9762,N_9393);
or UO_1359 (O_1359,N_8846,N_9848);
and UO_1360 (O_1360,N_7792,N_7653);
and UO_1361 (O_1361,N_9749,N_8779);
nor UO_1362 (O_1362,N_8640,N_9256);
or UO_1363 (O_1363,N_8913,N_7862);
nand UO_1364 (O_1364,N_9213,N_9593);
or UO_1365 (O_1365,N_9626,N_9206);
or UO_1366 (O_1366,N_9109,N_8076);
nor UO_1367 (O_1367,N_7507,N_8416);
or UO_1368 (O_1368,N_8476,N_7775);
nor UO_1369 (O_1369,N_8451,N_9855);
or UO_1370 (O_1370,N_9836,N_9755);
and UO_1371 (O_1371,N_8809,N_8572);
and UO_1372 (O_1372,N_9265,N_9436);
or UO_1373 (O_1373,N_9522,N_7757);
nand UO_1374 (O_1374,N_8196,N_8445);
nor UO_1375 (O_1375,N_9153,N_8238);
nand UO_1376 (O_1376,N_9180,N_7687);
nor UO_1377 (O_1377,N_7542,N_9596);
or UO_1378 (O_1378,N_8076,N_8838);
or UO_1379 (O_1379,N_9427,N_9128);
or UO_1380 (O_1380,N_8043,N_7876);
nor UO_1381 (O_1381,N_8429,N_9822);
or UO_1382 (O_1382,N_9437,N_9374);
nand UO_1383 (O_1383,N_7929,N_8264);
and UO_1384 (O_1384,N_9480,N_7936);
or UO_1385 (O_1385,N_9882,N_8258);
nand UO_1386 (O_1386,N_9242,N_8664);
nand UO_1387 (O_1387,N_9806,N_7524);
nor UO_1388 (O_1388,N_7548,N_9142);
nand UO_1389 (O_1389,N_9221,N_9549);
or UO_1390 (O_1390,N_9475,N_8190);
nand UO_1391 (O_1391,N_9393,N_8998);
nand UO_1392 (O_1392,N_8639,N_9482);
nand UO_1393 (O_1393,N_9494,N_7702);
and UO_1394 (O_1394,N_8215,N_9324);
nor UO_1395 (O_1395,N_7518,N_7792);
nor UO_1396 (O_1396,N_8302,N_9064);
or UO_1397 (O_1397,N_8920,N_7796);
nor UO_1398 (O_1398,N_9902,N_8323);
and UO_1399 (O_1399,N_8452,N_8886);
nand UO_1400 (O_1400,N_8965,N_8781);
and UO_1401 (O_1401,N_9739,N_8582);
nor UO_1402 (O_1402,N_9632,N_9502);
or UO_1403 (O_1403,N_9273,N_8679);
nor UO_1404 (O_1404,N_7994,N_8381);
and UO_1405 (O_1405,N_9505,N_9620);
or UO_1406 (O_1406,N_8313,N_8876);
nand UO_1407 (O_1407,N_7706,N_8215);
nand UO_1408 (O_1408,N_8624,N_7651);
nand UO_1409 (O_1409,N_9561,N_7758);
xor UO_1410 (O_1410,N_8372,N_8746);
nand UO_1411 (O_1411,N_8812,N_9210);
nand UO_1412 (O_1412,N_8233,N_8948);
and UO_1413 (O_1413,N_8831,N_8088);
nor UO_1414 (O_1414,N_7516,N_9036);
nor UO_1415 (O_1415,N_9621,N_9251);
nand UO_1416 (O_1416,N_8945,N_9845);
nor UO_1417 (O_1417,N_9736,N_9301);
nor UO_1418 (O_1418,N_8302,N_8813);
nor UO_1419 (O_1419,N_8706,N_9030);
or UO_1420 (O_1420,N_8544,N_7970);
and UO_1421 (O_1421,N_8301,N_9228);
nor UO_1422 (O_1422,N_8205,N_8996);
nor UO_1423 (O_1423,N_8929,N_7995);
nand UO_1424 (O_1424,N_8334,N_9092);
nor UO_1425 (O_1425,N_9593,N_8010);
nor UO_1426 (O_1426,N_8678,N_8125);
nand UO_1427 (O_1427,N_9100,N_8716);
nand UO_1428 (O_1428,N_8200,N_8916);
nor UO_1429 (O_1429,N_8865,N_9278);
or UO_1430 (O_1430,N_7778,N_9550);
nor UO_1431 (O_1431,N_8139,N_8214);
or UO_1432 (O_1432,N_7992,N_9396);
nor UO_1433 (O_1433,N_9978,N_9090);
and UO_1434 (O_1434,N_9822,N_9404);
nand UO_1435 (O_1435,N_7614,N_8502);
and UO_1436 (O_1436,N_8345,N_8760);
nand UO_1437 (O_1437,N_8191,N_9124);
and UO_1438 (O_1438,N_8480,N_9715);
nor UO_1439 (O_1439,N_9455,N_8404);
or UO_1440 (O_1440,N_8496,N_9013);
and UO_1441 (O_1441,N_8954,N_7523);
nor UO_1442 (O_1442,N_8236,N_8865);
nand UO_1443 (O_1443,N_7758,N_9281);
and UO_1444 (O_1444,N_7885,N_7638);
nor UO_1445 (O_1445,N_8542,N_9277);
and UO_1446 (O_1446,N_7964,N_9257);
and UO_1447 (O_1447,N_8157,N_9869);
or UO_1448 (O_1448,N_8965,N_8597);
and UO_1449 (O_1449,N_8507,N_9402);
and UO_1450 (O_1450,N_9156,N_9017);
nor UO_1451 (O_1451,N_7874,N_8946);
or UO_1452 (O_1452,N_8854,N_8291);
and UO_1453 (O_1453,N_9352,N_9128);
nor UO_1454 (O_1454,N_7542,N_9799);
nor UO_1455 (O_1455,N_8083,N_8703);
nand UO_1456 (O_1456,N_8786,N_8614);
and UO_1457 (O_1457,N_8066,N_9364);
xnor UO_1458 (O_1458,N_7671,N_9652);
nor UO_1459 (O_1459,N_9367,N_8038);
or UO_1460 (O_1460,N_8623,N_7800);
and UO_1461 (O_1461,N_9949,N_9543);
nand UO_1462 (O_1462,N_7509,N_8589);
nor UO_1463 (O_1463,N_8022,N_8332);
nor UO_1464 (O_1464,N_9695,N_8257);
nand UO_1465 (O_1465,N_7972,N_7878);
nor UO_1466 (O_1466,N_8486,N_8799);
nor UO_1467 (O_1467,N_8764,N_7719);
nor UO_1468 (O_1468,N_7622,N_7837);
nand UO_1469 (O_1469,N_9773,N_8380);
or UO_1470 (O_1470,N_9986,N_9660);
nor UO_1471 (O_1471,N_8842,N_8439);
nand UO_1472 (O_1472,N_8660,N_9592);
nor UO_1473 (O_1473,N_8938,N_8057);
and UO_1474 (O_1474,N_8641,N_8076);
or UO_1475 (O_1475,N_8605,N_8259);
nor UO_1476 (O_1476,N_7807,N_8628);
and UO_1477 (O_1477,N_7716,N_8292);
nand UO_1478 (O_1478,N_7959,N_7619);
or UO_1479 (O_1479,N_8447,N_8020);
nor UO_1480 (O_1480,N_8009,N_9440);
xor UO_1481 (O_1481,N_8467,N_7687);
or UO_1482 (O_1482,N_9321,N_9075);
xor UO_1483 (O_1483,N_7809,N_9752);
nor UO_1484 (O_1484,N_9394,N_9247);
nor UO_1485 (O_1485,N_7587,N_8613);
nand UO_1486 (O_1486,N_9069,N_7743);
nor UO_1487 (O_1487,N_7562,N_7685);
and UO_1488 (O_1488,N_8267,N_9381);
nor UO_1489 (O_1489,N_8238,N_7958);
nand UO_1490 (O_1490,N_9592,N_9214);
nor UO_1491 (O_1491,N_9096,N_7996);
and UO_1492 (O_1492,N_9343,N_8600);
or UO_1493 (O_1493,N_7659,N_9262);
or UO_1494 (O_1494,N_8986,N_9847);
xor UO_1495 (O_1495,N_9478,N_7895);
nand UO_1496 (O_1496,N_7618,N_7910);
nand UO_1497 (O_1497,N_9111,N_8262);
or UO_1498 (O_1498,N_8561,N_9172);
and UO_1499 (O_1499,N_8340,N_8274);
endmodule