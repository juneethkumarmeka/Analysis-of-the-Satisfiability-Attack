module basic_500_3000_500_4_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xor U0 (N_0,In_311,In_293);
nor U1 (N_1,In_7,In_199);
nand U2 (N_2,In_418,In_137);
nor U3 (N_3,In_61,In_236);
nand U4 (N_4,In_89,In_366);
and U5 (N_5,In_120,In_150);
nor U6 (N_6,In_456,In_361);
nor U7 (N_7,In_422,In_63);
and U8 (N_8,In_154,In_388);
and U9 (N_9,In_95,In_303);
nor U10 (N_10,In_281,In_9);
nand U11 (N_11,In_149,In_56);
nor U12 (N_12,In_110,In_255);
or U13 (N_13,In_104,In_486);
nor U14 (N_14,In_93,In_333);
and U15 (N_15,In_175,In_403);
or U16 (N_16,In_329,In_233);
or U17 (N_17,In_390,In_477);
nor U18 (N_18,In_379,In_2);
or U19 (N_19,In_256,In_392);
and U20 (N_20,In_204,In_259);
nand U21 (N_21,In_36,In_28);
nor U22 (N_22,In_44,In_444);
nand U23 (N_23,In_414,In_463);
or U24 (N_24,In_340,In_365);
nand U25 (N_25,In_373,In_319);
and U26 (N_26,In_29,In_399);
nor U27 (N_27,In_431,In_242);
and U28 (N_28,In_409,In_119);
or U29 (N_29,In_32,In_135);
nor U30 (N_30,In_84,In_107);
and U31 (N_31,In_5,In_467);
and U32 (N_32,In_35,In_201);
and U33 (N_33,In_100,In_453);
and U34 (N_34,In_45,In_384);
nor U35 (N_35,In_307,In_315);
nand U36 (N_36,In_429,In_24);
nand U37 (N_37,In_218,In_23);
nand U38 (N_38,In_219,In_326);
or U39 (N_39,In_336,In_332);
or U40 (N_40,In_142,In_160);
nand U41 (N_41,In_254,In_98);
or U42 (N_42,In_64,In_1);
and U43 (N_43,In_54,In_368);
nor U44 (N_44,In_72,In_216);
and U45 (N_45,In_251,In_480);
nand U46 (N_46,In_442,In_113);
nand U47 (N_47,In_260,In_277);
or U48 (N_48,In_447,In_144);
or U49 (N_49,In_434,In_435);
or U50 (N_50,In_286,In_33);
and U51 (N_51,In_300,In_128);
nor U52 (N_52,In_198,In_173);
nand U53 (N_53,In_401,In_306);
or U54 (N_54,In_168,In_481);
nand U55 (N_55,In_343,In_375);
and U56 (N_56,In_17,In_385);
or U57 (N_57,In_408,In_102);
or U58 (N_58,In_404,In_186);
nand U59 (N_59,In_237,In_147);
nand U60 (N_60,In_280,In_351);
nand U61 (N_61,In_499,In_289);
nand U62 (N_62,In_416,In_91);
xor U63 (N_63,In_158,In_202);
or U64 (N_64,In_490,In_352);
or U65 (N_65,In_164,In_125);
nor U66 (N_66,In_3,In_347);
and U67 (N_67,In_151,In_139);
or U68 (N_68,In_90,In_492);
and U69 (N_69,In_493,In_71);
and U70 (N_70,In_180,In_483);
and U71 (N_71,In_181,In_389);
or U72 (N_72,In_349,In_318);
nand U73 (N_73,In_275,In_417);
and U74 (N_74,In_439,In_288);
nand U75 (N_75,In_10,In_257);
and U76 (N_76,In_155,In_383);
nand U77 (N_77,In_121,In_213);
nor U78 (N_78,In_79,In_226);
nor U79 (N_79,In_356,In_443);
or U80 (N_80,In_305,In_245);
and U81 (N_81,In_203,In_126);
nor U82 (N_82,In_425,In_432);
nor U83 (N_83,In_327,In_75);
and U84 (N_84,In_469,In_210);
and U85 (N_85,In_369,In_274);
or U86 (N_86,In_264,In_331);
nor U87 (N_87,In_395,In_148);
nand U88 (N_88,In_458,In_362);
nor U89 (N_89,In_182,In_77);
nand U90 (N_90,In_38,In_393);
nor U91 (N_91,In_308,In_170);
nand U92 (N_92,In_448,In_382);
nand U93 (N_93,In_258,In_222);
xnor U94 (N_94,In_152,In_234);
nor U95 (N_95,In_65,In_421);
or U96 (N_96,In_212,In_470);
and U97 (N_97,In_420,In_178);
nand U98 (N_98,In_47,In_489);
nor U99 (N_99,In_83,In_140);
or U100 (N_100,In_114,In_192);
nor U101 (N_101,In_338,In_11);
nand U102 (N_102,In_159,In_252);
nor U103 (N_103,In_334,In_141);
nand U104 (N_104,In_122,In_111);
xor U105 (N_105,In_241,In_69);
or U106 (N_106,In_68,In_377);
nor U107 (N_107,In_13,In_200);
and U108 (N_108,In_482,In_92);
nor U109 (N_109,In_406,In_328);
or U110 (N_110,In_317,In_127);
or U111 (N_111,In_440,In_460);
nand U112 (N_112,In_94,In_209);
nand U113 (N_113,In_39,In_118);
or U114 (N_114,In_478,In_217);
and U115 (N_115,In_446,In_157);
nand U116 (N_116,In_455,In_55);
or U117 (N_117,In_487,In_342);
and U118 (N_118,In_80,In_302);
nand U119 (N_119,In_82,In_42);
nor U120 (N_120,In_358,In_415);
or U121 (N_121,In_103,In_250);
and U122 (N_122,In_166,In_441);
and U123 (N_123,In_312,In_454);
nor U124 (N_124,In_131,In_57);
nor U125 (N_125,In_413,In_272);
nor U126 (N_126,In_235,In_105);
and U127 (N_127,In_228,In_402);
xnor U128 (N_128,In_86,In_230);
or U129 (N_129,In_194,In_70);
xor U130 (N_130,In_207,In_348);
and U131 (N_131,In_253,In_0);
nor U132 (N_132,In_468,In_18);
and U133 (N_133,In_430,In_387);
or U134 (N_134,In_459,In_189);
nand U135 (N_135,In_324,In_183);
and U136 (N_136,In_249,In_278);
and U137 (N_137,In_364,In_161);
and U138 (N_138,In_134,In_464);
nor U139 (N_139,In_451,In_232);
nand U140 (N_140,In_262,In_223);
nor U141 (N_141,In_474,In_101);
nor U142 (N_142,In_290,In_339);
or U143 (N_143,In_437,In_381);
or U144 (N_144,In_309,In_283);
xnor U145 (N_145,In_145,In_14);
nor U146 (N_146,In_34,In_88);
xnor U147 (N_147,In_495,In_240);
or U148 (N_148,In_273,In_30);
or U149 (N_149,In_355,In_445);
nand U150 (N_150,In_363,In_452);
nor U151 (N_151,In_282,In_497);
and U152 (N_152,In_475,In_171);
or U153 (N_153,In_476,In_129);
or U154 (N_154,In_195,In_74);
nor U155 (N_155,In_52,In_325);
nor U156 (N_156,In_266,In_438);
and U157 (N_157,In_227,In_81);
and U158 (N_158,In_167,In_184);
nor U159 (N_159,In_269,In_238);
nand U160 (N_160,In_20,In_66);
nor U161 (N_161,In_287,In_208);
and U162 (N_162,In_136,In_472);
nor U163 (N_163,In_25,In_248);
and U164 (N_164,In_97,In_423);
or U165 (N_165,In_193,In_279);
nor U166 (N_166,In_270,In_176);
nand U167 (N_167,In_31,In_410);
nor U168 (N_168,In_313,In_398);
xnor U169 (N_169,In_76,In_58);
or U170 (N_170,In_466,In_163);
nor U171 (N_171,In_211,In_359);
nand U172 (N_172,In_8,In_457);
xnor U173 (N_173,In_27,In_19);
and U174 (N_174,In_344,In_427);
and U175 (N_175,In_40,In_360);
or U176 (N_176,In_191,In_304);
and U177 (N_177,In_60,In_78);
and U178 (N_178,In_112,In_323);
nand U179 (N_179,In_299,In_345);
nor U180 (N_180,In_426,In_172);
or U181 (N_181,In_354,In_411);
nand U182 (N_182,In_346,In_62);
or U183 (N_183,In_394,In_412);
or U184 (N_184,In_46,In_386);
nand U185 (N_185,In_51,In_214);
or U186 (N_186,In_108,In_205);
nor U187 (N_187,In_295,In_419);
or U188 (N_188,In_491,In_116);
nand U189 (N_189,In_156,In_138);
nand U190 (N_190,In_291,In_494);
nor U191 (N_191,In_169,In_73);
nor U192 (N_192,In_165,In_267);
nand U193 (N_193,In_407,In_292);
nor U194 (N_194,In_133,In_284);
xor U195 (N_195,In_461,In_433);
nand U196 (N_196,In_400,In_321);
and U197 (N_197,In_99,In_261);
and U198 (N_198,In_341,In_380);
nor U199 (N_199,In_353,In_188);
or U200 (N_200,In_330,In_22);
or U201 (N_201,In_12,In_96);
nand U202 (N_202,In_179,In_177);
nand U203 (N_203,In_471,In_316);
nor U204 (N_204,In_85,In_391);
nand U205 (N_205,In_436,In_174);
nand U206 (N_206,In_6,In_265);
and U207 (N_207,In_37,In_21);
and U208 (N_208,In_16,In_15);
nand U209 (N_209,In_106,In_484);
and U210 (N_210,In_115,In_196);
or U211 (N_211,In_124,In_298);
nand U212 (N_212,In_243,In_367);
nor U213 (N_213,In_320,In_215);
nand U214 (N_214,In_374,In_372);
xor U215 (N_215,In_268,In_67);
or U216 (N_216,In_296,In_335);
nand U217 (N_217,In_225,In_297);
and U218 (N_218,In_350,In_162);
nor U219 (N_219,In_53,In_496);
nand U220 (N_220,In_314,In_190);
nand U221 (N_221,In_371,In_271);
and U222 (N_222,In_294,In_485);
nand U223 (N_223,In_206,In_4);
and U224 (N_224,In_473,In_48);
and U225 (N_225,In_59,In_50);
nor U226 (N_226,In_132,In_428);
nor U227 (N_227,In_462,In_143);
and U228 (N_228,In_378,In_322);
or U229 (N_229,In_498,In_185);
nor U230 (N_230,In_221,In_123);
nor U231 (N_231,In_397,In_424);
nor U232 (N_232,In_43,In_197);
xor U233 (N_233,In_246,In_449);
or U234 (N_234,In_488,In_239);
or U235 (N_235,In_26,In_146);
nor U236 (N_236,In_247,In_465);
or U237 (N_237,In_224,In_301);
and U238 (N_238,In_479,In_337);
and U239 (N_239,In_117,In_130);
nand U240 (N_240,In_229,In_405);
and U241 (N_241,In_310,In_396);
xnor U242 (N_242,In_244,In_263);
nand U243 (N_243,In_187,In_370);
nand U244 (N_244,In_376,In_220);
or U245 (N_245,In_87,In_109);
nor U246 (N_246,In_41,In_285);
and U247 (N_247,In_153,In_276);
nand U248 (N_248,In_357,In_49);
nor U249 (N_249,In_231,In_450);
nor U250 (N_250,In_86,In_334);
or U251 (N_251,In_444,In_237);
or U252 (N_252,In_95,In_64);
xor U253 (N_253,In_95,In_326);
or U254 (N_254,In_487,In_402);
and U255 (N_255,In_27,In_82);
nor U256 (N_256,In_34,In_347);
and U257 (N_257,In_389,In_171);
nor U258 (N_258,In_39,In_227);
and U259 (N_259,In_105,In_65);
nor U260 (N_260,In_228,In_435);
and U261 (N_261,In_410,In_387);
nor U262 (N_262,In_20,In_121);
nand U263 (N_263,In_266,In_322);
xor U264 (N_264,In_213,In_112);
nor U265 (N_265,In_252,In_220);
and U266 (N_266,In_293,In_384);
and U267 (N_267,In_103,In_138);
and U268 (N_268,In_224,In_83);
nor U269 (N_269,In_457,In_246);
or U270 (N_270,In_468,In_146);
nor U271 (N_271,In_4,In_172);
and U272 (N_272,In_55,In_436);
or U273 (N_273,In_495,In_142);
and U274 (N_274,In_447,In_45);
and U275 (N_275,In_118,In_461);
and U276 (N_276,In_72,In_496);
nand U277 (N_277,In_307,In_333);
and U278 (N_278,In_309,In_166);
or U279 (N_279,In_129,In_91);
or U280 (N_280,In_270,In_361);
nor U281 (N_281,In_169,In_313);
nand U282 (N_282,In_109,In_481);
nand U283 (N_283,In_55,In_334);
and U284 (N_284,In_259,In_297);
nor U285 (N_285,In_110,In_354);
and U286 (N_286,In_177,In_465);
and U287 (N_287,In_389,In_314);
xnor U288 (N_288,In_191,In_162);
nor U289 (N_289,In_211,In_394);
nand U290 (N_290,In_264,In_257);
nand U291 (N_291,In_370,In_242);
nor U292 (N_292,In_496,In_18);
nand U293 (N_293,In_314,In_331);
or U294 (N_294,In_414,In_429);
nor U295 (N_295,In_30,In_254);
nand U296 (N_296,In_22,In_420);
and U297 (N_297,In_436,In_406);
nand U298 (N_298,In_186,In_3);
and U299 (N_299,In_379,In_8);
nand U300 (N_300,In_164,In_67);
and U301 (N_301,In_114,In_50);
nand U302 (N_302,In_157,In_416);
nor U303 (N_303,In_207,In_29);
nand U304 (N_304,In_149,In_107);
nor U305 (N_305,In_95,In_41);
nor U306 (N_306,In_51,In_454);
nand U307 (N_307,In_202,In_75);
nand U308 (N_308,In_160,In_294);
and U309 (N_309,In_9,In_487);
xor U310 (N_310,In_89,In_337);
nor U311 (N_311,In_488,In_318);
nor U312 (N_312,In_370,In_492);
nor U313 (N_313,In_285,In_378);
and U314 (N_314,In_4,In_174);
and U315 (N_315,In_436,In_52);
or U316 (N_316,In_392,In_305);
xnor U317 (N_317,In_480,In_472);
or U318 (N_318,In_487,In_152);
nor U319 (N_319,In_38,In_101);
nand U320 (N_320,In_292,In_103);
nand U321 (N_321,In_314,In_400);
or U322 (N_322,In_48,In_232);
and U323 (N_323,In_326,In_277);
nand U324 (N_324,In_312,In_263);
or U325 (N_325,In_5,In_277);
nand U326 (N_326,In_414,In_87);
nor U327 (N_327,In_60,In_329);
nand U328 (N_328,In_491,In_218);
nor U329 (N_329,In_210,In_381);
and U330 (N_330,In_21,In_319);
or U331 (N_331,In_71,In_81);
nand U332 (N_332,In_318,In_174);
nand U333 (N_333,In_180,In_153);
or U334 (N_334,In_125,In_345);
nand U335 (N_335,In_337,In_243);
nand U336 (N_336,In_206,In_152);
xor U337 (N_337,In_473,In_319);
nand U338 (N_338,In_201,In_48);
and U339 (N_339,In_490,In_152);
or U340 (N_340,In_139,In_487);
and U341 (N_341,In_267,In_42);
and U342 (N_342,In_88,In_94);
xnor U343 (N_343,In_66,In_347);
xor U344 (N_344,In_218,In_307);
nor U345 (N_345,In_428,In_70);
or U346 (N_346,In_428,In_191);
and U347 (N_347,In_244,In_16);
nand U348 (N_348,In_115,In_492);
and U349 (N_349,In_209,In_450);
nand U350 (N_350,In_207,In_210);
and U351 (N_351,In_260,In_403);
or U352 (N_352,In_455,In_4);
and U353 (N_353,In_359,In_231);
or U354 (N_354,In_54,In_380);
or U355 (N_355,In_215,In_496);
and U356 (N_356,In_202,In_197);
nor U357 (N_357,In_299,In_467);
nor U358 (N_358,In_319,In_374);
or U359 (N_359,In_172,In_335);
xnor U360 (N_360,In_107,In_62);
nand U361 (N_361,In_288,In_351);
nor U362 (N_362,In_497,In_392);
xor U363 (N_363,In_438,In_35);
nor U364 (N_364,In_285,In_164);
and U365 (N_365,In_133,In_113);
and U366 (N_366,In_160,In_208);
nand U367 (N_367,In_418,In_224);
nand U368 (N_368,In_427,In_34);
nor U369 (N_369,In_151,In_314);
nor U370 (N_370,In_290,In_173);
or U371 (N_371,In_358,In_194);
or U372 (N_372,In_279,In_36);
or U373 (N_373,In_475,In_57);
nand U374 (N_374,In_20,In_95);
xor U375 (N_375,In_75,In_70);
nor U376 (N_376,In_437,In_324);
nor U377 (N_377,In_406,In_9);
nand U378 (N_378,In_218,In_323);
and U379 (N_379,In_357,In_37);
or U380 (N_380,In_118,In_1);
xnor U381 (N_381,In_290,In_325);
nand U382 (N_382,In_494,In_18);
or U383 (N_383,In_416,In_51);
nor U384 (N_384,In_269,In_329);
or U385 (N_385,In_102,In_22);
or U386 (N_386,In_426,In_57);
and U387 (N_387,In_1,In_88);
and U388 (N_388,In_131,In_109);
and U389 (N_389,In_169,In_250);
and U390 (N_390,In_346,In_270);
xnor U391 (N_391,In_448,In_440);
nor U392 (N_392,In_80,In_419);
and U393 (N_393,In_339,In_147);
or U394 (N_394,In_477,In_155);
nand U395 (N_395,In_323,In_125);
nand U396 (N_396,In_181,In_443);
or U397 (N_397,In_301,In_261);
or U398 (N_398,In_341,In_115);
or U399 (N_399,In_155,In_81);
and U400 (N_400,In_185,In_163);
nand U401 (N_401,In_10,In_183);
or U402 (N_402,In_168,In_211);
or U403 (N_403,In_162,In_416);
nor U404 (N_404,In_315,In_411);
nand U405 (N_405,In_493,In_385);
nand U406 (N_406,In_323,In_377);
and U407 (N_407,In_455,In_119);
nand U408 (N_408,In_369,In_14);
or U409 (N_409,In_132,In_452);
xnor U410 (N_410,In_262,In_458);
xnor U411 (N_411,In_351,In_67);
nor U412 (N_412,In_261,In_346);
or U413 (N_413,In_183,In_392);
xnor U414 (N_414,In_143,In_178);
or U415 (N_415,In_138,In_267);
or U416 (N_416,In_172,In_415);
nor U417 (N_417,In_410,In_416);
nand U418 (N_418,In_114,In_296);
and U419 (N_419,In_64,In_228);
xnor U420 (N_420,In_366,In_450);
nor U421 (N_421,In_207,In_447);
nand U422 (N_422,In_361,In_491);
and U423 (N_423,In_243,In_60);
or U424 (N_424,In_192,In_264);
nor U425 (N_425,In_146,In_406);
or U426 (N_426,In_260,In_75);
and U427 (N_427,In_201,In_342);
or U428 (N_428,In_292,In_249);
or U429 (N_429,In_324,In_406);
xnor U430 (N_430,In_115,In_439);
xor U431 (N_431,In_253,In_44);
nor U432 (N_432,In_412,In_298);
xor U433 (N_433,In_126,In_162);
nand U434 (N_434,In_488,In_191);
nor U435 (N_435,In_430,In_393);
nor U436 (N_436,In_306,In_479);
nor U437 (N_437,In_368,In_281);
and U438 (N_438,In_194,In_481);
or U439 (N_439,In_237,In_365);
nand U440 (N_440,In_457,In_113);
and U441 (N_441,In_429,In_300);
nand U442 (N_442,In_123,In_335);
nor U443 (N_443,In_280,In_104);
and U444 (N_444,In_281,In_16);
nand U445 (N_445,In_204,In_382);
nand U446 (N_446,In_227,In_354);
and U447 (N_447,In_84,In_463);
nand U448 (N_448,In_393,In_240);
or U449 (N_449,In_81,In_253);
nand U450 (N_450,In_219,In_181);
xor U451 (N_451,In_315,In_58);
nor U452 (N_452,In_249,In_304);
nor U453 (N_453,In_96,In_76);
nor U454 (N_454,In_388,In_31);
or U455 (N_455,In_296,In_412);
nand U456 (N_456,In_187,In_490);
or U457 (N_457,In_376,In_108);
or U458 (N_458,In_101,In_388);
and U459 (N_459,In_215,In_333);
and U460 (N_460,In_2,In_432);
or U461 (N_461,In_332,In_234);
nand U462 (N_462,In_284,In_492);
nor U463 (N_463,In_409,In_370);
or U464 (N_464,In_384,In_428);
xnor U465 (N_465,In_145,In_236);
and U466 (N_466,In_461,In_401);
and U467 (N_467,In_270,In_408);
nor U468 (N_468,In_361,In_477);
and U469 (N_469,In_70,In_102);
and U470 (N_470,In_179,In_24);
nand U471 (N_471,In_173,In_34);
xnor U472 (N_472,In_265,In_159);
and U473 (N_473,In_467,In_379);
and U474 (N_474,In_434,In_124);
nor U475 (N_475,In_485,In_471);
nor U476 (N_476,In_339,In_359);
nor U477 (N_477,In_281,In_62);
nand U478 (N_478,In_88,In_412);
and U479 (N_479,In_303,In_376);
or U480 (N_480,In_70,In_340);
xnor U481 (N_481,In_213,In_415);
nor U482 (N_482,In_452,In_494);
nand U483 (N_483,In_70,In_191);
nor U484 (N_484,In_227,In_344);
nor U485 (N_485,In_403,In_415);
or U486 (N_486,In_123,In_34);
xnor U487 (N_487,In_317,In_72);
nand U488 (N_488,In_46,In_112);
or U489 (N_489,In_450,In_354);
nor U490 (N_490,In_219,In_109);
nand U491 (N_491,In_150,In_309);
or U492 (N_492,In_351,In_264);
nor U493 (N_493,In_296,In_455);
nor U494 (N_494,In_392,In_211);
nand U495 (N_495,In_158,In_189);
nor U496 (N_496,In_293,In_196);
and U497 (N_497,In_87,In_225);
nor U498 (N_498,In_109,In_112);
and U499 (N_499,In_288,In_275);
and U500 (N_500,In_335,In_425);
nor U501 (N_501,In_431,In_372);
nand U502 (N_502,In_358,In_442);
nand U503 (N_503,In_445,In_26);
or U504 (N_504,In_40,In_318);
nor U505 (N_505,In_349,In_444);
or U506 (N_506,In_115,In_173);
and U507 (N_507,In_497,In_310);
nor U508 (N_508,In_164,In_237);
nand U509 (N_509,In_133,In_369);
nand U510 (N_510,In_345,In_471);
nor U511 (N_511,In_417,In_420);
nand U512 (N_512,In_58,In_416);
xor U513 (N_513,In_417,In_297);
and U514 (N_514,In_222,In_450);
xor U515 (N_515,In_34,In_305);
xnor U516 (N_516,In_127,In_65);
nand U517 (N_517,In_308,In_374);
nor U518 (N_518,In_273,In_336);
nand U519 (N_519,In_496,In_50);
and U520 (N_520,In_37,In_457);
and U521 (N_521,In_333,In_60);
nor U522 (N_522,In_461,In_264);
or U523 (N_523,In_286,In_389);
or U524 (N_524,In_340,In_250);
nor U525 (N_525,In_473,In_335);
or U526 (N_526,In_80,In_159);
nand U527 (N_527,In_146,In_262);
nand U528 (N_528,In_34,In_485);
nand U529 (N_529,In_190,In_105);
and U530 (N_530,In_29,In_153);
nor U531 (N_531,In_340,In_45);
nand U532 (N_532,In_86,In_13);
and U533 (N_533,In_337,In_493);
or U534 (N_534,In_391,In_243);
xor U535 (N_535,In_449,In_228);
nor U536 (N_536,In_110,In_258);
or U537 (N_537,In_399,In_247);
or U538 (N_538,In_467,In_291);
or U539 (N_539,In_94,In_224);
or U540 (N_540,In_86,In_229);
nand U541 (N_541,In_467,In_391);
xor U542 (N_542,In_53,In_123);
and U543 (N_543,In_360,In_119);
nand U544 (N_544,In_231,In_119);
or U545 (N_545,In_110,In_85);
or U546 (N_546,In_19,In_296);
or U547 (N_547,In_345,In_55);
nand U548 (N_548,In_497,In_383);
and U549 (N_549,In_459,In_287);
nand U550 (N_550,In_486,In_350);
nand U551 (N_551,In_3,In_155);
xor U552 (N_552,In_423,In_416);
and U553 (N_553,In_159,In_196);
and U554 (N_554,In_266,In_327);
nor U555 (N_555,In_195,In_332);
or U556 (N_556,In_385,In_496);
nand U557 (N_557,In_34,In_331);
or U558 (N_558,In_146,In_68);
or U559 (N_559,In_391,In_92);
and U560 (N_560,In_347,In_151);
and U561 (N_561,In_25,In_56);
and U562 (N_562,In_34,In_85);
nand U563 (N_563,In_479,In_459);
or U564 (N_564,In_247,In_98);
nor U565 (N_565,In_313,In_456);
and U566 (N_566,In_22,In_346);
xnor U567 (N_567,In_217,In_438);
or U568 (N_568,In_247,In_267);
nor U569 (N_569,In_442,In_51);
or U570 (N_570,In_378,In_149);
nor U571 (N_571,In_190,In_110);
or U572 (N_572,In_426,In_147);
or U573 (N_573,In_158,In_159);
and U574 (N_574,In_47,In_356);
nand U575 (N_575,In_306,In_55);
xnor U576 (N_576,In_122,In_345);
or U577 (N_577,In_93,In_331);
nor U578 (N_578,In_210,In_76);
or U579 (N_579,In_203,In_473);
nand U580 (N_580,In_383,In_352);
xor U581 (N_581,In_202,In_156);
nor U582 (N_582,In_36,In_39);
nand U583 (N_583,In_222,In_153);
and U584 (N_584,In_288,In_66);
or U585 (N_585,In_253,In_466);
and U586 (N_586,In_499,In_303);
nand U587 (N_587,In_256,In_76);
nor U588 (N_588,In_148,In_154);
and U589 (N_589,In_374,In_345);
nand U590 (N_590,In_395,In_47);
and U591 (N_591,In_47,In_87);
and U592 (N_592,In_36,In_416);
or U593 (N_593,In_471,In_342);
nor U594 (N_594,In_73,In_309);
xor U595 (N_595,In_51,In_397);
xor U596 (N_596,In_149,In_270);
nor U597 (N_597,In_457,In_145);
or U598 (N_598,In_138,In_85);
and U599 (N_599,In_67,In_97);
or U600 (N_600,In_304,In_362);
or U601 (N_601,In_331,In_15);
nor U602 (N_602,In_188,In_164);
or U603 (N_603,In_219,In_281);
nor U604 (N_604,In_261,In_297);
nor U605 (N_605,In_288,In_424);
nand U606 (N_606,In_458,In_181);
nor U607 (N_607,In_252,In_353);
nand U608 (N_608,In_208,In_49);
nand U609 (N_609,In_75,In_195);
and U610 (N_610,In_163,In_177);
nor U611 (N_611,In_271,In_351);
and U612 (N_612,In_358,In_418);
nor U613 (N_613,In_348,In_256);
nand U614 (N_614,In_416,In_385);
nor U615 (N_615,In_70,In_128);
nor U616 (N_616,In_25,In_231);
and U617 (N_617,In_444,In_318);
or U618 (N_618,In_288,In_269);
or U619 (N_619,In_274,In_169);
nand U620 (N_620,In_471,In_211);
or U621 (N_621,In_49,In_61);
nand U622 (N_622,In_325,In_6);
nand U623 (N_623,In_310,In_65);
nand U624 (N_624,In_225,In_157);
or U625 (N_625,In_300,In_434);
nand U626 (N_626,In_121,In_12);
and U627 (N_627,In_412,In_195);
and U628 (N_628,In_412,In_234);
and U629 (N_629,In_181,In_393);
or U630 (N_630,In_60,In_434);
nor U631 (N_631,In_4,In_419);
nor U632 (N_632,In_13,In_460);
or U633 (N_633,In_479,In_35);
nor U634 (N_634,In_487,In_39);
or U635 (N_635,In_372,In_159);
or U636 (N_636,In_57,In_471);
nand U637 (N_637,In_249,In_285);
or U638 (N_638,In_475,In_177);
or U639 (N_639,In_96,In_251);
nand U640 (N_640,In_312,In_289);
nor U641 (N_641,In_72,In_428);
and U642 (N_642,In_108,In_393);
nand U643 (N_643,In_419,In_252);
and U644 (N_644,In_299,In_165);
or U645 (N_645,In_480,In_386);
or U646 (N_646,In_347,In_495);
nand U647 (N_647,In_10,In_406);
nor U648 (N_648,In_205,In_236);
or U649 (N_649,In_363,In_461);
nand U650 (N_650,In_343,In_457);
nor U651 (N_651,In_350,In_85);
nor U652 (N_652,In_284,In_33);
and U653 (N_653,In_375,In_288);
nand U654 (N_654,In_388,In_108);
nor U655 (N_655,In_297,In_249);
nor U656 (N_656,In_415,In_341);
and U657 (N_657,In_80,In_319);
and U658 (N_658,In_393,In_312);
or U659 (N_659,In_301,In_186);
nor U660 (N_660,In_460,In_323);
and U661 (N_661,In_168,In_389);
and U662 (N_662,In_157,In_73);
xor U663 (N_663,In_416,In_224);
or U664 (N_664,In_92,In_274);
or U665 (N_665,In_124,In_478);
nand U666 (N_666,In_355,In_387);
or U667 (N_667,In_43,In_460);
or U668 (N_668,In_484,In_186);
nand U669 (N_669,In_253,In_378);
and U670 (N_670,In_46,In_325);
nor U671 (N_671,In_388,In_120);
nor U672 (N_672,In_137,In_289);
and U673 (N_673,In_452,In_311);
nor U674 (N_674,In_15,In_92);
nor U675 (N_675,In_339,In_22);
or U676 (N_676,In_138,In_289);
and U677 (N_677,In_49,In_77);
nor U678 (N_678,In_204,In_229);
nor U679 (N_679,In_323,In_452);
nor U680 (N_680,In_82,In_33);
and U681 (N_681,In_351,In_469);
or U682 (N_682,In_413,In_295);
nor U683 (N_683,In_428,In_381);
nand U684 (N_684,In_165,In_213);
nor U685 (N_685,In_141,In_266);
nand U686 (N_686,In_392,In_74);
or U687 (N_687,In_277,In_327);
and U688 (N_688,In_60,In_142);
and U689 (N_689,In_378,In_37);
or U690 (N_690,In_379,In_168);
nand U691 (N_691,In_377,In_3);
nand U692 (N_692,In_437,In_7);
nand U693 (N_693,In_34,In_96);
nand U694 (N_694,In_101,In_8);
nand U695 (N_695,In_429,In_412);
or U696 (N_696,In_238,In_361);
nand U697 (N_697,In_134,In_90);
nor U698 (N_698,In_478,In_6);
or U699 (N_699,In_89,In_355);
or U700 (N_700,In_79,In_88);
nand U701 (N_701,In_92,In_97);
and U702 (N_702,In_258,In_163);
nor U703 (N_703,In_231,In_272);
xnor U704 (N_704,In_123,In_78);
nor U705 (N_705,In_95,In_53);
or U706 (N_706,In_118,In_484);
and U707 (N_707,In_124,In_112);
and U708 (N_708,In_344,In_435);
and U709 (N_709,In_178,In_70);
nand U710 (N_710,In_3,In_306);
or U711 (N_711,In_231,In_293);
nand U712 (N_712,In_417,In_461);
and U713 (N_713,In_116,In_193);
or U714 (N_714,In_417,In_475);
xnor U715 (N_715,In_223,In_479);
nand U716 (N_716,In_497,In_95);
xnor U717 (N_717,In_482,In_190);
nand U718 (N_718,In_198,In_278);
nand U719 (N_719,In_320,In_495);
nor U720 (N_720,In_438,In_374);
xnor U721 (N_721,In_200,In_330);
xor U722 (N_722,In_293,In_307);
and U723 (N_723,In_25,In_341);
and U724 (N_724,In_405,In_45);
nor U725 (N_725,In_262,In_449);
nor U726 (N_726,In_343,In_393);
nand U727 (N_727,In_151,In_444);
nand U728 (N_728,In_138,In_428);
and U729 (N_729,In_315,In_316);
and U730 (N_730,In_429,In_111);
nor U731 (N_731,In_290,In_354);
nor U732 (N_732,In_21,In_325);
or U733 (N_733,In_480,In_129);
or U734 (N_734,In_162,In_106);
nor U735 (N_735,In_329,In_258);
and U736 (N_736,In_255,In_78);
and U737 (N_737,In_431,In_404);
or U738 (N_738,In_415,In_330);
or U739 (N_739,In_459,In_440);
nand U740 (N_740,In_101,In_331);
nand U741 (N_741,In_2,In_320);
or U742 (N_742,In_45,In_192);
or U743 (N_743,In_363,In_475);
xor U744 (N_744,In_191,In_435);
and U745 (N_745,In_139,In_288);
or U746 (N_746,In_143,In_314);
and U747 (N_747,In_299,In_346);
nand U748 (N_748,In_48,In_447);
nand U749 (N_749,In_259,In_221);
nor U750 (N_750,N_416,N_295);
or U751 (N_751,N_272,N_713);
or U752 (N_752,N_392,N_580);
or U753 (N_753,N_68,N_180);
xor U754 (N_754,N_323,N_253);
nor U755 (N_755,N_142,N_429);
nor U756 (N_756,N_625,N_89);
and U757 (N_757,N_308,N_641);
nor U758 (N_758,N_65,N_197);
xor U759 (N_759,N_606,N_656);
nand U760 (N_760,N_48,N_244);
nor U761 (N_761,N_524,N_27);
or U762 (N_762,N_186,N_124);
nand U763 (N_763,N_296,N_623);
xnor U764 (N_764,N_703,N_569);
or U765 (N_765,N_330,N_163);
or U766 (N_766,N_629,N_47);
nand U767 (N_767,N_727,N_368);
and U768 (N_768,N_565,N_329);
and U769 (N_769,N_73,N_218);
nand U770 (N_770,N_682,N_100);
nand U771 (N_771,N_592,N_523);
and U772 (N_772,N_684,N_185);
and U773 (N_773,N_744,N_120);
and U774 (N_774,N_571,N_126);
nand U775 (N_775,N_576,N_42);
xor U776 (N_776,N_254,N_635);
nand U777 (N_777,N_675,N_663);
and U778 (N_778,N_551,N_265);
or U779 (N_779,N_209,N_603);
xor U780 (N_780,N_644,N_566);
or U781 (N_781,N_262,N_154);
nand U782 (N_782,N_510,N_707);
nor U783 (N_783,N_619,N_282);
nand U784 (N_784,N_87,N_591);
nor U785 (N_785,N_438,N_494);
xor U786 (N_786,N_229,N_122);
and U787 (N_787,N_749,N_177);
and U788 (N_788,N_22,N_364);
xor U789 (N_789,N_354,N_711);
xor U790 (N_790,N_672,N_431);
and U791 (N_791,N_317,N_595);
nor U792 (N_792,N_237,N_650);
nor U793 (N_793,N_532,N_144);
nand U794 (N_794,N_320,N_586);
or U795 (N_795,N_506,N_715);
and U796 (N_796,N_730,N_655);
nand U797 (N_797,N_125,N_183);
nand U798 (N_798,N_609,N_171);
or U799 (N_799,N_721,N_134);
nand U800 (N_800,N_77,N_455);
and U801 (N_801,N_246,N_212);
xor U802 (N_802,N_653,N_222);
or U803 (N_803,N_688,N_502);
and U804 (N_804,N_678,N_473);
or U805 (N_805,N_101,N_350);
nand U806 (N_806,N_79,N_718);
nand U807 (N_807,N_556,N_182);
nor U808 (N_808,N_430,N_632);
xor U809 (N_809,N_129,N_234);
or U810 (N_810,N_80,N_121);
nand U811 (N_811,N_585,N_386);
nor U812 (N_812,N_643,N_271);
or U813 (N_813,N_467,N_661);
xnor U814 (N_814,N_173,N_321);
nor U815 (N_815,N_333,N_151);
and U816 (N_816,N_81,N_270);
and U817 (N_817,N_492,N_176);
nor U818 (N_818,N_489,N_337);
nor U819 (N_819,N_360,N_287);
nor U820 (N_820,N_362,N_40);
nand U821 (N_821,N_33,N_373);
and U822 (N_822,N_470,N_106);
or U823 (N_823,N_353,N_227);
nor U824 (N_824,N_136,N_102);
or U825 (N_825,N_252,N_664);
nor U826 (N_826,N_546,N_402);
nand U827 (N_827,N_164,N_657);
nor U828 (N_828,N_640,N_153);
nand U829 (N_829,N_704,N_54);
or U830 (N_830,N_335,N_50);
nor U831 (N_831,N_395,N_626);
or U832 (N_832,N_497,N_61);
nor U833 (N_833,N_389,N_2);
nand U834 (N_834,N_319,N_292);
nor U835 (N_835,N_526,N_639);
or U836 (N_836,N_515,N_114);
nor U837 (N_837,N_452,N_652);
nand U838 (N_838,N_456,N_277);
xnor U839 (N_839,N_450,N_605);
and U840 (N_840,N_117,N_486);
nor U841 (N_841,N_235,N_531);
nand U842 (N_842,N_279,N_55);
and U843 (N_843,N_720,N_132);
nand U844 (N_844,N_522,N_458);
nor U845 (N_845,N_299,N_712);
nand U846 (N_846,N_342,N_747);
nor U847 (N_847,N_554,N_341);
nand U848 (N_848,N_128,N_230);
nand U849 (N_849,N_516,N_67);
or U850 (N_850,N_505,N_683);
nand U851 (N_851,N_86,N_7);
nor U852 (N_852,N_401,N_9);
nand U853 (N_853,N_484,N_427);
and U854 (N_854,N_278,N_92);
nor U855 (N_855,N_268,N_705);
nor U856 (N_856,N_10,N_243);
and U857 (N_857,N_118,N_194);
and U858 (N_858,N_340,N_525);
and U859 (N_859,N_167,N_57);
nand U860 (N_860,N_159,N_20);
nand U861 (N_861,N_385,N_71);
and U862 (N_862,N_620,N_84);
nand U863 (N_863,N_220,N_138);
or U864 (N_864,N_95,N_674);
or U865 (N_865,N_618,N_491);
xnor U866 (N_866,N_318,N_155);
and U867 (N_867,N_109,N_303);
and U868 (N_868,N_196,N_555);
nor U869 (N_869,N_19,N_701);
or U870 (N_870,N_729,N_610);
nand U871 (N_871,N_593,N_740);
nor U872 (N_872,N_251,N_149);
or U873 (N_873,N_614,N_700);
and U874 (N_874,N_748,N_174);
or U875 (N_875,N_432,N_192);
and U876 (N_876,N_734,N_400);
nor U877 (N_877,N_130,N_725);
or U878 (N_878,N_150,N_290);
and U879 (N_879,N_348,N_607);
and U880 (N_880,N_665,N_170);
or U881 (N_881,N_410,N_509);
xnor U882 (N_882,N_44,N_372);
or U883 (N_883,N_451,N_504);
or U884 (N_884,N_582,N_152);
nand U885 (N_885,N_313,N_517);
and U886 (N_886,N_572,N_286);
nor U887 (N_887,N_293,N_168);
or U888 (N_888,N_557,N_13);
and U889 (N_889,N_460,N_544);
xnor U890 (N_890,N_6,N_594);
and U891 (N_891,N_443,N_453);
nor U892 (N_892,N_3,N_336);
and U893 (N_893,N_175,N_23);
nand U894 (N_894,N_558,N_375);
xor U895 (N_895,N_420,N_198);
nand U896 (N_896,N_83,N_181);
and U897 (N_897,N_219,N_387);
and U898 (N_898,N_600,N_288);
and U899 (N_899,N_37,N_399);
nor U900 (N_900,N_356,N_108);
xor U901 (N_901,N_534,N_216);
xnor U902 (N_902,N_724,N_241);
and U903 (N_903,N_719,N_30);
nand U904 (N_904,N_28,N_257);
nand U905 (N_905,N_221,N_217);
nor U906 (N_906,N_479,N_99);
nor U907 (N_907,N_634,N_331);
xor U908 (N_908,N_559,N_38);
nand U909 (N_909,N_223,N_503);
and U910 (N_910,N_698,N_111);
or U911 (N_911,N_371,N_611);
nand U912 (N_912,N_127,N_495);
nor U913 (N_913,N_511,N_56);
and U914 (N_914,N_596,N_8);
or U915 (N_915,N_36,N_103);
or U916 (N_916,N_158,N_107);
nor U917 (N_917,N_72,N_647);
xor U918 (N_918,N_298,N_357);
nor U919 (N_919,N_543,N_706);
or U920 (N_920,N_457,N_541);
and U921 (N_921,N_327,N_475);
and U922 (N_922,N_94,N_263);
xnor U923 (N_923,N_404,N_39);
nand U924 (N_924,N_325,N_147);
nand U925 (N_925,N_692,N_530);
nor U926 (N_926,N_538,N_97);
nor U927 (N_927,N_273,N_670);
nand U928 (N_928,N_419,N_463);
or U929 (N_929,N_225,N_428);
nand U930 (N_930,N_454,N_487);
and U931 (N_931,N_642,N_16);
xor U932 (N_932,N_143,N_542);
nand U933 (N_933,N_91,N_723);
or U934 (N_934,N_417,N_694);
or U935 (N_935,N_204,N_338);
xnor U936 (N_936,N_302,N_501);
nand U937 (N_937,N_393,N_74);
nor U938 (N_938,N_379,N_178);
nand U939 (N_939,N_165,N_85);
xnor U940 (N_940,N_137,N_179);
or U941 (N_941,N_628,N_745);
nor U942 (N_942,N_322,N_476);
nand U943 (N_943,N_344,N_666);
nand U944 (N_944,N_201,N_280);
nor U945 (N_945,N_306,N_14);
nor U946 (N_946,N_660,N_224);
or U947 (N_947,N_45,N_579);
nand U948 (N_948,N_662,N_345);
nand U949 (N_949,N_377,N_374);
nand U950 (N_950,N_518,N_633);
nor U951 (N_951,N_309,N_25);
nor U952 (N_952,N_722,N_60);
nor U953 (N_953,N_119,N_738);
nor U954 (N_954,N_112,N_513);
nor U955 (N_955,N_211,N_423);
and U956 (N_956,N_261,N_528);
and U957 (N_957,N_560,N_184);
xnor U958 (N_958,N_242,N_613);
and U959 (N_959,N_671,N_187);
nor U960 (N_960,N_285,N_17);
or U961 (N_961,N_267,N_247);
nor U962 (N_962,N_250,N_18);
nand U963 (N_963,N_587,N_638);
and U964 (N_964,N_471,N_203);
xnor U965 (N_965,N_365,N_407);
nand U966 (N_966,N_695,N_414);
nor U967 (N_967,N_157,N_195);
xor U968 (N_968,N_256,N_258);
nor U969 (N_969,N_366,N_381);
nand U970 (N_970,N_202,N_343);
and U971 (N_971,N_361,N_355);
xor U972 (N_972,N_169,N_376);
nand U973 (N_973,N_358,N_75);
and U974 (N_974,N_474,N_346);
or U975 (N_975,N_500,N_11);
or U976 (N_976,N_307,N_440);
and U977 (N_977,N_115,N_351);
xnor U978 (N_978,N_496,N_394);
or U979 (N_979,N_462,N_679);
xnor U980 (N_980,N_326,N_239);
nand U981 (N_981,N_104,N_477);
nor U982 (N_982,N_617,N_677);
nand U983 (N_983,N_301,N_686);
nand U984 (N_984,N_575,N_564);
nor U985 (N_985,N_110,N_434);
xnor U986 (N_986,N_76,N_697);
nand U987 (N_987,N_191,N_260);
or U988 (N_988,N_412,N_391);
and U989 (N_989,N_349,N_232);
or U990 (N_990,N_469,N_676);
nand U991 (N_991,N_1,N_214);
nand U992 (N_992,N_669,N_472);
nand U993 (N_993,N_478,N_736);
nor U994 (N_994,N_645,N_589);
and U995 (N_995,N_733,N_29);
nand U996 (N_996,N_161,N_411);
nand U997 (N_997,N_396,N_21);
and U998 (N_998,N_300,N_584);
and U999 (N_999,N_269,N_654);
nor U1000 (N_1000,N_378,N_590);
nor U1001 (N_1001,N_446,N_418);
nor U1002 (N_1002,N_339,N_562);
nand U1003 (N_1003,N_464,N_608);
and U1004 (N_1004,N_577,N_488);
or U1005 (N_1005,N_41,N_685);
nor U1006 (N_1006,N_305,N_384);
nand U1007 (N_1007,N_166,N_441);
or U1008 (N_1008,N_59,N_616);
xor U1009 (N_1009,N_390,N_537);
nor U1010 (N_1010,N_693,N_46);
nor U1011 (N_1011,N_284,N_708);
and U1012 (N_1012,N_622,N_570);
or U1013 (N_1013,N_78,N_567);
and U1014 (N_1014,N_190,N_597);
nand U1015 (N_1015,N_294,N_421);
or U1016 (N_1016,N_156,N_690);
nor U1017 (N_1017,N_648,N_631);
xnor U1018 (N_1018,N_742,N_200);
nand U1019 (N_1019,N_12,N_636);
xnor U1020 (N_1020,N_621,N_553);
and U1021 (N_1021,N_370,N_24);
and U1022 (N_1022,N_409,N_714);
nor U1023 (N_1023,N_249,N_383);
and U1024 (N_1024,N_449,N_498);
nor U1025 (N_1025,N_521,N_709);
or U1026 (N_1026,N_172,N_435);
nand U1027 (N_1027,N_297,N_627);
xor U1028 (N_1028,N_604,N_444);
nor U1029 (N_1029,N_405,N_550);
nand U1030 (N_1030,N_116,N_480);
and U1031 (N_1031,N_328,N_687);
xor U1032 (N_1032,N_739,N_535);
nand U1033 (N_1033,N_332,N_601);
nand U1034 (N_1034,N_208,N_439);
and U1035 (N_1035,N_248,N_728);
and U1036 (N_1036,N_26,N_447);
and U1037 (N_1037,N_508,N_746);
nor U1038 (N_1038,N_64,N_363);
or U1039 (N_1039,N_649,N_731);
and U1040 (N_1040,N_4,N_66);
or U1041 (N_1041,N_563,N_716);
and U1042 (N_1042,N_437,N_88);
nor U1043 (N_1043,N_90,N_651);
nor U1044 (N_1044,N_231,N_275);
and U1045 (N_1045,N_732,N_424);
or U1046 (N_1046,N_380,N_549);
nand U1047 (N_1047,N_316,N_304);
or U1048 (N_1048,N_481,N_70);
nor U1049 (N_1049,N_573,N_259);
and U1050 (N_1050,N_545,N_291);
or U1051 (N_1051,N_667,N_352);
nor U1052 (N_1052,N_255,N_445);
nor U1053 (N_1053,N_367,N_717);
xnor U1054 (N_1054,N_561,N_612);
nand U1055 (N_1055,N_459,N_615);
nand U1056 (N_1056,N_448,N_62);
nand U1057 (N_1057,N_637,N_512);
nor U1058 (N_1058,N_281,N_98);
or U1059 (N_1059,N_141,N_735);
or U1060 (N_1060,N_568,N_743);
and U1061 (N_1061,N_696,N_240);
nand U1062 (N_1062,N_283,N_426);
xor U1063 (N_1063,N_311,N_213);
nand U1064 (N_1064,N_574,N_624);
and U1065 (N_1065,N_160,N_468);
nor U1066 (N_1066,N_397,N_51);
or U1067 (N_1067,N_413,N_403);
xor U1068 (N_1068,N_483,N_215);
nand U1069 (N_1069,N_96,N_461);
and U1070 (N_1070,N_135,N_581);
and U1071 (N_1071,N_206,N_266);
xnor U1072 (N_1072,N_433,N_69);
nand U1073 (N_1073,N_442,N_536);
xnor U1074 (N_1074,N_578,N_369);
nor U1075 (N_1075,N_123,N_689);
or U1076 (N_1076,N_646,N_314);
nand U1077 (N_1077,N_245,N_359);
nor U1078 (N_1078,N_533,N_140);
nand U1079 (N_1079,N_507,N_547);
and U1080 (N_1080,N_312,N_43);
nand U1081 (N_1081,N_274,N_465);
nand U1082 (N_1082,N_31,N_737);
nand U1083 (N_1083,N_58,N_334);
and U1084 (N_1084,N_131,N_15);
xor U1085 (N_1085,N_113,N_5);
nand U1086 (N_1086,N_681,N_276);
or U1087 (N_1087,N_189,N_146);
and U1088 (N_1088,N_702,N_82);
and U1089 (N_1089,N_148,N_34);
xnor U1090 (N_1090,N_398,N_726);
nor U1091 (N_1091,N_205,N_588);
nand U1092 (N_1092,N_741,N_691);
nand U1093 (N_1093,N_53,N_539);
xor U1094 (N_1094,N_188,N_199);
nand U1095 (N_1095,N_347,N_552);
or U1096 (N_1096,N_408,N_210);
nor U1097 (N_1097,N_673,N_63);
nor U1098 (N_1098,N_529,N_49);
xor U1099 (N_1099,N_659,N_485);
or U1100 (N_1100,N_193,N_527);
nor U1101 (N_1101,N_236,N_583);
nor U1102 (N_1102,N_315,N_226);
or U1103 (N_1103,N_32,N_490);
or U1104 (N_1104,N_310,N_499);
and U1105 (N_1105,N_436,N_207);
xnor U1106 (N_1106,N_93,N_145);
or U1107 (N_1107,N_548,N_540);
and U1108 (N_1108,N_630,N_425);
nand U1109 (N_1109,N_599,N_264);
or U1110 (N_1110,N_0,N_710);
nor U1111 (N_1111,N_382,N_514);
and U1112 (N_1112,N_289,N_680);
or U1113 (N_1113,N_519,N_658);
or U1114 (N_1114,N_520,N_699);
and U1115 (N_1115,N_422,N_238);
nand U1116 (N_1116,N_602,N_233);
and U1117 (N_1117,N_139,N_388);
or U1118 (N_1118,N_52,N_162);
nor U1119 (N_1119,N_105,N_324);
nor U1120 (N_1120,N_133,N_406);
or U1121 (N_1121,N_482,N_228);
nor U1122 (N_1122,N_35,N_598);
nand U1123 (N_1123,N_493,N_668);
and U1124 (N_1124,N_466,N_415);
and U1125 (N_1125,N_97,N_436);
nor U1126 (N_1126,N_242,N_483);
nand U1127 (N_1127,N_730,N_299);
nand U1128 (N_1128,N_613,N_59);
or U1129 (N_1129,N_395,N_163);
or U1130 (N_1130,N_42,N_715);
and U1131 (N_1131,N_716,N_492);
or U1132 (N_1132,N_462,N_88);
nand U1133 (N_1133,N_722,N_502);
nand U1134 (N_1134,N_64,N_309);
or U1135 (N_1135,N_663,N_707);
or U1136 (N_1136,N_221,N_180);
nand U1137 (N_1137,N_55,N_624);
nor U1138 (N_1138,N_365,N_94);
nand U1139 (N_1139,N_360,N_77);
nor U1140 (N_1140,N_451,N_373);
and U1141 (N_1141,N_732,N_400);
and U1142 (N_1142,N_516,N_466);
nand U1143 (N_1143,N_681,N_493);
xnor U1144 (N_1144,N_683,N_153);
xor U1145 (N_1145,N_170,N_703);
or U1146 (N_1146,N_79,N_218);
nand U1147 (N_1147,N_37,N_76);
nand U1148 (N_1148,N_457,N_42);
xor U1149 (N_1149,N_597,N_137);
xnor U1150 (N_1150,N_514,N_345);
or U1151 (N_1151,N_146,N_303);
xnor U1152 (N_1152,N_90,N_344);
nand U1153 (N_1153,N_640,N_536);
and U1154 (N_1154,N_386,N_138);
or U1155 (N_1155,N_195,N_380);
nor U1156 (N_1156,N_255,N_358);
or U1157 (N_1157,N_593,N_79);
nor U1158 (N_1158,N_189,N_465);
xnor U1159 (N_1159,N_99,N_241);
and U1160 (N_1160,N_440,N_703);
or U1161 (N_1161,N_164,N_707);
and U1162 (N_1162,N_150,N_254);
xnor U1163 (N_1163,N_339,N_705);
or U1164 (N_1164,N_475,N_59);
or U1165 (N_1165,N_571,N_397);
or U1166 (N_1166,N_591,N_510);
and U1167 (N_1167,N_665,N_630);
nor U1168 (N_1168,N_288,N_464);
xor U1169 (N_1169,N_118,N_110);
or U1170 (N_1170,N_669,N_150);
nand U1171 (N_1171,N_10,N_409);
or U1172 (N_1172,N_690,N_279);
nand U1173 (N_1173,N_676,N_478);
xnor U1174 (N_1174,N_587,N_378);
xnor U1175 (N_1175,N_317,N_296);
nor U1176 (N_1176,N_77,N_636);
or U1177 (N_1177,N_4,N_363);
nor U1178 (N_1178,N_440,N_578);
nand U1179 (N_1179,N_83,N_197);
and U1180 (N_1180,N_493,N_410);
nor U1181 (N_1181,N_194,N_541);
nand U1182 (N_1182,N_82,N_610);
and U1183 (N_1183,N_322,N_495);
xor U1184 (N_1184,N_192,N_288);
and U1185 (N_1185,N_413,N_224);
or U1186 (N_1186,N_43,N_449);
nor U1187 (N_1187,N_534,N_614);
or U1188 (N_1188,N_104,N_119);
and U1189 (N_1189,N_313,N_426);
nand U1190 (N_1190,N_199,N_343);
or U1191 (N_1191,N_495,N_340);
and U1192 (N_1192,N_574,N_399);
nand U1193 (N_1193,N_299,N_48);
nor U1194 (N_1194,N_481,N_578);
and U1195 (N_1195,N_577,N_525);
or U1196 (N_1196,N_99,N_585);
or U1197 (N_1197,N_174,N_444);
nor U1198 (N_1198,N_72,N_86);
and U1199 (N_1199,N_376,N_52);
and U1200 (N_1200,N_467,N_689);
nand U1201 (N_1201,N_452,N_115);
nor U1202 (N_1202,N_261,N_15);
and U1203 (N_1203,N_526,N_252);
and U1204 (N_1204,N_344,N_149);
or U1205 (N_1205,N_528,N_232);
nand U1206 (N_1206,N_685,N_559);
or U1207 (N_1207,N_344,N_631);
or U1208 (N_1208,N_27,N_467);
or U1209 (N_1209,N_659,N_524);
xnor U1210 (N_1210,N_289,N_301);
and U1211 (N_1211,N_259,N_381);
and U1212 (N_1212,N_260,N_703);
xnor U1213 (N_1213,N_402,N_383);
nand U1214 (N_1214,N_570,N_35);
and U1215 (N_1215,N_365,N_156);
nor U1216 (N_1216,N_516,N_457);
and U1217 (N_1217,N_168,N_476);
nor U1218 (N_1218,N_444,N_265);
xnor U1219 (N_1219,N_690,N_596);
nand U1220 (N_1220,N_670,N_253);
nor U1221 (N_1221,N_547,N_212);
nor U1222 (N_1222,N_607,N_728);
or U1223 (N_1223,N_316,N_113);
and U1224 (N_1224,N_711,N_609);
or U1225 (N_1225,N_243,N_603);
and U1226 (N_1226,N_474,N_235);
nor U1227 (N_1227,N_478,N_617);
nor U1228 (N_1228,N_72,N_137);
or U1229 (N_1229,N_246,N_606);
or U1230 (N_1230,N_397,N_7);
or U1231 (N_1231,N_299,N_427);
and U1232 (N_1232,N_738,N_344);
and U1233 (N_1233,N_471,N_455);
and U1234 (N_1234,N_151,N_730);
nor U1235 (N_1235,N_212,N_46);
xor U1236 (N_1236,N_222,N_380);
nor U1237 (N_1237,N_547,N_520);
and U1238 (N_1238,N_555,N_475);
and U1239 (N_1239,N_274,N_649);
or U1240 (N_1240,N_431,N_675);
nand U1241 (N_1241,N_488,N_417);
nand U1242 (N_1242,N_739,N_307);
nor U1243 (N_1243,N_401,N_639);
nor U1244 (N_1244,N_716,N_109);
and U1245 (N_1245,N_602,N_415);
and U1246 (N_1246,N_273,N_356);
and U1247 (N_1247,N_447,N_200);
or U1248 (N_1248,N_713,N_494);
or U1249 (N_1249,N_261,N_653);
nor U1250 (N_1250,N_565,N_348);
or U1251 (N_1251,N_275,N_615);
xnor U1252 (N_1252,N_621,N_69);
nor U1253 (N_1253,N_108,N_546);
nor U1254 (N_1254,N_665,N_699);
nand U1255 (N_1255,N_332,N_207);
or U1256 (N_1256,N_708,N_133);
or U1257 (N_1257,N_384,N_258);
nand U1258 (N_1258,N_2,N_675);
nor U1259 (N_1259,N_732,N_14);
xnor U1260 (N_1260,N_3,N_548);
and U1261 (N_1261,N_639,N_678);
nor U1262 (N_1262,N_457,N_259);
nand U1263 (N_1263,N_400,N_407);
nand U1264 (N_1264,N_597,N_293);
and U1265 (N_1265,N_507,N_655);
nor U1266 (N_1266,N_13,N_14);
nand U1267 (N_1267,N_287,N_682);
or U1268 (N_1268,N_322,N_178);
xnor U1269 (N_1269,N_126,N_166);
nor U1270 (N_1270,N_250,N_210);
nor U1271 (N_1271,N_21,N_557);
or U1272 (N_1272,N_722,N_439);
nand U1273 (N_1273,N_362,N_505);
or U1274 (N_1274,N_511,N_93);
or U1275 (N_1275,N_59,N_117);
nor U1276 (N_1276,N_313,N_370);
and U1277 (N_1277,N_276,N_136);
or U1278 (N_1278,N_479,N_55);
nor U1279 (N_1279,N_103,N_14);
or U1280 (N_1280,N_327,N_468);
xnor U1281 (N_1281,N_323,N_60);
and U1282 (N_1282,N_20,N_3);
and U1283 (N_1283,N_20,N_396);
and U1284 (N_1284,N_594,N_615);
or U1285 (N_1285,N_111,N_63);
or U1286 (N_1286,N_505,N_330);
xnor U1287 (N_1287,N_434,N_385);
nor U1288 (N_1288,N_517,N_476);
or U1289 (N_1289,N_17,N_731);
nand U1290 (N_1290,N_688,N_587);
nor U1291 (N_1291,N_342,N_746);
or U1292 (N_1292,N_688,N_147);
nand U1293 (N_1293,N_59,N_205);
and U1294 (N_1294,N_441,N_97);
nor U1295 (N_1295,N_542,N_671);
nor U1296 (N_1296,N_728,N_188);
nor U1297 (N_1297,N_535,N_351);
nand U1298 (N_1298,N_431,N_267);
or U1299 (N_1299,N_650,N_304);
and U1300 (N_1300,N_595,N_44);
nand U1301 (N_1301,N_587,N_692);
nor U1302 (N_1302,N_121,N_497);
nor U1303 (N_1303,N_147,N_53);
nor U1304 (N_1304,N_126,N_492);
and U1305 (N_1305,N_210,N_707);
nand U1306 (N_1306,N_331,N_580);
xor U1307 (N_1307,N_598,N_547);
nor U1308 (N_1308,N_566,N_201);
and U1309 (N_1309,N_595,N_33);
or U1310 (N_1310,N_630,N_520);
or U1311 (N_1311,N_364,N_291);
nor U1312 (N_1312,N_10,N_39);
nor U1313 (N_1313,N_161,N_572);
nor U1314 (N_1314,N_45,N_124);
and U1315 (N_1315,N_603,N_589);
nand U1316 (N_1316,N_154,N_617);
xnor U1317 (N_1317,N_560,N_411);
and U1318 (N_1318,N_442,N_712);
nor U1319 (N_1319,N_416,N_9);
nand U1320 (N_1320,N_624,N_70);
nor U1321 (N_1321,N_527,N_729);
and U1322 (N_1322,N_225,N_183);
nor U1323 (N_1323,N_551,N_427);
xnor U1324 (N_1324,N_562,N_397);
or U1325 (N_1325,N_357,N_339);
nand U1326 (N_1326,N_60,N_120);
nand U1327 (N_1327,N_85,N_576);
and U1328 (N_1328,N_669,N_592);
and U1329 (N_1329,N_6,N_73);
nor U1330 (N_1330,N_1,N_53);
or U1331 (N_1331,N_330,N_22);
or U1332 (N_1332,N_730,N_304);
nand U1333 (N_1333,N_309,N_459);
xor U1334 (N_1334,N_182,N_207);
nand U1335 (N_1335,N_724,N_501);
nand U1336 (N_1336,N_692,N_152);
and U1337 (N_1337,N_542,N_249);
nand U1338 (N_1338,N_467,N_91);
nand U1339 (N_1339,N_351,N_212);
and U1340 (N_1340,N_328,N_14);
nand U1341 (N_1341,N_519,N_364);
and U1342 (N_1342,N_643,N_374);
xor U1343 (N_1343,N_657,N_371);
nor U1344 (N_1344,N_651,N_443);
and U1345 (N_1345,N_490,N_96);
and U1346 (N_1346,N_71,N_187);
or U1347 (N_1347,N_431,N_101);
and U1348 (N_1348,N_610,N_108);
and U1349 (N_1349,N_134,N_425);
nand U1350 (N_1350,N_477,N_375);
or U1351 (N_1351,N_329,N_697);
nor U1352 (N_1352,N_749,N_94);
and U1353 (N_1353,N_265,N_419);
nor U1354 (N_1354,N_551,N_516);
or U1355 (N_1355,N_166,N_542);
or U1356 (N_1356,N_109,N_188);
nand U1357 (N_1357,N_357,N_378);
nand U1358 (N_1358,N_586,N_254);
nand U1359 (N_1359,N_182,N_269);
and U1360 (N_1360,N_318,N_502);
nand U1361 (N_1361,N_735,N_292);
and U1362 (N_1362,N_389,N_171);
nand U1363 (N_1363,N_232,N_106);
and U1364 (N_1364,N_741,N_635);
and U1365 (N_1365,N_155,N_530);
nor U1366 (N_1366,N_457,N_696);
nand U1367 (N_1367,N_713,N_281);
or U1368 (N_1368,N_254,N_147);
nand U1369 (N_1369,N_632,N_440);
and U1370 (N_1370,N_621,N_177);
nand U1371 (N_1371,N_674,N_225);
nor U1372 (N_1372,N_86,N_81);
nand U1373 (N_1373,N_31,N_599);
nor U1374 (N_1374,N_719,N_143);
nand U1375 (N_1375,N_323,N_466);
or U1376 (N_1376,N_496,N_536);
and U1377 (N_1377,N_602,N_472);
nor U1378 (N_1378,N_657,N_544);
or U1379 (N_1379,N_138,N_389);
and U1380 (N_1380,N_281,N_316);
nor U1381 (N_1381,N_541,N_603);
nor U1382 (N_1382,N_527,N_622);
nor U1383 (N_1383,N_555,N_46);
or U1384 (N_1384,N_252,N_644);
or U1385 (N_1385,N_588,N_687);
xnor U1386 (N_1386,N_709,N_347);
or U1387 (N_1387,N_500,N_663);
and U1388 (N_1388,N_219,N_92);
and U1389 (N_1389,N_684,N_294);
and U1390 (N_1390,N_303,N_524);
or U1391 (N_1391,N_637,N_618);
and U1392 (N_1392,N_180,N_187);
or U1393 (N_1393,N_411,N_198);
xnor U1394 (N_1394,N_336,N_400);
and U1395 (N_1395,N_566,N_592);
and U1396 (N_1396,N_168,N_61);
xor U1397 (N_1397,N_535,N_466);
nand U1398 (N_1398,N_305,N_548);
and U1399 (N_1399,N_624,N_686);
and U1400 (N_1400,N_70,N_306);
and U1401 (N_1401,N_14,N_542);
and U1402 (N_1402,N_405,N_474);
nor U1403 (N_1403,N_630,N_80);
and U1404 (N_1404,N_335,N_23);
or U1405 (N_1405,N_293,N_620);
nor U1406 (N_1406,N_364,N_92);
nand U1407 (N_1407,N_566,N_728);
or U1408 (N_1408,N_567,N_70);
and U1409 (N_1409,N_333,N_174);
and U1410 (N_1410,N_296,N_430);
nand U1411 (N_1411,N_548,N_640);
nand U1412 (N_1412,N_126,N_81);
and U1413 (N_1413,N_279,N_700);
nor U1414 (N_1414,N_705,N_744);
and U1415 (N_1415,N_705,N_299);
nor U1416 (N_1416,N_426,N_504);
and U1417 (N_1417,N_635,N_491);
nand U1418 (N_1418,N_387,N_479);
xor U1419 (N_1419,N_276,N_493);
or U1420 (N_1420,N_708,N_600);
or U1421 (N_1421,N_178,N_563);
nor U1422 (N_1422,N_503,N_175);
and U1423 (N_1423,N_626,N_131);
or U1424 (N_1424,N_85,N_683);
or U1425 (N_1425,N_82,N_388);
nor U1426 (N_1426,N_361,N_265);
nor U1427 (N_1427,N_19,N_78);
and U1428 (N_1428,N_140,N_218);
or U1429 (N_1429,N_365,N_2);
and U1430 (N_1430,N_497,N_708);
or U1431 (N_1431,N_40,N_648);
nor U1432 (N_1432,N_308,N_27);
and U1433 (N_1433,N_629,N_539);
and U1434 (N_1434,N_57,N_295);
nor U1435 (N_1435,N_469,N_206);
nand U1436 (N_1436,N_229,N_495);
nor U1437 (N_1437,N_669,N_734);
nand U1438 (N_1438,N_705,N_276);
nor U1439 (N_1439,N_657,N_411);
nor U1440 (N_1440,N_470,N_717);
or U1441 (N_1441,N_576,N_692);
xor U1442 (N_1442,N_497,N_113);
nor U1443 (N_1443,N_312,N_495);
or U1444 (N_1444,N_556,N_392);
and U1445 (N_1445,N_585,N_358);
nand U1446 (N_1446,N_130,N_459);
or U1447 (N_1447,N_128,N_651);
and U1448 (N_1448,N_716,N_259);
or U1449 (N_1449,N_32,N_148);
or U1450 (N_1450,N_661,N_17);
and U1451 (N_1451,N_22,N_683);
nand U1452 (N_1452,N_337,N_156);
nand U1453 (N_1453,N_6,N_334);
and U1454 (N_1454,N_372,N_82);
nand U1455 (N_1455,N_375,N_738);
and U1456 (N_1456,N_227,N_633);
nand U1457 (N_1457,N_447,N_105);
nand U1458 (N_1458,N_462,N_307);
xnor U1459 (N_1459,N_105,N_581);
xnor U1460 (N_1460,N_252,N_500);
nor U1461 (N_1461,N_358,N_389);
nor U1462 (N_1462,N_157,N_97);
nor U1463 (N_1463,N_338,N_343);
or U1464 (N_1464,N_164,N_554);
and U1465 (N_1465,N_105,N_234);
xnor U1466 (N_1466,N_137,N_432);
nand U1467 (N_1467,N_672,N_283);
or U1468 (N_1468,N_30,N_66);
or U1469 (N_1469,N_172,N_430);
nand U1470 (N_1470,N_234,N_374);
or U1471 (N_1471,N_572,N_442);
nor U1472 (N_1472,N_349,N_431);
or U1473 (N_1473,N_29,N_98);
nand U1474 (N_1474,N_672,N_645);
and U1475 (N_1475,N_331,N_153);
and U1476 (N_1476,N_416,N_187);
and U1477 (N_1477,N_568,N_46);
nand U1478 (N_1478,N_724,N_77);
nand U1479 (N_1479,N_567,N_648);
nor U1480 (N_1480,N_351,N_338);
xnor U1481 (N_1481,N_487,N_23);
nor U1482 (N_1482,N_190,N_169);
nand U1483 (N_1483,N_349,N_438);
nor U1484 (N_1484,N_297,N_522);
nand U1485 (N_1485,N_469,N_746);
nand U1486 (N_1486,N_13,N_389);
and U1487 (N_1487,N_506,N_31);
nand U1488 (N_1488,N_52,N_293);
or U1489 (N_1489,N_480,N_6);
nand U1490 (N_1490,N_493,N_375);
and U1491 (N_1491,N_112,N_651);
and U1492 (N_1492,N_603,N_705);
or U1493 (N_1493,N_387,N_128);
or U1494 (N_1494,N_260,N_333);
nand U1495 (N_1495,N_196,N_598);
nand U1496 (N_1496,N_107,N_160);
xnor U1497 (N_1497,N_432,N_280);
and U1498 (N_1498,N_476,N_224);
or U1499 (N_1499,N_408,N_549);
nor U1500 (N_1500,N_791,N_951);
nand U1501 (N_1501,N_811,N_877);
nand U1502 (N_1502,N_800,N_1378);
and U1503 (N_1503,N_1053,N_1266);
nand U1504 (N_1504,N_1223,N_1387);
nor U1505 (N_1505,N_1030,N_1054);
nor U1506 (N_1506,N_1166,N_850);
and U1507 (N_1507,N_1471,N_1091);
nand U1508 (N_1508,N_1434,N_1465);
nand U1509 (N_1509,N_944,N_1422);
and U1510 (N_1510,N_1095,N_873);
and U1511 (N_1511,N_1086,N_943);
xnor U1512 (N_1512,N_855,N_1288);
nor U1513 (N_1513,N_1483,N_1025);
and U1514 (N_1514,N_1308,N_1048);
nand U1515 (N_1515,N_960,N_1273);
nor U1516 (N_1516,N_1195,N_1251);
nor U1517 (N_1517,N_1010,N_1219);
nor U1518 (N_1518,N_1292,N_756);
nand U1519 (N_1519,N_1477,N_817);
nand U1520 (N_1520,N_1404,N_952);
and U1521 (N_1521,N_1302,N_1311);
nand U1522 (N_1522,N_1147,N_1359);
nor U1523 (N_1523,N_1338,N_1112);
nand U1524 (N_1524,N_1263,N_1397);
and U1525 (N_1525,N_782,N_985);
nor U1526 (N_1526,N_1021,N_1486);
or U1527 (N_1527,N_1320,N_1394);
or U1528 (N_1528,N_789,N_934);
nor U1529 (N_1529,N_939,N_1040);
xnor U1530 (N_1530,N_1125,N_1447);
nor U1531 (N_1531,N_771,N_1383);
xnor U1532 (N_1532,N_1200,N_786);
xor U1533 (N_1533,N_843,N_916);
and U1534 (N_1534,N_762,N_757);
xor U1535 (N_1535,N_930,N_1305);
and U1536 (N_1536,N_1293,N_793);
or U1537 (N_1537,N_1360,N_968);
and U1538 (N_1538,N_1051,N_864);
and U1539 (N_1539,N_941,N_976);
or U1540 (N_1540,N_1304,N_912);
xor U1541 (N_1541,N_888,N_1106);
or U1542 (N_1542,N_1371,N_1395);
nor U1543 (N_1543,N_809,N_846);
or U1544 (N_1544,N_1159,N_1211);
or U1545 (N_1545,N_1313,N_1415);
nor U1546 (N_1546,N_1409,N_1068);
and U1547 (N_1547,N_928,N_766);
xor U1548 (N_1548,N_1228,N_1358);
and U1549 (N_1549,N_796,N_1233);
and U1550 (N_1550,N_1188,N_1489);
nor U1551 (N_1551,N_1274,N_1231);
and U1552 (N_1552,N_1396,N_931);
nor U1553 (N_1553,N_1022,N_977);
and U1554 (N_1554,N_967,N_1303);
nor U1555 (N_1555,N_1239,N_848);
or U1556 (N_1556,N_849,N_1144);
nor U1557 (N_1557,N_1083,N_1016);
and U1558 (N_1558,N_1492,N_1407);
and U1559 (N_1559,N_1101,N_798);
or U1560 (N_1560,N_1041,N_1122);
nand U1561 (N_1561,N_1301,N_966);
or U1562 (N_1562,N_1045,N_1330);
or U1563 (N_1563,N_1150,N_1449);
and U1564 (N_1564,N_797,N_1000);
nor U1565 (N_1565,N_831,N_1009);
nand U1566 (N_1566,N_1116,N_1232);
nor U1567 (N_1567,N_1493,N_1044);
nor U1568 (N_1568,N_1463,N_993);
or U1569 (N_1569,N_1425,N_1323);
or U1570 (N_1570,N_1210,N_1250);
xor U1571 (N_1571,N_1270,N_1204);
nor U1572 (N_1572,N_1340,N_980);
nand U1573 (N_1573,N_962,N_861);
and U1574 (N_1574,N_955,N_1280);
and U1575 (N_1575,N_1442,N_1451);
nand U1576 (N_1576,N_1017,N_973);
nand U1577 (N_1577,N_1361,N_946);
or U1578 (N_1578,N_874,N_1355);
nor U1579 (N_1579,N_1418,N_1061);
and U1580 (N_1580,N_788,N_1373);
nand U1581 (N_1581,N_1152,N_910);
or U1582 (N_1582,N_1163,N_988);
nand U1583 (N_1583,N_872,N_1376);
nor U1584 (N_1584,N_1324,N_999);
nor U1585 (N_1585,N_979,N_1278);
xor U1586 (N_1586,N_914,N_1470);
or U1587 (N_1587,N_1146,N_965);
nor U1588 (N_1588,N_1084,N_1128);
and U1589 (N_1589,N_957,N_1184);
and U1590 (N_1590,N_866,N_1007);
nand U1591 (N_1591,N_1328,N_1435);
or U1592 (N_1592,N_913,N_1149);
nor U1593 (N_1593,N_984,N_1120);
nand U1594 (N_1594,N_1473,N_1260);
and U1595 (N_1595,N_936,N_1236);
or U1596 (N_1596,N_1458,N_1291);
or U1597 (N_1597,N_1105,N_803);
xnor U1598 (N_1598,N_1336,N_1464);
xor U1599 (N_1599,N_1490,N_1129);
nand U1600 (N_1600,N_1286,N_1310);
and U1601 (N_1601,N_1244,N_1156);
and U1602 (N_1602,N_1108,N_1354);
and U1603 (N_1603,N_1230,N_915);
nor U1604 (N_1604,N_1472,N_1158);
nand U1605 (N_1605,N_869,N_812);
or U1606 (N_1606,N_1182,N_1193);
xnor U1607 (N_1607,N_1454,N_1093);
nor U1608 (N_1608,N_1450,N_1332);
nand U1609 (N_1609,N_1057,N_1367);
and U1610 (N_1610,N_1365,N_1065);
and U1611 (N_1611,N_1099,N_1480);
nor U1612 (N_1612,N_1078,N_862);
and U1613 (N_1613,N_768,N_1300);
nor U1614 (N_1614,N_751,N_1350);
and U1615 (N_1615,N_838,N_794);
or U1616 (N_1616,N_958,N_1240);
nor U1617 (N_1617,N_863,N_895);
nor U1618 (N_1618,N_876,N_1269);
nor U1619 (N_1619,N_1491,N_1107);
nor U1620 (N_1620,N_887,N_1306);
nor U1621 (N_1621,N_975,N_1036);
xor U1622 (N_1622,N_889,N_1011);
nand U1623 (N_1623,N_1123,N_778);
and U1624 (N_1624,N_1117,N_1056);
and U1625 (N_1625,N_1275,N_1202);
nand U1626 (N_1626,N_1374,N_1111);
nor U1627 (N_1627,N_1089,N_902);
or U1628 (N_1628,N_1467,N_1224);
nand U1629 (N_1629,N_818,N_1218);
nand U1630 (N_1630,N_1460,N_1178);
nor U1631 (N_1631,N_1499,N_1031);
or U1632 (N_1632,N_1322,N_1419);
nor U1633 (N_1633,N_1189,N_1100);
or U1634 (N_1634,N_1001,N_1443);
nor U1635 (N_1635,N_1047,N_901);
or U1636 (N_1636,N_938,N_1353);
and U1637 (N_1637,N_1148,N_1438);
or U1638 (N_1638,N_1271,N_1253);
xor U1639 (N_1639,N_758,N_1363);
and U1640 (N_1640,N_997,N_808);
nand U1641 (N_1641,N_1186,N_1176);
nor U1642 (N_1642,N_926,N_1227);
nand U1643 (N_1643,N_1416,N_814);
xor U1644 (N_1644,N_1135,N_1071);
nor U1645 (N_1645,N_1362,N_1282);
xnor U1646 (N_1646,N_774,N_1364);
or U1647 (N_1647,N_1173,N_883);
or U1648 (N_1648,N_959,N_1343);
nand U1649 (N_1649,N_1018,N_1073);
nor U1650 (N_1650,N_1055,N_920);
and U1651 (N_1651,N_1479,N_1385);
and U1652 (N_1652,N_1319,N_1254);
or U1653 (N_1653,N_1075,N_1154);
xnor U1654 (N_1654,N_1206,N_835);
or U1655 (N_1655,N_799,N_1238);
or U1656 (N_1656,N_911,N_1290);
nor U1657 (N_1657,N_1118,N_1297);
nand U1658 (N_1658,N_1208,N_1437);
and U1659 (N_1659,N_945,N_853);
nand U1660 (N_1660,N_1344,N_1008);
nand U1661 (N_1661,N_1137,N_1015);
or U1662 (N_1662,N_998,N_776);
or U1663 (N_1663,N_825,N_1279);
xnor U1664 (N_1664,N_903,N_919);
or U1665 (N_1665,N_1205,N_969);
xnor U1666 (N_1666,N_1058,N_1348);
and U1667 (N_1667,N_832,N_1431);
and U1668 (N_1668,N_1289,N_907);
or U1669 (N_1669,N_1424,N_1352);
xor U1670 (N_1670,N_868,N_1023);
or U1671 (N_1671,N_1172,N_1393);
nand U1672 (N_1672,N_805,N_859);
nand U1673 (N_1673,N_1453,N_1430);
and U1674 (N_1674,N_819,N_1029);
and U1675 (N_1675,N_1398,N_1180);
nand U1676 (N_1676,N_1098,N_1375);
xnor U1677 (N_1677,N_840,N_1427);
nand U1678 (N_1678,N_767,N_1142);
nor U1679 (N_1679,N_1377,N_1024);
nor U1680 (N_1680,N_1114,N_765);
nand U1681 (N_1681,N_1062,N_896);
and U1682 (N_1682,N_1124,N_1247);
nor U1683 (N_1683,N_1222,N_1235);
nor U1684 (N_1684,N_1405,N_956);
and U1685 (N_1685,N_1441,N_1080);
and U1686 (N_1686,N_1256,N_856);
nand U1687 (N_1687,N_1487,N_801);
or U1688 (N_1688,N_898,N_1496);
xor U1689 (N_1689,N_815,N_858);
xnor U1690 (N_1690,N_1072,N_1046);
nor U1691 (N_1691,N_1207,N_995);
nor U1692 (N_1692,N_961,N_785);
nand U1693 (N_1693,N_1198,N_827);
or U1694 (N_1694,N_921,N_1259);
nor U1695 (N_1695,N_1334,N_1181);
and U1696 (N_1696,N_1432,N_1004);
or U1697 (N_1697,N_1455,N_894);
and U1698 (N_1698,N_1298,N_1255);
or U1699 (N_1699,N_802,N_884);
or U1700 (N_1700,N_1429,N_1452);
nor U1701 (N_1701,N_1468,N_1005);
xnor U1702 (N_1702,N_1194,N_1157);
nor U1703 (N_1703,N_1209,N_1070);
nand U1704 (N_1704,N_1171,N_1216);
nand U1705 (N_1705,N_1482,N_1433);
nor U1706 (N_1706,N_1356,N_852);
xnor U1707 (N_1707,N_1085,N_1333);
nor U1708 (N_1708,N_1267,N_890);
xor U1709 (N_1709,N_1342,N_1476);
xnor U1710 (N_1710,N_1478,N_940);
xnor U1711 (N_1711,N_1141,N_1076);
or U1712 (N_1712,N_841,N_1495);
and U1713 (N_1713,N_752,N_1131);
nand U1714 (N_1714,N_1140,N_1408);
or U1715 (N_1715,N_908,N_787);
nand U1716 (N_1716,N_935,N_1082);
and U1717 (N_1717,N_885,N_1299);
or U1718 (N_1718,N_1063,N_918);
or U1719 (N_1719,N_1258,N_1296);
or U1720 (N_1720,N_1134,N_1252);
or U1721 (N_1721,N_1444,N_1475);
or U1722 (N_1722,N_1337,N_759);
or U1723 (N_1723,N_1314,N_1345);
or U1724 (N_1724,N_833,N_1339);
or U1725 (N_1725,N_851,N_1246);
nand U1726 (N_1726,N_820,N_1032);
or U1727 (N_1727,N_1168,N_1215);
nor U1728 (N_1728,N_1446,N_996);
nor U1729 (N_1729,N_990,N_1428);
nor U1730 (N_1730,N_777,N_821);
xor U1731 (N_1731,N_1165,N_987);
and U1732 (N_1732,N_937,N_844);
and U1733 (N_1733,N_1382,N_1448);
xnor U1734 (N_1734,N_1102,N_1265);
nor U1735 (N_1735,N_1096,N_1064);
or U1736 (N_1736,N_826,N_1136);
and U1737 (N_1737,N_870,N_974);
and U1738 (N_1738,N_1160,N_772);
xor U1739 (N_1739,N_1317,N_1461);
nor U1740 (N_1740,N_764,N_875);
nor U1741 (N_1741,N_1121,N_1388);
nor U1742 (N_1742,N_1484,N_1104);
nor U1743 (N_1743,N_1321,N_1366);
or U1744 (N_1744,N_804,N_924);
and U1745 (N_1745,N_837,N_1097);
xnor U1746 (N_1746,N_1213,N_807);
xnor U1747 (N_1747,N_1392,N_1318);
nor U1748 (N_1748,N_1153,N_1012);
and U1749 (N_1749,N_1237,N_1315);
nand U1750 (N_1750,N_949,N_879);
nor U1751 (N_1751,N_978,N_836);
nor U1752 (N_1752,N_1220,N_783);
and U1753 (N_1753,N_1349,N_1167);
and U1754 (N_1754,N_1006,N_1217);
or U1755 (N_1755,N_1380,N_1411);
or U1756 (N_1756,N_834,N_839);
xor U1757 (N_1757,N_750,N_1049);
nor U1758 (N_1758,N_948,N_1133);
or U1759 (N_1759,N_854,N_781);
and U1760 (N_1760,N_992,N_904);
nand U1761 (N_1761,N_1069,N_1403);
and U1762 (N_1762,N_810,N_1196);
nand U1763 (N_1763,N_1326,N_1059);
nand U1764 (N_1764,N_1013,N_1488);
nand U1765 (N_1765,N_954,N_1185);
or U1766 (N_1766,N_1139,N_769);
nor U1767 (N_1767,N_1212,N_1423);
and U1768 (N_1768,N_1192,N_1113);
nand U1769 (N_1769,N_1203,N_1281);
nor U1770 (N_1770,N_1087,N_1119);
and U1771 (N_1771,N_1341,N_950);
and U1772 (N_1772,N_970,N_1042);
or U1773 (N_1773,N_1201,N_933);
nor U1774 (N_1774,N_830,N_753);
or U1775 (N_1775,N_770,N_878);
nor U1776 (N_1776,N_1440,N_1331);
and U1777 (N_1777,N_986,N_1115);
or U1778 (N_1778,N_1110,N_1079);
nor U1779 (N_1779,N_1191,N_1034);
or U1780 (N_1780,N_963,N_1028);
nand U1781 (N_1781,N_1081,N_1050);
or U1782 (N_1782,N_1389,N_1038);
or U1783 (N_1783,N_1417,N_1234);
nor U1784 (N_1784,N_981,N_1481);
and U1785 (N_1785,N_1088,N_1190);
nand U1786 (N_1786,N_1245,N_1109);
and U1787 (N_1787,N_1402,N_1027);
nand U1788 (N_1788,N_891,N_881);
and U1789 (N_1789,N_784,N_1439);
nor U1790 (N_1790,N_1020,N_1372);
and U1791 (N_1791,N_1307,N_1369);
and U1792 (N_1792,N_929,N_1052);
and U1793 (N_1793,N_1164,N_982);
xor U1794 (N_1794,N_1420,N_1400);
nand U1795 (N_1795,N_983,N_763);
nand U1796 (N_1796,N_1241,N_1312);
nand U1797 (N_1797,N_1357,N_1381);
nand U1798 (N_1798,N_1092,N_1284);
or U1799 (N_1799,N_1243,N_989);
or U1800 (N_1800,N_822,N_964);
nand U1801 (N_1801,N_971,N_1035);
or U1802 (N_1802,N_1414,N_1019);
nor U1803 (N_1803,N_1037,N_1261);
and U1804 (N_1804,N_1413,N_1268);
or U1805 (N_1805,N_1497,N_1127);
and U1806 (N_1806,N_1485,N_893);
nand U1807 (N_1807,N_886,N_1347);
or U1808 (N_1808,N_1169,N_1469);
or U1809 (N_1809,N_824,N_1264);
nor U1810 (N_1810,N_1410,N_867);
or U1811 (N_1811,N_1391,N_1187);
and U1812 (N_1812,N_1221,N_1401);
and U1813 (N_1813,N_847,N_925);
and U1814 (N_1814,N_760,N_1316);
or U1815 (N_1815,N_806,N_1043);
nand U1816 (N_1816,N_1346,N_1214);
or U1817 (N_1817,N_1248,N_1379);
or U1818 (N_1818,N_1351,N_1262);
xnor U1819 (N_1819,N_1177,N_1474);
and U1820 (N_1820,N_1276,N_1457);
or U1821 (N_1821,N_1456,N_1399);
nor U1822 (N_1822,N_1066,N_1151);
nand U1823 (N_1823,N_882,N_1033);
nor U1824 (N_1824,N_942,N_1014);
and U1825 (N_1825,N_892,N_972);
nor U1826 (N_1826,N_1003,N_828);
nor U1827 (N_1827,N_1295,N_1329);
nor U1828 (N_1828,N_905,N_1287);
and U1829 (N_1829,N_842,N_1384);
nand U1830 (N_1830,N_1094,N_1126);
nor U1831 (N_1831,N_1090,N_880);
and U1832 (N_1832,N_1170,N_1138);
or U1833 (N_1833,N_1074,N_1327);
or U1834 (N_1834,N_1294,N_1325);
or U1835 (N_1835,N_1175,N_1309);
and U1836 (N_1836,N_1406,N_1370);
xor U1837 (N_1837,N_1272,N_1277);
nand U1838 (N_1838,N_1077,N_900);
xor U1839 (N_1839,N_1412,N_860);
nand U1840 (N_1840,N_1229,N_1249);
nand U1841 (N_1841,N_927,N_780);
nand U1842 (N_1842,N_1390,N_1183);
xnor U1843 (N_1843,N_829,N_1459);
and U1844 (N_1844,N_779,N_953);
and U1845 (N_1845,N_1426,N_1002);
xnor U1846 (N_1846,N_790,N_1162);
and U1847 (N_1847,N_1462,N_1368);
or U1848 (N_1848,N_1466,N_773);
or U1849 (N_1849,N_1386,N_1155);
xor U1850 (N_1850,N_1421,N_1257);
and U1851 (N_1851,N_795,N_909);
and U1852 (N_1852,N_1335,N_871);
nor U1853 (N_1853,N_1199,N_994);
and U1854 (N_1854,N_899,N_754);
or U1855 (N_1855,N_1197,N_917);
nor U1856 (N_1856,N_761,N_1498);
xnor U1857 (N_1857,N_922,N_906);
nor U1858 (N_1858,N_1283,N_792);
nand U1859 (N_1859,N_1026,N_1445);
nor U1860 (N_1860,N_1494,N_865);
or U1861 (N_1861,N_755,N_1039);
nor U1862 (N_1862,N_1143,N_1130);
nand U1863 (N_1863,N_1067,N_1161);
nand U1864 (N_1864,N_1103,N_923);
and U1865 (N_1865,N_991,N_1060);
and U1866 (N_1866,N_1225,N_775);
and U1867 (N_1867,N_845,N_947);
and U1868 (N_1868,N_1145,N_1285);
nand U1869 (N_1869,N_823,N_1132);
nand U1870 (N_1870,N_1436,N_1242);
and U1871 (N_1871,N_813,N_897);
nand U1872 (N_1872,N_857,N_816);
and U1873 (N_1873,N_1174,N_932);
and U1874 (N_1874,N_1226,N_1179);
nor U1875 (N_1875,N_1428,N_1080);
or U1876 (N_1876,N_788,N_755);
or U1877 (N_1877,N_1143,N_1087);
or U1878 (N_1878,N_1499,N_802);
or U1879 (N_1879,N_950,N_1430);
or U1880 (N_1880,N_881,N_1485);
or U1881 (N_1881,N_960,N_778);
xnor U1882 (N_1882,N_816,N_870);
nor U1883 (N_1883,N_940,N_839);
xnor U1884 (N_1884,N_1124,N_1121);
nand U1885 (N_1885,N_974,N_1348);
and U1886 (N_1886,N_752,N_1266);
and U1887 (N_1887,N_812,N_882);
xnor U1888 (N_1888,N_1064,N_1366);
nor U1889 (N_1889,N_1098,N_901);
and U1890 (N_1890,N_785,N_1316);
xor U1891 (N_1891,N_1283,N_988);
and U1892 (N_1892,N_1360,N_1179);
nor U1893 (N_1893,N_1326,N_1240);
nand U1894 (N_1894,N_1190,N_958);
and U1895 (N_1895,N_1379,N_1044);
nand U1896 (N_1896,N_910,N_1333);
nor U1897 (N_1897,N_1027,N_1270);
nor U1898 (N_1898,N_973,N_1425);
and U1899 (N_1899,N_1426,N_762);
nand U1900 (N_1900,N_1010,N_1122);
or U1901 (N_1901,N_1014,N_1333);
or U1902 (N_1902,N_917,N_801);
and U1903 (N_1903,N_819,N_1348);
nand U1904 (N_1904,N_1213,N_886);
nand U1905 (N_1905,N_1241,N_1055);
or U1906 (N_1906,N_1097,N_831);
and U1907 (N_1907,N_1159,N_1415);
and U1908 (N_1908,N_990,N_1022);
and U1909 (N_1909,N_1025,N_942);
nand U1910 (N_1910,N_831,N_1116);
and U1911 (N_1911,N_1360,N_933);
and U1912 (N_1912,N_1437,N_1385);
and U1913 (N_1913,N_1016,N_967);
and U1914 (N_1914,N_802,N_1468);
or U1915 (N_1915,N_1360,N_1399);
and U1916 (N_1916,N_1086,N_1221);
nor U1917 (N_1917,N_1163,N_1410);
nand U1918 (N_1918,N_841,N_929);
nand U1919 (N_1919,N_1022,N_1402);
or U1920 (N_1920,N_1009,N_940);
and U1921 (N_1921,N_1467,N_1233);
xor U1922 (N_1922,N_1115,N_1140);
and U1923 (N_1923,N_1345,N_1305);
nand U1924 (N_1924,N_779,N_1059);
or U1925 (N_1925,N_1238,N_1070);
nand U1926 (N_1926,N_1254,N_1017);
nand U1927 (N_1927,N_1302,N_1168);
and U1928 (N_1928,N_958,N_1406);
xnor U1929 (N_1929,N_1315,N_1095);
and U1930 (N_1930,N_1083,N_930);
nor U1931 (N_1931,N_1439,N_806);
nor U1932 (N_1932,N_1051,N_1008);
nand U1933 (N_1933,N_1283,N_1388);
or U1934 (N_1934,N_778,N_906);
nor U1935 (N_1935,N_786,N_1298);
and U1936 (N_1936,N_815,N_1095);
or U1937 (N_1937,N_1239,N_1071);
nor U1938 (N_1938,N_904,N_1416);
or U1939 (N_1939,N_1460,N_1362);
nor U1940 (N_1940,N_1483,N_838);
and U1941 (N_1941,N_1484,N_1166);
nand U1942 (N_1942,N_1403,N_1240);
or U1943 (N_1943,N_962,N_969);
nand U1944 (N_1944,N_761,N_1207);
nor U1945 (N_1945,N_1024,N_1243);
and U1946 (N_1946,N_1317,N_1199);
or U1947 (N_1947,N_1246,N_1101);
nand U1948 (N_1948,N_846,N_1374);
nand U1949 (N_1949,N_1261,N_853);
xor U1950 (N_1950,N_1438,N_1431);
nor U1951 (N_1951,N_1127,N_1421);
and U1952 (N_1952,N_1152,N_1171);
xnor U1953 (N_1953,N_1005,N_1438);
nand U1954 (N_1954,N_1288,N_976);
or U1955 (N_1955,N_1452,N_774);
and U1956 (N_1956,N_1168,N_878);
or U1957 (N_1957,N_1478,N_1350);
nor U1958 (N_1958,N_1312,N_1166);
or U1959 (N_1959,N_1260,N_808);
nor U1960 (N_1960,N_1348,N_1219);
nand U1961 (N_1961,N_1080,N_1358);
nor U1962 (N_1962,N_1024,N_1256);
nor U1963 (N_1963,N_1364,N_1268);
xor U1964 (N_1964,N_943,N_1433);
nor U1965 (N_1965,N_1031,N_1444);
xnor U1966 (N_1966,N_1062,N_1323);
and U1967 (N_1967,N_1444,N_1228);
nand U1968 (N_1968,N_850,N_1481);
or U1969 (N_1969,N_908,N_1243);
nor U1970 (N_1970,N_1194,N_1329);
and U1971 (N_1971,N_1206,N_990);
nor U1972 (N_1972,N_806,N_802);
nor U1973 (N_1973,N_1478,N_1411);
or U1974 (N_1974,N_1285,N_926);
and U1975 (N_1975,N_1373,N_1048);
nand U1976 (N_1976,N_1444,N_1014);
xor U1977 (N_1977,N_1426,N_854);
and U1978 (N_1978,N_1277,N_1169);
xnor U1979 (N_1979,N_1008,N_1498);
or U1980 (N_1980,N_1150,N_1423);
or U1981 (N_1981,N_1005,N_1313);
nor U1982 (N_1982,N_1483,N_1263);
and U1983 (N_1983,N_1403,N_920);
and U1984 (N_1984,N_772,N_1312);
nor U1985 (N_1985,N_1121,N_807);
and U1986 (N_1986,N_1116,N_1227);
nor U1987 (N_1987,N_1367,N_792);
or U1988 (N_1988,N_796,N_1479);
xnor U1989 (N_1989,N_1216,N_1060);
nor U1990 (N_1990,N_1221,N_848);
or U1991 (N_1991,N_1121,N_1472);
or U1992 (N_1992,N_1085,N_768);
or U1993 (N_1993,N_1375,N_901);
and U1994 (N_1994,N_1085,N_1050);
or U1995 (N_1995,N_1247,N_962);
nand U1996 (N_1996,N_1178,N_1161);
and U1997 (N_1997,N_1175,N_1008);
nor U1998 (N_1998,N_1384,N_1383);
nor U1999 (N_1999,N_1101,N_1085);
nand U2000 (N_2000,N_857,N_1461);
and U2001 (N_2001,N_1023,N_814);
or U2002 (N_2002,N_1133,N_1225);
and U2003 (N_2003,N_758,N_1457);
nand U2004 (N_2004,N_1039,N_1405);
or U2005 (N_2005,N_1421,N_1142);
nand U2006 (N_2006,N_1011,N_1278);
or U2007 (N_2007,N_1245,N_1152);
nor U2008 (N_2008,N_1231,N_897);
and U2009 (N_2009,N_929,N_1015);
nor U2010 (N_2010,N_1022,N_889);
nand U2011 (N_2011,N_1066,N_798);
nor U2012 (N_2012,N_1329,N_1076);
nand U2013 (N_2013,N_1456,N_1075);
nor U2014 (N_2014,N_1392,N_1081);
and U2015 (N_2015,N_1171,N_1341);
or U2016 (N_2016,N_1345,N_857);
and U2017 (N_2017,N_1431,N_980);
xor U2018 (N_2018,N_936,N_790);
nand U2019 (N_2019,N_809,N_1483);
nand U2020 (N_2020,N_1311,N_1175);
and U2021 (N_2021,N_1082,N_1276);
nand U2022 (N_2022,N_816,N_1280);
or U2023 (N_2023,N_1222,N_1155);
or U2024 (N_2024,N_1454,N_1395);
nor U2025 (N_2025,N_1247,N_1413);
or U2026 (N_2026,N_1169,N_1305);
nand U2027 (N_2027,N_906,N_1022);
and U2028 (N_2028,N_880,N_1322);
nand U2029 (N_2029,N_944,N_1118);
xor U2030 (N_2030,N_1430,N_1213);
nor U2031 (N_2031,N_787,N_1317);
xor U2032 (N_2032,N_1342,N_1368);
or U2033 (N_2033,N_1422,N_1324);
and U2034 (N_2034,N_1166,N_1052);
nor U2035 (N_2035,N_1392,N_1101);
nand U2036 (N_2036,N_768,N_905);
or U2037 (N_2037,N_1114,N_934);
and U2038 (N_2038,N_884,N_1289);
or U2039 (N_2039,N_1424,N_1079);
nand U2040 (N_2040,N_768,N_1386);
xnor U2041 (N_2041,N_822,N_1257);
nor U2042 (N_2042,N_1033,N_1270);
and U2043 (N_2043,N_1106,N_1022);
and U2044 (N_2044,N_1125,N_1391);
nor U2045 (N_2045,N_1088,N_1369);
xnor U2046 (N_2046,N_929,N_885);
nor U2047 (N_2047,N_1156,N_1268);
nor U2048 (N_2048,N_1097,N_987);
nor U2049 (N_2049,N_1267,N_1298);
and U2050 (N_2050,N_817,N_976);
nand U2051 (N_2051,N_888,N_773);
nand U2052 (N_2052,N_1433,N_1200);
or U2053 (N_2053,N_757,N_1385);
and U2054 (N_2054,N_1452,N_1180);
nor U2055 (N_2055,N_1436,N_1142);
nand U2056 (N_2056,N_1441,N_1274);
nand U2057 (N_2057,N_783,N_1282);
or U2058 (N_2058,N_1064,N_796);
nand U2059 (N_2059,N_921,N_1463);
and U2060 (N_2060,N_1046,N_887);
xor U2061 (N_2061,N_1116,N_1308);
nor U2062 (N_2062,N_1092,N_750);
nor U2063 (N_2063,N_1103,N_795);
nand U2064 (N_2064,N_896,N_1041);
nor U2065 (N_2065,N_1170,N_1413);
nand U2066 (N_2066,N_1039,N_891);
and U2067 (N_2067,N_1185,N_1071);
xnor U2068 (N_2068,N_777,N_1044);
and U2069 (N_2069,N_1030,N_1033);
and U2070 (N_2070,N_1291,N_1269);
nand U2071 (N_2071,N_820,N_1013);
nand U2072 (N_2072,N_1277,N_903);
nor U2073 (N_2073,N_1314,N_1228);
and U2074 (N_2074,N_940,N_1286);
or U2075 (N_2075,N_935,N_1176);
and U2076 (N_2076,N_1334,N_1359);
nor U2077 (N_2077,N_1216,N_1263);
nand U2078 (N_2078,N_1429,N_1332);
nand U2079 (N_2079,N_1149,N_895);
xnor U2080 (N_2080,N_1189,N_1230);
nand U2081 (N_2081,N_1440,N_756);
or U2082 (N_2082,N_971,N_1009);
and U2083 (N_2083,N_1292,N_1047);
xor U2084 (N_2084,N_971,N_1277);
nand U2085 (N_2085,N_1255,N_943);
nor U2086 (N_2086,N_784,N_1483);
and U2087 (N_2087,N_1098,N_1207);
nand U2088 (N_2088,N_1457,N_1383);
and U2089 (N_2089,N_982,N_1123);
and U2090 (N_2090,N_764,N_1245);
and U2091 (N_2091,N_1473,N_1072);
or U2092 (N_2092,N_1490,N_1214);
or U2093 (N_2093,N_792,N_1178);
and U2094 (N_2094,N_803,N_1150);
xnor U2095 (N_2095,N_758,N_1145);
nand U2096 (N_2096,N_852,N_1495);
nand U2097 (N_2097,N_907,N_1360);
xnor U2098 (N_2098,N_934,N_778);
and U2099 (N_2099,N_1478,N_805);
nand U2100 (N_2100,N_1108,N_1078);
xnor U2101 (N_2101,N_1237,N_1295);
nand U2102 (N_2102,N_1347,N_1410);
nand U2103 (N_2103,N_1451,N_1424);
nor U2104 (N_2104,N_1241,N_793);
nor U2105 (N_2105,N_997,N_784);
nor U2106 (N_2106,N_1047,N_1167);
and U2107 (N_2107,N_870,N_1055);
nor U2108 (N_2108,N_916,N_1252);
nand U2109 (N_2109,N_820,N_1303);
or U2110 (N_2110,N_931,N_1103);
or U2111 (N_2111,N_1162,N_1084);
or U2112 (N_2112,N_1258,N_1478);
nor U2113 (N_2113,N_1333,N_1355);
or U2114 (N_2114,N_1352,N_913);
nand U2115 (N_2115,N_1037,N_1140);
nor U2116 (N_2116,N_956,N_1357);
or U2117 (N_2117,N_1093,N_1344);
xnor U2118 (N_2118,N_1470,N_1371);
nor U2119 (N_2119,N_1092,N_1083);
nor U2120 (N_2120,N_990,N_1491);
or U2121 (N_2121,N_1099,N_1359);
nand U2122 (N_2122,N_1140,N_949);
nand U2123 (N_2123,N_1352,N_1123);
or U2124 (N_2124,N_771,N_1059);
nor U2125 (N_2125,N_944,N_838);
nor U2126 (N_2126,N_1093,N_868);
nor U2127 (N_2127,N_1318,N_1211);
or U2128 (N_2128,N_1117,N_999);
nor U2129 (N_2129,N_1379,N_1345);
or U2130 (N_2130,N_1093,N_1265);
nor U2131 (N_2131,N_920,N_1427);
nor U2132 (N_2132,N_840,N_786);
and U2133 (N_2133,N_1064,N_1147);
nor U2134 (N_2134,N_1351,N_1045);
xnor U2135 (N_2135,N_1422,N_1459);
or U2136 (N_2136,N_1426,N_879);
xnor U2137 (N_2137,N_1470,N_1390);
nor U2138 (N_2138,N_1121,N_904);
or U2139 (N_2139,N_1069,N_1114);
nor U2140 (N_2140,N_867,N_1330);
or U2141 (N_2141,N_864,N_1303);
nor U2142 (N_2142,N_1343,N_929);
or U2143 (N_2143,N_1290,N_1367);
and U2144 (N_2144,N_897,N_1097);
nand U2145 (N_2145,N_798,N_1170);
and U2146 (N_2146,N_1345,N_901);
nand U2147 (N_2147,N_844,N_1104);
nor U2148 (N_2148,N_808,N_1302);
nor U2149 (N_2149,N_1015,N_1432);
nand U2150 (N_2150,N_1139,N_965);
nand U2151 (N_2151,N_849,N_786);
or U2152 (N_2152,N_1185,N_864);
nor U2153 (N_2153,N_1477,N_1422);
or U2154 (N_2154,N_1013,N_1238);
xor U2155 (N_2155,N_1418,N_1022);
nor U2156 (N_2156,N_1451,N_1392);
nor U2157 (N_2157,N_1413,N_1468);
or U2158 (N_2158,N_1243,N_863);
nand U2159 (N_2159,N_1115,N_1089);
nand U2160 (N_2160,N_1023,N_894);
nor U2161 (N_2161,N_1067,N_790);
nand U2162 (N_2162,N_1391,N_968);
and U2163 (N_2163,N_1071,N_769);
nor U2164 (N_2164,N_1304,N_947);
and U2165 (N_2165,N_1297,N_1162);
or U2166 (N_2166,N_1088,N_1443);
or U2167 (N_2167,N_1260,N_1098);
nand U2168 (N_2168,N_1059,N_1404);
nor U2169 (N_2169,N_981,N_1011);
nor U2170 (N_2170,N_944,N_1415);
or U2171 (N_2171,N_876,N_1195);
or U2172 (N_2172,N_1000,N_1406);
nand U2173 (N_2173,N_1105,N_824);
nand U2174 (N_2174,N_1338,N_1282);
nor U2175 (N_2175,N_1447,N_966);
or U2176 (N_2176,N_989,N_812);
or U2177 (N_2177,N_934,N_1129);
and U2178 (N_2178,N_1356,N_1488);
nand U2179 (N_2179,N_958,N_1431);
nand U2180 (N_2180,N_1017,N_1319);
nor U2181 (N_2181,N_1452,N_1351);
nand U2182 (N_2182,N_991,N_858);
nor U2183 (N_2183,N_769,N_1387);
and U2184 (N_2184,N_1357,N_1210);
nand U2185 (N_2185,N_1469,N_1413);
or U2186 (N_2186,N_984,N_1355);
nand U2187 (N_2187,N_1481,N_928);
and U2188 (N_2188,N_1461,N_1385);
and U2189 (N_2189,N_1378,N_1338);
and U2190 (N_2190,N_962,N_1037);
xor U2191 (N_2191,N_1102,N_1016);
and U2192 (N_2192,N_1163,N_1178);
nand U2193 (N_2193,N_1297,N_926);
and U2194 (N_2194,N_808,N_1301);
nand U2195 (N_2195,N_807,N_1134);
or U2196 (N_2196,N_1191,N_938);
and U2197 (N_2197,N_1143,N_1028);
nand U2198 (N_2198,N_1414,N_1108);
and U2199 (N_2199,N_1198,N_1255);
and U2200 (N_2200,N_1277,N_1021);
and U2201 (N_2201,N_1393,N_1073);
or U2202 (N_2202,N_1069,N_1079);
xnor U2203 (N_2203,N_1219,N_1423);
or U2204 (N_2204,N_1053,N_1245);
and U2205 (N_2205,N_828,N_1497);
or U2206 (N_2206,N_1031,N_1048);
or U2207 (N_2207,N_1086,N_1174);
nor U2208 (N_2208,N_1247,N_779);
and U2209 (N_2209,N_892,N_1357);
or U2210 (N_2210,N_953,N_972);
nand U2211 (N_2211,N_1123,N_787);
and U2212 (N_2212,N_1478,N_1107);
nor U2213 (N_2213,N_1416,N_1405);
nor U2214 (N_2214,N_989,N_1490);
and U2215 (N_2215,N_1025,N_1240);
or U2216 (N_2216,N_1187,N_1481);
or U2217 (N_2217,N_1289,N_1494);
and U2218 (N_2218,N_897,N_1474);
and U2219 (N_2219,N_1424,N_1080);
and U2220 (N_2220,N_1054,N_1036);
nand U2221 (N_2221,N_1043,N_1170);
and U2222 (N_2222,N_1239,N_1135);
nor U2223 (N_2223,N_1268,N_777);
and U2224 (N_2224,N_1247,N_1420);
nand U2225 (N_2225,N_1108,N_1148);
nor U2226 (N_2226,N_761,N_1454);
nand U2227 (N_2227,N_1188,N_1233);
and U2228 (N_2228,N_1217,N_1287);
or U2229 (N_2229,N_1292,N_1050);
and U2230 (N_2230,N_1358,N_1312);
xnor U2231 (N_2231,N_1099,N_1358);
xnor U2232 (N_2232,N_1073,N_751);
or U2233 (N_2233,N_827,N_1429);
or U2234 (N_2234,N_1444,N_1098);
nor U2235 (N_2235,N_1349,N_1469);
or U2236 (N_2236,N_1192,N_907);
and U2237 (N_2237,N_1275,N_1177);
and U2238 (N_2238,N_1111,N_1136);
nand U2239 (N_2239,N_799,N_1241);
or U2240 (N_2240,N_916,N_1451);
nor U2241 (N_2241,N_982,N_1487);
nor U2242 (N_2242,N_1167,N_1347);
nor U2243 (N_2243,N_1036,N_1317);
nand U2244 (N_2244,N_1189,N_1091);
or U2245 (N_2245,N_1026,N_939);
and U2246 (N_2246,N_1433,N_1397);
nand U2247 (N_2247,N_1011,N_1058);
nor U2248 (N_2248,N_1172,N_892);
nor U2249 (N_2249,N_1317,N_1074);
xor U2250 (N_2250,N_1786,N_1547);
nor U2251 (N_2251,N_2092,N_1843);
nor U2252 (N_2252,N_2103,N_2007);
or U2253 (N_2253,N_2175,N_1683);
or U2254 (N_2254,N_2183,N_2073);
or U2255 (N_2255,N_1893,N_1562);
xor U2256 (N_2256,N_2223,N_1984);
nor U2257 (N_2257,N_1540,N_1693);
and U2258 (N_2258,N_2070,N_1587);
or U2259 (N_2259,N_1785,N_1612);
nand U2260 (N_2260,N_1661,N_1765);
and U2261 (N_2261,N_1940,N_1981);
nand U2262 (N_2262,N_1628,N_2116);
nor U2263 (N_2263,N_2205,N_1791);
and U2264 (N_2264,N_2055,N_1611);
nor U2265 (N_2265,N_1688,N_1878);
nand U2266 (N_2266,N_1559,N_1677);
nand U2267 (N_2267,N_1952,N_2237);
nand U2268 (N_2268,N_1660,N_1966);
or U2269 (N_2269,N_2168,N_1859);
xor U2270 (N_2270,N_2090,N_2192);
and U2271 (N_2271,N_2082,N_2005);
nand U2272 (N_2272,N_1701,N_1871);
nand U2273 (N_2273,N_1608,N_2164);
nor U2274 (N_2274,N_2130,N_1741);
nand U2275 (N_2275,N_1576,N_1880);
or U2276 (N_2276,N_1938,N_1528);
nand U2277 (N_2277,N_2200,N_1899);
or U2278 (N_2278,N_1517,N_1697);
or U2279 (N_2279,N_1531,N_1971);
nand U2280 (N_2280,N_1963,N_1778);
and U2281 (N_2281,N_1854,N_1781);
and U2282 (N_2282,N_2064,N_2146);
or U2283 (N_2283,N_2131,N_1754);
or U2284 (N_2284,N_1584,N_1715);
nand U2285 (N_2285,N_1968,N_2085);
or U2286 (N_2286,N_1927,N_2127);
or U2287 (N_2287,N_1998,N_1507);
and U2288 (N_2288,N_1922,N_2136);
nor U2289 (N_2289,N_1732,N_1890);
nor U2290 (N_2290,N_1624,N_1919);
and U2291 (N_2291,N_2034,N_2129);
nand U2292 (N_2292,N_1513,N_1873);
nand U2293 (N_2293,N_1823,N_1947);
nand U2294 (N_2294,N_1616,N_1719);
and U2295 (N_2295,N_1831,N_2102);
nor U2296 (N_2296,N_1635,N_1597);
nand U2297 (N_2297,N_2194,N_1884);
and U2298 (N_2298,N_1995,N_2170);
and U2299 (N_2299,N_2144,N_1606);
xnor U2300 (N_2300,N_1949,N_2178);
and U2301 (N_2301,N_1595,N_2142);
nand U2302 (N_2302,N_1629,N_1681);
xnor U2303 (N_2303,N_2242,N_1652);
or U2304 (N_2304,N_1943,N_1936);
or U2305 (N_2305,N_2167,N_1742);
nor U2306 (N_2306,N_1596,N_1806);
nand U2307 (N_2307,N_1876,N_2246);
or U2308 (N_2308,N_1977,N_1802);
nor U2309 (N_2309,N_1664,N_2213);
nand U2310 (N_2310,N_2061,N_1603);
nand U2311 (N_2311,N_1905,N_2197);
or U2312 (N_2312,N_1735,N_2148);
nand U2313 (N_2313,N_2115,N_2062);
and U2314 (N_2314,N_1727,N_1694);
or U2315 (N_2315,N_2211,N_1812);
nand U2316 (N_2316,N_1544,N_1607);
xor U2317 (N_2317,N_1663,N_1510);
or U2318 (N_2318,N_1768,N_2228);
and U2319 (N_2319,N_1645,N_2180);
or U2320 (N_2320,N_1708,N_1976);
xor U2321 (N_2321,N_1865,N_2195);
xnor U2322 (N_2322,N_2235,N_2023);
xor U2323 (N_2323,N_1524,N_1924);
xnor U2324 (N_2324,N_2037,N_1944);
and U2325 (N_2325,N_1555,N_1901);
and U2326 (N_2326,N_1935,N_1948);
nor U2327 (N_2327,N_1994,N_2137);
nand U2328 (N_2328,N_1908,N_2248);
or U2329 (N_2329,N_2135,N_2222);
or U2330 (N_2330,N_1730,N_1522);
or U2331 (N_2331,N_1578,N_2011);
nor U2332 (N_2332,N_2077,N_2049);
and U2333 (N_2333,N_1717,N_2231);
or U2334 (N_2334,N_1591,N_1918);
nor U2335 (N_2335,N_1851,N_1632);
nand U2336 (N_2336,N_1993,N_1906);
or U2337 (N_2337,N_2145,N_1643);
or U2338 (N_2338,N_1803,N_2132);
nand U2339 (N_2339,N_1761,N_1642);
or U2340 (N_2340,N_1975,N_1511);
nor U2341 (N_2341,N_2100,N_2099);
and U2342 (N_2342,N_1500,N_1684);
xor U2343 (N_2343,N_1749,N_2229);
or U2344 (N_2344,N_2156,N_1996);
nand U2345 (N_2345,N_1932,N_2226);
and U2346 (N_2346,N_1852,N_2159);
nand U2347 (N_2347,N_1921,N_1813);
nor U2348 (N_2348,N_1516,N_1551);
nand U2349 (N_2349,N_2245,N_2191);
and U2350 (N_2350,N_1912,N_2057);
nand U2351 (N_2351,N_1991,N_1739);
nand U2352 (N_2352,N_1866,N_1707);
or U2353 (N_2353,N_1961,N_1759);
or U2354 (N_2354,N_1581,N_2187);
xnor U2355 (N_2355,N_1985,N_2113);
xor U2356 (N_2356,N_1610,N_1755);
xor U2357 (N_2357,N_1824,N_2204);
or U2358 (N_2358,N_1804,N_1667);
nand U2359 (N_2359,N_2009,N_1543);
and U2360 (N_2360,N_2134,N_2042);
nor U2361 (N_2361,N_1917,N_2059);
nand U2362 (N_2362,N_1891,N_1794);
and U2363 (N_2363,N_1712,N_1679);
nor U2364 (N_2364,N_2243,N_1572);
nand U2365 (N_2365,N_1585,N_1680);
nand U2366 (N_2366,N_2177,N_2081);
or U2367 (N_2367,N_1514,N_2190);
and U2368 (N_2368,N_1620,N_1575);
or U2369 (N_2369,N_1841,N_2122);
nor U2370 (N_2370,N_1766,N_2045);
or U2371 (N_2371,N_2174,N_1954);
nor U2372 (N_2372,N_1613,N_1832);
and U2373 (N_2373,N_1907,N_1850);
xor U2374 (N_2374,N_1953,N_1554);
or U2375 (N_2375,N_1594,N_1894);
and U2376 (N_2376,N_1509,N_1877);
and U2377 (N_2377,N_2032,N_2128);
or U2378 (N_2378,N_2214,N_1752);
or U2379 (N_2379,N_1666,N_1779);
nand U2380 (N_2380,N_1671,N_1923);
or U2381 (N_2381,N_2173,N_2014);
nor U2382 (N_2382,N_2186,N_1902);
and U2383 (N_2383,N_1518,N_1860);
nand U2384 (N_2384,N_1637,N_1839);
nor U2385 (N_2385,N_1969,N_2188);
or U2386 (N_2386,N_1973,N_1826);
nor U2387 (N_2387,N_2160,N_1784);
and U2388 (N_2388,N_1744,N_2196);
xor U2389 (N_2389,N_2083,N_2075);
nand U2390 (N_2390,N_2107,N_2120);
nand U2391 (N_2391,N_1598,N_1601);
or U2392 (N_2392,N_1777,N_2044);
and U2393 (N_2393,N_1979,N_1920);
nand U2394 (N_2394,N_1723,N_1974);
and U2395 (N_2395,N_1926,N_1548);
nand U2396 (N_2396,N_2001,N_2114);
or U2397 (N_2397,N_1626,N_2157);
nor U2398 (N_2398,N_2006,N_2105);
and U2399 (N_2399,N_1828,N_2234);
xnor U2400 (N_2400,N_1962,N_1937);
nor U2401 (N_2401,N_2000,N_1848);
xnor U2402 (N_2402,N_1706,N_1668);
and U2403 (N_2403,N_1872,N_1916);
or U2404 (N_2404,N_1763,N_2019);
nand U2405 (N_2405,N_1734,N_2010);
nand U2406 (N_2406,N_2069,N_1521);
xor U2407 (N_2407,N_1800,N_2166);
nand U2408 (N_2408,N_1825,N_1622);
xnor U2409 (N_2409,N_1776,N_1574);
and U2410 (N_2410,N_2236,N_1844);
nand U2411 (N_2411,N_1644,N_2093);
or U2412 (N_2412,N_2112,N_2106);
nor U2413 (N_2413,N_1753,N_1696);
or U2414 (N_2414,N_1900,N_2225);
nand U2415 (N_2415,N_2169,N_1691);
nand U2416 (N_2416,N_1702,N_2249);
xnor U2417 (N_2417,N_1821,N_2052);
nor U2418 (N_2418,N_1997,N_1656);
nand U2419 (N_2419,N_1714,N_1934);
and U2420 (N_2420,N_1711,N_1686);
nor U2421 (N_2421,N_2076,N_1960);
nor U2422 (N_2422,N_2030,N_1834);
nand U2423 (N_2423,N_2022,N_2152);
nor U2424 (N_2424,N_1858,N_2020);
nand U2425 (N_2425,N_1946,N_1563);
nand U2426 (N_2426,N_2218,N_1773);
and U2427 (N_2427,N_2172,N_1951);
xnor U2428 (N_2428,N_1930,N_1748);
nor U2429 (N_2429,N_1743,N_1928);
or U2430 (N_2430,N_2040,N_2054);
or U2431 (N_2431,N_2025,N_1546);
or U2432 (N_2432,N_2124,N_1809);
nor U2433 (N_2433,N_1992,N_2110);
or U2434 (N_2434,N_1810,N_1838);
nand U2435 (N_2435,N_1913,N_2161);
nor U2436 (N_2436,N_2071,N_1830);
nand U2437 (N_2437,N_1541,N_1721);
nor U2438 (N_2438,N_1816,N_1895);
nand U2439 (N_2439,N_2185,N_1835);
or U2440 (N_2440,N_1675,N_1552);
and U2441 (N_2441,N_1990,N_2043);
nor U2442 (N_2442,N_2068,N_1653);
nand U2443 (N_2443,N_1842,N_1700);
or U2444 (N_2444,N_2098,N_2151);
and U2445 (N_2445,N_2067,N_1758);
or U2446 (N_2446,N_1550,N_1530);
or U2447 (N_2447,N_1672,N_2119);
and U2448 (N_2448,N_1793,N_1945);
xnor U2449 (N_2449,N_2247,N_1669);
nand U2450 (N_2450,N_2095,N_2039);
nand U2451 (N_2451,N_2015,N_2028);
nor U2452 (N_2452,N_1967,N_1837);
or U2453 (N_2453,N_1657,N_1568);
nor U2454 (N_2454,N_1775,N_1790);
or U2455 (N_2455,N_1795,N_2215);
and U2456 (N_2456,N_1797,N_1904);
nor U2457 (N_2457,N_1534,N_1634);
nand U2458 (N_2458,N_1950,N_1955);
nor U2459 (N_2459,N_1957,N_1673);
and U2460 (N_2460,N_1845,N_1710);
xor U2461 (N_2461,N_1864,N_1623);
or U2462 (N_2462,N_1592,N_1720);
nor U2463 (N_2463,N_1988,N_1698);
nor U2464 (N_2464,N_1699,N_1986);
nand U2465 (N_2465,N_1737,N_1589);
or U2466 (N_2466,N_1853,N_1888);
and U2467 (N_2467,N_1636,N_1705);
xor U2468 (N_2468,N_2097,N_1978);
and U2469 (N_2469,N_1633,N_2027);
and U2470 (N_2470,N_1756,N_2193);
nand U2471 (N_2471,N_2024,N_2031);
nor U2472 (N_2472,N_1887,N_2241);
xnor U2473 (N_2473,N_1582,N_1615);
nand U2474 (N_2474,N_1716,N_1529);
nand U2475 (N_2475,N_2126,N_1855);
or U2476 (N_2476,N_1539,N_2003);
nor U2477 (N_2477,N_1814,N_2096);
nand U2478 (N_2478,N_1508,N_2171);
and U2479 (N_2479,N_1639,N_2141);
nand U2480 (N_2480,N_1586,N_1692);
or U2481 (N_2481,N_2084,N_1787);
xor U2482 (N_2482,N_2086,N_2091);
nor U2483 (N_2483,N_2079,N_1646);
nor U2484 (N_2484,N_2154,N_2143);
nand U2485 (N_2485,N_2181,N_2002);
nand U2486 (N_2486,N_1736,N_2118);
nand U2487 (N_2487,N_1502,N_1690);
nand U2488 (N_2488,N_1750,N_2080);
xor U2489 (N_2489,N_1774,N_1820);
nor U2490 (N_2490,N_1770,N_1964);
xnor U2491 (N_2491,N_1745,N_1941);
or U2492 (N_2492,N_2021,N_1857);
xnor U2493 (N_2493,N_1862,N_1801);
nand U2494 (N_2494,N_2150,N_1621);
xnor U2495 (N_2495,N_2117,N_1729);
nor U2496 (N_2496,N_2047,N_2212);
and U2497 (N_2497,N_2238,N_2088);
nand U2498 (N_2498,N_1618,N_1863);
and U2499 (N_2499,N_1833,N_1915);
nor U2500 (N_2500,N_1999,N_1771);
and U2501 (N_2501,N_2017,N_1896);
and U2502 (N_2502,N_1874,N_1604);
or U2503 (N_2503,N_2094,N_1815);
xor U2504 (N_2504,N_2038,N_1625);
nor U2505 (N_2505,N_1527,N_2056);
nor U2506 (N_2506,N_1760,N_1658);
and U2507 (N_2507,N_1780,N_2189);
xnor U2508 (N_2508,N_2220,N_1549);
nand U2509 (N_2509,N_1980,N_1783);
nor U2510 (N_2510,N_1535,N_2087);
or U2511 (N_2511,N_2198,N_2046);
nand U2512 (N_2512,N_1678,N_1867);
xnor U2513 (N_2513,N_2155,N_1569);
nor U2514 (N_2514,N_1641,N_1560);
nor U2515 (N_2515,N_2206,N_1757);
nor U2516 (N_2516,N_2140,N_1849);
nand U2517 (N_2517,N_2058,N_1911);
nand U2518 (N_2518,N_1769,N_1713);
or U2519 (N_2519,N_2066,N_1965);
nand U2520 (N_2520,N_1566,N_2012);
nor U2521 (N_2521,N_2230,N_1557);
or U2522 (N_2522,N_2013,N_1903);
and U2523 (N_2523,N_1807,N_1501);
nand U2524 (N_2524,N_1970,N_1879);
and U2525 (N_2525,N_1619,N_1817);
and U2526 (N_2526,N_1875,N_1738);
nand U2527 (N_2527,N_2089,N_1819);
and U2528 (N_2528,N_2208,N_1897);
nor U2529 (N_2529,N_1808,N_2240);
and U2530 (N_2530,N_2008,N_1532);
and U2531 (N_2531,N_1983,N_2125);
xnor U2532 (N_2532,N_2133,N_1818);
or U2533 (N_2533,N_2108,N_1939);
or U2534 (N_2534,N_1519,N_1931);
and U2535 (N_2535,N_1847,N_2176);
nand U2536 (N_2536,N_2139,N_2216);
nand U2537 (N_2537,N_1886,N_1506);
nand U2538 (N_2538,N_2033,N_1630);
nand U2539 (N_2539,N_1805,N_1868);
xnor U2540 (N_2540,N_1605,N_1722);
nand U2541 (N_2541,N_1840,N_2219);
nor U2542 (N_2542,N_1526,N_1685);
or U2543 (N_2543,N_2244,N_1651);
xnor U2544 (N_2544,N_1689,N_1792);
nand U2545 (N_2545,N_1882,N_1525);
nor U2546 (N_2546,N_1538,N_1515);
nor U2547 (N_2547,N_1829,N_2026);
nand U2548 (N_2548,N_1674,N_1798);
and U2549 (N_2549,N_1503,N_1709);
or U2550 (N_2550,N_1536,N_1558);
nand U2551 (N_2551,N_1933,N_1570);
and U2552 (N_2552,N_2153,N_2210);
nor U2553 (N_2553,N_1665,N_2203);
nor U2554 (N_2554,N_1659,N_1811);
nand U2555 (N_2555,N_1579,N_1573);
nand U2556 (N_2556,N_1767,N_1588);
nor U2557 (N_2557,N_1958,N_1987);
and U2558 (N_2558,N_1614,N_1728);
or U2559 (N_2559,N_1638,N_2060);
nor U2560 (N_2560,N_1910,N_2149);
and U2561 (N_2561,N_2065,N_1726);
nor U2562 (N_2562,N_2179,N_1599);
nor U2563 (N_2563,N_1567,N_2163);
and U2564 (N_2564,N_1856,N_1892);
or U2565 (N_2565,N_1670,N_2224);
nand U2566 (N_2566,N_2227,N_1654);
xor U2567 (N_2567,N_1740,N_1695);
and U2568 (N_2568,N_2018,N_1542);
nor U2569 (N_2569,N_1565,N_1898);
nand U2570 (N_2570,N_2078,N_1914);
nand U2571 (N_2571,N_1881,N_1650);
and U2572 (N_2572,N_2217,N_1662);
or U2573 (N_2573,N_1631,N_1883);
xnor U2574 (N_2574,N_1718,N_1782);
and U2575 (N_2575,N_1504,N_2104);
nor U2576 (N_2576,N_1772,N_1725);
or U2577 (N_2577,N_1577,N_1788);
nor U2578 (N_2578,N_1505,N_2111);
nand U2579 (N_2579,N_1982,N_1590);
xor U2580 (N_2580,N_1827,N_1799);
and U2581 (N_2581,N_2201,N_1602);
or U2582 (N_2582,N_2048,N_1989);
and U2583 (N_2583,N_1747,N_2109);
nor U2584 (N_2584,N_1956,N_1537);
xor U2585 (N_2585,N_2147,N_1942);
nand U2586 (N_2586,N_2184,N_1533);
nor U2587 (N_2587,N_1889,N_1731);
xor U2588 (N_2588,N_1593,N_1640);
nand U2589 (N_2589,N_1600,N_2101);
xor U2590 (N_2590,N_1676,N_1869);
nor U2591 (N_2591,N_2138,N_1861);
or U2592 (N_2592,N_1929,N_2209);
and U2593 (N_2593,N_2158,N_1609);
and U2594 (N_2594,N_2041,N_2202);
or U2595 (N_2595,N_1564,N_1520);
nor U2596 (N_2596,N_1647,N_2232);
nand U2597 (N_2597,N_1724,N_1836);
nor U2598 (N_2598,N_1580,N_1649);
nor U2599 (N_2599,N_2072,N_2233);
nand U2600 (N_2600,N_1870,N_1972);
and U2601 (N_2601,N_1909,N_1885);
nor U2602 (N_2602,N_2123,N_1655);
xnor U2603 (N_2603,N_2050,N_2053);
or U2604 (N_2604,N_2207,N_1512);
or U2605 (N_2605,N_1682,N_2162);
nor U2606 (N_2606,N_1617,N_2036);
or U2607 (N_2607,N_2029,N_1583);
or U2608 (N_2608,N_1703,N_1553);
nor U2609 (N_2609,N_1796,N_1545);
nor U2610 (N_2610,N_2074,N_1959);
or U2611 (N_2611,N_1556,N_2063);
or U2612 (N_2612,N_1925,N_1523);
nand U2613 (N_2613,N_2221,N_2121);
or U2614 (N_2614,N_2004,N_2016);
or U2615 (N_2615,N_1704,N_1687);
and U2616 (N_2616,N_1627,N_1648);
nor U2617 (N_2617,N_2165,N_1746);
nand U2618 (N_2618,N_1764,N_1561);
or U2619 (N_2619,N_2199,N_1571);
or U2620 (N_2620,N_2239,N_1733);
nor U2621 (N_2621,N_1762,N_1751);
nand U2622 (N_2622,N_1789,N_2182);
and U2623 (N_2623,N_1822,N_2051);
and U2624 (N_2624,N_1846,N_2035);
nor U2625 (N_2625,N_2130,N_1574);
and U2626 (N_2626,N_2151,N_1825);
nand U2627 (N_2627,N_1855,N_1959);
nand U2628 (N_2628,N_1641,N_2067);
and U2629 (N_2629,N_1886,N_1523);
or U2630 (N_2630,N_2121,N_1871);
xor U2631 (N_2631,N_1616,N_1543);
and U2632 (N_2632,N_1950,N_1579);
or U2633 (N_2633,N_1682,N_2089);
and U2634 (N_2634,N_1802,N_1665);
nor U2635 (N_2635,N_1570,N_1603);
xor U2636 (N_2636,N_1759,N_1706);
xnor U2637 (N_2637,N_2183,N_1637);
xor U2638 (N_2638,N_1990,N_2133);
xor U2639 (N_2639,N_1832,N_1503);
xor U2640 (N_2640,N_1830,N_2244);
nor U2641 (N_2641,N_1675,N_2242);
or U2642 (N_2642,N_2015,N_2202);
or U2643 (N_2643,N_1710,N_1904);
nand U2644 (N_2644,N_1625,N_1510);
nor U2645 (N_2645,N_1537,N_1501);
nand U2646 (N_2646,N_1502,N_1777);
and U2647 (N_2647,N_1564,N_1769);
and U2648 (N_2648,N_2140,N_1914);
or U2649 (N_2649,N_1609,N_1541);
and U2650 (N_2650,N_1775,N_1795);
nand U2651 (N_2651,N_1787,N_2162);
nand U2652 (N_2652,N_1969,N_1530);
xor U2653 (N_2653,N_1846,N_1661);
or U2654 (N_2654,N_1532,N_2065);
and U2655 (N_2655,N_2109,N_1824);
or U2656 (N_2656,N_2018,N_2002);
and U2657 (N_2657,N_2199,N_2065);
xor U2658 (N_2658,N_1530,N_2100);
nand U2659 (N_2659,N_2180,N_1911);
and U2660 (N_2660,N_1552,N_1764);
or U2661 (N_2661,N_1986,N_1619);
nand U2662 (N_2662,N_1818,N_1542);
nand U2663 (N_2663,N_1675,N_1853);
or U2664 (N_2664,N_1920,N_1700);
nand U2665 (N_2665,N_1978,N_1646);
nand U2666 (N_2666,N_2085,N_1665);
nand U2667 (N_2667,N_1516,N_1993);
nand U2668 (N_2668,N_1543,N_2186);
nand U2669 (N_2669,N_1505,N_1553);
and U2670 (N_2670,N_1922,N_2007);
and U2671 (N_2671,N_1789,N_1773);
nand U2672 (N_2672,N_2113,N_1845);
nand U2673 (N_2673,N_1928,N_1599);
and U2674 (N_2674,N_1723,N_1992);
and U2675 (N_2675,N_2087,N_1977);
nor U2676 (N_2676,N_1645,N_1640);
and U2677 (N_2677,N_1725,N_1693);
nor U2678 (N_2678,N_2045,N_1508);
xnor U2679 (N_2679,N_1850,N_1660);
or U2680 (N_2680,N_1735,N_1933);
and U2681 (N_2681,N_1514,N_1518);
nor U2682 (N_2682,N_1545,N_2127);
xnor U2683 (N_2683,N_2097,N_1862);
or U2684 (N_2684,N_1969,N_1579);
nor U2685 (N_2685,N_1919,N_1989);
nor U2686 (N_2686,N_1582,N_1601);
nor U2687 (N_2687,N_2236,N_1972);
xnor U2688 (N_2688,N_1700,N_1824);
nor U2689 (N_2689,N_1540,N_1847);
xor U2690 (N_2690,N_1592,N_1536);
or U2691 (N_2691,N_2004,N_1708);
and U2692 (N_2692,N_1610,N_2188);
nand U2693 (N_2693,N_1734,N_1910);
nor U2694 (N_2694,N_1793,N_1981);
nand U2695 (N_2695,N_2090,N_1743);
xor U2696 (N_2696,N_1654,N_1511);
nand U2697 (N_2697,N_1566,N_2249);
and U2698 (N_2698,N_1545,N_2208);
xnor U2699 (N_2699,N_2061,N_1779);
or U2700 (N_2700,N_1526,N_1521);
and U2701 (N_2701,N_2096,N_1805);
and U2702 (N_2702,N_1622,N_2229);
and U2703 (N_2703,N_2168,N_2134);
nand U2704 (N_2704,N_2191,N_1612);
nand U2705 (N_2705,N_1690,N_2033);
or U2706 (N_2706,N_1828,N_2159);
and U2707 (N_2707,N_2248,N_1580);
or U2708 (N_2708,N_1537,N_1708);
nor U2709 (N_2709,N_1698,N_1915);
nand U2710 (N_2710,N_1567,N_1864);
nor U2711 (N_2711,N_1947,N_1532);
nand U2712 (N_2712,N_2138,N_1725);
nand U2713 (N_2713,N_1510,N_1997);
and U2714 (N_2714,N_1544,N_1589);
xnor U2715 (N_2715,N_1689,N_1509);
xor U2716 (N_2716,N_1930,N_1510);
nor U2717 (N_2717,N_2009,N_1925);
and U2718 (N_2718,N_2141,N_1995);
or U2719 (N_2719,N_1602,N_1746);
nand U2720 (N_2720,N_2072,N_1719);
or U2721 (N_2721,N_1884,N_1786);
or U2722 (N_2722,N_2154,N_2218);
nor U2723 (N_2723,N_1841,N_1909);
and U2724 (N_2724,N_1674,N_1738);
nand U2725 (N_2725,N_1564,N_1704);
nand U2726 (N_2726,N_2197,N_1570);
nor U2727 (N_2727,N_1913,N_2139);
nand U2728 (N_2728,N_2100,N_1784);
nand U2729 (N_2729,N_1852,N_2122);
xor U2730 (N_2730,N_1592,N_1803);
xor U2731 (N_2731,N_1824,N_1539);
nor U2732 (N_2732,N_2029,N_1719);
and U2733 (N_2733,N_2243,N_1820);
and U2734 (N_2734,N_2163,N_2121);
nor U2735 (N_2735,N_1755,N_1835);
nor U2736 (N_2736,N_1725,N_1567);
and U2737 (N_2737,N_1525,N_1786);
or U2738 (N_2738,N_1820,N_1779);
nor U2739 (N_2739,N_1935,N_2213);
or U2740 (N_2740,N_2033,N_2182);
or U2741 (N_2741,N_1895,N_1943);
and U2742 (N_2742,N_1504,N_1598);
nor U2743 (N_2743,N_1647,N_2143);
xnor U2744 (N_2744,N_1777,N_1746);
xor U2745 (N_2745,N_1586,N_1526);
and U2746 (N_2746,N_1548,N_1581);
nor U2747 (N_2747,N_1735,N_1560);
or U2748 (N_2748,N_2063,N_1531);
xor U2749 (N_2749,N_1768,N_1951);
nand U2750 (N_2750,N_1818,N_2017);
nand U2751 (N_2751,N_2080,N_1790);
xnor U2752 (N_2752,N_1638,N_1663);
nand U2753 (N_2753,N_1619,N_1634);
nor U2754 (N_2754,N_1825,N_2169);
nand U2755 (N_2755,N_2223,N_1989);
and U2756 (N_2756,N_1893,N_2077);
or U2757 (N_2757,N_1564,N_1978);
and U2758 (N_2758,N_2059,N_1722);
or U2759 (N_2759,N_2197,N_1659);
and U2760 (N_2760,N_1863,N_1843);
and U2761 (N_2761,N_1702,N_2088);
and U2762 (N_2762,N_2017,N_1761);
xnor U2763 (N_2763,N_2008,N_1898);
nor U2764 (N_2764,N_1836,N_1695);
xor U2765 (N_2765,N_1690,N_2104);
xnor U2766 (N_2766,N_2113,N_1858);
nor U2767 (N_2767,N_2248,N_1568);
or U2768 (N_2768,N_2034,N_2043);
nor U2769 (N_2769,N_1887,N_1769);
or U2770 (N_2770,N_1543,N_2179);
xnor U2771 (N_2771,N_1714,N_2173);
and U2772 (N_2772,N_1723,N_2213);
and U2773 (N_2773,N_1818,N_1916);
or U2774 (N_2774,N_1797,N_2181);
nand U2775 (N_2775,N_2110,N_1776);
or U2776 (N_2776,N_2044,N_1699);
nor U2777 (N_2777,N_2021,N_1510);
nor U2778 (N_2778,N_1532,N_1962);
and U2779 (N_2779,N_2031,N_1583);
or U2780 (N_2780,N_1993,N_1730);
or U2781 (N_2781,N_2186,N_1707);
xor U2782 (N_2782,N_1960,N_1713);
or U2783 (N_2783,N_1977,N_2028);
or U2784 (N_2784,N_1922,N_1885);
xor U2785 (N_2785,N_1845,N_2012);
or U2786 (N_2786,N_1769,N_2111);
and U2787 (N_2787,N_1957,N_2233);
and U2788 (N_2788,N_2197,N_1820);
nor U2789 (N_2789,N_1690,N_1572);
and U2790 (N_2790,N_1882,N_2202);
and U2791 (N_2791,N_1955,N_2094);
nand U2792 (N_2792,N_1937,N_1592);
and U2793 (N_2793,N_1652,N_2165);
or U2794 (N_2794,N_1937,N_1689);
nand U2795 (N_2795,N_2200,N_2162);
and U2796 (N_2796,N_2243,N_2129);
nand U2797 (N_2797,N_2109,N_1901);
and U2798 (N_2798,N_1712,N_2103);
nor U2799 (N_2799,N_2138,N_2123);
nand U2800 (N_2800,N_1845,N_1869);
or U2801 (N_2801,N_1967,N_1506);
nand U2802 (N_2802,N_2071,N_1500);
nor U2803 (N_2803,N_1892,N_2048);
and U2804 (N_2804,N_2085,N_1897);
and U2805 (N_2805,N_2016,N_1537);
or U2806 (N_2806,N_1743,N_1579);
or U2807 (N_2807,N_1653,N_1599);
and U2808 (N_2808,N_2122,N_2142);
or U2809 (N_2809,N_1614,N_2170);
or U2810 (N_2810,N_2047,N_1521);
and U2811 (N_2811,N_1758,N_2153);
nand U2812 (N_2812,N_2005,N_1748);
or U2813 (N_2813,N_1775,N_1578);
or U2814 (N_2814,N_2101,N_2021);
or U2815 (N_2815,N_1727,N_1651);
xor U2816 (N_2816,N_1560,N_1714);
or U2817 (N_2817,N_1628,N_1977);
nand U2818 (N_2818,N_1736,N_2106);
nor U2819 (N_2819,N_1863,N_2067);
or U2820 (N_2820,N_1745,N_1778);
nand U2821 (N_2821,N_2132,N_1615);
nor U2822 (N_2822,N_1554,N_1803);
or U2823 (N_2823,N_1844,N_1645);
nand U2824 (N_2824,N_1919,N_2152);
xnor U2825 (N_2825,N_1539,N_2112);
and U2826 (N_2826,N_2083,N_1945);
nand U2827 (N_2827,N_1806,N_2220);
nor U2828 (N_2828,N_2241,N_1658);
xor U2829 (N_2829,N_2054,N_1887);
nor U2830 (N_2830,N_1528,N_2233);
nor U2831 (N_2831,N_1677,N_1886);
or U2832 (N_2832,N_1588,N_1816);
nor U2833 (N_2833,N_2216,N_1616);
nand U2834 (N_2834,N_1629,N_1643);
and U2835 (N_2835,N_2193,N_1725);
nor U2836 (N_2836,N_1642,N_1791);
xnor U2837 (N_2837,N_2074,N_2019);
xnor U2838 (N_2838,N_2064,N_1725);
nor U2839 (N_2839,N_1892,N_1730);
nand U2840 (N_2840,N_2242,N_1827);
xnor U2841 (N_2841,N_1816,N_1527);
and U2842 (N_2842,N_1582,N_1634);
nor U2843 (N_2843,N_1558,N_1671);
or U2844 (N_2844,N_2240,N_1663);
nor U2845 (N_2845,N_2211,N_2219);
or U2846 (N_2846,N_1987,N_1998);
nor U2847 (N_2847,N_2079,N_1601);
or U2848 (N_2848,N_1852,N_1505);
nor U2849 (N_2849,N_2145,N_2141);
nand U2850 (N_2850,N_1949,N_1807);
or U2851 (N_2851,N_1782,N_2081);
nand U2852 (N_2852,N_1924,N_1554);
xor U2853 (N_2853,N_2190,N_1612);
and U2854 (N_2854,N_2101,N_1912);
or U2855 (N_2855,N_1553,N_2201);
nand U2856 (N_2856,N_1768,N_1916);
and U2857 (N_2857,N_1767,N_1968);
nand U2858 (N_2858,N_1733,N_2073);
and U2859 (N_2859,N_1884,N_2093);
and U2860 (N_2860,N_1721,N_1612);
and U2861 (N_2861,N_2181,N_2140);
and U2862 (N_2862,N_2012,N_1825);
nor U2863 (N_2863,N_1891,N_1988);
and U2864 (N_2864,N_2116,N_1710);
and U2865 (N_2865,N_1550,N_2027);
nand U2866 (N_2866,N_1757,N_1636);
or U2867 (N_2867,N_1533,N_1743);
or U2868 (N_2868,N_1825,N_2062);
xnor U2869 (N_2869,N_2191,N_1833);
and U2870 (N_2870,N_1898,N_1878);
and U2871 (N_2871,N_2089,N_2059);
and U2872 (N_2872,N_1551,N_1940);
nor U2873 (N_2873,N_1720,N_2065);
and U2874 (N_2874,N_1555,N_1796);
nor U2875 (N_2875,N_2187,N_1899);
nand U2876 (N_2876,N_1994,N_1757);
and U2877 (N_2877,N_1920,N_1823);
and U2878 (N_2878,N_2040,N_1789);
xnor U2879 (N_2879,N_2210,N_1695);
nand U2880 (N_2880,N_1749,N_2156);
nand U2881 (N_2881,N_1599,N_1510);
nand U2882 (N_2882,N_2072,N_1769);
or U2883 (N_2883,N_1693,N_2011);
nor U2884 (N_2884,N_1721,N_2227);
nand U2885 (N_2885,N_1590,N_1988);
nor U2886 (N_2886,N_1505,N_2135);
xor U2887 (N_2887,N_1984,N_2221);
nor U2888 (N_2888,N_2230,N_1790);
or U2889 (N_2889,N_2056,N_2023);
nand U2890 (N_2890,N_1709,N_1548);
nand U2891 (N_2891,N_1524,N_1600);
nor U2892 (N_2892,N_1516,N_1973);
xor U2893 (N_2893,N_1867,N_1735);
or U2894 (N_2894,N_1742,N_2099);
or U2895 (N_2895,N_1846,N_2239);
nand U2896 (N_2896,N_1514,N_1570);
or U2897 (N_2897,N_2213,N_1677);
nor U2898 (N_2898,N_1873,N_1522);
nor U2899 (N_2899,N_2166,N_1788);
nor U2900 (N_2900,N_1775,N_2025);
and U2901 (N_2901,N_1551,N_1559);
and U2902 (N_2902,N_1711,N_1600);
nand U2903 (N_2903,N_2064,N_1664);
xor U2904 (N_2904,N_1937,N_2020);
and U2905 (N_2905,N_1584,N_1915);
nand U2906 (N_2906,N_2003,N_1886);
or U2907 (N_2907,N_1710,N_1655);
xor U2908 (N_2908,N_1878,N_1503);
and U2909 (N_2909,N_1698,N_2180);
and U2910 (N_2910,N_2111,N_2013);
nor U2911 (N_2911,N_2240,N_2136);
and U2912 (N_2912,N_2068,N_1789);
nor U2913 (N_2913,N_1758,N_1992);
nor U2914 (N_2914,N_1758,N_1576);
nor U2915 (N_2915,N_1877,N_2085);
xor U2916 (N_2916,N_1879,N_1540);
xor U2917 (N_2917,N_1622,N_1751);
nand U2918 (N_2918,N_2055,N_1680);
nor U2919 (N_2919,N_1907,N_2207);
nor U2920 (N_2920,N_1696,N_1903);
and U2921 (N_2921,N_1599,N_1604);
nor U2922 (N_2922,N_2144,N_1970);
and U2923 (N_2923,N_1830,N_1983);
nor U2924 (N_2924,N_2189,N_2063);
nor U2925 (N_2925,N_2164,N_1919);
and U2926 (N_2926,N_2056,N_1894);
and U2927 (N_2927,N_2073,N_2059);
and U2928 (N_2928,N_1633,N_1706);
and U2929 (N_2929,N_1702,N_2152);
nand U2930 (N_2930,N_2083,N_2080);
and U2931 (N_2931,N_2079,N_1703);
or U2932 (N_2932,N_2148,N_1581);
nor U2933 (N_2933,N_2176,N_1792);
and U2934 (N_2934,N_1819,N_1718);
or U2935 (N_2935,N_1749,N_1721);
and U2936 (N_2936,N_2064,N_1969);
or U2937 (N_2937,N_2022,N_1758);
and U2938 (N_2938,N_2035,N_2083);
and U2939 (N_2939,N_2184,N_1941);
nand U2940 (N_2940,N_1511,N_1602);
nand U2941 (N_2941,N_1511,N_1782);
and U2942 (N_2942,N_1735,N_1571);
nor U2943 (N_2943,N_1514,N_1993);
xor U2944 (N_2944,N_1995,N_1836);
nor U2945 (N_2945,N_1920,N_1531);
nand U2946 (N_2946,N_2012,N_1700);
nor U2947 (N_2947,N_1669,N_2085);
nand U2948 (N_2948,N_1828,N_2213);
xnor U2949 (N_2949,N_2143,N_1718);
nor U2950 (N_2950,N_1959,N_1840);
nor U2951 (N_2951,N_1607,N_2073);
nor U2952 (N_2952,N_1817,N_2001);
or U2953 (N_2953,N_1850,N_2207);
and U2954 (N_2954,N_1991,N_1830);
or U2955 (N_2955,N_1846,N_2034);
and U2956 (N_2956,N_2112,N_2082);
and U2957 (N_2957,N_1543,N_1968);
nand U2958 (N_2958,N_2133,N_2052);
nand U2959 (N_2959,N_2163,N_1670);
nand U2960 (N_2960,N_2111,N_1600);
and U2961 (N_2961,N_1754,N_1866);
or U2962 (N_2962,N_2210,N_1962);
or U2963 (N_2963,N_2090,N_1994);
nand U2964 (N_2964,N_2238,N_2235);
and U2965 (N_2965,N_2245,N_1945);
or U2966 (N_2966,N_1964,N_1527);
nand U2967 (N_2967,N_2177,N_1973);
and U2968 (N_2968,N_1546,N_1715);
nand U2969 (N_2969,N_1926,N_1563);
and U2970 (N_2970,N_1864,N_1945);
and U2971 (N_2971,N_1624,N_1731);
nand U2972 (N_2972,N_1636,N_1877);
and U2973 (N_2973,N_1828,N_1654);
and U2974 (N_2974,N_1722,N_1882);
nand U2975 (N_2975,N_2067,N_1539);
and U2976 (N_2976,N_2032,N_2183);
and U2977 (N_2977,N_2034,N_2209);
xor U2978 (N_2978,N_2247,N_1699);
nand U2979 (N_2979,N_1877,N_2162);
nor U2980 (N_2980,N_2244,N_1928);
nand U2981 (N_2981,N_1885,N_2050);
and U2982 (N_2982,N_2167,N_2133);
or U2983 (N_2983,N_1771,N_2112);
and U2984 (N_2984,N_1553,N_1664);
nor U2985 (N_2985,N_2187,N_2033);
or U2986 (N_2986,N_2176,N_2070);
nand U2987 (N_2987,N_2145,N_1624);
xor U2988 (N_2988,N_2113,N_2104);
or U2989 (N_2989,N_2170,N_1920);
xor U2990 (N_2990,N_1727,N_1940);
or U2991 (N_2991,N_1754,N_1742);
nand U2992 (N_2992,N_1501,N_1989);
and U2993 (N_2993,N_2242,N_2051);
or U2994 (N_2994,N_1846,N_2215);
and U2995 (N_2995,N_1618,N_2242);
nor U2996 (N_2996,N_1676,N_1569);
and U2997 (N_2997,N_1859,N_1986);
nor U2998 (N_2998,N_1547,N_1746);
or U2999 (N_2999,N_1610,N_2081);
nor UO_0 (O_0,N_2864,N_2951);
nor UO_1 (O_1,N_2858,N_2746);
nand UO_2 (O_2,N_2629,N_2299);
and UO_3 (O_3,N_2785,N_2833);
nand UO_4 (O_4,N_2582,N_2314);
and UO_5 (O_5,N_2732,N_2600);
xor UO_6 (O_6,N_2900,N_2980);
and UO_7 (O_7,N_2839,N_2856);
and UO_8 (O_8,N_2487,N_2430);
nor UO_9 (O_9,N_2550,N_2797);
xor UO_10 (O_10,N_2763,N_2283);
nand UO_11 (O_11,N_2310,N_2477);
and UO_12 (O_12,N_2613,N_2394);
or UO_13 (O_13,N_2981,N_2373);
or UO_14 (O_14,N_2846,N_2806);
xor UO_15 (O_15,N_2623,N_2948);
or UO_16 (O_16,N_2699,N_2376);
nor UO_17 (O_17,N_2952,N_2887);
nand UO_18 (O_18,N_2612,N_2554);
and UO_19 (O_19,N_2848,N_2758);
nor UO_20 (O_20,N_2653,N_2304);
nand UO_21 (O_21,N_2821,N_2319);
nor UO_22 (O_22,N_2744,N_2327);
nor UO_23 (O_23,N_2562,N_2463);
nor UO_24 (O_24,N_2320,N_2977);
or UO_25 (O_25,N_2606,N_2584);
nand UO_26 (O_26,N_2474,N_2497);
xnor UO_27 (O_27,N_2943,N_2740);
xor UO_28 (O_28,N_2725,N_2421);
or UO_29 (O_29,N_2647,N_2922);
xnor UO_30 (O_30,N_2380,N_2538);
and UO_31 (O_31,N_2597,N_2250);
xnor UO_32 (O_32,N_2336,N_2985);
and UO_33 (O_33,N_2636,N_2514);
nor UO_34 (O_34,N_2680,N_2339);
nor UO_35 (O_35,N_2891,N_2571);
or UO_36 (O_36,N_2372,N_2490);
and UO_37 (O_37,N_2726,N_2632);
and UO_38 (O_38,N_2999,N_2702);
xnor UO_39 (O_39,N_2860,N_2386);
or UO_40 (O_40,N_2536,N_2899);
and UO_41 (O_41,N_2272,N_2601);
and UO_42 (O_42,N_2989,N_2666);
nand UO_43 (O_43,N_2906,N_2638);
nor UO_44 (O_44,N_2604,N_2729);
or UO_45 (O_45,N_2573,N_2341);
and UO_46 (O_46,N_2302,N_2295);
or UO_47 (O_47,N_2893,N_2264);
xnor UO_48 (O_48,N_2709,N_2589);
nor UO_49 (O_49,N_2622,N_2418);
and UO_50 (O_50,N_2940,N_2649);
and UO_51 (O_51,N_2690,N_2280);
and UO_52 (O_52,N_2933,N_2478);
and UO_53 (O_53,N_2393,N_2834);
and UO_54 (O_54,N_2742,N_2741);
or UO_55 (O_55,N_2458,N_2377);
nand UO_56 (O_56,N_2397,N_2466);
and UO_57 (O_57,N_2930,N_2257);
nor UO_58 (O_58,N_2605,N_2683);
nor UO_59 (O_59,N_2626,N_2396);
and UO_60 (O_60,N_2801,N_2961);
nor UO_61 (O_61,N_2956,N_2455);
nor UO_62 (O_62,N_2531,N_2389);
or UO_63 (O_63,N_2449,N_2401);
xnor UO_64 (O_64,N_2697,N_2657);
or UO_65 (O_65,N_2370,N_2378);
nor UO_66 (O_66,N_2828,N_2588);
xnor UO_67 (O_67,N_2349,N_2585);
nor UO_68 (O_68,N_2820,N_2289);
and UO_69 (O_69,N_2644,N_2790);
and UO_70 (O_70,N_2464,N_2382);
and UO_71 (O_71,N_2306,N_2791);
nand UO_72 (O_72,N_2668,N_2442);
or UO_73 (O_73,N_2772,N_2537);
and UO_74 (O_74,N_2935,N_2390);
or UO_75 (O_75,N_2356,N_2326);
nor UO_76 (O_76,N_2512,N_2260);
nor UO_77 (O_77,N_2403,N_2625);
nor UO_78 (O_78,N_2841,N_2457);
nor UO_79 (O_79,N_2581,N_2851);
or UO_80 (O_80,N_2273,N_2984);
xnor UO_81 (O_81,N_2912,N_2628);
or UO_82 (O_82,N_2901,N_2492);
or UO_83 (O_83,N_2368,N_2574);
xor UO_84 (O_84,N_2794,N_2759);
nor UO_85 (O_85,N_2780,N_2364);
nor UO_86 (O_86,N_2516,N_2593);
nor UO_87 (O_87,N_2251,N_2778);
nor UO_88 (O_88,N_2795,N_2357);
xnor UO_89 (O_89,N_2889,N_2792);
or UO_90 (O_90,N_2722,N_2409);
nand UO_91 (O_91,N_2541,N_2936);
nor UO_92 (O_92,N_2494,N_2796);
xnor UO_93 (O_93,N_2350,N_2942);
and UO_94 (O_94,N_2716,N_2354);
and UO_95 (O_95,N_2934,N_2660);
or UO_96 (O_96,N_2454,N_2501);
and UO_97 (O_97,N_2405,N_2367);
nand UO_98 (O_98,N_2924,N_2361);
and UO_99 (O_99,N_2902,N_2555);
nor UO_100 (O_100,N_2603,N_2691);
nor UO_101 (O_101,N_2506,N_2276);
and UO_102 (O_102,N_2853,N_2640);
xor UO_103 (O_103,N_2460,N_2894);
and UO_104 (O_104,N_2278,N_2347);
xor UO_105 (O_105,N_2521,N_2826);
nor UO_106 (O_106,N_2358,N_2770);
xor UO_107 (O_107,N_2465,N_2342);
or UO_108 (O_108,N_2991,N_2946);
and UO_109 (O_109,N_2496,N_2334);
nor UO_110 (O_110,N_2750,N_2489);
or UO_111 (O_111,N_2570,N_2611);
or UO_112 (O_112,N_2727,N_2602);
or UO_113 (O_113,N_2798,N_2333);
xnor UO_114 (O_114,N_2845,N_2387);
and UO_115 (O_115,N_2534,N_2374);
or UO_116 (O_116,N_2335,N_2705);
nand UO_117 (O_117,N_2954,N_2311);
nor UO_118 (O_118,N_2700,N_2522);
or UO_119 (O_119,N_2544,N_2618);
nand UO_120 (O_120,N_2275,N_2769);
or UO_121 (O_121,N_2266,N_2282);
and UO_122 (O_122,N_2897,N_2486);
nor UO_123 (O_123,N_2712,N_2391);
nor UO_124 (O_124,N_2982,N_2915);
nor UO_125 (O_125,N_2437,N_2768);
xnor UO_126 (O_126,N_2682,N_2748);
nand UO_127 (O_127,N_2782,N_2621);
and UO_128 (O_128,N_2549,N_2929);
or UO_129 (O_129,N_2793,N_2616);
and UO_130 (O_130,N_2706,N_2650);
and UO_131 (O_131,N_2771,N_2484);
nand UO_132 (O_132,N_2819,N_2756);
and UO_133 (O_133,N_2467,N_2423);
xor UO_134 (O_134,N_2976,N_2614);
or UO_135 (O_135,N_2444,N_2656);
nor UO_136 (O_136,N_2747,N_2914);
nor UO_137 (O_137,N_2972,N_2947);
or UO_138 (O_138,N_2825,N_2411);
nor UO_139 (O_139,N_2523,N_2757);
or UO_140 (O_140,N_2329,N_2654);
and UO_141 (O_141,N_2784,N_2822);
and UO_142 (O_142,N_2955,N_2703);
or UO_143 (O_143,N_2526,N_2542);
nor UO_144 (O_144,N_2877,N_2440);
nor UO_145 (O_145,N_2535,N_2472);
nor UO_146 (O_146,N_2296,N_2619);
nor UO_147 (O_147,N_2944,N_2686);
nor UO_148 (O_148,N_2633,N_2662);
nor UO_149 (O_149,N_2525,N_2804);
nor UO_150 (O_150,N_2962,N_2767);
and UO_151 (O_151,N_2328,N_2499);
or UO_152 (O_152,N_2528,N_2736);
or UO_153 (O_153,N_2388,N_2776);
and UO_154 (O_154,N_2469,N_2254);
and UO_155 (O_155,N_2884,N_2590);
or UO_156 (O_156,N_2920,N_2470);
xnor UO_157 (O_157,N_2928,N_2262);
nor UO_158 (O_158,N_2369,N_2994);
nand UO_159 (O_159,N_2451,N_2607);
xor UO_160 (O_160,N_2859,N_2733);
nand UO_161 (O_161,N_2267,N_2321);
nor UO_162 (O_162,N_2745,N_2286);
xor UO_163 (O_163,N_2563,N_2443);
and UO_164 (O_164,N_2755,N_2711);
and UO_165 (O_165,N_2847,N_2849);
or UO_166 (O_166,N_2988,N_2572);
nor UO_167 (O_167,N_2762,N_2359);
or UO_168 (O_168,N_2883,N_2529);
nand UO_169 (O_169,N_2434,N_2840);
and UO_170 (O_170,N_2292,N_2315);
xor UO_171 (O_171,N_2425,N_2575);
or UO_172 (O_172,N_2398,N_2422);
nand UO_173 (O_173,N_2979,N_2500);
or UO_174 (O_174,N_2330,N_2701);
xor UO_175 (O_175,N_2395,N_2432);
nand UO_176 (O_176,N_2371,N_2971);
nand UO_177 (O_177,N_2441,N_2677);
nor UO_178 (O_178,N_2392,N_2363);
or UO_179 (O_179,N_2789,N_2927);
nand UO_180 (O_180,N_2524,N_2803);
or UO_181 (O_181,N_2406,N_2888);
or UO_182 (O_182,N_2865,N_2402);
nand UO_183 (O_183,N_2886,N_2546);
or UO_184 (O_184,N_2491,N_2693);
nand UO_185 (O_185,N_2509,N_2824);
and UO_186 (O_186,N_2399,N_2481);
nor UO_187 (O_187,N_2805,N_2873);
and UO_188 (O_188,N_2895,N_2766);
nor UO_189 (O_189,N_2635,N_2400);
nand UO_190 (O_190,N_2854,N_2268);
nor UO_191 (O_191,N_2688,N_2408);
nor UO_192 (O_192,N_2498,N_2997);
or UO_193 (O_193,N_2459,N_2560);
and UO_194 (O_194,N_2993,N_2527);
xor UO_195 (O_195,N_2714,N_2424);
or UO_196 (O_196,N_2921,N_2485);
nand UO_197 (O_197,N_2907,N_2539);
or UO_198 (O_198,N_2505,N_2713);
and UO_199 (O_199,N_2324,N_2431);
nand UO_200 (O_200,N_2595,N_2375);
and UO_201 (O_201,N_2909,N_2850);
nor UO_202 (O_202,N_2764,N_2673);
xor UO_203 (O_203,N_2968,N_2675);
xor UO_204 (O_204,N_2259,N_2837);
nor UO_205 (O_205,N_2918,N_2513);
nand UO_206 (O_206,N_2519,N_2910);
nand UO_207 (O_207,N_2468,N_2652);
or UO_208 (O_208,N_2631,N_2274);
or UO_209 (O_209,N_2404,N_2843);
or UO_210 (O_210,N_2671,N_2717);
and UO_211 (O_211,N_2303,N_2471);
nor UO_212 (O_212,N_2301,N_2863);
or UO_213 (O_213,N_2429,N_2723);
nor UO_214 (O_214,N_2777,N_2317);
xor UO_215 (O_215,N_2624,N_2724);
and UO_216 (O_216,N_2868,N_2694);
and UO_217 (O_217,N_2676,N_2802);
or UO_218 (O_218,N_2836,N_2645);
nand UO_219 (O_219,N_2473,N_2594);
nand UO_220 (O_220,N_2739,N_2510);
nor UO_221 (O_221,N_2779,N_2285);
nor UO_222 (O_222,N_2852,N_2360);
or UO_223 (O_223,N_2438,N_2617);
nor UO_224 (O_224,N_2291,N_2761);
nand UO_225 (O_225,N_2753,N_2637);
nand UO_226 (O_226,N_2809,N_2558);
nand UO_227 (O_227,N_2911,N_2351);
or UO_228 (O_228,N_2969,N_2577);
and UO_229 (O_229,N_2871,N_2453);
and UO_230 (O_230,N_2892,N_2503);
nor UO_231 (O_231,N_2307,N_2904);
or UO_232 (O_232,N_2446,N_2312);
nor UO_233 (O_233,N_2383,N_2987);
and UO_234 (O_234,N_2252,N_2787);
nor UO_235 (O_235,N_2518,N_2569);
and UO_236 (O_236,N_2659,N_2788);
or UO_237 (O_237,N_2479,N_2331);
or UO_238 (O_238,N_2343,N_2530);
nor UO_239 (O_239,N_2831,N_2931);
or UO_240 (O_240,N_2812,N_2692);
or UO_241 (O_241,N_2681,N_2567);
and UO_242 (O_242,N_2410,N_2881);
nand UO_243 (O_243,N_2832,N_2520);
nor UO_244 (O_244,N_2448,N_2433);
nand UO_245 (O_245,N_2737,N_2419);
nor UO_246 (O_246,N_2735,N_2256);
and UO_247 (O_247,N_2483,N_2258);
xor UO_248 (O_248,N_2811,N_2559);
nand UO_249 (O_249,N_2532,N_2730);
xor UO_250 (O_250,N_2651,N_2598);
and UO_251 (O_251,N_2511,N_2298);
nand UO_252 (O_252,N_2452,N_2835);
nor UO_253 (O_253,N_2810,N_2462);
and UO_254 (O_254,N_2669,N_2495);
nand UO_255 (O_255,N_2658,N_2507);
nand UO_256 (O_256,N_2561,N_2547);
or UO_257 (O_257,N_2332,N_2974);
or UO_258 (O_258,N_2908,N_2707);
and UO_259 (O_259,N_2866,N_2861);
and UO_260 (O_260,N_2905,N_2255);
or UO_261 (O_261,N_2978,N_2545);
and UO_262 (O_262,N_2941,N_2564);
xnor UO_263 (O_263,N_2316,N_2870);
nand UO_264 (O_264,N_2269,N_2667);
xnor UO_265 (O_265,N_2687,N_2456);
and UO_266 (O_266,N_2738,N_2355);
or UO_267 (O_267,N_2308,N_2872);
nand UO_268 (O_268,N_2447,N_2565);
or UO_269 (O_269,N_2879,N_2998);
or UO_270 (O_270,N_2290,N_2996);
and UO_271 (O_271,N_2731,N_2799);
nor UO_272 (O_272,N_2323,N_2715);
nand UO_273 (O_273,N_2695,N_2754);
or UO_274 (O_274,N_2305,N_2609);
or UO_275 (O_275,N_2818,N_2728);
or UO_276 (O_276,N_2678,N_2765);
and UO_277 (O_277,N_2428,N_2813);
and UO_278 (O_278,N_2752,N_2461);
xnor UO_279 (O_279,N_2838,N_2646);
nor UO_280 (O_280,N_2265,N_2566);
xor UO_281 (O_281,N_2515,N_2661);
xor UO_282 (O_282,N_2365,N_2412);
and UO_283 (O_283,N_2540,N_2480);
nand UO_284 (O_284,N_2720,N_2427);
nand UO_285 (O_285,N_2663,N_2482);
nor UO_286 (O_286,N_2953,N_2352);
or UO_287 (O_287,N_2385,N_2965);
nand UO_288 (O_288,N_2337,N_2439);
nand UO_289 (O_289,N_2829,N_2309);
xnor UO_290 (O_290,N_2751,N_2345);
or UO_291 (O_291,N_2346,N_2475);
or UO_292 (O_292,N_2288,N_2990);
xnor UO_293 (O_293,N_2966,N_2414);
nor UO_294 (O_294,N_2963,N_2517);
or UO_295 (O_295,N_2664,N_2689);
nand UO_296 (O_296,N_2708,N_2937);
nor UO_297 (O_297,N_2696,N_2983);
or UO_298 (O_298,N_2919,N_2366);
xor UO_299 (O_299,N_2610,N_2874);
and UO_300 (O_300,N_2344,N_2615);
nand UO_301 (O_301,N_2885,N_2823);
or UO_302 (O_302,N_2642,N_2420);
xor UO_303 (O_303,N_2591,N_2896);
and UO_304 (O_304,N_2719,N_2592);
or UO_305 (O_305,N_2348,N_2445);
or UO_306 (O_306,N_2986,N_2415);
or UO_307 (O_307,N_2816,N_2913);
nand UO_308 (O_308,N_2270,N_2679);
or UO_309 (O_309,N_2284,N_2808);
or UO_310 (O_310,N_2294,N_2533);
or UO_311 (O_311,N_2641,N_2557);
and UO_312 (O_312,N_2655,N_2807);
or UO_313 (O_313,N_2648,N_2760);
nor UO_314 (O_314,N_2923,N_2450);
or UO_315 (O_315,N_2551,N_2857);
and UO_316 (O_316,N_2975,N_2932);
nand UO_317 (O_317,N_2362,N_2734);
xor UO_318 (O_318,N_2970,N_2253);
nor UO_319 (O_319,N_2493,N_2890);
and UO_320 (O_320,N_2903,N_2685);
nor UO_321 (O_321,N_2957,N_2322);
nand UO_322 (O_322,N_2882,N_2880);
or UO_323 (O_323,N_2815,N_2416);
nand UO_324 (O_324,N_2842,N_2867);
nand UO_325 (O_325,N_2917,N_2436);
or UO_326 (O_326,N_2721,N_2973);
nand UO_327 (O_327,N_2381,N_2578);
nand UO_328 (O_328,N_2876,N_2576);
and UO_329 (O_329,N_2608,N_2277);
or UO_330 (O_330,N_2844,N_2587);
or UO_331 (O_331,N_2293,N_2898);
xnor UO_332 (O_332,N_2855,N_2926);
xor UO_333 (O_333,N_2774,N_2916);
nand UO_334 (O_334,N_2508,N_2297);
nor UO_335 (O_335,N_2488,N_2318);
nand UO_336 (O_336,N_2704,N_2639);
nor UO_337 (O_337,N_2586,N_2384);
nor UO_338 (O_338,N_2698,N_2556);
and UO_339 (O_339,N_2583,N_2949);
and UO_340 (O_340,N_2718,N_2814);
nand UO_341 (O_341,N_2543,N_2340);
or UO_342 (O_342,N_2964,N_2773);
and UO_343 (O_343,N_2775,N_2568);
nor UO_344 (O_344,N_2783,N_2261);
and UO_345 (O_345,N_2300,N_2630);
xnor UO_346 (O_346,N_2417,N_2579);
or UO_347 (O_347,N_2502,N_2413);
nand UO_348 (O_348,N_2967,N_2945);
nor UO_349 (O_349,N_2781,N_2670);
xnor UO_350 (O_350,N_2263,N_2875);
and UO_351 (O_351,N_2279,N_2800);
nand UO_352 (O_352,N_2939,N_2950);
and UO_353 (O_353,N_2992,N_2743);
xor UO_354 (O_354,N_2620,N_2960);
nor UO_355 (O_355,N_2684,N_2407);
or UO_356 (O_356,N_2580,N_2271);
or UO_357 (O_357,N_2426,N_2553);
or UO_358 (O_358,N_2338,N_2827);
nand UO_359 (O_359,N_2325,N_2599);
nand UO_360 (O_360,N_2749,N_2552);
and UO_361 (O_361,N_2596,N_2379);
or UO_362 (O_362,N_2817,N_2710);
and UO_363 (O_363,N_2313,N_2672);
and UO_364 (O_364,N_2878,N_2287);
nand UO_365 (O_365,N_2959,N_2958);
nand UO_366 (O_366,N_2627,N_2995);
nor UO_367 (O_367,N_2643,N_2938);
and UO_368 (O_368,N_2634,N_2435);
nand UO_369 (O_369,N_2353,N_2674);
or UO_370 (O_370,N_2869,N_2548);
and UO_371 (O_371,N_2476,N_2925);
xnor UO_372 (O_372,N_2504,N_2665);
nor UO_373 (O_373,N_2830,N_2786);
or UO_374 (O_374,N_2281,N_2862);
nand UO_375 (O_375,N_2519,N_2422);
or UO_376 (O_376,N_2835,N_2422);
nor UO_377 (O_377,N_2559,N_2534);
nand UO_378 (O_378,N_2972,N_2285);
nor UO_379 (O_379,N_2829,N_2364);
nor UO_380 (O_380,N_2263,N_2477);
and UO_381 (O_381,N_2580,N_2567);
or UO_382 (O_382,N_2899,N_2305);
and UO_383 (O_383,N_2399,N_2422);
and UO_384 (O_384,N_2314,N_2998);
nand UO_385 (O_385,N_2411,N_2659);
nand UO_386 (O_386,N_2513,N_2289);
xor UO_387 (O_387,N_2335,N_2310);
and UO_388 (O_388,N_2431,N_2545);
or UO_389 (O_389,N_2260,N_2455);
nand UO_390 (O_390,N_2703,N_2898);
or UO_391 (O_391,N_2250,N_2731);
or UO_392 (O_392,N_2938,N_2854);
and UO_393 (O_393,N_2742,N_2519);
and UO_394 (O_394,N_2882,N_2352);
and UO_395 (O_395,N_2937,N_2516);
nand UO_396 (O_396,N_2562,N_2991);
xnor UO_397 (O_397,N_2979,N_2900);
nor UO_398 (O_398,N_2712,N_2565);
and UO_399 (O_399,N_2631,N_2702);
nand UO_400 (O_400,N_2392,N_2747);
and UO_401 (O_401,N_2654,N_2759);
nor UO_402 (O_402,N_2776,N_2534);
nand UO_403 (O_403,N_2256,N_2850);
nor UO_404 (O_404,N_2982,N_2848);
or UO_405 (O_405,N_2294,N_2499);
or UO_406 (O_406,N_2633,N_2787);
nor UO_407 (O_407,N_2944,N_2510);
xor UO_408 (O_408,N_2772,N_2255);
nor UO_409 (O_409,N_2391,N_2714);
nor UO_410 (O_410,N_2794,N_2346);
and UO_411 (O_411,N_2816,N_2396);
and UO_412 (O_412,N_2474,N_2348);
nor UO_413 (O_413,N_2925,N_2505);
nor UO_414 (O_414,N_2756,N_2752);
or UO_415 (O_415,N_2594,N_2324);
nor UO_416 (O_416,N_2589,N_2480);
xor UO_417 (O_417,N_2382,N_2349);
and UO_418 (O_418,N_2325,N_2588);
nand UO_419 (O_419,N_2333,N_2526);
or UO_420 (O_420,N_2343,N_2253);
xnor UO_421 (O_421,N_2851,N_2709);
and UO_422 (O_422,N_2809,N_2276);
xnor UO_423 (O_423,N_2527,N_2455);
or UO_424 (O_424,N_2763,N_2504);
and UO_425 (O_425,N_2964,N_2625);
nor UO_426 (O_426,N_2954,N_2941);
nand UO_427 (O_427,N_2757,N_2672);
nand UO_428 (O_428,N_2642,N_2443);
or UO_429 (O_429,N_2459,N_2795);
nand UO_430 (O_430,N_2291,N_2943);
nor UO_431 (O_431,N_2691,N_2446);
or UO_432 (O_432,N_2474,N_2456);
or UO_433 (O_433,N_2848,N_2348);
nor UO_434 (O_434,N_2503,N_2312);
nand UO_435 (O_435,N_2773,N_2688);
and UO_436 (O_436,N_2966,N_2956);
xnor UO_437 (O_437,N_2781,N_2485);
nor UO_438 (O_438,N_2821,N_2804);
nand UO_439 (O_439,N_2974,N_2883);
and UO_440 (O_440,N_2758,N_2699);
nand UO_441 (O_441,N_2985,N_2424);
nand UO_442 (O_442,N_2654,N_2520);
or UO_443 (O_443,N_2601,N_2562);
nor UO_444 (O_444,N_2309,N_2416);
xor UO_445 (O_445,N_2984,N_2819);
nor UO_446 (O_446,N_2362,N_2732);
nor UO_447 (O_447,N_2997,N_2881);
nor UO_448 (O_448,N_2967,N_2990);
nor UO_449 (O_449,N_2803,N_2616);
nand UO_450 (O_450,N_2417,N_2442);
and UO_451 (O_451,N_2817,N_2842);
or UO_452 (O_452,N_2649,N_2447);
or UO_453 (O_453,N_2379,N_2943);
and UO_454 (O_454,N_2399,N_2488);
nand UO_455 (O_455,N_2589,N_2660);
and UO_456 (O_456,N_2570,N_2722);
nand UO_457 (O_457,N_2612,N_2978);
nor UO_458 (O_458,N_2400,N_2654);
and UO_459 (O_459,N_2529,N_2579);
nor UO_460 (O_460,N_2644,N_2635);
or UO_461 (O_461,N_2837,N_2953);
and UO_462 (O_462,N_2260,N_2312);
or UO_463 (O_463,N_2933,N_2312);
nor UO_464 (O_464,N_2459,N_2644);
nand UO_465 (O_465,N_2811,N_2382);
xnor UO_466 (O_466,N_2478,N_2712);
or UO_467 (O_467,N_2642,N_2457);
nand UO_468 (O_468,N_2274,N_2839);
or UO_469 (O_469,N_2439,N_2936);
or UO_470 (O_470,N_2275,N_2824);
nor UO_471 (O_471,N_2562,N_2330);
xor UO_472 (O_472,N_2707,N_2706);
nand UO_473 (O_473,N_2540,N_2687);
or UO_474 (O_474,N_2710,N_2440);
and UO_475 (O_475,N_2471,N_2307);
or UO_476 (O_476,N_2372,N_2903);
and UO_477 (O_477,N_2278,N_2502);
or UO_478 (O_478,N_2312,N_2401);
or UO_479 (O_479,N_2682,N_2845);
nor UO_480 (O_480,N_2664,N_2948);
and UO_481 (O_481,N_2257,N_2620);
nor UO_482 (O_482,N_2728,N_2611);
nor UO_483 (O_483,N_2981,N_2335);
nand UO_484 (O_484,N_2529,N_2422);
and UO_485 (O_485,N_2902,N_2443);
nand UO_486 (O_486,N_2755,N_2494);
xor UO_487 (O_487,N_2669,N_2373);
nor UO_488 (O_488,N_2560,N_2554);
nor UO_489 (O_489,N_2524,N_2722);
and UO_490 (O_490,N_2320,N_2469);
and UO_491 (O_491,N_2368,N_2641);
nor UO_492 (O_492,N_2735,N_2715);
xnor UO_493 (O_493,N_2820,N_2665);
xnor UO_494 (O_494,N_2594,N_2727);
nand UO_495 (O_495,N_2824,N_2651);
nand UO_496 (O_496,N_2339,N_2825);
nand UO_497 (O_497,N_2618,N_2436);
and UO_498 (O_498,N_2336,N_2318);
nor UO_499 (O_499,N_2871,N_2358);
endmodule