module basic_750_5000_1000_2_levels_2xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2512,N_2513,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2538,N_2539,N_2540,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2551,N_2552,N_2553,N_2555,N_2556,N_2558,N_2559,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2570,N_2572,N_2575,N_2576,N_2578,N_2580,N_2581,N_2583,N_2585,N_2587,N_2588,N_2590,N_2591,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2602,N_2603,N_2604,N_2605,N_2606,N_2610,N_2611,N_2612,N_2613,N_2615,N_2616,N_2619,N_2623,N_2624,N_2627,N_2628,N_2630,N_2633,N_2634,N_2636,N_2637,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2647,N_2648,N_2649,N_2650,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2664,N_2665,N_2666,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2719,N_2720,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2729,N_2731,N_2732,N_2733,N_2734,N_2735,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2749,N_2750,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2763,N_2765,N_2767,N_2769,N_2771,N_2772,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2791,N_2792,N_2793,N_2795,N_2796,N_2797,N_2800,N_2802,N_2803,N_2804,N_2805,N_2807,N_2808,N_2809,N_2810,N_2811,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2823,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2832,N_2833,N_2834,N_2836,N_2837,N_2838,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2852,N_2853,N_2856,N_2857,N_2858,N_2859,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2877,N_2878,N_2879,N_2880,N_2881,N_2884,N_2885,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2897,N_2898,N_2899,N_2900,N_2901,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2912,N_2913,N_2914,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2936,N_2937,N_2938,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2949,N_2950,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2959,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2973,N_2974,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2999,N_3000,N_3002,N_3003,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3019,N_3020,N_3021,N_3023,N_3024,N_3025,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3040,N_3043,N_3044,N_3045,N_3046,N_3048,N_3049,N_3050,N_3051,N_3052,N_3057,N_3058,N_3060,N_3062,N_3065,N_3066,N_3067,N_3069,N_3071,N_3072,N_3073,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3102,N_3103,N_3104,N_3105,N_3106,N_3108,N_3109,N_3110,N_3111,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3131,N_3132,N_3133,N_3134,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3146,N_3147,N_3148,N_3149,N_3152,N_3155,N_3156,N_3158,N_3159,N_3160,N_3161,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3172,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3188,N_3189,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3216,N_3217,N_3218,N_3220,N_3221,N_3222,N_3224,N_3226,N_3227,N_3228,N_3229,N_3232,N_3234,N_3235,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3244,N_3245,N_3246,N_3248,N_3249,N_3250,N_3252,N_3254,N_3255,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3273,N_3275,N_3276,N_3277,N_3278,N_3280,N_3281,N_3282,N_3284,N_3285,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3295,N_3297,N_3298,N_3299,N_3300,N_3301,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3321,N_3322,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3360,N_3362,N_3364,N_3365,N_3366,N_3367,N_3368,N_3370,N_3371,N_3372,N_3373,N_3375,N_3376,N_3377,N_3378,N_3380,N_3381,N_3383,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3396,N_3397,N_3399,N_3400,N_3402,N_3403,N_3404,N_3405,N_3407,N_3408,N_3409,N_3410,N_3412,N_3413,N_3414,N_3416,N_3418,N_3420,N_3421,N_3422,N_3423,N_3425,N_3426,N_3427,N_3428,N_3429,N_3431,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3442,N_3443,N_3444,N_3445,N_3446,N_3449,N_3450,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3462,N_3463,N_3465,N_3466,N_3467,N_3469,N_3470,N_3471,N_3472,N_3473,N_3475,N_3476,N_3477,N_3478,N_3480,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3502,N_3503,N_3504,N_3505,N_3506,N_3508,N_3509,N_3510,N_3512,N_3513,N_3514,N_3515,N_3516,N_3518,N_3519,N_3521,N_3522,N_3523,N_3525,N_3527,N_3528,N_3529,N_3530,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3540,N_3542,N_3543,N_3544,N_3546,N_3547,N_3548,N_3551,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3568,N_3569,N_3570,N_3571,N_3573,N_3574,N_3575,N_3576,N_3579,N_3580,N_3581,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3592,N_3593,N_3596,N_3597,N_3598,N_3599,N_3602,N_3604,N_3605,N_3606,N_3607,N_3608,N_3611,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3625,N_3626,N_3627,N_3628,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3647,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3672,N_3674,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3690,N_3691,N_3692,N_3693,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3703,N_3705,N_3706,N_3708,N_3709,N_3710,N_3714,N_3716,N_3717,N_3718,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3742,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3759,N_3760,N_3761,N_3762,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3783,N_3784,N_3785,N_3786,N_3787,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3807,N_3809,N_3810,N_3811,N_3813,N_3815,N_3816,N_3817,N_3820,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3842,N_3843,N_3844,N_3846,N_3847,N_3848,N_3849,N_3850,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3859,N_3860,N_3862,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3871,N_3872,N_3873,N_3875,N_3876,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3886,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3901,N_3902,N_3903,N_3904,N_3905,N_3907,N_3909,N_3910,N_3911,N_3912,N_3914,N_3915,N_3916,N_3917,N_3918,N_3920,N_3923,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3934,N_3935,N_3937,N_3938,N_3939,N_3940,N_3941,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3950,N_3951,N_3953,N_3954,N_3955,N_3956,N_3957,N_3959,N_3960,N_3961,N_3963,N_3964,N_3965,N_3966,N_3967,N_3969,N_3970,N_3971,N_3973,N_3974,N_3975,N_3976,N_3977,N_3979,N_3982,N_3984,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4013,N_4014,N_4015,N_4017,N_4018,N_4019,N_4020,N_4022,N_4023,N_4024,N_4025,N_4026,N_4028,N_4029,N_4030,N_4031,N_4033,N_4034,N_4035,N_4038,N_4039,N_4040,N_4041,N_4042,N_4044,N_4046,N_4047,N_4048,N_4049,N_4050,N_4052,N_4053,N_4054,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4066,N_4067,N_4068,N_4070,N_4071,N_4072,N_4074,N_4075,N_4076,N_4077,N_4079,N_4080,N_4081,N_4082,N_4083,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4102,N_4103,N_4104,N_4106,N_4107,N_4108,N_4109,N_4110,N_4113,N_4115,N_4116,N_4117,N_4118,N_4119,N_4121,N_4122,N_4123,N_4125,N_4128,N_4129,N_4130,N_4131,N_4133,N_4134,N_4136,N_4137,N_4138,N_4140,N_4141,N_4142,N_4144,N_4145,N_4146,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4160,N_4161,N_4164,N_4165,N_4166,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4186,N_4187,N_4188,N_4190,N_4192,N_4194,N_4195,N_4196,N_4197,N_4200,N_4202,N_4203,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4226,N_4227,N_4228,N_4229,N_4232,N_4233,N_4234,N_4235,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4262,N_4263,N_4265,N_4266,N_4267,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4280,N_4282,N_4283,N_4284,N_4285,N_4286,N_4288,N_4289,N_4290,N_4291,N_4292,N_4294,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4304,N_4305,N_4307,N_4309,N_4310,N_4311,N_4312,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4324,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4346,N_4347,N_4348,N_4349,N_4351,N_4352,N_4353,N_4354,N_4355,N_4357,N_4358,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4367,N_4368,N_4370,N_4371,N_4372,N_4375,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4385,N_4386,N_4387,N_4388,N_4390,N_4391,N_4392,N_4393,N_4394,N_4397,N_4398,N_4399,N_4400,N_4401,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4457,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4470,N_4472,N_4474,N_4475,N_4476,N_4477,N_4479,N_4480,N_4481,N_4482,N_4483,N_4485,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4534,N_4536,N_4538,N_4539,N_4540,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4563,N_4564,N_4566,N_4568,N_4569,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4584,N_4585,N_4587,N_4588,N_4591,N_4593,N_4594,N_4595,N_4596,N_4598,N_4600,N_4601,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4620,N_4621,N_4623,N_4624,N_4625,N_4628,N_4629,N_4631,N_4633,N_4634,N_4635,N_4637,N_4639,N_4641,N_4642,N_4643,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4679,N_4680,N_4681,N_4682,N_4683,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4698,N_4699,N_4701,N_4702,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4713,N_4714,N_4715,N_4716,N_4718,N_4720,N_4721,N_4723,N_4724,N_4725,N_4728,N_4729,N_4730,N_4732,N_4734,N_4735,N_4738,N_4739,N_4741,N_4743,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4756,N_4758,N_4759,N_4760,N_4761,N_4762,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4776,N_4777,N_4778,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4809,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4839,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4851,N_4852,N_4856,N_4857,N_4858,N_4859,N_4860,N_4862,N_4863,N_4864,N_4865,N_4867,N_4868,N_4870,N_4871,N_4872,N_4873,N_4875,N_4876,N_4877,N_4878,N_4880,N_4881,N_4883,N_4884,N_4885,N_4886,N_4888,N_4889,N_4890,N_4893,N_4894,N_4895,N_4896,N_4898,N_4899,N_4900,N_4901,N_4903,N_4904,N_4906,N_4907,N_4909,N_4910,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4939,N_4940,N_4941,N_4942,N_4943,N_4945,N_4946,N_4947,N_4948,N_4949,N_4951,N_4952,N_4953,N_4955,N_4956,N_4957,N_4958,N_4960,N_4961,N_4962,N_4963,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4973,N_4974,N_4975,N_4976,N_4977,N_4979,N_4980,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
and U0 (N_0,In_267,In_349);
or U1 (N_1,In_330,In_558);
and U2 (N_2,In_34,In_475);
and U3 (N_3,In_309,In_458);
nand U4 (N_4,In_727,In_742);
or U5 (N_5,In_235,In_142);
nor U6 (N_6,In_512,In_749);
nor U7 (N_7,In_269,In_470);
nor U8 (N_8,In_598,In_407);
or U9 (N_9,In_250,In_438);
or U10 (N_10,In_2,In_264);
and U11 (N_11,In_333,In_87);
and U12 (N_12,In_36,In_523);
and U13 (N_13,In_312,In_107);
or U14 (N_14,In_599,In_41);
nor U15 (N_15,In_383,In_204);
and U16 (N_16,In_467,In_553);
nand U17 (N_17,In_745,In_94);
nor U18 (N_18,In_251,In_108);
nand U19 (N_19,In_640,In_601);
or U20 (N_20,In_404,In_95);
or U21 (N_21,In_261,In_389);
nor U22 (N_22,In_741,In_189);
or U23 (N_23,In_221,In_284);
nor U24 (N_24,In_203,In_595);
nor U25 (N_25,In_89,In_588);
or U26 (N_26,In_700,In_431);
or U27 (N_27,In_303,In_670);
and U28 (N_28,In_155,In_535);
and U29 (N_29,In_394,In_217);
and U30 (N_30,In_265,In_65);
nand U31 (N_31,In_571,In_143);
nor U32 (N_32,In_564,In_707);
nand U33 (N_33,In_304,In_540);
or U34 (N_34,In_324,In_559);
nor U35 (N_35,In_660,In_659);
and U36 (N_36,In_332,In_583);
nand U37 (N_37,In_287,In_225);
nand U38 (N_38,In_694,In_735);
nand U39 (N_39,In_300,In_445);
nor U40 (N_40,In_328,In_630);
nand U41 (N_41,In_131,In_198);
nand U42 (N_42,In_563,In_657);
and U43 (N_43,In_231,In_684);
nand U44 (N_44,In_341,In_353);
or U45 (N_45,In_248,In_575);
nor U46 (N_46,In_104,In_704);
and U47 (N_47,In_562,In_10);
nand U48 (N_48,In_42,In_581);
nor U49 (N_49,In_151,In_663);
or U50 (N_50,In_413,In_200);
and U51 (N_51,In_127,In_162);
nor U52 (N_52,In_218,In_212);
nor U53 (N_53,In_323,In_592);
nand U54 (N_54,In_703,In_279);
and U55 (N_55,In_359,In_446);
xor U56 (N_56,In_585,In_711);
and U57 (N_57,In_40,In_129);
and U58 (N_58,In_271,In_75);
xnor U59 (N_59,In_292,In_435);
or U60 (N_60,In_488,In_12);
and U61 (N_61,In_568,In_125);
nand U62 (N_62,In_26,In_392);
or U63 (N_63,In_709,In_693);
xor U64 (N_64,In_652,In_105);
nand U65 (N_65,In_343,In_288);
or U66 (N_66,In_260,In_443);
and U67 (N_67,In_245,In_718);
nor U68 (N_68,In_406,In_723);
nand U69 (N_69,In_298,In_560);
or U70 (N_70,In_52,In_199);
nor U71 (N_71,In_0,In_422);
nor U72 (N_72,In_25,In_346);
and U73 (N_73,In_124,In_715);
or U74 (N_74,In_335,In_380);
or U75 (N_75,In_112,In_24);
nor U76 (N_76,In_364,In_465);
nor U77 (N_77,In_123,In_427);
and U78 (N_78,In_713,In_14);
nand U79 (N_79,In_132,In_172);
or U80 (N_80,In_209,In_355);
nand U81 (N_81,In_738,In_194);
xnor U82 (N_82,In_505,In_717);
nand U83 (N_83,In_450,In_229);
and U84 (N_84,In_669,In_702);
and U85 (N_85,In_520,In_545);
or U86 (N_86,In_536,In_532);
nor U87 (N_87,In_276,In_331);
and U88 (N_88,In_325,In_188);
or U89 (N_89,In_134,In_117);
nor U90 (N_90,In_401,In_593);
nand U91 (N_91,In_701,In_420);
nand U92 (N_92,In_487,In_442);
and U93 (N_93,In_495,In_395);
and U94 (N_94,In_186,In_529);
and U95 (N_95,In_626,In_734);
and U96 (N_96,In_725,In_430);
or U97 (N_97,In_469,In_187);
nor U98 (N_98,In_139,In_739);
nand U99 (N_99,In_351,In_339);
and U100 (N_100,In_531,In_586);
or U101 (N_101,In_432,In_482);
nor U102 (N_102,In_547,In_128);
nor U103 (N_103,In_297,In_522);
and U104 (N_104,In_354,In_211);
nand U105 (N_105,In_79,In_100);
and U106 (N_106,In_662,In_444);
nor U107 (N_107,In_732,In_414);
and U108 (N_108,In_140,In_681);
nor U109 (N_109,In_665,In_629);
nand U110 (N_110,In_290,In_255);
nand U111 (N_111,In_410,In_546);
and U112 (N_112,In_68,In_146);
nand U113 (N_113,In_476,In_381);
or U114 (N_114,In_173,In_180);
nor U115 (N_115,In_368,In_305);
and U116 (N_116,In_539,In_115);
and U117 (N_117,In_569,In_460);
and U118 (N_118,In_637,In_177);
nor U119 (N_119,In_471,In_83);
nor U120 (N_120,In_415,In_237);
xnor U121 (N_121,In_296,In_69);
nand U122 (N_122,In_405,In_463);
or U123 (N_123,In_602,In_39);
and U124 (N_124,In_480,In_13);
nor U125 (N_125,In_461,In_433);
or U126 (N_126,In_656,In_321);
and U127 (N_127,In_604,In_600);
xor U128 (N_128,In_508,In_295);
nand U129 (N_129,In_215,In_500);
nor U130 (N_130,In_90,In_348);
and U131 (N_131,In_737,In_277);
nor U132 (N_132,In_206,In_541);
and U133 (N_133,In_30,In_516);
nor U134 (N_134,In_257,In_137);
nor U135 (N_135,In_646,In_740);
nor U136 (N_136,In_518,In_426);
or U137 (N_137,In_572,In_506);
nor U138 (N_138,In_136,In_249);
nor U139 (N_139,In_399,In_289);
nand U140 (N_140,In_428,In_192);
and U141 (N_141,In_627,In_148);
and U142 (N_142,In_273,In_610);
and U143 (N_143,In_370,In_678);
and U144 (N_144,In_687,In_207);
or U145 (N_145,In_133,In_336);
and U146 (N_146,In_214,In_54);
and U147 (N_147,In_391,In_497);
and U148 (N_148,In_486,In_570);
and U149 (N_149,In_99,In_548);
and U150 (N_150,In_641,In_674);
or U151 (N_151,In_419,In_596);
nand U152 (N_152,In_538,In_376);
or U153 (N_153,In_719,In_113);
and U154 (N_154,In_159,In_603);
nor U155 (N_155,In_416,In_220);
nor U156 (N_156,In_167,In_526);
and U157 (N_157,In_474,In_576);
and U158 (N_158,In_153,In_165);
or U159 (N_159,In_286,In_650);
nand U160 (N_160,In_633,In_712);
xor U161 (N_161,In_55,In_521);
nor U162 (N_162,In_747,In_621);
xor U163 (N_163,In_233,In_18);
or U164 (N_164,In_57,In_126);
or U165 (N_165,In_110,In_92);
and U166 (N_166,In_574,In_258);
nor U167 (N_167,In_566,In_8);
nand U168 (N_168,In_385,In_350);
nand U169 (N_169,In_86,In_239);
or U170 (N_170,In_106,In_63);
and U171 (N_171,In_363,In_266);
and U172 (N_172,In_377,In_408);
nor U173 (N_173,In_197,In_565);
nand U174 (N_174,In_318,In_96);
and U175 (N_175,In_326,In_64);
xnor U176 (N_176,In_294,In_22);
and U177 (N_177,In_243,In_542);
nand U178 (N_178,In_32,In_623);
and U179 (N_179,In_356,In_44);
nand U180 (N_180,In_714,In_390);
nand U181 (N_181,In_116,In_418);
and U182 (N_182,In_4,In_334);
or U183 (N_183,In_421,In_149);
nand U184 (N_184,In_668,In_530);
and U185 (N_185,In_178,In_639);
or U186 (N_186,In_425,In_78);
and U187 (N_187,In_379,In_746);
nor U188 (N_188,In_283,In_384);
nor U189 (N_189,In_82,In_612);
nor U190 (N_190,In_7,In_317);
nand U191 (N_191,In_280,In_252);
nor U192 (N_192,In_454,In_160);
and U193 (N_193,In_347,In_679);
and U194 (N_194,In_56,In_31);
nand U195 (N_195,In_358,In_238);
nor U196 (N_196,In_77,In_468);
nand U197 (N_197,In_479,In_20);
nand U198 (N_198,In_477,In_1);
and U199 (N_199,In_120,In_372);
nor U200 (N_200,In_201,In_164);
nor U201 (N_201,In_683,In_176);
or U202 (N_202,In_278,In_281);
or U203 (N_203,In_247,In_424);
nand U204 (N_204,In_748,In_71);
and U205 (N_205,In_451,In_561);
or U206 (N_206,In_344,In_114);
or U207 (N_207,In_244,In_150);
or U208 (N_208,In_411,In_527);
nand U209 (N_209,In_169,In_550);
nor U210 (N_210,In_357,In_729);
nor U211 (N_211,In_316,In_447);
nor U212 (N_212,In_509,In_744);
and U213 (N_213,In_111,In_642);
and U214 (N_214,In_135,In_653);
nand U215 (N_215,In_622,In_644);
nor U216 (N_216,In_118,In_607);
or U217 (N_217,In_23,In_66);
and U218 (N_218,In_185,In_434);
and U219 (N_219,In_171,In_181);
nand U220 (N_220,In_49,In_70);
and U221 (N_221,In_613,In_27);
and U222 (N_222,In_726,In_489);
nor U223 (N_223,In_584,In_708);
or U224 (N_224,In_691,In_664);
or U225 (N_225,In_375,In_692);
and U226 (N_226,In_567,In_667);
nor U227 (N_227,In_360,In_609);
and U228 (N_228,In_525,In_190);
and U229 (N_229,In_624,In_382);
and U230 (N_230,In_21,In_170);
or U231 (N_231,In_645,In_671);
or U232 (N_232,In_589,In_606);
and U233 (N_233,In_308,In_174);
or U234 (N_234,In_80,In_224);
and U235 (N_235,In_722,In_412);
or U236 (N_236,In_195,In_322);
nor U237 (N_237,In_73,In_145);
or U238 (N_238,In_631,In_676);
nor U239 (N_239,In_661,In_436);
nor U240 (N_240,In_400,In_441);
nor U241 (N_241,In_483,In_282);
nor U242 (N_242,In_84,In_697);
nor U243 (N_243,In_647,In_590);
and U244 (N_244,In_594,In_302);
nand U245 (N_245,In_699,In_234);
nor U246 (N_246,In_716,In_440);
nand U247 (N_247,In_138,In_61);
nor U248 (N_248,In_98,In_50);
and U249 (N_249,In_614,In_329);
nand U250 (N_250,In_513,In_361);
or U251 (N_251,In_557,In_270);
or U252 (N_252,In_528,In_473);
and U253 (N_253,In_103,In_371);
or U254 (N_254,In_366,In_11);
and U255 (N_255,In_19,In_232);
and U256 (N_256,In_320,In_388);
nor U257 (N_257,In_97,In_580);
nand U258 (N_258,In_552,In_5);
nor U259 (N_259,In_449,In_362);
nand U260 (N_260,In_76,In_731);
or U261 (N_261,In_705,In_291);
and U262 (N_262,In_503,In_310);
nor U263 (N_263,In_152,In_398);
nor U264 (N_264,In_373,In_365);
nand U265 (N_265,In_462,In_58);
or U266 (N_266,In_109,In_119);
and U267 (N_267,In_240,In_511);
nor U268 (N_268,In_396,In_501);
or U269 (N_269,In_515,In_397);
or U270 (N_270,In_369,In_493);
and U271 (N_271,In_314,In_507);
nand U272 (N_272,In_675,In_534);
nand U273 (N_273,In_619,In_459);
nor U274 (N_274,In_611,In_367);
or U275 (N_275,In_578,In_274);
or U276 (N_276,In_638,In_43);
nor U277 (N_277,In_685,In_337);
nand U278 (N_278,In_268,In_253);
and U279 (N_279,In_48,In_196);
or U280 (N_280,In_182,In_743);
and U281 (N_281,In_72,In_494);
or U282 (N_282,In_677,In_386);
and U283 (N_283,In_45,In_736);
nor U284 (N_284,In_456,In_387);
and U285 (N_285,In_184,In_393);
and U286 (N_286,In_340,In_17);
nor U287 (N_287,In_689,In_625);
nor U288 (N_288,In_161,In_618);
or U289 (N_289,In_293,In_696);
or U290 (N_290,In_51,In_374);
or U291 (N_291,In_130,In_616);
and U292 (N_292,In_183,In_498);
nor U293 (N_293,In_88,In_33);
nor U294 (N_294,In_537,In_147);
nor U295 (N_295,In_591,In_556);
or U296 (N_296,In_299,In_551);
and U297 (N_297,In_35,In_236);
nand U298 (N_298,In_210,In_403);
xnor U299 (N_299,In_327,In_439);
nor U300 (N_300,In_643,In_524);
nor U301 (N_301,In_311,In_549);
nand U302 (N_302,In_423,In_554);
nor U303 (N_303,In_175,In_6);
nor U304 (N_304,In_59,In_216);
xnor U305 (N_305,In_533,In_122);
nor U306 (N_306,In_658,In_587);
or U307 (N_307,In_263,In_655);
nand U308 (N_308,In_491,In_227);
nor U309 (N_309,In_706,In_651);
or U310 (N_310,In_46,In_228);
or U311 (N_311,In_654,In_121);
nor U312 (N_312,In_648,In_85);
nand U313 (N_313,In_338,In_673);
nand U314 (N_314,In_695,In_345);
nor U315 (N_315,In_579,In_262);
nor U316 (N_316,In_16,In_466);
nor U317 (N_317,In_191,In_246);
nor U318 (N_318,In_60,In_499);
and U319 (N_319,In_455,In_710);
nor U320 (N_320,In_315,In_457);
or U321 (N_321,In_91,In_93);
or U322 (N_322,In_272,In_686);
or U323 (N_323,In_634,In_649);
or U324 (N_324,In_636,In_53);
or U325 (N_325,In_74,In_484);
and U326 (N_326,In_156,In_620);
and U327 (N_327,In_285,In_158);
or U328 (N_328,In_605,In_213);
nor U329 (N_329,In_666,In_29);
and U330 (N_330,In_730,In_28);
and U331 (N_331,In_259,In_519);
or U332 (N_332,In_573,In_492);
nor U333 (N_333,In_632,In_230);
and U334 (N_334,In_544,In_222);
or U335 (N_335,In_721,In_307);
or U336 (N_336,In_452,In_163);
and U337 (N_337,In_342,In_254);
nor U338 (N_338,In_485,In_608);
nor U339 (N_339,In_502,In_306);
and U340 (N_340,In_15,In_429);
nor U341 (N_341,In_223,In_226);
nor U342 (N_342,In_67,In_688);
or U343 (N_343,In_682,In_490);
nor U344 (N_344,In_219,In_417);
and U345 (N_345,In_378,In_680);
nand U346 (N_346,In_504,In_275);
and U347 (N_347,In_628,In_3);
nor U348 (N_348,In_193,In_38);
and U349 (N_349,In_478,In_733);
nor U350 (N_350,In_154,In_144);
nand U351 (N_351,In_179,In_101);
nand U352 (N_352,In_37,In_517);
nand U353 (N_353,In_690,In_448);
and U354 (N_354,In_352,In_555);
and U355 (N_355,In_319,In_481);
or U356 (N_356,In_205,In_464);
nand U357 (N_357,In_543,In_301);
nor U358 (N_358,In_672,In_81);
and U359 (N_359,In_166,In_9);
nor U360 (N_360,In_256,In_313);
or U361 (N_361,In_208,In_472);
or U362 (N_362,In_168,In_724);
nor U363 (N_363,In_202,In_242);
nand U364 (N_364,In_615,In_141);
or U365 (N_365,In_241,In_453);
nand U366 (N_366,In_402,In_409);
nor U367 (N_367,In_102,In_47);
and U368 (N_368,In_496,In_582);
nor U369 (N_369,In_157,In_577);
xor U370 (N_370,In_514,In_597);
or U371 (N_371,In_720,In_617);
or U372 (N_372,In_437,In_635);
and U373 (N_373,In_510,In_728);
or U374 (N_374,In_698,In_62);
nor U375 (N_375,In_486,In_496);
and U376 (N_376,In_228,In_449);
and U377 (N_377,In_240,In_428);
nand U378 (N_378,In_94,In_247);
or U379 (N_379,In_663,In_622);
nand U380 (N_380,In_200,In_280);
nor U381 (N_381,In_207,In_29);
or U382 (N_382,In_197,In_193);
nor U383 (N_383,In_292,In_431);
xnor U384 (N_384,In_735,In_2);
and U385 (N_385,In_735,In_367);
or U386 (N_386,In_154,In_233);
nand U387 (N_387,In_742,In_673);
nor U388 (N_388,In_25,In_140);
nand U389 (N_389,In_637,In_708);
and U390 (N_390,In_256,In_136);
and U391 (N_391,In_415,In_222);
or U392 (N_392,In_308,In_123);
or U393 (N_393,In_213,In_525);
and U394 (N_394,In_591,In_289);
and U395 (N_395,In_526,In_500);
nand U396 (N_396,In_602,In_616);
nor U397 (N_397,In_600,In_397);
and U398 (N_398,In_698,In_6);
and U399 (N_399,In_411,In_694);
nor U400 (N_400,In_647,In_83);
nor U401 (N_401,In_528,In_203);
nand U402 (N_402,In_719,In_597);
and U403 (N_403,In_185,In_80);
or U404 (N_404,In_564,In_315);
nand U405 (N_405,In_642,In_295);
nor U406 (N_406,In_649,In_420);
nor U407 (N_407,In_311,In_554);
and U408 (N_408,In_10,In_466);
nor U409 (N_409,In_317,In_219);
or U410 (N_410,In_188,In_496);
nor U411 (N_411,In_231,In_92);
and U412 (N_412,In_306,In_44);
and U413 (N_413,In_173,In_737);
or U414 (N_414,In_136,In_91);
or U415 (N_415,In_629,In_74);
nand U416 (N_416,In_709,In_23);
or U417 (N_417,In_611,In_143);
and U418 (N_418,In_375,In_744);
and U419 (N_419,In_66,In_136);
nand U420 (N_420,In_517,In_412);
nor U421 (N_421,In_664,In_735);
or U422 (N_422,In_589,In_347);
nor U423 (N_423,In_560,In_156);
nand U424 (N_424,In_145,In_175);
or U425 (N_425,In_150,In_363);
and U426 (N_426,In_748,In_458);
and U427 (N_427,In_729,In_77);
and U428 (N_428,In_134,In_407);
or U429 (N_429,In_589,In_310);
or U430 (N_430,In_671,In_490);
nand U431 (N_431,In_164,In_92);
and U432 (N_432,In_731,In_196);
and U433 (N_433,In_414,In_15);
nor U434 (N_434,In_253,In_244);
nand U435 (N_435,In_292,In_534);
xnor U436 (N_436,In_362,In_725);
or U437 (N_437,In_64,In_330);
or U438 (N_438,In_72,In_721);
nand U439 (N_439,In_490,In_381);
nor U440 (N_440,In_12,In_416);
and U441 (N_441,In_69,In_155);
or U442 (N_442,In_583,In_638);
nor U443 (N_443,In_716,In_681);
or U444 (N_444,In_690,In_108);
nand U445 (N_445,In_111,In_75);
or U446 (N_446,In_237,In_167);
and U447 (N_447,In_148,In_262);
nor U448 (N_448,In_569,In_522);
nand U449 (N_449,In_629,In_121);
nand U450 (N_450,In_197,In_574);
or U451 (N_451,In_568,In_104);
nor U452 (N_452,In_256,In_56);
and U453 (N_453,In_581,In_530);
or U454 (N_454,In_384,In_185);
and U455 (N_455,In_481,In_517);
and U456 (N_456,In_722,In_331);
nand U457 (N_457,In_657,In_265);
or U458 (N_458,In_711,In_502);
nor U459 (N_459,In_608,In_302);
and U460 (N_460,In_176,In_657);
nor U461 (N_461,In_746,In_477);
or U462 (N_462,In_710,In_363);
nor U463 (N_463,In_448,In_399);
nor U464 (N_464,In_655,In_65);
or U465 (N_465,In_430,In_324);
nand U466 (N_466,In_419,In_169);
xor U467 (N_467,In_401,In_149);
or U468 (N_468,In_312,In_496);
nor U469 (N_469,In_685,In_30);
nor U470 (N_470,In_608,In_145);
nor U471 (N_471,In_493,In_582);
nor U472 (N_472,In_575,In_140);
or U473 (N_473,In_657,In_483);
or U474 (N_474,In_596,In_492);
nand U475 (N_475,In_408,In_103);
or U476 (N_476,In_458,In_742);
and U477 (N_477,In_613,In_618);
nand U478 (N_478,In_288,In_364);
and U479 (N_479,In_444,In_212);
nand U480 (N_480,In_742,In_603);
nand U481 (N_481,In_640,In_274);
nor U482 (N_482,In_326,In_270);
nor U483 (N_483,In_276,In_581);
nand U484 (N_484,In_674,In_384);
or U485 (N_485,In_180,In_749);
or U486 (N_486,In_299,In_464);
or U487 (N_487,In_187,In_642);
and U488 (N_488,In_555,In_680);
and U489 (N_489,In_302,In_481);
nor U490 (N_490,In_125,In_122);
nand U491 (N_491,In_365,In_381);
nor U492 (N_492,In_437,In_241);
nor U493 (N_493,In_468,In_366);
nor U494 (N_494,In_289,In_1);
and U495 (N_495,In_34,In_127);
and U496 (N_496,In_558,In_222);
nand U497 (N_497,In_355,In_249);
nand U498 (N_498,In_331,In_105);
or U499 (N_499,In_612,In_552);
nor U500 (N_500,In_342,In_138);
or U501 (N_501,In_672,In_597);
and U502 (N_502,In_215,In_202);
nor U503 (N_503,In_143,In_374);
or U504 (N_504,In_581,In_738);
nand U505 (N_505,In_633,In_399);
nand U506 (N_506,In_339,In_408);
nor U507 (N_507,In_64,In_196);
or U508 (N_508,In_227,In_618);
or U509 (N_509,In_132,In_579);
and U510 (N_510,In_22,In_108);
nor U511 (N_511,In_21,In_599);
and U512 (N_512,In_612,In_202);
nor U513 (N_513,In_474,In_708);
nand U514 (N_514,In_664,In_413);
and U515 (N_515,In_142,In_614);
and U516 (N_516,In_555,In_35);
nand U517 (N_517,In_36,In_419);
and U518 (N_518,In_151,In_563);
xnor U519 (N_519,In_254,In_390);
or U520 (N_520,In_643,In_82);
and U521 (N_521,In_657,In_284);
or U522 (N_522,In_51,In_448);
or U523 (N_523,In_220,In_154);
nor U524 (N_524,In_539,In_247);
or U525 (N_525,In_96,In_44);
and U526 (N_526,In_44,In_449);
nor U527 (N_527,In_457,In_122);
nor U528 (N_528,In_739,In_601);
nand U529 (N_529,In_253,In_207);
nor U530 (N_530,In_392,In_617);
nand U531 (N_531,In_160,In_668);
xor U532 (N_532,In_104,In_736);
and U533 (N_533,In_529,In_679);
and U534 (N_534,In_427,In_582);
nor U535 (N_535,In_694,In_325);
or U536 (N_536,In_699,In_228);
or U537 (N_537,In_345,In_30);
nand U538 (N_538,In_466,In_590);
nand U539 (N_539,In_292,In_239);
or U540 (N_540,In_323,In_427);
and U541 (N_541,In_491,In_143);
or U542 (N_542,In_706,In_333);
nor U543 (N_543,In_658,In_732);
nor U544 (N_544,In_667,In_394);
nor U545 (N_545,In_80,In_662);
or U546 (N_546,In_417,In_561);
or U547 (N_547,In_321,In_71);
nor U548 (N_548,In_287,In_472);
nand U549 (N_549,In_521,In_182);
nor U550 (N_550,In_83,In_739);
nor U551 (N_551,In_64,In_434);
nor U552 (N_552,In_174,In_430);
or U553 (N_553,In_482,In_511);
nand U554 (N_554,In_731,In_212);
and U555 (N_555,In_554,In_700);
nand U556 (N_556,In_90,In_68);
nor U557 (N_557,In_121,In_275);
and U558 (N_558,In_5,In_645);
and U559 (N_559,In_391,In_543);
nor U560 (N_560,In_445,In_744);
nor U561 (N_561,In_401,In_704);
and U562 (N_562,In_559,In_63);
or U563 (N_563,In_1,In_705);
nor U564 (N_564,In_182,In_354);
nand U565 (N_565,In_539,In_648);
nor U566 (N_566,In_735,In_358);
nand U567 (N_567,In_101,In_620);
and U568 (N_568,In_211,In_204);
or U569 (N_569,In_710,In_401);
nand U570 (N_570,In_516,In_221);
and U571 (N_571,In_351,In_738);
nor U572 (N_572,In_136,In_543);
nand U573 (N_573,In_674,In_234);
nor U574 (N_574,In_244,In_709);
or U575 (N_575,In_566,In_24);
or U576 (N_576,In_75,In_69);
and U577 (N_577,In_127,In_148);
or U578 (N_578,In_443,In_195);
or U579 (N_579,In_387,In_511);
nor U580 (N_580,In_9,In_700);
and U581 (N_581,In_349,In_560);
nand U582 (N_582,In_170,In_210);
nand U583 (N_583,In_614,In_18);
nor U584 (N_584,In_367,In_343);
and U585 (N_585,In_665,In_689);
and U586 (N_586,In_153,In_283);
nor U587 (N_587,In_743,In_91);
nand U588 (N_588,In_76,In_301);
and U589 (N_589,In_293,In_635);
nor U590 (N_590,In_371,In_346);
nor U591 (N_591,In_151,In_386);
or U592 (N_592,In_172,In_289);
nor U593 (N_593,In_592,In_704);
nor U594 (N_594,In_677,In_579);
nand U595 (N_595,In_246,In_283);
nand U596 (N_596,In_692,In_209);
and U597 (N_597,In_332,In_351);
nor U598 (N_598,In_643,In_514);
or U599 (N_599,In_179,In_546);
xor U600 (N_600,In_447,In_252);
or U601 (N_601,In_391,In_719);
and U602 (N_602,In_279,In_613);
nand U603 (N_603,In_511,In_117);
nor U604 (N_604,In_143,In_286);
nor U605 (N_605,In_38,In_544);
or U606 (N_606,In_185,In_271);
nand U607 (N_607,In_201,In_349);
nor U608 (N_608,In_502,In_223);
and U609 (N_609,In_132,In_400);
nand U610 (N_610,In_588,In_57);
or U611 (N_611,In_340,In_137);
nand U612 (N_612,In_623,In_610);
nand U613 (N_613,In_475,In_339);
nor U614 (N_614,In_263,In_579);
or U615 (N_615,In_178,In_128);
or U616 (N_616,In_127,In_561);
and U617 (N_617,In_535,In_200);
or U618 (N_618,In_608,In_228);
and U619 (N_619,In_432,In_435);
and U620 (N_620,In_657,In_727);
or U621 (N_621,In_748,In_147);
nand U622 (N_622,In_53,In_297);
nand U623 (N_623,In_10,In_283);
and U624 (N_624,In_411,In_448);
and U625 (N_625,In_302,In_606);
or U626 (N_626,In_65,In_178);
nand U627 (N_627,In_500,In_175);
or U628 (N_628,In_100,In_305);
nand U629 (N_629,In_71,In_534);
or U630 (N_630,In_554,In_716);
and U631 (N_631,In_195,In_410);
nor U632 (N_632,In_461,In_722);
nand U633 (N_633,In_279,In_667);
and U634 (N_634,In_251,In_355);
nor U635 (N_635,In_8,In_673);
or U636 (N_636,In_145,In_722);
and U637 (N_637,In_178,In_511);
nand U638 (N_638,In_70,In_536);
nor U639 (N_639,In_100,In_230);
or U640 (N_640,In_566,In_279);
and U641 (N_641,In_732,In_333);
and U642 (N_642,In_657,In_45);
nor U643 (N_643,In_249,In_443);
nand U644 (N_644,In_204,In_704);
or U645 (N_645,In_501,In_631);
or U646 (N_646,In_357,In_545);
and U647 (N_647,In_97,In_25);
nand U648 (N_648,In_479,In_101);
nand U649 (N_649,In_160,In_60);
nand U650 (N_650,In_672,In_609);
nand U651 (N_651,In_622,In_88);
and U652 (N_652,In_353,In_671);
nor U653 (N_653,In_518,In_737);
and U654 (N_654,In_549,In_502);
and U655 (N_655,In_106,In_220);
nand U656 (N_656,In_231,In_374);
or U657 (N_657,In_108,In_732);
nor U658 (N_658,In_91,In_367);
nand U659 (N_659,In_185,In_317);
nand U660 (N_660,In_186,In_694);
nor U661 (N_661,In_48,In_505);
and U662 (N_662,In_520,In_590);
xnor U663 (N_663,In_740,In_341);
or U664 (N_664,In_216,In_395);
or U665 (N_665,In_747,In_211);
nor U666 (N_666,In_608,In_287);
or U667 (N_667,In_72,In_741);
nor U668 (N_668,In_353,In_735);
nand U669 (N_669,In_261,In_93);
or U670 (N_670,In_691,In_649);
and U671 (N_671,In_700,In_365);
or U672 (N_672,In_602,In_437);
nand U673 (N_673,In_72,In_33);
xor U674 (N_674,In_417,In_497);
or U675 (N_675,In_17,In_171);
nor U676 (N_676,In_300,In_2);
nor U677 (N_677,In_596,In_641);
nand U678 (N_678,In_451,In_358);
nand U679 (N_679,In_39,In_698);
and U680 (N_680,In_29,In_484);
or U681 (N_681,In_104,In_111);
nor U682 (N_682,In_181,In_185);
nand U683 (N_683,In_688,In_144);
and U684 (N_684,In_703,In_11);
and U685 (N_685,In_63,In_499);
or U686 (N_686,In_406,In_634);
nor U687 (N_687,In_240,In_72);
nand U688 (N_688,In_384,In_363);
and U689 (N_689,In_235,In_67);
nor U690 (N_690,In_486,In_239);
nor U691 (N_691,In_415,In_419);
nand U692 (N_692,In_163,In_365);
or U693 (N_693,In_730,In_420);
nor U694 (N_694,In_349,In_323);
nor U695 (N_695,In_701,In_0);
nor U696 (N_696,In_83,In_401);
and U697 (N_697,In_515,In_596);
and U698 (N_698,In_405,In_505);
nor U699 (N_699,In_368,In_551);
nor U700 (N_700,In_220,In_645);
nand U701 (N_701,In_601,In_244);
and U702 (N_702,In_707,In_672);
nor U703 (N_703,In_69,In_239);
and U704 (N_704,In_687,In_576);
and U705 (N_705,In_145,In_495);
or U706 (N_706,In_168,In_364);
or U707 (N_707,In_165,In_249);
and U708 (N_708,In_279,In_212);
nand U709 (N_709,In_205,In_229);
nand U710 (N_710,In_549,In_459);
nand U711 (N_711,In_312,In_5);
nor U712 (N_712,In_371,In_109);
nor U713 (N_713,In_235,In_374);
xnor U714 (N_714,In_745,In_376);
nand U715 (N_715,In_83,In_382);
and U716 (N_716,In_749,In_51);
nor U717 (N_717,In_25,In_585);
and U718 (N_718,In_508,In_322);
xor U719 (N_719,In_97,In_291);
or U720 (N_720,In_119,In_138);
nand U721 (N_721,In_17,In_277);
or U722 (N_722,In_0,In_662);
nand U723 (N_723,In_559,In_383);
and U724 (N_724,In_457,In_682);
nor U725 (N_725,In_667,In_661);
nor U726 (N_726,In_426,In_56);
nor U727 (N_727,In_314,In_359);
or U728 (N_728,In_70,In_187);
nor U729 (N_729,In_222,In_597);
nand U730 (N_730,In_384,In_270);
nand U731 (N_731,In_490,In_38);
nor U732 (N_732,In_719,In_403);
and U733 (N_733,In_422,In_368);
and U734 (N_734,In_437,In_576);
nor U735 (N_735,In_579,In_210);
nor U736 (N_736,In_615,In_1);
nor U737 (N_737,In_355,In_158);
and U738 (N_738,In_279,In_225);
and U739 (N_739,In_185,In_210);
or U740 (N_740,In_585,In_345);
and U741 (N_741,In_341,In_48);
nor U742 (N_742,In_392,In_281);
nand U743 (N_743,In_520,In_503);
or U744 (N_744,In_68,In_257);
or U745 (N_745,In_126,In_424);
nand U746 (N_746,In_728,In_558);
xnor U747 (N_747,In_124,In_630);
nand U748 (N_748,In_677,In_530);
and U749 (N_749,In_20,In_292);
nor U750 (N_750,In_297,In_82);
and U751 (N_751,In_638,In_61);
and U752 (N_752,In_244,In_266);
nor U753 (N_753,In_293,In_745);
and U754 (N_754,In_500,In_718);
or U755 (N_755,In_384,In_562);
nand U756 (N_756,In_642,In_560);
and U757 (N_757,In_165,In_48);
nand U758 (N_758,In_74,In_584);
or U759 (N_759,In_119,In_528);
or U760 (N_760,In_638,In_137);
nor U761 (N_761,In_31,In_723);
or U762 (N_762,In_86,In_230);
nor U763 (N_763,In_559,In_281);
nor U764 (N_764,In_519,In_38);
and U765 (N_765,In_693,In_96);
and U766 (N_766,In_42,In_481);
and U767 (N_767,In_656,In_359);
nor U768 (N_768,In_487,In_634);
nor U769 (N_769,In_2,In_381);
and U770 (N_770,In_554,In_615);
and U771 (N_771,In_275,In_4);
nor U772 (N_772,In_262,In_400);
nor U773 (N_773,In_174,In_577);
and U774 (N_774,In_695,In_376);
or U775 (N_775,In_604,In_642);
nand U776 (N_776,In_132,In_37);
and U777 (N_777,In_160,In_650);
nand U778 (N_778,In_150,In_615);
nor U779 (N_779,In_35,In_669);
or U780 (N_780,In_232,In_457);
nand U781 (N_781,In_590,In_446);
nor U782 (N_782,In_166,In_390);
or U783 (N_783,In_456,In_181);
and U784 (N_784,In_673,In_58);
and U785 (N_785,In_586,In_583);
or U786 (N_786,In_723,In_577);
nand U787 (N_787,In_574,In_453);
or U788 (N_788,In_22,In_585);
nand U789 (N_789,In_465,In_212);
nand U790 (N_790,In_720,In_646);
nor U791 (N_791,In_528,In_737);
nor U792 (N_792,In_407,In_344);
or U793 (N_793,In_35,In_126);
or U794 (N_794,In_242,In_650);
and U795 (N_795,In_505,In_360);
and U796 (N_796,In_56,In_429);
and U797 (N_797,In_112,In_570);
nor U798 (N_798,In_110,In_568);
nor U799 (N_799,In_95,In_546);
nand U800 (N_800,In_503,In_15);
or U801 (N_801,In_611,In_437);
and U802 (N_802,In_151,In_698);
and U803 (N_803,In_732,In_11);
nand U804 (N_804,In_473,In_317);
or U805 (N_805,In_128,In_236);
nand U806 (N_806,In_313,In_629);
nand U807 (N_807,In_517,In_325);
nor U808 (N_808,In_384,In_732);
or U809 (N_809,In_577,In_528);
nor U810 (N_810,In_217,In_565);
nand U811 (N_811,In_202,In_444);
nand U812 (N_812,In_433,In_163);
or U813 (N_813,In_402,In_364);
nor U814 (N_814,In_408,In_727);
nor U815 (N_815,In_45,In_81);
and U816 (N_816,In_508,In_664);
nand U817 (N_817,In_536,In_57);
nor U818 (N_818,In_375,In_487);
nor U819 (N_819,In_335,In_628);
nor U820 (N_820,In_30,In_553);
nand U821 (N_821,In_645,In_558);
or U822 (N_822,In_59,In_417);
and U823 (N_823,In_137,In_584);
and U824 (N_824,In_299,In_373);
or U825 (N_825,In_469,In_442);
and U826 (N_826,In_703,In_65);
and U827 (N_827,In_92,In_219);
nor U828 (N_828,In_366,In_152);
nor U829 (N_829,In_75,In_35);
or U830 (N_830,In_563,In_283);
nand U831 (N_831,In_216,In_517);
and U832 (N_832,In_614,In_16);
nor U833 (N_833,In_531,In_14);
or U834 (N_834,In_13,In_217);
or U835 (N_835,In_374,In_17);
or U836 (N_836,In_568,In_501);
and U837 (N_837,In_597,In_471);
nand U838 (N_838,In_327,In_574);
xor U839 (N_839,In_742,In_651);
nand U840 (N_840,In_645,In_639);
or U841 (N_841,In_698,In_302);
and U842 (N_842,In_163,In_84);
or U843 (N_843,In_59,In_163);
nand U844 (N_844,In_182,In_359);
nor U845 (N_845,In_743,In_331);
nand U846 (N_846,In_65,In_256);
nor U847 (N_847,In_530,In_680);
or U848 (N_848,In_388,In_725);
nor U849 (N_849,In_700,In_212);
and U850 (N_850,In_724,In_697);
nand U851 (N_851,In_730,In_155);
nor U852 (N_852,In_499,In_371);
and U853 (N_853,In_512,In_593);
and U854 (N_854,In_629,In_474);
or U855 (N_855,In_442,In_327);
nand U856 (N_856,In_204,In_162);
and U857 (N_857,In_36,In_617);
nor U858 (N_858,In_208,In_457);
and U859 (N_859,In_297,In_400);
and U860 (N_860,In_114,In_161);
nor U861 (N_861,In_459,In_545);
or U862 (N_862,In_156,In_523);
nand U863 (N_863,In_476,In_494);
and U864 (N_864,In_476,In_75);
or U865 (N_865,In_668,In_372);
or U866 (N_866,In_62,In_272);
nor U867 (N_867,In_238,In_48);
xnor U868 (N_868,In_481,In_231);
nand U869 (N_869,In_414,In_569);
nand U870 (N_870,In_532,In_126);
nand U871 (N_871,In_434,In_511);
and U872 (N_872,In_350,In_662);
and U873 (N_873,In_673,In_53);
or U874 (N_874,In_321,In_686);
nand U875 (N_875,In_540,In_473);
nor U876 (N_876,In_346,In_67);
or U877 (N_877,In_85,In_388);
nor U878 (N_878,In_464,In_627);
nand U879 (N_879,In_574,In_70);
and U880 (N_880,In_669,In_362);
or U881 (N_881,In_95,In_43);
and U882 (N_882,In_730,In_564);
xnor U883 (N_883,In_210,In_118);
or U884 (N_884,In_70,In_682);
or U885 (N_885,In_88,In_81);
or U886 (N_886,In_362,In_170);
and U887 (N_887,In_737,In_360);
and U888 (N_888,In_590,In_668);
nand U889 (N_889,In_702,In_609);
nand U890 (N_890,In_499,In_318);
or U891 (N_891,In_397,In_134);
nor U892 (N_892,In_30,In_744);
nand U893 (N_893,In_440,In_575);
and U894 (N_894,In_654,In_452);
or U895 (N_895,In_275,In_165);
nor U896 (N_896,In_424,In_519);
and U897 (N_897,In_358,In_27);
or U898 (N_898,In_465,In_681);
nor U899 (N_899,In_523,In_9);
and U900 (N_900,In_502,In_666);
nor U901 (N_901,In_683,In_143);
or U902 (N_902,In_210,In_676);
nor U903 (N_903,In_95,In_296);
nand U904 (N_904,In_743,In_267);
and U905 (N_905,In_387,In_520);
or U906 (N_906,In_5,In_223);
and U907 (N_907,In_23,In_56);
nor U908 (N_908,In_199,In_423);
nand U909 (N_909,In_88,In_318);
and U910 (N_910,In_482,In_544);
xnor U911 (N_911,In_610,In_673);
and U912 (N_912,In_140,In_618);
xor U913 (N_913,In_651,In_227);
nand U914 (N_914,In_617,In_568);
nor U915 (N_915,In_10,In_558);
nor U916 (N_916,In_408,In_591);
and U917 (N_917,In_242,In_160);
nor U918 (N_918,In_611,In_344);
nand U919 (N_919,In_612,In_517);
nand U920 (N_920,In_387,In_119);
or U921 (N_921,In_119,In_5);
nor U922 (N_922,In_706,In_95);
nand U923 (N_923,In_0,In_589);
xnor U924 (N_924,In_692,In_548);
nor U925 (N_925,In_145,In_749);
or U926 (N_926,In_524,In_400);
nor U927 (N_927,In_745,In_307);
xor U928 (N_928,In_712,In_281);
nor U929 (N_929,In_513,In_473);
nand U930 (N_930,In_343,In_80);
and U931 (N_931,In_275,In_510);
and U932 (N_932,In_477,In_317);
nor U933 (N_933,In_114,In_4);
nor U934 (N_934,In_376,In_474);
or U935 (N_935,In_108,In_408);
xor U936 (N_936,In_22,In_58);
nand U937 (N_937,In_174,In_61);
and U938 (N_938,In_736,In_340);
xnor U939 (N_939,In_539,In_198);
or U940 (N_940,In_218,In_528);
and U941 (N_941,In_505,In_168);
nor U942 (N_942,In_696,In_322);
nand U943 (N_943,In_397,In_107);
or U944 (N_944,In_20,In_438);
and U945 (N_945,In_315,In_612);
and U946 (N_946,In_237,In_642);
nand U947 (N_947,In_465,In_307);
or U948 (N_948,In_666,In_739);
nand U949 (N_949,In_571,In_274);
xor U950 (N_950,In_301,In_214);
or U951 (N_951,In_263,In_517);
nor U952 (N_952,In_251,In_260);
nand U953 (N_953,In_287,In_435);
or U954 (N_954,In_70,In_108);
xnor U955 (N_955,In_472,In_291);
nor U956 (N_956,In_79,In_235);
xor U957 (N_957,In_274,In_337);
nand U958 (N_958,In_326,In_6);
or U959 (N_959,In_474,In_71);
nor U960 (N_960,In_627,In_458);
and U961 (N_961,In_89,In_691);
and U962 (N_962,In_431,In_460);
or U963 (N_963,In_334,In_336);
and U964 (N_964,In_118,In_182);
and U965 (N_965,In_312,In_245);
nor U966 (N_966,In_557,In_371);
nor U967 (N_967,In_705,In_183);
nand U968 (N_968,In_565,In_409);
and U969 (N_969,In_676,In_75);
and U970 (N_970,In_151,In_124);
and U971 (N_971,In_144,In_109);
nand U972 (N_972,In_84,In_667);
and U973 (N_973,In_398,In_500);
xnor U974 (N_974,In_386,In_493);
nor U975 (N_975,In_677,In_151);
nand U976 (N_976,In_361,In_461);
nand U977 (N_977,In_711,In_450);
and U978 (N_978,In_708,In_502);
or U979 (N_979,In_6,In_638);
nand U980 (N_980,In_85,In_741);
xor U981 (N_981,In_564,In_593);
and U982 (N_982,In_171,In_18);
or U983 (N_983,In_236,In_92);
or U984 (N_984,In_229,In_335);
and U985 (N_985,In_299,In_629);
or U986 (N_986,In_122,In_591);
nor U987 (N_987,In_350,In_254);
nor U988 (N_988,In_71,In_59);
nor U989 (N_989,In_712,In_570);
or U990 (N_990,In_652,In_357);
nand U991 (N_991,In_56,In_213);
xnor U992 (N_992,In_706,In_33);
and U993 (N_993,In_529,In_218);
and U994 (N_994,In_665,In_621);
or U995 (N_995,In_104,In_194);
or U996 (N_996,In_404,In_481);
and U997 (N_997,In_545,In_74);
nor U998 (N_998,In_23,In_317);
nand U999 (N_999,In_294,In_246);
nor U1000 (N_1000,In_463,In_253);
and U1001 (N_1001,In_353,In_243);
nor U1002 (N_1002,In_447,In_564);
and U1003 (N_1003,In_641,In_438);
nor U1004 (N_1004,In_595,In_419);
and U1005 (N_1005,In_259,In_386);
nor U1006 (N_1006,In_579,In_530);
or U1007 (N_1007,In_236,In_170);
and U1008 (N_1008,In_696,In_248);
or U1009 (N_1009,In_179,In_708);
or U1010 (N_1010,In_439,In_733);
and U1011 (N_1011,In_511,In_646);
or U1012 (N_1012,In_746,In_175);
nand U1013 (N_1013,In_124,In_301);
nor U1014 (N_1014,In_502,In_67);
and U1015 (N_1015,In_658,In_505);
nand U1016 (N_1016,In_639,In_214);
and U1017 (N_1017,In_653,In_547);
nor U1018 (N_1018,In_368,In_549);
nand U1019 (N_1019,In_449,In_144);
nand U1020 (N_1020,In_719,In_431);
nand U1021 (N_1021,In_651,In_581);
or U1022 (N_1022,In_687,In_81);
or U1023 (N_1023,In_622,In_22);
nor U1024 (N_1024,In_202,In_222);
nand U1025 (N_1025,In_642,In_539);
and U1026 (N_1026,In_278,In_103);
or U1027 (N_1027,In_417,In_81);
and U1028 (N_1028,In_373,In_642);
nand U1029 (N_1029,In_734,In_525);
nand U1030 (N_1030,In_602,In_137);
or U1031 (N_1031,In_103,In_247);
and U1032 (N_1032,In_701,In_22);
and U1033 (N_1033,In_236,In_169);
nor U1034 (N_1034,In_96,In_500);
nor U1035 (N_1035,In_465,In_155);
or U1036 (N_1036,In_536,In_447);
nand U1037 (N_1037,In_260,In_286);
nand U1038 (N_1038,In_667,In_507);
and U1039 (N_1039,In_109,In_589);
or U1040 (N_1040,In_729,In_407);
nor U1041 (N_1041,In_747,In_264);
and U1042 (N_1042,In_465,In_310);
nand U1043 (N_1043,In_436,In_197);
or U1044 (N_1044,In_234,In_694);
or U1045 (N_1045,In_690,In_727);
or U1046 (N_1046,In_642,In_162);
and U1047 (N_1047,In_245,In_48);
or U1048 (N_1048,In_516,In_150);
xnor U1049 (N_1049,In_235,In_60);
nand U1050 (N_1050,In_420,In_98);
nand U1051 (N_1051,In_43,In_435);
and U1052 (N_1052,In_739,In_253);
and U1053 (N_1053,In_674,In_476);
or U1054 (N_1054,In_371,In_694);
and U1055 (N_1055,In_139,In_280);
and U1056 (N_1056,In_190,In_141);
and U1057 (N_1057,In_687,In_481);
nor U1058 (N_1058,In_18,In_57);
nor U1059 (N_1059,In_386,In_36);
nand U1060 (N_1060,In_81,In_610);
nor U1061 (N_1061,In_405,In_238);
nor U1062 (N_1062,In_320,In_231);
nor U1063 (N_1063,In_194,In_282);
nand U1064 (N_1064,In_547,In_631);
and U1065 (N_1065,In_599,In_600);
nand U1066 (N_1066,In_313,In_576);
nor U1067 (N_1067,In_6,In_660);
nand U1068 (N_1068,In_724,In_731);
nand U1069 (N_1069,In_703,In_2);
or U1070 (N_1070,In_721,In_430);
nor U1071 (N_1071,In_583,In_217);
nand U1072 (N_1072,In_441,In_284);
nand U1073 (N_1073,In_101,In_264);
nor U1074 (N_1074,In_460,In_68);
nor U1075 (N_1075,In_553,In_419);
and U1076 (N_1076,In_160,In_53);
nor U1077 (N_1077,In_433,In_43);
or U1078 (N_1078,In_332,In_324);
and U1079 (N_1079,In_659,In_534);
nor U1080 (N_1080,In_350,In_482);
and U1081 (N_1081,In_195,In_625);
and U1082 (N_1082,In_19,In_208);
or U1083 (N_1083,In_101,In_200);
or U1084 (N_1084,In_416,In_228);
and U1085 (N_1085,In_120,In_87);
or U1086 (N_1086,In_534,In_494);
and U1087 (N_1087,In_7,In_422);
and U1088 (N_1088,In_296,In_702);
nand U1089 (N_1089,In_57,In_606);
or U1090 (N_1090,In_113,In_690);
nor U1091 (N_1091,In_742,In_714);
nor U1092 (N_1092,In_279,In_425);
nor U1093 (N_1093,In_366,In_456);
nand U1094 (N_1094,In_274,In_81);
nor U1095 (N_1095,In_272,In_371);
nor U1096 (N_1096,In_131,In_180);
and U1097 (N_1097,In_422,In_726);
or U1098 (N_1098,In_389,In_102);
and U1099 (N_1099,In_466,In_68);
nor U1100 (N_1100,In_392,In_660);
and U1101 (N_1101,In_451,In_638);
nand U1102 (N_1102,In_69,In_95);
nor U1103 (N_1103,In_57,In_22);
or U1104 (N_1104,In_570,In_385);
nor U1105 (N_1105,In_598,In_512);
xnor U1106 (N_1106,In_290,In_334);
nor U1107 (N_1107,In_277,In_304);
and U1108 (N_1108,In_448,In_516);
nor U1109 (N_1109,In_309,In_406);
nor U1110 (N_1110,In_472,In_630);
nor U1111 (N_1111,In_304,In_345);
nor U1112 (N_1112,In_182,In_464);
or U1113 (N_1113,In_603,In_507);
nand U1114 (N_1114,In_698,In_44);
and U1115 (N_1115,In_661,In_416);
and U1116 (N_1116,In_382,In_461);
nor U1117 (N_1117,In_502,In_80);
and U1118 (N_1118,In_185,In_465);
and U1119 (N_1119,In_229,In_574);
or U1120 (N_1120,In_152,In_429);
or U1121 (N_1121,In_641,In_458);
or U1122 (N_1122,In_740,In_327);
or U1123 (N_1123,In_356,In_163);
and U1124 (N_1124,In_225,In_421);
and U1125 (N_1125,In_723,In_41);
and U1126 (N_1126,In_34,In_126);
and U1127 (N_1127,In_524,In_67);
nor U1128 (N_1128,In_192,In_551);
xor U1129 (N_1129,In_95,In_611);
and U1130 (N_1130,In_95,In_405);
nand U1131 (N_1131,In_510,In_660);
nor U1132 (N_1132,In_114,In_207);
nand U1133 (N_1133,In_537,In_641);
or U1134 (N_1134,In_577,In_223);
and U1135 (N_1135,In_329,In_594);
xnor U1136 (N_1136,In_157,In_698);
and U1137 (N_1137,In_292,In_250);
and U1138 (N_1138,In_590,In_421);
nand U1139 (N_1139,In_318,In_311);
or U1140 (N_1140,In_303,In_209);
nand U1141 (N_1141,In_102,In_709);
and U1142 (N_1142,In_164,In_74);
nor U1143 (N_1143,In_10,In_243);
nand U1144 (N_1144,In_146,In_261);
and U1145 (N_1145,In_641,In_276);
or U1146 (N_1146,In_241,In_418);
or U1147 (N_1147,In_659,In_2);
nor U1148 (N_1148,In_353,In_286);
nor U1149 (N_1149,In_113,In_49);
nand U1150 (N_1150,In_500,In_682);
nand U1151 (N_1151,In_132,In_321);
xnor U1152 (N_1152,In_579,In_101);
and U1153 (N_1153,In_307,In_515);
or U1154 (N_1154,In_484,In_306);
nor U1155 (N_1155,In_543,In_278);
nand U1156 (N_1156,In_510,In_274);
and U1157 (N_1157,In_2,In_366);
or U1158 (N_1158,In_671,In_229);
nand U1159 (N_1159,In_391,In_519);
and U1160 (N_1160,In_240,In_199);
and U1161 (N_1161,In_436,In_159);
xnor U1162 (N_1162,In_251,In_673);
nor U1163 (N_1163,In_530,In_19);
nand U1164 (N_1164,In_478,In_217);
nand U1165 (N_1165,In_558,In_398);
or U1166 (N_1166,In_89,In_659);
or U1167 (N_1167,In_479,In_525);
and U1168 (N_1168,In_467,In_156);
nand U1169 (N_1169,In_144,In_76);
nand U1170 (N_1170,In_307,In_529);
and U1171 (N_1171,In_436,In_48);
nor U1172 (N_1172,In_340,In_249);
and U1173 (N_1173,In_264,In_219);
nor U1174 (N_1174,In_364,In_109);
and U1175 (N_1175,In_578,In_87);
nor U1176 (N_1176,In_312,In_573);
nor U1177 (N_1177,In_375,In_497);
nor U1178 (N_1178,In_687,In_295);
or U1179 (N_1179,In_588,In_648);
nor U1180 (N_1180,In_27,In_2);
nor U1181 (N_1181,In_59,In_604);
nand U1182 (N_1182,In_144,In_413);
nand U1183 (N_1183,In_626,In_128);
nand U1184 (N_1184,In_149,In_506);
or U1185 (N_1185,In_535,In_581);
nand U1186 (N_1186,In_53,In_504);
and U1187 (N_1187,In_85,In_3);
nor U1188 (N_1188,In_655,In_629);
and U1189 (N_1189,In_561,In_183);
or U1190 (N_1190,In_362,In_272);
nand U1191 (N_1191,In_499,In_600);
or U1192 (N_1192,In_206,In_745);
nand U1193 (N_1193,In_673,In_638);
nor U1194 (N_1194,In_215,In_440);
nor U1195 (N_1195,In_81,In_501);
or U1196 (N_1196,In_295,In_595);
nor U1197 (N_1197,In_175,In_532);
nand U1198 (N_1198,In_575,In_652);
nand U1199 (N_1199,In_642,In_643);
nand U1200 (N_1200,In_449,In_276);
or U1201 (N_1201,In_160,In_121);
nand U1202 (N_1202,In_328,In_47);
nand U1203 (N_1203,In_582,In_109);
nand U1204 (N_1204,In_457,In_108);
and U1205 (N_1205,In_12,In_67);
or U1206 (N_1206,In_513,In_533);
or U1207 (N_1207,In_176,In_163);
nor U1208 (N_1208,In_98,In_307);
nand U1209 (N_1209,In_536,In_450);
and U1210 (N_1210,In_508,In_385);
or U1211 (N_1211,In_602,In_127);
and U1212 (N_1212,In_187,In_335);
and U1213 (N_1213,In_658,In_502);
nand U1214 (N_1214,In_104,In_471);
nor U1215 (N_1215,In_624,In_249);
nor U1216 (N_1216,In_640,In_318);
or U1217 (N_1217,In_558,In_740);
and U1218 (N_1218,In_631,In_219);
nor U1219 (N_1219,In_62,In_442);
nor U1220 (N_1220,In_686,In_639);
and U1221 (N_1221,In_276,In_231);
nor U1222 (N_1222,In_579,In_206);
nand U1223 (N_1223,In_495,In_466);
and U1224 (N_1224,In_299,In_493);
nand U1225 (N_1225,In_547,In_150);
nor U1226 (N_1226,In_609,In_100);
or U1227 (N_1227,In_409,In_632);
nand U1228 (N_1228,In_635,In_20);
nand U1229 (N_1229,In_570,In_244);
nor U1230 (N_1230,In_388,In_16);
nand U1231 (N_1231,In_374,In_703);
nand U1232 (N_1232,In_727,In_381);
and U1233 (N_1233,In_490,In_36);
and U1234 (N_1234,In_145,In_598);
or U1235 (N_1235,In_72,In_253);
nor U1236 (N_1236,In_718,In_668);
and U1237 (N_1237,In_232,In_555);
or U1238 (N_1238,In_686,In_4);
and U1239 (N_1239,In_719,In_333);
and U1240 (N_1240,In_718,In_107);
xor U1241 (N_1241,In_686,In_230);
or U1242 (N_1242,In_174,In_336);
nor U1243 (N_1243,In_363,In_420);
nand U1244 (N_1244,In_302,In_294);
nor U1245 (N_1245,In_535,In_2);
and U1246 (N_1246,In_640,In_261);
or U1247 (N_1247,In_734,In_378);
nor U1248 (N_1248,In_746,In_732);
nand U1249 (N_1249,In_502,In_438);
nor U1250 (N_1250,In_484,In_520);
nand U1251 (N_1251,In_560,In_657);
or U1252 (N_1252,In_297,In_552);
xor U1253 (N_1253,In_169,In_574);
and U1254 (N_1254,In_713,In_551);
nand U1255 (N_1255,In_339,In_197);
and U1256 (N_1256,In_232,In_441);
and U1257 (N_1257,In_192,In_672);
nor U1258 (N_1258,In_302,In_675);
nor U1259 (N_1259,In_69,In_138);
or U1260 (N_1260,In_677,In_551);
nand U1261 (N_1261,In_153,In_390);
nor U1262 (N_1262,In_246,In_547);
nor U1263 (N_1263,In_732,In_233);
and U1264 (N_1264,In_449,In_133);
nand U1265 (N_1265,In_447,In_678);
or U1266 (N_1266,In_157,In_222);
or U1267 (N_1267,In_367,In_674);
nand U1268 (N_1268,In_110,In_692);
or U1269 (N_1269,In_180,In_714);
and U1270 (N_1270,In_141,In_494);
nor U1271 (N_1271,In_726,In_340);
nor U1272 (N_1272,In_691,In_669);
or U1273 (N_1273,In_234,In_375);
and U1274 (N_1274,In_683,In_336);
xor U1275 (N_1275,In_380,In_419);
and U1276 (N_1276,In_682,In_621);
nor U1277 (N_1277,In_247,In_173);
and U1278 (N_1278,In_365,In_571);
nor U1279 (N_1279,In_386,In_297);
or U1280 (N_1280,In_141,In_58);
or U1281 (N_1281,In_163,In_109);
nor U1282 (N_1282,In_327,In_429);
or U1283 (N_1283,In_132,In_491);
xnor U1284 (N_1284,In_64,In_12);
nand U1285 (N_1285,In_319,In_532);
nor U1286 (N_1286,In_126,In_616);
xnor U1287 (N_1287,In_113,In_355);
nand U1288 (N_1288,In_290,In_477);
or U1289 (N_1289,In_478,In_205);
and U1290 (N_1290,In_307,In_668);
or U1291 (N_1291,In_173,In_41);
and U1292 (N_1292,In_433,In_231);
nor U1293 (N_1293,In_244,In_461);
xnor U1294 (N_1294,In_0,In_433);
xor U1295 (N_1295,In_367,In_73);
nor U1296 (N_1296,In_716,In_257);
and U1297 (N_1297,In_444,In_140);
nand U1298 (N_1298,In_257,In_487);
nor U1299 (N_1299,In_119,In_656);
nand U1300 (N_1300,In_661,In_223);
nor U1301 (N_1301,In_478,In_37);
nand U1302 (N_1302,In_532,In_8);
and U1303 (N_1303,In_122,In_422);
nor U1304 (N_1304,In_120,In_428);
nor U1305 (N_1305,In_649,In_536);
and U1306 (N_1306,In_138,In_534);
nand U1307 (N_1307,In_658,In_213);
nand U1308 (N_1308,In_643,In_626);
and U1309 (N_1309,In_667,In_309);
or U1310 (N_1310,In_362,In_229);
nor U1311 (N_1311,In_469,In_248);
nand U1312 (N_1312,In_79,In_564);
nand U1313 (N_1313,In_380,In_746);
or U1314 (N_1314,In_173,In_5);
nand U1315 (N_1315,In_144,In_266);
and U1316 (N_1316,In_22,In_273);
nand U1317 (N_1317,In_629,In_265);
nor U1318 (N_1318,In_346,In_263);
and U1319 (N_1319,In_532,In_25);
xnor U1320 (N_1320,In_485,In_481);
or U1321 (N_1321,In_20,In_538);
nor U1322 (N_1322,In_749,In_507);
and U1323 (N_1323,In_66,In_416);
or U1324 (N_1324,In_206,In_120);
or U1325 (N_1325,In_685,In_675);
nand U1326 (N_1326,In_12,In_183);
nor U1327 (N_1327,In_507,In_352);
or U1328 (N_1328,In_175,In_623);
nand U1329 (N_1329,In_749,In_525);
nor U1330 (N_1330,In_122,In_105);
nor U1331 (N_1331,In_242,In_337);
nand U1332 (N_1332,In_554,In_409);
nor U1333 (N_1333,In_253,In_293);
and U1334 (N_1334,In_334,In_248);
nor U1335 (N_1335,In_111,In_231);
nor U1336 (N_1336,In_187,In_51);
nor U1337 (N_1337,In_447,In_514);
nor U1338 (N_1338,In_57,In_708);
and U1339 (N_1339,In_312,In_271);
or U1340 (N_1340,In_702,In_285);
or U1341 (N_1341,In_157,In_278);
and U1342 (N_1342,In_353,In_487);
and U1343 (N_1343,In_377,In_47);
or U1344 (N_1344,In_152,In_551);
nand U1345 (N_1345,In_50,In_387);
and U1346 (N_1346,In_600,In_318);
and U1347 (N_1347,In_264,In_407);
and U1348 (N_1348,In_434,In_325);
and U1349 (N_1349,In_168,In_125);
and U1350 (N_1350,In_372,In_581);
and U1351 (N_1351,In_474,In_515);
nand U1352 (N_1352,In_366,In_494);
and U1353 (N_1353,In_600,In_381);
and U1354 (N_1354,In_467,In_421);
or U1355 (N_1355,In_213,In_221);
and U1356 (N_1356,In_366,In_281);
and U1357 (N_1357,In_583,In_119);
and U1358 (N_1358,In_176,In_178);
and U1359 (N_1359,In_428,In_244);
and U1360 (N_1360,In_65,In_332);
and U1361 (N_1361,In_128,In_517);
and U1362 (N_1362,In_176,In_181);
nor U1363 (N_1363,In_85,In_523);
nor U1364 (N_1364,In_377,In_466);
or U1365 (N_1365,In_204,In_647);
nand U1366 (N_1366,In_431,In_78);
nand U1367 (N_1367,In_316,In_515);
nor U1368 (N_1368,In_428,In_59);
nor U1369 (N_1369,In_450,In_717);
nor U1370 (N_1370,In_374,In_434);
or U1371 (N_1371,In_425,In_189);
nor U1372 (N_1372,In_103,In_487);
and U1373 (N_1373,In_90,In_98);
and U1374 (N_1374,In_125,In_729);
nand U1375 (N_1375,In_328,In_466);
and U1376 (N_1376,In_270,In_703);
nor U1377 (N_1377,In_576,In_429);
and U1378 (N_1378,In_714,In_271);
and U1379 (N_1379,In_400,In_583);
or U1380 (N_1380,In_446,In_222);
nor U1381 (N_1381,In_135,In_720);
or U1382 (N_1382,In_483,In_280);
and U1383 (N_1383,In_728,In_384);
nand U1384 (N_1384,In_246,In_126);
nand U1385 (N_1385,In_330,In_11);
or U1386 (N_1386,In_743,In_272);
nand U1387 (N_1387,In_207,In_438);
or U1388 (N_1388,In_641,In_455);
and U1389 (N_1389,In_38,In_275);
nand U1390 (N_1390,In_277,In_259);
or U1391 (N_1391,In_133,In_233);
or U1392 (N_1392,In_22,In_364);
or U1393 (N_1393,In_629,In_628);
or U1394 (N_1394,In_693,In_643);
or U1395 (N_1395,In_483,In_724);
and U1396 (N_1396,In_167,In_215);
and U1397 (N_1397,In_548,In_555);
nand U1398 (N_1398,In_411,In_531);
nand U1399 (N_1399,In_452,In_122);
nor U1400 (N_1400,In_208,In_299);
nor U1401 (N_1401,In_236,In_289);
or U1402 (N_1402,In_384,In_520);
nor U1403 (N_1403,In_179,In_633);
nor U1404 (N_1404,In_608,In_94);
or U1405 (N_1405,In_76,In_20);
and U1406 (N_1406,In_672,In_649);
nor U1407 (N_1407,In_648,In_477);
nor U1408 (N_1408,In_580,In_91);
and U1409 (N_1409,In_539,In_685);
or U1410 (N_1410,In_93,In_223);
nor U1411 (N_1411,In_69,In_354);
nor U1412 (N_1412,In_300,In_569);
nand U1413 (N_1413,In_335,In_533);
nand U1414 (N_1414,In_517,In_264);
nand U1415 (N_1415,In_345,In_464);
nand U1416 (N_1416,In_192,In_303);
nor U1417 (N_1417,In_696,In_128);
nor U1418 (N_1418,In_12,In_131);
nor U1419 (N_1419,In_585,In_415);
and U1420 (N_1420,In_699,In_636);
nand U1421 (N_1421,In_708,In_744);
and U1422 (N_1422,In_518,In_461);
xor U1423 (N_1423,In_597,In_80);
nand U1424 (N_1424,In_11,In_354);
or U1425 (N_1425,In_553,In_240);
nor U1426 (N_1426,In_361,In_404);
nor U1427 (N_1427,In_266,In_234);
or U1428 (N_1428,In_707,In_584);
or U1429 (N_1429,In_391,In_136);
nand U1430 (N_1430,In_414,In_675);
or U1431 (N_1431,In_552,In_493);
and U1432 (N_1432,In_220,In_370);
xor U1433 (N_1433,In_460,In_97);
nor U1434 (N_1434,In_571,In_336);
nand U1435 (N_1435,In_644,In_661);
nor U1436 (N_1436,In_93,In_353);
xnor U1437 (N_1437,In_147,In_24);
or U1438 (N_1438,In_714,In_389);
and U1439 (N_1439,In_642,In_749);
nor U1440 (N_1440,In_85,In_578);
nand U1441 (N_1441,In_101,In_688);
and U1442 (N_1442,In_543,In_375);
or U1443 (N_1443,In_265,In_233);
nand U1444 (N_1444,In_211,In_724);
or U1445 (N_1445,In_235,In_694);
or U1446 (N_1446,In_584,In_392);
nor U1447 (N_1447,In_352,In_12);
or U1448 (N_1448,In_312,In_285);
nand U1449 (N_1449,In_565,In_404);
nor U1450 (N_1450,In_161,In_23);
and U1451 (N_1451,In_15,In_275);
and U1452 (N_1452,In_35,In_181);
or U1453 (N_1453,In_41,In_522);
or U1454 (N_1454,In_29,In_572);
nor U1455 (N_1455,In_433,In_150);
nand U1456 (N_1456,In_471,In_440);
or U1457 (N_1457,In_201,In_199);
and U1458 (N_1458,In_493,In_298);
and U1459 (N_1459,In_168,In_78);
nand U1460 (N_1460,In_110,In_355);
nor U1461 (N_1461,In_352,In_739);
nand U1462 (N_1462,In_292,In_654);
nor U1463 (N_1463,In_127,In_529);
and U1464 (N_1464,In_557,In_563);
nand U1465 (N_1465,In_574,In_440);
and U1466 (N_1466,In_706,In_345);
nor U1467 (N_1467,In_211,In_27);
or U1468 (N_1468,In_16,In_217);
or U1469 (N_1469,In_562,In_672);
nor U1470 (N_1470,In_151,In_289);
nand U1471 (N_1471,In_295,In_264);
or U1472 (N_1472,In_131,In_172);
nor U1473 (N_1473,In_658,In_53);
nand U1474 (N_1474,In_580,In_725);
xor U1475 (N_1475,In_529,In_85);
nor U1476 (N_1476,In_748,In_115);
or U1477 (N_1477,In_301,In_638);
and U1478 (N_1478,In_436,In_354);
nand U1479 (N_1479,In_652,In_207);
nor U1480 (N_1480,In_173,In_228);
and U1481 (N_1481,In_410,In_402);
or U1482 (N_1482,In_302,In_433);
or U1483 (N_1483,In_690,In_342);
nor U1484 (N_1484,In_504,In_377);
or U1485 (N_1485,In_52,In_438);
nor U1486 (N_1486,In_70,In_597);
nand U1487 (N_1487,In_91,In_510);
nor U1488 (N_1488,In_315,In_566);
or U1489 (N_1489,In_343,In_402);
and U1490 (N_1490,In_317,In_703);
nand U1491 (N_1491,In_573,In_644);
and U1492 (N_1492,In_682,In_610);
and U1493 (N_1493,In_571,In_591);
and U1494 (N_1494,In_120,In_181);
and U1495 (N_1495,In_149,In_699);
nor U1496 (N_1496,In_402,In_619);
or U1497 (N_1497,In_643,In_638);
nor U1498 (N_1498,In_747,In_543);
and U1499 (N_1499,In_716,In_491);
and U1500 (N_1500,In_412,In_67);
nor U1501 (N_1501,In_573,In_261);
xor U1502 (N_1502,In_535,In_54);
xor U1503 (N_1503,In_248,In_52);
nand U1504 (N_1504,In_78,In_11);
nor U1505 (N_1505,In_502,In_693);
and U1506 (N_1506,In_481,In_466);
nand U1507 (N_1507,In_264,In_57);
or U1508 (N_1508,In_584,In_500);
nor U1509 (N_1509,In_436,In_597);
nor U1510 (N_1510,In_420,In_242);
nor U1511 (N_1511,In_493,In_585);
or U1512 (N_1512,In_549,In_569);
and U1513 (N_1513,In_417,In_358);
nand U1514 (N_1514,In_615,In_465);
and U1515 (N_1515,In_590,In_562);
nor U1516 (N_1516,In_552,In_365);
and U1517 (N_1517,In_465,In_585);
or U1518 (N_1518,In_667,In_216);
nand U1519 (N_1519,In_589,In_486);
nand U1520 (N_1520,In_291,In_50);
nand U1521 (N_1521,In_420,In_590);
xnor U1522 (N_1522,In_158,In_720);
nor U1523 (N_1523,In_240,In_720);
or U1524 (N_1524,In_358,In_619);
or U1525 (N_1525,In_223,In_266);
or U1526 (N_1526,In_213,In_393);
nor U1527 (N_1527,In_450,In_279);
or U1528 (N_1528,In_213,In_405);
nor U1529 (N_1529,In_275,In_183);
and U1530 (N_1530,In_71,In_539);
nor U1531 (N_1531,In_167,In_289);
nand U1532 (N_1532,In_70,In_517);
or U1533 (N_1533,In_661,In_117);
xor U1534 (N_1534,In_167,In_512);
xor U1535 (N_1535,In_327,In_572);
or U1536 (N_1536,In_370,In_627);
and U1537 (N_1537,In_641,In_506);
nor U1538 (N_1538,In_120,In_240);
and U1539 (N_1539,In_128,In_28);
or U1540 (N_1540,In_672,In_352);
or U1541 (N_1541,In_200,In_482);
nand U1542 (N_1542,In_643,In_736);
or U1543 (N_1543,In_679,In_184);
nand U1544 (N_1544,In_322,In_558);
or U1545 (N_1545,In_153,In_53);
nor U1546 (N_1546,In_288,In_331);
or U1547 (N_1547,In_596,In_247);
nand U1548 (N_1548,In_345,In_294);
or U1549 (N_1549,In_200,In_71);
or U1550 (N_1550,In_152,In_175);
and U1551 (N_1551,In_426,In_64);
and U1552 (N_1552,In_546,In_703);
xnor U1553 (N_1553,In_502,In_473);
nand U1554 (N_1554,In_136,In_127);
nor U1555 (N_1555,In_449,In_447);
nor U1556 (N_1556,In_111,In_237);
nand U1557 (N_1557,In_58,In_72);
and U1558 (N_1558,In_186,In_133);
or U1559 (N_1559,In_389,In_166);
nand U1560 (N_1560,In_700,In_243);
or U1561 (N_1561,In_81,In_262);
and U1562 (N_1562,In_21,In_268);
or U1563 (N_1563,In_537,In_663);
or U1564 (N_1564,In_527,In_444);
or U1565 (N_1565,In_20,In_247);
or U1566 (N_1566,In_191,In_97);
or U1567 (N_1567,In_133,In_255);
or U1568 (N_1568,In_237,In_23);
nor U1569 (N_1569,In_111,In_18);
or U1570 (N_1570,In_93,In_530);
or U1571 (N_1571,In_607,In_225);
and U1572 (N_1572,In_493,In_738);
nor U1573 (N_1573,In_91,In_192);
and U1574 (N_1574,In_436,In_644);
nor U1575 (N_1575,In_48,In_570);
nand U1576 (N_1576,In_209,In_733);
nor U1577 (N_1577,In_268,In_543);
and U1578 (N_1578,In_259,In_337);
or U1579 (N_1579,In_159,In_572);
and U1580 (N_1580,In_401,In_546);
nor U1581 (N_1581,In_295,In_540);
and U1582 (N_1582,In_502,In_579);
or U1583 (N_1583,In_561,In_636);
nand U1584 (N_1584,In_698,In_66);
or U1585 (N_1585,In_208,In_726);
or U1586 (N_1586,In_57,In_564);
nor U1587 (N_1587,In_346,In_326);
nand U1588 (N_1588,In_699,In_564);
and U1589 (N_1589,In_576,In_626);
nor U1590 (N_1590,In_672,In_199);
nor U1591 (N_1591,In_675,In_694);
nand U1592 (N_1592,In_313,In_746);
and U1593 (N_1593,In_509,In_391);
and U1594 (N_1594,In_667,In_669);
nand U1595 (N_1595,In_454,In_448);
and U1596 (N_1596,In_631,In_229);
or U1597 (N_1597,In_708,In_716);
and U1598 (N_1598,In_46,In_742);
and U1599 (N_1599,In_17,In_204);
nand U1600 (N_1600,In_184,In_592);
or U1601 (N_1601,In_225,In_238);
or U1602 (N_1602,In_271,In_349);
and U1603 (N_1603,In_219,In_490);
or U1604 (N_1604,In_385,In_88);
nand U1605 (N_1605,In_583,In_163);
or U1606 (N_1606,In_327,In_392);
and U1607 (N_1607,In_335,In_733);
or U1608 (N_1608,In_320,In_272);
and U1609 (N_1609,In_6,In_265);
and U1610 (N_1610,In_437,In_619);
and U1611 (N_1611,In_289,In_499);
nor U1612 (N_1612,In_419,In_414);
nand U1613 (N_1613,In_70,In_162);
or U1614 (N_1614,In_29,In_267);
or U1615 (N_1615,In_332,In_674);
nor U1616 (N_1616,In_307,In_703);
or U1617 (N_1617,In_558,In_442);
and U1618 (N_1618,In_307,In_285);
and U1619 (N_1619,In_654,In_239);
nor U1620 (N_1620,In_235,In_578);
and U1621 (N_1621,In_386,In_79);
and U1622 (N_1622,In_315,In_141);
and U1623 (N_1623,In_253,In_94);
or U1624 (N_1624,In_434,In_668);
nand U1625 (N_1625,In_481,In_562);
or U1626 (N_1626,In_590,In_224);
xor U1627 (N_1627,In_255,In_161);
nand U1628 (N_1628,In_332,In_278);
or U1629 (N_1629,In_307,In_564);
nand U1630 (N_1630,In_21,In_179);
and U1631 (N_1631,In_380,In_329);
or U1632 (N_1632,In_400,In_658);
nand U1633 (N_1633,In_389,In_99);
and U1634 (N_1634,In_244,In_486);
or U1635 (N_1635,In_273,In_583);
nor U1636 (N_1636,In_553,In_530);
nand U1637 (N_1637,In_328,In_568);
and U1638 (N_1638,In_699,In_419);
and U1639 (N_1639,In_335,In_440);
and U1640 (N_1640,In_670,In_26);
nand U1641 (N_1641,In_742,In_303);
or U1642 (N_1642,In_632,In_532);
nor U1643 (N_1643,In_390,In_291);
nor U1644 (N_1644,In_185,In_222);
nor U1645 (N_1645,In_457,In_619);
nor U1646 (N_1646,In_241,In_383);
and U1647 (N_1647,In_27,In_156);
nor U1648 (N_1648,In_693,In_454);
nor U1649 (N_1649,In_110,In_737);
or U1650 (N_1650,In_629,In_201);
or U1651 (N_1651,In_736,In_360);
nand U1652 (N_1652,In_493,In_52);
nor U1653 (N_1653,In_561,In_619);
or U1654 (N_1654,In_665,In_282);
or U1655 (N_1655,In_90,In_559);
or U1656 (N_1656,In_592,In_660);
and U1657 (N_1657,In_696,In_742);
and U1658 (N_1658,In_394,In_712);
and U1659 (N_1659,In_613,In_317);
nand U1660 (N_1660,In_9,In_24);
nor U1661 (N_1661,In_384,In_477);
or U1662 (N_1662,In_173,In_658);
nand U1663 (N_1663,In_516,In_350);
or U1664 (N_1664,In_311,In_406);
nand U1665 (N_1665,In_426,In_747);
nor U1666 (N_1666,In_703,In_694);
or U1667 (N_1667,In_424,In_41);
nor U1668 (N_1668,In_614,In_200);
nor U1669 (N_1669,In_739,In_304);
nor U1670 (N_1670,In_218,In_713);
or U1671 (N_1671,In_516,In_157);
or U1672 (N_1672,In_168,In_124);
nand U1673 (N_1673,In_256,In_422);
nor U1674 (N_1674,In_231,In_605);
or U1675 (N_1675,In_481,In_259);
xnor U1676 (N_1676,In_269,In_88);
and U1677 (N_1677,In_39,In_511);
or U1678 (N_1678,In_27,In_249);
and U1679 (N_1679,In_460,In_456);
and U1680 (N_1680,In_72,In_462);
nor U1681 (N_1681,In_345,In_256);
nor U1682 (N_1682,In_383,In_703);
nor U1683 (N_1683,In_694,In_379);
or U1684 (N_1684,In_331,In_177);
and U1685 (N_1685,In_712,In_684);
nor U1686 (N_1686,In_351,In_543);
nor U1687 (N_1687,In_212,In_713);
nand U1688 (N_1688,In_451,In_524);
or U1689 (N_1689,In_52,In_298);
or U1690 (N_1690,In_706,In_142);
nand U1691 (N_1691,In_180,In_581);
nand U1692 (N_1692,In_59,In_594);
nor U1693 (N_1693,In_454,In_700);
and U1694 (N_1694,In_100,In_354);
nor U1695 (N_1695,In_150,In_197);
nand U1696 (N_1696,In_497,In_295);
nand U1697 (N_1697,In_371,In_221);
and U1698 (N_1698,In_77,In_287);
and U1699 (N_1699,In_389,In_116);
or U1700 (N_1700,In_508,In_747);
and U1701 (N_1701,In_661,In_46);
and U1702 (N_1702,In_688,In_443);
nor U1703 (N_1703,In_401,In_29);
nor U1704 (N_1704,In_345,In_445);
nor U1705 (N_1705,In_644,In_582);
nor U1706 (N_1706,In_103,In_693);
and U1707 (N_1707,In_433,In_215);
nand U1708 (N_1708,In_161,In_463);
and U1709 (N_1709,In_714,In_319);
nand U1710 (N_1710,In_34,In_149);
and U1711 (N_1711,In_351,In_678);
or U1712 (N_1712,In_133,In_1);
or U1713 (N_1713,In_725,In_5);
or U1714 (N_1714,In_244,In_499);
and U1715 (N_1715,In_593,In_348);
and U1716 (N_1716,In_166,In_562);
or U1717 (N_1717,In_501,In_117);
and U1718 (N_1718,In_375,In_609);
or U1719 (N_1719,In_715,In_523);
nor U1720 (N_1720,In_31,In_595);
or U1721 (N_1721,In_729,In_391);
or U1722 (N_1722,In_481,In_113);
and U1723 (N_1723,In_66,In_166);
and U1724 (N_1724,In_65,In_357);
nand U1725 (N_1725,In_105,In_481);
nor U1726 (N_1726,In_512,In_156);
and U1727 (N_1727,In_482,In_297);
or U1728 (N_1728,In_615,In_352);
and U1729 (N_1729,In_275,In_90);
and U1730 (N_1730,In_336,In_34);
or U1731 (N_1731,In_25,In_138);
and U1732 (N_1732,In_181,In_376);
nor U1733 (N_1733,In_139,In_329);
and U1734 (N_1734,In_7,In_286);
nor U1735 (N_1735,In_296,In_647);
nor U1736 (N_1736,In_613,In_152);
nor U1737 (N_1737,In_236,In_137);
nor U1738 (N_1738,In_691,In_0);
or U1739 (N_1739,In_165,In_222);
nor U1740 (N_1740,In_356,In_385);
and U1741 (N_1741,In_730,In_184);
nor U1742 (N_1742,In_699,In_307);
nand U1743 (N_1743,In_335,In_24);
nor U1744 (N_1744,In_608,In_685);
nand U1745 (N_1745,In_683,In_450);
and U1746 (N_1746,In_519,In_596);
or U1747 (N_1747,In_154,In_247);
and U1748 (N_1748,In_585,In_430);
and U1749 (N_1749,In_642,In_496);
xnor U1750 (N_1750,In_47,In_176);
or U1751 (N_1751,In_80,In_309);
nand U1752 (N_1752,In_471,In_218);
and U1753 (N_1753,In_391,In_533);
nand U1754 (N_1754,In_675,In_690);
nand U1755 (N_1755,In_528,In_157);
nand U1756 (N_1756,In_29,In_522);
and U1757 (N_1757,In_13,In_565);
nand U1758 (N_1758,In_664,In_533);
and U1759 (N_1759,In_235,In_245);
nand U1760 (N_1760,In_233,In_314);
or U1761 (N_1761,In_505,In_308);
or U1762 (N_1762,In_11,In_33);
nand U1763 (N_1763,In_417,In_483);
nand U1764 (N_1764,In_244,In_229);
nor U1765 (N_1765,In_354,In_739);
and U1766 (N_1766,In_525,In_544);
nand U1767 (N_1767,In_261,In_676);
nand U1768 (N_1768,In_635,In_115);
nor U1769 (N_1769,In_623,In_689);
nand U1770 (N_1770,In_742,In_627);
nor U1771 (N_1771,In_62,In_119);
or U1772 (N_1772,In_383,In_505);
nand U1773 (N_1773,In_503,In_278);
nor U1774 (N_1774,In_453,In_429);
or U1775 (N_1775,In_343,In_57);
or U1776 (N_1776,In_48,In_536);
and U1777 (N_1777,In_430,In_102);
nand U1778 (N_1778,In_518,In_490);
or U1779 (N_1779,In_1,In_356);
or U1780 (N_1780,In_70,In_106);
nor U1781 (N_1781,In_333,In_538);
nand U1782 (N_1782,In_543,In_96);
and U1783 (N_1783,In_344,In_277);
and U1784 (N_1784,In_714,In_408);
and U1785 (N_1785,In_620,In_78);
nand U1786 (N_1786,In_65,In_742);
and U1787 (N_1787,In_388,In_360);
nand U1788 (N_1788,In_231,In_47);
nand U1789 (N_1789,In_659,In_259);
and U1790 (N_1790,In_661,In_106);
and U1791 (N_1791,In_393,In_489);
and U1792 (N_1792,In_100,In_303);
and U1793 (N_1793,In_264,In_128);
nor U1794 (N_1794,In_44,In_569);
nor U1795 (N_1795,In_530,In_148);
and U1796 (N_1796,In_460,In_318);
xnor U1797 (N_1797,In_535,In_380);
or U1798 (N_1798,In_301,In_432);
and U1799 (N_1799,In_749,In_357);
xor U1800 (N_1800,In_280,In_718);
nand U1801 (N_1801,In_145,In_469);
nor U1802 (N_1802,In_502,In_387);
nand U1803 (N_1803,In_274,In_425);
or U1804 (N_1804,In_38,In_160);
nand U1805 (N_1805,In_586,In_66);
or U1806 (N_1806,In_468,In_5);
or U1807 (N_1807,In_630,In_444);
nand U1808 (N_1808,In_647,In_250);
nand U1809 (N_1809,In_106,In_84);
and U1810 (N_1810,In_180,In_648);
nor U1811 (N_1811,In_117,In_396);
or U1812 (N_1812,In_15,In_658);
nor U1813 (N_1813,In_423,In_634);
nand U1814 (N_1814,In_330,In_265);
nand U1815 (N_1815,In_32,In_692);
nor U1816 (N_1816,In_654,In_472);
and U1817 (N_1817,In_620,In_735);
nand U1818 (N_1818,In_669,In_413);
nor U1819 (N_1819,In_685,In_433);
and U1820 (N_1820,In_526,In_542);
or U1821 (N_1821,In_555,In_604);
and U1822 (N_1822,In_674,In_165);
nand U1823 (N_1823,In_380,In_209);
and U1824 (N_1824,In_310,In_186);
or U1825 (N_1825,In_58,In_221);
nor U1826 (N_1826,In_169,In_206);
xnor U1827 (N_1827,In_26,In_665);
or U1828 (N_1828,In_278,In_78);
or U1829 (N_1829,In_555,In_644);
xnor U1830 (N_1830,In_82,In_481);
nor U1831 (N_1831,In_534,In_461);
nor U1832 (N_1832,In_665,In_729);
and U1833 (N_1833,In_346,In_14);
nor U1834 (N_1834,In_335,In_681);
or U1835 (N_1835,In_54,In_604);
or U1836 (N_1836,In_538,In_42);
nand U1837 (N_1837,In_377,In_716);
or U1838 (N_1838,In_277,In_204);
or U1839 (N_1839,In_248,In_388);
or U1840 (N_1840,In_157,In_683);
and U1841 (N_1841,In_159,In_280);
and U1842 (N_1842,In_589,In_602);
nor U1843 (N_1843,In_414,In_116);
and U1844 (N_1844,In_68,In_310);
nor U1845 (N_1845,In_636,In_525);
nand U1846 (N_1846,In_685,In_15);
and U1847 (N_1847,In_447,In_297);
nor U1848 (N_1848,In_46,In_625);
or U1849 (N_1849,In_129,In_735);
nor U1850 (N_1850,In_615,In_132);
and U1851 (N_1851,In_259,In_555);
and U1852 (N_1852,In_493,In_673);
or U1853 (N_1853,In_710,In_433);
nor U1854 (N_1854,In_242,In_387);
or U1855 (N_1855,In_501,In_622);
and U1856 (N_1856,In_227,In_323);
nand U1857 (N_1857,In_460,In_392);
nor U1858 (N_1858,In_224,In_306);
nor U1859 (N_1859,In_589,In_543);
xor U1860 (N_1860,In_95,In_312);
nor U1861 (N_1861,In_418,In_119);
nand U1862 (N_1862,In_260,In_740);
or U1863 (N_1863,In_479,In_649);
and U1864 (N_1864,In_288,In_401);
nand U1865 (N_1865,In_45,In_702);
nor U1866 (N_1866,In_202,In_208);
or U1867 (N_1867,In_550,In_399);
and U1868 (N_1868,In_225,In_101);
or U1869 (N_1869,In_45,In_247);
nand U1870 (N_1870,In_206,In_733);
or U1871 (N_1871,In_541,In_194);
nand U1872 (N_1872,In_247,In_493);
nand U1873 (N_1873,In_332,In_571);
or U1874 (N_1874,In_105,In_711);
or U1875 (N_1875,In_370,In_487);
and U1876 (N_1876,In_438,In_481);
or U1877 (N_1877,In_16,In_575);
or U1878 (N_1878,In_263,In_586);
or U1879 (N_1879,In_59,In_21);
or U1880 (N_1880,In_10,In_7);
nand U1881 (N_1881,In_192,In_88);
or U1882 (N_1882,In_356,In_698);
nor U1883 (N_1883,In_54,In_498);
nor U1884 (N_1884,In_274,In_308);
and U1885 (N_1885,In_121,In_135);
or U1886 (N_1886,In_168,In_147);
or U1887 (N_1887,In_253,In_102);
xnor U1888 (N_1888,In_609,In_590);
nand U1889 (N_1889,In_323,In_294);
or U1890 (N_1890,In_650,In_511);
nand U1891 (N_1891,In_687,In_525);
nand U1892 (N_1892,In_235,In_675);
or U1893 (N_1893,In_355,In_722);
and U1894 (N_1894,In_608,In_141);
and U1895 (N_1895,In_241,In_604);
nor U1896 (N_1896,In_277,In_415);
xnor U1897 (N_1897,In_289,In_336);
nor U1898 (N_1898,In_84,In_659);
nand U1899 (N_1899,In_658,In_652);
nand U1900 (N_1900,In_495,In_552);
or U1901 (N_1901,In_423,In_26);
or U1902 (N_1902,In_20,In_2);
or U1903 (N_1903,In_250,In_453);
nor U1904 (N_1904,In_398,In_155);
or U1905 (N_1905,In_146,In_163);
nor U1906 (N_1906,In_302,In_101);
nor U1907 (N_1907,In_595,In_186);
or U1908 (N_1908,In_249,In_221);
and U1909 (N_1909,In_138,In_580);
nand U1910 (N_1910,In_538,In_352);
nand U1911 (N_1911,In_141,In_732);
nor U1912 (N_1912,In_258,In_401);
nand U1913 (N_1913,In_402,In_603);
or U1914 (N_1914,In_69,In_262);
and U1915 (N_1915,In_739,In_301);
and U1916 (N_1916,In_727,In_682);
xnor U1917 (N_1917,In_69,In_76);
and U1918 (N_1918,In_114,In_75);
nand U1919 (N_1919,In_135,In_196);
and U1920 (N_1920,In_178,In_115);
nor U1921 (N_1921,In_235,In_89);
and U1922 (N_1922,In_424,In_85);
nor U1923 (N_1923,In_289,In_566);
and U1924 (N_1924,In_527,In_386);
xnor U1925 (N_1925,In_303,In_14);
and U1926 (N_1926,In_245,In_322);
and U1927 (N_1927,In_608,In_339);
and U1928 (N_1928,In_207,In_264);
or U1929 (N_1929,In_528,In_592);
or U1930 (N_1930,In_457,In_696);
or U1931 (N_1931,In_76,In_570);
nor U1932 (N_1932,In_353,In_214);
and U1933 (N_1933,In_428,In_351);
nand U1934 (N_1934,In_300,In_496);
and U1935 (N_1935,In_102,In_662);
and U1936 (N_1936,In_31,In_404);
nand U1937 (N_1937,In_369,In_463);
and U1938 (N_1938,In_9,In_70);
and U1939 (N_1939,In_651,In_118);
nor U1940 (N_1940,In_512,In_589);
nor U1941 (N_1941,In_473,In_247);
nand U1942 (N_1942,In_55,In_291);
or U1943 (N_1943,In_279,In_216);
or U1944 (N_1944,In_243,In_590);
or U1945 (N_1945,In_574,In_435);
nand U1946 (N_1946,In_640,In_636);
or U1947 (N_1947,In_628,In_720);
nor U1948 (N_1948,In_456,In_415);
and U1949 (N_1949,In_42,In_687);
nand U1950 (N_1950,In_50,In_82);
nor U1951 (N_1951,In_334,In_289);
and U1952 (N_1952,In_522,In_482);
or U1953 (N_1953,In_453,In_580);
and U1954 (N_1954,In_699,In_297);
xor U1955 (N_1955,In_748,In_665);
or U1956 (N_1956,In_346,In_473);
and U1957 (N_1957,In_11,In_378);
nand U1958 (N_1958,In_435,In_296);
or U1959 (N_1959,In_189,In_447);
nor U1960 (N_1960,In_310,In_77);
and U1961 (N_1961,In_287,In_510);
nor U1962 (N_1962,In_642,In_201);
or U1963 (N_1963,In_493,In_703);
nand U1964 (N_1964,In_276,In_500);
or U1965 (N_1965,In_76,In_335);
nor U1966 (N_1966,In_244,In_301);
or U1967 (N_1967,In_121,In_2);
nand U1968 (N_1968,In_646,In_395);
and U1969 (N_1969,In_610,In_668);
nor U1970 (N_1970,In_510,In_473);
and U1971 (N_1971,In_576,In_548);
and U1972 (N_1972,In_678,In_697);
and U1973 (N_1973,In_516,In_174);
nand U1974 (N_1974,In_298,In_21);
or U1975 (N_1975,In_347,In_246);
nand U1976 (N_1976,In_496,In_519);
and U1977 (N_1977,In_406,In_619);
and U1978 (N_1978,In_187,In_711);
and U1979 (N_1979,In_461,In_154);
nor U1980 (N_1980,In_8,In_109);
nand U1981 (N_1981,In_68,In_201);
or U1982 (N_1982,In_381,In_292);
nand U1983 (N_1983,In_339,In_580);
nor U1984 (N_1984,In_414,In_331);
nand U1985 (N_1985,In_416,In_104);
nand U1986 (N_1986,In_389,In_354);
and U1987 (N_1987,In_492,In_594);
nor U1988 (N_1988,In_361,In_520);
nor U1989 (N_1989,In_206,In_600);
xnor U1990 (N_1990,In_449,In_429);
xnor U1991 (N_1991,In_398,In_749);
nor U1992 (N_1992,In_447,In_669);
nand U1993 (N_1993,In_608,In_110);
and U1994 (N_1994,In_111,In_395);
and U1995 (N_1995,In_85,In_413);
or U1996 (N_1996,In_709,In_403);
nor U1997 (N_1997,In_559,In_16);
or U1998 (N_1998,In_156,In_606);
or U1999 (N_1999,In_39,In_441);
nor U2000 (N_2000,In_588,In_470);
xor U2001 (N_2001,In_55,In_684);
nand U2002 (N_2002,In_16,In_270);
or U2003 (N_2003,In_616,In_672);
or U2004 (N_2004,In_140,In_384);
or U2005 (N_2005,In_714,In_197);
and U2006 (N_2006,In_316,In_48);
nor U2007 (N_2007,In_509,In_716);
and U2008 (N_2008,In_157,In_297);
and U2009 (N_2009,In_40,In_466);
and U2010 (N_2010,In_34,In_238);
and U2011 (N_2011,In_252,In_326);
nor U2012 (N_2012,In_426,In_231);
and U2013 (N_2013,In_65,In_480);
nor U2014 (N_2014,In_228,In_131);
nor U2015 (N_2015,In_400,In_516);
or U2016 (N_2016,In_556,In_161);
nor U2017 (N_2017,In_651,In_479);
nor U2018 (N_2018,In_540,In_280);
or U2019 (N_2019,In_583,In_148);
nor U2020 (N_2020,In_481,In_448);
xor U2021 (N_2021,In_105,In_69);
or U2022 (N_2022,In_410,In_574);
nor U2023 (N_2023,In_424,In_667);
nor U2024 (N_2024,In_171,In_439);
nor U2025 (N_2025,In_559,In_146);
or U2026 (N_2026,In_509,In_205);
and U2027 (N_2027,In_120,In_691);
nand U2028 (N_2028,In_404,In_379);
or U2029 (N_2029,In_111,In_484);
nand U2030 (N_2030,In_194,In_513);
and U2031 (N_2031,In_440,In_731);
nand U2032 (N_2032,In_440,In_734);
nand U2033 (N_2033,In_187,In_93);
nand U2034 (N_2034,In_563,In_654);
xnor U2035 (N_2035,In_246,In_147);
nand U2036 (N_2036,In_14,In_435);
nand U2037 (N_2037,In_143,In_50);
nor U2038 (N_2038,In_91,In_408);
nand U2039 (N_2039,In_15,In_105);
and U2040 (N_2040,In_619,In_100);
nand U2041 (N_2041,In_112,In_85);
or U2042 (N_2042,In_224,In_460);
nand U2043 (N_2043,In_336,In_123);
and U2044 (N_2044,In_75,In_354);
nor U2045 (N_2045,In_644,In_4);
or U2046 (N_2046,In_486,In_165);
nand U2047 (N_2047,In_59,In_331);
or U2048 (N_2048,In_587,In_524);
or U2049 (N_2049,In_293,In_481);
xor U2050 (N_2050,In_624,In_97);
or U2051 (N_2051,In_90,In_379);
nand U2052 (N_2052,In_128,In_260);
nand U2053 (N_2053,In_620,In_165);
or U2054 (N_2054,In_492,In_340);
nor U2055 (N_2055,In_700,In_289);
and U2056 (N_2056,In_164,In_388);
nor U2057 (N_2057,In_462,In_54);
and U2058 (N_2058,In_496,In_411);
and U2059 (N_2059,In_440,In_344);
or U2060 (N_2060,In_465,In_654);
or U2061 (N_2061,In_319,In_102);
and U2062 (N_2062,In_632,In_98);
nand U2063 (N_2063,In_584,In_599);
or U2064 (N_2064,In_71,In_379);
nand U2065 (N_2065,In_239,In_726);
or U2066 (N_2066,In_410,In_686);
nor U2067 (N_2067,In_609,In_87);
nor U2068 (N_2068,In_92,In_213);
or U2069 (N_2069,In_154,In_329);
or U2070 (N_2070,In_61,In_131);
nor U2071 (N_2071,In_576,In_633);
nand U2072 (N_2072,In_189,In_2);
or U2073 (N_2073,In_241,In_481);
nand U2074 (N_2074,In_485,In_104);
nor U2075 (N_2075,In_725,In_85);
nand U2076 (N_2076,In_118,In_695);
nor U2077 (N_2077,In_135,In_357);
and U2078 (N_2078,In_597,In_740);
and U2079 (N_2079,In_288,In_732);
and U2080 (N_2080,In_513,In_140);
or U2081 (N_2081,In_529,In_118);
nand U2082 (N_2082,In_84,In_416);
or U2083 (N_2083,In_85,In_170);
and U2084 (N_2084,In_72,In_322);
xor U2085 (N_2085,In_215,In_252);
nand U2086 (N_2086,In_250,In_327);
nor U2087 (N_2087,In_485,In_197);
nor U2088 (N_2088,In_590,In_167);
or U2089 (N_2089,In_174,In_545);
or U2090 (N_2090,In_221,In_79);
or U2091 (N_2091,In_107,In_118);
and U2092 (N_2092,In_331,In_436);
or U2093 (N_2093,In_460,In_554);
nand U2094 (N_2094,In_588,In_39);
nor U2095 (N_2095,In_361,In_499);
nor U2096 (N_2096,In_258,In_606);
nand U2097 (N_2097,In_680,In_248);
nor U2098 (N_2098,In_573,In_332);
or U2099 (N_2099,In_665,In_20);
nor U2100 (N_2100,In_612,In_310);
nand U2101 (N_2101,In_147,In_417);
or U2102 (N_2102,In_266,In_310);
and U2103 (N_2103,In_698,In_37);
or U2104 (N_2104,In_175,In_264);
nand U2105 (N_2105,In_268,In_390);
and U2106 (N_2106,In_630,In_56);
or U2107 (N_2107,In_729,In_55);
nand U2108 (N_2108,In_227,In_659);
nor U2109 (N_2109,In_161,In_535);
or U2110 (N_2110,In_723,In_588);
or U2111 (N_2111,In_233,In_639);
nand U2112 (N_2112,In_641,In_3);
nor U2113 (N_2113,In_96,In_619);
or U2114 (N_2114,In_288,In_153);
nand U2115 (N_2115,In_499,In_130);
nor U2116 (N_2116,In_604,In_75);
nor U2117 (N_2117,In_650,In_682);
or U2118 (N_2118,In_594,In_427);
or U2119 (N_2119,In_467,In_335);
xor U2120 (N_2120,In_728,In_710);
nand U2121 (N_2121,In_114,In_634);
nor U2122 (N_2122,In_140,In_116);
and U2123 (N_2123,In_534,In_293);
and U2124 (N_2124,In_23,In_604);
or U2125 (N_2125,In_228,In_124);
nor U2126 (N_2126,In_414,In_220);
and U2127 (N_2127,In_487,In_478);
nand U2128 (N_2128,In_350,In_173);
nor U2129 (N_2129,In_708,In_164);
and U2130 (N_2130,In_274,In_412);
nor U2131 (N_2131,In_103,In_302);
nor U2132 (N_2132,In_188,In_654);
or U2133 (N_2133,In_13,In_330);
xnor U2134 (N_2134,In_27,In_427);
or U2135 (N_2135,In_248,In_28);
xnor U2136 (N_2136,In_241,In_685);
nand U2137 (N_2137,In_193,In_642);
and U2138 (N_2138,In_646,In_50);
nor U2139 (N_2139,In_184,In_128);
nand U2140 (N_2140,In_94,In_168);
or U2141 (N_2141,In_301,In_36);
or U2142 (N_2142,In_39,In_82);
or U2143 (N_2143,In_280,In_256);
nor U2144 (N_2144,In_539,In_83);
or U2145 (N_2145,In_29,In_67);
nor U2146 (N_2146,In_455,In_538);
or U2147 (N_2147,In_625,In_598);
and U2148 (N_2148,In_625,In_33);
nand U2149 (N_2149,In_514,In_665);
nor U2150 (N_2150,In_649,In_569);
and U2151 (N_2151,In_268,In_141);
nor U2152 (N_2152,In_227,In_133);
nand U2153 (N_2153,In_669,In_552);
and U2154 (N_2154,In_641,In_69);
nor U2155 (N_2155,In_321,In_125);
or U2156 (N_2156,In_336,In_163);
nor U2157 (N_2157,In_6,In_122);
nor U2158 (N_2158,In_302,In_690);
nand U2159 (N_2159,In_244,In_235);
or U2160 (N_2160,In_562,In_612);
nor U2161 (N_2161,In_489,In_641);
nor U2162 (N_2162,In_89,In_168);
and U2163 (N_2163,In_177,In_457);
nand U2164 (N_2164,In_198,In_435);
and U2165 (N_2165,In_415,In_351);
nand U2166 (N_2166,In_621,In_372);
nor U2167 (N_2167,In_163,In_107);
or U2168 (N_2168,In_568,In_635);
nor U2169 (N_2169,In_43,In_376);
and U2170 (N_2170,In_211,In_554);
or U2171 (N_2171,In_101,In_625);
xor U2172 (N_2172,In_648,In_407);
or U2173 (N_2173,In_357,In_270);
and U2174 (N_2174,In_77,In_645);
nor U2175 (N_2175,In_479,In_520);
nand U2176 (N_2176,In_527,In_553);
nor U2177 (N_2177,In_31,In_6);
and U2178 (N_2178,In_554,In_209);
and U2179 (N_2179,In_628,In_450);
nor U2180 (N_2180,In_23,In_525);
or U2181 (N_2181,In_315,In_394);
and U2182 (N_2182,In_705,In_306);
nor U2183 (N_2183,In_325,In_9);
nor U2184 (N_2184,In_450,In_246);
and U2185 (N_2185,In_231,In_572);
nand U2186 (N_2186,In_503,In_21);
and U2187 (N_2187,In_650,In_167);
or U2188 (N_2188,In_390,In_703);
nand U2189 (N_2189,In_611,In_151);
nor U2190 (N_2190,In_155,In_412);
nand U2191 (N_2191,In_232,In_371);
or U2192 (N_2192,In_490,In_115);
nand U2193 (N_2193,In_643,In_167);
nor U2194 (N_2194,In_456,In_504);
or U2195 (N_2195,In_375,In_694);
or U2196 (N_2196,In_360,In_511);
nor U2197 (N_2197,In_714,In_547);
nor U2198 (N_2198,In_334,In_139);
nor U2199 (N_2199,In_320,In_567);
nand U2200 (N_2200,In_222,In_340);
or U2201 (N_2201,In_604,In_92);
nand U2202 (N_2202,In_96,In_297);
or U2203 (N_2203,In_619,In_338);
or U2204 (N_2204,In_344,In_645);
or U2205 (N_2205,In_7,In_215);
nor U2206 (N_2206,In_475,In_612);
and U2207 (N_2207,In_741,In_434);
and U2208 (N_2208,In_481,In_157);
nand U2209 (N_2209,In_68,In_69);
and U2210 (N_2210,In_189,In_428);
or U2211 (N_2211,In_744,In_722);
or U2212 (N_2212,In_201,In_631);
nand U2213 (N_2213,In_213,In_73);
nand U2214 (N_2214,In_561,In_587);
nor U2215 (N_2215,In_11,In_365);
nand U2216 (N_2216,In_61,In_702);
nand U2217 (N_2217,In_116,In_654);
or U2218 (N_2218,In_306,In_441);
nand U2219 (N_2219,In_700,In_460);
xnor U2220 (N_2220,In_390,In_582);
or U2221 (N_2221,In_426,In_466);
or U2222 (N_2222,In_284,In_191);
or U2223 (N_2223,In_308,In_363);
nor U2224 (N_2224,In_275,In_151);
nor U2225 (N_2225,In_166,In_491);
or U2226 (N_2226,In_697,In_15);
and U2227 (N_2227,In_628,In_301);
nor U2228 (N_2228,In_531,In_288);
nand U2229 (N_2229,In_494,In_230);
and U2230 (N_2230,In_240,In_674);
and U2231 (N_2231,In_254,In_630);
nand U2232 (N_2232,In_362,In_99);
and U2233 (N_2233,In_135,In_500);
nand U2234 (N_2234,In_339,In_598);
nand U2235 (N_2235,In_107,In_513);
and U2236 (N_2236,In_506,In_570);
nand U2237 (N_2237,In_716,In_418);
and U2238 (N_2238,In_133,In_45);
nor U2239 (N_2239,In_6,In_264);
or U2240 (N_2240,In_568,In_512);
xor U2241 (N_2241,In_123,In_96);
or U2242 (N_2242,In_154,In_85);
nand U2243 (N_2243,In_14,In_439);
nand U2244 (N_2244,In_292,In_244);
nand U2245 (N_2245,In_679,In_357);
nor U2246 (N_2246,In_33,In_66);
nor U2247 (N_2247,In_592,In_616);
nor U2248 (N_2248,In_70,In_151);
and U2249 (N_2249,In_408,In_624);
and U2250 (N_2250,In_78,In_442);
xor U2251 (N_2251,In_637,In_56);
nand U2252 (N_2252,In_352,In_505);
nand U2253 (N_2253,In_220,In_656);
and U2254 (N_2254,In_94,In_697);
nor U2255 (N_2255,In_447,In_298);
nand U2256 (N_2256,In_386,In_330);
and U2257 (N_2257,In_86,In_640);
nand U2258 (N_2258,In_557,In_250);
nand U2259 (N_2259,In_386,In_361);
nor U2260 (N_2260,In_424,In_583);
and U2261 (N_2261,In_460,In_613);
nand U2262 (N_2262,In_694,In_689);
nor U2263 (N_2263,In_44,In_319);
nand U2264 (N_2264,In_657,In_1);
or U2265 (N_2265,In_651,In_538);
or U2266 (N_2266,In_501,In_624);
nor U2267 (N_2267,In_483,In_653);
nand U2268 (N_2268,In_505,In_489);
or U2269 (N_2269,In_73,In_117);
or U2270 (N_2270,In_17,In_472);
nand U2271 (N_2271,In_483,In_188);
nand U2272 (N_2272,In_348,In_566);
nor U2273 (N_2273,In_523,In_557);
or U2274 (N_2274,In_210,In_79);
or U2275 (N_2275,In_142,In_52);
nand U2276 (N_2276,In_298,In_717);
and U2277 (N_2277,In_410,In_75);
and U2278 (N_2278,In_739,In_327);
or U2279 (N_2279,In_414,In_227);
or U2280 (N_2280,In_637,In_510);
nor U2281 (N_2281,In_695,In_372);
or U2282 (N_2282,In_20,In_226);
xnor U2283 (N_2283,In_29,In_333);
and U2284 (N_2284,In_89,In_119);
nor U2285 (N_2285,In_710,In_252);
nand U2286 (N_2286,In_499,In_362);
and U2287 (N_2287,In_315,In_549);
and U2288 (N_2288,In_381,In_576);
nor U2289 (N_2289,In_44,In_222);
or U2290 (N_2290,In_659,In_97);
nand U2291 (N_2291,In_314,In_594);
nor U2292 (N_2292,In_165,In_199);
nand U2293 (N_2293,In_53,In_304);
and U2294 (N_2294,In_556,In_98);
nand U2295 (N_2295,In_254,In_21);
nand U2296 (N_2296,In_649,In_154);
nor U2297 (N_2297,In_726,In_613);
and U2298 (N_2298,In_701,In_282);
and U2299 (N_2299,In_517,In_238);
and U2300 (N_2300,In_190,In_381);
nand U2301 (N_2301,In_568,In_159);
nor U2302 (N_2302,In_28,In_662);
or U2303 (N_2303,In_373,In_443);
and U2304 (N_2304,In_207,In_582);
nor U2305 (N_2305,In_432,In_296);
nor U2306 (N_2306,In_98,In_243);
nor U2307 (N_2307,In_187,In_613);
and U2308 (N_2308,In_594,In_571);
xnor U2309 (N_2309,In_127,In_745);
nand U2310 (N_2310,In_83,In_209);
nor U2311 (N_2311,In_457,In_149);
nor U2312 (N_2312,In_318,In_302);
and U2313 (N_2313,In_620,In_42);
and U2314 (N_2314,In_426,In_93);
nor U2315 (N_2315,In_395,In_187);
or U2316 (N_2316,In_642,In_191);
or U2317 (N_2317,In_502,In_451);
and U2318 (N_2318,In_492,In_313);
nor U2319 (N_2319,In_341,In_189);
and U2320 (N_2320,In_371,In_281);
nor U2321 (N_2321,In_709,In_545);
nor U2322 (N_2322,In_400,In_286);
and U2323 (N_2323,In_459,In_528);
nand U2324 (N_2324,In_278,In_383);
or U2325 (N_2325,In_449,In_668);
xnor U2326 (N_2326,In_406,In_49);
nor U2327 (N_2327,In_503,In_496);
nor U2328 (N_2328,In_747,In_595);
and U2329 (N_2329,In_243,In_293);
nor U2330 (N_2330,In_643,In_721);
nor U2331 (N_2331,In_289,In_449);
or U2332 (N_2332,In_70,In_575);
and U2333 (N_2333,In_12,In_475);
or U2334 (N_2334,In_286,In_409);
nand U2335 (N_2335,In_235,In_699);
nor U2336 (N_2336,In_529,In_438);
or U2337 (N_2337,In_382,In_659);
or U2338 (N_2338,In_34,In_109);
nand U2339 (N_2339,In_39,In_717);
or U2340 (N_2340,In_132,In_515);
or U2341 (N_2341,In_624,In_536);
or U2342 (N_2342,In_34,In_575);
xnor U2343 (N_2343,In_239,In_646);
nand U2344 (N_2344,In_25,In_182);
and U2345 (N_2345,In_391,In_164);
xnor U2346 (N_2346,In_119,In_678);
and U2347 (N_2347,In_580,In_748);
nor U2348 (N_2348,In_716,In_463);
or U2349 (N_2349,In_351,In_26);
and U2350 (N_2350,In_389,In_159);
nor U2351 (N_2351,In_229,In_587);
and U2352 (N_2352,In_638,In_21);
nor U2353 (N_2353,In_71,In_34);
nand U2354 (N_2354,In_354,In_370);
nor U2355 (N_2355,In_749,In_81);
or U2356 (N_2356,In_627,In_254);
nor U2357 (N_2357,In_237,In_345);
or U2358 (N_2358,In_455,In_637);
or U2359 (N_2359,In_70,In_563);
and U2360 (N_2360,In_189,In_694);
and U2361 (N_2361,In_607,In_416);
nor U2362 (N_2362,In_155,In_690);
nand U2363 (N_2363,In_657,In_221);
nand U2364 (N_2364,In_558,In_171);
nand U2365 (N_2365,In_490,In_510);
or U2366 (N_2366,In_451,In_110);
and U2367 (N_2367,In_247,In_207);
or U2368 (N_2368,In_358,In_591);
and U2369 (N_2369,In_325,In_635);
or U2370 (N_2370,In_749,In_735);
and U2371 (N_2371,In_517,In_506);
nand U2372 (N_2372,In_270,In_306);
nor U2373 (N_2373,In_354,In_203);
or U2374 (N_2374,In_501,In_611);
nor U2375 (N_2375,In_633,In_537);
nor U2376 (N_2376,In_169,In_245);
nor U2377 (N_2377,In_158,In_601);
nor U2378 (N_2378,In_532,In_233);
or U2379 (N_2379,In_601,In_584);
nor U2380 (N_2380,In_48,In_595);
nor U2381 (N_2381,In_725,In_303);
nor U2382 (N_2382,In_145,In_191);
xor U2383 (N_2383,In_719,In_710);
or U2384 (N_2384,In_536,In_49);
nor U2385 (N_2385,In_581,In_677);
nand U2386 (N_2386,In_497,In_12);
or U2387 (N_2387,In_206,In_37);
nor U2388 (N_2388,In_0,In_169);
nand U2389 (N_2389,In_463,In_178);
or U2390 (N_2390,In_343,In_726);
nand U2391 (N_2391,In_67,In_293);
nor U2392 (N_2392,In_489,In_130);
and U2393 (N_2393,In_727,In_224);
and U2394 (N_2394,In_148,In_378);
nand U2395 (N_2395,In_371,In_257);
and U2396 (N_2396,In_207,In_134);
nand U2397 (N_2397,In_564,In_106);
xor U2398 (N_2398,In_516,In_296);
and U2399 (N_2399,In_547,In_414);
or U2400 (N_2400,In_600,In_561);
and U2401 (N_2401,In_34,In_282);
and U2402 (N_2402,In_350,In_600);
nor U2403 (N_2403,In_355,In_383);
or U2404 (N_2404,In_37,In_380);
nand U2405 (N_2405,In_642,In_392);
nor U2406 (N_2406,In_230,In_222);
nor U2407 (N_2407,In_211,In_498);
or U2408 (N_2408,In_651,In_4);
or U2409 (N_2409,In_286,In_475);
nor U2410 (N_2410,In_129,In_235);
and U2411 (N_2411,In_571,In_664);
nand U2412 (N_2412,In_63,In_107);
xnor U2413 (N_2413,In_180,In_299);
nor U2414 (N_2414,In_148,In_129);
xnor U2415 (N_2415,In_209,In_222);
xor U2416 (N_2416,In_256,In_38);
nand U2417 (N_2417,In_542,In_598);
nor U2418 (N_2418,In_519,In_732);
nand U2419 (N_2419,In_637,In_461);
nand U2420 (N_2420,In_501,In_548);
and U2421 (N_2421,In_448,In_207);
nor U2422 (N_2422,In_183,In_18);
nor U2423 (N_2423,In_159,In_449);
and U2424 (N_2424,In_724,In_392);
or U2425 (N_2425,In_309,In_335);
nand U2426 (N_2426,In_691,In_72);
nor U2427 (N_2427,In_603,In_711);
or U2428 (N_2428,In_291,In_122);
nor U2429 (N_2429,In_500,In_567);
nand U2430 (N_2430,In_533,In_585);
and U2431 (N_2431,In_194,In_407);
and U2432 (N_2432,In_394,In_224);
nor U2433 (N_2433,In_71,In_631);
nand U2434 (N_2434,In_566,In_361);
or U2435 (N_2435,In_195,In_65);
xnor U2436 (N_2436,In_53,In_281);
nor U2437 (N_2437,In_8,In_416);
nor U2438 (N_2438,In_642,In_383);
nor U2439 (N_2439,In_365,In_71);
and U2440 (N_2440,In_522,In_471);
and U2441 (N_2441,In_210,In_484);
nor U2442 (N_2442,In_80,In_209);
nor U2443 (N_2443,In_495,In_685);
or U2444 (N_2444,In_331,In_744);
nor U2445 (N_2445,In_316,In_452);
nand U2446 (N_2446,In_225,In_484);
or U2447 (N_2447,In_104,In_478);
nor U2448 (N_2448,In_29,In_165);
or U2449 (N_2449,In_603,In_208);
nand U2450 (N_2450,In_7,In_494);
and U2451 (N_2451,In_213,In_85);
nand U2452 (N_2452,In_140,In_150);
nor U2453 (N_2453,In_151,In_451);
nor U2454 (N_2454,In_372,In_633);
nand U2455 (N_2455,In_374,In_277);
nor U2456 (N_2456,In_581,In_78);
and U2457 (N_2457,In_490,In_434);
and U2458 (N_2458,In_645,In_298);
or U2459 (N_2459,In_37,In_116);
nand U2460 (N_2460,In_441,In_354);
or U2461 (N_2461,In_517,In_654);
xor U2462 (N_2462,In_497,In_747);
nor U2463 (N_2463,In_739,In_275);
or U2464 (N_2464,In_155,In_442);
nor U2465 (N_2465,In_295,In_528);
nand U2466 (N_2466,In_222,In_370);
nand U2467 (N_2467,In_731,In_589);
or U2468 (N_2468,In_624,In_85);
nor U2469 (N_2469,In_443,In_206);
nand U2470 (N_2470,In_493,In_747);
nor U2471 (N_2471,In_261,In_190);
and U2472 (N_2472,In_616,In_561);
and U2473 (N_2473,In_75,In_540);
nor U2474 (N_2474,In_55,In_209);
nor U2475 (N_2475,In_527,In_251);
nor U2476 (N_2476,In_4,In_708);
and U2477 (N_2477,In_655,In_87);
nor U2478 (N_2478,In_67,In_17);
nand U2479 (N_2479,In_522,In_63);
nor U2480 (N_2480,In_581,In_56);
or U2481 (N_2481,In_129,In_725);
or U2482 (N_2482,In_571,In_267);
or U2483 (N_2483,In_277,In_433);
and U2484 (N_2484,In_256,In_584);
nand U2485 (N_2485,In_158,In_740);
nor U2486 (N_2486,In_665,In_171);
or U2487 (N_2487,In_466,In_334);
nand U2488 (N_2488,In_566,In_113);
nor U2489 (N_2489,In_202,In_69);
nand U2490 (N_2490,In_549,In_553);
or U2491 (N_2491,In_152,In_212);
and U2492 (N_2492,In_445,In_302);
and U2493 (N_2493,In_18,In_23);
xnor U2494 (N_2494,In_636,In_586);
and U2495 (N_2495,In_686,In_414);
nor U2496 (N_2496,In_522,In_730);
nand U2497 (N_2497,In_210,In_312);
and U2498 (N_2498,In_49,In_428);
nand U2499 (N_2499,In_10,In_519);
or U2500 (N_2500,N_2498,N_131);
nand U2501 (N_2501,N_1525,N_340);
and U2502 (N_2502,N_1123,N_1826);
or U2503 (N_2503,N_1768,N_1865);
and U2504 (N_2504,N_1122,N_2428);
and U2505 (N_2505,N_1916,N_703);
nand U2506 (N_2506,N_1535,N_2257);
xor U2507 (N_2507,N_719,N_934);
nor U2508 (N_2508,N_269,N_11);
or U2509 (N_2509,N_621,N_90);
and U2510 (N_2510,N_1915,N_1978);
nor U2511 (N_2511,N_149,N_1508);
and U2512 (N_2512,N_1064,N_1977);
nor U2513 (N_2513,N_1721,N_1901);
or U2514 (N_2514,N_605,N_1043);
nand U2515 (N_2515,N_751,N_1181);
or U2516 (N_2516,N_157,N_1139);
and U2517 (N_2517,N_287,N_1247);
and U2518 (N_2518,N_4,N_481);
and U2519 (N_2519,N_811,N_1646);
or U2520 (N_2520,N_1930,N_1843);
nand U2521 (N_2521,N_2239,N_188);
and U2522 (N_2522,N_2312,N_1223);
and U2523 (N_2523,N_898,N_416);
nor U2524 (N_2524,N_1769,N_48);
nor U2525 (N_2525,N_1377,N_2468);
nand U2526 (N_2526,N_557,N_1649);
and U2527 (N_2527,N_1522,N_1288);
nand U2528 (N_2528,N_2180,N_1953);
or U2529 (N_2529,N_1531,N_1393);
or U2530 (N_2530,N_1324,N_1200);
nand U2531 (N_2531,N_492,N_683);
and U2532 (N_2532,N_1986,N_1255);
nor U2533 (N_2533,N_874,N_943);
nor U2534 (N_2534,N_349,N_2270);
and U2535 (N_2535,N_9,N_2456);
or U2536 (N_2536,N_235,N_1638);
nand U2537 (N_2537,N_2075,N_45);
and U2538 (N_2538,N_101,N_1215);
or U2539 (N_2539,N_54,N_2238);
nand U2540 (N_2540,N_896,N_1461);
nand U2541 (N_2541,N_726,N_2076);
and U2542 (N_2542,N_1902,N_1048);
nand U2543 (N_2543,N_440,N_1842);
and U2544 (N_2544,N_749,N_316);
nand U2545 (N_2545,N_200,N_845);
nand U2546 (N_2546,N_1702,N_1925);
nand U2547 (N_2547,N_789,N_1246);
nor U2548 (N_2548,N_232,N_1654);
or U2549 (N_2549,N_488,N_2092);
and U2550 (N_2550,N_1631,N_572);
nand U2551 (N_2551,N_530,N_2337);
and U2552 (N_2552,N_836,N_800);
and U2553 (N_2553,N_341,N_376);
nand U2554 (N_2554,N_6,N_2386);
nor U2555 (N_2555,N_1455,N_2083);
nand U2556 (N_2556,N_1801,N_458);
or U2557 (N_2557,N_599,N_1680);
nand U2558 (N_2558,N_46,N_2318);
or U2559 (N_2559,N_1292,N_1671);
or U2560 (N_2560,N_2380,N_705);
xor U2561 (N_2561,N_987,N_296);
nor U2562 (N_2562,N_190,N_1162);
nand U2563 (N_2563,N_533,N_1530);
or U2564 (N_2564,N_1211,N_788);
nand U2565 (N_2565,N_402,N_1808);
and U2566 (N_2566,N_1078,N_975);
or U2567 (N_2567,N_741,N_1841);
nor U2568 (N_2568,N_2465,N_1598);
nor U2569 (N_2569,N_1354,N_1956);
nor U2570 (N_2570,N_833,N_2302);
or U2571 (N_2571,N_1759,N_2101);
nand U2572 (N_2572,N_2137,N_1148);
or U2573 (N_2573,N_1551,N_2426);
or U2574 (N_2574,N_1846,N_2474);
and U2575 (N_2575,N_191,N_1490);
nand U2576 (N_2576,N_756,N_2469);
or U2577 (N_2577,N_1595,N_920);
and U2578 (N_2578,N_1844,N_202);
and U2579 (N_2579,N_2209,N_445);
nand U2580 (N_2580,N_728,N_2371);
or U2581 (N_2581,N_1960,N_291);
and U2582 (N_2582,N_392,N_1491);
and U2583 (N_2583,N_328,N_1295);
and U2584 (N_2584,N_2353,N_1198);
or U2585 (N_2585,N_2344,N_733);
nand U2586 (N_2586,N_56,N_1378);
xnor U2587 (N_2587,N_2268,N_245);
nand U2588 (N_2588,N_638,N_565);
nand U2589 (N_2589,N_1875,N_700);
or U2590 (N_2590,N_2422,N_140);
nor U2591 (N_2591,N_2043,N_978);
and U2592 (N_2592,N_531,N_1413);
xor U2593 (N_2593,N_2154,N_2414);
or U2594 (N_2594,N_448,N_2390);
and U2595 (N_2595,N_817,N_2105);
xor U2596 (N_2596,N_1163,N_1066);
and U2597 (N_2597,N_867,N_2225);
nor U2598 (N_2598,N_249,N_160);
and U2599 (N_2599,N_2367,N_1992);
and U2600 (N_2600,N_1624,N_1691);
nor U2601 (N_2601,N_1806,N_1283);
nor U2602 (N_2602,N_1094,N_429);
nor U2603 (N_2603,N_842,N_1890);
and U2604 (N_2604,N_1934,N_2454);
or U2605 (N_2605,N_216,N_1035);
and U2606 (N_2606,N_274,N_945);
and U2607 (N_2607,N_569,N_1274);
or U2608 (N_2608,N_753,N_1429);
or U2609 (N_2609,N_133,N_2319);
and U2610 (N_2610,N_2335,N_1884);
nor U2611 (N_2611,N_1002,N_2152);
or U2612 (N_2612,N_1710,N_2280);
xnor U2613 (N_2613,N_49,N_1906);
nor U2614 (N_2614,N_351,N_2094);
nor U2615 (N_2615,N_2132,N_171);
nor U2616 (N_2616,N_805,N_1542);
or U2617 (N_2617,N_1052,N_1502);
or U2618 (N_2618,N_1336,N_2356);
xor U2619 (N_2619,N_776,N_1171);
nand U2620 (N_2620,N_750,N_44);
or U2621 (N_2621,N_2014,N_497);
or U2622 (N_2622,N_248,N_865);
or U2623 (N_2623,N_2072,N_2451);
nor U2624 (N_2624,N_1154,N_1819);
or U2625 (N_2625,N_2099,N_1729);
nor U2626 (N_2626,N_2106,N_709);
nor U2627 (N_2627,N_2003,N_1672);
or U2628 (N_2628,N_32,N_593);
nor U2629 (N_2629,N_1424,N_727);
or U2630 (N_2630,N_1487,N_170);
or U2631 (N_2631,N_224,N_434);
nand U2632 (N_2632,N_682,N_352);
nor U2633 (N_2633,N_1384,N_632);
nand U2634 (N_2634,N_453,N_2261);
and U2635 (N_2635,N_860,N_648);
or U2636 (N_2636,N_1838,N_1892);
nand U2637 (N_2637,N_1626,N_78);
or U2638 (N_2638,N_1118,N_1824);
and U2639 (N_2639,N_1999,N_2299);
or U2640 (N_2640,N_1766,N_2057);
and U2641 (N_2641,N_1818,N_2275);
and U2642 (N_2642,N_424,N_110);
or U2643 (N_2643,N_1505,N_596);
nand U2644 (N_2644,N_1544,N_1785);
nor U2645 (N_2645,N_470,N_1722);
nand U2646 (N_2646,N_1360,N_72);
and U2647 (N_2647,N_1226,N_169);
or U2648 (N_2648,N_597,N_1788);
nor U2649 (N_2649,N_1972,N_483);
or U2650 (N_2650,N_2224,N_1618);
and U2651 (N_2651,N_1021,N_490);
nand U2652 (N_2652,N_1003,N_1833);
nor U2653 (N_2653,N_18,N_172);
nand U2654 (N_2654,N_685,N_163);
or U2655 (N_2655,N_1194,N_322);
nor U2656 (N_2656,N_911,N_426);
and U2657 (N_2657,N_2402,N_2282);
xnor U2658 (N_2658,N_2085,N_982);
or U2659 (N_2659,N_125,N_1299);
or U2660 (N_2660,N_2020,N_459);
nand U2661 (N_2661,N_946,N_1664);
nor U2662 (N_2662,N_696,N_423);
or U2663 (N_2663,N_427,N_559);
nand U2664 (N_2664,N_1371,N_937);
nor U2665 (N_2665,N_2493,N_981);
nor U2666 (N_2666,N_1132,N_745);
nand U2667 (N_2667,N_1744,N_1367);
nor U2668 (N_2668,N_894,N_852);
nand U2669 (N_2669,N_2011,N_283);
and U2670 (N_2670,N_684,N_761);
nand U2671 (N_2671,N_1013,N_1850);
and U2672 (N_2672,N_2452,N_305);
or U2673 (N_2673,N_823,N_510);
and U2674 (N_2674,N_534,N_1903);
nand U2675 (N_2675,N_1178,N_2144);
or U2676 (N_2676,N_1106,N_1789);
nor U2677 (N_2677,N_1187,N_1580);
or U2678 (N_2678,N_2449,N_1770);
nand U2679 (N_2679,N_329,N_815);
and U2680 (N_2680,N_7,N_936);
nand U2681 (N_2681,N_536,N_1589);
nand U2682 (N_2682,N_109,N_551);
or U2683 (N_2683,N_93,N_636);
nor U2684 (N_2684,N_1623,N_1600);
and U2685 (N_2685,N_2055,N_1305);
nand U2686 (N_2686,N_1289,N_135);
or U2687 (N_2687,N_1945,N_517);
nor U2688 (N_2688,N_2162,N_525);
nor U2689 (N_2689,N_1866,N_2482);
nand U2690 (N_2690,N_1650,N_1817);
or U2691 (N_2691,N_1209,N_73);
nand U2692 (N_2692,N_962,N_906);
and U2693 (N_2693,N_891,N_1804);
and U2694 (N_2694,N_2462,N_1428);
and U2695 (N_2695,N_725,N_618);
xor U2696 (N_2696,N_2287,N_71);
nand U2697 (N_2697,N_1912,N_1813);
nor U2698 (N_2698,N_890,N_256);
or U2699 (N_2699,N_1946,N_1694);
or U2700 (N_2700,N_2019,N_374);
or U2701 (N_2701,N_1238,N_591);
and U2702 (N_2702,N_637,N_2096);
and U2703 (N_2703,N_1792,N_1837);
nand U2704 (N_2704,N_2120,N_1863);
or U2705 (N_2705,N_2119,N_2317);
or U2706 (N_2706,N_2093,N_122);
or U2707 (N_2707,N_760,N_1379);
and U2708 (N_2708,N_782,N_1655);
or U2709 (N_2709,N_59,N_1938);
and U2710 (N_2710,N_1730,N_1007);
nor U2711 (N_2711,N_1908,N_785);
nor U2712 (N_2712,N_691,N_1253);
and U2713 (N_2713,N_903,N_438);
nand U2714 (N_2714,N_1553,N_1860);
and U2715 (N_2715,N_623,N_1703);
and U2716 (N_2716,N_2159,N_883);
nor U2717 (N_2717,N_344,N_1558);
nor U2718 (N_2718,N_630,N_347);
or U2719 (N_2719,N_1287,N_1337);
nand U2720 (N_2720,N_1620,N_1658);
nand U2721 (N_2721,N_635,N_1244);
or U2722 (N_2722,N_315,N_335);
or U2723 (N_2723,N_1800,N_578);
nand U2724 (N_2724,N_406,N_2095);
and U2725 (N_2725,N_277,N_1566);
nor U2726 (N_2726,N_607,N_1167);
nor U2727 (N_2727,N_964,N_239);
nor U2728 (N_2728,N_1389,N_79);
and U2729 (N_2729,N_735,N_1666);
nor U2730 (N_2730,N_1232,N_1290);
or U2731 (N_2731,N_610,N_2483);
nor U2732 (N_2732,N_1536,N_612);
or U2733 (N_2733,N_1332,N_1913);
nor U2734 (N_2734,N_1909,N_1188);
or U2735 (N_2735,N_680,N_795);
nand U2736 (N_2736,N_114,N_1414);
and U2737 (N_2737,N_1086,N_396);
or U2738 (N_2738,N_1227,N_1513);
and U2739 (N_2739,N_1684,N_1764);
or U2740 (N_2740,N_1988,N_851);
nor U2741 (N_2741,N_1834,N_549);
or U2742 (N_2742,N_583,N_1587);
or U2743 (N_2743,N_614,N_1027);
or U2744 (N_2744,N_1660,N_1370);
nand U2745 (N_2745,N_579,N_1060);
nand U2746 (N_2746,N_333,N_1485);
nand U2747 (N_2747,N_872,N_1460);
or U2748 (N_2748,N_1932,N_1811);
nor U2749 (N_2749,N_1998,N_1041);
and U2750 (N_2750,N_480,N_690);
and U2751 (N_2751,N_778,N_238);
and U2752 (N_2752,N_2073,N_871);
or U2753 (N_2753,N_2068,N_1750);
nor U2754 (N_2754,N_555,N_1894);
and U2755 (N_2755,N_43,N_1474);
and U2756 (N_2756,N_222,N_2084);
and U2757 (N_2757,N_729,N_1281);
xnor U2758 (N_2758,N_1459,N_2080);
or U2759 (N_2759,N_332,N_308);
nor U2760 (N_2760,N_954,N_372);
nand U2761 (N_2761,N_780,N_460);
and U2762 (N_2762,N_451,N_2392);
or U2763 (N_2763,N_877,N_507);
or U2764 (N_2764,N_2197,N_1562);
nor U2765 (N_2765,N_1543,N_659);
and U2766 (N_2766,N_2488,N_587);
or U2767 (N_2767,N_2334,N_276);
and U2768 (N_2768,N_1886,N_411);
nor U2769 (N_2769,N_100,N_174);
nor U2770 (N_2770,N_951,N_499);
and U2771 (N_2771,N_757,N_1179);
nor U2772 (N_2772,N_1628,N_2439);
and U2773 (N_2773,N_1076,N_2363);
nand U2774 (N_2774,N_1751,N_1780);
and U2775 (N_2775,N_1991,N_1310);
nand U2776 (N_2776,N_13,N_2231);
nor U2777 (N_2777,N_826,N_754);
nor U2778 (N_2778,N_2023,N_1321);
and U2779 (N_2779,N_363,N_1432);
and U2780 (N_2780,N_2229,N_2342);
nand U2781 (N_2781,N_1368,N_651);
nand U2782 (N_2782,N_2485,N_1509);
and U2783 (N_2783,N_2258,N_1113);
or U2784 (N_2784,N_882,N_1854);
and U2785 (N_2785,N_435,N_1517);
nor U2786 (N_2786,N_1775,N_2037);
xnor U2787 (N_2787,N_688,N_2423);
and U2788 (N_2788,N_19,N_1495);
nand U2789 (N_2789,N_1112,N_893);
and U2790 (N_2790,N_526,N_1594);
nand U2791 (N_2791,N_236,N_2198);
nor U2792 (N_2792,N_2174,N_132);
and U2793 (N_2793,N_1071,N_1773);
nor U2794 (N_2794,N_1114,N_1207);
or U2795 (N_2795,N_1778,N_1173);
nand U2796 (N_2796,N_2150,N_1404);
nor U2797 (N_2797,N_2427,N_939);
and U2798 (N_2798,N_2283,N_1920);
or U2799 (N_2799,N_2338,N_1345);
or U2800 (N_2800,N_1492,N_2113);
or U2801 (N_2801,N_2354,N_1153);
and U2802 (N_2802,N_595,N_1823);
xor U2803 (N_2803,N_547,N_1527);
and U2804 (N_2804,N_957,N_1315);
nand U2805 (N_2805,N_2115,N_505);
or U2806 (N_2806,N_2138,N_2167);
or U2807 (N_2807,N_1411,N_1254);
nand U2808 (N_2808,N_2059,N_2286);
and U2809 (N_2809,N_1058,N_1133);
and U2810 (N_2810,N_2271,N_1774);
nand U2811 (N_2811,N_1358,N_1771);
nor U2812 (N_2812,N_1149,N_2406);
nor U2813 (N_2813,N_2408,N_1239);
and U2814 (N_2814,N_699,N_1196);
xor U2815 (N_2815,N_2012,N_123);
xor U2816 (N_2816,N_1549,N_1067);
and U2817 (N_2817,N_1166,N_2273);
and U2818 (N_2818,N_2002,N_1302);
nand U2819 (N_2819,N_1947,N_2213);
and U2820 (N_2820,N_2021,N_1291);
nor U2821 (N_2821,N_1425,N_1462);
nor U2822 (N_2822,N_1169,N_989);
nand U2823 (N_2823,N_2036,N_1520);
or U2824 (N_2824,N_1607,N_592);
and U2825 (N_2825,N_314,N_506);
and U2826 (N_2826,N_1718,N_2348);
and U2827 (N_2827,N_62,N_724);
and U2828 (N_2828,N_217,N_970);
and U2829 (N_2829,N_972,N_2421);
and U2830 (N_2830,N_1000,N_442);
nand U2831 (N_2831,N_410,N_74);
nand U2832 (N_2832,N_10,N_2425);
nand U2833 (N_2833,N_950,N_1008);
nand U2834 (N_2834,N_1142,N_1627);
nor U2835 (N_2835,N_879,N_1791);
nor U2836 (N_2836,N_995,N_1723);
nand U2837 (N_2837,N_1403,N_1482);
or U2838 (N_2838,N_1610,N_2383);
and U2839 (N_2839,N_2031,N_2330);
or U2840 (N_2840,N_1784,N_1540);
or U2841 (N_2841,N_849,N_394);
and U2842 (N_2842,N_444,N_1301);
and U2843 (N_2843,N_606,N_734);
xnor U2844 (N_2844,N_1264,N_334);
nand U2845 (N_2845,N_141,N_1852);
nor U2846 (N_2846,N_676,N_1634);
xnor U2847 (N_2847,N_1476,N_1256);
nand U2848 (N_2848,N_1511,N_1588);
nor U2849 (N_2849,N_2446,N_75);
nor U2850 (N_2850,N_2089,N_475);
nand U2851 (N_2851,N_1599,N_963);
or U2852 (N_2852,N_1061,N_552);
or U2853 (N_2853,N_67,N_1574);
nor U2854 (N_2854,N_2110,N_1969);
nor U2855 (N_2855,N_731,N_966);
or U2856 (N_2856,N_1240,N_2434);
and U2857 (N_2857,N_1539,N_223);
nand U2858 (N_2858,N_252,N_1342);
or U2859 (N_2859,N_837,N_1706);
nor U2860 (N_2860,N_1409,N_2191);
and U2861 (N_2861,N_838,N_2416);
xor U2862 (N_2862,N_96,N_983);
or U2863 (N_2863,N_948,N_771);
or U2864 (N_2864,N_298,N_2081);
nor U2865 (N_2865,N_752,N_1612);
nand U2866 (N_2866,N_870,N_293);
nor U2867 (N_2867,N_590,N_2166);
and U2868 (N_2868,N_1355,N_2424);
or U2869 (N_2869,N_2188,N_437);
nand U2870 (N_2870,N_542,N_289);
nand U2871 (N_2871,N_147,N_1447);
nor U2872 (N_2872,N_1268,N_1144);
nand U2873 (N_2873,N_652,N_504);
or U2874 (N_2874,N_382,N_1883);
nor U2875 (N_2875,N_1349,N_177);
or U2876 (N_2876,N_658,N_2108);
nand U2877 (N_2877,N_1097,N_1897);
nor U2878 (N_2878,N_1559,N_998);
xor U2879 (N_2879,N_1961,N_829);
nor U2880 (N_2880,N_1557,N_2433);
or U2881 (N_2881,N_1943,N_1224);
or U2882 (N_2882,N_1847,N_1929);
or U2883 (N_2883,N_1435,N_2123);
nand U2884 (N_2884,N_885,N_1421);
nor U2885 (N_2885,N_1625,N_116);
nor U2886 (N_2886,N_1306,N_447);
nand U2887 (N_2887,N_88,N_1713);
and U2888 (N_2888,N_391,N_2480);
and U2889 (N_2889,N_647,N_518);
or U2890 (N_2890,N_790,N_566);
nor U2891 (N_2891,N_2496,N_461);
or U2892 (N_2892,N_1176,N_866);
nor U2893 (N_2893,N_1401,N_138);
nor U2894 (N_2894,N_303,N_2304);
nor U2895 (N_2895,N_2418,N_921);
nor U2896 (N_2896,N_2314,N_2495);
and U2897 (N_2897,N_1867,N_2364);
or U2898 (N_2898,N_1155,N_1592);
xor U2899 (N_2899,N_1616,N_330);
and U2900 (N_2900,N_1339,N_1640);
and U2901 (N_2901,N_548,N_1463);
or U2902 (N_2902,N_1236,N_1701);
nand U2903 (N_2903,N_1,N_2475);
nand U2904 (N_2904,N_986,N_253);
and U2905 (N_2905,N_2373,N_2291);
or U2906 (N_2906,N_1590,N_1395);
nand U2907 (N_2907,N_2463,N_2388);
or U2908 (N_2908,N_1025,N_1575);
or U2909 (N_2909,N_1190,N_581);
and U2910 (N_2910,N_1888,N_2127);
or U2911 (N_2911,N_2403,N_68);
nor U2912 (N_2912,N_1796,N_430);
and U2913 (N_2913,N_360,N_1601);
xnor U2914 (N_2914,N_422,N_687);
nor U2915 (N_2915,N_467,N_2399);
or U2916 (N_2916,N_2444,N_1031);
nor U2917 (N_2917,N_1406,N_1045);
nor U2918 (N_2918,N_234,N_988);
or U2919 (N_2919,N_1245,N_875);
or U2920 (N_2920,N_2220,N_1662);
or U2921 (N_2921,N_500,N_2432);
or U2922 (N_2922,N_1830,N_111);
nor U2923 (N_2923,N_1068,N_482);
and U2924 (N_2924,N_1152,N_205);
nand U2925 (N_2925,N_41,N_2048);
nor U2926 (N_2926,N_1790,N_994);
nor U2927 (N_2927,N_1164,N_1102);
or U2928 (N_2928,N_227,N_2254);
and U2929 (N_2929,N_2369,N_1159);
and U2930 (N_2930,N_1083,N_2443);
or U2931 (N_2931,N_2058,N_2400);
nand U2932 (N_2932,N_929,N_927);
and U2933 (N_2933,N_2,N_1156);
or U2934 (N_2934,N_1935,N_1080);
and U2935 (N_2935,N_2064,N_450);
nand U2936 (N_2936,N_2461,N_2226);
nand U2937 (N_2937,N_859,N_1096);
or U2938 (N_2938,N_908,N_613);
or U2939 (N_2939,N_2333,N_1091);
nand U2940 (N_2940,N_2217,N_1974);
or U2941 (N_2941,N_1265,N_1392);
or U2942 (N_2942,N_2232,N_1758);
or U2943 (N_2943,N_1944,N_1203);
and U2944 (N_2944,N_2289,N_1017);
and U2945 (N_2945,N_2328,N_763);
nor U2946 (N_2946,N_711,N_1719);
nand U2947 (N_2947,N_1259,N_1250);
and U2948 (N_2948,N_1656,N_575);
nand U2949 (N_2949,N_2121,N_1644);
nand U2950 (N_2950,N_180,N_370);
nor U2951 (N_2951,N_2184,N_1488);
nand U2952 (N_2952,N_649,N_1220);
xnor U2953 (N_2953,N_1712,N_2397);
nor U2954 (N_2954,N_965,N_1964);
or U2955 (N_2955,N_1262,N_1347);
or U2956 (N_2956,N_2103,N_993);
nor U2957 (N_2957,N_917,N_1018);
nand U2958 (N_2958,N_242,N_601);
nand U2959 (N_2959,N_97,N_1327);
nor U2960 (N_2960,N_431,N_1569);
nand U2961 (N_2961,N_387,N_1093);
or U2962 (N_2962,N_1394,N_1251);
or U2963 (N_2963,N_1016,N_1416);
nor U2964 (N_2964,N_197,N_1603);
nand U2965 (N_2965,N_474,N_747);
or U2966 (N_2966,N_389,N_611);
nand U2967 (N_2967,N_759,N_2247);
and U2968 (N_2968,N_794,N_1252);
and U2969 (N_2969,N_466,N_765);
and U2970 (N_2970,N_388,N_1523);
nor U2971 (N_2971,N_22,N_973);
and U2972 (N_2972,N_617,N_830);
or U2973 (N_2973,N_1975,N_1285);
and U2974 (N_2974,N_1326,N_1891);
and U2975 (N_2975,N_1716,N_1145);
nor U2976 (N_2976,N_1896,N_1449);
nor U2977 (N_2977,N_1341,N_1911);
nand U2978 (N_2978,N_924,N_631);
nand U2979 (N_2979,N_2478,N_1516);
nor U2980 (N_2980,N_1519,N_1936);
or U2981 (N_2981,N_449,N_2118);
and U2982 (N_2982,N_1352,N_425);
or U2983 (N_2983,N_1518,N_1538);
nand U2984 (N_2984,N_2378,N_1776);
nand U2985 (N_2985,N_2201,N_589);
xor U2986 (N_2986,N_1604,N_1258);
nor U2987 (N_2987,N_626,N_2491);
and U2988 (N_2988,N_1848,N_201);
or U2989 (N_2989,N_2389,N_1772);
or U2990 (N_2990,N_675,N_841);
or U2991 (N_2991,N_2368,N_878);
or U2992 (N_2992,N_2376,N_1478);
xor U2993 (N_2993,N_2460,N_2343);
nand U2994 (N_2994,N_1278,N_2029);
or U2995 (N_2995,N_1271,N_1514);
nor U2996 (N_2996,N_1698,N_1231);
nand U2997 (N_2997,N_650,N_2172);
nand U2998 (N_2998,N_1827,N_38);
or U2999 (N_2999,N_1637,N_777);
and U3000 (N_3000,N_2212,N_1917);
nor U3001 (N_3001,N_271,N_2207);
and U3002 (N_3002,N_1431,N_1351);
or U3003 (N_3003,N_755,N_1415);
or U3004 (N_3004,N_799,N_2295);
nor U3005 (N_3005,N_113,N_343);
nor U3006 (N_3006,N_1746,N_2494);
and U3007 (N_3007,N_2061,N_83);
nor U3008 (N_3008,N_1552,N_2404);
or U3009 (N_3009,N_1554,N_2079);
nand U3010 (N_3010,N_1593,N_887);
and U3011 (N_3011,N_899,N_2320);
nor U3012 (N_3012,N_1328,N_60);
and U3013 (N_3013,N_432,N_456);
nor U3014 (N_3014,N_336,N_2026);
nand U3015 (N_3015,N_925,N_50);
or U3016 (N_3016,N_373,N_1304);
nor U3017 (N_3017,N_1137,N_2297);
and U3018 (N_3018,N_165,N_1905);
or U3019 (N_3019,N_1642,N_1717);
or U3020 (N_3020,N_5,N_905);
nand U3021 (N_3021,N_421,N_511);
nand U3022 (N_3022,N_1099,N_2185);
and U3023 (N_3023,N_813,N_1261);
nand U3024 (N_3024,N_1690,N_1748);
and U3025 (N_3025,N_1700,N_1633);
and U3026 (N_3026,N_1125,N_1201);
and U3027 (N_3027,N_2240,N_20);
or U3028 (N_3028,N_1950,N_1380);
or U3029 (N_3029,N_1397,N_713);
nor U3030 (N_3030,N_1985,N_1507);
nand U3031 (N_3031,N_524,N_2340);
and U3032 (N_3032,N_812,N_2200);
or U3033 (N_3033,N_1388,N_1454);
nand U3034 (N_3034,N_2006,N_2267);
nor U3035 (N_3035,N_571,N_58);
and U3036 (N_3036,N_2306,N_1054);
nor U3037 (N_3037,N_1275,N_708);
nand U3038 (N_3038,N_484,N_828);
nand U3039 (N_3039,N_281,N_1498);
nand U3040 (N_3040,N_1100,N_2413);
or U3041 (N_3041,N_620,N_237);
and U3042 (N_3042,N_573,N_1387);
and U3043 (N_3043,N_668,N_76);
and U3044 (N_3044,N_2417,N_1731);
nand U3045 (N_3045,N_1427,N_2412);
and U3046 (N_3046,N_1329,N_1128);
and U3047 (N_3047,N_1065,N_1859);
nor U3048 (N_3048,N_2134,N_1313);
nand U3049 (N_3049,N_1526,N_931);
nand U3050 (N_3050,N_401,N_2035);
nand U3051 (N_3051,N_1444,N_624);
or U3052 (N_3052,N_2146,N_809);
and U3053 (N_3053,N_119,N_2010);
and U3054 (N_3054,N_2042,N_145);
nand U3055 (N_3055,N_2265,N_539);
nand U3056 (N_3056,N_784,N_1191);
nand U3057 (N_3057,N_2358,N_707);
and U3058 (N_3058,N_1165,N_868);
nand U3059 (N_3059,N_1276,N_831);
xor U3060 (N_3060,N_1874,N_1222);
nand U3061 (N_3061,N_1343,N_928);
or U3062 (N_3062,N_971,N_1742);
nand U3063 (N_3063,N_383,N_2250);
or U3064 (N_3064,N_619,N_189);
or U3065 (N_3065,N_522,N_1849);
or U3066 (N_3066,N_1033,N_585);
nor U3067 (N_3067,N_586,N_2324);
nor U3068 (N_3068,N_2448,N_1087);
or U3069 (N_3069,N_909,N_2431);
and U3070 (N_3070,N_857,N_358);
nor U3071 (N_3071,N_808,N_266);
nand U3072 (N_3072,N_1204,N_904);
and U3073 (N_3073,N_226,N_1237);
nand U3074 (N_3074,N_1647,N_2109);
or U3075 (N_3075,N_2453,N_584);
or U3076 (N_3076,N_3,N_468);
or U3077 (N_3077,N_2419,N_692);
or U3078 (N_3078,N_1386,N_974);
nand U3079 (N_3079,N_1798,N_732);
nand U3080 (N_3080,N_509,N_600);
and U3081 (N_3081,N_673,N_310);
nand U3082 (N_3082,N_2442,N_816);
or U3083 (N_3083,N_2393,N_1243);
and U3084 (N_3084,N_1996,N_1410);
nand U3085 (N_3085,N_1762,N_736);
or U3086 (N_3086,N_546,N_1967);
nand U3087 (N_3087,N_2303,N_472);
or U3088 (N_3088,N_2017,N_2411);
nand U3089 (N_3089,N_2228,N_2457);
and U3090 (N_3090,N_112,N_2051);
and U3091 (N_3091,N_1545,N_1810);
nor U3092 (N_3092,N_689,N_2294);
nor U3093 (N_3093,N_179,N_669);
or U3094 (N_3094,N_2125,N_2049);
nor U3095 (N_3095,N_1407,N_1445);
or U3096 (N_3096,N_1895,N_1877);
and U3097 (N_3097,N_290,N_1012);
and U3098 (N_3098,N_339,N_212);
nor U3099 (N_3099,N_665,N_2053);
or U3100 (N_3100,N_220,N_134);
or U3101 (N_3101,N_1697,N_99);
and U3102 (N_3102,N_553,N_2398);
and U3103 (N_3103,N_653,N_791);
and U3104 (N_3104,N_1466,N_2045);
nor U3105 (N_3105,N_2429,N_1405);
and U3106 (N_3106,N_105,N_2445);
nor U3107 (N_3107,N_36,N_1032);
nor U3108 (N_3108,N_366,N_1103);
and U3109 (N_3109,N_2251,N_1699);
nor U3110 (N_3110,N_1311,N_670);
and U3111 (N_3111,N_543,N_1669);
nor U3112 (N_3112,N_284,N_1024);
and U3113 (N_3113,N_2479,N_309);
and U3114 (N_3114,N_1676,N_2346);
xnor U3115 (N_3115,N_1465,N_2301);
and U3116 (N_3116,N_1186,N_2322);
and U3117 (N_3117,N_323,N_1753);
nand U3118 (N_3118,N_1212,N_722);
nand U3119 (N_3119,N_1995,N_1479);
or U3120 (N_3120,N_562,N_1374);
nor U3121 (N_3121,N_561,N_1714);
nand U3122 (N_3122,N_603,N_471);
or U3123 (N_3123,N_2276,N_1815);
or U3124 (N_3124,N_1752,N_2069);
nor U3125 (N_3125,N_889,N_1170);
or U3126 (N_3126,N_1111,N_822);
nor U3127 (N_3127,N_1635,N_2292);
and U3128 (N_3128,N_2236,N_1418);
and U3129 (N_3129,N_2088,N_835);
nand U3130 (N_3130,N_1889,N_337);
and U3131 (N_3131,N_1812,N_1257);
nor U3132 (N_3132,N_47,N_302);
and U3133 (N_3133,N_1715,N_318);
nor U3134 (N_3134,N_1303,N_629);
nor U3135 (N_3135,N_942,N_1597);
nor U3136 (N_3136,N_312,N_1537);
and U3137 (N_3137,N_1885,N_1399);
nand U3138 (N_3138,N_30,N_1085);
nor U3139 (N_3139,N_661,N_463);
or U3140 (N_3140,N_1221,N_1057);
or U3141 (N_3141,N_540,N_1591);
nor U3142 (N_3142,N_2362,N_902);
nor U3143 (N_3143,N_1182,N_1861);
nand U3144 (N_3144,N_1119,N_2311);
or U3145 (N_3145,N_523,N_2143);
nor U3146 (N_3146,N_634,N_1862);
and U3147 (N_3147,N_953,N_2215);
or U3148 (N_3148,N_2202,N_2395);
nand U3149 (N_3149,N_1362,N_856);
and U3150 (N_3150,N_935,N_1734);
nor U3151 (N_3151,N_465,N_1596);
or U3152 (N_3152,N_1582,N_1450);
nor U3153 (N_3153,N_2117,N_80);
or U3154 (N_3154,N_282,N_2153);
or U3155 (N_3155,N_1583,N_2194);
or U3156 (N_3156,N_263,N_2259);
nand U3157 (N_3157,N_1151,N_1140);
or U3158 (N_3158,N_2170,N_770);
or U3159 (N_3159,N_968,N_1483);
nand U3160 (N_3160,N_807,N_2242);
or U3161 (N_3161,N_1063,N_796);
and U3162 (N_3162,N_1300,N_231);
nor U3163 (N_3163,N_1348,N_311);
and U3164 (N_3164,N_1668,N_528);
and U3165 (N_3165,N_720,N_992);
or U3166 (N_3166,N_199,N_1185);
nand U3167 (N_3167,N_2481,N_2107);
and U3168 (N_3168,N_1745,N_545);
and U3169 (N_3169,N_1228,N_2307);
and U3170 (N_3170,N_1500,N_386);
and U3171 (N_3171,N_1469,N_1506);
nor U3172 (N_3172,N_2401,N_362);
and U3173 (N_3173,N_1131,N_932);
nor U3174 (N_3174,N_1423,N_847);
nor U3175 (N_3175,N_1019,N_1869);
nor U3176 (N_3176,N_1997,N_1331);
nand U3177 (N_3177,N_1737,N_2052);
nand U3178 (N_3178,N_538,N_115);
nor U3179 (N_3179,N_824,N_1828);
nor U3180 (N_3180,N_55,N_991);
nand U3181 (N_3181,N_895,N_1309);
and U3182 (N_3182,N_2187,N_1267);
nand U3183 (N_3183,N_839,N_967);
or U3184 (N_3184,N_2347,N_628);
nand U3185 (N_3185,N_1678,N_2219);
and U3186 (N_3186,N_486,N_858);
or U3187 (N_3187,N_1079,N_1216);
nand U3188 (N_3188,N_285,N_301);
or U3189 (N_3189,N_377,N_783);
nor U3190 (N_3190,N_2394,N_353);
and U3191 (N_3191,N_2189,N_1437);
nor U3192 (N_3192,N_714,N_1396);
nand U3193 (N_3193,N_208,N_1088);
or U3194 (N_3194,N_2135,N_81);
and U3195 (N_3195,N_1266,N_2223);
xor U3196 (N_3196,N_2160,N_494);
and U3197 (N_3197,N_241,N_1736);
nor U3198 (N_3198,N_1942,N_681);
or U3199 (N_3199,N_2210,N_103);
nor U3200 (N_3200,N_1652,N_148);
nand U3201 (N_3201,N_1208,N_2235);
nand U3202 (N_3202,N_2490,N_1585);
or U3203 (N_3203,N_556,N_2140);
or U3204 (N_3204,N_1757,N_873);
and U3205 (N_3205,N_1160,N_996);
nor U3206 (N_3206,N_1458,N_1904);
or U3207 (N_3207,N_574,N_1047);
nor U3208 (N_3208,N_1009,N_1317);
nand U3209 (N_3209,N_65,N_259);
nand U3210 (N_3210,N_1001,N_1197);
nor U3211 (N_3211,N_627,N_2284);
nand U3212 (N_3212,N_1937,N_35);
and U3213 (N_3213,N_643,N_1448);
or U3214 (N_3214,N_260,N_639);
and U3215 (N_3215,N_1322,N_1515);
and U3216 (N_3216,N_1955,N_1548);
nand U3217 (N_3217,N_622,N_1728);
or U3218 (N_3218,N_454,N_327);
or U3219 (N_3219,N_2151,N_1689);
nor U3220 (N_3220,N_1787,N_715);
and U3221 (N_3221,N_2366,N_1193);
nand U3222 (N_3222,N_1966,N_1177);
nand U3223 (N_3223,N_737,N_1056);
nand U3224 (N_3224,N_1366,N_1783);
nor U3225 (N_3225,N_979,N_2139);
nor U3226 (N_3226,N_1682,N_1475);
nor U3227 (N_3227,N_1420,N_439);
xnor U3228 (N_3228,N_863,N_1641);
and U3229 (N_3229,N_743,N_1576);
and U3230 (N_3230,N_265,N_1821);
nor U3231 (N_3231,N_1412,N_2141);
nand U3232 (N_3232,N_602,N_850);
and U3233 (N_3233,N_2377,N_1359);
or U3234 (N_3234,N_2128,N_1696);
or U3235 (N_3235,N_717,N_82);
nand U3236 (N_3236,N_1980,N_1034);
nand U3237 (N_3237,N_107,N_1755);
nor U3238 (N_3238,N_51,N_914);
or U3239 (N_3239,N_136,N_1971);
and U3240 (N_3240,N_295,N_1674);
or U3241 (N_3241,N_464,N_487);
or U3242 (N_3242,N_2471,N_881);
nand U3243 (N_3243,N_697,N_28);
or U3244 (N_3244,N_2149,N_861);
nand U3245 (N_3245,N_2436,N_1486);
and U3246 (N_3246,N_2447,N_744);
or U3247 (N_3247,N_198,N_640);
or U3248 (N_3248,N_1286,N_195);
or U3249 (N_3249,N_1130,N_1629);
nor U3250 (N_3250,N_1335,N_550);
nor U3251 (N_3251,N_1098,N_832);
xor U3252 (N_3252,N_1928,N_739);
nor U3253 (N_3253,N_1615,N_997);
nand U3254 (N_3254,N_1363,N_1398);
and U3255 (N_3255,N_646,N_1738);
or U3256 (N_3256,N_541,N_633);
nand U3257 (N_3257,N_436,N_2030);
nor U3258 (N_3258,N_1879,N_1779);
nand U3259 (N_3259,N_834,N_1782);
or U3260 (N_3260,N_2136,N_264);
nor U3261 (N_3261,N_1686,N_92);
nor U3262 (N_3262,N_2409,N_959);
or U3263 (N_3263,N_1039,N_2067);
nor U3264 (N_3264,N_1124,N_1174);
or U3265 (N_3265,N_884,N_1858);
and U3266 (N_3266,N_403,N_1503);
nor U3267 (N_3267,N_2233,N_2308);
nor U3268 (N_3268,N_1369,N_1073);
nand U3269 (N_3269,N_129,N_85);
nand U3270 (N_3270,N_657,N_320);
nand U3271 (N_3271,N_408,N_1754);
nor U3272 (N_3272,N_1881,N_489);
nand U3273 (N_3273,N_250,N_1857);
or U3274 (N_3274,N_2183,N_1029);
and U3275 (N_3275,N_2168,N_1464);
nand U3276 (N_3276,N_1081,N_1981);
nand U3277 (N_3277,N_1338,N_1472);
nand U3278 (N_3278,N_1101,N_577);
nor U3279 (N_3279,N_1430,N_233);
nand U3280 (N_3280,N_535,N_521);
nand U3281 (N_3281,N_2044,N_1584);
and U3282 (N_3282,N_1108,N_515);
and U3283 (N_3283,N_609,N_1129);
nor U3284 (N_3284,N_532,N_2182);
and U3285 (N_3285,N_2384,N_2489);
or U3286 (N_3286,N_2375,N_2077);
or U3287 (N_3287,N_768,N_184);
or U3288 (N_3288,N_294,N_146);
nand U3289 (N_3289,N_1822,N_1344);
nand U3290 (N_3290,N_1314,N_207);
or U3291 (N_3291,N_960,N_1075);
nand U3292 (N_3292,N_2246,N_2336);
nor U3293 (N_3293,N_399,N_1484);
nand U3294 (N_3294,N_1747,N_2033);
or U3295 (N_3295,N_1353,N_892);
nand U3296 (N_3296,N_1382,N_1146);
nand U3297 (N_3297,N_2361,N_2309);
or U3298 (N_3298,N_25,N_1835);
nand U3299 (N_3299,N_469,N_1532);
nor U3300 (N_3300,N_949,N_594);
and U3301 (N_3301,N_192,N_1667);
nor U3302 (N_3302,N_748,N_1471);
nor U3303 (N_3303,N_213,N_2175);
or U3304 (N_3304,N_2305,N_491);
nand U3305 (N_3305,N_876,N_142);
and U3306 (N_3306,N_764,N_368);
nor U3307 (N_3307,N_1206,N_2196);
nor U3308 (N_3308,N_175,N_1104);
and U3309 (N_3309,N_1192,N_307);
and U3310 (N_3310,N_1534,N_2065);
or U3311 (N_3311,N_2156,N_1659);
nor U3312 (N_3312,N_247,N_2279);
and U3313 (N_3313,N_1050,N_2391);
nand U3314 (N_3314,N_1364,N_1681);
nor U3315 (N_3315,N_121,N_1880);
or U3316 (N_3316,N_196,N_1307);
and U3317 (N_3317,N_418,N_2486);
nand U3318 (N_3318,N_2034,N_958);
nor U3319 (N_3319,N_2173,N_1442);
nand U3320 (N_3320,N_348,N_1832);
and U3321 (N_3321,N_1931,N_1077);
xnor U3322 (N_3322,N_1158,N_2396);
or U3323 (N_3323,N_2015,N_2326);
and U3324 (N_3324,N_2163,N_409);
or U3325 (N_3325,N_159,N_1372);
nand U3326 (N_3326,N_452,N_194);
or U3327 (N_3327,N_1578,N_1965);
nand U3328 (N_3328,N_182,N_1825);
nand U3329 (N_3329,N_1794,N_209);
and U3330 (N_3330,N_94,N_956);
and U3331 (N_3331,N_1434,N_1577);
or U3332 (N_3332,N_2078,N_130);
nand U3333 (N_3333,N_730,N_2157);
and U3334 (N_3334,N_1443,N_1856);
or U3335 (N_3335,N_1611,N_1053);
nand U3336 (N_3336,N_2321,N_1436);
or U3337 (N_3337,N_1298,N_2100);
nand U3338 (N_3338,N_913,N_225);
and U3339 (N_3339,N_1233,N_984);
nor U3340 (N_3340,N_1294,N_297);
nand U3341 (N_3341,N_1685,N_1136);
nor U3342 (N_3342,N_385,N_384);
nor U3343 (N_3343,N_1653,N_1573);
or U3344 (N_3344,N_1117,N_1116);
or U3345 (N_3345,N_128,N_1277);
or U3346 (N_3346,N_124,N_1383);
nor U3347 (N_3347,N_2430,N_1038);
and U3348 (N_3348,N_2155,N_1675);
nor U3349 (N_3349,N_1550,N_2176);
and U3350 (N_3350,N_1864,N_2126);
nor U3351 (N_3351,N_272,N_1189);
nor U3352 (N_3352,N_848,N_798);
and U3353 (N_3353,N_2039,N_286);
or U3354 (N_3354,N_2492,N_1951);
or U3355 (N_3355,N_2204,N_167);
nor U3356 (N_3356,N_1665,N_1630);
and U3357 (N_3357,N_686,N_2407);
nand U3358 (N_3358,N_299,N_1683);
and U3359 (N_3359,N_1602,N_397);
and U3360 (N_3360,N_1319,N_187);
or U3361 (N_3361,N_369,N_2435);
and U3362 (N_3362,N_1456,N_1581);
or U3363 (N_3363,N_1062,N_1878);
or U3364 (N_3364,N_1183,N_244);
or U3365 (N_3365,N_2112,N_86);
and U3366 (N_3366,N_1026,N_615);
and U3367 (N_3367,N_2016,N_1473);
and U3368 (N_3368,N_395,N_1870);
nor U3369 (N_3369,N_1011,N_1648);
and U3370 (N_3370,N_455,N_446);
nor U3371 (N_3371,N_787,N_1643);
nand U3372 (N_3372,N_762,N_2007);
nand U3373 (N_3373,N_2355,N_2263);
xor U3374 (N_3374,N_853,N_679);
xor U3375 (N_3375,N_361,N_2114);
nand U3376 (N_3376,N_738,N_1632);
or U3377 (N_3377,N_1121,N_656);
and U3378 (N_3378,N_1092,N_193);
and U3379 (N_3379,N_2190,N_1356);
nor U3380 (N_3380,N_183,N_278);
nor U3381 (N_3381,N_1350,N_2090);
or U3382 (N_3382,N_1340,N_2437);
or U3383 (N_3383,N_2142,N_2313);
nand U3384 (N_3384,N_2274,N_1807);
nor U3385 (N_3385,N_1175,N_1107);
or U3386 (N_3386,N_2071,N_2315);
nor U3387 (N_3387,N_645,N_2216);
nand U3388 (N_3388,N_139,N_1512);
and U3389 (N_3389,N_2264,N_356);
nand U3390 (N_3390,N_12,N_1014);
nand U3391 (N_3391,N_821,N_1426);
nor U3392 (N_3392,N_598,N_2255);
or U3393 (N_3393,N_1876,N_2464);
nor U3394 (N_3394,N_462,N_2296);
nor U3395 (N_3395,N_797,N_153);
and U3396 (N_3396,N_321,N_1765);
and U3397 (N_3397,N_2472,N_1249);
or U3398 (N_3398,N_1272,N_1150);
or U3399 (N_3399,N_2352,N_1028);
and U3400 (N_3400,N_810,N_1919);
and U3401 (N_3401,N_2122,N_1839);
nor U3402 (N_3402,N_1004,N_2323);
and U3403 (N_3403,N_1489,N_666);
nor U3404 (N_3404,N_221,N_1330);
and U3405 (N_3405,N_2310,N_1541);
or U3406 (N_3406,N_1688,N_1433);
and U3407 (N_3407,N_1809,N_1987);
and U3408 (N_3408,N_1417,N_1134);
or U3409 (N_3409,N_1082,N_1907);
nor U3410 (N_3410,N_1439,N_1422);
and U3411 (N_3411,N_767,N_2459);
nand U3412 (N_3412,N_1524,N_537);
nor U3413 (N_3413,N_1241,N_846);
nand U3414 (N_3414,N_704,N_2381);
nor U3415 (N_3415,N_2372,N_2199);
nor U3416 (N_3416,N_2004,N_1385);
nor U3417 (N_3417,N_1663,N_1127);
nor U3418 (N_3418,N_16,N_1419);
nand U3419 (N_3419,N_1933,N_1962);
nand U3420 (N_3420,N_742,N_1831);
nand U3421 (N_3421,N_825,N_803);
nand U3422 (N_3422,N_2018,N_2050);
or U3423 (N_3423,N_144,N_1900);
or U3424 (N_3424,N_1280,N_1563);
and U3425 (N_3425,N_42,N_1708);
or U3426 (N_3426,N_87,N_152);
nor U3427 (N_3427,N_2357,N_229);
nand U3428 (N_3428,N_897,N_678);
or U3429 (N_3429,N_2124,N_941);
nor U3430 (N_3430,N_2476,N_1609);
nand U3431 (N_3431,N_1741,N_2009);
or U3432 (N_3432,N_1055,N_2027);
or U3433 (N_3433,N_1391,N_267);
nand U3434 (N_3434,N_1470,N_2466);
and U3435 (N_3435,N_2091,N_558);
or U3436 (N_3436,N_2063,N_1836);
and U3437 (N_3437,N_2203,N_985);
and U3438 (N_3438,N_306,N_375);
xor U3439 (N_3439,N_381,N_2382);
nor U3440 (N_3440,N_1777,N_2458);
and U3441 (N_3441,N_2230,N_485);
or U3442 (N_3442,N_1670,N_1560);
or U3443 (N_3443,N_502,N_746);
or U3444 (N_3444,N_1940,N_2327);
or U3445 (N_3445,N_2477,N_1376);
nand U3446 (N_3446,N_1720,N_940);
nand U3447 (N_3447,N_802,N_1899);
nand U3448 (N_3448,N_886,N_324);
nand U3449 (N_3449,N_417,N_554);
or U3450 (N_3450,N_1242,N_1893);
or U3451 (N_3451,N_412,N_1984);
nor U3452 (N_3452,N_1234,N_2208);
or U3453 (N_3453,N_2179,N_270);
nor U3454 (N_3454,N_1036,N_479);
nand U3455 (N_3455,N_1408,N_1297);
or U3456 (N_3456,N_84,N_1293);
and U3457 (N_3457,N_2056,N_313);
or U3458 (N_3458,N_2192,N_1269);
and U3459 (N_3459,N_1493,N_393);
and U3460 (N_3460,N_2032,N_1521);
or U3461 (N_3461,N_900,N_154);
nor U3462 (N_3462,N_1260,N_1957);
or U3463 (N_3463,N_1090,N_89);
nor U3464 (N_3464,N_1726,N_1989);
xnor U3465 (N_3465,N_254,N_1724);
nand U3466 (N_3466,N_1651,N_2130);
nor U3467 (N_3467,N_1556,N_520);
xor U3468 (N_3468,N_1205,N_2262);
nand U3469 (N_3469,N_1141,N_944);
or U3470 (N_3470,N_1037,N_1761);
and U3471 (N_3471,N_918,N_1586);
nand U3472 (N_3472,N_1440,N_61);
nand U3473 (N_3473,N_288,N_1816);
or U3474 (N_3474,N_2087,N_844);
and U3475 (N_3475,N_1606,N_2104);
nor U3476 (N_3476,N_1400,N_1845);
nand U3477 (N_3477,N_2193,N_53);
or U3478 (N_3478,N_1235,N_1927);
nor U3479 (N_3479,N_2066,N_2145);
and U3480 (N_3480,N_168,N_1983);
and U3481 (N_3481,N_2186,N_1468);
nor U3482 (N_3482,N_1452,N_801);
nor U3483 (N_3483,N_888,N_1095);
or U3484 (N_3484,N_26,N_27);
and U3485 (N_3485,N_2177,N_2484);
nand U3486 (N_3486,N_215,N_568);
and U3487 (N_3487,N_1756,N_947);
or U3488 (N_3488,N_2098,N_331);
and U3489 (N_3489,N_930,N_2206);
nor U3490 (N_3490,N_910,N_428);
nor U3491 (N_3491,N_644,N_1568);
nor U3492 (N_3492,N_2038,N_1739);
and U3493 (N_3493,N_642,N_1390);
xor U3494 (N_3494,N_1561,N_2441);
and U3495 (N_3495,N_317,N_2097);
or U3496 (N_3496,N_473,N_2260);
and U3497 (N_3497,N_1213,N_52);
or U3498 (N_3498,N_1763,N_2147);
nor U3499 (N_3499,N_1608,N_952);
and U3500 (N_3500,N_2164,N_1069);
or U3501 (N_3501,N_2005,N_758);
or U3502 (N_3502,N_1346,N_66);
nor U3503 (N_3503,N_120,N_1225);
or U3504 (N_3504,N_214,N_173);
or U3505 (N_3505,N_1749,N_203);
or U3506 (N_3506,N_457,N_922);
and U3507 (N_3507,N_2288,N_980);
or U3508 (N_3508,N_258,N_2277);
or U3509 (N_3509,N_1496,N_2470);
and U3510 (N_3510,N_2022,N_1882);
nor U3511 (N_3511,N_2499,N_1799);
and U3512 (N_3512,N_280,N_419);
nand U3513 (N_3513,N_364,N_775);
nand U3514 (N_3514,N_2086,N_1357);
xor U3515 (N_3515,N_2281,N_1248);
or U3516 (N_3516,N_1973,N_926);
and U3517 (N_3517,N_1499,N_2040);
nor U3518 (N_3518,N_1803,N_1693);
nand U3519 (N_3519,N_1497,N_862);
nand U3520 (N_3520,N_1147,N_1918);
nand U3521 (N_3521,N_2316,N_1707);
and U3522 (N_3522,N_2161,N_2171);
or U3523 (N_3523,N_912,N_915);
or U3524 (N_3524,N_1970,N_2148);
xnor U3525 (N_3525,N_240,N_1015);
and U3526 (N_3526,N_104,N_304);
or U3527 (N_3527,N_1282,N_773);
nand U3528 (N_3528,N_664,N_1855);
nand U3529 (N_3529,N_77,N_766);
nand U3530 (N_3530,N_1022,N_2178);
nand U3531 (N_3531,N_2497,N_378);
nor U3532 (N_3532,N_1564,N_1924);
and U3533 (N_3533,N_261,N_1679);
nand U3534 (N_3534,N_655,N_34);
or U3535 (N_3535,N_529,N_2331);
or U3536 (N_3536,N_1871,N_1711);
nor U3537 (N_3537,N_2024,N_210);
nand U3538 (N_3538,N_503,N_2272);
nor U3539 (N_3539,N_1820,N_1546);
or U3540 (N_3540,N_106,N_740);
nand U3541 (N_3541,N_1994,N_1161);
or U3542 (N_3542,N_977,N_2205);
nand U3543 (N_3543,N_1070,N_1273);
and U3544 (N_3544,N_1781,N_102);
or U3545 (N_3545,N_1567,N_354);
or U3546 (N_3546,N_990,N_292);
or U3547 (N_3547,N_694,N_781);
or U3548 (N_3548,N_1120,N_1049);
nand U3549 (N_3549,N_365,N_901);
and U3550 (N_3550,N_818,N_1501);
nor U3551 (N_3551,N_1732,N_1453);
nand U3552 (N_3552,N_443,N_1195);
and U3553 (N_3553,N_496,N_2450);
nor U3554 (N_3554,N_923,N_1760);
and U3555 (N_3555,N_1143,N_2046);
nand U3556 (N_3556,N_576,N_477);
and U3557 (N_3557,N_2062,N_2041);
nor U3558 (N_3558,N_1072,N_880);
nand U3559 (N_3559,N_1795,N_2278);
nor U3560 (N_3560,N_40,N_2374);
nor U3561 (N_3561,N_1963,N_1645);
or U3562 (N_3562,N_2243,N_786);
or U3563 (N_3563,N_793,N_1923);
and U3564 (N_3564,N_1939,N_1528);
or U3565 (N_3565,N_519,N_1381);
nand U3566 (N_3566,N_1727,N_359);
nand U3567 (N_3567,N_2298,N_1284);
or U3568 (N_3568,N_156,N_2218);
nand U3569 (N_3569,N_1733,N_355);
nor U3570 (N_3570,N_95,N_721);
and U3571 (N_3571,N_1572,N_1547);
and U3572 (N_3572,N_1579,N_933);
and U3573 (N_3573,N_1705,N_1296);
and U3574 (N_3574,N_560,N_433);
and U3575 (N_3575,N_2054,N_161);
or U3576 (N_3576,N_279,N_1571);
or U3577 (N_3577,N_2060,N_2131);
nor U3578 (N_3578,N_2241,N_127);
nor U3579 (N_3579,N_1210,N_1910);
nor U3580 (N_3580,N_2415,N_158);
and U3581 (N_3581,N_854,N_1504);
nor U3582 (N_3582,N_969,N_1373);
nor U3583 (N_3583,N_916,N_404);
or U3584 (N_3584,N_2116,N_1138);
or U3585 (N_3585,N_723,N_390);
or U3586 (N_3586,N_804,N_1157);
nand U3587 (N_3587,N_1555,N_855);
or U3588 (N_3588,N_1477,N_204);
or U3589 (N_3589,N_493,N_1126);
nand U3590 (N_3590,N_2221,N_660);
nand U3591 (N_3591,N_2214,N_976);
and U3592 (N_3592,N_1767,N_1214);
or U3593 (N_3593,N_1695,N_1115);
nand U3594 (N_3594,N_1613,N_1786);
or U3595 (N_3595,N_1802,N_2290);
nor U3596 (N_3596,N_1829,N_1510);
or U3597 (N_3597,N_2266,N_98);
xnor U3598 (N_3598,N_1110,N_570);
or U3599 (N_3599,N_33,N_2237);
and U3600 (N_3600,N_407,N_185);
and U3601 (N_3601,N_2370,N_1325);
nor U3602 (N_3602,N_1184,N_814);
or U3603 (N_3603,N_2181,N_654);
nor U3604 (N_3604,N_1814,N_1202);
nand U3605 (N_3605,N_840,N_275);
or U3606 (N_3606,N_2252,N_1565);
or U3607 (N_3607,N_1333,N_1042);
and U3608 (N_3608,N_2360,N_1617);
nor U3609 (N_3609,N_869,N_1692);
or U3610 (N_3610,N_792,N_1533);
xnor U3611 (N_3611,N_350,N_143);
xnor U3612 (N_3612,N_1467,N_1480);
nor U3613 (N_3613,N_1005,N_1230);
and U3614 (N_3614,N_677,N_273);
nor U3615 (N_3615,N_582,N_230);
or U3616 (N_3616,N_1217,N_2211);
and U3617 (N_3617,N_827,N_1263);
nand U3618 (N_3618,N_2008,N_961);
and U3619 (N_3619,N_1725,N_246);
or U3620 (N_3620,N_63,N_2410);
nor U3621 (N_3621,N_1361,N_769);
or U3622 (N_3622,N_1926,N_39);
nor U3623 (N_3623,N_1168,N_2339);
nor U3624 (N_3624,N_166,N_1887);
and U3625 (N_3625,N_1954,N_1010);
nand U3626 (N_3626,N_2351,N_513);
nand U3627 (N_3627,N_346,N_1441);
or U3628 (N_3628,N_512,N_21);
and U3629 (N_3629,N_514,N_441);
nor U3630 (N_3630,N_162,N_325);
and U3631 (N_3631,N_588,N_70);
nand U3632 (N_3632,N_1673,N_702);
nor U3633 (N_3633,N_2227,N_1365);
or U3634 (N_3634,N_2440,N_151);
nand U3635 (N_3635,N_1941,N_1105);
and U3636 (N_3636,N_508,N_176);
nor U3637 (N_3637,N_1334,N_1740);
and U3638 (N_3638,N_300,N_1402);
or U3639 (N_3639,N_819,N_2379);
nor U3640 (N_3640,N_1636,N_413);
or U3641 (N_3641,N_357,N_498);
and U3642 (N_3642,N_1639,N_1051);
nand U3643 (N_3643,N_907,N_1979);
and U3644 (N_3644,N_405,N_2455);
and U3645 (N_3645,N_1968,N_2365);
nand U3646 (N_3646,N_701,N_1952);
and U3647 (N_3647,N_1958,N_1570);
and U3648 (N_3648,N_1446,N_1840);
or U3649 (N_3649,N_695,N_8);
or U3650 (N_3650,N_1312,N_400);
or U3651 (N_3651,N_2133,N_2000);
and U3652 (N_3652,N_345,N_23);
nor U3653 (N_3653,N_1030,N_1873);
or U3654 (N_3654,N_1199,N_1089);
nand U3655 (N_3655,N_625,N_712);
and U3656 (N_3656,N_2234,N_1709);
nand U3657 (N_3657,N_1229,N_2341);
nor U3658 (N_3658,N_2473,N_1993);
nor U3659 (N_3659,N_1914,N_544);
or U3660 (N_3660,N_1868,N_0);
nor U3661 (N_3661,N_663,N_604);
nor U3662 (N_3662,N_641,N_1621);
or U3663 (N_3663,N_2387,N_1622);
or U3664 (N_3664,N_218,N_1323);
and U3665 (N_3665,N_1657,N_64);
nand U3666 (N_3666,N_718,N_2350);
nand U3667 (N_3667,N_108,N_820);
and U3668 (N_3668,N_1805,N_1949);
nand U3669 (N_3669,N_1074,N_243);
or U3670 (N_3670,N_1661,N_14);
or U3671 (N_3671,N_2082,N_2300);
or U3672 (N_3672,N_476,N_367);
and U3673 (N_3673,N_2487,N_1135);
and U3674 (N_3674,N_1059,N_1922);
or U3675 (N_3675,N_955,N_1793);
nand U3676 (N_3676,N_69,N_91);
nand U3677 (N_3677,N_228,N_2102);
nor U3678 (N_3678,N_1735,N_420);
and U3679 (N_3679,N_774,N_1023);
or U3680 (N_3680,N_118,N_1687);
nor U3681 (N_3681,N_563,N_2111);
nor U3682 (N_3682,N_31,N_1921);
nor U3683 (N_3683,N_1320,N_1180);
xor U3684 (N_3684,N_501,N_126);
or U3685 (N_3685,N_1219,N_2129);
nor U3686 (N_3686,N_1318,N_1976);
nand U3687 (N_3687,N_24,N_2158);
nand U3688 (N_3688,N_567,N_268);
nor U3689 (N_3689,N_1982,N_1438);
or U3690 (N_3690,N_1872,N_1040);
or U3691 (N_3691,N_414,N_772);
nor U3692 (N_3692,N_1704,N_706);
and U3693 (N_3693,N_2222,N_219);
or U3694 (N_3694,N_150,N_206);
nand U3695 (N_3695,N_2405,N_2025);
xnor U3696 (N_3696,N_1109,N_164);
nand U3697 (N_3697,N_379,N_2269);
and U3698 (N_3698,N_919,N_17);
nor U3699 (N_3699,N_1959,N_2332);
nor U3700 (N_3700,N_2385,N_667);
nor U3701 (N_3701,N_57,N_137);
nor U3702 (N_3702,N_1853,N_2345);
or U3703 (N_3703,N_806,N_672);
xnor U3704 (N_3704,N_178,N_2359);
or U3705 (N_3705,N_319,N_1619);
nand U3706 (N_3706,N_999,N_674);
and U3707 (N_3707,N_371,N_255);
or U3708 (N_3708,N_211,N_2293);
and U3709 (N_3709,N_1529,N_415);
nor U3710 (N_3710,N_1172,N_15);
or U3711 (N_3711,N_262,N_843);
or U3712 (N_3712,N_2248,N_1677);
nand U3713 (N_3713,N_2013,N_2256);
or U3714 (N_3714,N_1797,N_495);
nor U3715 (N_3715,N_779,N_2249);
and U3716 (N_3716,N_257,N_1457);
nor U3717 (N_3717,N_1046,N_1218);
nor U3718 (N_3718,N_338,N_2028);
and U3719 (N_3719,N_1044,N_2329);
or U3720 (N_3720,N_1451,N_1605);
and U3721 (N_3721,N_2245,N_710);
or U3722 (N_3722,N_2420,N_864);
and U3723 (N_3723,N_580,N_186);
and U3724 (N_3724,N_2438,N_251);
and U3725 (N_3725,N_2070,N_2195);
or U3726 (N_3726,N_716,N_155);
xnor U3727 (N_3727,N_2285,N_1481);
nor U3728 (N_3728,N_1084,N_342);
and U3729 (N_3729,N_1948,N_2253);
and U3730 (N_3730,N_181,N_698);
and U3731 (N_3731,N_693,N_1375);
nor U3732 (N_3732,N_1279,N_2074);
and U3733 (N_3733,N_2325,N_1006);
nand U3734 (N_3734,N_2349,N_398);
nand U3735 (N_3735,N_1743,N_1020);
nor U3736 (N_3736,N_1990,N_117);
nand U3737 (N_3737,N_2165,N_938);
nor U3738 (N_3738,N_527,N_2001);
or U3739 (N_3739,N_516,N_326);
and U3740 (N_3740,N_1270,N_380);
nand U3741 (N_3741,N_616,N_1316);
nand U3742 (N_3742,N_29,N_37);
or U3743 (N_3743,N_478,N_1308);
or U3744 (N_3744,N_1494,N_2244);
nand U3745 (N_3745,N_1898,N_608);
and U3746 (N_3746,N_671,N_662);
nor U3747 (N_3747,N_1851,N_1614);
nand U3748 (N_3748,N_564,N_2169);
and U3749 (N_3749,N_2047,N_2467);
nand U3750 (N_3750,N_2325,N_587);
and U3751 (N_3751,N_840,N_473);
or U3752 (N_3752,N_130,N_504);
nor U3753 (N_3753,N_1392,N_1230);
and U3754 (N_3754,N_1916,N_2363);
and U3755 (N_3755,N_1643,N_693);
and U3756 (N_3756,N_938,N_919);
or U3757 (N_3757,N_1844,N_1465);
and U3758 (N_3758,N_265,N_1789);
or U3759 (N_3759,N_2316,N_2039);
nand U3760 (N_3760,N_2178,N_1850);
or U3761 (N_3761,N_2483,N_1074);
or U3762 (N_3762,N_498,N_995);
or U3763 (N_3763,N_1405,N_240);
nand U3764 (N_3764,N_1858,N_763);
xor U3765 (N_3765,N_1699,N_610);
and U3766 (N_3766,N_2362,N_2460);
nor U3767 (N_3767,N_2345,N_2236);
nand U3768 (N_3768,N_153,N_110);
and U3769 (N_3769,N_2167,N_185);
nor U3770 (N_3770,N_1847,N_2470);
or U3771 (N_3771,N_1631,N_2390);
nand U3772 (N_3772,N_1907,N_25);
and U3773 (N_3773,N_1203,N_1813);
and U3774 (N_3774,N_836,N_2420);
xor U3775 (N_3775,N_2117,N_2077);
nor U3776 (N_3776,N_458,N_1219);
and U3777 (N_3777,N_1300,N_2129);
nor U3778 (N_3778,N_1046,N_2161);
nor U3779 (N_3779,N_1303,N_686);
or U3780 (N_3780,N_1025,N_141);
nor U3781 (N_3781,N_2370,N_1376);
and U3782 (N_3782,N_393,N_397);
and U3783 (N_3783,N_2094,N_1368);
or U3784 (N_3784,N_2195,N_84);
nand U3785 (N_3785,N_1095,N_766);
nor U3786 (N_3786,N_2060,N_2377);
nand U3787 (N_3787,N_295,N_778);
and U3788 (N_3788,N_969,N_13);
and U3789 (N_3789,N_1498,N_2018);
nand U3790 (N_3790,N_2445,N_425);
or U3791 (N_3791,N_823,N_2132);
nor U3792 (N_3792,N_2032,N_2081);
nand U3793 (N_3793,N_1153,N_436);
nand U3794 (N_3794,N_2034,N_1467);
or U3795 (N_3795,N_28,N_1313);
or U3796 (N_3796,N_1357,N_1680);
nor U3797 (N_3797,N_556,N_549);
and U3798 (N_3798,N_390,N_830);
and U3799 (N_3799,N_1495,N_682);
and U3800 (N_3800,N_337,N_668);
nand U3801 (N_3801,N_2062,N_2074);
and U3802 (N_3802,N_1971,N_214);
or U3803 (N_3803,N_991,N_1463);
or U3804 (N_3804,N_672,N_488);
nand U3805 (N_3805,N_2213,N_240);
nor U3806 (N_3806,N_1899,N_2425);
and U3807 (N_3807,N_1945,N_678);
nor U3808 (N_3808,N_639,N_1915);
and U3809 (N_3809,N_2286,N_2195);
or U3810 (N_3810,N_1302,N_966);
and U3811 (N_3811,N_1315,N_733);
nand U3812 (N_3812,N_570,N_966);
or U3813 (N_3813,N_670,N_1152);
and U3814 (N_3814,N_336,N_1869);
and U3815 (N_3815,N_57,N_1711);
nand U3816 (N_3816,N_1186,N_2364);
nor U3817 (N_3817,N_2156,N_1662);
and U3818 (N_3818,N_1234,N_694);
nor U3819 (N_3819,N_1606,N_770);
and U3820 (N_3820,N_2070,N_1583);
or U3821 (N_3821,N_257,N_1626);
nand U3822 (N_3822,N_1496,N_991);
nor U3823 (N_3823,N_2272,N_1410);
or U3824 (N_3824,N_790,N_2138);
nor U3825 (N_3825,N_436,N_1831);
and U3826 (N_3826,N_2239,N_781);
nor U3827 (N_3827,N_595,N_2257);
or U3828 (N_3828,N_1450,N_79);
nand U3829 (N_3829,N_449,N_994);
nand U3830 (N_3830,N_1364,N_556);
nor U3831 (N_3831,N_2499,N_1324);
nand U3832 (N_3832,N_1012,N_792);
and U3833 (N_3833,N_1212,N_1661);
xnor U3834 (N_3834,N_2164,N_1553);
nand U3835 (N_3835,N_2282,N_810);
or U3836 (N_3836,N_859,N_2075);
nor U3837 (N_3837,N_1437,N_95);
nor U3838 (N_3838,N_957,N_752);
nand U3839 (N_3839,N_1343,N_2175);
nand U3840 (N_3840,N_1410,N_43);
nor U3841 (N_3841,N_2415,N_2288);
nor U3842 (N_3842,N_1997,N_2162);
nand U3843 (N_3843,N_2394,N_2342);
or U3844 (N_3844,N_120,N_878);
or U3845 (N_3845,N_473,N_2092);
or U3846 (N_3846,N_902,N_2482);
or U3847 (N_3847,N_1378,N_2001);
and U3848 (N_3848,N_701,N_1169);
nor U3849 (N_3849,N_113,N_2201);
or U3850 (N_3850,N_1758,N_1521);
and U3851 (N_3851,N_2260,N_667);
or U3852 (N_3852,N_1117,N_2329);
nor U3853 (N_3853,N_927,N_647);
nand U3854 (N_3854,N_189,N_2470);
nand U3855 (N_3855,N_1612,N_1780);
or U3856 (N_3856,N_1657,N_577);
nand U3857 (N_3857,N_1553,N_961);
and U3858 (N_3858,N_678,N_729);
xnor U3859 (N_3859,N_850,N_336);
or U3860 (N_3860,N_1215,N_288);
or U3861 (N_3861,N_926,N_585);
and U3862 (N_3862,N_1474,N_1823);
and U3863 (N_3863,N_880,N_2096);
and U3864 (N_3864,N_1266,N_2067);
nor U3865 (N_3865,N_1460,N_115);
and U3866 (N_3866,N_888,N_2295);
and U3867 (N_3867,N_425,N_2358);
nand U3868 (N_3868,N_884,N_2052);
nand U3869 (N_3869,N_2260,N_584);
and U3870 (N_3870,N_2326,N_245);
nand U3871 (N_3871,N_1244,N_1939);
nand U3872 (N_3872,N_1358,N_1870);
nand U3873 (N_3873,N_1613,N_0);
nand U3874 (N_3874,N_2280,N_2484);
nor U3875 (N_3875,N_2360,N_332);
nand U3876 (N_3876,N_2067,N_269);
or U3877 (N_3877,N_1146,N_2174);
or U3878 (N_3878,N_920,N_1650);
or U3879 (N_3879,N_654,N_1543);
nor U3880 (N_3880,N_701,N_1355);
nor U3881 (N_3881,N_307,N_465);
and U3882 (N_3882,N_1894,N_1841);
nor U3883 (N_3883,N_661,N_446);
or U3884 (N_3884,N_1855,N_1885);
nor U3885 (N_3885,N_1964,N_2302);
nand U3886 (N_3886,N_2277,N_308);
and U3887 (N_3887,N_2310,N_526);
or U3888 (N_3888,N_471,N_124);
nand U3889 (N_3889,N_726,N_1521);
or U3890 (N_3890,N_1159,N_1900);
or U3891 (N_3891,N_2215,N_1900);
nor U3892 (N_3892,N_2185,N_1000);
nand U3893 (N_3893,N_2424,N_1189);
and U3894 (N_3894,N_443,N_1611);
nand U3895 (N_3895,N_500,N_1359);
or U3896 (N_3896,N_1027,N_1247);
or U3897 (N_3897,N_1557,N_20);
nor U3898 (N_3898,N_1663,N_2271);
or U3899 (N_3899,N_1691,N_1231);
and U3900 (N_3900,N_876,N_666);
nor U3901 (N_3901,N_683,N_1589);
or U3902 (N_3902,N_281,N_1066);
or U3903 (N_3903,N_711,N_803);
nand U3904 (N_3904,N_612,N_2349);
and U3905 (N_3905,N_1303,N_1117);
or U3906 (N_3906,N_1715,N_1802);
nand U3907 (N_3907,N_479,N_1229);
nand U3908 (N_3908,N_2113,N_2367);
nand U3909 (N_3909,N_896,N_1963);
and U3910 (N_3910,N_781,N_420);
nor U3911 (N_3911,N_807,N_2018);
or U3912 (N_3912,N_567,N_1772);
or U3913 (N_3913,N_381,N_2419);
nand U3914 (N_3914,N_1422,N_948);
nand U3915 (N_3915,N_1161,N_1991);
nor U3916 (N_3916,N_1339,N_1469);
nor U3917 (N_3917,N_2359,N_2444);
and U3918 (N_3918,N_1709,N_651);
nor U3919 (N_3919,N_408,N_1344);
and U3920 (N_3920,N_127,N_1656);
or U3921 (N_3921,N_934,N_506);
or U3922 (N_3922,N_955,N_2372);
and U3923 (N_3923,N_1426,N_942);
and U3924 (N_3924,N_1557,N_600);
and U3925 (N_3925,N_1544,N_1596);
and U3926 (N_3926,N_1797,N_1299);
or U3927 (N_3927,N_1961,N_2431);
nand U3928 (N_3928,N_1820,N_1582);
and U3929 (N_3929,N_688,N_2374);
or U3930 (N_3930,N_1934,N_1029);
nor U3931 (N_3931,N_405,N_1292);
nand U3932 (N_3932,N_2475,N_1408);
nor U3933 (N_3933,N_2478,N_916);
nand U3934 (N_3934,N_1166,N_1427);
nand U3935 (N_3935,N_1379,N_516);
nor U3936 (N_3936,N_1606,N_1301);
nand U3937 (N_3937,N_2379,N_943);
or U3938 (N_3938,N_467,N_656);
or U3939 (N_3939,N_196,N_976);
nor U3940 (N_3940,N_2028,N_13);
or U3941 (N_3941,N_2481,N_24);
or U3942 (N_3942,N_409,N_2346);
and U3943 (N_3943,N_369,N_236);
nor U3944 (N_3944,N_1058,N_1912);
nor U3945 (N_3945,N_2178,N_855);
nor U3946 (N_3946,N_1538,N_1272);
or U3947 (N_3947,N_1760,N_65);
nor U3948 (N_3948,N_882,N_778);
and U3949 (N_3949,N_2331,N_783);
and U3950 (N_3950,N_287,N_2290);
nor U3951 (N_3951,N_1545,N_894);
nor U3952 (N_3952,N_349,N_1809);
and U3953 (N_3953,N_1630,N_1572);
or U3954 (N_3954,N_2445,N_1949);
or U3955 (N_3955,N_257,N_1824);
or U3956 (N_3956,N_585,N_1214);
and U3957 (N_3957,N_2444,N_2259);
or U3958 (N_3958,N_564,N_2239);
nor U3959 (N_3959,N_234,N_956);
nand U3960 (N_3960,N_1116,N_1450);
or U3961 (N_3961,N_9,N_1794);
nand U3962 (N_3962,N_514,N_962);
nor U3963 (N_3963,N_2274,N_430);
nand U3964 (N_3964,N_2458,N_2033);
nand U3965 (N_3965,N_1375,N_1563);
nand U3966 (N_3966,N_2221,N_1630);
or U3967 (N_3967,N_345,N_1516);
and U3968 (N_3968,N_2231,N_923);
nand U3969 (N_3969,N_728,N_832);
nor U3970 (N_3970,N_1108,N_1188);
and U3971 (N_3971,N_1775,N_176);
or U3972 (N_3972,N_1521,N_1930);
xor U3973 (N_3973,N_1745,N_1037);
or U3974 (N_3974,N_1626,N_1966);
or U3975 (N_3975,N_2145,N_638);
or U3976 (N_3976,N_2325,N_1130);
nand U3977 (N_3977,N_1104,N_2369);
or U3978 (N_3978,N_643,N_1736);
nand U3979 (N_3979,N_1638,N_1081);
and U3980 (N_3980,N_2333,N_1674);
nor U3981 (N_3981,N_1799,N_2148);
nor U3982 (N_3982,N_1228,N_77);
or U3983 (N_3983,N_456,N_1751);
and U3984 (N_3984,N_421,N_2461);
or U3985 (N_3985,N_1121,N_2430);
nor U3986 (N_3986,N_1431,N_272);
or U3987 (N_3987,N_498,N_1653);
nor U3988 (N_3988,N_1677,N_1168);
nand U3989 (N_3989,N_1039,N_450);
and U3990 (N_3990,N_2001,N_1899);
and U3991 (N_3991,N_933,N_1047);
nand U3992 (N_3992,N_1911,N_1768);
nand U3993 (N_3993,N_2427,N_955);
nor U3994 (N_3994,N_196,N_284);
nor U3995 (N_3995,N_2348,N_1158);
or U3996 (N_3996,N_1153,N_932);
nor U3997 (N_3997,N_727,N_99);
and U3998 (N_3998,N_271,N_566);
nand U3999 (N_3999,N_740,N_1777);
and U4000 (N_4000,N_635,N_1826);
or U4001 (N_4001,N_1150,N_108);
xor U4002 (N_4002,N_264,N_1045);
and U4003 (N_4003,N_1378,N_1867);
and U4004 (N_4004,N_504,N_149);
or U4005 (N_4005,N_1647,N_113);
or U4006 (N_4006,N_292,N_1123);
nand U4007 (N_4007,N_880,N_1246);
nand U4008 (N_4008,N_2130,N_147);
nor U4009 (N_4009,N_595,N_510);
nand U4010 (N_4010,N_1505,N_1332);
or U4011 (N_4011,N_1603,N_142);
nand U4012 (N_4012,N_359,N_2466);
and U4013 (N_4013,N_1524,N_2391);
and U4014 (N_4014,N_436,N_1461);
nand U4015 (N_4015,N_1253,N_803);
and U4016 (N_4016,N_1601,N_228);
nand U4017 (N_4017,N_610,N_857);
nand U4018 (N_4018,N_537,N_2127);
and U4019 (N_4019,N_1533,N_1129);
and U4020 (N_4020,N_1638,N_1628);
and U4021 (N_4021,N_1059,N_1084);
or U4022 (N_4022,N_1768,N_1353);
nor U4023 (N_4023,N_1881,N_285);
nand U4024 (N_4024,N_2185,N_1831);
nor U4025 (N_4025,N_1652,N_2359);
nor U4026 (N_4026,N_2181,N_1025);
nor U4027 (N_4027,N_1659,N_394);
nor U4028 (N_4028,N_2350,N_877);
or U4029 (N_4029,N_592,N_528);
or U4030 (N_4030,N_269,N_1193);
or U4031 (N_4031,N_696,N_285);
and U4032 (N_4032,N_1818,N_531);
or U4033 (N_4033,N_493,N_2002);
or U4034 (N_4034,N_728,N_2443);
and U4035 (N_4035,N_2452,N_1703);
and U4036 (N_4036,N_2275,N_504);
nand U4037 (N_4037,N_2311,N_1833);
or U4038 (N_4038,N_1330,N_2266);
nor U4039 (N_4039,N_1159,N_1417);
and U4040 (N_4040,N_2204,N_1581);
and U4041 (N_4041,N_2365,N_1195);
or U4042 (N_4042,N_1831,N_1744);
nor U4043 (N_4043,N_1394,N_1388);
nand U4044 (N_4044,N_1717,N_1109);
nand U4045 (N_4045,N_1183,N_1663);
or U4046 (N_4046,N_1240,N_934);
nor U4047 (N_4047,N_814,N_1051);
or U4048 (N_4048,N_368,N_287);
nor U4049 (N_4049,N_319,N_604);
or U4050 (N_4050,N_2375,N_2018);
or U4051 (N_4051,N_1814,N_1273);
or U4052 (N_4052,N_418,N_1979);
nand U4053 (N_4053,N_83,N_1525);
or U4054 (N_4054,N_1049,N_2015);
nor U4055 (N_4055,N_2386,N_1046);
or U4056 (N_4056,N_1437,N_2275);
nand U4057 (N_4057,N_1902,N_49);
xor U4058 (N_4058,N_531,N_520);
or U4059 (N_4059,N_1557,N_1561);
nor U4060 (N_4060,N_2456,N_1559);
xnor U4061 (N_4061,N_1927,N_2296);
nand U4062 (N_4062,N_2092,N_1792);
nor U4063 (N_4063,N_1613,N_1098);
or U4064 (N_4064,N_580,N_2498);
or U4065 (N_4065,N_2387,N_2150);
nand U4066 (N_4066,N_2208,N_1956);
and U4067 (N_4067,N_219,N_1090);
nand U4068 (N_4068,N_2239,N_1700);
nor U4069 (N_4069,N_1125,N_1235);
nor U4070 (N_4070,N_1957,N_999);
or U4071 (N_4071,N_1075,N_1115);
or U4072 (N_4072,N_2090,N_710);
nand U4073 (N_4073,N_2419,N_2339);
nand U4074 (N_4074,N_1512,N_945);
nor U4075 (N_4075,N_2146,N_1064);
or U4076 (N_4076,N_2430,N_2051);
or U4077 (N_4077,N_626,N_398);
and U4078 (N_4078,N_612,N_753);
or U4079 (N_4079,N_1896,N_628);
or U4080 (N_4080,N_819,N_1255);
or U4081 (N_4081,N_411,N_2158);
and U4082 (N_4082,N_279,N_325);
nor U4083 (N_4083,N_913,N_712);
or U4084 (N_4084,N_1627,N_728);
nor U4085 (N_4085,N_2008,N_431);
or U4086 (N_4086,N_502,N_1917);
or U4087 (N_4087,N_452,N_2432);
and U4088 (N_4088,N_640,N_852);
nor U4089 (N_4089,N_1431,N_2306);
nand U4090 (N_4090,N_241,N_1771);
nor U4091 (N_4091,N_382,N_709);
nor U4092 (N_4092,N_879,N_2001);
nand U4093 (N_4093,N_1969,N_738);
nand U4094 (N_4094,N_900,N_2098);
nor U4095 (N_4095,N_1268,N_60);
and U4096 (N_4096,N_112,N_1900);
nand U4097 (N_4097,N_532,N_870);
or U4098 (N_4098,N_2268,N_863);
nand U4099 (N_4099,N_1107,N_2037);
or U4100 (N_4100,N_729,N_1194);
nor U4101 (N_4101,N_528,N_1489);
or U4102 (N_4102,N_405,N_1377);
and U4103 (N_4103,N_662,N_1068);
or U4104 (N_4104,N_2159,N_1835);
or U4105 (N_4105,N_1478,N_893);
or U4106 (N_4106,N_2249,N_1000);
nor U4107 (N_4107,N_2407,N_1126);
and U4108 (N_4108,N_713,N_1171);
nor U4109 (N_4109,N_2490,N_1560);
and U4110 (N_4110,N_1886,N_1837);
nand U4111 (N_4111,N_659,N_394);
and U4112 (N_4112,N_1140,N_1905);
nand U4113 (N_4113,N_451,N_949);
or U4114 (N_4114,N_1023,N_85);
nand U4115 (N_4115,N_1642,N_2273);
nand U4116 (N_4116,N_802,N_2425);
nor U4117 (N_4117,N_369,N_1987);
and U4118 (N_4118,N_1443,N_1685);
nor U4119 (N_4119,N_857,N_1431);
or U4120 (N_4120,N_2031,N_2432);
and U4121 (N_4121,N_1882,N_1417);
and U4122 (N_4122,N_1603,N_706);
and U4123 (N_4123,N_1319,N_791);
nor U4124 (N_4124,N_822,N_2165);
nand U4125 (N_4125,N_842,N_239);
and U4126 (N_4126,N_152,N_2133);
nor U4127 (N_4127,N_2133,N_2162);
or U4128 (N_4128,N_1478,N_295);
nor U4129 (N_4129,N_793,N_2138);
nand U4130 (N_4130,N_1973,N_1803);
nand U4131 (N_4131,N_519,N_1985);
nor U4132 (N_4132,N_1563,N_201);
and U4133 (N_4133,N_426,N_505);
nand U4134 (N_4134,N_1656,N_1688);
nand U4135 (N_4135,N_858,N_69);
or U4136 (N_4136,N_363,N_834);
nand U4137 (N_4137,N_189,N_2275);
and U4138 (N_4138,N_1806,N_595);
xor U4139 (N_4139,N_1028,N_2431);
nand U4140 (N_4140,N_843,N_77);
or U4141 (N_4141,N_2065,N_950);
nand U4142 (N_4142,N_1320,N_1398);
nor U4143 (N_4143,N_1580,N_2203);
or U4144 (N_4144,N_2435,N_1386);
or U4145 (N_4145,N_177,N_1203);
nor U4146 (N_4146,N_434,N_225);
and U4147 (N_4147,N_895,N_110);
nor U4148 (N_4148,N_1290,N_2481);
nor U4149 (N_4149,N_1680,N_1653);
nand U4150 (N_4150,N_499,N_677);
nand U4151 (N_4151,N_2073,N_824);
nand U4152 (N_4152,N_1108,N_2185);
nor U4153 (N_4153,N_1254,N_2246);
or U4154 (N_4154,N_1833,N_92);
or U4155 (N_4155,N_1245,N_394);
nor U4156 (N_4156,N_2086,N_103);
nor U4157 (N_4157,N_2147,N_1654);
nand U4158 (N_4158,N_55,N_1828);
and U4159 (N_4159,N_498,N_1105);
nor U4160 (N_4160,N_1796,N_1442);
nor U4161 (N_4161,N_2048,N_2454);
or U4162 (N_4162,N_1842,N_964);
or U4163 (N_4163,N_2497,N_943);
or U4164 (N_4164,N_321,N_347);
nand U4165 (N_4165,N_2143,N_172);
or U4166 (N_4166,N_2083,N_177);
nand U4167 (N_4167,N_308,N_2269);
nand U4168 (N_4168,N_1436,N_1184);
nand U4169 (N_4169,N_17,N_801);
nand U4170 (N_4170,N_2159,N_691);
and U4171 (N_4171,N_2280,N_898);
nor U4172 (N_4172,N_998,N_972);
or U4173 (N_4173,N_2301,N_1084);
or U4174 (N_4174,N_1973,N_1385);
and U4175 (N_4175,N_1437,N_784);
or U4176 (N_4176,N_437,N_1368);
nand U4177 (N_4177,N_1817,N_826);
and U4178 (N_4178,N_76,N_1113);
nor U4179 (N_4179,N_47,N_1750);
nor U4180 (N_4180,N_320,N_2301);
or U4181 (N_4181,N_1252,N_1890);
and U4182 (N_4182,N_329,N_1776);
nor U4183 (N_4183,N_1169,N_704);
and U4184 (N_4184,N_1808,N_1350);
nand U4185 (N_4185,N_2328,N_858);
or U4186 (N_4186,N_282,N_1311);
or U4187 (N_4187,N_2193,N_2270);
or U4188 (N_4188,N_2436,N_556);
or U4189 (N_4189,N_2318,N_146);
and U4190 (N_4190,N_227,N_2456);
or U4191 (N_4191,N_249,N_1028);
nand U4192 (N_4192,N_979,N_1182);
or U4193 (N_4193,N_2140,N_101);
and U4194 (N_4194,N_1108,N_2464);
nand U4195 (N_4195,N_2453,N_33);
nor U4196 (N_4196,N_1981,N_2019);
nor U4197 (N_4197,N_1346,N_1219);
or U4198 (N_4198,N_756,N_1848);
nor U4199 (N_4199,N_1842,N_94);
nor U4200 (N_4200,N_1543,N_19);
nor U4201 (N_4201,N_2378,N_434);
and U4202 (N_4202,N_2005,N_196);
nor U4203 (N_4203,N_1030,N_2004);
or U4204 (N_4204,N_1997,N_1639);
nor U4205 (N_4205,N_1450,N_637);
nand U4206 (N_4206,N_1691,N_942);
nand U4207 (N_4207,N_2360,N_1394);
or U4208 (N_4208,N_1527,N_165);
xnor U4209 (N_4209,N_342,N_2217);
nor U4210 (N_4210,N_1656,N_52);
and U4211 (N_4211,N_84,N_1808);
and U4212 (N_4212,N_1053,N_2262);
and U4213 (N_4213,N_571,N_1195);
or U4214 (N_4214,N_1124,N_482);
or U4215 (N_4215,N_790,N_177);
and U4216 (N_4216,N_935,N_1414);
nor U4217 (N_4217,N_1275,N_40);
nor U4218 (N_4218,N_1376,N_2445);
or U4219 (N_4219,N_1585,N_358);
and U4220 (N_4220,N_362,N_1957);
nand U4221 (N_4221,N_1103,N_1547);
and U4222 (N_4222,N_2267,N_2127);
and U4223 (N_4223,N_1981,N_2011);
or U4224 (N_4224,N_419,N_2259);
or U4225 (N_4225,N_2242,N_1814);
nand U4226 (N_4226,N_757,N_2475);
nor U4227 (N_4227,N_1830,N_1080);
nor U4228 (N_4228,N_701,N_731);
or U4229 (N_4229,N_1868,N_219);
and U4230 (N_4230,N_1891,N_1040);
nand U4231 (N_4231,N_1384,N_448);
nand U4232 (N_4232,N_2371,N_909);
nand U4233 (N_4233,N_2451,N_2420);
or U4234 (N_4234,N_140,N_1828);
and U4235 (N_4235,N_829,N_2411);
and U4236 (N_4236,N_2249,N_309);
nor U4237 (N_4237,N_899,N_2403);
xor U4238 (N_4238,N_2474,N_252);
nor U4239 (N_4239,N_2282,N_1106);
and U4240 (N_4240,N_1527,N_838);
nand U4241 (N_4241,N_590,N_686);
nor U4242 (N_4242,N_1473,N_2441);
xor U4243 (N_4243,N_201,N_1798);
nand U4244 (N_4244,N_1210,N_573);
nand U4245 (N_4245,N_118,N_2291);
or U4246 (N_4246,N_82,N_1683);
or U4247 (N_4247,N_2173,N_429);
or U4248 (N_4248,N_869,N_902);
or U4249 (N_4249,N_1573,N_1443);
nor U4250 (N_4250,N_1756,N_1784);
nand U4251 (N_4251,N_2167,N_1085);
and U4252 (N_4252,N_1585,N_2067);
nor U4253 (N_4253,N_2330,N_2100);
nand U4254 (N_4254,N_2395,N_1220);
nor U4255 (N_4255,N_145,N_878);
or U4256 (N_4256,N_2415,N_211);
or U4257 (N_4257,N_2342,N_1747);
nor U4258 (N_4258,N_2045,N_1478);
or U4259 (N_4259,N_189,N_1559);
nor U4260 (N_4260,N_1551,N_459);
nand U4261 (N_4261,N_1964,N_1038);
and U4262 (N_4262,N_1232,N_1680);
and U4263 (N_4263,N_2475,N_1113);
or U4264 (N_4264,N_2086,N_1782);
nand U4265 (N_4265,N_1863,N_1426);
nor U4266 (N_4266,N_559,N_2080);
nand U4267 (N_4267,N_179,N_1952);
nand U4268 (N_4268,N_71,N_2240);
and U4269 (N_4269,N_789,N_1688);
nor U4270 (N_4270,N_2059,N_908);
and U4271 (N_4271,N_2215,N_1091);
nor U4272 (N_4272,N_1294,N_1490);
or U4273 (N_4273,N_1293,N_682);
nor U4274 (N_4274,N_1947,N_1284);
nand U4275 (N_4275,N_465,N_1249);
nor U4276 (N_4276,N_1979,N_1331);
nand U4277 (N_4277,N_1026,N_1335);
or U4278 (N_4278,N_911,N_566);
nand U4279 (N_4279,N_317,N_1312);
and U4280 (N_4280,N_763,N_505);
nor U4281 (N_4281,N_1489,N_1589);
or U4282 (N_4282,N_1342,N_1811);
nand U4283 (N_4283,N_150,N_1424);
or U4284 (N_4284,N_1612,N_1896);
xor U4285 (N_4285,N_851,N_2370);
nand U4286 (N_4286,N_1051,N_226);
nand U4287 (N_4287,N_1546,N_567);
or U4288 (N_4288,N_2141,N_72);
or U4289 (N_4289,N_2370,N_344);
and U4290 (N_4290,N_1433,N_437);
nor U4291 (N_4291,N_967,N_1551);
nand U4292 (N_4292,N_2084,N_1638);
or U4293 (N_4293,N_49,N_1605);
or U4294 (N_4294,N_263,N_2105);
nor U4295 (N_4295,N_553,N_767);
nand U4296 (N_4296,N_121,N_2187);
and U4297 (N_4297,N_373,N_901);
or U4298 (N_4298,N_1453,N_874);
and U4299 (N_4299,N_240,N_14);
nor U4300 (N_4300,N_1046,N_343);
and U4301 (N_4301,N_1118,N_913);
xnor U4302 (N_4302,N_26,N_298);
nand U4303 (N_4303,N_102,N_1682);
nor U4304 (N_4304,N_2477,N_2478);
or U4305 (N_4305,N_1457,N_214);
nand U4306 (N_4306,N_855,N_2040);
or U4307 (N_4307,N_1090,N_1927);
or U4308 (N_4308,N_1571,N_2191);
and U4309 (N_4309,N_1473,N_1885);
or U4310 (N_4310,N_2226,N_1470);
nand U4311 (N_4311,N_1969,N_453);
nor U4312 (N_4312,N_2090,N_47);
nor U4313 (N_4313,N_447,N_281);
and U4314 (N_4314,N_267,N_655);
nor U4315 (N_4315,N_292,N_605);
or U4316 (N_4316,N_2217,N_1858);
nand U4317 (N_4317,N_1760,N_683);
and U4318 (N_4318,N_1791,N_619);
nand U4319 (N_4319,N_2115,N_642);
and U4320 (N_4320,N_2287,N_1697);
nor U4321 (N_4321,N_1839,N_2276);
nand U4322 (N_4322,N_1929,N_841);
nand U4323 (N_4323,N_1649,N_2201);
nor U4324 (N_4324,N_651,N_1348);
or U4325 (N_4325,N_1710,N_1932);
nand U4326 (N_4326,N_518,N_1907);
or U4327 (N_4327,N_2367,N_2268);
xnor U4328 (N_4328,N_1320,N_687);
or U4329 (N_4329,N_2384,N_834);
and U4330 (N_4330,N_1981,N_790);
and U4331 (N_4331,N_467,N_734);
or U4332 (N_4332,N_1543,N_2360);
and U4333 (N_4333,N_1491,N_179);
nand U4334 (N_4334,N_18,N_1551);
or U4335 (N_4335,N_1916,N_1375);
nor U4336 (N_4336,N_1546,N_1488);
and U4337 (N_4337,N_154,N_355);
nor U4338 (N_4338,N_313,N_382);
or U4339 (N_4339,N_2436,N_68);
or U4340 (N_4340,N_2006,N_365);
and U4341 (N_4341,N_2376,N_1311);
and U4342 (N_4342,N_1040,N_1324);
nor U4343 (N_4343,N_738,N_1470);
or U4344 (N_4344,N_185,N_2372);
nand U4345 (N_4345,N_1995,N_358);
nor U4346 (N_4346,N_2413,N_1105);
or U4347 (N_4347,N_1071,N_2219);
and U4348 (N_4348,N_2275,N_1266);
or U4349 (N_4349,N_617,N_560);
xor U4350 (N_4350,N_1337,N_787);
nand U4351 (N_4351,N_1948,N_856);
nor U4352 (N_4352,N_924,N_1137);
or U4353 (N_4353,N_1356,N_24);
nor U4354 (N_4354,N_1268,N_2287);
and U4355 (N_4355,N_469,N_326);
nand U4356 (N_4356,N_2402,N_253);
nor U4357 (N_4357,N_151,N_954);
or U4358 (N_4358,N_2413,N_1605);
nand U4359 (N_4359,N_961,N_1119);
or U4360 (N_4360,N_2229,N_1952);
and U4361 (N_4361,N_560,N_1555);
nor U4362 (N_4362,N_580,N_334);
nor U4363 (N_4363,N_1325,N_2002);
or U4364 (N_4364,N_1752,N_336);
nand U4365 (N_4365,N_1635,N_1520);
nor U4366 (N_4366,N_2462,N_1261);
and U4367 (N_4367,N_767,N_2411);
and U4368 (N_4368,N_1574,N_2229);
or U4369 (N_4369,N_1812,N_304);
and U4370 (N_4370,N_750,N_241);
nor U4371 (N_4371,N_2044,N_86);
nand U4372 (N_4372,N_1382,N_236);
nand U4373 (N_4373,N_1825,N_1622);
nand U4374 (N_4374,N_187,N_935);
nor U4375 (N_4375,N_1542,N_1248);
or U4376 (N_4376,N_1139,N_1590);
or U4377 (N_4377,N_853,N_1358);
and U4378 (N_4378,N_727,N_1568);
nor U4379 (N_4379,N_864,N_1167);
nor U4380 (N_4380,N_1436,N_1886);
or U4381 (N_4381,N_1090,N_1955);
nand U4382 (N_4382,N_699,N_1309);
nand U4383 (N_4383,N_37,N_1923);
nor U4384 (N_4384,N_586,N_2350);
and U4385 (N_4385,N_384,N_2036);
and U4386 (N_4386,N_1537,N_1482);
nand U4387 (N_4387,N_2176,N_247);
or U4388 (N_4388,N_492,N_974);
and U4389 (N_4389,N_1425,N_2143);
nor U4390 (N_4390,N_1365,N_1149);
or U4391 (N_4391,N_701,N_456);
and U4392 (N_4392,N_1540,N_1896);
or U4393 (N_4393,N_136,N_1578);
nand U4394 (N_4394,N_1433,N_804);
or U4395 (N_4395,N_2231,N_365);
or U4396 (N_4396,N_782,N_1577);
nor U4397 (N_4397,N_1827,N_670);
nand U4398 (N_4398,N_1516,N_252);
and U4399 (N_4399,N_633,N_1946);
nand U4400 (N_4400,N_2420,N_744);
nor U4401 (N_4401,N_1585,N_2244);
nand U4402 (N_4402,N_1456,N_644);
nand U4403 (N_4403,N_2311,N_785);
and U4404 (N_4404,N_2304,N_390);
nor U4405 (N_4405,N_1798,N_886);
nand U4406 (N_4406,N_1987,N_1989);
nand U4407 (N_4407,N_37,N_1643);
xor U4408 (N_4408,N_473,N_1397);
or U4409 (N_4409,N_2116,N_1467);
nor U4410 (N_4410,N_1847,N_1388);
or U4411 (N_4411,N_252,N_2247);
nor U4412 (N_4412,N_2363,N_2345);
nor U4413 (N_4413,N_304,N_1601);
nor U4414 (N_4414,N_633,N_1663);
and U4415 (N_4415,N_647,N_1504);
nand U4416 (N_4416,N_125,N_2397);
and U4417 (N_4417,N_1914,N_1327);
or U4418 (N_4418,N_1501,N_2176);
or U4419 (N_4419,N_202,N_353);
and U4420 (N_4420,N_1687,N_1389);
nand U4421 (N_4421,N_103,N_2399);
nor U4422 (N_4422,N_2056,N_2434);
and U4423 (N_4423,N_768,N_983);
or U4424 (N_4424,N_491,N_474);
nand U4425 (N_4425,N_1591,N_1636);
or U4426 (N_4426,N_2069,N_1839);
nor U4427 (N_4427,N_1731,N_2495);
nand U4428 (N_4428,N_804,N_1597);
nor U4429 (N_4429,N_16,N_92);
nor U4430 (N_4430,N_2317,N_1046);
nor U4431 (N_4431,N_1414,N_582);
nand U4432 (N_4432,N_1185,N_1952);
or U4433 (N_4433,N_717,N_801);
nor U4434 (N_4434,N_474,N_2242);
nor U4435 (N_4435,N_1994,N_2066);
or U4436 (N_4436,N_2310,N_409);
or U4437 (N_4437,N_2114,N_286);
or U4438 (N_4438,N_1085,N_845);
nor U4439 (N_4439,N_2086,N_841);
nand U4440 (N_4440,N_2409,N_2006);
nor U4441 (N_4441,N_1869,N_2312);
nand U4442 (N_4442,N_894,N_1745);
and U4443 (N_4443,N_1462,N_580);
and U4444 (N_4444,N_1676,N_1628);
nor U4445 (N_4445,N_1806,N_1971);
or U4446 (N_4446,N_336,N_205);
and U4447 (N_4447,N_1253,N_889);
nor U4448 (N_4448,N_310,N_2106);
nand U4449 (N_4449,N_97,N_1966);
nand U4450 (N_4450,N_1541,N_2335);
xor U4451 (N_4451,N_1494,N_1079);
nand U4452 (N_4452,N_1050,N_1502);
nor U4453 (N_4453,N_1323,N_961);
and U4454 (N_4454,N_1487,N_1410);
nor U4455 (N_4455,N_2362,N_440);
and U4456 (N_4456,N_879,N_2177);
and U4457 (N_4457,N_1784,N_2040);
nor U4458 (N_4458,N_172,N_1017);
and U4459 (N_4459,N_1384,N_908);
or U4460 (N_4460,N_906,N_57);
and U4461 (N_4461,N_214,N_839);
nand U4462 (N_4462,N_646,N_444);
nor U4463 (N_4463,N_271,N_1640);
and U4464 (N_4464,N_35,N_309);
and U4465 (N_4465,N_1684,N_845);
xor U4466 (N_4466,N_947,N_39);
nor U4467 (N_4467,N_217,N_951);
nor U4468 (N_4468,N_2308,N_1251);
nor U4469 (N_4469,N_2186,N_1663);
nand U4470 (N_4470,N_1331,N_1632);
xnor U4471 (N_4471,N_1388,N_2400);
nor U4472 (N_4472,N_1306,N_973);
or U4473 (N_4473,N_1361,N_2249);
nor U4474 (N_4474,N_1075,N_2238);
and U4475 (N_4475,N_1294,N_354);
or U4476 (N_4476,N_346,N_1488);
and U4477 (N_4477,N_817,N_2280);
nand U4478 (N_4478,N_726,N_1740);
or U4479 (N_4479,N_1173,N_2151);
nor U4480 (N_4480,N_123,N_760);
and U4481 (N_4481,N_290,N_2496);
xnor U4482 (N_4482,N_418,N_852);
nor U4483 (N_4483,N_1528,N_201);
nor U4484 (N_4484,N_2172,N_872);
nand U4485 (N_4485,N_1092,N_1589);
nor U4486 (N_4486,N_882,N_2322);
xor U4487 (N_4487,N_1084,N_1446);
nand U4488 (N_4488,N_74,N_2018);
nor U4489 (N_4489,N_232,N_920);
nand U4490 (N_4490,N_942,N_2070);
or U4491 (N_4491,N_1877,N_882);
nand U4492 (N_4492,N_750,N_2185);
nor U4493 (N_4493,N_772,N_2467);
nor U4494 (N_4494,N_750,N_402);
nor U4495 (N_4495,N_2318,N_2489);
or U4496 (N_4496,N_1591,N_557);
nor U4497 (N_4497,N_594,N_146);
and U4498 (N_4498,N_975,N_1360);
nand U4499 (N_4499,N_2114,N_253);
or U4500 (N_4500,N_117,N_1835);
or U4501 (N_4501,N_917,N_1285);
or U4502 (N_4502,N_2450,N_1071);
nand U4503 (N_4503,N_1503,N_660);
and U4504 (N_4504,N_2047,N_270);
nor U4505 (N_4505,N_1405,N_271);
and U4506 (N_4506,N_206,N_271);
or U4507 (N_4507,N_906,N_1512);
or U4508 (N_4508,N_1500,N_576);
nand U4509 (N_4509,N_2329,N_1485);
or U4510 (N_4510,N_754,N_1617);
nand U4511 (N_4511,N_545,N_1852);
nand U4512 (N_4512,N_863,N_2399);
or U4513 (N_4513,N_528,N_958);
or U4514 (N_4514,N_36,N_2011);
nand U4515 (N_4515,N_1121,N_1600);
and U4516 (N_4516,N_941,N_182);
or U4517 (N_4517,N_244,N_1347);
nor U4518 (N_4518,N_2266,N_397);
nand U4519 (N_4519,N_2174,N_2202);
and U4520 (N_4520,N_1761,N_1823);
nor U4521 (N_4521,N_1116,N_1648);
or U4522 (N_4522,N_223,N_521);
nand U4523 (N_4523,N_1134,N_808);
and U4524 (N_4524,N_694,N_864);
nor U4525 (N_4525,N_1327,N_1504);
nor U4526 (N_4526,N_1782,N_2483);
nand U4527 (N_4527,N_598,N_2142);
and U4528 (N_4528,N_1443,N_1739);
nand U4529 (N_4529,N_732,N_2464);
or U4530 (N_4530,N_2392,N_2042);
nor U4531 (N_4531,N_2429,N_873);
and U4532 (N_4532,N_1454,N_719);
nand U4533 (N_4533,N_2136,N_787);
nand U4534 (N_4534,N_1625,N_1533);
nand U4535 (N_4535,N_1985,N_1577);
and U4536 (N_4536,N_197,N_1698);
and U4537 (N_4537,N_1835,N_1007);
and U4538 (N_4538,N_673,N_2024);
or U4539 (N_4539,N_42,N_464);
nand U4540 (N_4540,N_2129,N_1666);
or U4541 (N_4541,N_1615,N_2129);
nand U4542 (N_4542,N_1796,N_1265);
or U4543 (N_4543,N_2326,N_426);
or U4544 (N_4544,N_2296,N_316);
nor U4545 (N_4545,N_2421,N_919);
nor U4546 (N_4546,N_987,N_1054);
nand U4547 (N_4547,N_2274,N_1229);
nand U4548 (N_4548,N_1653,N_1758);
nand U4549 (N_4549,N_723,N_22);
nor U4550 (N_4550,N_542,N_922);
nand U4551 (N_4551,N_57,N_2465);
or U4552 (N_4552,N_1200,N_1098);
nand U4553 (N_4553,N_1158,N_2009);
or U4554 (N_4554,N_1756,N_474);
and U4555 (N_4555,N_1695,N_14);
xnor U4556 (N_4556,N_1580,N_1827);
nand U4557 (N_4557,N_2244,N_1390);
and U4558 (N_4558,N_958,N_1256);
or U4559 (N_4559,N_1416,N_2005);
or U4560 (N_4560,N_274,N_801);
and U4561 (N_4561,N_23,N_963);
nand U4562 (N_4562,N_2374,N_302);
and U4563 (N_4563,N_385,N_1729);
and U4564 (N_4564,N_305,N_2133);
xor U4565 (N_4565,N_1499,N_384);
or U4566 (N_4566,N_1168,N_2060);
or U4567 (N_4567,N_397,N_1822);
nand U4568 (N_4568,N_1101,N_218);
nor U4569 (N_4569,N_146,N_69);
nand U4570 (N_4570,N_897,N_294);
nor U4571 (N_4571,N_2191,N_148);
nand U4572 (N_4572,N_793,N_803);
or U4573 (N_4573,N_207,N_1751);
nor U4574 (N_4574,N_2083,N_538);
nor U4575 (N_4575,N_1064,N_380);
nor U4576 (N_4576,N_849,N_915);
and U4577 (N_4577,N_1354,N_1143);
nand U4578 (N_4578,N_2273,N_1057);
nand U4579 (N_4579,N_1748,N_1007);
nand U4580 (N_4580,N_2235,N_1343);
and U4581 (N_4581,N_2372,N_2128);
xnor U4582 (N_4582,N_861,N_1087);
nand U4583 (N_4583,N_496,N_1043);
nor U4584 (N_4584,N_288,N_1359);
nand U4585 (N_4585,N_274,N_1064);
and U4586 (N_4586,N_893,N_1371);
nand U4587 (N_4587,N_284,N_1962);
nand U4588 (N_4588,N_1923,N_116);
xnor U4589 (N_4589,N_143,N_327);
and U4590 (N_4590,N_308,N_2281);
or U4591 (N_4591,N_772,N_1858);
xor U4592 (N_4592,N_2128,N_1046);
nor U4593 (N_4593,N_1557,N_496);
or U4594 (N_4594,N_1163,N_1303);
or U4595 (N_4595,N_2381,N_1927);
or U4596 (N_4596,N_807,N_519);
nand U4597 (N_4597,N_2499,N_2423);
nor U4598 (N_4598,N_748,N_190);
xor U4599 (N_4599,N_363,N_281);
nor U4600 (N_4600,N_381,N_1161);
or U4601 (N_4601,N_928,N_520);
nand U4602 (N_4602,N_2455,N_516);
or U4603 (N_4603,N_1361,N_2328);
xor U4604 (N_4604,N_2423,N_968);
nand U4605 (N_4605,N_1766,N_1529);
xnor U4606 (N_4606,N_2185,N_272);
and U4607 (N_4607,N_1785,N_1715);
or U4608 (N_4608,N_184,N_681);
nor U4609 (N_4609,N_917,N_25);
nor U4610 (N_4610,N_1470,N_295);
nor U4611 (N_4611,N_263,N_1838);
nor U4612 (N_4612,N_2406,N_1498);
nand U4613 (N_4613,N_48,N_449);
nor U4614 (N_4614,N_2125,N_1766);
or U4615 (N_4615,N_1752,N_2468);
nand U4616 (N_4616,N_935,N_1874);
xnor U4617 (N_4617,N_1408,N_2335);
or U4618 (N_4618,N_53,N_380);
nand U4619 (N_4619,N_1585,N_1711);
or U4620 (N_4620,N_1286,N_2242);
or U4621 (N_4621,N_1950,N_942);
nor U4622 (N_4622,N_1805,N_2179);
or U4623 (N_4623,N_2405,N_1556);
or U4624 (N_4624,N_1091,N_1470);
nor U4625 (N_4625,N_2199,N_1514);
nor U4626 (N_4626,N_2218,N_1148);
and U4627 (N_4627,N_1748,N_315);
or U4628 (N_4628,N_789,N_1540);
nand U4629 (N_4629,N_2173,N_133);
and U4630 (N_4630,N_2464,N_1895);
and U4631 (N_4631,N_1192,N_160);
and U4632 (N_4632,N_2409,N_2342);
and U4633 (N_4633,N_1123,N_567);
or U4634 (N_4634,N_1135,N_321);
and U4635 (N_4635,N_930,N_1810);
nor U4636 (N_4636,N_1867,N_1820);
and U4637 (N_4637,N_1254,N_1558);
nor U4638 (N_4638,N_410,N_333);
or U4639 (N_4639,N_2168,N_1998);
nand U4640 (N_4640,N_330,N_1803);
or U4641 (N_4641,N_1432,N_2295);
nand U4642 (N_4642,N_1999,N_1849);
or U4643 (N_4643,N_2408,N_926);
nor U4644 (N_4644,N_1496,N_2203);
nand U4645 (N_4645,N_1979,N_2018);
and U4646 (N_4646,N_1208,N_108);
or U4647 (N_4647,N_443,N_2346);
or U4648 (N_4648,N_1601,N_1065);
or U4649 (N_4649,N_238,N_1150);
nor U4650 (N_4650,N_2134,N_1201);
nand U4651 (N_4651,N_2238,N_519);
nand U4652 (N_4652,N_693,N_620);
or U4653 (N_4653,N_1360,N_1002);
nor U4654 (N_4654,N_607,N_1134);
and U4655 (N_4655,N_2419,N_2483);
nand U4656 (N_4656,N_484,N_2243);
nor U4657 (N_4657,N_2480,N_462);
and U4658 (N_4658,N_697,N_2496);
nand U4659 (N_4659,N_553,N_1510);
and U4660 (N_4660,N_2448,N_908);
nor U4661 (N_4661,N_626,N_2099);
and U4662 (N_4662,N_1222,N_1244);
nand U4663 (N_4663,N_2399,N_548);
nand U4664 (N_4664,N_2321,N_735);
nor U4665 (N_4665,N_1893,N_1290);
or U4666 (N_4666,N_1956,N_1287);
nor U4667 (N_4667,N_179,N_152);
nor U4668 (N_4668,N_1320,N_322);
nand U4669 (N_4669,N_1251,N_1677);
nor U4670 (N_4670,N_879,N_2033);
nor U4671 (N_4671,N_516,N_882);
xnor U4672 (N_4672,N_2278,N_2151);
or U4673 (N_4673,N_577,N_959);
and U4674 (N_4674,N_40,N_206);
nor U4675 (N_4675,N_1065,N_431);
and U4676 (N_4676,N_2223,N_1165);
and U4677 (N_4677,N_2182,N_136);
nor U4678 (N_4678,N_1779,N_2375);
nor U4679 (N_4679,N_335,N_1758);
nand U4680 (N_4680,N_1416,N_1767);
and U4681 (N_4681,N_2345,N_1985);
and U4682 (N_4682,N_2020,N_530);
and U4683 (N_4683,N_1222,N_1996);
nor U4684 (N_4684,N_1456,N_2076);
and U4685 (N_4685,N_1433,N_1920);
and U4686 (N_4686,N_1393,N_1534);
nor U4687 (N_4687,N_981,N_880);
or U4688 (N_4688,N_335,N_1166);
or U4689 (N_4689,N_1110,N_788);
or U4690 (N_4690,N_287,N_60);
nand U4691 (N_4691,N_926,N_2053);
or U4692 (N_4692,N_1918,N_975);
and U4693 (N_4693,N_1240,N_1561);
nand U4694 (N_4694,N_495,N_2089);
nor U4695 (N_4695,N_1519,N_1421);
and U4696 (N_4696,N_1062,N_149);
nor U4697 (N_4697,N_1406,N_437);
nand U4698 (N_4698,N_657,N_1941);
xnor U4699 (N_4699,N_1369,N_2417);
nor U4700 (N_4700,N_1487,N_1250);
or U4701 (N_4701,N_1028,N_533);
nand U4702 (N_4702,N_1982,N_617);
nand U4703 (N_4703,N_1348,N_428);
nor U4704 (N_4704,N_587,N_1064);
and U4705 (N_4705,N_269,N_1588);
nor U4706 (N_4706,N_1516,N_2315);
nor U4707 (N_4707,N_189,N_2069);
or U4708 (N_4708,N_2128,N_1684);
and U4709 (N_4709,N_2230,N_881);
or U4710 (N_4710,N_2235,N_1859);
or U4711 (N_4711,N_703,N_341);
nor U4712 (N_4712,N_2047,N_1792);
nand U4713 (N_4713,N_2227,N_1613);
nor U4714 (N_4714,N_574,N_1745);
nand U4715 (N_4715,N_1404,N_2278);
or U4716 (N_4716,N_1173,N_2215);
and U4717 (N_4717,N_918,N_1832);
or U4718 (N_4718,N_132,N_1353);
and U4719 (N_4719,N_765,N_2269);
and U4720 (N_4720,N_2291,N_2164);
nand U4721 (N_4721,N_260,N_1542);
nor U4722 (N_4722,N_2404,N_1674);
nor U4723 (N_4723,N_2225,N_216);
nand U4724 (N_4724,N_679,N_1024);
and U4725 (N_4725,N_295,N_2152);
or U4726 (N_4726,N_251,N_914);
or U4727 (N_4727,N_169,N_2249);
and U4728 (N_4728,N_742,N_1626);
and U4729 (N_4729,N_1183,N_366);
or U4730 (N_4730,N_787,N_1243);
nor U4731 (N_4731,N_1168,N_2163);
nand U4732 (N_4732,N_50,N_1894);
nand U4733 (N_4733,N_1817,N_997);
nor U4734 (N_4734,N_2297,N_1143);
or U4735 (N_4735,N_1724,N_53);
nor U4736 (N_4736,N_481,N_902);
nor U4737 (N_4737,N_1574,N_183);
or U4738 (N_4738,N_1049,N_324);
and U4739 (N_4739,N_1970,N_925);
and U4740 (N_4740,N_597,N_1295);
and U4741 (N_4741,N_2310,N_1471);
or U4742 (N_4742,N_500,N_1862);
or U4743 (N_4743,N_876,N_204);
nor U4744 (N_4744,N_294,N_870);
or U4745 (N_4745,N_402,N_1588);
xnor U4746 (N_4746,N_943,N_19);
and U4747 (N_4747,N_1870,N_1252);
and U4748 (N_4748,N_1058,N_711);
nor U4749 (N_4749,N_2416,N_635);
or U4750 (N_4750,N_668,N_1975);
or U4751 (N_4751,N_613,N_1036);
nand U4752 (N_4752,N_500,N_799);
nor U4753 (N_4753,N_645,N_1324);
and U4754 (N_4754,N_281,N_939);
nand U4755 (N_4755,N_337,N_2208);
and U4756 (N_4756,N_1288,N_1146);
nor U4757 (N_4757,N_963,N_547);
and U4758 (N_4758,N_2446,N_1618);
nor U4759 (N_4759,N_1006,N_736);
and U4760 (N_4760,N_2254,N_345);
xor U4761 (N_4761,N_1970,N_2320);
or U4762 (N_4762,N_1166,N_2370);
or U4763 (N_4763,N_2172,N_564);
nor U4764 (N_4764,N_354,N_2135);
and U4765 (N_4765,N_2345,N_301);
nor U4766 (N_4766,N_1724,N_409);
and U4767 (N_4767,N_1855,N_2216);
nor U4768 (N_4768,N_1912,N_1067);
nor U4769 (N_4769,N_796,N_1192);
nor U4770 (N_4770,N_1181,N_619);
and U4771 (N_4771,N_751,N_2367);
or U4772 (N_4772,N_850,N_499);
nor U4773 (N_4773,N_1724,N_1430);
and U4774 (N_4774,N_668,N_715);
nor U4775 (N_4775,N_1797,N_660);
nor U4776 (N_4776,N_2331,N_1627);
and U4777 (N_4777,N_1887,N_193);
nand U4778 (N_4778,N_1995,N_586);
and U4779 (N_4779,N_1917,N_2381);
nand U4780 (N_4780,N_1634,N_938);
or U4781 (N_4781,N_829,N_2222);
nand U4782 (N_4782,N_1773,N_1947);
nor U4783 (N_4783,N_1777,N_649);
nor U4784 (N_4784,N_2490,N_1665);
and U4785 (N_4785,N_853,N_918);
nor U4786 (N_4786,N_2155,N_1624);
nand U4787 (N_4787,N_1957,N_857);
and U4788 (N_4788,N_2186,N_2086);
and U4789 (N_4789,N_606,N_344);
nor U4790 (N_4790,N_747,N_1506);
nor U4791 (N_4791,N_2117,N_570);
nand U4792 (N_4792,N_680,N_1746);
nor U4793 (N_4793,N_785,N_854);
or U4794 (N_4794,N_2142,N_1321);
nand U4795 (N_4795,N_2425,N_421);
nand U4796 (N_4796,N_685,N_2136);
xnor U4797 (N_4797,N_527,N_504);
and U4798 (N_4798,N_848,N_1711);
and U4799 (N_4799,N_557,N_9);
nor U4800 (N_4800,N_1473,N_1849);
nand U4801 (N_4801,N_778,N_1614);
and U4802 (N_4802,N_135,N_2165);
and U4803 (N_4803,N_1174,N_683);
nand U4804 (N_4804,N_1470,N_2104);
nor U4805 (N_4805,N_291,N_756);
nor U4806 (N_4806,N_1845,N_488);
nand U4807 (N_4807,N_1584,N_1272);
or U4808 (N_4808,N_294,N_333);
nor U4809 (N_4809,N_1390,N_1511);
and U4810 (N_4810,N_2281,N_155);
xor U4811 (N_4811,N_263,N_748);
or U4812 (N_4812,N_1636,N_1611);
nor U4813 (N_4813,N_1161,N_1090);
or U4814 (N_4814,N_2243,N_1961);
or U4815 (N_4815,N_729,N_2497);
or U4816 (N_4816,N_245,N_817);
xor U4817 (N_4817,N_1229,N_295);
and U4818 (N_4818,N_401,N_209);
nor U4819 (N_4819,N_2496,N_536);
nand U4820 (N_4820,N_512,N_692);
nand U4821 (N_4821,N_1346,N_2113);
nand U4822 (N_4822,N_759,N_910);
or U4823 (N_4823,N_1924,N_636);
nand U4824 (N_4824,N_1048,N_1233);
nand U4825 (N_4825,N_2213,N_1432);
and U4826 (N_4826,N_748,N_1039);
and U4827 (N_4827,N_1294,N_907);
xor U4828 (N_4828,N_226,N_2357);
or U4829 (N_4829,N_1591,N_47);
nand U4830 (N_4830,N_507,N_838);
nand U4831 (N_4831,N_1243,N_1184);
nor U4832 (N_4832,N_1965,N_1864);
or U4833 (N_4833,N_1884,N_2323);
or U4834 (N_4834,N_1901,N_1186);
xnor U4835 (N_4835,N_187,N_1387);
nor U4836 (N_4836,N_274,N_622);
or U4837 (N_4837,N_2213,N_2375);
nand U4838 (N_4838,N_2009,N_1268);
nor U4839 (N_4839,N_2184,N_1490);
nand U4840 (N_4840,N_1373,N_2486);
or U4841 (N_4841,N_1541,N_648);
and U4842 (N_4842,N_1166,N_2139);
and U4843 (N_4843,N_894,N_958);
and U4844 (N_4844,N_1495,N_1311);
and U4845 (N_4845,N_910,N_1979);
nor U4846 (N_4846,N_619,N_1219);
nand U4847 (N_4847,N_642,N_1347);
and U4848 (N_4848,N_4,N_217);
or U4849 (N_4849,N_1420,N_619);
nand U4850 (N_4850,N_92,N_1430);
and U4851 (N_4851,N_2209,N_2085);
and U4852 (N_4852,N_1329,N_52);
nor U4853 (N_4853,N_1801,N_2361);
or U4854 (N_4854,N_983,N_154);
and U4855 (N_4855,N_1914,N_2101);
or U4856 (N_4856,N_2054,N_767);
or U4857 (N_4857,N_2144,N_571);
and U4858 (N_4858,N_910,N_1802);
or U4859 (N_4859,N_2126,N_839);
or U4860 (N_4860,N_2299,N_1701);
or U4861 (N_4861,N_1890,N_1733);
nand U4862 (N_4862,N_1551,N_1320);
nand U4863 (N_4863,N_2432,N_2427);
or U4864 (N_4864,N_1731,N_2126);
nand U4865 (N_4865,N_2083,N_187);
and U4866 (N_4866,N_2000,N_865);
xor U4867 (N_4867,N_2211,N_2333);
or U4868 (N_4868,N_1431,N_53);
nor U4869 (N_4869,N_2244,N_994);
or U4870 (N_4870,N_890,N_950);
nand U4871 (N_4871,N_1816,N_1842);
or U4872 (N_4872,N_1530,N_2002);
or U4873 (N_4873,N_391,N_1048);
nor U4874 (N_4874,N_93,N_1707);
xnor U4875 (N_4875,N_285,N_1602);
and U4876 (N_4876,N_2336,N_1118);
nand U4877 (N_4877,N_246,N_755);
nand U4878 (N_4878,N_2311,N_128);
nand U4879 (N_4879,N_926,N_1495);
xnor U4880 (N_4880,N_689,N_2197);
or U4881 (N_4881,N_1871,N_2181);
nand U4882 (N_4882,N_2344,N_168);
xor U4883 (N_4883,N_1738,N_661);
nand U4884 (N_4884,N_1143,N_242);
and U4885 (N_4885,N_1838,N_2057);
and U4886 (N_4886,N_1981,N_1280);
nand U4887 (N_4887,N_1810,N_410);
nor U4888 (N_4888,N_2084,N_1366);
and U4889 (N_4889,N_1721,N_84);
xor U4890 (N_4890,N_296,N_1592);
nand U4891 (N_4891,N_2003,N_1165);
nand U4892 (N_4892,N_673,N_2226);
and U4893 (N_4893,N_498,N_774);
or U4894 (N_4894,N_576,N_56);
and U4895 (N_4895,N_1020,N_816);
xor U4896 (N_4896,N_1515,N_776);
nand U4897 (N_4897,N_853,N_1355);
and U4898 (N_4898,N_1274,N_330);
nand U4899 (N_4899,N_811,N_18);
nand U4900 (N_4900,N_747,N_62);
or U4901 (N_4901,N_501,N_287);
nor U4902 (N_4902,N_642,N_197);
nor U4903 (N_4903,N_2346,N_1055);
nor U4904 (N_4904,N_1959,N_1924);
nor U4905 (N_4905,N_1667,N_1081);
and U4906 (N_4906,N_1604,N_958);
and U4907 (N_4907,N_302,N_647);
and U4908 (N_4908,N_359,N_1259);
or U4909 (N_4909,N_2112,N_1088);
and U4910 (N_4910,N_2355,N_2397);
nor U4911 (N_4911,N_268,N_211);
nand U4912 (N_4912,N_1785,N_905);
nand U4913 (N_4913,N_1536,N_1806);
and U4914 (N_4914,N_1486,N_539);
and U4915 (N_4915,N_1856,N_1832);
nor U4916 (N_4916,N_69,N_2178);
and U4917 (N_4917,N_546,N_1155);
or U4918 (N_4918,N_1952,N_980);
nor U4919 (N_4919,N_1353,N_312);
or U4920 (N_4920,N_1824,N_2416);
nor U4921 (N_4921,N_1751,N_2487);
nand U4922 (N_4922,N_1053,N_1852);
nand U4923 (N_4923,N_2067,N_449);
or U4924 (N_4924,N_192,N_2364);
xor U4925 (N_4925,N_1627,N_1580);
or U4926 (N_4926,N_1410,N_1779);
nor U4927 (N_4927,N_181,N_1392);
nor U4928 (N_4928,N_1623,N_374);
or U4929 (N_4929,N_1262,N_354);
or U4930 (N_4930,N_1585,N_1567);
nand U4931 (N_4931,N_1197,N_1029);
or U4932 (N_4932,N_95,N_108);
and U4933 (N_4933,N_494,N_907);
or U4934 (N_4934,N_993,N_417);
nand U4935 (N_4935,N_58,N_1473);
and U4936 (N_4936,N_813,N_591);
and U4937 (N_4937,N_1746,N_7);
or U4938 (N_4938,N_225,N_1640);
or U4939 (N_4939,N_622,N_773);
nor U4940 (N_4940,N_2316,N_67);
and U4941 (N_4941,N_881,N_1377);
nor U4942 (N_4942,N_239,N_120);
or U4943 (N_4943,N_2457,N_117);
or U4944 (N_4944,N_1808,N_1689);
xor U4945 (N_4945,N_129,N_1102);
or U4946 (N_4946,N_477,N_2203);
nand U4947 (N_4947,N_1080,N_2);
or U4948 (N_4948,N_1768,N_1089);
or U4949 (N_4949,N_1235,N_1155);
nand U4950 (N_4950,N_2011,N_889);
nor U4951 (N_4951,N_2336,N_487);
nand U4952 (N_4952,N_1438,N_436);
or U4953 (N_4953,N_1896,N_1419);
nor U4954 (N_4954,N_633,N_1376);
nor U4955 (N_4955,N_2212,N_1807);
nor U4956 (N_4956,N_2023,N_137);
nor U4957 (N_4957,N_2133,N_2220);
or U4958 (N_4958,N_1666,N_144);
and U4959 (N_4959,N_610,N_1679);
xor U4960 (N_4960,N_2379,N_1272);
nand U4961 (N_4961,N_131,N_1299);
or U4962 (N_4962,N_1095,N_539);
nand U4963 (N_4963,N_206,N_1801);
nor U4964 (N_4964,N_309,N_257);
or U4965 (N_4965,N_757,N_321);
and U4966 (N_4966,N_1306,N_1935);
and U4967 (N_4967,N_273,N_418);
or U4968 (N_4968,N_281,N_858);
and U4969 (N_4969,N_1994,N_2028);
nand U4970 (N_4970,N_2056,N_169);
or U4971 (N_4971,N_765,N_1486);
and U4972 (N_4972,N_1383,N_547);
or U4973 (N_4973,N_1226,N_2176);
nor U4974 (N_4974,N_445,N_2174);
and U4975 (N_4975,N_216,N_1667);
and U4976 (N_4976,N_1218,N_962);
or U4977 (N_4977,N_1960,N_1161);
and U4978 (N_4978,N_1920,N_1483);
nand U4979 (N_4979,N_1177,N_2038);
nor U4980 (N_4980,N_1764,N_2064);
or U4981 (N_4981,N_438,N_1532);
nand U4982 (N_4982,N_1312,N_3);
and U4983 (N_4983,N_434,N_90);
xor U4984 (N_4984,N_192,N_349);
and U4985 (N_4985,N_1885,N_1670);
or U4986 (N_4986,N_503,N_754);
nor U4987 (N_4987,N_462,N_1415);
nor U4988 (N_4988,N_1801,N_54);
or U4989 (N_4989,N_1720,N_1173);
or U4990 (N_4990,N_1687,N_1579);
and U4991 (N_4991,N_52,N_2440);
nor U4992 (N_4992,N_1094,N_1000);
nor U4993 (N_4993,N_341,N_1114);
or U4994 (N_4994,N_156,N_917);
and U4995 (N_4995,N_2021,N_748);
nand U4996 (N_4996,N_1922,N_1187);
nand U4997 (N_4997,N_859,N_468);
nand U4998 (N_4998,N_1272,N_2019);
and U4999 (N_4999,N_2213,N_2455);
or UO_0 (O_0,N_2973,N_3164);
and UO_1 (O_1,N_3453,N_4463);
nor UO_2 (O_2,N_2870,N_3969);
nand UO_3 (O_3,N_3540,N_2686);
or UO_4 (O_4,N_4414,N_4310);
or UO_5 (O_5,N_4046,N_3998);
and UO_6 (O_6,N_4649,N_2700);
nor UO_7 (O_7,N_4430,N_3040);
nand UO_8 (O_8,N_2580,N_3810);
and UO_9 (O_9,N_4391,N_3852);
nor UO_10 (O_10,N_4081,N_4425);
and UO_11 (O_11,N_2938,N_4062);
xnor UO_12 (O_12,N_4003,N_4017);
nor UO_13 (O_13,N_2908,N_2819);
and UO_14 (O_14,N_4915,N_4080);
or UO_15 (O_15,N_3977,N_4213);
nand UO_16 (O_16,N_3273,N_4260);
nand UO_17 (O_17,N_3071,N_3510);
nor UO_18 (O_18,N_4556,N_2567);
nand UO_19 (O_19,N_4488,N_4336);
and UO_20 (O_20,N_4658,N_3298);
nor UO_21 (O_21,N_2564,N_4661);
nand UO_22 (O_22,N_3099,N_2500);
or UO_23 (O_23,N_4795,N_2941);
nor UO_24 (O_24,N_4949,N_3950);
nor UO_25 (O_25,N_3518,N_4573);
nand UO_26 (O_26,N_4595,N_4115);
nand UO_27 (O_27,N_4449,N_4778);
and UO_28 (O_28,N_4734,N_2692);
or UO_29 (O_29,N_2967,N_3669);
or UO_30 (O_30,N_3014,N_2701);
nor UO_31 (O_31,N_3761,N_3159);
nand UO_32 (O_32,N_3770,N_2615);
nor UO_33 (O_33,N_4472,N_3897);
and UO_34 (O_34,N_4651,N_4292);
or UO_35 (O_35,N_3709,N_4404);
or UO_36 (O_36,N_4354,N_2805);
or UO_37 (O_37,N_2556,N_3804);
or UO_38 (O_38,N_3679,N_3559);
or UO_39 (O_39,N_4769,N_4802);
nor UO_40 (O_40,N_3477,N_2610);
nor UO_41 (O_41,N_3766,N_3005);
nor UO_42 (O_42,N_4888,N_4137);
and UO_43 (O_43,N_4910,N_4208);
nor UO_44 (O_44,N_3779,N_2964);
nand UO_45 (O_45,N_2983,N_4005);
or UO_46 (O_46,N_2750,N_2989);
and UO_47 (O_47,N_3185,N_4913);
nor UO_48 (O_48,N_3255,N_3824);
nor UO_49 (O_49,N_3748,N_4989);
nor UO_50 (O_50,N_4852,N_3557);
nand UO_51 (O_51,N_4130,N_3044);
or UO_52 (O_52,N_3108,N_4681);
nand UO_53 (O_53,N_3090,N_3635);
nor UO_54 (O_54,N_2504,N_4419);
nand UO_55 (O_55,N_3844,N_3241);
and UO_56 (O_56,N_2703,N_3025);
and UO_57 (O_57,N_2520,N_3516);
nand UO_58 (O_58,N_3495,N_4841);
nor UO_59 (O_59,N_2644,N_4848);
nand UO_60 (O_60,N_4221,N_3338);
or UO_61 (O_61,N_4955,N_3747);
xor UO_62 (O_62,N_4593,N_3322);
nor UO_63 (O_63,N_2914,N_2991);
nor UO_64 (O_64,N_3126,N_4890);
and UO_65 (O_65,N_4935,N_4762);
and UO_66 (O_66,N_4546,N_3944);
and UO_67 (O_67,N_4859,N_4772);
nand UO_68 (O_68,N_3306,N_4993);
nor UO_69 (O_69,N_4233,N_2687);
and UO_70 (O_70,N_4611,N_4098);
nand UO_71 (O_71,N_4028,N_3794);
or UO_72 (O_72,N_4280,N_3078);
nand UO_73 (O_73,N_2953,N_4650);
or UO_74 (O_74,N_4059,N_4429);
or UO_75 (O_75,N_4453,N_3200);
and UO_76 (O_76,N_4401,N_4489);
and UO_77 (O_77,N_4986,N_4491);
or UO_78 (O_78,N_3413,N_4904);
or UO_79 (O_79,N_4785,N_2597);
nor UO_80 (O_80,N_2753,N_2714);
nand UO_81 (O_81,N_4945,N_4097);
or UO_82 (O_82,N_3458,N_3067);
nor UO_83 (O_83,N_3716,N_3206);
nand UO_84 (O_84,N_3940,N_3848);
nand UO_85 (O_85,N_2719,N_4591);
and UO_86 (O_86,N_3203,N_4219);
nand UO_87 (O_87,N_3915,N_3585);
and UO_88 (O_88,N_3875,N_3811);
or UO_89 (O_89,N_4975,N_3073);
nand UO_90 (O_90,N_3665,N_4040);
nand UO_91 (O_91,N_4079,N_4492);
and UO_92 (O_92,N_3509,N_3471);
or UO_93 (O_93,N_3544,N_3611);
nand UO_94 (O_94,N_2776,N_3888);
nor UO_95 (O_95,N_4104,N_4660);
or UO_96 (O_96,N_3584,N_3573);
or UO_97 (O_97,N_4107,N_3929);
nand UO_98 (O_98,N_3890,N_4857);
nand UO_99 (O_99,N_4603,N_4416);
or UO_100 (O_100,N_4467,N_3708);
nand UO_101 (O_101,N_4914,N_3696);
and UO_102 (O_102,N_4701,N_4305);
nor UO_103 (O_103,N_3434,N_3472);
nor UO_104 (O_104,N_4202,N_2977);
nand UO_105 (O_105,N_2804,N_3082);
nor UO_106 (O_106,N_2924,N_4946);
nand UO_107 (O_107,N_3214,N_2857);
nor UO_108 (O_108,N_3703,N_4642);
or UO_109 (O_109,N_3764,N_4931);
nor UO_110 (O_110,N_3258,N_4362);
nand UO_111 (O_111,N_4424,N_2678);
or UO_112 (O_112,N_2884,N_3291);
or UO_113 (O_113,N_3480,N_3334);
nor UO_114 (O_114,N_3827,N_2833);
and UO_115 (O_115,N_2710,N_4476);
nor UO_116 (O_116,N_4344,N_4151);
or UO_117 (O_117,N_3400,N_3866);
and UO_118 (O_118,N_4691,N_3776);
or UO_119 (O_119,N_4758,N_2809);
or UO_120 (O_120,N_4728,N_3790);
or UO_121 (O_121,N_4883,N_2928);
nand UO_122 (O_122,N_4714,N_4527);
nor UO_123 (O_123,N_4628,N_3912);
or UO_124 (O_124,N_2845,N_4207);
nor UO_125 (O_125,N_3649,N_3543);
nand UO_126 (O_126,N_4510,N_3909);
and UO_127 (O_127,N_4187,N_3558);
nand UO_128 (O_128,N_3988,N_2942);
xor UO_129 (O_129,N_4794,N_4706);
nand UO_130 (O_130,N_4771,N_4582);
or UO_131 (O_131,N_2842,N_3745);
or UO_132 (O_132,N_3050,N_4049);
or UO_133 (O_133,N_3871,N_4784);
and UO_134 (O_134,N_2743,N_3537);
nand UO_135 (O_135,N_4276,N_3607);
nand UO_136 (O_136,N_4520,N_4405);
nor UO_137 (O_137,N_3692,N_4335);
and UO_138 (O_138,N_3892,N_4631);
or UO_139 (O_139,N_4621,N_2756);
nand UO_140 (O_140,N_2623,N_3659);
nand UO_141 (O_141,N_4893,N_3194);
or UO_142 (O_142,N_3647,N_4695);
nor UO_143 (O_143,N_2716,N_2931);
xor UO_144 (O_144,N_3928,N_4932);
nor UO_145 (O_145,N_4513,N_4704);
nand UO_146 (O_146,N_4668,N_3956);
nand UO_147 (O_147,N_4930,N_2598);
nand UO_148 (O_148,N_3807,N_4629);
and UO_149 (O_149,N_2503,N_4131);
nor UO_150 (O_150,N_2769,N_4188);
nor UO_151 (O_151,N_4176,N_2543);
and UO_152 (O_152,N_3881,N_3248);
nor UO_153 (O_153,N_2791,N_4171);
nand UO_154 (O_154,N_4540,N_4092);
nor UO_155 (O_155,N_4365,N_3846);
nand UO_156 (O_156,N_4381,N_3115);
or UO_157 (O_157,N_2649,N_2988);
nor UO_158 (O_158,N_4690,N_3538);
and UO_159 (O_159,N_3795,N_4474);
or UO_160 (O_160,N_2666,N_3043);
or UO_161 (O_161,N_4172,N_3309);
nor UO_162 (O_162,N_3297,N_3282);
or UO_163 (O_163,N_2837,N_4947);
or UO_164 (O_164,N_3227,N_4625);
nor UO_165 (O_165,N_4657,N_4534);
nor UO_166 (O_166,N_3843,N_2604);
xnor UO_167 (O_167,N_3269,N_3514);
nand UO_168 (O_168,N_3324,N_3343);
nand UO_169 (O_169,N_3570,N_3140);
and UO_170 (O_170,N_3974,N_3639);
and UO_171 (O_171,N_4122,N_4501);
nand UO_172 (O_172,N_4756,N_4206);
or UO_173 (O_173,N_4000,N_4633);
nor UO_174 (O_174,N_3860,N_3473);
nand UO_175 (O_175,N_2529,N_4466);
nand UO_176 (O_176,N_3033,N_3321);
or UO_177 (O_177,N_2954,N_2746);
and UO_178 (O_178,N_3110,N_2696);
nand UO_179 (O_179,N_3080,N_3902);
nand UO_180 (O_180,N_4824,N_3167);
or UO_181 (O_181,N_3394,N_2950);
and UO_182 (O_182,N_4006,N_2995);
or UO_183 (O_183,N_2881,N_4117);
nor UO_184 (O_184,N_2685,N_4380);
or UO_185 (O_185,N_4431,N_4542);
nor UO_186 (O_186,N_3781,N_4239);
nor UO_187 (O_187,N_3259,N_2534);
and UO_188 (O_188,N_4994,N_4519);
or UO_189 (O_189,N_3426,N_4584);
or UO_190 (O_190,N_4600,N_4161);
or UO_191 (O_191,N_2603,N_3657);
nand UO_192 (O_192,N_3318,N_3358);
or UO_193 (O_193,N_4786,N_4110);
nand UO_194 (O_194,N_4123,N_3268);
nor UO_195 (O_195,N_3530,N_2771);
nand UO_196 (O_196,N_3450,N_3160);
nand UO_197 (O_197,N_4789,N_3681);
or UO_198 (O_198,N_2506,N_2717);
or UO_199 (O_199,N_2725,N_3729);
nor UO_200 (O_200,N_4103,N_4504);
and UO_201 (O_201,N_4317,N_4035);
nor UO_202 (O_202,N_3722,N_3264);
nor UO_203 (O_203,N_4992,N_3975);
or UO_204 (O_204,N_3486,N_4495);
nand UO_205 (O_205,N_4348,N_3459);
nor UO_206 (O_206,N_4751,N_3534);
or UO_207 (O_207,N_3094,N_2742);
and UO_208 (O_208,N_4274,N_3616);
nor UO_209 (O_209,N_2729,N_2501);
and UO_210 (O_210,N_3777,N_3373);
nand UO_211 (O_211,N_3971,N_3934);
and UO_212 (O_212,N_4766,N_4417);
xnor UO_213 (O_213,N_4999,N_3701);
and UO_214 (O_214,N_2925,N_3615);
nand UO_215 (O_215,N_2866,N_2937);
or UO_216 (O_216,N_2957,N_4470);
and UO_217 (O_217,N_3880,N_2897);
nor UO_218 (O_218,N_3354,N_4262);
and UO_219 (O_219,N_4361,N_4352);
nand UO_220 (O_220,N_4494,N_3684);
and UO_221 (O_221,N_4421,N_2611);
and UO_222 (O_222,N_4783,N_3246);
nand UO_223 (O_223,N_3086,N_4805);
and UO_224 (O_224,N_3346,N_4141);
or UO_225 (O_225,N_3571,N_3721);
or UO_226 (O_226,N_4809,N_4828);
and UO_227 (O_227,N_4316,N_4067);
and UO_228 (O_228,N_3889,N_4443);
or UO_229 (O_229,N_2843,N_4030);
or UO_230 (O_230,N_3650,N_3997);
or UO_231 (O_231,N_4780,N_3491);
and UO_232 (O_232,N_4441,N_3823);
nor UO_233 (O_233,N_3667,N_3386);
nand UO_234 (O_234,N_2637,N_4083);
and UO_235 (O_235,N_3300,N_4654);
nor UO_236 (O_236,N_4604,N_4683);
and UO_237 (O_237,N_3964,N_3731);
nor UO_238 (O_238,N_4745,N_2559);
nor UO_239 (O_239,N_4058,N_4039);
or UO_240 (O_240,N_3328,N_2680);
or UO_241 (O_241,N_2679,N_3966);
or UO_242 (O_242,N_2927,N_2658);
nand UO_243 (O_243,N_4738,N_3007);
or UO_244 (O_244,N_3008,N_4002);
and UO_245 (O_245,N_3831,N_4355);
and UO_246 (O_246,N_2913,N_4368);
nor UO_247 (O_247,N_3065,N_4749);
nor UO_248 (O_248,N_4249,N_4623);
and UO_249 (O_249,N_4246,N_4928);
nand UO_250 (O_250,N_2539,N_3801);
nor UO_251 (O_251,N_4118,N_4145);
and UO_252 (O_252,N_2785,N_4620);
nor UO_253 (O_253,N_4457,N_3965);
nor UO_254 (O_254,N_3213,N_3271);
and UO_255 (O_255,N_4294,N_2640);
nand UO_256 (O_256,N_4272,N_2517);
and UO_257 (O_257,N_4291,N_4906);
nor UO_258 (O_258,N_3628,N_3515);
nand UO_259 (O_259,N_4029,N_3528);
nand UO_260 (O_260,N_2826,N_2772);
and UO_261 (O_261,N_4210,N_2782);
nand UO_262 (O_262,N_3726,N_4076);
nor UO_263 (O_263,N_3945,N_3855);
nand UO_264 (O_264,N_4064,N_2909);
or UO_265 (O_265,N_4635,N_4068);
and UO_266 (O_266,N_4830,N_4451);
nor UO_267 (O_267,N_4108,N_3617);
xnor UO_268 (O_268,N_4340,N_4089);
and UO_269 (O_269,N_4833,N_4656);
or UO_270 (O_270,N_2655,N_4426);
nand UO_271 (O_271,N_4663,N_2869);
or UO_272 (O_272,N_4517,N_4829);
or UO_273 (O_273,N_2966,N_4579);
or UO_274 (O_274,N_4987,N_2802);
or UO_275 (O_275,N_3131,N_4200);
nor UO_276 (O_276,N_2568,N_4933);
or UO_277 (O_277,N_2627,N_3626);
nand UO_278 (O_278,N_2732,N_3762);
nor UO_279 (O_279,N_4875,N_4251);
or UO_280 (O_280,N_2693,N_3497);
nor UO_281 (O_281,N_3587,N_2906);
nand UO_282 (O_282,N_3148,N_3381);
or UO_283 (O_283,N_4015,N_4514);
nand UO_284 (O_284,N_2536,N_2828);
nor UO_285 (O_285,N_4735,N_2675);
and UO_286 (O_286,N_4224,N_4832);
nor UO_287 (O_287,N_2561,N_4211);
nand UO_288 (O_288,N_4326,N_3045);
and UO_289 (O_289,N_4259,N_3092);
nor UO_290 (O_290,N_3813,N_2653);
nand UO_291 (O_291,N_4371,N_3188);
and UO_292 (O_292,N_3052,N_4136);
or UO_293 (O_293,N_4912,N_4707);
nand UO_294 (O_294,N_3666,N_3668);
nand UO_295 (O_295,N_4662,N_2786);
nor UO_296 (O_296,N_3589,N_4982);
or UO_297 (O_297,N_4334,N_4612);
nand UO_298 (O_298,N_3404,N_2745);
nor UO_299 (O_299,N_4962,N_2919);
nand UO_300 (O_300,N_4816,N_4922);
nand UO_301 (O_301,N_4382,N_3238);
nand UO_302 (O_302,N_4997,N_3914);
nor UO_303 (O_303,N_2549,N_4776);
and UO_304 (O_304,N_3979,N_4587);
nor UO_305 (O_305,N_3498,N_2639);
or UO_306 (O_306,N_2522,N_2645);
and UO_307 (O_307,N_3116,N_4552);
and UO_308 (O_308,N_4082,N_4370);
and UO_309 (O_309,N_3493,N_4008);
nor UO_310 (O_310,N_2733,N_4140);
nor UO_311 (O_311,N_4899,N_4525);
nor UO_312 (O_312,N_4164,N_4613);
or UO_313 (O_313,N_4843,N_3370);
nand UO_314 (O_314,N_4498,N_4284);
nand UO_315 (O_315,N_4422,N_4351);
and UO_316 (O_316,N_2705,N_4399);
nor UO_317 (O_317,N_3872,N_4521);
and UO_318 (O_318,N_3266,N_3139);
and UO_319 (O_319,N_3583,N_4605);
and UO_320 (O_320,N_4041,N_4858);
and UO_321 (O_321,N_4709,N_2558);
nand UO_322 (O_322,N_3536,N_3469);
nor UO_323 (O_323,N_4315,N_3249);
nor UO_324 (O_324,N_4580,N_3973);
xor UO_325 (O_325,N_3433,N_2669);
nand UO_326 (O_326,N_2563,N_4452);
nor UO_327 (O_327,N_3636,N_4528);
xnor UO_328 (O_328,N_3062,N_4967);
or UO_329 (O_329,N_4235,N_3020);
and UO_330 (O_330,N_3177,N_3676);
or UO_331 (O_331,N_3519,N_3754);
nand UO_332 (O_332,N_3847,N_3767);
or UO_333 (O_333,N_3329,N_2647);
nor UO_334 (O_334,N_4970,N_4741);
or UO_335 (O_335,N_3125,N_4054);
nand UO_336 (O_336,N_3478,N_3027);
or UO_337 (O_337,N_4506,N_4109);
and UO_338 (O_338,N_4886,N_4637);
and UO_339 (O_339,N_3387,N_2668);
nand UO_340 (O_340,N_2508,N_2984);
nand UO_341 (O_341,N_3691,N_3079);
and UO_342 (O_342,N_2648,N_2523);
nand UO_343 (O_343,N_2841,N_3372);
and UO_344 (O_344,N_3161,N_4375);
nor UO_345 (O_345,N_3752,N_3986);
or UO_346 (O_346,N_2811,N_2918);
or UO_347 (O_347,N_4071,N_4066);
or UO_348 (O_348,N_4415,N_4461);
nand UO_349 (O_349,N_3857,N_4245);
nor UO_350 (O_350,N_3484,N_2661);
and UO_351 (O_351,N_3326,N_3948);
nor UO_352 (O_352,N_3319,N_2917);
or UO_353 (O_353,N_2929,N_3402);
nor UO_354 (O_354,N_2850,N_4197);
or UO_355 (O_355,N_3211,N_4974);
and UO_356 (O_356,N_4312,N_4273);
xor UO_357 (O_357,N_2723,N_4223);
nand UO_358 (O_358,N_2540,N_3580);
nor UO_359 (O_359,N_4705,N_3209);
nand UO_360 (O_360,N_4831,N_3654);
and UO_361 (O_361,N_4085,N_3438);
nor UO_362 (O_362,N_2981,N_3891);
or UO_363 (O_363,N_2982,N_3347);
nand UO_364 (O_364,N_3771,N_3038);
nand UO_365 (O_365,N_4400,N_4432);
and UO_366 (O_366,N_4177,N_4634);
nand UO_367 (O_367,N_2755,N_2820);
or UO_368 (O_368,N_4748,N_3385);
nor UO_369 (O_369,N_2528,N_4574);
nor UO_370 (O_370,N_4867,N_3586);
nor UO_371 (O_371,N_3368,N_4018);
or UO_372 (O_372,N_4653,N_2861);
and UO_373 (O_373,N_3425,N_2665);
and UO_374 (O_374,N_3562,N_3376);
and UO_375 (O_375,N_4782,N_3903);
and UO_376 (O_376,N_2744,N_3868);
and UO_377 (O_377,N_2760,N_3604);
xor UO_378 (O_378,N_2858,N_4240);
nor UO_379 (O_379,N_3365,N_4996);
and UO_380 (O_380,N_3100,N_4332);
nor UO_381 (O_381,N_4138,N_3512);
nand UO_382 (O_382,N_2821,N_3699);
nand UO_383 (O_383,N_3802,N_3267);
and UO_384 (O_384,N_3792,N_4507);
or UO_385 (O_385,N_3723,N_4877);
and UO_386 (O_386,N_3228,N_4884);
or UO_387 (O_387,N_3784,N_2979);
nand UO_388 (O_388,N_3299,N_4606);
or UO_389 (O_389,N_3183,N_2599);
and UO_390 (O_390,N_4050,N_4610);
or UO_391 (O_391,N_4614,N_4196);
and UO_392 (O_392,N_4937,N_3732);
and UO_393 (O_393,N_4764,N_4919);
nand UO_394 (O_394,N_2636,N_2535);
or UO_395 (O_395,N_2552,N_2694);
nor UO_396 (O_396,N_4343,N_2712);
or UO_397 (O_397,N_4182,N_3310);
nor UO_398 (O_398,N_2783,N_3097);
nand UO_399 (O_399,N_4671,N_3658);
and UO_400 (O_400,N_4965,N_4544);
nand UO_401 (O_401,N_4217,N_4881);
or UO_402 (O_402,N_3833,N_2934);
and UO_403 (O_403,N_3787,N_4522);
nand UO_404 (O_404,N_4724,N_4647);
or UO_405 (O_405,N_4314,N_3618);
nand UO_406 (O_406,N_2634,N_4842);
nand UO_407 (O_407,N_3506,N_4346);
or UO_408 (O_408,N_3734,N_2664);
nand UO_409 (O_409,N_3366,N_4234);
and UO_410 (O_410,N_2848,N_2555);
nand UO_411 (O_411,N_3278,N_4512);
nand UO_412 (O_412,N_2659,N_3350);
or UO_413 (O_413,N_4418,N_3742);
xor UO_414 (O_414,N_2670,N_3378);
and UO_415 (O_415,N_2581,N_4086);
nor UO_416 (O_416,N_2532,N_2997);
and UO_417 (O_417,N_4725,N_4718);
nand UO_418 (O_418,N_3377,N_3621);
nor UO_419 (O_419,N_3653,N_4266);
nand UO_420 (O_420,N_2551,N_4100);
nand UO_421 (O_421,N_4942,N_4929);
xnor UO_422 (O_422,N_4607,N_4566);
or UO_423 (O_423,N_3275,N_2616);
xor UO_424 (O_424,N_3797,N_3642);
or UO_425 (O_425,N_3925,N_2803);
nand UO_426 (O_426,N_2505,N_2650);
or UO_427 (O_427,N_3634,N_4847);
and UO_428 (O_428,N_3619,N_2513);
or UO_429 (O_429,N_4827,N_2633);
nand UO_430 (O_430,N_2872,N_4895);
xor UO_431 (O_431,N_2952,N_3017);
nor UO_432 (O_432,N_4152,N_4732);
nor UO_433 (O_433,N_3409,N_4518);
nand UO_434 (O_434,N_2588,N_2978);
or UO_435 (O_435,N_3895,N_4674);
nor UO_436 (O_436,N_2697,N_4288);
or UO_437 (O_437,N_3380,N_2778);
nor UO_438 (O_438,N_3192,N_3412);
nor UO_439 (O_439,N_4289,N_3348);
and UO_440 (O_440,N_3146,N_4958);
or UO_441 (O_441,N_3717,N_4397);
and UO_442 (O_442,N_2734,N_4125);
or UO_443 (O_443,N_4770,N_2788);
or UO_444 (O_444,N_4433,N_4483);
nor UO_445 (O_445,N_3263,N_4750);
and UO_446 (O_446,N_3523,N_4901);
or UO_447 (O_447,N_4353,N_4252);
nor UO_448 (O_448,N_2943,N_4339);
nand UO_449 (O_449,N_3935,N_3527);
nand UO_450 (O_450,N_4985,N_4720);
nor UO_451 (O_451,N_3706,N_3104);
nor UO_452 (O_452,N_2814,N_4228);
nor UO_453 (O_453,N_4588,N_4057);
nand UO_454 (O_454,N_3886,N_3485);
nand UO_455 (O_455,N_3023,N_4413);
nand UO_456 (O_456,N_4007,N_3593);
nand UO_457 (O_457,N_4420,N_2671);
nor UO_458 (O_458,N_4237,N_4232);
or UO_459 (O_459,N_2830,N_4968);
and UO_460 (O_460,N_3024,N_4508);
nand UO_461 (O_461,N_4227,N_4702);
and UO_462 (O_462,N_3134,N_4411);
or UO_463 (O_463,N_3397,N_4862);
and UO_464 (O_464,N_4423,N_2740);
and UO_465 (O_465,N_2724,N_4025);
nor UO_466 (O_466,N_4977,N_3555);
xor UO_467 (O_467,N_3504,N_3905);
or UO_468 (O_468,N_2970,N_3867);
and UO_469 (O_469,N_2955,N_2565);
nor UO_470 (O_470,N_3660,N_2643);
and UO_471 (O_471,N_2656,N_2509);
and UO_472 (O_472,N_2530,N_3439);
or UO_473 (O_473,N_4920,N_4839);
or UO_474 (O_474,N_3765,N_2922);
and UO_475 (O_475,N_2907,N_4601);
nand UO_476 (O_476,N_3422,N_4953);
and UO_477 (O_477,N_3217,N_4013);
nand UO_478 (O_478,N_2916,N_4686);
nand UO_479 (O_479,N_4909,N_3124);
nor UO_480 (O_480,N_3662,N_3287);
nand UO_481 (O_481,N_4328,N_4927);
nand UO_482 (O_482,N_4047,N_3499);
xnor UO_483 (O_483,N_4821,N_2630);
nand UO_484 (O_484,N_4070,N_3799);
or UO_485 (O_485,N_3632,N_3176);
nor UO_486 (O_486,N_2808,N_3907);
and UO_487 (O_487,N_2832,N_3590);
nor UO_488 (O_488,N_3443,N_3746);
nor UO_489 (O_489,N_2672,N_3449);
nand UO_490 (O_490,N_2515,N_2781);
and UO_491 (O_491,N_2727,N_4667);
and UO_492 (O_492,N_3569,N_3028);
and UO_493 (O_493,N_2602,N_2956);
nand UO_494 (O_494,N_3260,N_4282);
nand UO_495 (O_495,N_4257,N_4133);
nor UO_496 (O_496,N_2545,N_4106);
or UO_497 (O_497,N_2930,N_3293);
and UO_498 (O_498,N_3838,N_3927);
nand UO_499 (O_499,N_3546,N_3393);
and UO_500 (O_500,N_3465,N_4568);
or UO_501 (O_501,N_4768,N_4983);
or UO_502 (O_502,N_3842,N_4860);
and UO_503 (O_503,N_2683,N_4563);
nor UO_504 (O_504,N_3898,N_4575);
nor UO_505 (O_505,N_3218,N_3700);
xnor UO_506 (O_506,N_3496,N_3229);
or UO_507 (O_507,N_2946,N_4479);
nor UO_508 (O_508,N_3288,N_4019);
or UO_509 (O_509,N_3995,N_4490);
and UO_510 (O_510,N_3733,N_3627);
or UO_511 (O_511,N_2605,N_2871);
nor UO_512 (O_512,N_2936,N_3009);
nor UO_513 (O_513,N_3235,N_4477);
and UO_514 (O_514,N_2596,N_4304);
or UO_515 (O_515,N_3087,N_3961);
and UO_516 (O_516,N_4165,N_2932);
or UO_517 (O_517,N_3714,N_4526);
or UO_518 (O_518,N_4812,N_3237);
nand UO_519 (O_519,N_3084,N_4090);
and UO_520 (O_520,N_4338,N_4991);
nand UO_521 (O_521,N_3353,N_3357);
and UO_522 (O_522,N_3989,N_2846);
and UO_523 (O_523,N_4943,N_3602);
nor UO_524 (O_524,N_3193,N_2784);
nand UO_525 (O_525,N_4386,N_3738);
nand UO_526 (O_526,N_3553,N_4088);
or UO_527 (O_527,N_2654,N_4437);
nor UO_528 (O_528,N_3137,N_4547);
and UO_529 (O_529,N_2905,N_4248);
nand UO_530 (O_530,N_4564,N_4265);
and UO_531 (O_531,N_4271,N_3508);
or UO_532 (O_532,N_3575,N_4713);
and UO_533 (O_533,N_3820,N_2895);
or UO_534 (O_534,N_4774,N_4459);
nor UO_535 (O_535,N_4643,N_4435);
or UO_536 (O_536,N_4646,N_4516);
nor UO_537 (O_537,N_4192,N_4889);
nand UO_538 (O_538,N_3170,N_4585);
or UO_539 (O_539,N_3012,N_2795);
xnor UO_540 (O_540,N_3118,N_3013);
nand UO_541 (O_541,N_3865,N_4960);
nor UO_542 (O_542,N_3031,N_3780);
nand UO_543 (O_543,N_3548,N_3436);
and UO_544 (O_544,N_3250,N_4183);
and UO_545 (O_545,N_2815,N_4349);
nor UO_546 (O_546,N_2793,N_3502);
or UO_547 (O_547,N_4390,N_4063);
nand UO_548 (O_548,N_4798,N_4190);
nor UO_549 (O_549,N_4557,N_2904);
or UO_550 (O_550,N_2920,N_2591);
or UO_551 (O_551,N_4333,N_3873);
nor UO_552 (O_552,N_2877,N_3705);
nor UO_553 (O_553,N_4863,N_4011);
nor UO_554 (O_554,N_3489,N_3351);
and UO_555 (O_555,N_3490,N_4408);
or UO_556 (O_556,N_3680,N_3242);
or UO_557 (O_557,N_2684,N_3184);
nand UO_558 (O_558,N_4870,N_2698);
or UO_559 (O_559,N_3076,N_3786);
nor UO_560 (O_560,N_4216,N_4226);
and UO_561 (O_561,N_4581,N_2807);
and UO_562 (O_562,N_3760,N_4708);
nand UO_563 (O_563,N_3596,N_4900);
or UO_564 (O_564,N_4173,N_4158);
nor UO_565 (O_565,N_4229,N_4648);
nor UO_566 (O_566,N_2899,N_3261);
and UO_567 (O_567,N_4896,N_2933);
nor UO_568 (O_568,N_3421,N_3407);
nand UO_569 (O_569,N_3492,N_3389);
nor UO_570 (O_570,N_3197,N_4729);
nand UO_571 (O_571,N_2987,N_3859);
nor UO_572 (O_572,N_2709,N_4551);
or UO_573 (O_573,N_4578,N_2996);
nor UO_574 (O_574,N_3625,N_3109);
or UO_575 (O_575,N_2706,N_4676);
or UO_576 (O_576,N_3976,N_4392);
nor UO_577 (O_577,N_2823,N_4480);
nand UO_578 (O_578,N_4448,N_3303);
and UO_579 (O_579,N_4309,N_4675);
nor UO_580 (O_580,N_3010,N_4267);
nor UO_581 (O_581,N_2926,N_3342);
nand UO_582 (O_582,N_4455,N_2887);
nand UO_583 (O_583,N_2590,N_3355);
nand UO_584 (O_584,N_4868,N_4301);
or UO_585 (O_585,N_4009,N_3003);
and UO_586 (O_586,N_3277,N_2662);
or UO_587 (O_587,N_3753,N_3085);
or UO_588 (O_588,N_2570,N_2980);
nand UO_589 (O_589,N_3216,N_3744);
and UO_590 (O_590,N_4538,N_4438);
nor UO_591 (O_591,N_2974,N_3403);
nand UO_592 (O_592,N_3360,N_3487);
nand UO_593 (O_593,N_4445,N_2587);
nand UO_594 (O_594,N_2994,N_3947);
and UO_595 (O_595,N_3829,N_4450);
and UO_596 (O_596,N_4500,N_3333);
or UO_597 (O_597,N_2856,N_4218);
or UO_598 (O_598,N_3994,N_3239);
nand UO_599 (O_599,N_4205,N_3568);
or UO_600 (O_600,N_2562,N_4555);
nand UO_601 (O_601,N_4666,N_3672);
or UO_602 (O_602,N_2578,N_4212);
and UO_603 (O_603,N_2959,N_3724);
or UO_604 (O_604,N_4095,N_3123);
and UO_605 (O_605,N_4615,N_3252);
nor UO_606 (O_606,N_3685,N_2512);
nand UO_607 (O_607,N_3683,N_2767);
nor UO_608 (O_608,N_4641,N_2676);
nor UO_609 (O_609,N_3655,N_4388);
or UO_610 (O_610,N_3457,N_3463);
nand UO_611 (O_611,N_2708,N_4596);
nor UO_612 (O_612,N_4363,N_3835);
and UO_613 (O_613,N_3918,N_3623);
or UO_614 (O_614,N_4119,N_3437);
xnor UO_615 (O_615,N_4244,N_2947);
nand UO_616 (O_616,N_4148,N_2524);
nor UO_617 (O_617,N_4918,N_4836);
and UO_618 (O_618,N_3147,N_2553);
and UO_619 (O_619,N_4856,N_3051);
and UO_620 (O_620,N_4444,N_4166);
nand UO_621 (O_621,N_3839,N_3456);
or UO_622 (O_622,N_4743,N_3289);
nor UO_623 (O_623,N_2572,N_3535);
nand UO_624 (O_624,N_4296,N_4243);
and UO_625 (O_625,N_3175,N_4385);
xor UO_626 (O_626,N_3371,N_3926);
nand UO_627 (O_627,N_4077,N_3301);
nor UO_628 (O_628,N_3029,N_2673);
or UO_629 (O_629,N_4024,N_2518);
or UO_630 (O_630,N_3482,N_2780);
nor UO_631 (O_631,N_3652,N_2628);
or UO_632 (O_632,N_4903,N_4761);
and UO_633 (O_633,N_4403,N_4885);
and UO_634 (O_634,N_3598,N_3690);
and UO_635 (O_635,N_4263,N_4948);
and UO_636 (O_636,N_2779,N_3444);
or UO_637 (O_637,N_3718,N_3210);
and UO_638 (O_638,N_3181,N_2538);
or UO_639 (O_639,N_3284,N_3542);
nor UO_640 (O_640,N_4342,N_4670);
or UO_641 (O_641,N_3330,N_4979);
nand UO_642 (O_642,N_4976,N_3356);
nor UO_643 (O_643,N_4730,N_3494);
and UO_644 (O_644,N_4184,N_2969);
nor UO_645 (O_645,N_4523,N_3416);
nand UO_646 (O_646,N_2711,N_2502);
nor UO_647 (O_647,N_2912,N_3315);
and UO_648 (O_648,N_4995,N_3308);
nand UO_649 (O_649,N_4846,N_2758);
or UO_650 (O_650,N_4872,N_3854);
nor UO_651 (O_651,N_3939,N_2759);
and UO_652 (O_652,N_4806,N_3138);
nand UO_653 (O_653,N_3036,N_4531);
nand UO_654 (O_654,N_3622,N_3189);
or UO_655 (O_655,N_3664,N_2583);
and UO_656 (O_656,N_4524,N_3117);
nor UO_657 (O_657,N_2695,N_4969);
nand UO_658 (O_658,N_3423,N_3106);
nor UO_659 (O_659,N_3678,N_3946);
nand UO_660 (O_660,N_3442,N_3462);
nor UO_661 (O_661,N_2722,N_4984);
nand UO_662 (O_662,N_4815,N_3335);
nor UO_663 (O_663,N_3896,N_3576);
xor UO_664 (O_664,N_2547,N_3021);
nor UO_665 (O_665,N_3856,N_3698);
nor UO_666 (O_666,N_4134,N_4072);
nor UO_667 (O_667,N_3735,N_3884);
and UO_668 (O_668,N_3414,N_3391);
and UO_669 (O_669,N_4096,N_3165);
and UO_670 (O_670,N_2510,N_2704);
or UO_671 (O_671,N_3111,N_3920);
nand UO_672 (O_672,N_4536,N_4258);
nand UO_673 (O_673,N_3783,N_4241);
nor UO_674 (O_674,N_4924,N_4285);
or UO_675 (O_675,N_3993,N_2674);
or UO_676 (O_676,N_4864,N_4487);
or UO_677 (O_677,N_3876,N_2792);
xor UO_678 (O_678,N_4876,N_3798);
nand UO_679 (O_679,N_3750,N_4952);
nor UO_680 (O_680,N_3103,N_3179);
nand UO_681 (O_681,N_4936,N_3470);
nand UO_682 (O_682,N_3620,N_4680);
or UO_683 (O_683,N_4060,N_4797);
nand UO_684 (O_684,N_3996,N_2844);
and UO_685 (O_685,N_4826,N_4765);
or UO_686 (O_686,N_3953,N_4677);
xor UO_687 (O_687,N_2600,N_4791);
or UO_688 (O_688,N_2689,N_4558);
and UO_689 (O_689,N_3505,N_3826);
or UO_690 (O_690,N_4364,N_3035);
xnor UO_691 (O_691,N_4576,N_2613);
nand UO_692 (O_692,N_2642,N_4270);
or UO_693 (O_693,N_4509,N_3212);
nor UO_694 (O_694,N_4379,N_3196);
or UO_695 (O_695,N_4102,N_3345);
and UO_696 (O_696,N_2731,N_2707);
and UO_697 (O_697,N_4767,N_4598);
and UO_698 (O_698,N_3513,N_3503);
and UO_699 (O_699,N_4269,N_4121);
xnor UO_700 (O_700,N_3069,N_4144);
and UO_701 (O_701,N_2660,N_2829);
nor UO_702 (O_702,N_4916,N_4721);
and UO_703 (O_703,N_4099,N_4020);
nor UO_704 (O_704,N_3693,N_4254);
or UO_705 (O_705,N_4307,N_4835);
nand UO_706 (O_706,N_2516,N_3883);
nor UO_707 (O_707,N_3049,N_2548);
nor UO_708 (O_708,N_4023,N_4961);
nor UO_709 (O_709,N_3133,N_3608);
xnor UO_710 (O_710,N_3911,N_4327);
or UO_711 (O_711,N_3208,N_2893);
nand UO_712 (O_712,N_3987,N_3677);
and UO_713 (O_713,N_4898,N_3755);
nand UO_714 (O_714,N_2738,N_4645);
or UO_715 (O_715,N_3475,N_3093);
or UO_716 (O_716,N_2874,N_4154);
xnor UO_717 (O_717,N_3521,N_3431);
and UO_718 (O_718,N_4481,N_3240);
nand UO_719 (O_719,N_3169,N_3869);
or UO_720 (O_720,N_4004,N_3817);
and UO_721 (O_721,N_4010,N_3991);
or UO_722 (O_722,N_3375,N_4800);
nand UO_723 (O_723,N_4819,N_2891);
and UO_724 (O_724,N_4699,N_4907);
or UO_725 (O_725,N_3077,N_4811);
nand UO_726 (O_726,N_4790,N_4988);
nand UO_727 (O_727,N_4014,N_3113);
and UO_728 (O_728,N_4407,N_4286);
or UO_729 (O_729,N_4174,N_3882);
nand UO_730 (O_730,N_3466,N_3180);
nor UO_731 (O_731,N_2544,N_4624);
nor UO_732 (O_732,N_4696,N_2546);
nand UO_733 (O_733,N_2836,N_2566);
nand UO_734 (O_734,N_3445,N_4175);
or UO_735 (O_735,N_3893,N_4673);
nand UO_736 (O_736,N_4639,N_3757);
nor UO_737 (O_737,N_3201,N_3816);
or UO_738 (O_738,N_3435,N_3440);
nor UO_739 (O_739,N_4042,N_4331);
nand UO_740 (O_740,N_3533,N_3522);
nor UO_741 (O_741,N_3383,N_3149);
or UO_742 (O_742,N_2688,N_4468);
or UO_743 (O_743,N_4446,N_3155);
xnor UO_744 (O_744,N_4973,N_3032);
nor UO_745 (O_745,N_2834,N_3687);
nand UO_746 (O_746,N_3815,N_3566);
and UO_747 (O_747,N_3984,N_4026);
nand UO_748 (O_748,N_3803,N_2735);
or UO_749 (O_749,N_3254,N_3862);
nand UO_750 (O_750,N_4692,N_4220);
nor UO_751 (O_751,N_3245,N_3556);
or UO_752 (O_752,N_3574,N_3202);
or UO_753 (O_753,N_3006,N_3102);
xnor UO_754 (O_754,N_4990,N_3830);
nor UO_755 (O_755,N_3011,N_2531);
nor UO_756 (O_756,N_4957,N_3967);
or UO_757 (O_757,N_3825,N_2624);
or UO_758 (O_758,N_3091,N_2741);
or UO_759 (O_759,N_2971,N_3396);
nand UO_760 (O_760,N_3633,N_4322);
nand UO_761 (O_761,N_3785,N_2963);
nor UO_762 (O_762,N_4048,N_4186);
xnor UO_763 (O_763,N_2774,N_3483);
and UO_764 (O_764,N_2810,N_2944);
nand UO_765 (O_765,N_2817,N_3959);
nand UO_766 (O_766,N_4150,N_2965);
xnor UO_767 (O_767,N_4687,N_3019);
nor UO_768 (O_768,N_4146,N_2749);
and UO_769 (O_769,N_2527,N_4410);
and UO_770 (O_770,N_4951,N_3864);
nand UO_771 (O_771,N_2827,N_4113);
or UO_772 (O_772,N_3262,N_2765);
nand UO_773 (O_773,N_3132,N_4160);
nor UO_774 (O_774,N_3141,N_2889);
and UO_775 (O_775,N_3127,N_3943);
nor UO_776 (O_776,N_2859,N_3114);
nand UO_777 (O_777,N_4195,N_3778);
or UO_778 (O_778,N_3931,N_4033);
nor UO_779 (O_779,N_2691,N_4759);
and UO_780 (O_780,N_4170,N_3809);
and UO_781 (O_781,N_4311,N_3960);
and UO_782 (O_782,N_3606,N_4693);
or UO_783 (O_783,N_3643,N_3894);
and UO_784 (O_784,N_3312,N_2888);
nor UO_785 (O_785,N_4543,N_3992);
nand UO_786 (O_786,N_3276,N_3178);
nand UO_787 (O_787,N_3163,N_3878);
xnor UO_788 (O_788,N_3244,N_2862);
and UO_789 (O_789,N_4398,N_4880);
and UO_790 (O_790,N_4934,N_3597);
or UO_791 (O_791,N_3046,N_2825);
nand UO_792 (O_792,N_3588,N_4116);
nor UO_793 (O_793,N_4128,N_4053);
nor UO_794 (O_794,N_4406,N_2852);
nor UO_795 (O_795,N_3800,N_3554);
or UO_796 (O_796,N_4956,N_3605);
or UO_797 (O_797,N_3198,N_2900);
nor UO_798 (O_798,N_4689,N_3791);
nor UO_799 (O_799,N_3982,N_3156);
and UO_800 (O_800,N_4807,N_2594);
and UO_801 (O_801,N_4515,N_4454);
or UO_802 (O_802,N_4329,N_3327);
xor UO_803 (O_803,N_4283,N_2641);
and UO_804 (O_804,N_2726,N_3640);
nand UO_805 (O_805,N_4873,N_3637);
xnor UO_806 (O_806,N_2853,N_2576);
or UO_807 (O_807,N_4298,N_3581);
or UO_808 (O_808,N_4923,N_4669);
nor UO_809 (O_809,N_4865,N_4694);
nor UO_810 (O_810,N_3736,N_4155);
nor UO_811 (O_811,N_2921,N_3280);
or UO_812 (O_812,N_3015,N_3182);
or UO_813 (O_813,N_3836,N_4894);
or UO_814 (O_814,N_4616,N_4685);
nand UO_815 (O_815,N_3222,N_2796);
and UO_816 (O_816,N_3265,N_3186);
nand UO_817 (O_817,N_3656,N_3128);
xor UO_818 (O_818,N_3143,N_3930);
or UO_819 (O_819,N_2910,N_4529);
and UO_820 (O_820,N_3057,N_4792);
and UO_821 (O_821,N_4357,N_4367);
nand UO_822 (O_822,N_4803,N_4917);
xnor UO_823 (O_823,N_2752,N_4493);
and UO_824 (O_824,N_2593,N_4440);
nand UO_825 (O_825,N_4549,N_3332);
and UO_826 (O_826,N_4179,N_3418);
and UO_827 (O_827,N_2682,N_3158);
nor UO_828 (O_828,N_3774,N_3963);
or UO_829 (O_829,N_3388,N_4372);
nand UO_830 (O_830,N_4760,N_2992);
and UO_831 (O_831,N_3467,N_4715);
nor UO_832 (O_832,N_4091,N_3500);
nor UO_833 (O_833,N_3098,N_3454);
or UO_834 (O_834,N_4688,N_4553);
or UO_835 (O_835,N_4290,N_3564);
or UO_836 (O_836,N_3710,N_3232);
or UO_837 (O_837,N_4087,N_3759);
nor UO_838 (O_838,N_3446,N_4061);
nand UO_839 (O_839,N_2894,N_2949);
nand UO_840 (O_840,N_2542,N_3455);
nor UO_841 (O_841,N_4844,N_4652);
or UO_842 (O_842,N_3427,N_2885);
nor UO_843 (O_843,N_2720,N_3362);
or UO_844 (O_844,N_4723,N_2606);
or UO_845 (O_845,N_3000,N_3429);
and UO_846 (O_846,N_2507,N_3725);
nand UO_847 (O_847,N_3592,N_4377);
or UO_848 (O_848,N_3737,N_3756);
and UO_849 (O_849,N_3270,N_3174);
nand UO_850 (O_850,N_3796,N_4921);
nand UO_851 (O_851,N_2993,N_2612);
nand UO_852 (O_852,N_3910,N_4939);
nor UO_853 (O_853,N_2868,N_3307);
nand UO_854 (O_854,N_3037,N_3075);
or UO_855 (O_855,N_2816,N_4482);
xor UO_856 (O_856,N_3613,N_4813);
nand UO_857 (O_857,N_3340,N_4447);
xnor UO_858 (O_858,N_4814,N_3168);
nand UO_859 (O_859,N_2533,N_4358);
or UO_860 (O_860,N_4300,N_4548);
or UO_861 (O_861,N_3916,N_3205);
nor UO_862 (O_862,N_4672,N_3083);
and UO_863 (O_863,N_2787,N_3476);
nand UO_864 (O_864,N_3834,N_3644);
nand UO_865 (O_865,N_4659,N_2777);
nor UO_866 (O_866,N_4442,N_3352);
nor UO_867 (O_867,N_3290,N_4330);
or UO_868 (O_868,N_4142,N_4360);
or UO_869 (O_869,N_3314,N_3405);
nor UO_870 (O_870,N_4299,N_3579);
and UO_871 (O_871,N_2864,N_4324);
and UO_872 (O_872,N_2519,N_4439);
or UO_873 (O_873,N_3285,N_2763);
and UO_874 (O_874,N_3805,N_4247);
nor UO_875 (O_875,N_3749,N_4530);
nand UO_876 (O_876,N_3428,N_3488);
or UO_877 (O_877,N_3410,N_4347);
nand UO_878 (O_878,N_4250,N_2595);
nor UO_879 (O_879,N_3234,N_3932);
and UO_880 (O_880,N_2525,N_4075);
nor UO_881 (O_881,N_4539,N_3663);
xor UO_882 (O_882,N_3563,N_4275);
nor UO_883 (O_883,N_3923,N_3970);
nand UO_884 (O_884,N_2898,N_4022);
nor UO_885 (O_885,N_3525,N_2968);
or UO_886 (O_886,N_3768,N_2878);
nor UO_887 (O_887,N_4093,N_2999);
nor UO_888 (O_888,N_4320,N_3957);
or UO_889 (O_889,N_3917,N_4209);
nand UO_890 (O_890,N_4851,N_4577);
or UO_891 (O_891,N_3904,N_3341);
or UO_892 (O_892,N_3166,N_4318);
or UO_893 (O_893,N_4253,N_4679);
and UO_894 (O_894,N_4238,N_2699);
and UO_895 (O_895,N_3030,N_3367);
or UO_896 (O_896,N_3331,N_3561);
and UO_897 (O_897,N_3060,N_4698);
nand UO_898 (O_898,N_4496,N_4256);
and UO_899 (O_899,N_3529,N_4464);
nand UO_900 (O_900,N_3191,N_4545);
nor UO_901 (O_901,N_4462,N_4777);
or UO_902 (O_902,N_3121,N_4682);
nor UO_903 (O_903,N_4941,N_4980);
nor UO_904 (O_904,N_4594,N_3257);
or UO_905 (O_905,N_2677,N_3034);
or UO_906 (O_906,N_2863,N_3195);
and UO_907 (O_907,N_3955,N_3837);
or UO_908 (O_908,N_2789,N_3849);
nand UO_909 (O_909,N_3119,N_3999);
nand UO_910 (O_910,N_2962,N_3199);
and UO_911 (O_911,N_4773,N_4394);
or UO_912 (O_912,N_4038,N_4393);
or UO_913 (O_913,N_3364,N_3730);
nand UO_914 (O_914,N_4222,N_3420);
or UO_915 (O_915,N_4747,N_2521);
and UO_916 (O_916,N_3088,N_3002);
and UO_917 (O_917,N_2713,N_2879);
nor UO_918 (O_918,N_3089,N_4998);
nor UO_919 (O_919,N_3954,N_4149);
and UO_920 (O_920,N_2800,N_4746);
and UO_921 (O_921,N_4845,N_4409);
nor UO_922 (O_922,N_4242,N_4716);
nor UO_923 (O_923,N_3879,N_2945);
nand UO_924 (O_924,N_3937,N_3144);
nor UO_925 (O_925,N_4820,N_3651);
or UO_926 (O_926,N_3853,N_3172);
nand UO_927 (O_927,N_4793,N_3048);
nor UO_928 (O_928,N_3224,N_4277);
nor UO_929 (O_929,N_4963,N_3951);
nor UO_930 (O_930,N_3220,N_2976);
nand UO_931 (O_931,N_2901,N_3599);
nor UO_932 (O_932,N_4569,N_3682);
nand UO_933 (O_933,N_4278,N_4710);
nor UO_934 (O_934,N_4665,N_2873);
or UO_935 (O_935,N_2757,N_4156);
nor UO_936 (O_936,N_3720,N_3058);
nor UO_937 (O_937,N_2797,N_4297);
and UO_938 (O_938,N_2526,N_3337);
and UO_939 (O_939,N_4337,N_3066);
nand UO_940 (O_940,N_3295,N_3840);
and UO_941 (O_941,N_4940,N_4804);
nor UO_942 (O_942,N_4387,N_3316);
nor UO_943 (O_943,N_4034,N_4664);
or UO_944 (O_944,N_3399,N_3901);
and UO_945 (O_945,N_3775,N_3204);
nand UO_946 (O_946,N_3325,N_4203);
nor UO_947 (O_947,N_4180,N_2775);
xor UO_948 (O_948,N_4153,N_3281);
nor UO_949 (O_949,N_3641,N_2838);
nor UO_950 (O_950,N_4460,N_4781);
nand UO_951 (O_951,N_2715,N_2890);
nor UO_952 (O_952,N_4823,N_3392);
or UO_953 (O_953,N_3390,N_4505);
nand UO_954 (O_954,N_3016,N_4559);
nor UO_955 (O_955,N_4511,N_3095);
nand UO_956 (O_956,N_2575,N_4319);
and UO_957 (O_957,N_3292,N_2657);
and UO_958 (O_958,N_4799,N_3096);
nand UO_959 (O_959,N_4560,N_3532);
and UO_960 (O_960,N_2818,N_2754);
nand UO_961 (O_961,N_4321,N_3850);
and UO_962 (O_962,N_3221,N_3822);
or UO_963 (O_963,N_3072,N_2880);
nor UO_964 (O_964,N_4834,N_3832);
or UO_965 (O_965,N_4194,N_4031);
nor UO_966 (O_966,N_4255,N_4822);
nand UO_967 (O_967,N_3305,N_3313);
or UO_968 (O_968,N_2892,N_2865);
and UO_969 (O_969,N_2739,N_4341);
nand UO_970 (O_970,N_3408,N_3226);
or UO_971 (O_971,N_4428,N_3697);
nor UO_972 (O_972,N_2585,N_3990);
nor UO_973 (O_973,N_4966,N_3674);
and UO_974 (O_974,N_3105,N_4502);
and UO_975 (O_975,N_4871,N_3551);
nand UO_976 (O_976,N_4378,N_2985);
nand UO_977 (O_977,N_3547,N_4052);
nand UO_978 (O_978,N_4475,N_4129);
nand UO_979 (O_979,N_3793,N_4465);
and UO_980 (O_980,N_4801,N_4436);
nand UO_981 (O_981,N_4485,N_3938);
nand UO_982 (O_982,N_4044,N_3317);
nand UO_983 (O_983,N_3452,N_4849);
and UO_984 (O_984,N_4608,N_4178);
nor UO_985 (O_985,N_4739,N_3304);
nor UO_986 (O_986,N_3142,N_3614);
xnor UO_987 (O_987,N_3152,N_4074);
and UO_988 (O_988,N_3344,N_4181);
nor UO_989 (O_989,N_2961,N_4499);
nand UO_990 (O_990,N_4561,N_3686);
or UO_991 (O_991,N_2849,N_3565);
and UO_992 (O_992,N_3122,N_4214);
xnor UO_993 (O_993,N_2619,N_4971);
or UO_994 (O_994,N_4157,N_2867);
or UO_995 (O_995,N_4550,N_4818);
nor UO_996 (O_996,N_4878,N_3339);
or UO_997 (O_997,N_3941,N_2847);
nor UO_998 (O_998,N_3769,N_4497);
or UO_999 (O_999,N_3460,N_2990);
endmodule