module basic_1000_10000_1500_2_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5001,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5019,N_5021,N_5022,N_5025,N_5028,N_5030,N_5035,N_5036,N_5039,N_5041,N_5043,N_5044,N_5045,N_5046,N_5050,N_5051,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5061,N_5062,N_5065,N_5067,N_5070,N_5071,N_5072,N_5075,N_5076,N_5078,N_5080,N_5081,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5097,N_5102,N_5105,N_5106,N_5107,N_5108,N_5110,N_5111,N_5112,N_5113,N_5117,N_5118,N_5119,N_5120,N_5121,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5138,N_5139,N_5140,N_5142,N_5143,N_5144,N_5145,N_5147,N_5148,N_5150,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5159,N_5160,N_5163,N_5164,N_5166,N_5169,N_5170,N_5171,N_5173,N_5175,N_5177,N_5179,N_5180,N_5181,N_5184,N_5187,N_5188,N_5190,N_5192,N_5193,N_5195,N_5196,N_5198,N_5200,N_5201,N_5202,N_5204,N_5205,N_5207,N_5212,N_5214,N_5216,N_5217,N_5218,N_5220,N_5221,N_5222,N_5223,N_5225,N_5226,N_5230,N_5231,N_5237,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5246,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5258,N_5261,N_5262,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5274,N_5276,N_5278,N_5279,N_5281,N_5284,N_5285,N_5286,N_5289,N_5290,N_5291,N_5293,N_5295,N_5296,N_5297,N_5299,N_5300,N_5302,N_5304,N_5306,N_5307,N_5309,N_5312,N_5314,N_5315,N_5317,N_5319,N_5320,N_5321,N_5324,N_5325,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5334,N_5335,N_5340,N_5343,N_5345,N_5348,N_5349,N_5354,N_5357,N_5358,N_5360,N_5361,N_5362,N_5363,N_5365,N_5366,N_5367,N_5371,N_5372,N_5374,N_5375,N_5376,N_5377,N_5379,N_5382,N_5385,N_5386,N_5390,N_5391,N_5392,N_5394,N_5395,N_5397,N_5399,N_5400,N_5401,N_5402,N_5403,N_5405,N_5409,N_5412,N_5415,N_5416,N_5417,N_5418,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5427,N_5430,N_5431,N_5432,N_5435,N_5437,N_5438,N_5439,N_5442,N_5443,N_5444,N_5445,N_5448,N_5454,N_5455,N_5457,N_5458,N_5459,N_5462,N_5466,N_5467,N_5468,N_5469,N_5470,N_5472,N_5476,N_5477,N_5479,N_5482,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5493,N_5495,N_5502,N_5504,N_5505,N_5506,N_5508,N_5512,N_5515,N_5518,N_5519,N_5521,N_5522,N_5524,N_5526,N_5527,N_5528,N_5529,N_5531,N_5532,N_5534,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5544,N_5545,N_5546,N_5547,N_5549,N_5550,N_5552,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5561,N_5563,N_5565,N_5568,N_5569,N_5570,N_5571,N_5573,N_5576,N_5577,N_5581,N_5582,N_5583,N_5585,N_5587,N_5589,N_5591,N_5592,N_5593,N_5594,N_5597,N_5600,N_5601,N_5602,N_5603,N_5608,N_5610,N_5611,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5621,N_5622,N_5624,N_5625,N_5627,N_5629,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5646,N_5647,N_5648,N_5652,N_5653,N_5657,N_5659,N_5661,N_5663,N_5666,N_5668,N_5670,N_5671,N_5672,N_5676,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5705,N_5707,N_5709,N_5710,N_5712,N_5714,N_5715,N_5716,N_5718,N_5719,N_5720,N_5721,N_5724,N_5726,N_5727,N_5728,N_5729,N_5731,N_5733,N_5735,N_5736,N_5741,N_5743,N_5746,N_5747,N_5749,N_5752,N_5753,N_5754,N_5756,N_5759,N_5766,N_5768,N_5769,N_5772,N_5773,N_5774,N_5775,N_5777,N_5778,N_5779,N_5782,N_5783,N_5786,N_5787,N_5789,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5804,N_5806,N_5807,N_5808,N_5810,N_5811,N_5812,N_5815,N_5816,N_5817,N_5818,N_5819,N_5821,N_5824,N_5828,N_5829,N_5830,N_5834,N_5835,N_5836,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5847,N_5850,N_5852,N_5853,N_5855,N_5856,N_5859,N_5860,N_5861,N_5863,N_5868,N_5870,N_5873,N_5874,N_5875,N_5876,N_5880,N_5883,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5892,N_5893,N_5894,N_5895,N_5898,N_5900,N_5901,N_5903,N_5905,N_5906,N_5907,N_5910,N_5916,N_5917,N_5918,N_5920,N_5921,N_5923,N_5925,N_5926,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5939,N_5940,N_5942,N_5943,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5953,N_5954,N_5956,N_5957,N_5959,N_5967,N_5969,N_5972,N_5973,N_5974,N_5975,N_5976,N_5979,N_5982,N_5983,N_5984,N_5986,N_5988,N_5992,N_5993,N_5994,N_5996,N_5997,N_5999,N_6002,N_6005,N_6010,N_6011,N_6012,N_6013,N_6017,N_6018,N_6020,N_6021,N_6022,N_6023,N_6025,N_6027,N_6028,N_6029,N_6030,N_6033,N_6035,N_6036,N_6037,N_6038,N_6040,N_6041,N_6042,N_6043,N_6045,N_6048,N_6050,N_6051,N_6052,N_6053,N_6054,N_6057,N_6058,N_6060,N_6061,N_6062,N_6063,N_6065,N_6067,N_6069,N_6073,N_6074,N_6076,N_6077,N_6080,N_6081,N_6083,N_6085,N_6086,N_6087,N_6088,N_6089,N_6091,N_6092,N_6093,N_6094,N_6095,N_6097,N_6098,N_6100,N_6102,N_6105,N_6106,N_6108,N_6109,N_6110,N_6111,N_6113,N_6115,N_6116,N_6118,N_6120,N_6121,N_6123,N_6125,N_6126,N_6128,N_6129,N_6131,N_6132,N_6133,N_6134,N_6135,N_6139,N_6140,N_6143,N_6145,N_6146,N_6148,N_6149,N_6151,N_6152,N_6154,N_6156,N_6159,N_6160,N_6161,N_6164,N_6165,N_6167,N_6168,N_6169,N_6170,N_6172,N_6174,N_6176,N_6177,N_6180,N_6182,N_6183,N_6185,N_6188,N_6190,N_6192,N_6194,N_6200,N_6203,N_6204,N_6205,N_6207,N_6208,N_6209,N_6210,N_6213,N_6214,N_6215,N_6216,N_6217,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6226,N_6227,N_6230,N_6231,N_6232,N_6233,N_6235,N_6237,N_6238,N_6241,N_6244,N_6245,N_6248,N_6249,N_6250,N_6251,N_6253,N_6257,N_6259,N_6262,N_6263,N_6264,N_6267,N_6268,N_6269,N_6271,N_6272,N_6274,N_6275,N_6278,N_6279,N_6284,N_6285,N_6286,N_6287,N_6290,N_6292,N_6293,N_6294,N_6296,N_6297,N_6298,N_6300,N_6302,N_6304,N_6305,N_6307,N_6309,N_6310,N_6313,N_6315,N_6316,N_6319,N_6320,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6335,N_6336,N_6338,N_6340,N_6341,N_6342,N_6345,N_6346,N_6347,N_6348,N_6349,N_6352,N_6353,N_6354,N_6355,N_6359,N_6361,N_6362,N_6363,N_6367,N_6368,N_6369,N_6370,N_6372,N_6373,N_6374,N_6376,N_6377,N_6378,N_6380,N_6381,N_6382,N_6384,N_6385,N_6386,N_6388,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6401,N_6402,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6412,N_6414,N_6416,N_6419,N_6421,N_6422,N_6423,N_6425,N_6426,N_6427,N_6429,N_6430,N_6432,N_6434,N_6435,N_6436,N_6438,N_6441,N_6442,N_6443,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6457,N_6459,N_6461,N_6462,N_6463,N_6464,N_6466,N_6468,N_6470,N_6471,N_6472,N_6475,N_6479,N_6480,N_6481,N_6482,N_6483,N_6486,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6498,N_6499,N_6504,N_6506,N_6507,N_6508,N_6510,N_6512,N_6513,N_6516,N_6517,N_6519,N_6520,N_6521,N_6525,N_6526,N_6528,N_6529,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6545,N_6547,N_6550,N_6551,N_6554,N_6555,N_6557,N_6558,N_6560,N_6561,N_6562,N_6563,N_6564,N_6570,N_6571,N_6572,N_6573,N_6574,N_6578,N_6579,N_6580,N_6583,N_6584,N_6585,N_6586,N_6588,N_6589,N_6591,N_6592,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6614,N_6615,N_6620,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6631,N_6633,N_6634,N_6638,N_6639,N_6640,N_6641,N_6643,N_6645,N_6647,N_6657,N_6658,N_6659,N_6662,N_6665,N_6666,N_6667,N_6668,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6684,N_6685,N_6686,N_6688,N_6690,N_6691,N_6694,N_6695,N_6698,N_6699,N_6700,N_6702,N_6707,N_6708,N_6709,N_6712,N_6713,N_6714,N_6715,N_6718,N_6721,N_6723,N_6724,N_6725,N_6727,N_6729,N_6730,N_6733,N_6740,N_6741,N_6742,N_6743,N_6745,N_6748,N_6749,N_6750,N_6752,N_6753,N_6755,N_6756,N_6757,N_6758,N_6760,N_6763,N_6764,N_6765,N_6766,N_6768,N_6770,N_6773,N_6774,N_6776,N_6777,N_6781,N_6782,N_6783,N_6784,N_6785,N_6787,N_6788,N_6789,N_6792,N_6793,N_6795,N_6797,N_6798,N_6799,N_6800,N_6802,N_6803,N_6804,N_6807,N_6808,N_6809,N_6810,N_6812,N_6813,N_6814,N_6816,N_6817,N_6819,N_6821,N_6822,N_6826,N_6834,N_6836,N_6838,N_6839,N_6841,N_6844,N_6845,N_6847,N_6849,N_6850,N_6853,N_6854,N_6856,N_6861,N_6862,N_6863,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6875,N_6876,N_6877,N_6879,N_6880,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6890,N_6894,N_6895,N_6896,N_6898,N_6899,N_6903,N_6905,N_6906,N_6907,N_6909,N_6910,N_6911,N_6912,N_6915,N_6916,N_6917,N_6920,N_6921,N_6922,N_6923,N_6927,N_6929,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6951,N_6952,N_6956,N_6958,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6970,N_6972,N_6974,N_6975,N_6980,N_6983,N_6984,N_6985,N_6987,N_6988,N_6989,N_6990,N_6993,N_6996,N_7000,N_7002,N_7003,N_7006,N_7008,N_7009,N_7012,N_7013,N_7016,N_7018,N_7019,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7029,N_7030,N_7031,N_7034,N_7035,N_7037,N_7038,N_7040,N_7042,N_7044,N_7046,N_7047,N_7049,N_7050,N_7052,N_7054,N_7055,N_7057,N_7059,N_7062,N_7063,N_7064,N_7066,N_7067,N_7068,N_7069,N_7070,N_7072,N_7073,N_7076,N_7077,N_7078,N_7079,N_7080,N_7082,N_7084,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7097,N_7098,N_7101,N_7102,N_7104,N_7105,N_7111,N_7112,N_7114,N_7120,N_7121,N_7122,N_7123,N_7125,N_7126,N_7127,N_7128,N_7130,N_7131,N_7135,N_7136,N_7137,N_7142,N_7143,N_7145,N_7146,N_7147,N_7148,N_7150,N_7151,N_7152,N_7153,N_7157,N_7158,N_7160,N_7165,N_7166,N_7172,N_7178,N_7181,N_7182,N_7183,N_7184,N_7185,N_7187,N_7189,N_7192,N_7199,N_7200,N_7202,N_7204,N_7206,N_7207,N_7208,N_7211,N_7212,N_7213,N_7214,N_7215,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7225,N_7226,N_7229,N_7230,N_7231,N_7232,N_7233,N_7238,N_7239,N_7240,N_7241,N_7247,N_7248,N_7249,N_7250,N_7251,N_7253,N_7254,N_7260,N_7261,N_7262,N_7264,N_7266,N_7269,N_7271,N_7272,N_7273,N_7274,N_7276,N_7277,N_7278,N_7280,N_7282,N_7283,N_7284,N_7285,N_7288,N_7289,N_7290,N_7293,N_7294,N_7295,N_7296,N_7297,N_7300,N_7301,N_7303,N_7304,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7326,N_7329,N_7331,N_7332,N_7334,N_7335,N_7336,N_7337,N_7339,N_7340,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7349,N_7350,N_7352,N_7355,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7367,N_7368,N_7371,N_7372,N_7375,N_7378,N_7380,N_7383,N_7384,N_7385,N_7386,N_7388,N_7390,N_7392,N_7395,N_7398,N_7402,N_7403,N_7404,N_7405,N_7406,N_7408,N_7411,N_7412,N_7414,N_7416,N_7417,N_7418,N_7419,N_7421,N_7424,N_7427,N_7429,N_7430,N_7433,N_7434,N_7435,N_7438,N_7439,N_7440,N_7441,N_7446,N_7448,N_7450,N_7451,N_7452,N_7454,N_7459,N_7461,N_7463,N_7465,N_7466,N_7468,N_7472,N_7473,N_7474,N_7475,N_7476,N_7479,N_7481,N_7483,N_7485,N_7488,N_7489,N_7490,N_7491,N_7492,N_7494,N_7495,N_7498,N_7499,N_7500,N_7502,N_7505,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7515,N_7516,N_7518,N_7519,N_7522,N_7524,N_7527,N_7528,N_7530,N_7531,N_7532,N_7533,N_7535,N_7536,N_7537,N_7538,N_7539,N_7543,N_7544,N_7546,N_7550,N_7551,N_7553,N_7554,N_7555,N_7556,N_7559,N_7560,N_7561,N_7562,N_7564,N_7565,N_7566,N_7567,N_7568,N_7570,N_7571,N_7572,N_7575,N_7576,N_7577,N_7581,N_7584,N_7585,N_7586,N_7587,N_7588,N_7590,N_7592,N_7593,N_7594,N_7596,N_7597,N_7598,N_7603,N_7606,N_7607,N_7608,N_7613,N_7614,N_7615,N_7619,N_7620,N_7623,N_7624,N_7626,N_7629,N_7630,N_7633,N_7635,N_7636,N_7637,N_7638,N_7642,N_7643,N_7645,N_7646,N_7647,N_7651,N_7652,N_7653,N_7654,N_7655,N_7657,N_7658,N_7661,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7672,N_7673,N_7674,N_7677,N_7678,N_7680,N_7681,N_7683,N_7685,N_7686,N_7690,N_7692,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7702,N_7703,N_7704,N_7705,N_7707,N_7709,N_7711,N_7714,N_7715,N_7716,N_7717,N_7718,N_7720,N_7721,N_7722,N_7723,N_7726,N_7728,N_7729,N_7730,N_7732,N_7733,N_7734,N_7735,N_7736,N_7738,N_7743,N_7745,N_7747,N_7748,N_7750,N_7752,N_7753,N_7754,N_7755,N_7756,N_7759,N_7760,N_7761,N_7764,N_7765,N_7767,N_7768,N_7774,N_7775,N_7781,N_7783,N_7784,N_7786,N_7787,N_7788,N_7790,N_7791,N_7795,N_7796,N_7797,N_7799,N_7800,N_7801,N_7803,N_7804,N_7806,N_7807,N_7808,N_7810,N_7811,N_7812,N_7813,N_7817,N_7818,N_7821,N_7825,N_7827,N_7828,N_7829,N_7831,N_7832,N_7835,N_7837,N_7840,N_7841,N_7842,N_7843,N_7844,N_7847,N_7848,N_7850,N_7851,N_7852,N_7857,N_7860,N_7861,N_7862,N_7863,N_7864,N_7866,N_7867,N_7869,N_7872,N_7873,N_7875,N_7880,N_7882,N_7883,N_7884,N_7885,N_7888,N_7890,N_7891,N_7892,N_7895,N_7896,N_7897,N_7898,N_7901,N_7902,N_7906,N_7908,N_7909,N_7910,N_7912,N_7915,N_7916,N_7918,N_7919,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7928,N_7930,N_7932,N_7933,N_7934,N_7937,N_7940,N_7941,N_7942,N_7943,N_7945,N_7946,N_7947,N_7948,N_7950,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7961,N_7964,N_7965,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7975,N_7977,N_7978,N_7979,N_7980,N_7982,N_7985,N_7986,N_7991,N_7992,N_7993,N_7996,N_8000,N_8002,N_8005,N_8006,N_8007,N_8011,N_8013,N_8017,N_8018,N_8020,N_8022,N_8024,N_8025,N_8026,N_8027,N_8030,N_8031,N_8032,N_8034,N_8035,N_8038,N_8042,N_8044,N_8047,N_8048,N_8050,N_8053,N_8054,N_8055,N_8056,N_8057,N_8060,N_8061,N_8063,N_8065,N_8066,N_8068,N_8069,N_8070,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8080,N_8084,N_8086,N_8088,N_8089,N_8091,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8100,N_8101,N_8103,N_8104,N_8105,N_8107,N_8109,N_8110,N_8111,N_8113,N_8115,N_8116,N_8118,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8133,N_8134,N_8137,N_8138,N_8140,N_8141,N_8143,N_8148,N_8150,N_8151,N_8155,N_8156,N_8159,N_8160,N_8161,N_8162,N_8166,N_8167,N_8170,N_8171,N_8173,N_8177,N_8181,N_8183,N_8184,N_8186,N_8187,N_8189,N_8190,N_8192,N_8193,N_8197,N_8198,N_8201,N_8202,N_8204,N_8205,N_8206,N_8207,N_8208,N_8210,N_8211,N_8213,N_8214,N_8216,N_8217,N_8218,N_8219,N_8220,N_8222,N_8223,N_8224,N_8225,N_8227,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8241,N_8243,N_8244,N_8245,N_8246,N_8248,N_8249,N_8252,N_8253,N_8254,N_8255,N_8260,N_8261,N_8263,N_8265,N_8267,N_8268,N_8269,N_8272,N_8274,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8294,N_8295,N_8297,N_8298,N_8300,N_8301,N_8303,N_8305,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8320,N_8321,N_8322,N_8324,N_8325,N_8326,N_8327,N_8330,N_8331,N_8332,N_8333,N_8334,N_8337,N_8338,N_8340,N_8343,N_8344,N_8345,N_8348,N_8349,N_8350,N_8351,N_8354,N_8355,N_8357,N_8358,N_8359,N_8360,N_8361,N_8363,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8380,N_8382,N_8383,N_8384,N_8385,N_8387,N_8388,N_8389,N_8392,N_8394,N_8395,N_8396,N_8399,N_8400,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8409,N_8411,N_8413,N_8414,N_8415,N_8416,N_8417,N_8420,N_8421,N_8422,N_8424,N_8427,N_8428,N_8432,N_8433,N_8434,N_8435,N_8438,N_8440,N_8442,N_8444,N_8446,N_8447,N_8452,N_8453,N_8455,N_8456,N_8459,N_8461,N_8462,N_8463,N_8465,N_8466,N_8467,N_8468,N_8469,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8479,N_8480,N_8481,N_8482,N_8483,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8493,N_8495,N_8496,N_8498,N_8500,N_8502,N_8504,N_8506,N_8507,N_8509,N_8512,N_8513,N_8514,N_8517,N_8518,N_8525,N_8532,N_8533,N_8534,N_8535,N_8537,N_8539,N_8541,N_8542,N_8543,N_8544,N_8546,N_8549,N_8551,N_8555,N_8558,N_8559,N_8560,N_8561,N_8563,N_8565,N_8566,N_8568,N_8569,N_8571,N_8572,N_8573,N_8575,N_8577,N_8578,N_8580,N_8581,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8594,N_8599,N_8600,N_8603,N_8605,N_8606,N_8607,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8619,N_8620,N_8622,N_8625,N_8628,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8654,N_8655,N_8656,N_8657,N_8661,N_8663,N_8664,N_8666,N_8667,N_8671,N_8673,N_8674,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8683,N_8684,N_8685,N_8687,N_8688,N_8689,N_8690,N_8692,N_8695,N_8696,N_8697,N_8698,N_8700,N_8702,N_8703,N_8706,N_8707,N_8709,N_8711,N_8712,N_8713,N_8714,N_8715,N_8717,N_8720,N_8721,N_8723,N_8724,N_8726,N_8727,N_8729,N_8730,N_8732,N_8735,N_8737,N_8738,N_8740,N_8747,N_8748,N_8749,N_8750,N_8753,N_8757,N_8758,N_8759,N_8762,N_8763,N_8764,N_8765,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8777,N_8779,N_8780,N_8783,N_8784,N_8785,N_8786,N_8787,N_8789,N_8790,N_8792,N_8795,N_8796,N_8798,N_8801,N_8802,N_8803,N_8804,N_8806,N_8807,N_8808,N_8809,N_8810,N_8812,N_8815,N_8817,N_8818,N_8820,N_8821,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8833,N_8834,N_8838,N_8839,N_8840,N_8841,N_8842,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8853,N_8854,N_8855,N_8856,N_8859,N_8860,N_8861,N_8863,N_8864,N_8865,N_8866,N_8868,N_8869,N_8872,N_8875,N_8879,N_8880,N_8882,N_8884,N_8885,N_8886,N_8888,N_8889,N_8891,N_8895,N_8897,N_8898,N_8900,N_8902,N_8904,N_8905,N_8906,N_8907,N_8909,N_8911,N_8912,N_8914,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8926,N_8927,N_8928,N_8932,N_8933,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8956,N_8958,N_8959,N_8960,N_8962,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8978,N_8979,N_8980,N_8986,N_8987,N_8988,N_8991,N_8992,N_8993,N_8996,N_8998,N_8999,N_9002,N_9003,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9018,N_9019,N_9020,N_9021,N_9024,N_9026,N_9027,N_9028,N_9029,N_9030,N_9033,N_9036,N_9038,N_9039,N_9040,N_9041,N_9045,N_9049,N_9051,N_9053,N_9056,N_9057,N_9059,N_9061,N_9065,N_9066,N_9067,N_9068,N_9069,N_9072,N_9073,N_9075,N_9076,N_9078,N_9079,N_9080,N_9083,N_9084,N_9086,N_9087,N_9088,N_9089,N_9091,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9104,N_9107,N_9109,N_9110,N_9111,N_9113,N_9114,N_9115,N_9118,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9129,N_9130,N_9133,N_9135,N_9136,N_9137,N_9139,N_9141,N_9143,N_9144,N_9145,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9158,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9167,N_9169,N_9170,N_9171,N_9172,N_9174,N_9176,N_9177,N_9178,N_9179,N_9180,N_9182,N_9183,N_9184,N_9186,N_9187,N_9189,N_9190,N_9192,N_9193,N_9194,N_9196,N_9197,N_9198,N_9202,N_9203,N_9205,N_9207,N_9208,N_9209,N_9211,N_9213,N_9214,N_9215,N_9217,N_9218,N_9220,N_9222,N_9223,N_9224,N_9225,N_9227,N_9228,N_9229,N_9230,N_9232,N_9234,N_9235,N_9236,N_9237,N_9241,N_9243,N_9245,N_9246,N_9248,N_9249,N_9250,N_9253,N_9254,N_9255,N_9256,N_9257,N_9260,N_9261,N_9263,N_9264,N_9268,N_9269,N_9270,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9279,N_9281,N_9282,N_9285,N_9288,N_9289,N_9290,N_9294,N_9295,N_9297,N_9298,N_9301,N_9302,N_9305,N_9306,N_9309,N_9310,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9323,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9332,N_9335,N_9336,N_9338,N_9341,N_9342,N_9343,N_9345,N_9347,N_9348,N_9349,N_9352,N_9353,N_9354,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9367,N_9368,N_9369,N_9370,N_9371,N_9375,N_9376,N_9377,N_9379,N_9381,N_9382,N_9383,N_9386,N_9387,N_9390,N_9391,N_9392,N_9395,N_9396,N_9399,N_9402,N_9404,N_9406,N_9407,N_9410,N_9411,N_9412,N_9414,N_9415,N_9419,N_9422,N_9423,N_9424,N_9425,N_9427,N_9428,N_9429,N_9430,N_9431,N_9436,N_9437,N_9439,N_9444,N_9445,N_9446,N_9447,N_9449,N_9451,N_9452,N_9453,N_9456,N_9457,N_9459,N_9460,N_9461,N_9464,N_9465,N_9466,N_9468,N_9470,N_9473,N_9477,N_9479,N_9481,N_9482,N_9484,N_9485,N_9487,N_9488,N_9489,N_9490,N_9492,N_9494,N_9495,N_9497,N_9499,N_9502,N_9503,N_9504,N_9507,N_9508,N_9509,N_9510,N_9512,N_9513,N_9514,N_9515,N_9516,N_9519,N_9520,N_9522,N_9523,N_9525,N_9527,N_9528,N_9529,N_9530,N_9532,N_9536,N_9537,N_9538,N_9541,N_9542,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9551,N_9552,N_9553,N_9555,N_9556,N_9560,N_9563,N_9564,N_9565,N_9566,N_9567,N_9570,N_9573,N_9574,N_9576,N_9577,N_9578,N_9580,N_9581,N_9583,N_9588,N_9589,N_9590,N_9593,N_9596,N_9597,N_9598,N_9599,N_9601,N_9602,N_9603,N_9605,N_9606,N_9607,N_9608,N_9610,N_9614,N_9617,N_9618,N_9621,N_9623,N_9624,N_9626,N_9627,N_9628,N_9630,N_9632,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9641,N_9642,N_9643,N_9646,N_9648,N_9649,N_9652,N_9653,N_9654,N_9655,N_9657,N_9658,N_9659,N_9660,N_9662,N_9663,N_9665,N_9666,N_9667,N_9668,N_9670,N_9671,N_9674,N_9675,N_9678,N_9679,N_9680,N_9682,N_9683,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9693,N_9695,N_9697,N_9698,N_9700,N_9702,N_9708,N_9710,N_9711,N_9712,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9722,N_9724,N_9725,N_9727,N_9729,N_9730,N_9733,N_9735,N_9736,N_9737,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9780,N_9781,N_9782,N_9783,N_9784,N_9787,N_9791,N_9792,N_9793,N_9794,N_9795,N_9799,N_9800,N_9802,N_9803,N_9804,N_9805,N_9808,N_9809,N_9810,N_9811,N_9814,N_9815,N_9818,N_9820,N_9821,N_9822,N_9824,N_9825,N_9826,N_9827,N_9830,N_9832,N_9833,N_9834,N_9835,N_9838,N_9839,N_9841,N_9842,N_9846,N_9847,N_9849,N_9852,N_9855,N_9856,N_9862,N_9864,N_9865,N_9866,N_9867,N_9870,N_9871,N_9876,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9891,N_9892,N_9893,N_9895,N_9897,N_9899,N_9902,N_9904,N_9905,N_9906,N_9912,N_9914,N_9918,N_9919,N_9921,N_9922,N_9923,N_9924,N_9929,N_9930,N_9932,N_9935,N_9936,N_9940,N_9941,N_9942,N_9943,N_9945,N_9948,N_9950,N_9951,N_9952,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9962,N_9963,N_9964,N_9966,N_9968,N_9969,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9978,N_9988,N_9990,N_9993,N_9994,N_9995,N_9997,N_9998;
nand U0 (N_0,In_939,In_497);
xnor U1 (N_1,In_673,In_638);
nand U2 (N_2,In_137,In_754);
nand U3 (N_3,In_354,In_614);
and U4 (N_4,In_559,In_398);
or U5 (N_5,In_345,In_310);
nor U6 (N_6,In_613,In_883);
nor U7 (N_7,In_427,In_29);
nand U8 (N_8,In_641,In_402);
nor U9 (N_9,In_218,In_950);
and U10 (N_10,In_549,In_831);
or U11 (N_11,In_653,In_867);
and U12 (N_12,In_180,In_57);
nor U13 (N_13,In_32,In_174);
or U14 (N_14,In_448,In_335);
xnor U15 (N_15,In_666,In_557);
and U16 (N_16,In_251,In_708);
xor U17 (N_17,In_213,In_717);
and U18 (N_18,In_524,In_927);
or U19 (N_19,In_633,In_678);
nor U20 (N_20,In_445,In_346);
or U21 (N_21,In_479,In_366);
nor U22 (N_22,In_98,In_45);
nand U23 (N_23,In_483,In_709);
nor U24 (N_24,In_914,In_327);
or U25 (N_25,In_101,In_278);
nand U26 (N_26,In_547,In_753);
and U27 (N_27,In_150,In_201);
nand U28 (N_28,In_906,In_655);
or U29 (N_29,In_772,In_509);
xor U30 (N_30,In_735,In_811);
and U31 (N_31,In_338,In_15);
nand U32 (N_32,In_241,In_486);
and U33 (N_33,In_897,In_853);
and U34 (N_34,In_788,In_570);
nand U35 (N_35,In_349,In_211);
nand U36 (N_36,In_224,In_341);
nor U37 (N_37,In_615,In_191);
and U38 (N_38,In_250,In_287);
and U39 (N_39,In_563,In_551);
nand U40 (N_40,In_108,In_798);
or U41 (N_41,In_83,In_706);
nand U42 (N_42,In_409,In_473);
nand U43 (N_43,In_314,In_694);
nor U44 (N_44,In_890,In_151);
or U45 (N_45,In_520,In_422);
xor U46 (N_46,In_755,In_431);
nor U47 (N_47,In_229,In_234);
nand U48 (N_48,In_836,In_702);
nor U49 (N_49,In_693,In_809);
nor U50 (N_50,In_107,In_386);
nand U51 (N_51,In_685,In_919);
nor U52 (N_52,In_256,In_160);
nor U53 (N_53,In_604,In_19);
nor U54 (N_54,In_730,In_36);
nor U55 (N_55,In_987,In_624);
or U56 (N_56,In_627,In_301);
nand U57 (N_57,In_665,In_710);
nor U58 (N_58,In_235,In_356);
nand U59 (N_59,In_54,In_724);
and U60 (N_60,In_6,In_149);
and U61 (N_61,In_109,In_536);
or U62 (N_62,In_767,In_962);
and U63 (N_63,In_843,In_253);
or U64 (N_64,In_630,In_46);
nor U65 (N_65,In_552,In_106);
nor U66 (N_66,In_857,In_421);
nand U67 (N_67,In_806,In_320);
xnor U68 (N_68,In_865,In_646);
nor U69 (N_69,In_472,In_779);
and U70 (N_70,In_24,In_134);
nand U71 (N_71,In_50,In_114);
nor U72 (N_72,In_839,In_858);
and U73 (N_73,In_662,In_171);
xnor U74 (N_74,In_924,In_1);
and U75 (N_75,In_949,In_203);
and U76 (N_76,In_823,In_654);
nand U77 (N_77,In_944,In_429);
nand U78 (N_78,In_566,In_896);
nor U79 (N_79,In_885,In_78);
xnor U80 (N_80,In_959,In_980);
nor U81 (N_81,In_734,In_447);
nor U82 (N_82,In_585,In_481);
nand U83 (N_83,In_827,In_935);
and U84 (N_84,In_740,In_277);
or U85 (N_85,In_202,In_406);
nor U86 (N_86,In_417,In_308);
nor U87 (N_87,In_657,In_321);
and U88 (N_88,In_367,In_494);
xor U89 (N_89,In_501,In_131);
xnor U90 (N_90,In_842,In_999);
nand U91 (N_91,In_936,In_122);
and U92 (N_92,In_758,In_153);
nor U93 (N_93,In_855,In_219);
nor U94 (N_94,In_197,In_969);
nand U95 (N_95,In_726,In_640);
nand U96 (N_96,In_616,In_993);
nand U97 (N_97,In_820,In_254);
nand U98 (N_98,In_928,In_30);
and U99 (N_99,In_922,In_991);
nand U100 (N_100,In_818,In_263);
and U101 (N_101,In_355,In_701);
nand U102 (N_102,In_182,In_350);
and U103 (N_103,In_739,In_911);
or U104 (N_104,In_597,In_59);
or U105 (N_105,In_112,In_787);
or U106 (N_106,In_157,In_455);
nand U107 (N_107,In_282,In_230);
and U108 (N_108,In_903,In_410);
nand U109 (N_109,In_53,In_246);
nand U110 (N_110,In_485,In_220);
and U111 (N_111,In_889,In_783);
and U112 (N_112,In_271,In_871);
nand U113 (N_113,In_348,In_847);
or U114 (N_114,In_439,In_824);
nand U115 (N_115,In_718,In_393);
nand U116 (N_116,In_69,In_281);
nor U117 (N_117,In_713,In_937);
and U118 (N_118,In_893,In_913);
nand U119 (N_119,In_103,In_420);
or U120 (N_120,In_637,In_72);
nand U121 (N_121,In_407,In_769);
and U122 (N_122,In_631,In_199);
nor U123 (N_123,In_676,In_155);
nor U124 (N_124,In_66,In_68);
nand U125 (N_125,In_961,In_626);
or U126 (N_126,In_189,In_298);
and U127 (N_127,In_623,In_248);
nor U128 (N_128,In_568,In_216);
xnor U129 (N_129,In_771,In_403);
nor U130 (N_130,In_21,In_309);
nor U131 (N_131,In_698,In_791);
and U132 (N_132,In_304,In_786);
nand U133 (N_133,In_877,In_533);
nor U134 (N_134,In_195,In_577);
or U135 (N_135,In_147,In_292);
and U136 (N_136,In_430,In_644);
and U137 (N_137,In_848,In_516);
nor U138 (N_138,In_729,In_784);
and U139 (N_139,In_840,In_469);
nand U140 (N_140,In_981,In_505);
nor U141 (N_141,In_280,In_880);
and U142 (N_142,In_405,In_428);
nand U143 (N_143,In_440,In_800);
nor U144 (N_144,In_661,In_359);
or U145 (N_145,In_61,In_764);
or U146 (N_146,In_766,In_863);
and U147 (N_147,In_506,In_663);
and U148 (N_148,In_221,In_602);
nor U149 (N_149,In_84,In_968);
and U150 (N_150,In_841,In_294);
nor U151 (N_151,In_44,In_580);
nand U152 (N_152,In_144,In_25);
nor U153 (N_153,In_521,In_894);
and U154 (N_154,In_443,In_782);
and U155 (N_155,In_650,In_917);
xnor U156 (N_156,In_139,In_869);
or U157 (N_157,In_777,In_289);
nand U158 (N_158,In_920,In_601);
or U159 (N_159,In_90,In_468);
and U160 (N_160,In_974,In_165);
or U161 (N_161,In_99,In_682);
or U162 (N_162,In_105,In_11);
or U163 (N_163,In_873,In_528);
nand U164 (N_164,In_965,In_493);
or U165 (N_165,In_462,In_146);
or U166 (N_166,In_856,In_373);
or U167 (N_167,In_138,In_38);
nand U168 (N_168,In_378,In_530);
or U169 (N_169,In_882,In_612);
or U170 (N_170,In_502,In_91);
and U171 (N_171,In_63,In_778);
nand U172 (N_172,In_985,In_870);
nand U173 (N_173,In_757,In_140);
or U174 (N_174,In_934,In_408);
and U175 (N_175,In_544,In_929);
or U176 (N_176,In_744,In_411);
or U177 (N_177,In_37,In_542);
nand U178 (N_178,In_243,In_947);
nand U179 (N_179,In_82,In_802);
or U180 (N_180,In_244,In_908);
nor U181 (N_181,In_994,In_433);
or U182 (N_182,In_187,In_941);
nand U183 (N_183,In_982,In_697);
nor U184 (N_184,In_353,In_184);
nand U185 (N_185,In_384,In_515);
and U186 (N_186,In_56,In_326);
nand U187 (N_187,In_635,In_838);
nor U188 (N_188,In_340,In_450);
or U189 (N_189,In_303,In_539);
nor U190 (N_190,In_988,In_854);
or U191 (N_191,In_311,In_441);
and U192 (N_192,In_900,In_330);
nand U193 (N_193,In_383,In_196);
nand U194 (N_194,In_984,In_691);
nand U195 (N_195,In_275,In_526);
or U196 (N_196,In_826,In_159);
and U197 (N_197,In_859,In_487);
nand U198 (N_198,In_902,In_476);
or U199 (N_199,In_537,In_651);
xnor U200 (N_200,In_747,In_992);
nor U201 (N_201,In_997,In_742);
or U202 (N_202,In_933,In_971);
nor U203 (N_203,In_47,In_266);
nor U204 (N_204,In_290,In_168);
and U205 (N_205,In_972,In_491);
xnor U206 (N_206,In_674,In_901);
nor U207 (N_207,In_156,In_833);
and U208 (N_208,In_344,In_531);
nand U209 (N_209,In_444,In_609);
nor U210 (N_210,In_495,In_436);
xnor U211 (N_211,In_286,In_619);
or U212 (N_212,In_267,In_372);
or U213 (N_213,In_368,In_329);
or U214 (N_214,In_86,In_352);
nand U215 (N_215,In_212,In_273);
nor U216 (N_216,In_943,In_336);
nand U217 (N_217,In_181,In_252);
nor U218 (N_218,In_318,In_208);
xnor U219 (N_219,In_423,In_459);
nand U220 (N_220,In_194,In_860);
or U221 (N_221,In_104,In_895);
xnor U222 (N_222,In_162,In_652);
and U223 (N_223,In_228,In_500);
nor U224 (N_224,In_279,In_775);
nand U225 (N_225,In_915,In_357);
nand U226 (N_226,In_283,In_42);
nand U227 (N_227,In_371,In_300);
nor U228 (N_228,In_804,In_231);
nand U229 (N_229,In_39,In_593);
nand U230 (N_230,In_781,In_334);
xnor U231 (N_231,In_611,In_770);
nor U232 (N_232,In_7,In_686);
or U233 (N_233,In_70,In_498);
nand U234 (N_234,In_822,In_31);
xor U235 (N_235,In_790,In_888);
and U236 (N_236,In_206,In_288);
and U237 (N_237,In_799,In_741);
or U238 (N_238,In_930,In_97);
nor U239 (N_239,In_28,In_389);
or U240 (N_240,In_600,In_55);
nor U241 (N_241,In_369,In_51);
nand U242 (N_242,In_511,In_222);
and U243 (N_243,In_8,In_617);
and U244 (N_244,In_2,In_148);
or U245 (N_245,In_390,In_412);
xor U246 (N_246,In_503,In_392);
nor U247 (N_247,In_100,In_690);
or U248 (N_248,In_80,In_795);
or U249 (N_249,In_164,In_245);
nor U250 (N_250,In_9,In_377);
and U251 (N_251,In_425,In_746);
nor U252 (N_252,In_451,In_482);
nand U253 (N_253,In_722,In_810);
or U254 (N_254,In_591,In_830);
xnor U255 (N_255,In_305,In_170);
or U256 (N_256,In_794,In_875);
xor U257 (N_257,In_912,In_948);
nand U258 (N_258,In_796,In_967);
nand U259 (N_259,In_845,In_513);
and U260 (N_260,In_884,In_264);
xnor U261 (N_261,In_262,In_608);
nand U262 (N_262,In_26,In_480);
xnor U263 (N_263,In_517,In_133);
nor U264 (N_264,In_215,In_89);
nand U265 (N_265,In_898,In_382);
nand U266 (N_266,In_93,In_743);
or U267 (N_267,In_270,In_233);
nand U268 (N_268,In_177,In_761);
or U269 (N_269,In_669,In_565);
or U270 (N_270,In_175,In_508);
or U271 (N_271,In_65,In_360);
or U272 (N_272,In_34,In_71);
nand U273 (N_273,In_79,In_16);
or U274 (N_274,In_970,In_548);
and U275 (N_275,In_899,In_124);
nand U276 (N_276,In_477,In_257);
nand U277 (N_277,In_966,In_603);
nor U278 (N_278,In_169,In_695);
and U279 (N_279,In_453,In_258);
and U280 (N_280,In_188,In_276);
xor U281 (N_281,In_200,In_861);
or U282 (N_282,In_622,In_123);
or U283 (N_283,In_328,In_681);
and U284 (N_284,In_571,In_475);
xnor U285 (N_285,In_752,In_538);
and U286 (N_286,In_337,In_499);
nor U287 (N_287,In_945,In_470);
nor U288 (N_288,In_76,In_395);
and U289 (N_289,In_478,In_269);
and U290 (N_290,In_699,In_20);
nand U291 (N_291,In_550,In_291);
or U292 (N_292,In_963,In_192);
and U293 (N_293,In_522,In_639);
or U294 (N_294,In_413,In_995);
and U295 (N_295,In_738,In_573);
xnor U296 (N_296,In_998,In_926);
nand U297 (N_297,In_376,In_683);
nand U298 (N_298,In_135,In_117);
and U299 (N_299,In_714,In_307);
nor U300 (N_300,In_973,In_774);
or U301 (N_301,In_768,In_620);
nor U302 (N_302,In_904,In_362);
or U303 (N_303,In_813,In_582);
nand U304 (N_304,In_572,In_595);
and U305 (N_305,In_154,In_143);
or U306 (N_306,In_780,In_465);
and U307 (N_307,In_649,In_725);
nand U308 (N_308,In_862,In_596);
or U309 (N_309,In_918,In_696);
nor U310 (N_310,In_598,In_461);
nor U311 (N_311,In_272,In_750);
or U312 (N_312,In_977,In_553);
xor U313 (N_313,In_989,In_113);
and U314 (N_314,In_299,In_887);
and U315 (N_315,In_789,In_414);
xor U316 (N_316,In_496,In_715);
and U317 (N_317,In_932,In_592);
and U318 (N_318,In_792,In_460);
nand U319 (N_319,In_689,In_575);
and U320 (N_320,In_74,In_940);
xnor U321 (N_321,In_825,In_910);
or U322 (N_322,In_864,In_958);
xnor U323 (N_323,In_656,In_532);
or U324 (N_324,In_95,In_556);
or U325 (N_325,In_688,In_751);
nor U326 (N_326,In_529,In_81);
or U327 (N_327,In_849,In_343);
nor U328 (N_328,In_952,In_17);
nor U329 (N_329,In_721,In_178);
and U330 (N_330,In_803,In_832);
or U331 (N_331,In_293,In_437);
nor U332 (N_332,In_642,In_466);
and U333 (N_333,In_748,In_645);
and U334 (N_334,In_161,In_942);
nand U335 (N_335,In_546,In_921);
nand U336 (N_336,In_331,In_527);
and U337 (N_337,In_534,In_363);
and U338 (N_338,In_332,In_675);
and U339 (N_339,In_142,In_816);
xor U340 (N_340,In_834,In_578);
nand U341 (N_341,In_956,In_878);
nor U342 (N_342,In_664,In_679);
xor U343 (N_343,In_40,In_247);
or U344 (N_344,In_687,In_285);
xnor U345 (N_345,In_115,In_760);
nor U346 (N_346,In_850,In_732);
or U347 (N_347,In_110,In_35);
nand U348 (N_348,In_576,In_765);
or U349 (N_349,In_454,In_589);
nor U350 (N_350,In_558,In_306);
nand U351 (N_351,In_628,In_381);
nor U352 (N_352,In_385,In_23);
and U353 (N_353,In_166,In_957);
nand U354 (N_354,In_773,In_905);
or U355 (N_355,In_916,In_951);
xnor U356 (N_356,In_4,In_255);
or U357 (N_357,In_3,In_567);
or U358 (N_358,In_835,In_435);
and U359 (N_359,In_733,In_446);
and U360 (N_360,In_313,In_274);
nand U361 (N_361,In_677,In_866);
nor U362 (N_362,In_130,In_605);
nor U363 (N_363,In_400,In_172);
or U364 (N_364,In_762,In_519);
and U365 (N_365,In_312,In_490);
or U366 (N_366,In_394,In_464);
nor U367 (N_367,In_955,In_643);
nand U368 (N_368,In_684,In_574);
nand U369 (N_369,In_260,In_805);
nor U370 (N_370,In_126,In_886);
nor U371 (N_371,In_418,In_284);
nor U372 (N_372,In_720,In_756);
and U373 (N_373,In_672,In_152);
nand U374 (N_374,In_88,In_380);
xor U375 (N_375,In_671,In_632);
and U376 (N_376,In_12,In_27);
nor U377 (N_377,In_296,In_43);
and U378 (N_378,In_660,In_295);
and U379 (N_379,In_227,In_561);
nand U380 (N_380,In_909,In_358);
or U381 (N_381,In_562,In_815);
nand U382 (N_382,In_236,In_10);
and U383 (N_383,In_116,In_237);
or U384 (N_384,In_938,In_586);
nand U385 (N_385,In_323,In_749);
nand U386 (N_386,In_62,In_587);
nand U387 (N_387,In_793,In_302);
xor U388 (N_388,In_173,In_731);
and U389 (N_389,In_210,In_317);
and U390 (N_390,In_463,In_183);
nand U391 (N_391,In_179,In_193);
nand U392 (N_392,In_77,In_18);
and U393 (N_393,In_512,In_401);
and U394 (N_394,In_960,In_983);
nand U395 (N_395,In_259,In_419);
and U396 (N_396,In_484,In_555);
nor U397 (N_397,In_351,In_703);
nand U398 (N_398,In_426,In_396);
and U399 (N_399,In_370,In_723);
and U400 (N_400,In_121,In_711);
and U401 (N_401,In_606,In_978);
nand U402 (N_402,In_700,In_759);
and U403 (N_403,In_523,In_892);
or U404 (N_404,In_996,In_667);
or U405 (N_405,In_239,In_541);
or U406 (N_406,In_658,In_207);
nor U407 (N_407,In_821,In_41);
nor U408 (N_408,In_391,In_986);
nand U409 (N_409,In_96,In_119);
or U410 (N_410,In_670,In_881);
nor U411 (N_411,In_594,In_388);
nand U412 (N_412,In_876,In_205);
or U413 (N_413,In_668,In_797);
nor U414 (N_414,In_190,In_891);
or U415 (N_415,In_648,In_434);
nor U416 (N_416,In_58,In_564);
nor U417 (N_417,In_238,In_879);
nor U418 (N_418,In_158,In_492);
xor U419 (N_419,In_33,In_315);
and U420 (N_420,In_136,In_52);
nand U421 (N_421,In_535,In_727);
nand U422 (N_422,In_471,In_814);
nand U423 (N_423,In_223,In_785);
and U424 (N_424,In_925,In_186);
nor U425 (N_425,In_584,In_680);
and U426 (N_426,In_375,In_73);
or U427 (N_427,In_120,In_75);
nand U428 (N_428,In_510,In_736);
nand U429 (N_429,In_504,In_416);
or U430 (N_430,In_449,In_812);
and U431 (N_431,In_339,In_452);
nor U432 (N_432,In_704,In_808);
or U433 (N_433,In_198,In_325);
xnor U434 (N_434,In_514,In_242);
nor U435 (N_435,In_923,In_716);
and U436 (N_436,In_111,In_705);
nor U437 (N_437,In_852,In_127);
and U438 (N_438,In_387,In_581);
nor U439 (N_439,In_217,In_85);
or U440 (N_440,In_692,In_456);
or U441 (N_441,In_129,In_844);
or U442 (N_442,In_240,In_379);
nand U443 (N_443,In_361,In_953);
nand U444 (N_444,In_322,In_851);
and U445 (N_445,In_364,In_232);
nand U446 (N_446,In_518,In_268);
nand U447 (N_447,In_979,In_457);
nor U448 (N_448,In_807,In_817);
nor U449 (N_449,In_946,In_399);
nand U450 (N_450,In_588,In_990);
and U451 (N_451,In_347,In_209);
and U452 (N_452,In_297,In_261);
nor U453 (N_453,In_931,In_625);
and U454 (N_454,In_226,In_907);
and U455 (N_455,In_14,In_975);
and U456 (N_456,In_543,In_560);
and U457 (N_457,In_607,In_488);
nand U458 (N_458,In_438,In_442);
nor U459 (N_459,In_801,In_319);
nand U460 (N_460,In_67,In_404);
nand U461 (N_461,In_432,In_13);
xnor U462 (N_462,In_728,In_87);
or U463 (N_463,In_540,In_397);
nand U464 (N_464,In_610,In_636);
and U465 (N_465,In_819,In_874);
or U466 (N_466,In_964,In_48);
and U467 (N_467,In_265,In_145);
nand U468 (N_468,In_94,In_324);
and U469 (N_469,In_204,In_763);
nand U470 (N_470,In_333,In_141);
xnor U471 (N_471,In_176,In_629);
or U472 (N_472,In_22,In_976);
nand U473 (N_473,In_132,In_92);
or U474 (N_474,In_5,In_374);
or U475 (N_475,In_554,In_424);
or U476 (N_476,In_128,In_525);
and U477 (N_477,In_474,In_583);
nand U478 (N_478,In_64,In_829);
and U479 (N_479,In_249,In_569);
xnor U480 (N_480,In_828,In_214);
nand U481 (N_481,In_846,In_125);
and U482 (N_482,In_467,In_621);
and U483 (N_483,In_719,In_545);
nand U484 (N_484,In_60,In_167);
nor U485 (N_485,In_590,In_837);
or U486 (N_486,In_415,In_225);
nor U487 (N_487,In_163,In_647);
and U488 (N_488,In_634,In_342);
xnor U489 (N_489,In_365,In_712);
nor U490 (N_490,In_489,In_707);
nor U491 (N_491,In_599,In_872);
nor U492 (N_492,In_507,In_745);
and U493 (N_493,In_737,In_579);
and U494 (N_494,In_316,In_185);
nor U495 (N_495,In_618,In_776);
nor U496 (N_496,In_868,In_0);
nand U497 (N_497,In_458,In_49);
nand U498 (N_498,In_118,In_102);
and U499 (N_499,In_659,In_954);
or U500 (N_500,In_50,In_693);
nor U501 (N_501,In_284,In_16);
and U502 (N_502,In_727,In_963);
or U503 (N_503,In_262,In_477);
and U504 (N_504,In_711,In_577);
or U505 (N_505,In_920,In_412);
and U506 (N_506,In_292,In_347);
and U507 (N_507,In_165,In_458);
or U508 (N_508,In_331,In_568);
xnor U509 (N_509,In_616,In_86);
nor U510 (N_510,In_10,In_348);
nand U511 (N_511,In_776,In_428);
nor U512 (N_512,In_356,In_853);
and U513 (N_513,In_181,In_646);
or U514 (N_514,In_812,In_954);
and U515 (N_515,In_15,In_420);
and U516 (N_516,In_511,In_271);
and U517 (N_517,In_402,In_180);
and U518 (N_518,In_120,In_335);
or U519 (N_519,In_150,In_292);
or U520 (N_520,In_285,In_404);
or U521 (N_521,In_456,In_888);
or U522 (N_522,In_711,In_583);
or U523 (N_523,In_962,In_948);
nor U524 (N_524,In_859,In_755);
nor U525 (N_525,In_748,In_241);
or U526 (N_526,In_117,In_975);
nor U527 (N_527,In_81,In_600);
or U528 (N_528,In_379,In_985);
or U529 (N_529,In_226,In_170);
nand U530 (N_530,In_727,In_700);
or U531 (N_531,In_196,In_444);
nor U532 (N_532,In_232,In_225);
and U533 (N_533,In_815,In_982);
nor U534 (N_534,In_463,In_19);
nand U535 (N_535,In_478,In_188);
nand U536 (N_536,In_743,In_834);
and U537 (N_537,In_296,In_495);
nor U538 (N_538,In_852,In_583);
nor U539 (N_539,In_571,In_942);
nand U540 (N_540,In_824,In_698);
or U541 (N_541,In_191,In_3);
nand U542 (N_542,In_969,In_217);
nand U543 (N_543,In_605,In_988);
xnor U544 (N_544,In_32,In_677);
nor U545 (N_545,In_417,In_130);
or U546 (N_546,In_532,In_600);
or U547 (N_547,In_764,In_196);
and U548 (N_548,In_110,In_703);
nor U549 (N_549,In_672,In_712);
nand U550 (N_550,In_619,In_341);
and U551 (N_551,In_63,In_188);
nand U552 (N_552,In_273,In_927);
nor U553 (N_553,In_150,In_334);
nand U554 (N_554,In_326,In_281);
and U555 (N_555,In_845,In_120);
nand U556 (N_556,In_142,In_844);
and U557 (N_557,In_232,In_473);
nor U558 (N_558,In_691,In_446);
and U559 (N_559,In_461,In_415);
nor U560 (N_560,In_219,In_689);
or U561 (N_561,In_398,In_156);
nor U562 (N_562,In_307,In_20);
nor U563 (N_563,In_389,In_476);
xor U564 (N_564,In_552,In_507);
and U565 (N_565,In_398,In_753);
nand U566 (N_566,In_987,In_234);
and U567 (N_567,In_585,In_223);
and U568 (N_568,In_789,In_132);
xnor U569 (N_569,In_908,In_39);
nor U570 (N_570,In_47,In_66);
or U571 (N_571,In_412,In_641);
nand U572 (N_572,In_595,In_389);
nand U573 (N_573,In_344,In_179);
nor U574 (N_574,In_508,In_243);
and U575 (N_575,In_340,In_537);
nand U576 (N_576,In_22,In_746);
or U577 (N_577,In_225,In_313);
or U578 (N_578,In_419,In_745);
and U579 (N_579,In_759,In_256);
and U580 (N_580,In_444,In_882);
or U581 (N_581,In_999,In_584);
or U582 (N_582,In_153,In_391);
and U583 (N_583,In_854,In_524);
nand U584 (N_584,In_266,In_93);
or U585 (N_585,In_620,In_698);
or U586 (N_586,In_434,In_235);
nand U587 (N_587,In_815,In_976);
nor U588 (N_588,In_129,In_31);
nand U589 (N_589,In_991,In_944);
and U590 (N_590,In_751,In_503);
nand U591 (N_591,In_445,In_590);
nor U592 (N_592,In_512,In_694);
or U593 (N_593,In_621,In_557);
nor U594 (N_594,In_932,In_931);
nand U595 (N_595,In_634,In_549);
nand U596 (N_596,In_846,In_840);
nor U597 (N_597,In_74,In_15);
or U598 (N_598,In_134,In_241);
or U599 (N_599,In_300,In_199);
nor U600 (N_600,In_261,In_577);
or U601 (N_601,In_134,In_381);
nand U602 (N_602,In_71,In_395);
and U603 (N_603,In_432,In_726);
nor U604 (N_604,In_884,In_792);
nor U605 (N_605,In_119,In_77);
nand U606 (N_606,In_966,In_255);
nor U607 (N_607,In_449,In_333);
or U608 (N_608,In_421,In_593);
nand U609 (N_609,In_173,In_955);
or U610 (N_610,In_564,In_925);
or U611 (N_611,In_729,In_270);
nor U612 (N_612,In_469,In_403);
and U613 (N_613,In_179,In_568);
nor U614 (N_614,In_907,In_853);
nand U615 (N_615,In_109,In_195);
xor U616 (N_616,In_198,In_341);
nor U617 (N_617,In_393,In_225);
nor U618 (N_618,In_211,In_28);
and U619 (N_619,In_705,In_486);
xnor U620 (N_620,In_720,In_40);
and U621 (N_621,In_685,In_469);
nor U622 (N_622,In_390,In_993);
or U623 (N_623,In_555,In_827);
nand U624 (N_624,In_660,In_559);
and U625 (N_625,In_910,In_311);
nand U626 (N_626,In_588,In_403);
nor U627 (N_627,In_904,In_619);
nor U628 (N_628,In_149,In_648);
and U629 (N_629,In_315,In_22);
xor U630 (N_630,In_266,In_805);
or U631 (N_631,In_147,In_797);
xor U632 (N_632,In_439,In_108);
nand U633 (N_633,In_707,In_476);
or U634 (N_634,In_607,In_230);
and U635 (N_635,In_910,In_65);
nand U636 (N_636,In_977,In_14);
or U637 (N_637,In_853,In_975);
nand U638 (N_638,In_125,In_672);
and U639 (N_639,In_219,In_41);
or U640 (N_640,In_815,In_69);
xnor U641 (N_641,In_560,In_275);
or U642 (N_642,In_281,In_567);
nand U643 (N_643,In_692,In_995);
nor U644 (N_644,In_273,In_791);
and U645 (N_645,In_354,In_281);
and U646 (N_646,In_605,In_853);
nor U647 (N_647,In_282,In_900);
or U648 (N_648,In_287,In_264);
nor U649 (N_649,In_170,In_117);
or U650 (N_650,In_540,In_468);
and U651 (N_651,In_322,In_304);
nor U652 (N_652,In_378,In_114);
nor U653 (N_653,In_801,In_629);
nand U654 (N_654,In_79,In_954);
nand U655 (N_655,In_238,In_79);
nor U656 (N_656,In_775,In_584);
and U657 (N_657,In_902,In_972);
nand U658 (N_658,In_820,In_106);
or U659 (N_659,In_458,In_17);
nand U660 (N_660,In_210,In_576);
and U661 (N_661,In_323,In_900);
and U662 (N_662,In_982,In_424);
and U663 (N_663,In_354,In_680);
or U664 (N_664,In_17,In_249);
nor U665 (N_665,In_777,In_103);
and U666 (N_666,In_204,In_934);
nor U667 (N_667,In_239,In_752);
nand U668 (N_668,In_277,In_831);
and U669 (N_669,In_471,In_376);
and U670 (N_670,In_628,In_355);
nand U671 (N_671,In_939,In_466);
nand U672 (N_672,In_788,In_4);
or U673 (N_673,In_871,In_502);
and U674 (N_674,In_316,In_409);
or U675 (N_675,In_896,In_795);
and U676 (N_676,In_666,In_562);
and U677 (N_677,In_313,In_644);
nor U678 (N_678,In_793,In_92);
nand U679 (N_679,In_685,In_566);
nand U680 (N_680,In_737,In_802);
nor U681 (N_681,In_370,In_336);
or U682 (N_682,In_515,In_661);
and U683 (N_683,In_836,In_745);
and U684 (N_684,In_32,In_426);
or U685 (N_685,In_644,In_823);
xor U686 (N_686,In_893,In_81);
nand U687 (N_687,In_960,In_148);
nor U688 (N_688,In_832,In_892);
nand U689 (N_689,In_716,In_806);
nor U690 (N_690,In_166,In_191);
nor U691 (N_691,In_662,In_888);
or U692 (N_692,In_655,In_757);
xnor U693 (N_693,In_385,In_486);
xor U694 (N_694,In_319,In_663);
and U695 (N_695,In_359,In_644);
xor U696 (N_696,In_890,In_472);
nand U697 (N_697,In_633,In_916);
or U698 (N_698,In_364,In_259);
xor U699 (N_699,In_664,In_558);
nand U700 (N_700,In_838,In_224);
and U701 (N_701,In_145,In_761);
nor U702 (N_702,In_727,In_100);
or U703 (N_703,In_643,In_875);
nor U704 (N_704,In_486,In_756);
and U705 (N_705,In_433,In_127);
nand U706 (N_706,In_71,In_670);
nor U707 (N_707,In_765,In_55);
nand U708 (N_708,In_53,In_44);
nand U709 (N_709,In_952,In_13);
or U710 (N_710,In_104,In_134);
nand U711 (N_711,In_899,In_240);
nand U712 (N_712,In_881,In_932);
or U713 (N_713,In_907,In_373);
xor U714 (N_714,In_208,In_876);
nand U715 (N_715,In_906,In_419);
or U716 (N_716,In_626,In_702);
and U717 (N_717,In_803,In_251);
or U718 (N_718,In_169,In_663);
and U719 (N_719,In_255,In_330);
and U720 (N_720,In_422,In_515);
nor U721 (N_721,In_179,In_994);
nor U722 (N_722,In_382,In_31);
nand U723 (N_723,In_717,In_77);
xnor U724 (N_724,In_565,In_7);
nand U725 (N_725,In_48,In_710);
xor U726 (N_726,In_368,In_488);
and U727 (N_727,In_73,In_781);
nand U728 (N_728,In_467,In_611);
nor U729 (N_729,In_449,In_480);
and U730 (N_730,In_301,In_203);
nand U731 (N_731,In_950,In_663);
or U732 (N_732,In_956,In_160);
and U733 (N_733,In_325,In_44);
nand U734 (N_734,In_293,In_168);
or U735 (N_735,In_205,In_30);
and U736 (N_736,In_554,In_334);
and U737 (N_737,In_412,In_191);
or U738 (N_738,In_474,In_105);
or U739 (N_739,In_819,In_781);
nor U740 (N_740,In_782,In_172);
nor U741 (N_741,In_342,In_869);
nand U742 (N_742,In_238,In_427);
nor U743 (N_743,In_936,In_178);
nor U744 (N_744,In_374,In_187);
nand U745 (N_745,In_994,In_380);
nor U746 (N_746,In_945,In_454);
nand U747 (N_747,In_799,In_962);
and U748 (N_748,In_521,In_670);
nand U749 (N_749,In_369,In_228);
nand U750 (N_750,In_140,In_917);
nor U751 (N_751,In_222,In_149);
xor U752 (N_752,In_663,In_647);
nor U753 (N_753,In_557,In_488);
nor U754 (N_754,In_602,In_37);
nand U755 (N_755,In_203,In_536);
nand U756 (N_756,In_314,In_355);
nand U757 (N_757,In_276,In_55);
nand U758 (N_758,In_970,In_439);
and U759 (N_759,In_173,In_986);
nand U760 (N_760,In_662,In_568);
or U761 (N_761,In_843,In_479);
and U762 (N_762,In_834,In_598);
nand U763 (N_763,In_913,In_617);
xnor U764 (N_764,In_102,In_141);
or U765 (N_765,In_571,In_744);
xnor U766 (N_766,In_308,In_598);
and U767 (N_767,In_759,In_407);
nor U768 (N_768,In_730,In_994);
xor U769 (N_769,In_920,In_9);
xnor U770 (N_770,In_535,In_435);
or U771 (N_771,In_605,In_566);
nand U772 (N_772,In_392,In_72);
and U773 (N_773,In_203,In_218);
nand U774 (N_774,In_754,In_624);
and U775 (N_775,In_340,In_59);
nand U776 (N_776,In_918,In_281);
or U777 (N_777,In_27,In_307);
nor U778 (N_778,In_892,In_605);
and U779 (N_779,In_385,In_779);
and U780 (N_780,In_424,In_710);
and U781 (N_781,In_632,In_920);
and U782 (N_782,In_257,In_505);
and U783 (N_783,In_531,In_733);
or U784 (N_784,In_253,In_364);
nor U785 (N_785,In_887,In_440);
xor U786 (N_786,In_927,In_944);
and U787 (N_787,In_443,In_398);
nor U788 (N_788,In_649,In_652);
or U789 (N_789,In_202,In_189);
and U790 (N_790,In_423,In_763);
nor U791 (N_791,In_0,In_25);
nand U792 (N_792,In_372,In_962);
or U793 (N_793,In_652,In_40);
nand U794 (N_794,In_299,In_36);
nand U795 (N_795,In_841,In_150);
or U796 (N_796,In_442,In_363);
or U797 (N_797,In_114,In_755);
and U798 (N_798,In_752,In_777);
or U799 (N_799,In_839,In_476);
nand U800 (N_800,In_739,In_661);
or U801 (N_801,In_631,In_575);
nor U802 (N_802,In_114,In_355);
or U803 (N_803,In_401,In_133);
nand U804 (N_804,In_915,In_548);
xnor U805 (N_805,In_34,In_691);
nand U806 (N_806,In_622,In_86);
nor U807 (N_807,In_837,In_926);
or U808 (N_808,In_718,In_365);
xnor U809 (N_809,In_615,In_185);
xor U810 (N_810,In_96,In_880);
nand U811 (N_811,In_180,In_806);
nand U812 (N_812,In_612,In_852);
or U813 (N_813,In_831,In_458);
xor U814 (N_814,In_491,In_755);
or U815 (N_815,In_658,In_927);
nor U816 (N_816,In_924,In_905);
xor U817 (N_817,In_17,In_914);
nand U818 (N_818,In_818,In_599);
or U819 (N_819,In_439,In_698);
nand U820 (N_820,In_556,In_694);
or U821 (N_821,In_871,In_288);
and U822 (N_822,In_362,In_927);
nand U823 (N_823,In_357,In_751);
or U824 (N_824,In_137,In_569);
nor U825 (N_825,In_659,In_936);
or U826 (N_826,In_643,In_658);
and U827 (N_827,In_99,In_710);
nand U828 (N_828,In_873,In_628);
and U829 (N_829,In_699,In_183);
and U830 (N_830,In_448,In_518);
nand U831 (N_831,In_484,In_32);
and U832 (N_832,In_847,In_916);
and U833 (N_833,In_354,In_282);
or U834 (N_834,In_412,In_856);
or U835 (N_835,In_121,In_702);
nand U836 (N_836,In_976,In_43);
nand U837 (N_837,In_116,In_773);
nand U838 (N_838,In_959,In_881);
or U839 (N_839,In_1,In_433);
xnor U840 (N_840,In_16,In_538);
and U841 (N_841,In_99,In_387);
or U842 (N_842,In_188,In_47);
nand U843 (N_843,In_922,In_860);
xor U844 (N_844,In_274,In_215);
or U845 (N_845,In_928,In_106);
and U846 (N_846,In_778,In_737);
or U847 (N_847,In_567,In_568);
or U848 (N_848,In_956,In_546);
and U849 (N_849,In_610,In_952);
or U850 (N_850,In_593,In_344);
or U851 (N_851,In_560,In_447);
and U852 (N_852,In_860,In_385);
nor U853 (N_853,In_944,In_45);
nand U854 (N_854,In_372,In_39);
nor U855 (N_855,In_744,In_178);
and U856 (N_856,In_377,In_677);
or U857 (N_857,In_72,In_142);
nand U858 (N_858,In_666,In_821);
nand U859 (N_859,In_105,In_383);
and U860 (N_860,In_738,In_110);
nand U861 (N_861,In_832,In_246);
or U862 (N_862,In_588,In_20);
nor U863 (N_863,In_703,In_825);
and U864 (N_864,In_929,In_337);
nor U865 (N_865,In_949,In_358);
nand U866 (N_866,In_237,In_257);
or U867 (N_867,In_320,In_380);
and U868 (N_868,In_171,In_915);
xor U869 (N_869,In_814,In_154);
nor U870 (N_870,In_844,In_218);
nor U871 (N_871,In_495,In_892);
nand U872 (N_872,In_42,In_93);
nor U873 (N_873,In_186,In_132);
or U874 (N_874,In_304,In_386);
or U875 (N_875,In_635,In_259);
nand U876 (N_876,In_300,In_410);
or U877 (N_877,In_191,In_207);
nor U878 (N_878,In_976,In_515);
nand U879 (N_879,In_4,In_140);
or U880 (N_880,In_458,In_962);
or U881 (N_881,In_133,In_959);
or U882 (N_882,In_234,In_685);
nor U883 (N_883,In_926,In_493);
xnor U884 (N_884,In_978,In_359);
and U885 (N_885,In_383,In_432);
xor U886 (N_886,In_441,In_908);
or U887 (N_887,In_842,In_782);
or U888 (N_888,In_562,In_501);
xnor U889 (N_889,In_407,In_897);
and U890 (N_890,In_907,In_827);
xnor U891 (N_891,In_447,In_450);
and U892 (N_892,In_348,In_845);
nand U893 (N_893,In_415,In_335);
or U894 (N_894,In_580,In_666);
nor U895 (N_895,In_554,In_966);
or U896 (N_896,In_409,In_119);
and U897 (N_897,In_417,In_429);
nor U898 (N_898,In_472,In_595);
and U899 (N_899,In_58,In_422);
and U900 (N_900,In_557,In_830);
nor U901 (N_901,In_142,In_740);
and U902 (N_902,In_895,In_116);
or U903 (N_903,In_382,In_630);
nand U904 (N_904,In_734,In_626);
nand U905 (N_905,In_404,In_357);
or U906 (N_906,In_177,In_146);
xor U907 (N_907,In_446,In_695);
nor U908 (N_908,In_843,In_598);
and U909 (N_909,In_636,In_539);
nor U910 (N_910,In_757,In_726);
or U911 (N_911,In_752,In_6);
xnor U912 (N_912,In_483,In_455);
or U913 (N_913,In_227,In_358);
nor U914 (N_914,In_890,In_162);
nor U915 (N_915,In_852,In_453);
nand U916 (N_916,In_780,In_284);
or U917 (N_917,In_129,In_343);
nor U918 (N_918,In_898,In_146);
nand U919 (N_919,In_809,In_819);
nor U920 (N_920,In_243,In_207);
and U921 (N_921,In_662,In_8);
nor U922 (N_922,In_235,In_668);
or U923 (N_923,In_54,In_616);
nand U924 (N_924,In_448,In_87);
nand U925 (N_925,In_469,In_634);
and U926 (N_926,In_950,In_257);
nor U927 (N_927,In_608,In_190);
or U928 (N_928,In_546,In_411);
nor U929 (N_929,In_472,In_164);
or U930 (N_930,In_66,In_233);
or U931 (N_931,In_272,In_263);
nand U932 (N_932,In_966,In_79);
or U933 (N_933,In_212,In_282);
nor U934 (N_934,In_177,In_498);
and U935 (N_935,In_658,In_142);
nor U936 (N_936,In_45,In_835);
and U937 (N_937,In_750,In_798);
and U938 (N_938,In_626,In_748);
nand U939 (N_939,In_962,In_138);
or U940 (N_940,In_301,In_925);
nor U941 (N_941,In_69,In_146);
nand U942 (N_942,In_615,In_30);
nand U943 (N_943,In_296,In_14);
or U944 (N_944,In_488,In_326);
nor U945 (N_945,In_105,In_744);
nand U946 (N_946,In_381,In_113);
nor U947 (N_947,In_201,In_723);
nor U948 (N_948,In_263,In_664);
nand U949 (N_949,In_804,In_290);
nand U950 (N_950,In_236,In_830);
nor U951 (N_951,In_367,In_565);
nand U952 (N_952,In_808,In_132);
and U953 (N_953,In_373,In_930);
or U954 (N_954,In_883,In_429);
nand U955 (N_955,In_739,In_531);
nor U956 (N_956,In_984,In_843);
and U957 (N_957,In_157,In_366);
or U958 (N_958,In_97,In_317);
xor U959 (N_959,In_853,In_902);
nor U960 (N_960,In_248,In_646);
nor U961 (N_961,In_915,In_494);
xor U962 (N_962,In_924,In_996);
nor U963 (N_963,In_511,In_290);
or U964 (N_964,In_553,In_747);
and U965 (N_965,In_940,In_6);
nand U966 (N_966,In_292,In_695);
and U967 (N_967,In_941,In_754);
and U968 (N_968,In_903,In_643);
or U969 (N_969,In_339,In_508);
nor U970 (N_970,In_912,In_941);
or U971 (N_971,In_263,In_310);
and U972 (N_972,In_391,In_135);
nor U973 (N_973,In_849,In_631);
and U974 (N_974,In_713,In_781);
or U975 (N_975,In_180,In_454);
nor U976 (N_976,In_831,In_550);
and U977 (N_977,In_717,In_422);
nand U978 (N_978,In_287,In_19);
or U979 (N_979,In_116,In_618);
xnor U980 (N_980,In_450,In_401);
nand U981 (N_981,In_930,In_981);
and U982 (N_982,In_896,In_276);
nor U983 (N_983,In_651,In_975);
nor U984 (N_984,In_861,In_226);
xnor U985 (N_985,In_851,In_248);
nor U986 (N_986,In_254,In_517);
nor U987 (N_987,In_760,In_850);
nor U988 (N_988,In_739,In_569);
and U989 (N_989,In_842,In_107);
nand U990 (N_990,In_993,In_123);
and U991 (N_991,In_14,In_425);
and U992 (N_992,In_328,In_51);
and U993 (N_993,In_205,In_864);
or U994 (N_994,In_923,In_204);
and U995 (N_995,In_250,In_352);
xor U996 (N_996,In_250,In_409);
and U997 (N_997,In_40,In_179);
or U998 (N_998,In_977,In_602);
and U999 (N_999,In_636,In_0);
and U1000 (N_1000,In_107,In_981);
nand U1001 (N_1001,In_963,In_740);
and U1002 (N_1002,In_216,In_560);
nor U1003 (N_1003,In_739,In_767);
nand U1004 (N_1004,In_748,In_136);
xnor U1005 (N_1005,In_803,In_973);
and U1006 (N_1006,In_272,In_512);
and U1007 (N_1007,In_935,In_533);
or U1008 (N_1008,In_11,In_183);
nor U1009 (N_1009,In_712,In_720);
nor U1010 (N_1010,In_730,In_647);
or U1011 (N_1011,In_233,In_603);
or U1012 (N_1012,In_572,In_291);
nor U1013 (N_1013,In_643,In_380);
and U1014 (N_1014,In_663,In_332);
nor U1015 (N_1015,In_31,In_535);
or U1016 (N_1016,In_170,In_494);
nand U1017 (N_1017,In_136,In_938);
and U1018 (N_1018,In_490,In_755);
nand U1019 (N_1019,In_61,In_31);
and U1020 (N_1020,In_79,In_97);
xnor U1021 (N_1021,In_994,In_811);
nor U1022 (N_1022,In_269,In_761);
nand U1023 (N_1023,In_600,In_803);
nand U1024 (N_1024,In_975,In_681);
nand U1025 (N_1025,In_246,In_943);
nand U1026 (N_1026,In_237,In_880);
and U1027 (N_1027,In_701,In_533);
or U1028 (N_1028,In_889,In_110);
nand U1029 (N_1029,In_168,In_761);
and U1030 (N_1030,In_986,In_947);
nand U1031 (N_1031,In_981,In_636);
xor U1032 (N_1032,In_597,In_533);
and U1033 (N_1033,In_455,In_480);
xnor U1034 (N_1034,In_95,In_772);
nand U1035 (N_1035,In_514,In_303);
or U1036 (N_1036,In_318,In_608);
and U1037 (N_1037,In_732,In_432);
nand U1038 (N_1038,In_868,In_103);
nor U1039 (N_1039,In_420,In_728);
nor U1040 (N_1040,In_793,In_374);
nor U1041 (N_1041,In_459,In_219);
xnor U1042 (N_1042,In_298,In_392);
or U1043 (N_1043,In_697,In_301);
nor U1044 (N_1044,In_311,In_39);
nand U1045 (N_1045,In_288,In_375);
or U1046 (N_1046,In_440,In_756);
or U1047 (N_1047,In_785,In_261);
and U1048 (N_1048,In_586,In_267);
nor U1049 (N_1049,In_79,In_137);
nor U1050 (N_1050,In_447,In_536);
nor U1051 (N_1051,In_842,In_49);
or U1052 (N_1052,In_323,In_612);
or U1053 (N_1053,In_607,In_833);
nor U1054 (N_1054,In_674,In_366);
nand U1055 (N_1055,In_407,In_3);
xnor U1056 (N_1056,In_980,In_28);
nand U1057 (N_1057,In_607,In_162);
nor U1058 (N_1058,In_365,In_551);
or U1059 (N_1059,In_923,In_981);
nand U1060 (N_1060,In_418,In_105);
or U1061 (N_1061,In_869,In_826);
nand U1062 (N_1062,In_700,In_332);
xnor U1063 (N_1063,In_224,In_707);
nand U1064 (N_1064,In_929,In_261);
or U1065 (N_1065,In_486,In_696);
and U1066 (N_1066,In_695,In_997);
nor U1067 (N_1067,In_26,In_590);
nand U1068 (N_1068,In_863,In_69);
nor U1069 (N_1069,In_59,In_43);
nor U1070 (N_1070,In_225,In_974);
or U1071 (N_1071,In_150,In_527);
nand U1072 (N_1072,In_404,In_914);
nor U1073 (N_1073,In_191,In_99);
xnor U1074 (N_1074,In_932,In_987);
nand U1075 (N_1075,In_833,In_166);
nor U1076 (N_1076,In_863,In_848);
or U1077 (N_1077,In_346,In_116);
or U1078 (N_1078,In_826,In_559);
nor U1079 (N_1079,In_223,In_409);
and U1080 (N_1080,In_521,In_485);
nand U1081 (N_1081,In_933,In_188);
nor U1082 (N_1082,In_285,In_424);
nor U1083 (N_1083,In_496,In_4);
nor U1084 (N_1084,In_463,In_687);
and U1085 (N_1085,In_26,In_184);
nor U1086 (N_1086,In_129,In_900);
nor U1087 (N_1087,In_372,In_411);
or U1088 (N_1088,In_987,In_11);
nor U1089 (N_1089,In_63,In_749);
or U1090 (N_1090,In_797,In_238);
nor U1091 (N_1091,In_302,In_718);
nand U1092 (N_1092,In_91,In_828);
or U1093 (N_1093,In_557,In_236);
nand U1094 (N_1094,In_109,In_798);
and U1095 (N_1095,In_825,In_830);
and U1096 (N_1096,In_143,In_308);
nor U1097 (N_1097,In_655,In_482);
xor U1098 (N_1098,In_634,In_539);
nor U1099 (N_1099,In_186,In_504);
and U1100 (N_1100,In_185,In_823);
or U1101 (N_1101,In_746,In_904);
and U1102 (N_1102,In_304,In_824);
nand U1103 (N_1103,In_987,In_520);
nand U1104 (N_1104,In_840,In_904);
and U1105 (N_1105,In_708,In_949);
or U1106 (N_1106,In_509,In_902);
nand U1107 (N_1107,In_385,In_957);
or U1108 (N_1108,In_359,In_771);
and U1109 (N_1109,In_278,In_379);
and U1110 (N_1110,In_706,In_459);
nand U1111 (N_1111,In_433,In_204);
nand U1112 (N_1112,In_373,In_11);
nor U1113 (N_1113,In_885,In_805);
xnor U1114 (N_1114,In_476,In_209);
or U1115 (N_1115,In_309,In_417);
nor U1116 (N_1116,In_709,In_986);
nand U1117 (N_1117,In_865,In_124);
nor U1118 (N_1118,In_58,In_496);
nor U1119 (N_1119,In_850,In_362);
and U1120 (N_1120,In_701,In_139);
nand U1121 (N_1121,In_748,In_226);
nand U1122 (N_1122,In_123,In_501);
nand U1123 (N_1123,In_76,In_143);
xnor U1124 (N_1124,In_713,In_79);
or U1125 (N_1125,In_830,In_169);
xor U1126 (N_1126,In_975,In_393);
nor U1127 (N_1127,In_474,In_295);
and U1128 (N_1128,In_772,In_636);
or U1129 (N_1129,In_734,In_975);
and U1130 (N_1130,In_756,In_229);
and U1131 (N_1131,In_183,In_608);
or U1132 (N_1132,In_236,In_651);
or U1133 (N_1133,In_963,In_470);
nand U1134 (N_1134,In_897,In_597);
and U1135 (N_1135,In_682,In_205);
nor U1136 (N_1136,In_106,In_207);
nor U1137 (N_1137,In_487,In_695);
or U1138 (N_1138,In_540,In_272);
nand U1139 (N_1139,In_408,In_18);
nor U1140 (N_1140,In_612,In_213);
nor U1141 (N_1141,In_471,In_955);
nand U1142 (N_1142,In_618,In_433);
or U1143 (N_1143,In_866,In_983);
and U1144 (N_1144,In_29,In_417);
nor U1145 (N_1145,In_137,In_859);
nor U1146 (N_1146,In_392,In_57);
or U1147 (N_1147,In_700,In_109);
nor U1148 (N_1148,In_330,In_761);
or U1149 (N_1149,In_523,In_951);
and U1150 (N_1150,In_839,In_445);
or U1151 (N_1151,In_755,In_984);
nand U1152 (N_1152,In_230,In_251);
xnor U1153 (N_1153,In_349,In_862);
nand U1154 (N_1154,In_985,In_237);
nand U1155 (N_1155,In_682,In_922);
and U1156 (N_1156,In_985,In_998);
nand U1157 (N_1157,In_248,In_25);
or U1158 (N_1158,In_740,In_509);
xnor U1159 (N_1159,In_229,In_480);
or U1160 (N_1160,In_89,In_323);
nand U1161 (N_1161,In_511,In_49);
nor U1162 (N_1162,In_484,In_294);
nor U1163 (N_1163,In_463,In_752);
nor U1164 (N_1164,In_362,In_291);
xor U1165 (N_1165,In_214,In_689);
and U1166 (N_1166,In_523,In_654);
and U1167 (N_1167,In_382,In_216);
nand U1168 (N_1168,In_632,In_842);
and U1169 (N_1169,In_989,In_328);
nand U1170 (N_1170,In_73,In_644);
or U1171 (N_1171,In_661,In_769);
nor U1172 (N_1172,In_191,In_812);
or U1173 (N_1173,In_44,In_165);
nand U1174 (N_1174,In_821,In_770);
or U1175 (N_1175,In_673,In_426);
nand U1176 (N_1176,In_758,In_939);
nand U1177 (N_1177,In_469,In_263);
and U1178 (N_1178,In_890,In_384);
or U1179 (N_1179,In_913,In_644);
and U1180 (N_1180,In_420,In_331);
nor U1181 (N_1181,In_693,In_24);
or U1182 (N_1182,In_11,In_884);
xor U1183 (N_1183,In_476,In_904);
xnor U1184 (N_1184,In_437,In_371);
and U1185 (N_1185,In_745,In_136);
and U1186 (N_1186,In_415,In_658);
and U1187 (N_1187,In_536,In_205);
nand U1188 (N_1188,In_909,In_630);
nand U1189 (N_1189,In_951,In_920);
and U1190 (N_1190,In_397,In_503);
nand U1191 (N_1191,In_722,In_697);
nor U1192 (N_1192,In_864,In_679);
and U1193 (N_1193,In_23,In_458);
and U1194 (N_1194,In_950,In_902);
nor U1195 (N_1195,In_336,In_832);
nand U1196 (N_1196,In_437,In_948);
or U1197 (N_1197,In_490,In_625);
or U1198 (N_1198,In_538,In_104);
nand U1199 (N_1199,In_316,In_712);
nand U1200 (N_1200,In_709,In_480);
nand U1201 (N_1201,In_713,In_168);
or U1202 (N_1202,In_440,In_498);
nand U1203 (N_1203,In_232,In_514);
nor U1204 (N_1204,In_340,In_805);
and U1205 (N_1205,In_660,In_323);
xnor U1206 (N_1206,In_34,In_805);
or U1207 (N_1207,In_253,In_434);
or U1208 (N_1208,In_193,In_901);
nor U1209 (N_1209,In_618,In_781);
nor U1210 (N_1210,In_470,In_835);
or U1211 (N_1211,In_151,In_107);
or U1212 (N_1212,In_748,In_683);
nor U1213 (N_1213,In_878,In_719);
xnor U1214 (N_1214,In_190,In_520);
or U1215 (N_1215,In_712,In_184);
or U1216 (N_1216,In_821,In_985);
and U1217 (N_1217,In_91,In_124);
nor U1218 (N_1218,In_498,In_669);
or U1219 (N_1219,In_301,In_55);
and U1220 (N_1220,In_382,In_829);
nor U1221 (N_1221,In_557,In_487);
and U1222 (N_1222,In_676,In_67);
and U1223 (N_1223,In_348,In_699);
or U1224 (N_1224,In_486,In_498);
xnor U1225 (N_1225,In_696,In_381);
or U1226 (N_1226,In_933,In_621);
xor U1227 (N_1227,In_220,In_99);
or U1228 (N_1228,In_523,In_745);
nand U1229 (N_1229,In_217,In_208);
nor U1230 (N_1230,In_862,In_715);
or U1231 (N_1231,In_831,In_755);
and U1232 (N_1232,In_899,In_528);
nor U1233 (N_1233,In_314,In_434);
nand U1234 (N_1234,In_2,In_250);
and U1235 (N_1235,In_217,In_10);
or U1236 (N_1236,In_190,In_686);
nand U1237 (N_1237,In_988,In_855);
or U1238 (N_1238,In_777,In_971);
or U1239 (N_1239,In_102,In_768);
nand U1240 (N_1240,In_857,In_161);
xnor U1241 (N_1241,In_124,In_146);
and U1242 (N_1242,In_547,In_550);
or U1243 (N_1243,In_260,In_38);
nor U1244 (N_1244,In_555,In_868);
or U1245 (N_1245,In_733,In_617);
or U1246 (N_1246,In_473,In_395);
nand U1247 (N_1247,In_445,In_48);
nand U1248 (N_1248,In_737,In_750);
nand U1249 (N_1249,In_11,In_856);
and U1250 (N_1250,In_854,In_501);
and U1251 (N_1251,In_924,In_512);
and U1252 (N_1252,In_678,In_592);
or U1253 (N_1253,In_152,In_671);
or U1254 (N_1254,In_51,In_172);
or U1255 (N_1255,In_776,In_70);
or U1256 (N_1256,In_777,In_198);
and U1257 (N_1257,In_265,In_234);
or U1258 (N_1258,In_772,In_267);
nand U1259 (N_1259,In_542,In_762);
or U1260 (N_1260,In_849,In_9);
nor U1261 (N_1261,In_566,In_558);
nand U1262 (N_1262,In_449,In_174);
and U1263 (N_1263,In_39,In_168);
or U1264 (N_1264,In_269,In_621);
or U1265 (N_1265,In_798,In_316);
or U1266 (N_1266,In_612,In_678);
or U1267 (N_1267,In_761,In_713);
and U1268 (N_1268,In_258,In_431);
nand U1269 (N_1269,In_157,In_511);
or U1270 (N_1270,In_523,In_485);
and U1271 (N_1271,In_94,In_521);
and U1272 (N_1272,In_973,In_607);
nor U1273 (N_1273,In_730,In_109);
or U1274 (N_1274,In_573,In_454);
nor U1275 (N_1275,In_553,In_299);
nand U1276 (N_1276,In_598,In_175);
and U1277 (N_1277,In_468,In_476);
or U1278 (N_1278,In_975,In_69);
and U1279 (N_1279,In_992,In_792);
or U1280 (N_1280,In_367,In_201);
nor U1281 (N_1281,In_774,In_780);
nand U1282 (N_1282,In_228,In_382);
nand U1283 (N_1283,In_122,In_540);
xor U1284 (N_1284,In_242,In_224);
nand U1285 (N_1285,In_596,In_133);
or U1286 (N_1286,In_475,In_336);
nor U1287 (N_1287,In_842,In_613);
or U1288 (N_1288,In_331,In_71);
or U1289 (N_1289,In_593,In_594);
and U1290 (N_1290,In_991,In_94);
and U1291 (N_1291,In_727,In_16);
and U1292 (N_1292,In_690,In_12);
or U1293 (N_1293,In_748,In_298);
or U1294 (N_1294,In_13,In_158);
xor U1295 (N_1295,In_395,In_284);
or U1296 (N_1296,In_462,In_248);
and U1297 (N_1297,In_72,In_885);
nor U1298 (N_1298,In_400,In_642);
xor U1299 (N_1299,In_624,In_439);
xnor U1300 (N_1300,In_571,In_992);
nor U1301 (N_1301,In_379,In_727);
nor U1302 (N_1302,In_682,In_355);
nand U1303 (N_1303,In_109,In_310);
nand U1304 (N_1304,In_78,In_954);
and U1305 (N_1305,In_496,In_79);
xor U1306 (N_1306,In_534,In_813);
nand U1307 (N_1307,In_184,In_327);
nor U1308 (N_1308,In_528,In_249);
nand U1309 (N_1309,In_158,In_326);
or U1310 (N_1310,In_619,In_73);
or U1311 (N_1311,In_632,In_184);
or U1312 (N_1312,In_79,In_897);
or U1313 (N_1313,In_422,In_463);
or U1314 (N_1314,In_116,In_709);
xnor U1315 (N_1315,In_179,In_646);
or U1316 (N_1316,In_458,In_270);
or U1317 (N_1317,In_854,In_93);
or U1318 (N_1318,In_806,In_941);
xor U1319 (N_1319,In_583,In_660);
or U1320 (N_1320,In_274,In_718);
and U1321 (N_1321,In_768,In_438);
or U1322 (N_1322,In_475,In_513);
nand U1323 (N_1323,In_533,In_518);
and U1324 (N_1324,In_632,In_393);
and U1325 (N_1325,In_123,In_675);
or U1326 (N_1326,In_141,In_899);
nor U1327 (N_1327,In_732,In_656);
and U1328 (N_1328,In_595,In_806);
or U1329 (N_1329,In_397,In_182);
xor U1330 (N_1330,In_626,In_647);
and U1331 (N_1331,In_736,In_565);
and U1332 (N_1332,In_432,In_249);
or U1333 (N_1333,In_838,In_12);
and U1334 (N_1334,In_493,In_58);
nand U1335 (N_1335,In_663,In_112);
or U1336 (N_1336,In_396,In_109);
nor U1337 (N_1337,In_380,In_319);
or U1338 (N_1338,In_777,In_417);
or U1339 (N_1339,In_644,In_322);
or U1340 (N_1340,In_33,In_639);
nand U1341 (N_1341,In_995,In_742);
nor U1342 (N_1342,In_410,In_836);
nand U1343 (N_1343,In_771,In_207);
or U1344 (N_1344,In_30,In_328);
nor U1345 (N_1345,In_38,In_640);
or U1346 (N_1346,In_605,In_766);
nand U1347 (N_1347,In_335,In_111);
or U1348 (N_1348,In_562,In_672);
nand U1349 (N_1349,In_585,In_346);
and U1350 (N_1350,In_688,In_616);
nand U1351 (N_1351,In_843,In_432);
nand U1352 (N_1352,In_441,In_635);
nand U1353 (N_1353,In_284,In_19);
nor U1354 (N_1354,In_662,In_533);
xnor U1355 (N_1355,In_613,In_533);
xor U1356 (N_1356,In_96,In_255);
xnor U1357 (N_1357,In_113,In_734);
xor U1358 (N_1358,In_506,In_567);
nor U1359 (N_1359,In_358,In_549);
and U1360 (N_1360,In_628,In_468);
nand U1361 (N_1361,In_806,In_952);
or U1362 (N_1362,In_530,In_474);
nand U1363 (N_1363,In_108,In_637);
nand U1364 (N_1364,In_738,In_918);
or U1365 (N_1365,In_808,In_718);
nand U1366 (N_1366,In_550,In_894);
or U1367 (N_1367,In_567,In_279);
xor U1368 (N_1368,In_727,In_403);
nand U1369 (N_1369,In_13,In_152);
xnor U1370 (N_1370,In_426,In_729);
nor U1371 (N_1371,In_129,In_823);
and U1372 (N_1372,In_893,In_360);
and U1373 (N_1373,In_73,In_613);
and U1374 (N_1374,In_301,In_519);
nand U1375 (N_1375,In_948,In_800);
xnor U1376 (N_1376,In_813,In_927);
and U1377 (N_1377,In_130,In_74);
nor U1378 (N_1378,In_630,In_944);
and U1379 (N_1379,In_294,In_914);
nand U1380 (N_1380,In_905,In_268);
or U1381 (N_1381,In_278,In_441);
nor U1382 (N_1382,In_737,In_551);
nor U1383 (N_1383,In_169,In_730);
or U1384 (N_1384,In_609,In_17);
nand U1385 (N_1385,In_285,In_161);
and U1386 (N_1386,In_963,In_349);
nor U1387 (N_1387,In_57,In_962);
nand U1388 (N_1388,In_209,In_464);
or U1389 (N_1389,In_955,In_254);
nor U1390 (N_1390,In_636,In_74);
or U1391 (N_1391,In_134,In_456);
nand U1392 (N_1392,In_227,In_669);
xor U1393 (N_1393,In_919,In_803);
and U1394 (N_1394,In_230,In_664);
or U1395 (N_1395,In_161,In_27);
and U1396 (N_1396,In_627,In_479);
nand U1397 (N_1397,In_235,In_413);
and U1398 (N_1398,In_538,In_29);
nor U1399 (N_1399,In_154,In_593);
and U1400 (N_1400,In_959,In_737);
nor U1401 (N_1401,In_98,In_661);
or U1402 (N_1402,In_538,In_91);
and U1403 (N_1403,In_670,In_444);
or U1404 (N_1404,In_322,In_23);
and U1405 (N_1405,In_261,In_722);
and U1406 (N_1406,In_15,In_475);
or U1407 (N_1407,In_884,In_712);
nand U1408 (N_1408,In_481,In_417);
and U1409 (N_1409,In_970,In_761);
nor U1410 (N_1410,In_345,In_184);
and U1411 (N_1411,In_956,In_69);
nand U1412 (N_1412,In_16,In_752);
or U1413 (N_1413,In_800,In_592);
nor U1414 (N_1414,In_957,In_906);
xnor U1415 (N_1415,In_467,In_116);
or U1416 (N_1416,In_773,In_520);
and U1417 (N_1417,In_776,In_846);
or U1418 (N_1418,In_96,In_639);
nor U1419 (N_1419,In_807,In_833);
nor U1420 (N_1420,In_465,In_649);
and U1421 (N_1421,In_146,In_187);
nor U1422 (N_1422,In_125,In_664);
or U1423 (N_1423,In_769,In_160);
and U1424 (N_1424,In_698,In_453);
nand U1425 (N_1425,In_451,In_394);
or U1426 (N_1426,In_987,In_499);
and U1427 (N_1427,In_694,In_877);
and U1428 (N_1428,In_276,In_605);
and U1429 (N_1429,In_800,In_246);
or U1430 (N_1430,In_144,In_607);
nand U1431 (N_1431,In_669,In_372);
nand U1432 (N_1432,In_368,In_454);
nand U1433 (N_1433,In_197,In_462);
nand U1434 (N_1434,In_512,In_812);
nor U1435 (N_1435,In_914,In_895);
nor U1436 (N_1436,In_577,In_444);
or U1437 (N_1437,In_357,In_356);
nor U1438 (N_1438,In_660,In_655);
xnor U1439 (N_1439,In_405,In_209);
or U1440 (N_1440,In_829,In_635);
and U1441 (N_1441,In_184,In_365);
or U1442 (N_1442,In_317,In_364);
nand U1443 (N_1443,In_996,In_27);
nor U1444 (N_1444,In_832,In_6);
nor U1445 (N_1445,In_721,In_982);
xor U1446 (N_1446,In_717,In_153);
nand U1447 (N_1447,In_763,In_9);
or U1448 (N_1448,In_774,In_618);
nor U1449 (N_1449,In_107,In_1);
nor U1450 (N_1450,In_443,In_567);
and U1451 (N_1451,In_435,In_909);
and U1452 (N_1452,In_136,In_527);
nand U1453 (N_1453,In_168,In_148);
nor U1454 (N_1454,In_598,In_530);
or U1455 (N_1455,In_715,In_858);
and U1456 (N_1456,In_835,In_611);
nor U1457 (N_1457,In_452,In_927);
nand U1458 (N_1458,In_738,In_704);
nor U1459 (N_1459,In_191,In_50);
xnor U1460 (N_1460,In_947,In_704);
nand U1461 (N_1461,In_474,In_668);
or U1462 (N_1462,In_817,In_710);
xor U1463 (N_1463,In_270,In_859);
nand U1464 (N_1464,In_175,In_995);
nand U1465 (N_1465,In_805,In_788);
or U1466 (N_1466,In_632,In_558);
or U1467 (N_1467,In_897,In_828);
nand U1468 (N_1468,In_857,In_519);
or U1469 (N_1469,In_285,In_532);
or U1470 (N_1470,In_279,In_537);
and U1471 (N_1471,In_364,In_540);
nand U1472 (N_1472,In_953,In_275);
and U1473 (N_1473,In_575,In_915);
nor U1474 (N_1474,In_597,In_258);
nor U1475 (N_1475,In_195,In_88);
and U1476 (N_1476,In_105,In_230);
or U1477 (N_1477,In_554,In_342);
nor U1478 (N_1478,In_644,In_330);
or U1479 (N_1479,In_264,In_182);
nor U1480 (N_1480,In_547,In_309);
and U1481 (N_1481,In_36,In_720);
or U1482 (N_1482,In_519,In_930);
xnor U1483 (N_1483,In_774,In_244);
nand U1484 (N_1484,In_274,In_987);
xnor U1485 (N_1485,In_14,In_496);
or U1486 (N_1486,In_98,In_137);
or U1487 (N_1487,In_195,In_153);
nand U1488 (N_1488,In_786,In_476);
xor U1489 (N_1489,In_22,In_583);
xor U1490 (N_1490,In_849,In_669);
nor U1491 (N_1491,In_112,In_85);
and U1492 (N_1492,In_46,In_586);
nor U1493 (N_1493,In_115,In_655);
or U1494 (N_1494,In_628,In_495);
and U1495 (N_1495,In_966,In_924);
or U1496 (N_1496,In_949,In_139);
nor U1497 (N_1497,In_886,In_100);
xnor U1498 (N_1498,In_846,In_837);
and U1499 (N_1499,In_199,In_725);
nor U1500 (N_1500,In_486,In_593);
nor U1501 (N_1501,In_570,In_324);
or U1502 (N_1502,In_718,In_945);
or U1503 (N_1503,In_350,In_584);
or U1504 (N_1504,In_648,In_796);
nor U1505 (N_1505,In_317,In_41);
nor U1506 (N_1506,In_524,In_899);
and U1507 (N_1507,In_317,In_400);
nor U1508 (N_1508,In_723,In_614);
or U1509 (N_1509,In_739,In_272);
or U1510 (N_1510,In_418,In_515);
nand U1511 (N_1511,In_490,In_330);
nand U1512 (N_1512,In_157,In_739);
nand U1513 (N_1513,In_765,In_386);
xnor U1514 (N_1514,In_982,In_333);
xor U1515 (N_1515,In_381,In_291);
nand U1516 (N_1516,In_359,In_113);
xor U1517 (N_1517,In_784,In_224);
nor U1518 (N_1518,In_579,In_969);
or U1519 (N_1519,In_704,In_129);
or U1520 (N_1520,In_771,In_561);
nand U1521 (N_1521,In_463,In_513);
nand U1522 (N_1522,In_865,In_609);
and U1523 (N_1523,In_404,In_329);
or U1524 (N_1524,In_209,In_256);
nand U1525 (N_1525,In_844,In_514);
or U1526 (N_1526,In_159,In_418);
nor U1527 (N_1527,In_298,In_122);
or U1528 (N_1528,In_386,In_840);
and U1529 (N_1529,In_822,In_761);
and U1530 (N_1530,In_871,In_557);
or U1531 (N_1531,In_152,In_516);
nand U1532 (N_1532,In_564,In_748);
nor U1533 (N_1533,In_666,In_294);
nor U1534 (N_1534,In_136,In_763);
xnor U1535 (N_1535,In_762,In_47);
or U1536 (N_1536,In_609,In_176);
or U1537 (N_1537,In_461,In_565);
nand U1538 (N_1538,In_205,In_492);
nor U1539 (N_1539,In_373,In_924);
nor U1540 (N_1540,In_258,In_947);
nor U1541 (N_1541,In_388,In_590);
nand U1542 (N_1542,In_657,In_551);
nor U1543 (N_1543,In_311,In_905);
and U1544 (N_1544,In_403,In_312);
nor U1545 (N_1545,In_95,In_941);
nand U1546 (N_1546,In_540,In_230);
nor U1547 (N_1547,In_262,In_239);
or U1548 (N_1548,In_293,In_627);
nor U1549 (N_1549,In_621,In_970);
or U1550 (N_1550,In_390,In_693);
and U1551 (N_1551,In_95,In_894);
nor U1552 (N_1552,In_464,In_359);
nor U1553 (N_1553,In_652,In_593);
nor U1554 (N_1554,In_204,In_456);
and U1555 (N_1555,In_825,In_523);
nand U1556 (N_1556,In_757,In_313);
and U1557 (N_1557,In_68,In_307);
and U1558 (N_1558,In_374,In_338);
or U1559 (N_1559,In_987,In_991);
nor U1560 (N_1560,In_141,In_2);
nand U1561 (N_1561,In_215,In_241);
nand U1562 (N_1562,In_818,In_106);
nand U1563 (N_1563,In_483,In_334);
nand U1564 (N_1564,In_602,In_814);
nor U1565 (N_1565,In_712,In_804);
or U1566 (N_1566,In_170,In_285);
nand U1567 (N_1567,In_170,In_986);
nor U1568 (N_1568,In_137,In_26);
nor U1569 (N_1569,In_624,In_592);
and U1570 (N_1570,In_963,In_311);
nor U1571 (N_1571,In_600,In_898);
nand U1572 (N_1572,In_144,In_321);
or U1573 (N_1573,In_118,In_129);
nor U1574 (N_1574,In_319,In_588);
nand U1575 (N_1575,In_0,In_114);
nand U1576 (N_1576,In_105,In_207);
nand U1577 (N_1577,In_405,In_501);
and U1578 (N_1578,In_18,In_572);
and U1579 (N_1579,In_372,In_59);
nand U1580 (N_1580,In_616,In_171);
nor U1581 (N_1581,In_357,In_702);
nand U1582 (N_1582,In_808,In_147);
nor U1583 (N_1583,In_111,In_853);
nor U1584 (N_1584,In_297,In_563);
xor U1585 (N_1585,In_610,In_893);
or U1586 (N_1586,In_792,In_512);
and U1587 (N_1587,In_936,In_435);
and U1588 (N_1588,In_220,In_325);
nor U1589 (N_1589,In_414,In_31);
and U1590 (N_1590,In_722,In_371);
xnor U1591 (N_1591,In_758,In_851);
or U1592 (N_1592,In_556,In_50);
nor U1593 (N_1593,In_926,In_951);
nor U1594 (N_1594,In_288,In_620);
nor U1595 (N_1595,In_424,In_944);
nor U1596 (N_1596,In_451,In_466);
or U1597 (N_1597,In_262,In_586);
and U1598 (N_1598,In_392,In_619);
xor U1599 (N_1599,In_685,In_405);
or U1600 (N_1600,In_475,In_558);
nor U1601 (N_1601,In_159,In_968);
or U1602 (N_1602,In_448,In_523);
or U1603 (N_1603,In_578,In_549);
or U1604 (N_1604,In_467,In_233);
and U1605 (N_1605,In_350,In_837);
or U1606 (N_1606,In_733,In_176);
or U1607 (N_1607,In_892,In_326);
and U1608 (N_1608,In_897,In_298);
nor U1609 (N_1609,In_3,In_846);
nor U1610 (N_1610,In_896,In_261);
and U1611 (N_1611,In_836,In_112);
nand U1612 (N_1612,In_141,In_727);
nor U1613 (N_1613,In_367,In_746);
nand U1614 (N_1614,In_972,In_931);
and U1615 (N_1615,In_82,In_684);
nand U1616 (N_1616,In_239,In_645);
nor U1617 (N_1617,In_653,In_770);
nor U1618 (N_1618,In_414,In_506);
nor U1619 (N_1619,In_218,In_813);
and U1620 (N_1620,In_360,In_177);
nor U1621 (N_1621,In_200,In_270);
nor U1622 (N_1622,In_468,In_561);
nor U1623 (N_1623,In_74,In_913);
or U1624 (N_1624,In_691,In_393);
nand U1625 (N_1625,In_165,In_527);
and U1626 (N_1626,In_405,In_470);
xor U1627 (N_1627,In_588,In_138);
nor U1628 (N_1628,In_846,In_352);
nor U1629 (N_1629,In_237,In_722);
or U1630 (N_1630,In_847,In_515);
or U1631 (N_1631,In_0,In_354);
nor U1632 (N_1632,In_599,In_866);
or U1633 (N_1633,In_871,In_733);
nor U1634 (N_1634,In_482,In_78);
nor U1635 (N_1635,In_217,In_75);
and U1636 (N_1636,In_673,In_916);
or U1637 (N_1637,In_581,In_434);
nor U1638 (N_1638,In_202,In_691);
nand U1639 (N_1639,In_183,In_666);
xnor U1640 (N_1640,In_870,In_168);
xnor U1641 (N_1641,In_374,In_239);
and U1642 (N_1642,In_245,In_391);
and U1643 (N_1643,In_99,In_347);
nand U1644 (N_1644,In_680,In_409);
nor U1645 (N_1645,In_780,In_779);
xnor U1646 (N_1646,In_999,In_495);
nand U1647 (N_1647,In_176,In_344);
nor U1648 (N_1648,In_242,In_662);
and U1649 (N_1649,In_621,In_978);
or U1650 (N_1650,In_563,In_794);
and U1651 (N_1651,In_66,In_865);
nand U1652 (N_1652,In_117,In_648);
nor U1653 (N_1653,In_451,In_705);
nand U1654 (N_1654,In_710,In_668);
or U1655 (N_1655,In_62,In_750);
nand U1656 (N_1656,In_124,In_707);
or U1657 (N_1657,In_915,In_221);
nand U1658 (N_1658,In_394,In_953);
nor U1659 (N_1659,In_785,In_679);
nor U1660 (N_1660,In_975,In_885);
xnor U1661 (N_1661,In_681,In_281);
nand U1662 (N_1662,In_413,In_3);
or U1663 (N_1663,In_577,In_139);
or U1664 (N_1664,In_934,In_151);
nand U1665 (N_1665,In_242,In_429);
nor U1666 (N_1666,In_87,In_329);
xor U1667 (N_1667,In_640,In_130);
nand U1668 (N_1668,In_535,In_772);
nand U1669 (N_1669,In_499,In_325);
nor U1670 (N_1670,In_110,In_224);
and U1671 (N_1671,In_716,In_405);
and U1672 (N_1672,In_830,In_612);
and U1673 (N_1673,In_552,In_776);
nand U1674 (N_1674,In_759,In_101);
or U1675 (N_1675,In_474,In_623);
and U1676 (N_1676,In_312,In_482);
nand U1677 (N_1677,In_952,In_767);
or U1678 (N_1678,In_879,In_100);
or U1679 (N_1679,In_250,In_970);
nor U1680 (N_1680,In_917,In_141);
nand U1681 (N_1681,In_604,In_40);
nor U1682 (N_1682,In_889,In_12);
nand U1683 (N_1683,In_508,In_183);
nand U1684 (N_1684,In_388,In_445);
nor U1685 (N_1685,In_793,In_663);
nand U1686 (N_1686,In_429,In_195);
and U1687 (N_1687,In_758,In_442);
or U1688 (N_1688,In_515,In_504);
and U1689 (N_1689,In_173,In_402);
nand U1690 (N_1690,In_493,In_474);
and U1691 (N_1691,In_158,In_985);
or U1692 (N_1692,In_228,In_180);
and U1693 (N_1693,In_207,In_199);
and U1694 (N_1694,In_550,In_797);
nor U1695 (N_1695,In_184,In_784);
nor U1696 (N_1696,In_660,In_403);
nand U1697 (N_1697,In_629,In_327);
and U1698 (N_1698,In_17,In_324);
or U1699 (N_1699,In_774,In_202);
nor U1700 (N_1700,In_151,In_544);
and U1701 (N_1701,In_729,In_347);
nor U1702 (N_1702,In_579,In_478);
and U1703 (N_1703,In_363,In_948);
or U1704 (N_1704,In_532,In_237);
xor U1705 (N_1705,In_126,In_736);
nand U1706 (N_1706,In_497,In_286);
nand U1707 (N_1707,In_365,In_36);
and U1708 (N_1708,In_347,In_195);
and U1709 (N_1709,In_972,In_92);
nor U1710 (N_1710,In_142,In_271);
and U1711 (N_1711,In_959,In_503);
xor U1712 (N_1712,In_938,In_737);
or U1713 (N_1713,In_633,In_798);
or U1714 (N_1714,In_32,In_431);
or U1715 (N_1715,In_842,In_339);
or U1716 (N_1716,In_773,In_609);
nor U1717 (N_1717,In_237,In_816);
nor U1718 (N_1718,In_841,In_13);
nor U1719 (N_1719,In_892,In_538);
or U1720 (N_1720,In_769,In_952);
or U1721 (N_1721,In_408,In_735);
nor U1722 (N_1722,In_2,In_457);
or U1723 (N_1723,In_3,In_206);
nand U1724 (N_1724,In_937,In_495);
and U1725 (N_1725,In_813,In_78);
nor U1726 (N_1726,In_84,In_108);
nand U1727 (N_1727,In_386,In_192);
nand U1728 (N_1728,In_781,In_288);
or U1729 (N_1729,In_988,In_267);
xnor U1730 (N_1730,In_951,In_265);
xor U1731 (N_1731,In_812,In_889);
and U1732 (N_1732,In_940,In_618);
nand U1733 (N_1733,In_276,In_834);
or U1734 (N_1734,In_724,In_642);
or U1735 (N_1735,In_915,In_217);
nand U1736 (N_1736,In_805,In_42);
and U1737 (N_1737,In_48,In_955);
and U1738 (N_1738,In_136,In_70);
nand U1739 (N_1739,In_259,In_576);
and U1740 (N_1740,In_884,In_995);
or U1741 (N_1741,In_629,In_618);
and U1742 (N_1742,In_708,In_948);
or U1743 (N_1743,In_237,In_403);
and U1744 (N_1744,In_769,In_131);
nand U1745 (N_1745,In_734,In_80);
or U1746 (N_1746,In_351,In_69);
and U1747 (N_1747,In_499,In_956);
nand U1748 (N_1748,In_688,In_855);
nor U1749 (N_1749,In_395,In_909);
nand U1750 (N_1750,In_223,In_927);
nor U1751 (N_1751,In_332,In_215);
or U1752 (N_1752,In_341,In_951);
xor U1753 (N_1753,In_797,In_281);
and U1754 (N_1754,In_359,In_479);
or U1755 (N_1755,In_416,In_413);
nor U1756 (N_1756,In_18,In_379);
nand U1757 (N_1757,In_774,In_185);
or U1758 (N_1758,In_488,In_283);
nand U1759 (N_1759,In_317,In_958);
or U1760 (N_1760,In_386,In_590);
nand U1761 (N_1761,In_969,In_109);
nor U1762 (N_1762,In_378,In_0);
nor U1763 (N_1763,In_372,In_368);
nor U1764 (N_1764,In_764,In_955);
nand U1765 (N_1765,In_156,In_888);
or U1766 (N_1766,In_758,In_330);
nand U1767 (N_1767,In_677,In_221);
nor U1768 (N_1768,In_761,In_924);
and U1769 (N_1769,In_264,In_403);
or U1770 (N_1770,In_892,In_464);
nand U1771 (N_1771,In_828,In_346);
and U1772 (N_1772,In_543,In_185);
nand U1773 (N_1773,In_362,In_900);
or U1774 (N_1774,In_994,In_574);
nor U1775 (N_1775,In_58,In_958);
nand U1776 (N_1776,In_556,In_997);
and U1777 (N_1777,In_617,In_372);
nand U1778 (N_1778,In_860,In_6);
or U1779 (N_1779,In_113,In_598);
and U1780 (N_1780,In_243,In_749);
nand U1781 (N_1781,In_241,In_522);
nand U1782 (N_1782,In_34,In_470);
nand U1783 (N_1783,In_909,In_988);
or U1784 (N_1784,In_516,In_631);
and U1785 (N_1785,In_489,In_176);
nand U1786 (N_1786,In_650,In_965);
nand U1787 (N_1787,In_423,In_473);
xor U1788 (N_1788,In_666,In_82);
nand U1789 (N_1789,In_259,In_209);
or U1790 (N_1790,In_375,In_879);
and U1791 (N_1791,In_593,In_885);
nor U1792 (N_1792,In_493,In_626);
or U1793 (N_1793,In_396,In_917);
nor U1794 (N_1794,In_976,In_527);
nor U1795 (N_1795,In_630,In_470);
nand U1796 (N_1796,In_919,In_152);
and U1797 (N_1797,In_349,In_586);
nand U1798 (N_1798,In_855,In_143);
or U1799 (N_1799,In_546,In_628);
and U1800 (N_1800,In_581,In_400);
and U1801 (N_1801,In_719,In_304);
and U1802 (N_1802,In_106,In_648);
or U1803 (N_1803,In_46,In_689);
nand U1804 (N_1804,In_203,In_91);
nor U1805 (N_1805,In_378,In_472);
or U1806 (N_1806,In_902,In_472);
xor U1807 (N_1807,In_601,In_784);
and U1808 (N_1808,In_999,In_522);
or U1809 (N_1809,In_935,In_642);
and U1810 (N_1810,In_762,In_647);
and U1811 (N_1811,In_981,In_171);
nand U1812 (N_1812,In_131,In_126);
nor U1813 (N_1813,In_274,In_307);
nor U1814 (N_1814,In_547,In_995);
nand U1815 (N_1815,In_225,In_421);
nor U1816 (N_1816,In_620,In_322);
xnor U1817 (N_1817,In_344,In_948);
nor U1818 (N_1818,In_850,In_514);
nand U1819 (N_1819,In_517,In_9);
nor U1820 (N_1820,In_88,In_624);
and U1821 (N_1821,In_565,In_581);
and U1822 (N_1822,In_965,In_506);
xor U1823 (N_1823,In_71,In_149);
nand U1824 (N_1824,In_450,In_890);
or U1825 (N_1825,In_411,In_464);
and U1826 (N_1826,In_17,In_338);
xor U1827 (N_1827,In_174,In_137);
and U1828 (N_1828,In_702,In_402);
or U1829 (N_1829,In_632,In_334);
or U1830 (N_1830,In_732,In_497);
nor U1831 (N_1831,In_962,In_705);
and U1832 (N_1832,In_86,In_26);
nor U1833 (N_1833,In_591,In_635);
and U1834 (N_1834,In_792,In_843);
and U1835 (N_1835,In_429,In_962);
xor U1836 (N_1836,In_496,In_717);
nor U1837 (N_1837,In_879,In_209);
xnor U1838 (N_1838,In_776,In_532);
nand U1839 (N_1839,In_654,In_509);
nor U1840 (N_1840,In_188,In_544);
nand U1841 (N_1841,In_725,In_323);
nand U1842 (N_1842,In_523,In_96);
or U1843 (N_1843,In_741,In_238);
nand U1844 (N_1844,In_80,In_46);
or U1845 (N_1845,In_377,In_77);
and U1846 (N_1846,In_113,In_843);
or U1847 (N_1847,In_603,In_355);
nand U1848 (N_1848,In_763,In_4);
or U1849 (N_1849,In_300,In_375);
or U1850 (N_1850,In_497,In_80);
and U1851 (N_1851,In_949,In_441);
nor U1852 (N_1852,In_536,In_427);
or U1853 (N_1853,In_363,In_919);
nand U1854 (N_1854,In_342,In_990);
or U1855 (N_1855,In_378,In_168);
nor U1856 (N_1856,In_930,In_284);
and U1857 (N_1857,In_240,In_510);
or U1858 (N_1858,In_584,In_970);
and U1859 (N_1859,In_195,In_670);
nor U1860 (N_1860,In_249,In_400);
or U1861 (N_1861,In_883,In_46);
nand U1862 (N_1862,In_610,In_768);
nand U1863 (N_1863,In_522,In_389);
and U1864 (N_1864,In_593,In_49);
nor U1865 (N_1865,In_178,In_685);
or U1866 (N_1866,In_465,In_512);
nand U1867 (N_1867,In_41,In_10);
nor U1868 (N_1868,In_717,In_629);
nand U1869 (N_1869,In_625,In_85);
nor U1870 (N_1870,In_629,In_680);
xnor U1871 (N_1871,In_75,In_642);
and U1872 (N_1872,In_634,In_30);
xor U1873 (N_1873,In_249,In_768);
nor U1874 (N_1874,In_269,In_865);
or U1875 (N_1875,In_719,In_741);
nor U1876 (N_1876,In_162,In_701);
and U1877 (N_1877,In_97,In_739);
xnor U1878 (N_1878,In_83,In_252);
or U1879 (N_1879,In_891,In_654);
or U1880 (N_1880,In_55,In_489);
nor U1881 (N_1881,In_334,In_578);
or U1882 (N_1882,In_490,In_461);
and U1883 (N_1883,In_540,In_255);
and U1884 (N_1884,In_565,In_47);
or U1885 (N_1885,In_987,In_389);
nand U1886 (N_1886,In_610,In_709);
nand U1887 (N_1887,In_737,In_392);
nand U1888 (N_1888,In_776,In_484);
nor U1889 (N_1889,In_694,In_545);
or U1890 (N_1890,In_498,In_129);
xnor U1891 (N_1891,In_714,In_836);
nand U1892 (N_1892,In_588,In_631);
or U1893 (N_1893,In_176,In_241);
xor U1894 (N_1894,In_78,In_763);
nand U1895 (N_1895,In_296,In_706);
or U1896 (N_1896,In_934,In_247);
nor U1897 (N_1897,In_189,In_374);
nand U1898 (N_1898,In_430,In_453);
nor U1899 (N_1899,In_503,In_23);
and U1900 (N_1900,In_821,In_5);
nand U1901 (N_1901,In_283,In_722);
and U1902 (N_1902,In_864,In_655);
nor U1903 (N_1903,In_278,In_146);
and U1904 (N_1904,In_690,In_420);
xnor U1905 (N_1905,In_178,In_675);
nor U1906 (N_1906,In_510,In_769);
and U1907 (N_1907,In_144,In_449);
nor U1908 (N_1908,In_270,In_274);
or U1909 (N_1909,In_163,In_611);
xnor U1910 (N_1910,In_991,In_766);
and U1911 (N_1911,In_291,In_312);
nand U1912 (N_1912,In_574,In_552);
nor U1913 (N_1913,In_446,In_301);
nand U1914 (N_1914,In_161,In_212);
and U1915 (N_1915,In_775,In_116);
nand U1916 (N_1916,In_366,In_421);
or U1917 (N_1917,In_484,In_628);
and U1918 (N_1918,In_801,In_218);
or U1919 (N_1919,In_79,In_492);
or U1920 (N_1920,In_709,In_472);
or U1921 (N_1921,In_125,In_46);
and U1922 (N_1922,In_365,In_610);
and U1923 (N_1923,In_296,In_927);
and U1924 (N_1924,In_343,In_68);
nand U1925 (N_1925,In_241,In_715);
nand U1926 (N_1926,In_937,In_293);
and U1927 (N_1927,In_719,In_138);
nand U1928 (N_1928,In_614,In_738);
nand U1929 (N_1929,In_855,In_929);
xnor U1930 (N_1930,In_391,In_274);
nor U1931 (N_1931,In_370,In_783);
nor U1932 (N_1932,In_513,In_866);
or U1933 (N_1933,In_327,In_961);
nand U1934 (N_1934,In_889,In_463);
or U1935 (N_1935,In_248,In_192);
xnor U1936 (N_1936,In_480,In_328);
xor U1937 (N_1937,In_144,In_215);
nor U1938 (N_1938,In_82,In_539);
nand U1939 (N_1939,In_823,In_938);
nand U1940 (N_1940,In_340,In_189);
and U1941 (N_1941,In_553,In_783);
or U1942 (N_1942,In_814,In_236);
nor U1943 (N_1943,In_118,In_695);
nor U1944 (N_1944,In_559,In_472);
and U1945 (N_1945,In_693,In_344);
or U1946 (N_1946,In_439,In_549);
and U1947 (N_1947,In_508,In_960);
nand U1948 (N_1948,In_473,In_281);
and U1949 (N_1949,In_376,In_888);
xor U1950 (N_1950,In_380,In_329);
or U1951 (N_1951,In_236,In_675);
or U1952 (N_1952,In_131,In_543);
and U1953 (N_1953,In_946,In_792);
nand U1954 (N_1954,In_870,In_449);
nand U1955 (N_1955,In_128,In_702);
and U1956 (N_1956,In_84,In_605);
or U1957 (N_1957,In_574,In_956);
or U1958 (N_1958,In_10,In_68);
and U1959 (N_1959,In_954,In_340);
or U1960 (N_1960,In_355,In_423);
xor U1961 (N_1961,In_196,In_974);
nor U1962 (N_1962,In_315,In_496);
xnor U1963 (N_1963,In_62,In_931);
xor U1964 (N_1964,In_854,In_372);
or U1965 (N_1965,In_929,In_776);
or U1966 (N_1966,In_678,In_430);
or U1967 (N_1967,In_69,In_425);
nor U1968 (N_1968,In_765,In_56);
nand U1969 (N_1969,In_782,In_755);
and U1970 (N_1970,In_304,In_909);
or U1971 (N_1971,In_91,In_549);
and U1972 (N_1972,In_718,In_682);
nor U1973 (N_1973,In_999,In_118);
xnor U1974 (N_1974,In_173,In_659);
nor U1975 (N_1975,In_323,In_767);
or U1976 (N_1976,In_110,In_506);
or U1977 (N_1977,In_663,In_500);
nand U1978 (N_1978,In_234,In_415);
nor U1979 (N_1979,In_799,In_614);
or U1980 (N_1980,In_235,In_420);
nor U1981 (N_1981,In_932,In_697);
and U1982 (N_1982,In_290,In_113);
nand U1983 (N_1983,In_740,In_148);
or U1984 (N_1984,In_623,In_552);
and U1985 (N_1985,In_219,In_743);
nor U1986 (N_1986,In_268,In_464);
and U1987 (N_1987,In_417,In_575);
and U1988 (N_1988,In_36,In_164);
or U1989 (N_1989,In_498,In_800);
xnor U1990 (N_1990,In_407,In_240);
nand U1991 (N_1991,In_486,In_267);
nand U1992 (N_1992,In_855,In_783);
nor U1993 (N_1993,In_105,In_36);
nand U1994 (N_1994,In_149,In_669);
and U1995 (N_1995,In_343,In_903);
nand U1996 (N_1996,In_398,In_854);
or U1997 (N_1997,In_73,In_736);
and U1998 (N_1998,In_743,In_384);
and U1999 (N_1999,In_705,In_612);
and U2000 (N_2000,In_125,In_443);
xor U2001 (N_2001,In_13,In_141);
nand U2002 (N_2002,In_489,In_204);
or U2003 (N_2003,In_745,In_30);
and U2004 (N_2004,In_987,In_879);
nor U2005 (N_2005,In_707,In_54);
nand U2006 (N_2006,In_578,In_533);
or U2007 (N_2007,In_634,In_755);
or U2008 (N_2008,In_610,In_469);
or U2009 (N_2009,In_934,In_716);
nand U2010 (N_2010,In_13,In_720);
xnor U2011 (N_2011,In_121,In_462);
nand U2012 (N_2012,In_379,In_24);
nand U2013 (N_2013,In_298,In_757);
xor U2014 (N_2014,In_639,In_401);
nand U2015 (N_2015,In_141,In_21);
nand U2016 (N_2016,In_471,In_355);
nor U2017 (N_2017,In_788,In_89);
nand U2018 (N_2018,In_984,In_382);
and U2019 (N_2019,In_996,In_338);
or U2020 (N_2020,In_853,In_649);
or U2021 (N_2021,In_41,In_200);
nor U2022 (N_2022,In_564,In_837);
nand U2023 (N_2023,In_379,In_502);
nand U2024 (N_2024,In_610,In_464);
or U2025 (N_2025,In_706,In_888);
nand U2026 (N_2026,In_893,In_225);
and U2027 (N_2027,In_674,In_937);
nand U2028 (N_2028,In_329,In_360);
and U2029 (N_2029,In_189,In_647);
and U2030 (N_2030,In_200,In_838);
nand U2031 (N_2031,In_757,In_320);
nor U2032 (N_2032,In_573,In_732);
nor U2033 (N_2033,In_470,In_872);
nor U2034 (N_2034,In_264,In_333);
nor U2035 (N_2035,In_442,In_5);
or U2036 (N_2036,In_689,In_859);
nand U2037 (N_2037,In_976,In_780);
and U2038 (N_2038,In_562,In_726);
and U2039 (N_2039,In_73,In_500);
and U2040 (N_2040,In_769,In_175);
xnor U2041 (N_2041,In_170,In_26);
nor U2042 (N_2042,In_836,In_341);
or U2043 (N_2043,In_815,In_365);
nand U2044 (N_2044,In_313,In_955);
nor U2045 (N_2045,In_625,In_432);
or U2046 (N_2046,In_95,In_878);
nand U2047 (N_2047,In_408,In_828);
and U2048 (N_2048,In_798,In_800);
xnor U2049 (N_2049,In_453,In_644);
nand U2050 (N_2050,In_365,In_604);
nor U2051 (N_2051,In_691,In_433);
nand U2052 (N_2052,In_832,In_51);
and U2053 (N_2053,In_462,In_195);
nor U2054 (N_2054,In_401,In_931);
nor U2055 (N_2055,In_72,In_376);
nor U2056 (N_2056,In_373,In_346);
and U2057 (N_2057,In_190,In_696);
nor U2058 (N_2058,In_345,In_660);
nor U2059 (N_2059,In_526,In_675);
nand U2060 (N_2060,In_912,In_421);
or U2061 (N_2061,In_766,In_737);
xor U2062 (N_2062,In_13,In_618);
and U2063 (N_2063,In_656,In_985);
xnor U2064 (N_2064,In_797,In_952);
or U2065 (N_2065,In_380,In_292);
and U2066 (N_2066,In_792,In_342);
nor U2067 (N_2067,In_844,In_72);
nor U2068 (N_2068,In_937,In_516);
and U2069 (N_2069,In_672,In_812);
nor U2070 (N_2070,In_664,In_836);
nand U2071 (N_2071,In_297,In_682);
or U2072 (N_2072,In_145,In_418);
or U2073 (N_2073,In_352,In_550);
nor U2074 (N_2074,In_27,In_620);
and U2075 (N_2075,In_823,In_897);
nand U2076 (N_2076,In_327,In_167);
nor U2077 (N_2077,In_336,In_459);
xnor U2078 (N_2078,In_563,In_912);
and U2079 (N_2079,In_430,In_700);
nand U2080 (N_2080,In_94,In_474);
nor U2081 (N_2081,In_898,In_98);
nor U2082 (N_2082,In_541,In_906);
or U2083 (N_2083,In_532,In_710);
nor U2084 (N_2084,In_529,In_916);
nand U2085 (N_2085,In_935,In_491);
nor U2086 (N_2086,In_898,In_432);
and U2087 (N_2087,In_376,In_863);
nand U2088 (N_2088,In_123,In_68);
nand U2089 (N_2089,In_609,In_776);
and U2090 (N_2090,In_671,In_990);
or U2091 (N_2091,In_195,In_816);
nor U2092 (N_2092,In_641,In_799);
and U2093 (N_2093,In_514,In_782);
nand U2094 (N_2094,In_404,In_989);
nand U2095 (N_2095,In_44,In_378);
nor U2096 (N_2096,In_315,In_450);
or U2097 (N_2097,In_179,In_349);
and U2098 (N_2098,In_699,In_261);
nand U2099 (N_2099,In_123,In_401);
nand U2100 (N_2100,In_524,In_596);
nand U2101 (N_2101,In_147,In_168);
nand U2102 (N_2102,In_207,In_202);
or U2103 (N_2103,In_584,In_533);
nor U2104 (N_2104,In_117,In_859);
or U2105 (N_2105,In_929,In_689);
nor U2106 (N_2106,In_461,In_856);
and U2107 (N_2107,In_674,In_233);
nor U2108 (N_2108,In_930,In_754);
nor U2109 (N_2109,In_215,In_444);
nand U2110 (N_2110,In_433,In_366);
nor U2111 (N_2111,In_149,In_238);
and U2112 (N_2112,In_191,In_214);
or U2113 (N_2113,In_963,In_274);
nand U2114 (N_2114,In_508,In_203);
or U2115 (N_2115,In_187,In_803);
nor U2116 (N_2116,In_54,In_730);
nor U2117 (N_2117,In_545,In_733);
or U2118 (N_2118,In_305,In_315);
nand U2119 (N_2119,In_682,In_902);
xor U2120 (N_2120,In_879,In_477);
nand U2121 (N_2121,In_199,In_435);
nor U2122 (N_2122,In_280,In_751);
and U2123 (N_2123,In_595,In_819);
nor U2124 (N_2124,In_61,In_652);
nand U2125 (N_2125,In_310,In_240);
nand U2126 (N_2126,In_333,In_92);
and U2127 (N_2127,In_569,In_852);
nor U2128 (N_2128,In_373,In_685);
and U2129 (N_2129,In_938,In_33);
and U2130 (N_2130,In_239,In_831);
or U2131 (N_2131,In_66,In_846);
and U2132 (N_2132,In_872,In_180);
xor U2133 (N_2133,In_555,In_39);
nor U2134 (N_2134,In_483,In_701);
or U2135 (N_2135,In_547,In_631);
nand U2136 (N_2136,In_83,In_120);
nor U2137 (N_2137,In_704,In_616);
or U2138 (N_2138,In_651,In_522);
and U2139 (N_2139,In_736,In_61);
and U2140 (N_2140,In_917,In_572);
xor U2141 (N_2141,In_269,In_834);
or U2142 (N_2142,In_471,In_219);
and U2143 (N_2143,In_890,In_803);
nand U2144 (N_2144,In_849,In_540);
and U2145 (N_2145,In_46,In_138);
xor U2146 (N_2146,In_732,In_875);
nor U2147 (N_2147,In_98,In_964);
nor U2148 (N_2148,In_845,In_904);
nor U2149 (N_2149,In_392,In_283);
nor U2150 (N_2150,In_151,In_454);
nor U2151 (N_2151,In_252,In_601);
and U2152 (N_2152,In_459,In_540);
xnor U2153 (N_2153,In_150,In_356);
xor U2154 (N_2154,In_148,In_477);
nand U2155 (N_2155,In_162,In_505);
nor U2156 (N_2156,In_534,In_787);
nand U2157 (N_2157,In_965,In_366);
nor U2158 (N_2158,In_229,In_623);
or U2159 (N_2159,In_615,In_910);
and U2160 (N_2160,In_67,In_885);
nand U2161 (N_2161,In_330,In_457);
or U2162 (N_2162,In_151,In_440);
nor U2163 (N_2163,In_440,In_375);
xnor U2164 (N_2164,In_558,In_322);
xnor U2165 (N_2165,In_464,In_43);
or U2166 (N_2166,In_570,In_265);
or U2167 (N_2167,In_270,In_598);
or U2168 (N_2168,In_851,In_931);
xnor U2169 (N_2169,In_150,In_751);
or U2170 (N_2170,In_466,In_765);
and U2171 (N_2171,In_552,In_23);
or U2172 (N_2172,In_154,In_964);
nand U2173 (N_2173,In_944,In_249);
or U2174 (N_2174,In_578,In_545);
and U2175 (N_2175,In_590,In_594);
or U2176 (N_2176,In_833,In_384);
or U2177 (N_2177,In_584,In_714);
nor U2178 (N_2178,In_533,In_781);
nor U2179 (N_2179,In_550,In_818);
xnor U2180 (N_2180,In_368,In_246);
or U2181 (N_2181,In_818,In_928);
nand U2182 (N_2182,In_433,In_345);
xnor U2183 (N_2183,In_450,In_142);
nand U2184 (N_2184,In_534,In_779);
or U2185 (N_2185,In_855,In_330);
xnor U2186 (N_2186,In_719,In_517);
and U2187 (N_2187,In_40,In_651);
and U2188 (N_2188,In_969,In_465);
or U2189 (N_2189,In_647,In_259);
or U2190 (N_2190,In_458,In_141);
or U2191 (N_2191,In_77,In_54);
or U2192 (N_2192,In_73,In_632);
nor U2193 (N_2193,In_780,In_230);
and U2194 (N_2194,In_472,In_338);
or U2195 (N_2195,In_981,In_736);
nand U2196 (N_2196,In_548,In_700);
and U2197 (N_2197,In_59,In_804);
nand U2198 (N_2198,In_178,In_794);
and U2199 (N_2199,In_744,In_727);
or U2200 (N_2200,In_621,In_561);
and U2201 (N_2201,In_845,In_666);
xnor U2202 (N_2202,In_959,In_256);
nor U2203 (N_2203,In_221,In_42);
or U2204 (N_2204,In_186,In_528);
or U2205 (N_2205,In_561,In_447);
and U2206 (N_2206,In_472,In_780);
nand U2207 (N_2207,In_924,In_496);
nand U2208 (N_2208,In_777,In_609);
nand U2209 (N_2209,In_664,In_356);
or U2210 (N_2210,In_357,In_769);
xor U2211 (N_2211,In_445,In_142);
and U2212 (N_2212,In_285,In_835);
or U2213 (N_2213,In_508,In_250);
nand U2214 (N_2214,In_448,In_384);
nand U2215 (N_2215,In_404,In_621);
or U2216 (N_2216,In_789,In_520);
nand U2217 (N_2217,In_399,In_715);
nand U2218 (N_2218,In_157,In_500);
and U2219 (N_2219,In_223,In_702);
nor U2220 (N_2220,In_325,In_88);
or U2221 (N_2221,In_961,In_239);
nand U2222 (N_2222,In_545,In_660);
and U2223 (N_2223,In_230,In_373);
nor U2224 (N_2224,In_461,In_967);
nor U2225 (N_2225,In_412,In_762);
and U2226 (N_2226,In_424,In_147);
xnor U2227 (N_2227,In_661,In_612);
or U2228 (N_2228,In_94,In_25);
nor U2229 (N_2229,In_762,In_152);
and U2230 (N_2230,In_622,In_49);
xnor U2231 (N_2231,In_120,In_812);
nor U2232 (N_2232,In_406,In_472);
nor U2233 (N_2233,In_219,In_13);
nand U2234 (N_2234,In_402,In_622);
and U2235 (N_2235,In_300,In_239);
or U2236 (N_2236,In_156,In_237);
or U2237 (N_2237,In_620,In_460);
nand U2238 (N_2238,In_657,In_837);
nand U2239 (N_2239,In_306,In_896);
or U2240 (N_2240,In_235,In_426);
and U2241 (N_2241,In_636,In_483);
or U2242 (N_2242,In_607,In_705);
or U2243 (N_2243,In_903,In_773);
or U2244 (N_2244,In_37,In_482);
or U2245 (N_2245,In_962,In_177);
and U2246 (N_2246,In_123,In_876);
nand U2247 (N_2247,In_43,In_284);
nand U2248 (N_2248,In_921,In_977);
or U2249 (N_2249,In_166,In_716);
or U2250 (N_2250,In_589,In_358);
nand U2251 (N_2251,In_466,In_205);
nor U2252 (N_2252,In_242,In_215);
nand U2253 (N_2253,In_172,In_612);
nor U2254 (N_2254,In_780,In_500);
and U2255 (N_2255,In_809,In_523);
or U2256 (N_2256,In_490,In_339);
or U2257 (N_2257,In_138,In_349);
nor U2258 (N_2258,In_430,In_898);
nor U2259 (N_2259,In_784,In_997);
and U2260 (N_2260,In_186,In_32);
nor U2261 (N_2261,In_527,In_81);
nand U2262 (N_2262,In_253,In_26);
nand U2263 (N_2263,In_563,In_627);
nand U2264 (N_2264,In_41,In_878);
nor U2265 (N_2265,In_443,In_942);
nor U2266 (N_2266,In_449,In_299);
nor U2267 (N_2267,In_708,In_170);
nor U2268 (N_2268,In_956,In_436);
or U2269 (N_2269,In_903,In_670);
nand U2270 (N_2270,In_353,In_357);
xor U2271 (N_2271,In_153,In_135);
xor U2272 (N_2272,In_402,In_995);
nand U2273 (N_2273,In_428,In_811);
nand U2274 (N_2274,In_214,In_960);
xnor U2275 (N_2275,In_793,In_379);
and U2276 (N_2276,In_312,In_268);
nand U2277 (N_2277,In_300,In_81);
and U2278 (N_2278,In_330,In_230);
nor U2279 (N_2279,In_426,In_793);
nand U2280 (N_2280,In_187,In_634);
and U2281 (N_2281,In_6,In_12);
xor U2282 (N_2282,In_872,In_257);
or U2283 (N_2283,In_233,In_439);
xor U2284 (N_2284,In_469,In_707);
and U2285 (N_2285,In_42,In_278);
nand U2286 (N_2286,In_129,In_101);
nor U2287 (N_2287,In_977,In_197);
and U2288 (N_2288,In_195,In_76);
nor U2289 (N_2289,In_754,In_226);
xnor U2290 (N_2290,In_478,In_773);
xnor U2291 (N_2291,In_626,In_765);
or U2292 (N_2292,In_661,In_808);
nand U2293 (N_2293,In_535,In_647);
or U2294 (N_2294,In_383,In_530);
xnor U2295 (N_2295,In_894,In_232);
nor U2296 (N_2296,In_870,In_487);
xor U2297 (N_2297,In_369,In_442);
and U2298 (N_2298,In_9,In_323);
and U2299 (N_2299,In_266,In_853);
nand U2300 (N_2300,In_796,In_487);
nand U2301 (N_2301,In_436,In_842);
nand U2302 (N_2302,In_727,In_983);
or U2303 (N_2303,In_83,In_628);
nand U2304 (N_2304,In_106,In_690);
or U2305 (N_2305,In_551,In_861);
xnor U2306 (N_2306,In_478,In_294);
or U2307 (N_2307,In_95,In_500);
nor U2308 (N_2308,In_691,In_373);
nand U2309 (N_2309,In_655,In_678);
xnor U2310 (N_2310,In_502,In_52);
or U2311 (N_2311,In_774,In_431);
nand U2312 (N_2312,In_705,In_221);
and U2313 (N_2313,In_442,In_880);
nor U2314 (N_2314,In_97,In_723);
and U2315 (N_2315,In_207,In_33);
nor U2316 (N_2316,In_22,In_885);
and U2317 (N_2317,In_778,In_73);
xor U2318 (N_2318,In_293,In_495);
nor U2319 (N_2319,In_662,In_924);
and U2320 (N_2320,In_14,In_62);
nand U2321 (N_2321,In_731,In_726);
nand U2322 (N_2322,In_433,In_539);
nand U2323 (N_2323,In_830,In_312);
or U2324 (N_2324,In_52,In_116);
xor U2325 (N_2325,In_465,In_43);
nor U2326 (N_2326,In_317,In_101);
nand U2327 (N_2327,In_943,In_392);
nor U2328 (N_2328,In_731,In_737);
nor U2329 (N_2329,In_401,In_785);
xnor U2330 (N_2330,In_23,In_693);
nand U2331 (N_2331,In_557,In_171);
xnor U2332 (N_2332,In_324,In_858);
and U2333 (N_2333,In_156,In_188);
nor U2334 (N_2334,In_286,In_469);
nor U2335 (N_2335,In_803,In_184);
nor U2336 (N_2336,In_158,In_702);
and U2337 (N_2337,In_488,In_252);
or U2338 (N_2338,In_192,In_560);
and U2339 (N_2339,In_861,In_225);
or U2340 (N_2340,In_53,In_372);
nand U2341 (N_2341,In_119,In_659);
and U2342 (N_2342,In_210,In_126);
nor U2343 (N_2343,In_413,In_154);
nand U2344 (N_2344,In_110,In_405);
or U2345 (N_2345,In_163,In_84);
or U2346 (N_2346,In_370,In_930);
and U2347 (N_2347,In_135,In_870);
nor U2348 (N_2348,In_853,In_351);
and U2349 (N_2349,In_256,In_332);
nand U2350 (N_2350,In_423,In_285);
or U2351 (N_2351,In_211,In_525);
or U2352 (N_2352,In_959,In_59);
or U2353 (N_2353,In_627,In_598);
nand U2354 (N_2354,In_452,In_446);
nor U2355 (N_2355,In_526,In_986);
nand U2356 (N_2356,In_439,In_64);
or U2357 (N_2357,In_981,In_321);
and U2358 (N_2358,In_523,In_958);
or U2359 (N_2359,In_84,In_500);
xnor U2360 (N_2360,In_842,In_748);
and U2361 (N_2361,In_123,In_164);
xor U2362 (N_2362,In_680,In_725);
or U2363 (N_2363,In_498,In_598);
and U2364 (N_2364,In_717,In_177);
or U2365 (N_2365,In_482,In_969);
nand U2366 (N_2366,In_789,In_649);
and U2367 (N_2367,In_41,In_935);
xor U2368 (N_2368,In_60,In_629);
nor U2369 (N_2369,In_991,In_413);
nor U2370 (N_2370,In_12,In_505);
or U2371 (N_2371,In_633,In_483);
nand U2372 (N_2372,In_377,In_717);
xor U2373 (N_2373,In_173,In_516);
nor U2374 (N_2374,In_564,In_668);
or U2375 (N_2375,In_444,In_944);
or U2376 (N_2376,In_290,In_602);
or U2377 (N_2377,In_17,In_849);
nor U2378 (N_2378,In_304,In_20);
or U2379 (N_2379,In_807,In_323);
nand U2380 (N_2380,In_856,In_580);
and U2381 (N_2381,In_404,In_838);
xor U2382 (N_2382,In_32,In_798);
or U2383 (N_2383,In_480,In_707);
and U2384 (N_2384,In_986,In_326);
nand U2385 (N_2385,In_694,In_885);
or U2386 (N_2386,In_285,In_754);
nand U2387 (N_2387,In_771,In_470);
nand U2388 (N_2388,In_519,In_878);
nand U2389 (N_2389,In_821,In_135);
nor U2390 (N_2390,In_996,In_817);
nor U2391 (N_2391,In_793,In_276);
or U2392 (N_2392,In_202,In_911);
or U2393 (N_2393,In_783,In_351);
or U2394 (N_2394,In_854,In_842);
nor U2395 (N_2395,In_246,In_192);
nand U2396 (N_2396,In_368,In_233);
nor U2397 (N_2397,In_218,In_385);
and U2398 (N_2398,In_140,In_518);
nor U2399 (N_2399,In_768,In_223);
and U2400 (N_2400,In_972,In_508);
nand U2401 (N_2401,In_161,In_511);
or U2402 (N_2402,In_818,In_525);
and U2403 (N_2403,In_642,In_84);
and U2404 (N_2404,In_249,In_931);
nor U2405 (N_2405,In_192,In_195);
and U2406 (N_2406,In_799,In_154);
nand U2407 (N_2407,In_722,In_305);
and U2408 (N_2408,In_806,In_799);
and U2409 (N_2409,In_545,In_661);
xnor U2410 (N_2410,In_412,In_537);
or U2411 (N_2411,In_166,In_218);
or U2412 (N_2412,In_226,In_644);
nand U2413 (N_2413,In_416,In_483);
and U2414 (N_2414,In_137,In_614);
xnor U2415 (N_2415,In_712,In_493);
and U2416 (N_2416,In_275,In_26);
nand U2417 (N_2417,In_466,In_523);
and U2418 (N_2418,In_937,In_838);
nand U2419 (N_2419,In_868,In_224);
nor U2420 (N_2420,In_620,In_151);
nand U2421 (N_2421,In_111,In_18);
nor U2422 (N_2422,In_964,In_472);
and U2423 (N_2423,In_931,In_185);
or U2424 (N_2424,In_300,In_314);
xor U2425 (N_2425,In_954,In_783);
xor U2426 (N_2426,In_105,In_282);
or U2427 (N_2427,In_762,In_371);
or U2428 (N_2428,In_92,In_289);
nor U2429 (N_2429,In_157,In_943);
and U2430 (N_2430,In_11,In_265);
nand U2431 (N_2431,In_961,In_445);
nor U2432 (N_2432,In_900,In_238);
nor U2433 (N_2433,In_962,In_605);
and U2434 (N_2434,In_228,In_944);
nand U2435 (N_2435,In_162,In_620);
or U2436 (N_2436,In_366,In_179);
and U2437 (N_2437,In_611,In_953);
nor U2438 (N_2438,In_985,In_895);
and U2439 (N_2439,In_841,In_945);
nand U2440 (N_2440,In_941,In_714);
xnor U2441 (N_2441,In_727,In_204);
nor U2442 (N_2442,In_484,In_928);
and U2443 (N_2443,In_978,In_658);
or U2444 (N_2444,In_495,In_688);
nor U2445 (N_2445,In_911,In_204);
or U2446 (N_2446,In_988,In_313);
and U2447 (N_2447,In_627,In_25);
and U2448 (N_2448,In_950,In_532);
or U2449 (N_2449,In_855,In_895);
nor U2450 (N_2450,In_2,In_156);
and U2451 (N_2451,In_653,In_882);
and U2452 (N_2452,In_190,In_841);
or U2453 (N_2453,In_964,In_603);
nor U2454 (N_2454,In_156,In_179);
and U2455 (N_2455,In_126,In_597);
nor U2456 (N_2456,In_438,In_596);
and U2457 (N_2457,In_290,In_477);
and U2458 (N_2458,In_803,In_106);
nor U2459 (N_2459,In_873,In_187);
nand U2460 (N_2460,In_495,In_92);
or U2461 (N_2461,In_880,In_145);
nor U2462 (N_2462,In_471,In_945);
nand U2463 (N_2463,In_124,In_689);
xnor U2464 (N_2464,In_36,In_130);
or U2465 (N_2465,In_994,In_141);
nand U2466 (N_2466,In_576,In_325);
or U2467 (N_2467,In_942,In_981);
nor U2468 (N_2468,In_347,In_323);
and U2469 (N_2469,In_454,In_192);
or U2470 (N_2470,In_543,In_737);
or U2471 (N_2471,In_494,In_652);
nand U2472 (N_2472,In_62,In_251);
nor U2473 (N_2473,In_596,In_76);
nand U2474 (N_2474,In_669,In_529);
nand U2475 (N_2475,In_845,In_398);
or U2476 (N_2476,In_406,In_145);
nand U2477 (N_2477,In_553,In_101);
nand U2478 (N_2478,In_100,In_453);
xor U2479 (N_2479,In_246,In_962);
and U2480 (N_2480,In_798,In_392);
nor U2481 (N_2481,In_823,In_965);
or U2482 (N_2482,In_486,In_18);
and U2483 (N_2483,In_425,In_388);
xnor U2484 (N_2484,In_249,In_729);
nand U2485 (N_2485,In_473,In_198);
nand U2486 (N_2486,In_220,In_116);
nand U2487 (N_2487,In_999,In_143);
or U2488 (N_2488,In_263,In_193);
nor U2489 (N_2489,In_217,In_955);
nand U2490 (N_2490,In_760,In_114);
or U2491 (N_2491,In_356,In_444);
nand U2492 (N_2492,In_910,In_652);
nand U2493 (N_2493,In_217,In_861);
nand U2494 (N_2494,In_120,In_392);
xor U2495 (N_2495,In_90,In_420);
or U2496 (N_2496,In_923,In_748);
or U2497 (N_2497,In_10,In_414);
or U2498 (N_2498,In_883,In_840);
or U2499 (N_2499,In_536,In_69);
or U2500 (N_2500,In_73,In_109);
and U2501 (N_2501,In_256,In_253);
nor U2502 (N_2502,In_715,In_167);
xor U2503 (N_2503,In_986,In_717);
or U2504 (N_2504,In_876,In_137);
and U2505 (N_2505,In_367,In_281);
or U2506 (N_2506,In_383,In_843);
or U2507 (N_2507,In_922,In_492);
and U2508 (N_2508,In_547,In_430);
nand U2509 (N_2509,In_241,In_340);
or U2510 (N_2510,In_467,In_502);
and U2511 (N_2511,In_228,In_798);
nand U2512 (N_2512,In_939,In_137);
nand U2513 (N_2513,In_196,In_783);
nor U2514 (N_2514,In_135,In_889);
and U2515 (N_2515,In_888,In_278);
nand U2516 (N_2516,In_815,In_491);
and U2517 (N_2517,In_892,In_303);
xor U2518 (N_2518,In_557,In_273);
xor U2519 (N_2519,In_390,In_466);
nand U2520 (N_2520,In_175,In_211);
nor U2521 (N_2521,In_890,In_931);
xor U2522 (N_2522,In_860,In_187);
nor U2523 (N_2523,In_407,In_537);
nor U2524 (N_2524,In_716,In_659);
xor U2525 (N_2525,In_406,In_835);
and U2526 (N_2526,In_312,In_757);
or U2527 (N_2527,In_932,In_933);
nor U2528 (N_2528,In_23,In_416);
and U2529 (N_2529,In_269,In_534);
and U2530 (N_2530,In_937,In_758);
nand U2531 (N_2531,In_362,In_574);
nor U2532 (N_2532,In_312,In_452);
or U2533 (N_2533,In_298,In_401);
and U2534 (N_2534,In_574,In_104);
nor U2535 (N_2535,In_130,In_813);
and U2536 (N_2536,In_352,In_90);
nand U2537 (N_2537,In_384,In_441);
and U2538 (N_2538,In_282,In_716);
nor U2539 (N_2539,In_631,In_201);
nor U2540 (N_2540,In_412,In_182);
or U2541 (N_2541,In_946,In_701);
nor U2542 (N_2542,In_911,In_770);
nor U2543 (N_2543,In_447,In_333);
or U2544 (N_2544,In_835,In_775);
nand U2545 (N_2545,In_444,In_425);
and U2546 (N_2546,In_115,In_473);
or U2547 (N_2547,In_880,In_949);
xnor U2548 (N_2548,In_118,In_204);
or U2549 (N_2549,In_383,In_45);
or U2550 (N_2550,In_523,In_103);
and U2551 (N_2551,In_697,In_273);
nor U2552 (N_2552,In_497,In_176);
xor U2553 (N_2553,In_520,In_246);
nor U2554 (N_2554,In_291,In_831);
nor U2555 (N_2555,In_521,In_92);
nor U2556 (N_2556,In_9,In_411);
or U2557 (N_2557,In_706,In_997);
or U2558 (N_2558,In_620,In_3);
and U2559 (N_2559,In_138,In_492);
and U2560 (N_2560,In_96,In_616);
nor U2561 (N_2561,In_660,In_698);
or U2562 (N_2562,In_969,In_517);
and U2563 (N_2563,In_659,In_521);
and U2564 (N_2564,In_855,In_590);
and U2565 (N_2565,In_658,In_65);
nand U2566 (N_2566,In_684,In_564);
nand U2567 (N_2567,In_482,In_589);
and U2568 (N_2568,In_438,In_535);
xnor U2569 (N_2569,In_37,In_756);
or U2570 (N_2570,In_280,In_894);
nor U2571 (N_2571,In_374,In_629);
nor U2572 (N_2572,In_188,In_690);
or U2573 (N_2573,In_566,In_523);
and U2574 (N_2574,In_381,In_25);
or U2575 (N_2575,In_226,In_372);
or U2576 (N_2576,In_601,In_114);
or U2577 (N_2577,In_852,In_975);
nand U2578 (N_2578,In_199,In_528);
nand U2579 (N_2579,In_569,In_624);
nor U2580 (N_2580,In_75,In_807);
nor U2581 (N_2581,In_403,In_445);
or U2582 (N_2582,In_843,In_119);
nand U2583 (N_2583,In_937,In_699);
and U2584 (N_2584,In_0,In_98);
or U2585 (N_2585,In_491,In_400);
nand U2586 (N_2586,In_356,In_403);
nor U2587 (N_2587,In_390,In_237);
or U2588 (N_2588,In_46,In_660);
nand U2589 (N_2589,In_417,In_319);
nor U2590 (N_2590,In_413,In_825);
or U2591 (N_2591,In_114,In_497);
and U2592 (N_2592,In_465,In_75);
and U2593 (N_2593,In_868,In_91);
nand U2594 (N_2594,In_613,In_66);
and U2595 (N_2595,In_996,In_884);
and U2596 (N_2596,In_129,In_678);
or U2597 (N_2597,In_710,In_800);
or U2598 (N_2598,In_562,In_191);
xor U2599 (N_2599,In_833,In_817);
and U2600 (N_2600,In_774,In_990);
or U2601 (N_2601,In_669,In_690);
or U2602 (N_2602,In_227,In_529);
nand U2603 (N_2603,In_718,In_229);
nor U2604 (N_2604,In_555,In_758);
nand U2605 (N_2605,In_142,In_957);
and U2606 (N_2606,In_88,In_622);
and U2607 (N_2607,In_51,In_73);
nor U2608 (N_2608,In_887,In_977);
and U2609 (N_2609,In_256,In_124);
and U2610 (N_2610,In_948,In_85);
and U2611 (N_2611,In_832,In_330);
and U2612 (N_2612,In_397,In_370);
xor U2613 (N_2613,In_18,In_523);
nor U2614 (N_2614,In_522,In_448);
or U2615 (N_2615,In_633,In_613);
and U2616 (N_2616,In_456,In_71);
or U2617 (N_2617,In_647,In_594);
and U2618 (N_2618,In_55,In_490);
xnor U2619 (N_2619,In_238,In_855);
or U2620 (N_2620,In_387,In_758);
xnor U2621 (N_2621,In_304,In_352);
and U2622 (N_2622,In_743,In_340);
or U2623 (N_2623,In_13,In_398);
nor U2624 (N_2624,In_117,In_79);
and U2625 (N_2625,In_990,In_797);
or U2626 (N_2626,In_657,In_444);
and U2627 (N_2627,In_56,In_713);
nor U2628 (N_2628,In_655,In_716);
or U2629 (N_2629,In_687,In_587);
xor U2630 (N_2630,In_249,In_868);
nand U2631 (N_2631,In_437,In_831);
nand U2632 (N_2632,In_552,In_727);
or U2633 (N_2633,In_601,In_291);
nor U2634 (N_2634,In_291,In_5);
nand U2635 (N_2635,In_280,In_657);
and U2636 (N_2636,In_893,In_840);
nand U2637 (N_2637,In_428,In_774);
nor U2638 (N_2638,In_516,In_733);
nor U2639 (N_2639,In_99,In_527);
and U2640 (N_2640,In_124,In_207);
nor U2641 (N_2641,In_191,In_880);
or U2642 (N_2642,In_61,In_66);
or U2643 (N_2643,In_379,In_98);
nor U2644 (N_2644,In_436,In_474);
nor U2645 (N_2645,In_940,In_158);
xor U2646 (N_2646,In_847,In_200);
nor U2647 (N_2647,In_90,In_981);
nand U2648 (N_2648,In_627,In_148);
or U2649 (N_2649,In_301,In_131);
or U2650 (N_2650,In_797,In_976);
nor U2651 (N_2651,In_693,In_356);
xor U2652 (N_2652,In_229,In_34);
and U2653 (N_2653,In_630,In_718);
xor U2654 (N_2654,In_733,In_605);
or U2655 (N_2655,In_288,In_187);
nor U2656 (N_2656,In_401,In_267);
nor U2657 (N_2657,In_381,In_106);
and U2658 (N_2658,In_170,In_1);
and U2659 (N_2659,In_64,In_628);
or U2660 (N_2660,In_660,In_414);
nand U2661 (N_2661,In_595,In_818);
nor U2662 (N_2662,In_705,In_650);
and U2663 (N_2663,In_605,In_977);
or U2664 (N_2664,In_178,In_129);
nor U2665 (N_2665,In_148,In_176);
xnor U2666 (N_2666,In_165,In_424);
or U2667 (N_2667,In_580,In_338);
nor U2668 (N_2668,In_495,In_599);
nand U2669 (N_2669,In_220,In_57);
or U2670 (N_2670,In_357,In_479);
and U2671 (N_2671,In_308,In_393);
nor U2672 (N_2672,In_306,In_816);
xnor U2673 (N_2673,In_232,In_562);
nand U2674 (N_2674,In_71,In_522);
and U2675 (N_2675,In_12,In_793);
nor U2676 (N_2676,In_816,In_881);
xor U2677 (N_2677,In_370,In_921);
nand U2678 (N_2678,In_598,In_67);
or U2679 (N_2679,In_830,In_579);
or U2680 (N_2680,In_346,In_426);
and U2681 (N_2681,In_64,In_701);
nand U2682 (N_2682,In_506,In_888);
nor U2683 (N_2683,In_605,In_713);
nor U2684 (N_2684,In_782,In_135);
or U2685 (N_2685,In_596,In_669);
or U2686 (N_2686,In_92,In_806);
nand U2687 (N_2687,In_491,In_386);
and U2688 (N_2688,In_390,In_88);
and U2689 (N_2689,In_437,In_826);
or U2690 (N_2690,In_714,In_123);
and U2691 (N_2691,In_323,In_260);
xor U2692 (N_2692,In_306,In_503);
or U2693 (N_2693,In_541,In_106);
and U2694 (N_2694,In_896,In_158);
or U2695 (N_2695,In_148,In_656);
nor U2696 (N_2696,In_922,In_208);
and U2697 (N_2697,In_865,In_872);
and U2698 (N_2698,In_673,In_192);
and U2699 (N_2699,In_579,In_624);
nand U2700 (N_2700,In_550,In_653);
nor U2701 (N_2701,In_491,In_603);
or U2702 (N_2702,In_808,In_179);
and U2703 (N_2703,In_560,In_557);
and U2704 (N_2704,In_787,In_527);
and U2705 (N_2705,In_949,In_899);
xnor U2706 (N_2706,In_864,In_53);
nor U2707 (N_2707,In_73,In_658);
and U2708 (N_2708,In_225,In_9);
nor U2709 (N_2709,In_518,In_337);
and U2710 (N_2710,In_974,In_777);
nor U2711 (N_2711,In_403,In_368);
nand U2712 (N_2712,In_344,In_189);
and U2713 (N_2713,In_73,In_969);
or U2714 (N_2714,In_771,In_104);
nor U2715 (N_2715,In_251,In_583);
nand U2716 (N_2716,In_36,In_417);
or U2717 (N_2717,In_166,In_915);
or U2718 (N_2718,In_648,In_694);
nand U2719 (N_2719,In_853,In_603);
and U2720 (N_2720,In_620,In_377);
nor U2721 (N_2721,In_523,In_248);
xor U2722 (N_2722,In_360,In_848);
nor U2723 (N_2723,In_619,In_570);
nand U2724 (N_2724,In_388,In_467);
nand U2725 (N_2725,In_177,In_154);
and U2726 (N_2726,In_179,In_734);
nand U2727 (N_2727,In_686,In_661);
or U2728 (N_2728,In_969,In_94);
and U2729 (N_2729,In_490,In_857);
and U2730 (N_2730,In_593,In_755);
nand U2731 (N_2731,In_866,In_663);
nand U2732 (N_2732,In_419,In_717);
and U2733 (N_2733,In_587,In_916);
or U2734 (N_2734,In_756,In_950);
and U2735 (N_2735,In_265,In_302);
nor U2736 (N_2736,In_129,In_543);
nand U2737 (N_2737,In_526,In_32);
or U2738 (N_2738,In_379,In_394);
nand U2739 (N_2739,In_107,In_771);
nand U2740 (N_2740,In_990,In_539);
or U2741 (N_2741,In_497,In_366);
and U2742 (N_2742,In_153,In_500);
nand U2743 (N_2743,In_449,In_246);
or U2744 (N_2744,In_46,In_957);
xnor U2745 (N_2745,In_504,In_359);
or U2746 (N_2746,In_458,In_780);
xor U2747 (N_2747,In_798,In_350);
and U2748 (N_2748,In_680,In_29);
and U2749 (N_2749,In_234,In_642);
or U2750 (N_2750,In_196,In_864);
or U2751 (N_2751,In_718,In_867);
nand U2752 (N_2752,In_924,In_819);
nor U2753 (N_2753,In_314,In_977);
xor U2754 (N_2754,In_498,In_923);
and U2755 (N_2755,In_738,In_988);
xnor U2756 (N_2756,In_877,In_671);
nand U2757 (N_2757,In_153,In_582);
xnor U2758 (N_2758,In_423,In_336);
or U2759 (N_2759,In_853,In_884);
nor U2760 (N_2760,In_345,In_0);
or U2761 (N_2761,In_100,In_83);
and U2762 (N_2762,In_845,In_966);
or U2763 (N_2763,In_476,In_144);
and U2764 (N_2764,In_580,In_987);
nor U2765 (N_2765,In_830,In_41);
or U2766 (N_2766,In_577,In_682);
and U2767 (N_2767,In_360,In_690);
nor U2768 (N_2768,In_872,In_341);
nor U2769 (N_2769,In_885,In_283);
nand U2770 (N_2770,In_394,In_627);
nor U2771 (N_2771,In_978,In_680);
xor U2772 (N_2772,In_784,In_239);
xor U2773 (N_2773,In_51,In_846);
and U2774 (N_2774,In_566,In_412);
xor U2775 (N_2775,In_416,In_694);
nand U2776 (N_2776,In_458,In_196);
xnor U2777 (N_2777,In_876,In_105);
nand U2778 (N_2778,In_718,In_785);
and U2779 (N_2779,In_858,In_869);
and U2780 (N_2780,In_894,In_430);
nor U2781 (N_2781,In_179,In_173);
nor U2782 (N_2782,In_951,In_561);
and U2783 (N_2783,In_668,In_615);
or U2784 (N_2784,In_48,In_891);
or U2785 (N_2785,In_787,In_373);
nand U2786 (N_2786,In_777,In_784);
nor U2787 (N_2787,In_830,In_549);
nand U2788 (N_2788,In_513,In_579);
and U2789 (N_2789,In_887,In_607);
and U2790 (N_2790,In_155,In_415);
nor U2791 (N_2791,In_739,In_184);
or U2792 (N_2792,In_600,In_475);
or U2793 (N_2793,In_738,In_449);
xor U2794 (N_2794,In_555,In_531);
nand U2795 (N_2795,In_57,In_205);
and U2796 (N_2796,In_501,In_692);
and U2797 (N_2797,In_946,In_540);
xor U2798 (N_2798,In_735,In_907);
and U2799 (N_2799,In_900,In_141);
nor U2800 (N_2800,In_22,In_731);
and U2801 (N_2801,In_688,In_258);
nor U2802 (N_2802,In_170,In_224);
and U2803 (N_2803,In_840,In_473);
nor U2804 (N_2804,In_423,In_591);
nand U2805 (N_2805,In_49,In_998);
nor U2806 (N_2806,In_902,In_203);
nor U2807 (N_2807,In_287,In_378);
and U2808 (N_2808,In_971,In_652);
and U2809 (N_2809,In_425,In_740);
and U2810 (N_2810,In_724,In_467);
and U2811 (N_2811,In_645,In_909);
nand U2812 (N_2812,In_43,In_831);
and U2813 (N_2813,In_411,In_823);
nor U2814 (N_2814,In_835,In_540);
and U2815 (N_2815,In_451,In_108);
nor U2816 (N_2816,In_641,In_243);
xnor U2817 (N_2817,In_353,In_780);
nand U2818 (N_2818,In_763,In_166);
nand U2819 (N_2819,In_496,In_157);
nor U2820 (N_2820,In_315,In_250);
nor U2821 (N_2821,In_558,In_472);
nor U2822 (N_2822,In_61,In_587);
nand U2823 (N_2823,In_279,In_428);
nor U2824 (N_2824,In_142,In_194);
nor U2825 (N_2825,In_644,In_311);
nand U2826 (N_2826,In_940,In_655);
or U2827 (N_2827,In_121,In_295);
or U2828 (N_2828,In_879,In_182);
xor U2829 (N_2829,In_208,In_476);
xor U2830 (N_2830,In_86,In_123);
nor U2831 (N_2831,In_395,In_944);
nand U2832 (N_2832,In_96,In_675);
and U2833 (N_2833,In_539,In_79);
and U2834 (N_2834,In_691,In_892);
nand U2835 (N_2835,In_618,In_258);
and U2836 (N_2836,In_903,In_160);
nor U2837 (N_2837,In_544,In_565);
or U2838 (N_2838,In_233,In_418);
and U2839 (N_2839,In_442,In_636);
nor U2840 (N_2840,In_718,In_574);
or U2841 (N_2841,In_607,In_783);
nor U2842 (N_2842,In_545,In_532);
xnor U2843 (N_2843,In_265,In_904);
and U2844 (N_2844,In_467,In_130);
nor U2845 (N_2845,In_259,In_229);
xor U2846 (N_2846,In_237,In_187);
and U2847 (N_2847,In_220,In_314);
nor U2848 (N_2848,In_580,In_336);
nor U2849 (N_2849,In_404,In_665);
nand U2850 (N_2850,In_423,In_682);
nor U2851 (N_2851,In_564,In_718);
nand U2852 (N_2852,In_364,In_433);
nor U2853 (N_2853,In_319,In_156);
and U2854 (N_2854,In_43,In_924);
nor U2855 (N_2855,In_232,In_610);
nor U2856 (N_2856,In_697,In_696);
or U2857 (N_2857,In_916,In_359);
nand U2858 (N_2858,In_380,In_644);
nand U2859 (N_2859,In_70,In_956);
nor U2860 (N_2860,In_86,In_362);
xor U2861 (N_2861,In_356,In_55);
and U2862 (N_2862,In_498,In_551);
nand U2863 (N_2863,In_250,In_943);
and U2864 (N_2864,In_999,In_67);
or U2865 (N_2865,In_469,In_90);
nand U2866 (N_2866,In_702,In_406);
nor U2867 (N_2867,In_703,In_750);
and U2868 (N_2868,In_192,In_406);
nand U2869 (N_2869,In_385,In_280);
or U2870 (N_2870,In_172,In_163);
nand U2871 (N_2871,In_148,In_428);
nor U2872 (N_2872,In_807,In_506);
and U2873 (N_2873,In_160,In_85);
nand U2874 (N_2874,In_620,In_585);
nor U2875 (N_2875,In_585,In_623);
nor U2876 (N_2876,In_897,In_215);
or U2877 (N_2877,In_441,In_316);
nand U2878 (N_2878,In_112,In_680);
nand U2879 (N_2879,In_7,In_253);
nor U2880 (N_2880,In_283,In_212);
nor U2881 (N_2881,In_353,In_21);
nor U2882 (N_2882,In_207,In_880);
or U2883 (N_2883,In_391,In_614);
and U2884 (N_2884,In_532,In_232);
xnor U2885 (N_2885,In_262,In_29);
and U2886 (N_2886,In_223,In_870);
or U2887 (N_2887,In_140,In_780);
or U2888 (N_2888,In_362,In_344);
and U2889 (N_2889,In_846,In_281);
xor U2890 (N_2890,In_196,In_612);
and U2891 (N_2891,In_444,In_873);
or U2892 (N_2892,In_932,In_730);
nor U2893 (N_2893,In_407,In_461);
and U2894 (N_2894,In_718,In_159);
and U2895 (N_2895,In_697,In_155);
or U2896 (N_2896,In_641,In_70);
nand U2897 (N_2897,In_35,In_209);
xnor U2898 (N_2898,In_573,In_364);
nand U2899 (N_2899,In_972,In_658);
and U2900 (N_2900,In_480,In_662);
nor U2901 (N_2901,In_268,In_237);
or U2902 (N_2902,In_424,In_476);
nor U2903 (N_2903,In_198,In_654);
nand U2904 (N_2904,In_967,In_381);
and U2905 (N_2905,In_900,In_150);
xor U2906 (N_2906,In_43,In_437);
xor U2907 (N_2907,In_336,In_601);
or U2908 (N_2908,In_980,In_306);
nand U2909 (N_2909,In_315,In_197);
nand U2910 (N_2910,In_627,In_473);
nand U2911 (N_2911,In_352,In_909);
xor U2912 (N_2912,In_43,In_12);
nor U2913 (N_2913,In_867,In_246);
xnor U2914 (N_2914,In_584,In_445);
or U2915 (N_2915,In_764,In_507);
nand U2916 (N_2916,In_827,In_234);
nor U2917 (N_2917,In_634,In_981);
nor U2918 (N_2918,In_698,In_159);
nand U2919 (N_2919,In_308,In_710);
nor U2920 (N_2920,In_604,In_234);
nor U2921 (N_2921,In_62,In_937);
or U2922 (N_2922,In_774,In_991);
and U2923 (N_2923,In_942,In_386);
and U2924 (N_2924,In_223,In_17);
and U2925 (N_2925,In_278,In_61);
or U2926 (N_2926,In_608,In_364);
and U2927 (N_2927,In_669,In_844);
nand U2928 (N_2928,In_911,In_813);
and U2929 (N_2929,In_664,In_561);
xnor U2930 (N_2930,In_887,In_783);
nand U2931 (N_2931,In_619,In_87);
nor U2932 (N_2932,In_821,In_201);
nand U2933 (N_2933,In_167,In_757);
nand U2934 (N_2934,In_624,In_751);
nor U2935 (N_2935,In_58,In_693);
and U2936 (N_2936,In_585,In_728);
nand U2937 (N_2937,In_841,In_554);
nand U2938 (N_2938,In_444,In_936);
or U2939 (N_2939,In_531,In_534);
nor U2940 (N_2940,In_883,In_798);
nor U2941 (N_2941,In_801,In_392);
nand U2942 (N_2942,In_545,In_284);
and U2943 (N_2943,In_710,In_527);
xor U2944 (N_2944,In_518,In_585);
xnor U2945 (N_2945,In_583,In_856);
nor U2946 (N_2946,In_34,In_860);
nor U2947 (N_2947,In_327,In_861);
nand U2948 (N_2948,In_688,In_92);
or U2949 (N_2949,In_30,In_819);
xor U2950 (N_2950,In_337,In_762);
nand U2951 (N_2951,In_753,In_0);
xor U2952 (N_2952,In_542,In_617);
nor U2953 (N_2953,In_883,In_570);
nor U2954 (N_2954,In_529,In_711);
nand U2955 (N_2955,In_193,In_615);
or U2956 (N_2956,In_858,In_120);
and U2957 (N_2957,In_775,In_522);
and U2958 (N_2958,In_750,In_924);
or U2959 (N_2959,In_65,In_113);
xor U2960 (N_2960,In_689,In_337);
or U2961 (N_2961,In_892,In_818);
or U2962 (N_2962,In_495,In_38);
nor U2963 (N_2963,In_299,In_173);
nand U2964 (N_2964,In_713,In_441);
or U2965 (N_2965,In_141,In_78);
nand U2966 (N_2966,In_453,In_551);
nand U2967 (N_2967,In_833,In_772);
or U2968 (N_2968,In_48,In_407);
or U2969 (N_2969,In_229,In_305);
or U2970 (N_2970,In_969,In_525);
nor U2971 (N_2971,In_5,In_366);
or U2972 (N_2972,In_633,In_609);
nand U2973 (N_2973,In_682,In_882);
nor U2974 (N_2974,In_783,In_415);
nor U2975 (N_2975,In_603,In_480);
nand U2976 (N_2976,In_369,In_970);
and U2977 (N_2977,In_785,In_127);
xnor U2978 (N_2978,In_389,In_2);
nand U2979 (N_2979,In_452,In_740);
nor U2980 (N_2980,In_894,In_631);
nand U2981 (N_2981,In_26,In_203);
nand U2982 (N_2982,In_264,In_276);
or U2983 (N_2983,In_904,In_190);
or U2984 (N_2984,In_133,In_235);
and U2985 (N_2985,In_498,In_423);
nand U2986 (N_2986,In_625,In_179);
nor U2987 (N_2987,In_781,In_236);
xnor U2988 (N_2988,In_338,In_905);
nor U2989 (N_2989,In_729,In_553);
nor U2990 (N_2990,In_180,In_736);
or U2991 (N_2991,In_577,In_446);
nand U2992 (N_2992,In_764,In_793);
and U2993 (N_2993,In_200,In_146);
nor U2994 (N_2994,In_346,In_313);
or U2995 (N_2995,In_455,In_214);
and U2996 (N_2996,In_124,In_620);
nand U2997 (N_2997,In_865,In_986);
or U2998 (N_2998,In_608,In_209);
nor U2999 (N_2999,In_669,In_316);
nor U3000 (N_3000,In_628,In_386);
and U3001 (N_3001,In_921,In_854);
nor U3002 (N_3002,In_10,In_141);
and U3003 (N_3003,In_340,In_61);
nor U3004 (N_3004,In_264,In_703);
nor U3005 (N_3005,In_371,In_365);
or U3006 (N_3006,In_488,In_625);
nor U3007 (N_3007,In_957,In_841);
or U3008 (N_3008,In_812,In_41);
nand U3009 (N_3009,In_374,In_940);
or U3010 (N_3010,In_483,In_813);
nand U3011 (N_3011,In_830,In_987);
and U3012 (N_3012,In_436,In_3);
or U3013 (N_3013,In_56,In_652);
nor U3014 (N_3014,In_827,In_392);
xnor U3015 (N_3015,In_869,In_394);
or U3016 (N_3016,In_561,In_807);
nand U3017 (N_3017,In_555,In_151);
or U3018 (N_3018,In_146,In_160);
or U3019 (N_3019,In_936,In_358);
nand U3020 (N_3020,In_412,In_551);
and U3021 (N_3021,In_651,In_415);
or U3022 (N_3022,In_825,In_23);
nand U3023 (N_3023,In_787,In_100);
or U3024 (N_3024,In_599,In_335);
nand U3025 (N_3025,In_171,In_722);
and U3026 (N_3026,In_99,In_878);
or U3027 (N_3027,In_134,In_607);
and U3028 (N_3028,In_922,In_103);
nand U3029 (N_3029,In_183,In_468);
nor U3030 (N_3030,In_535,In_185);
and U3031 (N_3031,In_590,In_182);
and U3032 (N_3032,In_455,In_13);
nor U3033 (N_3033,In_956,In_14);
or U3034 (N_3034,In_599,In_922);
nand U3035 (N_3035,In_11,In_535);
and U3036 (N_3036,In_679,In_242);
or U3037 (N_3037,In_965,In_289);
nor U3038 (N_3038,In_897,In_361);
nand U3039 (N_3039,In_742,In_337);
and U3040 (N_3040,In_884,In_596);
nor U3041 (N_3041,In_361,In_844);
nand U3042 (N_3042,In_809,In_222);
and U3043 (N_3043,In_522,In_703);
nand U3044 (N_3044,In_413,In_689);
and U3045 (N_3045,In_420,In_650);
or U3046 (N_3046,In_544,In_846);
nor U3047 (N_3047,In_886,In_358);
nor U3048 (N_3048,In_365,In_817);
or U3049 (N_3049,In_41,In_615);
xnor U3050 (N_3050,In_176,In_164);
or U3051 (N_3051,In_185,In_228);
nand U3052 (N_3052,In_439,In_538);
and U3053 (N_3053,In_83,In_828);
nor U3054 (N_3054,In_841,In_448);
nand U3055 (N_3055,In_125,In_508);
nor U3056 (N_3056,In_346,In_97);
and U3057 (N_3057,In_215,In_646);
and U3058 (N_3058,In_269,In_507);
or U3059 (N_3059,In_862,In_495);
and U3060 (N_3060,In_341,In_774);
or U3061 (N_3061,In_479,In_757);
nand U3062 (N_3062,In_460,In_219);
and U3063 (N_3063,In_799,In_72);
nand U3064 (N_3064,In_475,In_921);
or U3065 (N_3065,In_637,In_886);
nand U3066 (N_3066,In_91,In_245);
nor U3067 (N_3067,In_681,In_79);
and U3068 (N_3068,In_572,In_250);
nand U3069 (N_3069,In_565,In_393);
and U3070 (N_3070,In_853,In_122);
nor U3071 (N_3071,In_586,In_579);
nand U3072 (N_3072,In_948,In_81);
or U3073 (N_3073,In_408,In_604);
or U3074 (N_3074,In_54,In_560);
xor U3075 (N_3075,In_816,In_287);
nor U3076 (N_3076,In_595,In_826);
or U3077 (N_3077,In_68,In_663);
nand U3078 (N_3078,In_903,In_626);
nor U3079 (N_3079,In_777,In_684);
nor U3080 (N_3080,In_156,In_800);
nor U3081 (N_3081,In_115,In_384);
nor U3082 (N_3082,In_978,In_96);
nand U3083 (N_3083,In_585,In_425);
nand U3084 (N_3084,In_432,In_436);
nor U3085 (N_3085,In_609,In_115);
or U3086 (N_3086,In_828,In_286);
nor U3087 (N_3087,In_352,In_347);
nor U3088 (N_3088,In_459,In_351);
and U3089 (N_3089,In_794,In_882);
xnor U3090 (N_3090,In_791,In_122);
or U3091 (N_3091,In_716,In_470);
or U3092 (N_3092,In_446,In_905);
xor U3093 (N_3093,In_582,In_143);
nand U3094 (N_3094,In_745,In_885);
or U3095 (N_3095,In_55,In_975);
and U3096 (N_3096,In_513,In_90);
and U3097 (N_3097,In_490,In_216);
nor U3098 (N_3098,In_936,In_673);
nand U3099 (N_3099,In_962,In_914);
and U3100 (N_3100,In_490,In_847);
and U3101 (N_3101,In_445,In_368);
xor U3102 (N_3102,In_557,In_239);
and U3103 (N_3103,In_563,In_894);
and U3104 (N_3104,In_206,In_942);
and U3105 (N_3105,In_20,In_59);
and U3106 (N_3106,In_181,In_918);
or U3107 (N_3107,In_904,In_44);
nand U3108 (N_3108,In_254,In_950);
or U3109 (N_3109,In_841,In_7);
or U3110 (N_3110,In_922,In_785);
or U3111 (N_3111,In_272,In_379);
or U3112 (N_3112,In_454,In_890);
xor U3113 (N_3113,In_959,In_757);
xor U3114 (N_3114,In_15,In_694);
xor U3115 (N_3115,In_110,In_754);
nand U3116 (N_3116,In_633,In_22);
and U3117 (N_3117,In_733,In_227);
nor U3118 (N_3118,In_591,In_688);
nand U3119 (N_3119,In_325,In_566);
or U3120 (N_3120,In_428,In_879);
nand U3121 (N_3121,In_261,In_283);
or U3122 (N_3122,In_545,In_102);
or U3123 (N_3123,In_891,In_750);
and U3124 (N_3124,In_78,In_797);
nand U3125 (N_3125,In_87,In_678);
and U3126 (N_3126,In_102,In_383);
xnor U3127 (N_3127,In_823,In_980);
nand U3128 (N_3128,In_294,In_399);
and U3129 (N_3129,In_358,In_547);
or U3130 (N_3130,In_193,In_61);
or U3131 (N_3131,In_923,In_547);
and U3132 (N_3132,In_408,In_486);
nand U3133 (N_3133,In_754,In_26);
nor U3134 (N_3134,In_710,In_9);
nand U3135 (N_3135,In_201,In_246);
nand U3136 (N_3136,In_295,In_930);
nor U3137 (N_3137,In_216,In_871);
or U3138 (N_3138,In_385,In_343);
nor U3139 (N_3139,In_674,In_902);
or U3140 (N_3140,In_13,In_512);
xnor U3141 (N_3141,In_206,In_851);
nand U3142 (N_3142,In_322,In_447);
nand U3143 (N_3143,In_748,In_32);
or U3144 (N_3144,In_663,In_353);
nor U3145 (N_3145,In_825,In_425);
nand U3146 (N_3146,In_875,In_216);
nand U3147 (N_3147,In_764,In_189);
or U3148 (N_3148,In_851,In_962);
nor U3149 (N_3149,In_209,In_601);
and U3150 (N_3150,In_488,In_903);
or U3151 (N_3151,In_16,In_61);
and U3152 (N_3152,In_865,In_283);
nand U3153 (N_3153,In_837,In_832);
and U3154 (N_3154,In_100,In_820);
xor U3155 (N_3155,In_934,In_268);
nor U3156 (N_3156,In_669,In_260);
or U3157 (N_3157,In_358,In_703);
nand U3158 (N_3158,In_304,In_211);
xor U3159 (N_3159,In_122,In_538);
or U3160 (N_3160,In_227,In_209);
and U3161 (N_3161,In_476,In_98);
or U3162 (N_3162,In_363,In_285);
or U3163 (N_3163,In_935,In_889);
xor U3164 (N_3164,In_414,In_871);
and U3165 (N_3165,In_752,In_397);
and U3166 (N_3166,In_181,In_616);
and U3167 (N_3167,In_717,In_40);
nor U3168 (N_3168,In_310,In_988);
xnor U3169 (N_3169,In_442,In_694);
nand U3170 (N_3170,In_26,In_103);
nor U3171 (N_3171,In_979,In_789);
xor U3172 (N_3172,In_343,In_187);
or U3173 (N_3173,In_734,In_856);
nor U3174 (N_3174,In_169,In_46);
nor U3175 (N_3175,In_373,In_374);
nand U3176 (N_3176,In_259,In_585);
or U3177 (N_3177,In_436,In_818);
or U3178 (N_3178,In_856,In_62);
nand U3179 (N_3179,In_849,In_155);
nand U3180 (N_3180,In_304,In_846);
nand U3181 (N_3181,In_287,In_687);
and U3182 (N_3182,In_692,In_7);
nor U3183 (N_3183,In_683,In_648);
and U3184 (N_3184,In_124,In_629);
nand U3185 (N_3185,In_554,In_179);
nor U3186 (N_3186,In_495,In_336);
or U3187 (N_3187,In_882,In_875);
or U3188 (N_3188,In_775,In_523);
and U3189 (N_3189,In_172,In_160);
nand U3190 (N_3190,In_213,In_488);
and U3191 (N_3191,In_253,In_796);
nor U3192 (N_3192,In_400,In_253);
and U3193 (N_3193,In_132,In_430);
or U3194 (N_3194,In_421,In_694);
nand U3195 (N_3195,In_176,In_483);
nand U3196 (N_3196,In_787,In_321);
and U3197 (N_3197,In_312,In_154);
nand U3198 (N_3198,In_506,In_666);
and U3199 (N_3199,In_984,In_469);
xor U3200 (N_3200,In_133,In_420);
nor U3201 (N_3201,In_645,In_638);
and U3202 (N_3202,In_221,In_615);
xor U3203 (N_3203,In_353,In_222);
or U3204 (N_3204,In_866,In_652);
and U3205 (N_3205,In_132,In_845);
nor U3206 (N_3206,In_982,In_512);
or U3207 (N_3207,In_785,In_215);
and U3208 (N_3208,In_480,In_393);
nand U3209 (N_3209,In_450,In_91);
and U3210 (N_3210,In_613,In_621);
or U3211 (N_3211,In_951,In_99);
nand U3212 (N_3212,In_352,In_773);
nand U3213 (N_3213,In_743,In_980);
and U3214 (N_3214,In_332,In_375);
nand U3215 (N_3215,In_482,In_923);
and U3216 (N_3216,In_230,In_861);
and U3217 (N_3217,In_807,In_600);
nor U3218 (N_3218,In_457,In_427);
nand U3219 (N_3219,In_924,In_122);
nor U3220 (N_3220,In_443,In_316);
nor U3221 (N_3221,In_454,In_897);
xor U3222 (N_3222,In_236,In_230);
or U3223 (N_3223,In_862,In_719);
nand U3224 (N_3224,In_725,In_703);
or U3225 (N_3225,In_228,In_215);
or U3226 (N_3226,In_424,In_75);
or U3227 (N_3227,In_405,In_513);
xor U3228 (N_3228,In_536,In_333);
and U3229 (N_3229,In_407,In_59);
nor U3230 (N_3230,In_193,In_594);
nand U3231 (N_3231,In_759,In_160);
nor U3232 (N_3232,In_290,In_216);
nand U3233 (N_3233,In_546,In_533);
nand U3234 (N_3234,In_685,In_411);
or U3235 (N_3235,In_33,In_626);
nor U3236 (N_3236,In_184,In_196);
nor U3237 (N_3237,In_593,In_435);
or U3238 (N_3238,In_770,In_341);
or U3239 (N_3239,In_826,In_684);
or U3240 (N_3240,In_494,In_798);
and U3241 (N_3241,In_409,In_108);
nor U3242 (N_3242,In_264,In_518);
or U3243 (N_3243,In_687,In_292);
or U3244 (N_3244,In_586,In_36);
nor U3245 (N_3245,In_431,In_44);
or U3246 (N_3246,In_539,In_544);
nand U3247 (N_3247,In_247,In_154);
nor U3248 (N_3248,In_350,In_748);
or U3249 (N_3249,In_672,In_457);
nand U3250 (N_3250,In_253,In_992);
nor U3251 (N_3251,In_473,In_221);
or U3252 (N_3252,In_956,In_107);
nand U3253 (N_3253,In_854,In_58);
and U3254 (N_3254,In_612,In_113);
or U3255 (N_3255,In_718,In_758);
nand U3256 (N_3256,In_464,In_605);
or U3257 (N_3257,In_349,In_628);
and U3258 (N_3258,In_720,In_625);
nor U3259 (N_3259,In_625,In_612);
nand U3260 (N_3260,In_335,In_807);
or U3261 (N_3261,In_511,In_267);
and U3262 (N_3262,In_950,In_37);
xnor U3263 (N_3263,In_37,In_541);
or U3264 (N_3264,In_96,In_384);
nor U3265 (N_3265,In_566,In_8);
and U3266 (N_3266,In_99,In_608);
xnor U3267 (N_3267,In_760,In_677);
nor U3268 (N_3268,In_95,In_339);
or U3269 (N_3269,In_959,In_958);
nand U3270 (N_3270,In_229,In_457);
xnor U3271 (N_3271,In_459,In_764);
or U3272 (N_3272,In_320,In_737);
nand U3273 (N_3273,In_539,In_953);
nand U3274 (N_3274,In_541,In_540);
and U3275 (N_3275,In_880,In_466);
and U3276 (N_3276,In_987,In_39);
nand U3277 (N_3277,In_106,In_481);
or U3278 (N_3278,In_5,In_681);
and U3279 (N_3279,In_829,In_407);
nor U3280 (N_3280,In_658,In_687);
or U3281 (N_3281,In_219,In_362);
nor U3282 (N_3282,In_166,In_922);
and U3283 (N_3283,In_415,In_191);
nand U3284 (N_3284,In_250,In_669);
nand U3285 (N_3285,In_374,In_155);
nand U3286 (N_3286,In_238,In_802);
or U3287 (N_3287,In_568,In_852);
and U3288 (N_3288,In_572,In_181);
xnor U3289 (N_3289,In_672,In_700);
nand U3290 (N_3290,In_565,In_291);
nand U3291 (N_3291,In_825,In_664);
or U3292 (N_3292,In_870,In_888);
or U3293 (N_3293,In_791,In_37);
nor U3294 (N_3294,In_776,In_475);
and U3295 (N_3295,In_887,In_105);
nor U3296 (N_3296,In_722,In_955);
nor U3297 (N_3297,In_405,In_805);
nor U3298 (N_3298,In_616,In_258);
xnor U3299 (N_3299,In_533,In_437);
nor U3300 (N_3300,In_790,In_703);
and U3301 (N_3301,In_930,In_949);
nand U3302 (N_3302,In_398,In_922);
or U3303 (N_3303,In_107,In_505);
nor U3304 (N_3304,In_575,In_269);
nand U3305 (N_3305,In_314,In_409);
nand U3306 (N_3306,In_299,In_339);
and U3307 (N_3307,In_192,In_726);
nor U3308 (N_3308,In_980,In_923);
or U3309 (N_3309,In_985,In_836);
nor U3310 (N_3310,In_377,In_945);
nor U3311 (N_3311,In_629,In_934);
xnor U3312 (N_3312,In_949,In_686);
nand U3313 (N_3313,In_64,In_862);
nor U3314 (N_3314,In_960,In_962);
xor U3315 (N_3315,In_907,In_712);
and U3316 (N_3316,In_474,In_930);
xor U3317 (N_3317,In_360,In_552);
and U3318 (N_3318,In_483,In_310);
or U3319 (N_3319,In_985,In_826);
or U3320 (N_3320,In_708,In_240);
nand U3321 (N_3321,In_299,In_682);
xor U3322 (N_3322,In_849,In_623);
and U3323 (N_3323,In_613,In_598);
and U3324 (N_3324,In_90,In_444);
or U3325 (N_3325,In_570,In_262);
or U3326 (N_3326,In_858,In_427);
nor U3327 (N_3327,In_608,In_468);
xor U3328 (N_3328,In_422,In_497);
and U3329 (N_3329,In_520,In_367);
nand U3330 (N_3330,In_14,In_157);
nand U3331 (N_3331,In_993,In_794);
or U3332 (N_3332,In_500,In_790);
nor U3333 (N_3333,In_427,In_480);
and U3334 (N_3334,In_543,In_966);
or U3335 (N_3335,In_26,In_402);
or U3336 (N_3336,In_614,In_729);
nand U3337 (N_3337,In_168,In_358);
nand U3338 (N_3338,In_708,In_174);
nor U3339 (N_3339,In_265,In_846);
or U3340 (N_3340,In_624,In_683);
and U3341 (N_3341,In_280,In_639);
nor U3342 (N_3342,In_28,In_320);
nand U3343 (N_3343,In_172,In_636);
nor U3344 (N_3344,In_844,In_547);
nand U3345 (N_3345,In_516,In_310);
nor U3346 (N_3346,In_738,In_326);
nor U3347 (N_3347,In_268,In_39);
nand U3348 (N_3348,In_339,In_685);
or U3349 (N_3349,In_96,In_768);
and U3350 (N_3350,In_497,In_770);
or U3351 (N_3351,In_128,In_920);
or U3352 (N_3352,In_690,In_646);
nand U3353 (N_3353,In_668,In_765);
or U3354 (N_3354,In_603,In_654);
nand U3355 (N_3355,In_237,In_964);
nor U3356 (N_3356,In_999,In_729);
nor U3357 (N_3357,In_41,In_785);
or U3358 (N_3358,In_515,In_170);
nand U3359 (N_3359,In_592,In_339);
nor U3360 (N_3360,In_514,In_328);
nand U3361 (N_3361,In_554,In_901);
or U3362 (N_3362,In_100,In_736);
xnor U3363 (N_3363,In_296,In_618);
nor U3364 (N_3364,In_108,In_633);
and U3365 (N_3365,In_522,In_605);
nor U3366 (N_3366,In_79,In_166);
nor U3367 (N_3367,In_670,In_458);
nor U3368 (N_3368,In_730,In_818);
and U3369 (N_3369,In_479,In_633);
and U3370 (N_3370,In_223,In_165);
nor U3371 (N_3371,In_102,In_462);
nor U3372 (N_3372,In_306,In_959);
nand U3373 (N_3373,In_891,In_304);
or U3374 (N_3374,In_383,In_538);
or U3375 (N_3375,In_197,In_522);
or U3376 (N_3376,In_931,In_783);
nor U3377 (N_3377,In_455,In_721);
or U3378 (N_3378,In_504,In_916);
or U3379 (N_3379,In_962,In_631);
or U3380 (N_3380,In_60,In_196);
xnor U3381 (N_3381,In_295,In_171);
and U3382 (N_3382,In_576,In_212);
or U3383 (N_3383,In_685,In_815);
and U3384 (N_3384,In_874,In_201);
and U3385 (N_3385,In_252,In_509);
or U3386 (N_3386,In_403,In_609);
xor U3387 (N_3387,In_687,In_379);
or U3388 (N_3388,In_42,In_673);
and U3389 (N_3389,In_515,In_114);
or U3390 (N_3390,In_951,In_60);
or U3391 (N_3391,In_513,In_379);
or U3392 (N_3392,In_955,In_109);
and U3393 (N_3393,In_100,In_592);
nor U3394 (N_3394,In_612,In_305);
or U3395 (N_3395,In_598,In_2);
or U3396 (N_3396,In_557,In_164);
and U3397 (N_3397,In_199,In_681);
nand U3398 (N_3398,In_801,In_811);
and U3399 (N_3399,In_382,In_515);
or U3400 (N_3400,In_257,In_301);
nand U3401 (N_3401,In_391,In_695);
xor U3402 (N_3402,In_127,In_619);
nand U3403 (N_3403,In_981,In_884);
nor U3404 (N_3404,In_614,In_113);
or U3405 (N_3405,In_470,In_182);
xor U3406 (N_3406,In_174,In_159);
and U3407 (N_3407,In_978,In_36);
nor U3408 (N_3408,In_622,In_490);
and U3409 (N_3409,In_456,In_192);
and U3410 (N_3410,In_609,In_430);
and U3411 (N_3411,In_897,In_890);
nor U3412 (N_3412,In_302,In_664);
and U3413 (N_3413,In_128,In_95);
nand U3414 (N_3414,In_305,In_905);
or U3415 (N_3415,In_238,In_111);
nand U3416 (N_3416,In_319,In_285);
or U3417 (N_3417,In_90,In_232);
or U3418 (N_3418,In_938,In_742);
nand U3419 (N_3419,In_639,In_293);
and U3420 (N_3420,In_495,In_641);
nand U3421 (N_3421,In_124,In_513);
and U3422 (N_3422,In_459,In_89);
nand U3423 (N_3423,In_202,In_78);
nor U3424 (N_3424,In_509,In_574);
nor U3425 (N_3425,In_333,In_103);
xor U3426 (N_3426,In_691,In_936);
or U3427 (N_3427,In_367,In_961);
and U3428 (N_3428,In_847,In_670);
and U3429 (N_3429,In_213,In_665);
nor U3430 (N_3430,In_385,In_995);
nor U3431 (N_3431,In_977,In_653);
nand U3432 (N_3432,In_614,In_31);
nor U3433 (N_3433,In_750,In_103);
nand U3434 (N_3434,In_893,In_680);
or U3435 (N_3435,In_73,In_274);
nand U3436 (N_3436,In_0,In_381);
or U3437 (N_3437,In_853,In_727);
nand U3438 (N_3438,In_29,In_729);
or U3439 (N_3439,In_414,In_395);
nand U3440 (N_3440,In_540,In_728);
or U3441 (N_3441,In_606,In_101);
nor U3442 (N_3442,In_25,In_706);
or U3443 (N_3443,In_555,In_586);
nor U3444 (N_3444,In_146,In_287);
and U3445 (N_3445,In_247,In_877);
nand U3446 (N_3446,In_202,In_604);
and U3447 (N_3447,In_888,In_510);
nor U3448 (N_3448,In_888,In_984);
and U3449 (N_3449,In_530,In_137);
nand U3450 (N_3450,In_590,In_811);
nor U3451 (N_3451,In_23,In_542);
or U3452 (N_3452,In_419,In_24);
or U3453 (N_3453,In_585,In_935);
nand U3454 (N_3454,In_660,In_61);
nor U3455 (N_3455,In_380,In_616);
nor U3456 (N_3456,In_413,In_412);
or U3457 (N_3457,In_385,In_758);
and U3458 (N_3458,In_669,In_776);
xor U3459 (N_3459,In_398,In_212);
and U3460 (N_3460,In_26,In_327);
nor U3461 (N_3461,In_335,In_45);
nand U3462 (N_3462,In_219,In_917);
nor U3463 (N_3463,In_301,In_967);
nor U3464 (N_3464,In_847,In_324);
and U3465 (N_3465,In_227,In_58);
nand U3466 (N_3466,In_594,In_214);
xor U3467 (N_3467,In_680,In_510);
or U3468 (N_3468,In_5,In_887);
nand U3469 (N_3469,In_715,In_215);
nand U3470 (N_3470,In_183,In_784);
xnor U3471 (N_3471,In_159,In_549);
or U3472 (N_3472,In_129,In_742);
and U3473 (N_3473,In_50,In_374);
xnor U3474 (N_3474,In_447,In_545);
and U3475 (N_3475,In_934,In_964);
nor U3476 (N_3476,In_406,In_604);
nor U3477 (N_3477,In_546,In_465);
and U3478 (N_3478,In_811,In_700);
nand U3479 (N_3479,In_567,In_364);
nor U3480 (N_3480,In_261,In_733);
and U3481 (N_3481,In_652,In_117);
xor U3482 (N_3482,In_571,In_177);
and U3483 (N_3483,In_409,In_356);
nor U3484 (N_3484,In_853,In_130);
nand U3485 (N_3485,In_85,In_711);
nand U3486 (N_3486,In_986,In_968);
nor U3487 (N_3487,In_763,In_305);
or U3488 (N_3488,In_438,In_874);
nor U3489 (N_3489,In_470,In_339);
nand U3490 (N_3490,In_15,In_667);
and U3491 (N_3491,In_234,In_660);
and U3492 (N_3492,In_271,In_483);
or U3493 (N_3493,In_313,In_441);
and U3494 (N_3494,In_504,In_95);
or U3495 (N_3495,In_394,In_568);
nand U3496 (N_3496,In_169,In_322);
or U3497 (N_3497,In_193,In_943);
nor U3498 (N_3498,In_121,In_66);
nand U3499 (N_3499,In_931,In_339);
and U3500 (N_3500,In_208,In_541);
nor U3501 (N_3501,In_384,In_474);
xnor U3502 (N_3502,In_642,In_190);
nand U3503 (N_3503,In_12,In_313);
and U3504 (N_3504,In_534,In_62);
nand U3505 (N_3505,In_808,In_161);
nor U3506 (N_3506,In_837,In_501);
nand U3507 (N_3507,In_1,In_783);
nor U3508 (N_3508,In_201,In_825);
nor U3509 (N_3509,In_889,In_192);
and U3510 (N_3510,In_980,In_664);
and U3511 (N_3511,In_884,In_305);
nand U3512 (N_3512,In_291,In_839);
or U3513 (N_3513,In_998,In_885);
nor U3514 (N_3514,In_771,In_294);
and U3515 (N_3515,In_104,In_224);
nand U3516 (N_3516,In_794,In_252);
nor U3517 (N_3517,In_721,In_973);
or U3518 (N_3518,In_105,In_169);
and U3519 (N_3519,In_556,In_999);
nand U3520 (N_3520,In_71,In_647);
and U3521 (N_3521,In_501,In_325);
or U3522 (N_3522,In_682,In_775);
nand U3523 (N_3523,In_655,In_557);
xor U3524 (N_3524,In_529,In_643);
nand U3525 (N_3525,In_353,In_9);
and U3526 (N_3526,In_777,In_636);
xnor U3527 (N_3527,In_942,In_96);
and U3528 (N_3528,In_117,In_51);
or U3529 (N_3529,In_190,In_122);
or U3530 (N_3530,In_756,In_674);
nand U3531 (N_3531,In_760,In_981);
nand U3532 (N_3532,In_930,In_743);
nor U3533 (N_3533,In_745,In_105);
and U3534 (N_3534,In_63,In_407);
or U3535 (N_3535,In_171,In_250);
nand U3536 (N_3536,In_174,In_185);
nor U3537 (N_3537,In_243,In_234);
and U3538 (N_3538,In_25,In_789);
and U3539 (N_3539,In_545,In_700);
nor U3540 (N_3540,In_228,In_664);
nand U3541 (N_3541,In_70,In_939);
or U3542 (N_3542,In_946,In_909);
and U3543 (N_3543,In_493,In_872);
nand U3544 (N_3544,In_590,In_606);
xor U3545 (N_3545,In_671,In_858);
or U3546 (N_3546,In_334,In_457);
or U3547 (N_3547,In_772,In_567);
and U3548 (N_3548,In_379,In_878);
or U3549 (N_3549,In_223,In_939);
nand U3550 (N_3550,In_576,In_277);
nand U3551 (N_3551,In_557,In_476);
nand U3552 (N_3552,In_143,In_647);
nand U3553 (N_3553,In_565,In_240);
and U3554 (N_3554,In_668,In_826);
nor U3555 (N_3555,In_856,In_565);
or U3556 (N_3556,In_371,In_677);
or U3557 (N_3557,In_348,In_904);
and U3558 (N_3558,In_436,In_942);
nor U3559 (N_3559,In_564,In_495);
nand U3560 (N_3560,In_904,In_129);
or U3561 (N_3561,In_210,In_769);
nand U3562 (N_3562,In_655,In_986);
and U3563 (N_3563,In_967,In_871);
nor U3564 (N_3564,In_264,In_692);
nand U3565 (N_3565,In_837,In_823);
or U3566 (N_3566,In_884,In_108);
nand U3567 (N_3567,In_349,In_430);
and U3568 (N_3568,In_855,In_516);
and U3569 (N_3569,In_908,In_902);
and U3570 (N_3570,In_671,In_81);
nand U3571 (N_3571,In_833,In_614);
nand U3572 (N_3572,In_328,In_431);
nand U3573 (N_3573,In_370,In_866);
or U3574 (N_3574,In_72,In_502);
or U3575 (N_3575,In_429,In_888);
and U3576 (N_3576,In_314,In_351);
xor U3577 (N_3577,In_75,In_623);
nor U3578 (N_3578,In_62,In_364);
and U3579 (N_3579,In_183,In_420);
or U3580 (N_3580,In_331,In_89);
and U3581 (N_3581,In_960,In_275);
nand U3582 (N_3582,In_531,In_163);
nor U3583 (N_3583,In_40,In_619);
or U3584 (N_3584,In_131,In_178);
or U3585 (N_3585,In_575,In_391);
or U3586 (N_3586,In_239,In_923);
nor U3587 (N_3587,In_835,In_196);
nand U3588 (N_3588,In_419,In_876);
and U3589 (N_3589,In_73,In_395);
nor U3590 (N_3590,In_908,In_774);
and U3591 (N_3591,In_455,In_906);
nor U3592 (N_3592,In_640,In_600);
nand U3593 (N_3593,In_624,In_274);
and U3594 (N_3594,In_663,In_96);
nand U3595 (N_3595,In_482,In_848);
nor U3596 (N_3596,In_323,In_946);
xnor U3597 (N_3597,In_142,In_267);
xnor U3598 (N_3598,In_440,In_624);
xor U3599 (N_3599,In_284,In_528);
nor U3600 (N_3600,In_185,In_924);
nand U3601 (N_3601,In_135,In_284);
and U3602 (N_3602,In_961,In_178);
and U3603 (N_3603,In_639,In_83);
and U3604 (N_3604,In_97,In_341);
or U3605 (N_3605,In_730,In_883);
or U3606 (N_3606,In_33,In_728);
nand U3607 (N_3607,In_761,In_645);
and U3608 (N_3608,In_444,In_92);
nand U3609 (N_3609,In_438,In_720);
or U3610 (N_3610,In_470,In_289);
nor U3611 (N_3611,In_778,In_78);
xnor U3612 (N_3612,In_326,In_549);
xnor U3613 (N_3613,In_504,In_357);
nand U3614 (N_3614,In_978,In_340);
and U3615 (N_3615,In_363,In_609);
nor U3616 (N_3616,In_205,In_254);
and U3617 (N_3617,In_740,In_45);
nor U3618 (N_3618,In_417,In_633);
and U3619 (N_3619,In_797,In_581);
nor U3620 (N_3620,In_404,In_913);
nor U3621 (N_3621,In_476,In_372);
or U3622 (N_3622,In_102,In_991);
and U3623 (N_3623,In_26,In_287);
xnor U3624 (N_3624,In_391,In_885);
nor U3625 (N_3625,In_637,In_290);
and U3626 (N_3626,In_716,In_146);
and U3627 (N_3627,In_439,In_825);
nor U3628 (N_3628,In_371,In_817);
or U3629 (N_3629,In_767,In_148);
xor U3630 (N_3630,In_763,In_710);
nand U3631 (N_3631,In_679,In_849);
and U3632 (N_3632,In_443,In_378);
nor U3633 (N_3633,In_968,In_777);
xor U3634 (N_3634,In_140,In_405);
or U3635 (N_3635,In_135,In_597);
nor U3636 (N_3636,In_795,In_794);
and U3637 (N_3637,In_182,In_854);
or U3638 (N_3638,In_153,In_620);
nand U3639 (N_3639,In_248,In_0);
or U3640 (N_3640,In_435,In_865);
nand U3641 (N_3641,In_335,In_122);
nand U3642 (N_3642,In_779,In_681);
and U3643 (N_3643,In_963,In_120);
or U3644 (N_3644,In_889,In_965);
xnor U3645 (N_3645,In_587,In_173);
or U3646 (N_3646,In_220,In_838);
and U3647 (N_3647,In_55,In_493);
and U3648 (N_3648,In_979,In_533);
nand U3649 (N_3649,In_587,In_725);
and U3650 (N_3650,In_941,In_655);
or U3651 (N_3651,In_888,In_110);
or U3652 (N_3652,In_733,In_667);
and U3653 (N_3653,In_726,In_781);
nand U3654 (N_3654,In_473,In_577);
xor U3655 (N_3655,In_216,In_992);
nand U3656 (N_3656,In_12,In_739);
or U3657 (N_3657,In_240,In_632);
or U3658 (N_3658,In_173,In_247);
nand U3659 (N_3659,In_367,In_24);
and U3660 (N_3660,In_65,In_432);
xnor U3661 (N_3661,In_556,In_674);
nor U3662 (N_3662,In_111,In_900);
nor U3663 (N_3663,In_389,In_128);
xor U3664 (N_3664,In_943,In_469);
xor U3665 (N_3665,In_608,In_552);
and U3666 (N_3666,In_618,In_405);
nor U3667 (N_3667,In_831,In_690);
or U3668 (N_3668,In_288,In_437);
nor U3669 (N_3669,In_220,In_135);
nor U3670 (N_3670,In_57,In_943);
nor U3671 (N_3671,In_586,In_189);
and U3672 (N_3672,In_911,In_345);
nand U3673 (N_3673,In_243,In_51);
nor U3674 (N_3674,In_939,In_804);
nand U3675 (N_3675,In_52,In_239);
xor U3676 (N_3676,In_583,In_552);
and U3677 (N_3677,In_509,In_54);
nor U3678 (N_3678,In_963,In_16);
nand U3679 (N_3679,In_964,In_160);
and U3680 (N_3680,In_262,In_205);
nand U3681 (N_3681,In_507,In_340);
nor U3682 (N_3682,In_191,In_273);
or U3683 (N_3683,In_615,In_812);
and U3684 (N_3684,In_139,In_864);
nor U3685 (N_3685,In_731,In_195);
nor U3686 (N_3686,In_313,In_558);
and U3687 (N_3687,In_353,In_629);
and U3688 (N_3688,In_359,In_845);
or U3689 (N_3689,In_218,In_264);
nor U3690 (N_3690,In_401,In_612);
and U3691 (N_3691,In_648,In_847);
nor U3692 (N_3692,In_578,In_653);
or U3693 (N_3693,In_703,In_916);
nand U3694 (N_3694,In_817,In_109);
and U3695 (N_3695,In_806,In_576);
and U3696 (N_3696,In_897,In_513);
nor U3697 (N_3697,In_353,In_76);
and U3698 (N_3698,In_23,In_71);
xor U3699 (N_3699,In_792,In_686);
or U3700 (N_3700,In_505,In_345);
nor U3701 (N_3701,In_340,In_470);
nor U3702 (N_3702,In_568,In_526);
nor U3703 (N_3703,In_924,In_599);
nor U3704 (N_3704,In_921,In_88);
and U3705 (N_3705,In_174,In_35);
and U3706 (N_3706,In_221,In_926);
and U3707 (N_3707,In_254,In_799);
and U3708 (N_3708,In_778,In_522);
or U3709 (N_3709,In_192,In_176);
nor U3710 (N_3710,In_232,In_754);
and U3711 (N_3711,In_75,In_68);
nand U3712 (N_3712,In_952,In_190);
and U3713 (N_3713,In_821,In_60);
or U3714 (N_3714,In_436,In_851);
nor U3715 (N_3715,In_62,In_763);
nor U3716 (N_3716,In_772,In_23);
nor U3717 (N_3717,In_225,In_626);
xnor U3718 (N_3718,In_296,In_143);
nand U3719 (N_3719,In_221,In_806);
or U3720 (N_3720,In_605,In_784);
or U3721 (N_3721,In_416,In_737);
nand U3722 (N_3722,In_225,In_131);
and U3723 (N_3723,In_747,In_583);
nand U3724 (N_3724,In_812,In_713);
nand U3725 (N_3725,In_486,In_424);
xor U3726 (N_3726,In_844,In_559);
nand U3727 (N_3727,In_374,In_397);
or U3728 (N_3728,In_648,In_859);
nor U3729 (N_3729,In_676,In_221);
and U3730 (N_3730,In_974,In_85);
nand U3731 (N_3731,In_168,In_181);
nor U3732 (N_3732,In_686,In_877);
nand U3733 (N_3733,In_97,In_914);
or U3734 (N_3734,In_171,In_780);
nand U3735 (N_3735,In_216,In_672);
nand U3736 (N_3736,In_222,In_540);
nor U3737 (N_3737,In_645,In_9);
nand U3738 (N_3738,In_963,In_553);
xor U3739 (N_3739,In_608,In_396);
nor U3740 (N_3740,In_99,In_534);
or U3741 (N_3741,In_608,In_88);
nor U3742 (N_3742,In_361,In_513);
nor U3743 (N_3743,In_522,In_949);
nor U3744 (N_3744,In_54,In_845);
or U3745 (N_3745,In_205,In_909);
nor U3746 (N_3746,In_708,In_655);
nand U3747 (N_3747,In_368,In_439);
nand U3748 (N_3748,In_790,In_530);
or U3749 (N_3749,In_950,In_549);
nand U3750 (N_3750,In_549,In_762);
nor U3751 (N_3751,In_256,In_69);
and U3752 (N_3752,In_747,In_621);
nand U3753 (N_3753,In_245,In_484);
and U3754 (N_3754,In_476,In_976);
xnor U3755 (N_3755,In_599,In_492);
and U3756 (N_3756,In_768,In_537);
nand U3757 (N_3757,In_880,In_952);
nor U3758 (N_3758,In_7,In_579);
nor U3759 (N_3759,In_774,In_916);
nor U3760 (N_3760,In_785,In_780);
and U3761 (N_3761,In_120,In_753);
nor U3762 (N_3762,In_553,In_917);
and U3763 (N_3763,In_337,In_193);
and U3764 (N_3764,In_587,In_568);
and U3765 (N_3765,In_429,In_701);
and U3766 (N_3766,In_92,In_660);
nand U3767 (N_3767,In_574,In_52);
nand U3768 (N_3768,In_288,In_669);
nor U3769 (N_3769,In_784,In_545);
nor U3770 (N_3770,In_229,In_455);
nand U3771 (N_3771,In_385,In_683);
nand U3772 (N_3772,In_529,In_787);
nor U3773 (N_3773,In_972,In_744);
or U3774 (N_3774,In_735,In_109);
nor U3775 (N_3775,In_603,In_620);
and U3776 (N_3776,In_677,In_690);
and U3777 (N_3777,In_95,In_145);
nor U3778 (N_3778,In_945,In_883);
or U3779 (N_3779,In_463,In_197);
or U3780 (N_3780,In_283,In_771);
nor U3781 (N_3781,In_318,In_90);
nand U3782 (N_3782,In_836,In_547);
and U3783 (N_3783,In_222,In_908);
and U3784 (N_3784,In_433,In_901);
xnor U3785 (N_3785,In_804,In_135);
nand U3786 (N_3786,In_183,In_243);
xor U3787 (N_3787,In_864,In_994);
nor U3788 (N_3788,In_797,In_800);
or U3789 (N_3789,In_135,In_69);
and U3790 (N_3790,In_37,In_221);
and U3791 (N_3791,In_970,In_952);
nor U3792 (N_3792,In_41,In_69);
and U3793 (N_3793,In_453,In_682);
and U3794 (N_3794,In_490,In_100);
nand U3795 (N_3795,In_273,In_688);
and U3796 (N_3796,In_755,In_839);
or U3797 (N_3797,In_903,In_170);
nor U3798 (N_3798,In_366,In_322);
nand U3799 (N_3799,In_195,In_386);
nor U3800 (N_3800,In_38,In_695);
or U3801 (N_3801,In_202,In_20);
nand U3802 (N_3802,In_285,In_993);
xnor U3803 (N_3803,In_42,In_280);
nand U3804 (N_3804,In_318,In_769);
xnor U3805 (N_3805,In_716,In_689);
nand U3806 (N_3806,In_528,In_997);
nand U3807 (N_3807,In_221,In_384);
nor U3808 (N_3808,In_123,In_487);
nor U3809 (N_3809,In_646,In_642);
xnor U3810 (N_3810,In_571,In_375);
or U3811 (N_3811,In_25,In_263);
xor U3812 (N_3812,In_936,In_27);
and U3813 (N_3813,In_150,In_21);
nand U3814 (N_3814,In_142,In_201);
nand U3815 (N_3815,In_650,In_641);
nand U3816 (N_3816,In_252,In_309);
and U3817 (N_3817,In_502,In_337);
xor U3818 (N_3818,In_385,In_251);
nand U3819 (N_3819,In_632,In_407);
nand U3820 (N_3820,In_295,In_906);
nor U3821 (N_3821,In_778,In_708);
or U3822 (N_3822,In_868,In_839);
and U3823 (N_3823,In_387,In_972);
nor U3824 (N_3824,In_870,In_485);
nor U3825 (N_3825,In_176,In_10);
or U3826 (N_3826,In_310,In_309);
and U3827 (N_3827,In_747,In_286);
nand U3828 (N_3828,In_688,In_712);
xor U3829 (N_3829,In_645,In_28);
or U3830 (N_3830,In_876,In_549);
nor U3831 (N_3831,In_669,In_233);
nor U3832 (N_3832,In_320,In_991);
xor U3833 (N_3833,In_329,In_263);
nor U3834 (N_3834,In_412,In_264);
nand U3835 (N_3835,In_572,In_472);
nor U3836 (N_3836,In_686,In_788);
or U3837 (N_3837,In_578,In_92);
nor U3838 (N_3838,In_723,In_439);
nor U3839 (N_3839,In_808,In_982);
nor U3840 (N_3840,In_768,In_363);
nand U3841 (N_3841,In_672,In_577);
nand U3842 (N_3842,In_529,In_134);
or U3843 (N_3843,In_744,In_358);
nand U3844 (N_3844,In_318,In_151);
nand U3845 (N_3845,In_134,In_889);
nand U3846 (N_3846,In_522,In_137);
nor U3847 (N_3847,In_294,In_429);
nand U3848 (N_3848,In_268,In_507);
nor U3849 (N_3849,In_75,In_409);
nand U3850 (N_3850,In_620,In_913);
nand U3851 (N_3851,In_160,In_411);
or U3852 (N_3852,In_945,In_725);
and U3853 (N_3853,In_692,In_469);
and U3854 (N_3854,In_677,In_336);
nand U3855 (N_3855,In_27,In_376);
and U3856 (N_3856,In_391,In_410);
xnor U3857 (N_3857,In_170,In_84);
and U3858 (N_3858,In_58,In_473);
and U3859 (N_3859,In_241,In_467);
and U3860 (N_3860,In_295,In_631);
and U3861 (N_3861,In_113,In_617);
nor U3862 (N_3862,In_951,In_358);
or U3863 (N_3863,In_526,In_628);
nand U3864 (N_3864,In_136,In_155);
nand U3865 (N_3865,In_183,In_828);
and U3866 (N_3866,In_732,In_272);
and U3867 (N_3867,In_406,In_379);
nand U3868 (N_3868,In_852,In_575);
nand U3869 (N_3869,In_12,In_227);
or U3870 (N_3870,In_878,In_127);
nand U3871 (N_3871,In_454,In_416);
xnor U3872 (N_3872,In_20,In_328);
and U3873 (N_3873,In_646,In_561);
or U3874 (N_3874,In_724,In_356);
nand U3875 (N_3875,In_884,In_713);
or U3876 (N_3876,In_445,In_540);
nand U3877 (N_3877,In_475,In_250);
and U3878 (N_3878,In_51,In_718);
nand U3879 (N_3879,In_336,In_837);
or U3880 (N_3880,In_562,In_277);
and U3881 (N_3881,In_987,In_694);
xor U3882 (N_3882,In_559,In_952);
nor U3883 (N_3883,In_500,In_655);
nand U3884 (N_3884,In_200,In_621);
and U3885 (N_3885,In_969,In_370);
and U3886 (N_3886,In_249,In_386);
nor U3887 (N_3887,In_961,In_513);
or U3888 (N_3888,In_225,In_632);
and U3889 (N_3889,In_709,In_816);
and U3890 (N_3890,In_42,In_739);
or U3891 (N_3891,In_401,In_649);
xor U3892 (N_3892,In_326,In_126);
xnor U3893 (N_3893,In_676,In_167);
nand U3894 (N_3894,In_859,In_924);
or U3895 (N_3895,In_709,In_121);
and U3896 (N_3896,In_631,In_866);
and U3897 (N_3897,In_78,In_215);
nand U3898 (N_3898,In_391,In_913);
nand U3899 (N_3899,In_729,In_276);
nand U3900 (N_3900,In_903,In_797);
nand U3901 (N_3901,In_23,In_899);
xor U3902 (N_3902,In_340,In_781);
nor U3903 (N_3903,In_350,In_62);
nand U3904 (N_3904,In_106,In_912);
nor U3905 (N_3905,In_334,In_350);
and U3906 (N_3906,In_362,In_436);
or U3907 (N_3907,In_87,In_600);
and U3908 (N_3908,In_471,In_4);
or U3909 (N_3909,In_120,In_700);
nor U3910 (N_3910,In_848,In_355);
nand U3911 (N_3911,In_555,In_723);
and U3912 (N_3912,In_523,In_244);
and U3913 (N_3913,In_98,In_562);
and U3914 (N_3914,In_956,In_8);
nor U3915 (N_3915,In_867,In_141);
and U3916 (N_3916,In_313,In_984);
nand U3917 (N_3917,In_591,In_513);
xnor U3918 (N_3918,In_545,In_266);
and U3919 (N_3919,In_584,In_611);
nand U3920 (N_3920,In_932,In_815);
nor U3921 (N_3921,In_629,In_814);
xor U3922 (N_3922,In_821,In_220);
or U3923 (N_3923,In_212,In_572);
nand U3924 (N_3924,In_913,In_677);
and U3925 (N_3925,In_251,In_498);
xnor U3926 (N_3926,In_982,In_7);
nand U3927 (N_3927,In_926,In_664);
or U3928 (N_3928,In_491,In_558);
or U3929 (N_3929,In_982,In_755);
nor U3930 (N_3930,In_365,In_387);
xnor U3931 (N_3931,In_260,In_103);
and U3932 (N_3932,In_864,In_993);
nand U3933 (N_3933,In_765,In_720);
nor U3934 (N_3934,In_611,In_144);
and U3935 (N_3935,In_342,In_273);
or U3936 (N_3936,In_898,In_554);
or U3937 (N_3937,In_396,In_502);
and U3938 (N_3938,In_862,In_360);
or U3939 (N_3939,In_937,In_149);
xnor U3940 (N_3940,In_499,In_469);
and U3941 (N_3941,In_689,In_908);
and U3942 (N_3942,In_62,In_231);
or U3943 (N_3943,In_612,In_72);
nand U3944 (N_3944,In_349,In_264);
and U3945 (N_3945,In_566,In_406);
nor U3946 (N_3946,In_556,In_395);
nand U3947 (N_3947,In_38,In_988);
nand U3948 (N_3948,In_512,In_921);
nand U3949 (N_3949,In_691,In_377);
nand U3950 (N_3950,In_894,In_379);
xnor U3951 (N_3951,In_256,In_897);
and U3952 (N_3952,In_14,In_116);
and U3953 (N_3953,In_676,In_767);
or U3954 (N_3954,In_761,In_580);
and U3955 (N_3955,In_610,In_77);
nor U3956 (N_3956,In_477,In_665);
and U3957 (N_3957,In_449,In_587);
and U3958 (N_3958,In_292,In_556);
xor U3959 (N_3959,In_535,In_418);
and U3960 (N_3960,In_851,In_131);
or U3961 (N_3961,In_830,In_938);
nor U3962 (N_3962,In_448,In_496);
nand U3963 (N_3963,In_594,In_235);
nor U3964 (N_3964,In_495,In_111);
nand U3965 (N_3965,In_862,In_435);
and U3966 (N_3966,In_906,In_103);
nor U3967 (N_3967,In_188,In_810);
xor U3968 (N_3968,In_353,In_120);
and U3969 (N_3969,In_383,In_12);
nand U3970 (N_3970,In_690,In_901);
nor U3971 (N_3971,In_870,In_444);
nor U3972 (N_3972,In_382,In_341);
or U3973 (N_3973,In_487,In_468);
and U3974 (N_3974,In_858,In_863);
and U3975 (N_3975,In_142,In_330);
nor U3976 (N_3976,In_848,In_820);
and U3977 (N_3977,In_592,In_517);
or U3978 (N_3978,In_875,In_187);
and U3979 (N_3979,In_675,In_827);
nor U3980 (N_3980,In_333,In_485);
or U3981 (N_3981,In_936,In_510);
nor U3982 (N_3982,In_333,In_218);
nand U3983 (N_3983,In_651,In_23);
and U3984 (N_3984,In_852,In_862);
or U3985 (N_3985,In_51,In_691);
and U3986 (N_3986,In_202,In_868);
or U3987 (N_3987,In_601,In_221);
xor U3988 (N_3988,In_371,In_899);
nand U3989 (N_3989,In_281,In_816);
nor U3990 (N_3990,In_879,In_959);
nand U3991 (N_3991,In_354,In_54);
xnor U3992 (N_3992,In_957,In_719);
or U3993 (N_3993,In_465,In_878);
nor U3994 (N_3994,In_181,In_362);
or U3995 (N_3995,In_621,In_638);
nor U3996 (N_3996,In_516,In_849);
or U3997 (N_3997,In_776,In_35);
nor U3998 (N_3998,In_691,In_248);
nor U3999 (N_3999,In_310,In_177);
and U4000 (N_4000,In_356,In_433);
nand U4001 (N_4001,In_701,In_96);
and U4002 (N_4002,In_895,In_649);
or U4003 (N_4003,In_727,In_399);
nor U4004 (N_4004,In_196,In_993);
or U4005 (N_4005,In_298,In_424);
or U4006 (N_4006,In_824,In_232);
and U4007 (N_4007,In_274,In_125);
and U4008 (N_4008,In_886,In_154);
nor U4009 (N_4009,In_31,In_633);
nand U4010 (N_4010,In_424,In_430);
nand U4011 (N_4011,In_684,In_988);
nand U4012 (N_4012,In_211,In_837);
and U4013 (N_4013,In_452,In_265);
nor U4014 (N_4014,In_466,In_793);
nor U4015 (N_4015,In_178,In_155);
xor U4016 (N_4016,In_761,In_260);
and U4017 (N_4017,In_906,In_996);
xor U4018 (N_4018,In_873,In_511);
and U4019 (N_4019,In_157,In_810);
xor U4020 (N_4020,In_885,In_349);
or U4021 (N_4021,In_638,In_686);
nand U4022 (N_4022,In_625,In_411);
and U4023 (N_4023,In_578,In_955);
and U4024 (N_4024,In_1,In_628);
nand U4025 (N_4025,In_404,In_579);
and U4026 (N_4026,In_995,In_535);
nor U4027 (N_4027,In_827,In_423);
or U4028 (N_4028,In_8,In_232);
and U4029 (N_4029,In_657,In_780);
and U4030 (N_4030,In_684,In_980);
nor U4031 (N_4031,In_408,In_750);
and U4032 (N_4032,In_781,In_861);
or U4033 (N_4033,In_482,In_681);
xor U4034 (N_4034,In_613,In_299);
and U4035 (N_4035,In_979,In_281);
nand U4036 (N_4036,In_416,In_278);
nor U4037 (N_4037,In_149,In_692);
xor U4038 (N_4038,In_234,In_641);
xor U4039 (N_4039,In_478,In_454);
and U4040 (N_4040,In_773,In_879);
nor U4041 (N_4041,In_345,In_261);
or U4042 (N_4042,In_99,In_819);
nand U4043 (N_4043,In_139,In_33);
nor U4044 (N_4044,In_876,In_739);
nand U4045 (N_4045,In_624,In_899);
or U4046 (N_4046,In_266,In_194);
nor U4047 (N_4047,In_469,In_834);
or U4048 (N_4048,In_44,In_25);
nand U4049 (N_4049,In_641,In_273);
nand U4050 (N_4050,In_619,In_973);
and U4051 (N_4051,In_877,In_561);
or U4052 (N_4052,In_957,In_284);
xnor U4053 (N_4053,In_525,In_533);
and U4054 (N_4054,In_335,In_233);
nand U4055 (N_4055,In_117,In_306);
nand U4056 (N_4056,In_661,In_820);
nand U4057 (N_4057,In_544,In_96);
xnor U4058 (N_4058,In_664,In_421);
or U4059 (N_4059,In_901,In_811);
or U4060 (N_4060,In_37,In_837);
nor U4061 (N_4061,In_943,In_650);
or U4062 (N_4062,In_773,In_32);
xor U4063 (N_4063,In_775,In_987);
or U4064 (N_4064,In_370,In_430);
or U4065 (N_4065,In_395,In_746);
and U4066 (N_4066,In_804,In_838);
xor U4067 (N_4067,In_688,In_662);
nor U4068 (N_4068,In_366,In_794);
or U4069 (N_4069,In_130,In_636);
nand U4070 (N_4070,In_717,In_556);
nand U4071 (N_4071,In_575,In_962);
nand U4072 (N_4072,In_864,In_860);
xor U4073 (N_4073,In_207,In_879);
nor U4074 (N_4074,In_762,In_408);
or U4075 (N_4075,In_4,In_170);
xnor U4076 (N_4076,In_387,In_888);
or U4077 (N_4077,In_122,In_939);
nand U4078 (N_4078,In_305,In_30);
nand U4079 (N_4079,In_235,In_194);
and U4080 (N_4080,In_259,In_205);
nand U4081 (N_4081,In_645,In_966);
xor U4082 (N_4082,In_275,In_937);
nand U4083 (N_4083,In_132,In_380);
nand U4084 (N_4084,In_609,In_629);
or U4085 (N_4085,In_453,In_224);
and U4086 (N_4086,In_787,In_176);
nand U4087 (N_4087,In_449,In_750);
and U4088 (N_4088,In_372,In_210);
nor U4089 (N_4089,In_683,In_414);
or U4090 (N_4090,In_158,In_328);
nor U4091 (N_4091,In_42,In_268);
nor U4092 (N_4092,In_628,In_205);
or U4093 (N_4093,In_855,In_499);
nor U4094 (N_4094,In_486,In_816);
or U4095 (N_4095,In_726,In_533);
nor U4096 (N_4096,In_702,In_77);
nor U4097 (N_4097,In_735,In_395);
and U4098 (N_4098,In_193,In_757);
xnor U4099 (N_4099,In_788,In_376);
or U4100 (N_4100,In_137,In_92);
nand U4101 (N_4101,In_37,In_32);
nor U4102 (N_4102,In_503,In_694);
nand U4103 (N_4103,In_579,In_982);
nand U4104 (N_4104,In_513,In_943);
and U4105 (N_4105,In_612,In_379);
xnor U4106 (N_4106,In_719,In_876);
and U4107 (N_4107,In_739,In_614);
nand U4108 (N_4108,In_257,In_986);
and U4109 (N_4109,In_313,In_847);
or U4110 (N_4110,In_759,In_227);
nand U4111 (N_4111,In_863,In_467);
and U4112 (N_4112,In_638,In_170);
xor U4113 (N_4113,In_822,In_2);
and U4114 (N_4114,In_793,In_732);
nor U4115 (N_4115,In_41,In_901);
or U4116 (N_4116,In_532,In_376);
nand U4117 (N_4117,In_442,In_202);
or U4118 (N_4118,In_935,In_322);
or U4119 (N_4119,In_694,In_619);
xnor U4120 (N_4120,In_174,In_573);
and U4121 (N_4121,In_82,In_838);
nor U4122 (N_4122,In_109,In_514);
xor U4123 (N_4123,In_795,In_289);
or U4124 (N_4124,In_992,In_658);
or U4125 (N_4125,In_724,In_427);
and U4126 (N_4126,In_715,In_347);
and U4127 (N_4127,In_354,In_822);
or U4128 (N_4128,In_427,In_135);
nand U4129 (N_4129,In_656,In_59);
nand U4130 (N_4130,In_998,In_650);
nor U4131 (N_4131,In_565,In_0);
xor U4132 (N_4132,In_819,In_835);
nand U4133 (N_4133,In_904,In_279);
or U4134 (N_4134,In_78,In_153);
and U4135 (N_4135,In_9,In_203);
xnor U4136 (N_4136,In_942,In_144);
and U4137 (N_4137,In_552,In_795);
or U4138 (N_4138,In_881,In_748);
xnor U4139 (N_4139,In_614,In_158);
nor U4140 (N_4140,In_577,In_587);
nor U4141 (N_4141,In_984,In_535);
nor U4142 (N_4142,In_164,In_589);
nand U4143 (N_4143,In_131,In_743);
nand U4144 (N_4144,In_403,In_81);
nand U4145 (N_4145,In_754,In_622);
and U4146 (N_4146,In_484,In_100);
and U4147 (N_4147,In_544,In_895);
nand U4148 (N_4148,In_425,In_680);
and U4149 (N_4149,In_633,In_467);
nor U4150 (N_4150,In_794,In_83);
xnor U4151 (N_4151,In_73,In_964);
nor U4152 (N_4152,In_573,In_348);
nor U4153 (N_4153,In_217,In_515);
nand U4154 (N_4154,In_569,In_63);
and U4155 (N_4155,In_192,In_680);
or U4156 (N_4156,In_527,In_670);
nand U4157 (N_4157,In_391,In_513);
or U4158 (N_4158,In_93,In_198);
or U4159 (N_4159,In_788,In_635);
nor U4160 (N_4160,In_771,In_78);
or U4161 (N_4161,In_477,In_850);
nor U4162 (N_4162,In_470,In_667);
and U4163 (N_4163,In_803,In_599);
nand U4164 (N_4164,In_14,In_187);
or U4165 (N_4165,In_438,In_87);
nand U4166 (N_4166,In_819,In_940);
xnor U4167 (N_4167,In_172,In_196);
and U4168 (N_4168,In_640,In_294);
nor U4169 (N_4169,In_251,In_450);
and U4170 (N_4170,In_927,In_656);
nand U4171 (N_4171,In_407,In_312);
nand U4172 (N_4172,In_298,In_483);
or U4173 (N_4173,In_356,In_479);
nor U4174 (N_4174,In_309,In_919);
nand U4175 (N_4175,In_63,In_152);
nand U4176 (N_4176,In_255,In_83);
and U4177 (N_4177,In_491,In_555);
and U4178 (N_4178,In_519,In_433);
nand U4179 (N_4179,In_867,In_635);
nand U4180 (N_4180,In_363,In_946);
or U4181 (N_4181,In_935,In_836);
nor U4182 (N_4182,In_792,In_201);
nor U4183 (N_4183,In_579,In_659);
xor U4184 (N_4184,In_323,In_142);
or U4185 (N_4185,In_743,In_861);
and U4186 (N_4186,In_952,In_831);
or U4187 (N_4187,In_77,In_670);
or U4188 (N_4188,In_48,In_472);
xnor U4189 (N_4189,In_744,In_264);
nor U4190 (N_4190,In_838,In_996);
nand U4191 (N_4191,In_258,In_895);
nor U4192 (N_4192,In_73,In_544);
xnor U4193 (N_4193,In_304,In_52);
xnor U4194 (N_4194,In_281,In_341);
xor U4195 (N_4195,In_668,In_775);
and U4196 (N_4196,In_80,In_298);
or U4197 (N_4197,In_994,In_295);
nor U4198 (N_4198,In_238,In_91);
and U4199 (N_4199,In_146,In_792);
xnor U4200 (N_4200,In_38,In_984);
nand U4201 (N_4201,In_110,In_725);
nand U4202 (N_4202,In_955,In_506);
or U4203 (N_4203,In_959,In_322);
and U4204 (N_4204,In_136,In_218);
or U4205 (N_4205,In_260,In_622);
nor U4206 (N_4206,In_113,In_434);
and U4207 (N_4207,In_420,In_703);
nor U4208 (N_4208,In_373,In_893);
xnor U4209 (N_4209,In_889,In_807);
or U4210 (N_4210,In_724,In_364);
or U4211 (N_4211,In_749,In_722);
or U4212 (N_4212,In_471,In_144);
or U4213 (N_4213,In_926,In_893);
nand U4214 (N_4214,In_627,In_60);
and U4215 (N_4215,In_16,In_667);
xor U4216 (N_4216,In_312,In_322);
or U4217 (N_4217,In_113,In_496);
and U4218 (N_4218,In_86,In_886);
and U4219 (N_4219,In_480,In_994);
and U4220 (N_4220,In_208,In_834);
and U4221 (N_4221,In_302,In_934);
nand U4222 (N_4222,In_901,In_253);
xnor U4223 (N_4223,In_544,In_818);
or U4224 (N_4224,In_893,In_654);
and U4225 (N_4225,In_350,In_557);
nor U4226 (N_4226,In_736,In_123);
xor U4227 (N_4227,In_628,In_844);
or U4228 (N_4228,In_931,In_769);
or U4229 (N_4229,In_607,In_224);
nand U4230 (N_4230,In_949,In_295);
nand U4231 (N_4231,In_858,In_159);
nand U4232 (N_4232,In_919,In_579);
and U4233 (N_4233,In_777,In_723);
nor U4234 (N_4234,In_684,In_258);
nor U4235 (N_4235,In_540,In_1);
nand U4236 (N_4236,In_82,In_361);
or U4237 (N_4237,In_923,In_709);
and U4238 (N_4238,In_238,In_663);
nor U4239 (N_4239,In_575,In_975);
nor U4240 (N_4240,In_920,In_423);
and U4241 (N_4241,In_380,In_714);
nand U4242 (N_4242,In_491,In_451);
or U4243 (N_4243,In_509,In_948);
nor U4244 (N_4244,In_641,In_385);
and U4245 (N_4245,In_632,In_781);
and U4246 (N_4246,In_38,In_813);
and U4247 (N_4247,In_494,In_900);
nor U4248 (N_4248,In_72,In_301);
nor U4249 (N_4249,In_956,In_873);
nor U4250 (N_4250,In_720,In_99);
nand U4251 (N_4251,In_676,In_481);
nor U4252 (N_4252,In_708,In_537);
or U4253 (N_4253,In_343,In_799);
nand U4254 (N_4254,In_208,In_296);
nor U4255 (N_4255,In_494,In_375);
nand U4256 (N_4256,In_148,In_116);
or U4257 (N_4257,In_67,In_216);
and U4258 (N_4258,In_548,In_342);
nor U4259 (N_4259,In_455,In_468);
nor U4260 (N_4260,In_305,In_840);
and U4261 (N_4261,In_318,In_393);
nand U4262 (N_4262,In_114,In_669);
or U4263 (N_4263,In_39,In_470);
nand U4264 (N_4264,In_475,In_224);
or U4265 (N_4265,In_409,In_569);
nand U4266 (N_4266,In_5,In_709);
nand U4267 (N_4267,In_215,In_595);
or U4268 (N_4268,In_982,In_485);
xor U4269 (N_4269,In_101,In_314);
nor U4270 (N_4270,In_898,In_141);
nor U4271 (N_4271,In_530,In_121);
xor U4272 (N_4272,In_978,In_434);
and U4273 (N_4273,In_0,In_300);
or U4274 (N_4274,In_851,In_421);
and U4275 (N_4275,In_105,In_600);
xor U4276 (N_4276,In_870,In_461);
or U4277 (N_4277,In_46,In_302);
and U4278 (N_4278,In_195,In_769);
and U4279 (N_4279,In_492,In_153);
and U4280 (N_4280,In_126,In_351);
and U4281 (N_4281,In_824,In_592);
nor U4282 (N_4282,In_546,In_681);
and U4283 (N_4283,In_487,In_121);
xnor U4284 (N_4284,In_346,In_936);
or U4285 (N_4285,In_963,In_953);
and U4286 (N_4286,In_570,In_396);
nand U4287 (N_4287,In_377,In_768);
and U4288 (N_4288,In_612,In_837);
and U4289 (N_4289,In_93,In_813);
nand U4290 (N_4290,In_921,In_502);
nor U4291 (N_4291,In_112,In_432);
or U4292 (N_4292,In_466,In_760);
nand U4293 (N_4293,In_163,In_629);
or U4294 (N_4294,In_173,In_168);
nand U4295 (N_4295,In_555,In_823);
and U4296 (N_4296,In_514,In_268);
nand U4297 (N_4297,In_720,In_217);
nor U4298 (N_4298,In_285,In_146);
nor U4299 (N_4299,In_452,In_752);
or U4300 (N_4300,In_268,In_136);
or U4301 (N_4301,In_189,In_509);
and U4302 (N_4302,In_643,In_424);
and U4303 (N_4303,In_502,In_46);
nand U4304 (N_4304,In_856,In_216);
or U4305 (N_4305,In_947,In_998);
xnor U4306 (N_4306,In_858,In_453);
xor U4307 (N_4307,In_640,In_334);
nand U4308 (N_4308,In_758,In_199);
nand U4309 (N_4309,In_705,In_569);
and U4310 (N_4310,In_752,In_690);
or U4311 (N_4311,In_9,In_857);
nand U4312 (N_4312,In_148,In_152);
nor U4313 (N_4313,In_862,In_189);
nor U4314 (N_4314,In_713,In_542);
or U4315 (N_4315,In_237,In_196);
xnor U4316 (N_4316,In_156,In_13);
nor U4317 (N_4317,In_127,In_880);
or U4318 (N_4318,In_418,In_815);
nand U4319 (N_4319,In_546,In_853);
or U4320 (N_4320,In_15,In_996);
and U4321 (N_4321,In_545,In_222);
or U4322 (N_4322,In_371,In_821);
or U4323 (N_4323,In_451,In_406);
and U4324 (N_4324,In_741,In_208);
or U4325 (N_4325,In_115,In_287);
or U4326 (N_4326,In_590,In_797);
and U4327 (N_4327,In_15,In_20);
nand U4328 (N_4328,In_246,In_788);
nand U4329 (N_4329,In_593,In_774);
or U4330 (N_4330,In_215,In_536);
or U4331 (N_4331,In_72,In_987);
and U4332 (N_4332,In_427,In_275);
nor U4333 (N_4333,In_789,In_593);
nand U4334 (N_4334,In_378,In_314);
and U4335 (N_4335,In_713,In_986);
nor U4336 (N_4336,In_176,In_243);
nand U4337 (N_4337,In_459,In_136);
nand U4338 (N_4338,In_772,In_361);
nor U4339 (N_4339,In_386,In_55);
nor U4340 (N_4340,In_889,In_670);
nand U4341 (N_4341,In_778,In_109);
or U4342 (N_4342,In_960,In_315);
xnor U4343 (N_4343,In_883,In_555);
or U4344 (N_4344,In_895,In_257);
and U4345 (N_4345,In_506,In_778);
and U4346 (N_4346,In_982,In_344);
or U4347 (N_4347,In_246,In_596);
and U4348 (N_4348,In_837,In_416);
and U4349 (N_4349,In_929,In_446);
and U4350 (N_4350,In_511,In_235);
or U4351 (N_4351,In_23,In_562);
nor U4352 (N_4352,In_409,In_617);
nand U4353 (N_4353,In_859,In_688);
or U4354 (N_4354,In_535,In_388);
and U4355 (N_4355,In_705,In_159);
or U4356 (N_4356,In_402,In_265);
nor U4357 (N_4357,In_685,In_317);
nor U4358 (N_4358,In_903,In_78);
xor U4359 (N_4359,In_442,In_117);
or U4360 (N_4360,In_396,In_84);
and U4361 (N_4361,In_354,In_194);
or U4362 (N_4362,In_105,In_68);
nand U4363 (N_4363,In_325,In_417);
or U4364 (N_4364,In_543,In_62);
nor U4365 (N_4365,In_440,In_748);
nor U4366 (N_4366,In_459,In_520);
nand U4367 (N_4367,In_876,In_729);
and U4368 (N_4368,In_173,In_124);
and U4369 (N_4369,In_407,In_519);
xnor U4370 (N_4370,In_544,In_630);
and U4371 (N_4371,In_479,In_675);
nor U4372 (N_4372,In_336,In_230);
nor U4373 (N_4373,In_227,In_588);
nand U4374 (N_4374,In_873,In_48);
xor U4375 (N_4375,In_769,In_47);
nor U4376 (N_4376,In_642,In_845);
nand U4377 (N_4377,In_313,In_650);
xnor U4378 (N_4378,In_569,In_929);
and U4379 (N_4379,In_905,In_555);
nor U4380 (N_4380,In_455,In_286);
and U4381 (N_4381,In_151,In_300);
nand U4382 (N_4382,In_50,In_233);
or U4383 (N_4383,In_329,In_167);
or U4384 (N_4384,In_645,In_775);
and U4385 (N_4385,In_890,In_160);
or U4386 (N_4386,In_747,In_979);
or U4387 (N_4387,In_3,In_36);
or U4388 (N_4388,In_992,In_62);
or U4389 (N_4389,In_340,In_31);
xor U4390 (N_4390,In_770,In_875);
or U4391 (N_4391,In_548,In_623);
nand U4392 (N_4392,In_990,In_487);
nor U4393 (N_4393,In_147,In_20);
and U4394 (N_4394,In_365,In_910);
nor U4395 (N_4395,In_655,In_433);
and U4396 (N_4396,In_275,In_598);
or U4397 (N_4397,In_374,In_769);
and U4398 (N_4398,In_355,In_237);
or U4399 (N_4399,In_120,In_349);
nor U4400 (N_4400,In_485,In_75);
and U4401 (N_4401,In_902,In_606);
or U4402 (N_4402,In_433,In_993);
xnor U4403 (N_4403,In_782,In_445);
nand U4404 (N_4404,In_190,In_743);
nor U4405 (N_4405,In_114,In_955);
nor U4406 (N_4406,In_160,In_922);
and U4407 (N_4407,In_312,In_21);
and U4408 (N_4408,In_455,In_969);
and U4409 (N_4409,In_156,In_332);
nor U4410 (N_4410,In_52,In_278);
or U4411 (N_4411,In_817,In_778);
nand U4412 (N_4412,In_896,In_104);
nand U4413 (N_4413,In_667,In_414);
or U4414 (N_4414,In_75,In_512);
xnor U4415 (N_4415,In_443,In_728);
nor U4416 (N_4416,In_217,In_347);
or U4417 (N_4417,In_567,In_558);
nor U4418 (N_4418,In_825,In_8);
and U4419 (N_4419,In_194,In_724);
and U4420 (N_4420,In_471,In_545);
nand U4421 (N_4421,In_389,In_92);
nor U4422 (N_4422,In_291,In_154);
xor U4423 (N_4423,In_352,In_588);
nand U4424 (N_4424,In_299,In_549);
xor U4425 (N_4425,In_618,In_228);
nor U4426 (N_4426,In_142,In_252);
nor U4427 (N_4427,In_331,In_176);
nor U4428 (N_4428,In_989,In_196);
xnor U4429 (N_4429,In_877,In_161);
and U4430 (N_4430,In_466,In_74);
nand U4431 (N_4431,In_255,In_560);
or U4432 (N_4432,In_847,In_760);
and U4433 (N_4433,In_20,In_704);
nand U4434 (N_4434,In_430,In_135);
nand U4435 (N_4435,In_811,In_366);
nor U4436 (N_4436,In_956,In_276);
and U4437 (N_4437,In_274,In_698);
nor U4438 (N_4438,In_453,In_552);
nand U4439 (N_4439,In_232,In_642);
xnor U4440 (N_4440,In_380,In_855);
and U4441 (N_4441,In_117,In_320);
and U4442 (N_4442,In_841,In_544);
nand U4443 (N_4443,In_282,In_373);
or U4444 (N_4444,In_186,In_653);
nand U4445 (N_4445,In_229,In_456);
nor U4446 (N_4446,In_160,In_202);
nand U4447 (N_4447,In_819,In_968);
nor U4448 (N_4448,In_899,In_377);
and U4449 (N_4449,In_190,In_124);
nand U4450 (N_4450,In_42,In_345);
nor U4451 (N_4451,In_924,In_46);
xor U4452 (N_4452,In_156,In_210);
nor U4453 (N_4453,In_718,In_571);
or U4454 (N_4454,In_20,In_542);
and U4455 (N_4455,In_275,In_124);
nand U4456 (N_4456,In_772,In_497);
nor U4457 (N_4457,In_717,In_852);
and U4458 (N_4458,In_777,In_773);
and U4459 (N_4459,In_531,In_512);
xnor U4460 (N_4460,In_162,In_186);
nand U4461 (N_4461,In_548,In_62);
nor U4462 (N_4462,In_203,In_21);
and U4463 (N_4463,In_525,In_580);
or U4464 (N_4464,In_326,In_318);
nand U4465 (N_4465,In_24,In_883);
nor U4466 (N_4466,In_415,In_473);
and U4467 (N_4467,In_987,In_332);
nand U4468 (N_4468,In_37,In_82);
or U4469 (N_4469,In_697,In_940);
nand U4470 (N_4470,In_530,In_982);
nand U4471 (N_4471,In_848,In_181);
nand U4472 (N_4472,In_245,In_692);
nand U4473 (N_4473,In_35,In_80);
and U4474 (N_4474,In_70,In_532);
xor U4475 (N_4475,In_63,In_380);
nor U4476 (N_4476,In_917,In_65);
or U4477 (N_4477,In_994,In_605);
xnor U4478 (N_4478,In_119,In_338);
and U4479 (N_4479,In_530,In_467);
and U4480 (N_4480,In_595,In_874);
or U4481 (N_4481,In_161,In_543);
nand U4482 (N_4482,In_990,In_229);
and U4483 (N_4483,In_157,In_533);
or U4484 (N_4484,In_680,In_125);
nand U4485 (N_4485,In_177,In_11);
nand U4486 (N_4486,In_253,In_104);
or U4487 (N_4487,In_987,In_740);
and U4488 (N_4488,In_566,In_256);
nor U4489 (N_4489,In_769,In_461);
or U4490 (N_4490,In_103,In_810);
xor U4491 (N_4491,In_265,In_53);
nand U4492 (N_4492,In_166,In_766);
nor U4493 (N_4493,In_348,In_701);
nand U4494 (N_4494,In_446,In_794);
and U4495 (N_4495,In_799,In_725);
nor U4496 (N_4496,In_39,In_435);
nand U4497 (N_4497,In_227,In_284);
and U4498 (N_4498,In_128,In_788);
nand U4499 (N_4499,In_228,In_407);
nor U4500 (N_4500,In_47,In_844);
nor U4501 (N_4501,In_86,In_920);
nand U4502 (N_4502,In_489,In_535);
and U4503 (N_4503,In_505,In_943);
and U4504 (N_4504,In_11,In_686);
and U4505 (N_4505,In_891,In_878);
nor U4506 (N_4506,In_801,In_29);
or U4507 (N_4507,In_530,In_738);
nand U4508 (N_4508,In_883,In_678);
and U4509 (N_4509,In_638,In_993);
or U4510 (N_4510,In_625,In_834);
and U4511 (N_4511,In_238,In_387);
nand U4512 (N_4512,In_747,In_945);
nor U4513 (N_4513,In_306,In_396);
xor U4514 (N_4514,In_105,In_904);
xnor U4515 (N_4515,In_846,In_145);
or U4516 (N_4516,In_105,In_152);
or U4517 (N_4517,In_112,In_197);
or U4518 (N_4518,In_22,In_476);
nand U4519 (N_4519,In_424,In_896);
nor U4520 (N_4520,In_504,In_953);
or U4521 (N_4521,In_107,In_453);
and U4522 (N_4522,In_489,In_222);
or U4523 (N_4523,In_401,In_904);
and U4524 (N_4524,In_62,In_809);
and U4525 (N_4525,In_540,In_270);
nor U4526 (N_4526,In_237,In_745);
and U4527 (N_4527,In_103,In_416);
or U4528 (N_4528,In_69,In_703);
or U4529 (N_4529,In_471,In_76);
or U4530 (N_4530,In_700,In_15);
nor U4531 (N_4531,In_207,In_739);
nand U4532 (N_4532,In_899,In_472);
nor U4533 (N_4533,In_323,In_804);
or U4534 (N_4534,In_824,In_436);
or U4535 (N_4535,In_479,In_88);
or U4536 (N_4536,In_179,In_162);
or U4537 (N_4537,In_21,In_509);
xnor U4538 (N_4538,In_761,In_406);
nand U4539 (N_4539,In_535,In_645);
and U4540 (N_4540,In_232,In_990);
or U4541 (N_4541,In_781,In_742);
and U4542 (N_4542,In_68,In_997);
or U4543 (N_4543,In_997,In_854);
or U4544 (N_4544,In_331,In_721);
xor U4545 (N_4545,In_265,In_633);
xor U4546 (N_4546,In_921,In_668);
nand U4547 (N_4547,In_286,In_536);
and U4548 (N_4548,In_860,In_915);
and U4549 (N_4549,In_566,In_543);
nand U4550 (N_4550,In_108,In_597);
nand U4551 (N_4551,In_457,In_55);
or U4552 (N_4552,In_434,In_259);
nand U4553 (N_4553,In_844,In_704);
and U4554 (N_4554,In_729,In_73);
nand U4555 (N_4555,In_870,In_782);
nand U4556 (N_4556,In_145,In_454);
and U4557 (N_4557,In_598,In_651);
nand U4558 (N_4558,In_943,In_794);
nand U4559 (N_4559,In_278,In_741);
xor U4560 (N_4560,In_349,In_208);
or U4561 (N_4561,In_303,In_808);
nor U4562 (N_4562,In_469,In_964);
and U4563 (N_4563,In_318,In_955);
nand U4564 (N_4564,In_297,In_502);
xor U4565 (N_4565,In_742,In_359);
and U4566 (N_4566,In_141,In_143);
nor U4567 (N_4567,In_972,In_164);
and U4568 (N_4568,In_518,In_620);
nor U4569 (N_4569,In_279,In_419);
nand U4570 (N_4570,In_779,In_48);
nand U4571 (N_4571,In_508,In_901);
nand U4572 (N_4572,In_301,In_84);
nor U4573 (N_4573,In_216,In_692);
and U4574 (N_4574,In_938,In_789);
xnor U4575 (N_4575,In_69,In_432);
nor U4576 (N_4576,In_719,In_968);
or U4577 (N_4577,In_273,In_914);
nor U4578 (N_4578,In_721,In_620);
nand U4579 (N_4579,In_849,In_750);
nor U4580 (N_4580,In_44,In_685);
and U4581 (N_4581,In_922,In_680);
or U4582 (N_4582,In_423,In_67);
nand U4583 (N_4583,In_609,In_877);
or U4584 (N_4584,In_185,In_683);
nand U4585 (N_4585,In_52,In_609);
and U4586 (N_4586,In_15,In_300);
and U4587 (N_4587,In_795,In_749);
nand U4588 (N_4588,In_898,In_224);
or U4589 (N_4589,In_931,In_806);
nand U4590 (N_4590,In_108,In_258);
or U4591 (N_4591,In_551,In_356);
and U4592 (N_4592,In_258,In_522);
or U4593 (N_4593,In_328,In_667);
xor U4594 (N_4594,In_674,In_381);
or U4595 (N_4595,In_632,In_323);
nor U4596 (N_4596,In_993,In_352);
nand U4597 (N_4597,In_601,In_433);
nand U4598 (N_4598,In_535,In_316);
and U4599 (N_4599,In_158,In_863);
nor U4600 (N_4600,In_915,In_675);
nand U4601 (N_4601,In_16,In_866);
and U4602 (N_4602,In_734,In_864);
xor U4603 (N_4603,In_884,In_567);
xnor U4604 (N_4604,In_74,In_238);
nor U4605 (N_4605,In_434,In_168);
and U4606 (N_4606,In_750,In_526);
nand U4607 (N_4607,In_894,In_799);
or U4608 (N_4608,In_413,In_881);
and U4609 (N_4609,In_823,In_496);
or U4610 (N_4610,In_735,In_774);
nand U4611 (N_4611,In_872,In_774);
nor U4612 (N_4612,In_111,In_763);
nand U4613 (N_4613,In_595,In_781);
nand U4614 (N_4614,In_542,In_992);
nand U4615 (N_4615,In_157,In_249);
or U4616 (N_4616,In_734,In_28);
nor U4617 (N_4617,In_372,In_742);
and U4618 (N_4618,In_880,In_353);
nor U4619 (N_4619,In_47,In_226);
xnor U4620 (N_4620,In_718,In_616);
and U4621 (N_4621,In_671,In_643);
xor U4622 (N_4622,In_873,In_337);
or U4623 (N_4623,In_833,In_815);
or U4624 (N_4624,In_922,In_974);
nand U4625 (N_4625,In_282,In_173);
nor U4626 (N_4626,In_1,In_986);
or U4627 (N_4627,In_842,In_62);
nand U4628 (N_4628,In_655,In_71);
or U4629 (N_4629,In_646,In_994);
or U4630 (N_4630,In_461,In_372);
nand U4631 (N_4631,In_967,In_417);
or U4632 (N_4632,In_300,In_905);
or U4633 (N_4633,In_532,In_938);
or U4634 (N_4634,In_491,In_762);
and U4635 (N_4635,In_611,In_465);
xor U4636 (N_4636,In_338,In_747);
nor U4637 (N_4637,In_933,In_770);
nor U4638 (N_4638,In_643,In_757);
and U4639 (N_4639,In_95,In_846);
or U4640 (N_4640,In_648,In_947);
nand U4641 (N_4641,In_983,In_805);
xnor U4642 (N_4642,In_268,In_319);
xor U4643 (N_4643,In_694,In_142);
and U4644 (N_4644,In_320,In_682);
nor U4645 (N_4645,In_540,In_669);
or U4646 (N_4646,In_649,In_756);
xnor U4647 (N_4647,In_454,In_757);
and U4648 (N_4648,In_693,In_234);
or U4649 (N_4649,In_913,In_32);
nor U4650 (N_4650,In_961,In_846);
and U4651 (N_4651,In_731,In_436);
and U4652 (N_4652,In_656,In_78);
nor U4653 (N_4653,In_347,In_164);
nand U4654 (N_4654,In_977,In_134);
nand U4655 (N_4655,In_941,In_280);
nand U4656 (N_4656,In_28,In_318);
xor U4657 (N_4657,In_58,In_29);
nor U4658 (N_4658,In_988,In_857);
xor U4659 (N_4659,In_705,In_908);
or U4660 (N_4660,In_749,In_720);
nor U4661 (N_4661,In_158,In_910);
nand U4662 (N_4662,In_108,In_447);
and U4663 (N_4663,In_969,In_862);
xor U4664 (N_4664,In_746,In_760);
nor U4665 (N_4665,In_874,In_921);
nor U4666 (N_4666,In_811,In_731);
or U4667 (N_4667,In_365,In_41);
and U4668 (N_4668,In_230,In_551);
xnor U4669 (N_4669,In_518,In_191);
or U4670 (N_4670,In_495,In_474);
nand U4671 (N_4671,In_149,In_860);
nand U4672 (N_4672,In_524,In_89);
nor U4673 (N_4673,In_915,In_684);
nand U4674 (N_4674,In_475,In_772);
nand U4675 (N_4675,In_578,In_667);
nor U4676 (N_4676,In_752,In_317);
nor U4677 (N_4677,In_599,In_817);
or U4678 (N_4678,In_779,In_291);
nor U4679 (N_4679,In_172,In_541);
xor U4680 (N_4680,In_502,In_343);
nand U4681 (N_4681,In_731,In_340);
nand U4682 (N_4682,In_55,In_190);
nor U4683 (N_4683,In_444,In_194);
and U4684 (N_4684,In_837,In_504);
nand U4685 (N_4685,In_546,In_407);
and U4686 (N_4686,In_223,In_919);
nand U4687 (N_4687,In_428,In_653);
and U4688 (N_4688,In_815,In_722);
xnor U4689 (N_4689,In_738,In_425);
nor U4690 (N_4690,In_277,In_658);
and U4691 (N_4691,In_891,In_805);
xor U4692 (N_4692,In_288,In_845);
nand U4693 (N_4693,In_537,In_301);
xor U4694 (N_4694,In_417,In_389);
nand U4695 (N_4695,In_783,In_19);
nand U4696 (N_4696,In_27,In_872);
and U4697 (N_4697,In_308,In_633);
or U4698 (N_4698,In_786,In_624);
and U4699 (N_4699,In_680,In_386);
and U4700 (N_4700,In_631,In_137);
nor U4701 (N_4701,In_517,In_477);
nor U4702 (N_4702,In_669,In_483);
or U4703 (N_4703,In_916,In_223);
nand U4704 (N_4704,In_418,In_526);
or U4705 (N_4705,In_535,In_949);
and U4706 (N_4706,In_215,In_396);
nand U4707 (N_4707,In_439,In_503);
nand U4708 (N_4708,In_106,In_509);
xnor U4709 (N_4709,In_111,In_835);
nor U4710 (N_4710,In_795,In_933);
nor U4711 (N_4711,In_675,In_839);
nand U4712 (N_4712,In_571,In_616);
xor U4713 (N_4713,In_914,In_826);
or U4714 (N_4714,In_313,In_450);
or U4715 (N_4715,In_972,In_557);
or U4716 (N_4716,In_167,In_654);
and U4717 (N_4717,In_832,In_224);
and U4718 (N_4718,In_2,In_850);
nand U4719 (N_4719,In_216,In_465);
and U4720 (N_4720,In_926,In_45);
nor U4721 (N_4721,In_465,In_111);
or U4722 (N_4722,In_925,In_127);
nand U4723 (N_4723,In_792,In_905);
nor U4724 (N_4724,In_484,In_200);
or U4725 (N_4725,In_54,In_835);
or U4726 (N_4726,In_281,In_948);
or U4727 (N_4727,In_739,In_940);
or U4728 (N_4728,In_319,In_968);
xor U4729 (N_4729,In_102,In_659);
or U4730 (N_4730,In_480,In_729);
or U4731 (N_4731,In_76,In_458);
or U4732 (N_4732,In_728,In_742);
and U4733 (N_4733,In_397,In_318);
xor U4734 (N_4734,In_7,In_900);
nand U4735 (N_4735,In_304,In_416);
and U4736 (N_4736,In_584,In_402);
nor U4737 (N_4737,In_360,In_930);
nand U4738 (N_4738,In_68,In_849);
nor U4739 (N_4739,In_40,In_77);
and U4740 (N_4740,In_440,In_586);
nor U4741 (N_4741,In_299,In_641);
and U4742 (N_4742,In_252,In_416);
nor U4743 (N_4743,In_154,In_912);
nor U4744 (N_4744,In_849,In_393);
or U4745 (N_4745,In_813,In_885);
and U4746 (N_4746,In_101,In_627);
and U4747 (N_4747,In_925,In_991);
or U4748 (N_4748,In_231,In_845);
nor U4749 (N_4749,In_933,In_200);
xnor U4750 (N_4750,In_256,In_290);
or U4751 (N_4751,In_708,In_386);
and U4752 (N_4752,In_233,In_888);
or U4753 (N_4753,In_935,In_489);
and U4754 (N_4754,In_159,In_15);
and U4755 (N_4755,In_896,In_50);
nor U4756 (N_4756,In_326,In_576);
and U4757 (N_4757,In_242,In_210);
nand U4758 (N_4758,In_286,In_105);
nand U4759 (N_4759,In_928,In_729);
xor U4760 (N_4760,In_572,In_891);
nor U4761 (N_4761,In_170,In_446);
and U4762 (N_4762,In_44,In_970);
and U4763 (N_4763,In_966,In_103);
nand U4764 (N_4764,In_66,In_798);
xnor U4765 (N_4765,In_653,In_534);
nor U4766 (N_4766,In_76,In_943);
and U4767 (N_4767,In_636,In_436);
or U4768 (N_4768,In_861,In_862);
nand U4769 (N_4769,In_798,In_614);
nand U4770 (N_4770,In_313,In_881);
and U4771 (N_4771,In_835,In_375);
nor U4772 (N_4772,In_504,In_608);
nor U4773 (N_4773,In_697,In_764);
nand U4774 (N_4774,In_519,In_796);
and U4775 (N_4775,In_958,In_853);
and U4776 (N_4776,In_53,In_230);
nor U4777 (N_4777,In_946,In_142);
nand U4778 (N_4778,In_250,In_98);
or U4779 (N_4779,In_673,In_779);
or U4780 (N_4780,In_329,In_28);
or U4781 (N_4781,In_771,In_275);
nand U4782 (N_4782,In_993,In_270);
nor U4783 (N_4783,In_579,In_453);
xnor U4784 (N_4784,In_871,In_788);
and U4785 (N_4785,In_490,In_168);
or U4786 (N_4786,In_224,In_488);
nand U4787 (N_4787,In_729,In_492);
nor U4788 (N_4788,In_787,In_880);
nand U4789 (N_4789,In_863,In_208);
or U4790 (N_4790,In_137,In_772);
or U4791 (N_4791,In_739,In_750);
nand U4792 (N_4792,In_454,In_167);
or U4793 (N_4793,In_198,In_983);
and U4794 (N_4794,In_916,In_794);
xnor U4795 (N_4795,In_79,In_309);
nor U4796 (N_4796,In_141,In_452);
nor U4797 (N_4797,In_84,In_58);
or U4798 (N_4798,In_935,In_551);
and U4799 (N_4799,In_322,In_566);
or U4800 (N_4800,In_752,In_479);
or U4801 (N_4801,In_932,In_26);
and U4802 (N_4802,In_492,In_548);
or U4803 (N_4803,In_87,In_757);
and U4804 (N_4804,In_694,In_354);
or U4805 (N_4805,In_520,In_608);
nor U4806 (N_4806,In_378,In_156);
nand U4807 (N_4807,In_72,In_771);
or U4808 (N_4808,In_300,In_288);
nand U4809 (N_4809,In_917,In_61);
nand U4810 (N_4810,In_818,In_188);
nand U4811 (N_4811,In_179,In_551);
nor U4812 (N_4812,In_253,In_82);
or U4813 (N_4813,In_519,In_363);
or U4814 (N_4814,In_518,In_771);
nor U4815 (N_4815,In_357,In_813);
nor U4816 (N_4816,In_934,In_582);
nand U4817 (N_4817,In_157,In_857);
and U4818 (N_4818,In_932,In_782);
or U4819 (N_4819,In_641,In_444);
xor U4820 (N_4820,In_468,In_651);
nand U4821 (N_4821,In_504,In_65);
nand U4822 (N_4822,In_396,In_750);
nand U4823 (N_4823,In_497,In_444);
nor U4824 (N_4824,In_329,In_51);
nand U4825 (N_4825,In_355,In_441);
nor U4826 (N_4826,In_312,In_2);
or U4827 (N_4827,In_836,In_793);
nand U4828 (N_4828,In_768,In_669);
xnor U4829 (N_4829,In_831,In_515);
nor U4830 (N_4830,In_900,In_280);
and U4831 (N_4831,In_438,In_636);
nor U4832 (N_4832,In_265,In_983);
nand U4833 (N_4833,In_944,In_130);
nor U4834 (N_4834,In_208,In_701);
or U4835 (N_4835,In_392,In_103);
and U4836 (N_4836,In_788,In_706);
nor U4837 (N_4837,In_720,In_564);
nor U4838 (N_4838,In_298,In_373);
and U4839 (N_4839,In_110,In_97);
nor U4840 (N_4840,In_438,In_483);
or U4841 (N_4841,In_33,In_158);
or U4842 (N_4842,In_436,In_689);
nor U4843 (N_4843,In_783,In_551);
nor U4844 (N_4844,In_770,In_420);
nor U4845 (N_4845,In_861,In_683);
nand U4846 (N_4846,In_91,In_541);
and U4847 (N_4847,In_298,In_188);
nor U4848 (N_4848,In_486,In_780);
nor U4849 (N_4849,In_837,In_545);
xor U4850 (N_4850,In_532,In_870);
and U4851 (N_4851,In_677,In_724);
nor U4852 (N_4852,In_962,In_115);
nor U4853 (N_4853,In_778,In_432);
or U4854 (N_4854,In_818,In_868);
xor U4855 (N_4855,In_150,In_567);
nor U4856 (N_4856,In_231,In_559);
and U4857 (N_4857,In_835,In_198);
and U4858 (N_4858,In_660,In_799);
nor U4859 (N_4859,In_107,In_576);
and U4860 (N_4860,In_729,In_749);
or U4861 (N_4861,In_93,In_719);
nand U4862 (N_4862,In_575,In_716);
nor U4863 (N_4863,In_59,In_774);
and U4864 (N_4864,In_971,In_69);
nand U4865 (N_4865,In_4,In_598);
nor U4866 (N_4866,In_220,In_363);
nand U4867 (N_4867,In_649,In_561);
and U4868 (N_4868,In_71,In_180);
nand U4869 (N_4869,In_530,In_863);
and U4870 (N_4870,In_117,In_384);
nand U4871 (N_4871,In_498,In_374);
or U4872 (N_4872,In_40,In_869);
and U4873 (N_4873,In_130,In_312);
nor U4874 (N_4874,In_465,In_871);
nand U4875 (N_4875,In_796,In_543);
nand U4876 (N_4876,In_339,In_847);
or U4877 (N_4877,In_991,In_338);
nor U4878 (N_4878,In_699,In_363);
nor U4879 (N_4879,In_387,In_598);
and U4880 (N_4880,In_208,In_890);
and U4881 (N_4881,In_781,In_888);
nor U4882 (N_4882,In_863,In_312);
and U4883 (N_4883,In_683,In_524);
nor U4884 (N_4884,In_475,In_648);
xor U4885 (N_4885,In_246,In_107);
and U4886 (N_4886,In_960,In_299);
nand U4887 (N_4887,In_594,In_939);
xnor U4888 (N_4888,In_144,In_757);
or U4889 (N_4889,In_379,In_500);
nor U4890 (N_4890,In_885,In_490);
xor U4891 (N_4891,In_57,In_548);
and U4892 (N_4892,In_883,In_794);
xnor U4893 (N_4893,In_809,In_247);
and U4894 (N_4894,In_456,In_408);
and U4895 (N_4895,In_565,In_316);
nand U4896 (N_4896,In_309,In_997);
or U4897 (N_4897,In_537,In_283);
or U4898 (N_4898,In_400,In_593);
and U4899 (N_4899,In_22,In_199);
nand U4900 (N_4900,In_156,In_417);
and U4901 (N_4901,In_892,In_528);
or U4902 (N_4902,In_161,In_723);
and U4903 (N_4903,In_956,In_82);
and U4904 (N_4904,In_801,In_255);
or U4905 (N_4905,In_392,In_49);
nor U4906 (N_4906,In_697,In_840);
and U4907 (N_4907,In_135,In_795);
nand U4908 (N_4908,In_447,In_811);
and U4909 (N_4909,In_741,In_204);
and U4910 (N_4910,In_227,In_430);
xnor U4911 (N_4911,In_181,In_568);
nand U4912 (N_4912,In_84,In_363);
or U4913 (N_4913,In_537,In_663);
or U4914 (N_4914,In_717,In_383);
nor U4915 (N_4915,In_204,In_328);
or U4916 (N_4916,In_808,In_109);
nor U4917 (N_4917,In_300,In_61);
or U4918 (N_4918,In_746,In_94);
nor U4919 (N_4919,In_285,In_960);
and U4920 (N_4920,In_106,In_223);
nor U4921 (N_4921,In_868,In_250);
and U4922 (N_4922,In_821,In_243);
or U4923 (N_4923,In_609,In_540);
nor U4924 (N_4924,In_540,In_949);
nand U4925 (N_4925,In_112,In_609);
and U4926 (N_4926,In_814,In_257);
nor U4927 (N_4927,In_164,In_803);
nand U4928 (N_4928,In_4,In_153);
nand U4929 (N_4929,In_527,In_986);
nor U4930 (N_4930,In_992,In_933);
and U4931 (N_4931,In_478,In_266);
nor U4932 (N_4932,In_903,In_808);
or U4933 (N_4933,In_442,In_548);
nand U4934 (N_4934,In_485,In_867);
or U4935 (N_4935,In_159,In_251);
nor U4936 (N_4936,In_467,In_277);
nor U4937 (N_4937,In_0,In_747);
and U4938 (N_4938,In_26,In_644);
nand U4939 (N_4939,In_581,In_65);
or U4940 (N_4940,In_715,In_240);
and U4941 (N_4941,In_129,In_235);
nand U4942 (N_4942,In_910,In_732);
and U4943 (N_4943,In_249,In_766);
or U4944 (N_4944,In_516,In_60);
or U4945 (N_4945,In_772,In_172);
and U4946 (N_4946,In_474,In_217);
nand U4947 (N_4947,In_33,In_719);
and U4948 (N_4948,In_189,In_577);
and U4949 (N_4949,In_186,In_518);
nor U4950 (N_4950,In_736,In_23);
nor U4951 (N_4951,In_155,In_128);
nand U4952 (N_4952,In_444,In_368);
nor U4953 (N_4953,In_408,In_876);
xnor U4954 (N_4954,In_299,In_554);
nor U4955 (N_4955,In_376,In_409);
nor U4956 (N_4956,In_751,In_151);
nand U4957 (N_4957,In_998,In_148);
or U4958 (N_4958,In_135,In_349);
nand U4959 (N_4959,In_766,In_721);
or U4960 (N_4960,In_471,In_688);
or U4961 (N_4961,In_195,In_176);
nand U4962 (N_4962,In_38,In_131);
and U4963 (N_4963,In_31,In_934);
nor U4964 (N_4964,In_574,In_443);
or U4965 (N_4965,In_377,In_177);
nor U4966 (N_4966,In_292,In_349);
nand U4967 (N_4967,In_437,In_496);
nand U4968 (N_4968,In_322,In_297);
xnor U4969 (N_4969,In_845,In_358);
nand U4970 (N_4970,In_389,In_665);
nand U4971 (N_4971,In_730,In_431);
or U4972 (N_4972,In_249,In_578);
nand U4973 (N_4973,In_620,In_165);
xnor U4974 (N_4974,In_759,In_384);
nor U4975 (N_4975,In_471,In_825);
and U4976 (N_4976,In_772,In_762);
and U4977 (N_4977,In_702,In_981);
or U4978 (N_4978,In_602,In_383);
nor U4979 (N_4979,In_444,In_710);
xnor U4980 (N_4980,In_898,In_97);
nand U4981 (N_4981,In_568,In_366);
nand U4982 (N_4982,In_920,In_466);
xnor U4983 (N_4983,In_550,In_623);
nand U4984 (N_4984,In_270,In_823);
xor U4985 (N_4985,In_104,In_93);
nand U4986 (N_4986,In_161,In_339);
nor U4987 (N_4987,In_507,In_863);
or U4988 (N_4988,In_818,In_393);
or U4989 (N_4989,In_77,In_104);
and U4990 (N_4990,In_654,In_498);
and U4991 (N_4991,In_489,In_753);
nor U4992 (N_4992,In_537,In_718);
xor U4993 (N_4993,In_414,In_479);
nor U4994 (N_4994,In_86,In_523);
and U4995 (N_4995,In_758,In_743);
nor U4996 (N_4996,In_588,In_670);
nor U4997 (N_4997,In_201,In_803);
nor U4998 (N_4998,In_365,In_374);
nor U4999 (N_4999,In_356,In_842);
and U5000 (N_5000,N_20,N_1109);
nand U5001 (N_5001,N_4857,N_2651);
xor U5002 (N_5002,N_557,N_2285);
nor U5003 (N_5003,N_3759,N_3395);
and U5004 (N_5004,N_875,N_4202);
nand U5005 (N_5005,N_3958,N_191);
xor U5006 (N_5006,N_3504,N_3540);
nand U5007 (N_5007,N_4988,N_4523);
and U5008 (N_5008,N_3358,N_1878);
nand U5009 (N_5009,N_1500,N_2238);
nor U5010 (N_5010,N_4760,N_1208);
and U5011 (N_5011,N_989,N_2184);
nand U5012 (N_5012,N_3848,N_1005);
or U5013 (N_5013,N_1909,N_828);
nor U5014 (N_5014,N_1711,N_4963);
or U5015 (N_5015,N_4500,N_1624);
and U5016 (N_5016,N_4862,N_1563);
nor U5017 (N_5017,N_4582,N_2542);
nor U5018 (N_5018,N_838,N_592);
nor U5019 (N_5019,N_2514,N_2933);
nor U5020 (N_5020,N_4553,N_220);
or U5021 (N_5021,N_1873,N_3565);
and U5022 (N_5022,N_3310,N_2856);
or U5023 (N_5023,N_744,N_4761);
and U5024 (N_5024,N_2773,N_387);
nor U5025 (N_5025,N_4890,N_2469);
xor U5026 (N_5026,N_4133,N_1185);
nor U5027 (N_5027,N_4797,N_1453);
nand U5028 (N_5028,N_4660,N_4);
or U5029 (N_5029,N_3263,N_4893);
and U5030 (N_5030,N_1324,N_1600);
and U5031 (N_5031,N_4437,N_139);
nand U5032 (N_5032,N_3538,N_621);
and U5033 (N_5033,N_1629,N_1896);
or U5034 (N_5034,N_885,N_2154);
nor U5035 (N_5035,N_1206,N_4615);
or U5036 (N_5036,N_3706,N_2897);
nor U5037 (N_5037,N_1780,N_4846);
nor U5038 (N_5038,N_4006,N_2090);
xor U5039 (N_5039,N_553,N_3340);
xor U5040 (N_5040,N_4560,N_1698);
or U5041 (N_5041,N_1008,N_1728);
nor U5042 (N_5042,N_115,N_3393);
or U5043 (N_5043,N_2286,N_27);
and U5044 (N_5044,N_2440,N_1228);
or U5045 (N_5045,N_3619,N_2415);
nand U5046 (N_5046,N_4197,N_3626);
nor U5047 (N_5047,N_4678,N_4685);
nor U5048 (N_5048,N_2637,N_822);
and U5049 (N_5049,N_2189,N_4337);
nand U5050 (N_5050,N_3284,N_4892);
xor U5051 (N_5051,N_2211,N_510);
xnor U5052 (N_5052,N_4896,N_2853);
xnor U5053 (N_5053,N_231,N_4220);
nor U5054 (N_5054,N_3857,N_4096);
xor U5055 (N_5055,N_2413,N_2341);
and U5056 (N_5056,N_1571,N_455);
or U5057 (N_5057,N_3063,N_3029);
nor U5058 (N_5058,N_2338,N_3233);
or U5059 (N_5059,N_1236,N_692);
or U5060 (N_5060,N_4820,N_718);
nor U5061 (N_5061,N_371,N_771);
nand U5062 (N_5062,N_476,N_3246);
or U5063 (N_5063,N_4454,N_4294);
nand U5064 (N_5064,N_1884,N_1916);
nand U5065 (N_5065,N_4422,N_3144);
xnor U5066 (N_5066,N_799,N_4719);
or U5067 (N_5067,N_4885,N_1582);
nand U5068 (N_5068,N_1486,N_2546);
nor U5069 (N_5069,N_4526,N_4246);
nor U5070 (N_5070,N_1238,N_1601);
or U5071 (N_5071,N_925,N_3396);
nand U5072 (N_5072,N_2385,N_205);
xnor U5073 (N_5073,N_1432,N_3131);
xor U5074 (N_5074,N_4874,N_2234);
nand U5075 (N_5075,N_159,N_541);
and U5076 (N_5076,N_1815,N_2598);
or U5077 (N_5077,N_2509,N_1576);
nand U5078 (N_5078,N_2359,N_2859);
and U5079 (N_5079,N_1021,N_289);
nand U5080 (N_5080,N_4871,N_4101);
nand U5081 (N_5081,N_1555,N_1076);
nor U5082 (N_5082,N_4625,N_1213);
and U5083 (N_5083,N_3556,N_1050);
or U5084 (N_5084,N_4591,N_1508);
or U5085 (N_5085,N_3946,N_3579);
or U5086 (N_5086,N_279,N_4020);
nor U5087 (N_5087,N_1464,N_2122);
and U5088 (N_5088,N_1424,N_2851);
nor U5089 (N_5089,N_3043,N_1932);
xnor U5090 (N_5090,N_851,N_4858);
and U5091 (N_5091,N_4714,N_3594);
or U5092 (N_5092,N_2436,N_315);
or U5093 (N_5093,N_1748,N_4470);
nand U5094 (N_5094,N_207,N_4784);
or U5095 (N_5095,N_4914,N_4711);
nor U5096 (N_5096,N_3306,N_3321);
nor U5097 (N_5097,N_3792,N_1811);
nand U5098 (N_5098,N_4190,N_3980);
xor U5099 (N_5099,N_853,N_2091);
or U5100 (N_5100,N_3894,N_4795);
nand U5101 (N_5101,N_1348,N_9);
nand U5102 (N_5102,N_2582,N_1176);
nand U5103 (N_5103,N_1712,N_4045);
nand U5104 (N_5104,N_3803,N_3229);
nand U5105 (N_5105,N_1817,N_3106);
nand U5106 (N_5106,N_2621,N_1144);
and U5107 (N_5107,N_2929,N_767);
and U5108 (N_5108,N_3884,N_1983);
or U5109 (N_5109,N_3937,N_1247);
xor U5110 (N_5110,N_2317,N_4116);
or U5111 (N_5111,N_2610,N_2980);
or U5112 (N_5112,N_2841,N_1919);
nand U5113 (N_5113,N_3702,N_4441);
xnor U5114 (N_5114,N_2024,N_993);
or U5115 (N_5115,N_3788,N_3075);
and U5116 (N_5116,N_2903,N_697);
xor U5117 (N_5117,N_43,N_2734);
or U5118 (N_5118,N_1099,N_4524);
and U5119 (N_5119,N_34,N_3123);
nand U5120 (N_5120,N_731,N_3282);
and U5121 (N_5121,N_3648,N_2443);
xor U5122 (N_5122,N_3835,N_1357);
nand U5123 (N_5123,N_129,N_3241);
nand U5124 (N_5124,N_2923,N_3247);
and U5125 (N_5125,N_4731,N_1141);
nor U5126 (N_5126,N_3189,N_317);
or U5127 (N_5127,N_4284,N_1869);
or U5128 (N_5128,N_2603,N_1297);
nor U5129 (N_5129,N_458,N_492);
nor U5130 (N_5130,N_4600,N_1781);
or U5131 (N_5131,N_1730,N_4255);
and U5132 (N_5132,N_1598,N_66);
and U5133 (N_5133,N_2937,N_2043);
or U5134 (N_5134,N_4200,N_4161);
nand U5135 (N_5135,N_1446,N_4712);
or U5136 (N_5136,N_609,N_1386);
nor U5137 (N_5137,N_1652,N_3056);
and U5138 (N_5138,N_1110,N_2074);
and U5139 (N_5139,N_942,N_1742);
nand U5140 (N_5140,N_4499,N_477);
and U5141 (N_5141,N_947,N_740);
nor U5142 (N_5142,N_3447,N_2535);
or U5143 (N_5143,N_1310,N_1737);
or U5144 (N_5144,N_2494,N_201);
nand U5145 (N_5145,N_1830,N_1749);
xor U5146 (N_5146,N_2505,N_4473);
or U5147 (N_5147,N_3492,N_446);
nor U5148 (N_5148,N_2308,N_359);
and U5149 (N_5149,N_486,N_2206);
and U5150 (N_5150,N_880,N_3858);
or U5151 (N_5151,N_4413,N_4387);
or U5152 (N_5152,N_3372,N_2792);
nor U5153 (N_5153,N_11,N_1644);
xnor U5154 (N_5154,N_4392,N_61);
nor U5155 (N_5155,N_4996,N_2177);
and U5156 (N_5156,N_3335,N_4718);
or U5157 (N_5157,N_1540,N_399);
and U5158 (N_5158,N_3834,N_4429);
and U5159 (N_5159,N_1963,N_1788);
nand U5160 (N_5160,N_2462,N_223);
and U5161 (N_5161,N_3789,N_3181);
or U5162 (N_5162,N_779,N_3547);
and U5163 (N_5163,N_271,N_1530);
or U5164 (N_5164,N_1263,N_2783);
xor U5165 (N_5165,N_4703,N_1999);
or U5166 (N_5166,N_1783,N_1);
nor U5167 (N_5167,N_2791,N_2798);
nand U5168 (N_5168,N_3260,N_3208);
nor U5169 (N_5169,N_3728,N_4014);
and U5170 (N_5170,N_1189,N_3672);
and U5171 (N_5171,N_1603,N_4036);
nand U5172 (N_5172,N_2070,N_2650);
or U5173 (N_5173,N_2021,N_4142);
and U5174 (N_5174,N_3090,N_1077);
nand U5175 (N_5175,N_530,N_4292);
xor U5176 (N_5176,N_1244,N_3201);
or U5177 (N_5177,N_631,N_2455);
and U5178 (N_5178,N_1370,N_257);
and U5179 (N_5179,N_2155,N_2183);
and U5180 (N_5180,N_3976,N_3343);
and U5181 (N_5181,N_1816,N_4395);
and U5182 (N_5182,N_3132,N_1019);
nor U5183 (N_5183,N_4082,N_670);
nand U5184 (N_5184,N_2662,N_3527);
xnor U5185 (N_5185,N_4657,N_3899);
nor U5186 (N_5186,N_2930,N_3066);
nand U5187 (N_5187,N_2906,N_354);
xor U5188 (N_5188,N_1597,N_3995);
or U5189 (N_5189,N_883,N_4332);
nand U5190 (N_5190,N_1086,N_1856);
nor U5191 (N_5191,N_556,N_3071);
nand U5192 (N_5192,N_2876,N_1205);
and U5193 (N_5193,N_295,N_368);
and U5194 (N_5194,N_4044,N_3637);
and U5195 (N_5195,N_4920,N_1908);
nand U5196 (N_5196,N_3,N_3555);
or U5197 (N_5197,N_4706,N_1560);
xnor U5198 (N_5198,N_847,N_3366);
or U5199 (N_5199,N_1281,N_3756);
nor U5200 (N_5200,N_4715,N_1806);
nor U5201 (N_5201,N_1275,N_902);
nand U5202 (N_5202,N_1317,N_2523);
and U5203 (N_5203,N_730,N_1162);
xnor U5204 (N_5204,N_3156,N_346);
nand U5205 (N_5205,N_4381,N_780);
nor U5206 (N_5206,N_3838,N_1580);
or U5207 (N_5207,N_2971,N_3367);
nand U5208 (N_5208,N_385,N_1814);
xnor U5209 (N_5209,N_2038,N_249);
nand U5210 (N_5210,N_2294,N_375);
nor U5211 (N_5211,N_107,N_1677);
nor U5212 (N_5212,N_3486,N_1537);
nor U5213 (N_5213,N_2617,N_3709);
or U5214 (N_5214,N_4145,N_4938);
nor U5215 (N_5215,N_1572,N_2247);
nor U5216 (N_5216,N_961,N_4434);
nand U5217 (N_5217,N_2404,N_2053);
and U5218 (N_5218,N_4602,N_4681);
nand U5219 (N_5219,N_2967,N_4496);
and U5220 (N_5220,N_4269,N_3970);
xnor U5221 (N_5221,N_3313,N_753);
nor U5222 (N_5222,N_3778,N_401);
nor U5223 (N_5223,N_3687,N_1328);
xnor U5224 (N_5224,N_4031,N_4416);
nand U5225 (N_5225,N_1025,N_4119);
and U5226 (N_5226,N_1336,N_392);
nor U5227 (N_5227,N_1651,N_3133);
nor U5228 (N_5228,N_4541,N_1477);
xor U5229 (N_5229,N_45,N_3191);
nor U5230 (N_5230,N_485,N_723);
or U5231 (N_5231,N_994,N_1637);
and U5232 (N_5232,N_4057,N_1163);
or U5233 (N_5233,N_4138,N_160);
and U5234 (N_5234,N_4595,N_4735);
nor U5235 (N_5235,N_871,N_3117);
nand U5236 (N_5236,N_2764,N_4873);
nand U5237 (N_5237,N_3328,N_4330);
xnor U5238 (N_5238,N_3537,N_876);
and U5239 (N_5239,N_2035,N_269);
and U5240 (N_5240,N_4682,N_152);
nand U5241 (N_5241,N_1051,N_4471);
nand U5242 (N_5242,N_2302,N_4386);
or U5243 (N_5243,N_2866,N_1871);
and U5244 (N_5244,N_4286,N_2188);
nor U5245 (N_5245,N_1532,N_3808);
or U5246 (N_5246,N_4830,N_1949);
nand U5247 (N_5247,N_3010,N_3120);
and U5248 (N_5248,N_1590,N_4828);
or U5249 (N_5249,N_2497,N_2327);
nor U5250 (N_5250,N_4863,N_841);
and U5251 (N_5251,N_4594,N_1858);
nor U5252 (N_5252,N_3409,N_3715);
and U5253 (N_5253,N_4618,N_217);
nand U5254 (N_5254,N_4160,N_4669);
and U5255 (N_5255,N_302,N_2533);
and U5256 (N_5256,N_2988,N_1450);
and U5257 (N_5257,N_4433,N_3007);
nand U5258 (N_5258,N_684,N_1294);
nor U5259 (N_5259,N_4225,N_2862);
nor U5260 (N_5260,N_877,N_900);
and U5261 (N_5261,N_1301,N_24);
and U5262 (N_5262,N_2312,N_4383);
xnor U5263 (N_5263,N_4492,N_1914);
and U5264 (N_5264,N_1994,N_3327);
nand U5265 (N_5265,N_538,N_1329);
or U5266 (N_5266,N_590,N_1030);
and U5267 (N_5267,N_4995,N_4936);
and U5268 (N_5268,N_3603,N_1408);
nor U5269 (N_5269,N_4501,N_2171);
or U5270 (N_5270,N_4550,N_4280);
and U5271 (N_5271,N_215,N_4878);
xnor U5272 (N_5272,N_698,N_2536);
and U5273 (N_5273,N_4358,N_2526);
nand U5274 (N_5274,N_3250,N_4001);
or U5275 (N_5275,N_1258,N_1948);
nor U5276 (N_5276,N_1291,N_2374);
nand U5277 (N_5277,N_364,N_2337);
xnor U5278 (N_5278,N_2356,N_351);
nor U5279 (N_5279,N_1380,N_1718);
or U5280 (N_5280,N_3587,N_85);
nor U5281 (N_5281,N_266,N_408);
nand U5282 (N_5282,N_1655,N_1633);
xnor U5283 (N_5283,N_1196,N_2647);
or U5284 (N_5284,N_2136,N_4066);
or U5285 (N_5285,N_2867,N_2805);
nor U5286 (N_5286,N_1314,N_789);
or U5287 (N_5287,N_383,N_845);
nor U5288 (N_5288,N_2687,N_2037);
and U5289 (N_5289,N_221,N_2379);
nand U5290 (N_5290,N_4046,N_4465);
nand U5291 (N_5291,N_3476,N_4884);
nor U5292 (N_5292,N_2215,N_2027);
nor U5293 (N_5293,N_4662,N_572);
xor U5294 (N_5294,N_274,N_3274);
xor U5295 (N_5295,N_4870,N_1851);
nand U5296 (N_5296,N_4729,N_4491);
or U5297 (N_5297,N_3523,N_3815);
and U5298 (N_5298,N_657,N_3719);
xnor U5299 (N_5299,N_641,N_2995);
and U5300 (N_5300,N_1501,N_1569);
or U5301 (N_5301,N_2977,N_3597);
and U5302 (N_5302,N_998,N_1992);
nor U5303 (N_5303,N_2575,N_2697);
or U5304 (N_5304,N_1470,N_4580);
nor U5305 (N_5305,N_382,N_3601);
nand U5306 (N_5306,N_2186,N_3549);
nand U5307 (N_5307,N_3929,N_1483);
nand U5308 (N_5308,N_2591,N_1564);
nand U5309 (N_5309,N_4185,N_2778);
and U5310 (N_5310,N_4782,N_4520);
nor U5311 (N_5311,N_16,N_122);
or U5312 (N_5312,N_1395,N_2417);
and U5313 (N_5313,N_921,N_1415);
xor U5314 (N_5314,N_2444,N_2124);
nor U5315 (N_5315,N_4047,N_4080);
or U5316 (N_5316,N_4274,N_1853);
nor U5317 (N_5317,N_3230,N_1354);
xnor U5318 (N_5318,N_2987,N_437);
nor U5319 (N_5319,N_4037,N_1197);
or U5320 (N_5320,N_4403,N_2467);
and U5321 (N_5321,N_3403,N_2508);
nand U5322 (N_5322,N_3501,N_3998);
nor U5323 (N_5323,N_4021,N_209);
or U5324 (N_5324,N_4069,N_4781);
nor U5325 (N_5325,N_688,N_3375);
xor U5326 (N_5326,N_897,N_335);
nand U5327 (N_5327,N_827,N_1107);
or U5328 (N_5328,N_562,N_3726);
or U5329 (N_5329,N_980,N_2813);
xor U5330 (N_5330,N_1476,N_2589);
or U5331 (N_5331,N_4813,N_4778);
nor U5332 (N_5332,N_873,N_1968);
nand U5333 (N_5333,N_1429,N_3798);
or U5334 (N_5334,N_4724,N_282);
and U5335 (N_5335,N_2130,N_814);
nor U5336 (N_5336,N_337,N_601);
nand U5337 (N_5337,N_842,N_2081);
or U5338 (N_5338,N_3140,N_4306);
nand U5339 (N_5339,N_4048,N_3979);
nor U5340 (N_5340,N_3913,N_1982);
and U5341 (N_5341,N_1523,N_3267);
nand U5342 (N_5342,N_3302,N_4456);
and U5343 (N_5343,N_3800,N_4616);
nand U5344 (N_5344,N_1610,N_1877);
or U5345 (N_5345,N_1414,N_3787);
and U5346 (N_5346,N_4460,N_100);
and U5347 (N_5347,N_2682,N_1355);
nor U5348 (N_5348,N_1670,N_3158);
nor U5349 (N_5349,N_4687,N_272);
nor U5350 (N_5350,N_4567,N_3017);
nor U5351 (N_5351,N_3794,N_433);
or U5352 (N_5352,N_276,N_3177);
or U5353 (N_5353,N_482,N_4800);
and U5354 (N_5354,N_4475,N_132);
nand U5355 (N_5355,N_4446,N_1122);
and U5356 (N_5356,N_3157,N_2103);
and U5357 (N_5357,N_2948,N_3077);
nand U5358 (N_5358,N_3548,N_1112);
and U5359 (N_5359,N_1663,N_1960);
and U5360 (N_5360,N_4421,N_2039);
nor U5361 (N_5361,N_2222,N_4307);
xnor U5362 (N_5362,N_3341,N_1678);
nand U5363 (N_5363,N_1116,N_472);
and U5364 (N_5364,N_3977,N_3425);
nand U5365 (N_5365,N_2611,N_1625);
nand U5366 (N_5366,N_839,N_3087);
nor U5367 (N_5367,N_981,N_3498);
or U5368 (N_5368,N_1409,N_3967);
or U5369 (N_5369,N_941,N_861);
or U5370 (N_5370,N_393,N_4585);
or U5371 (N_5371,N_588,N_977);
and U5372 (N_5372,N_1438,N_3497);
and U5373 (N_5373,N_1680,N_3399);
nor U5374 (N_5374,N_912,N_2838);
xnor U5375 (N_5375,N_2968,N_1936);
and U5376 (N_5376,N_75,N_3949);
nor U5377 (N_5377,N_4390,N_574);
nand U5378 (N_5378,N_3145,N_3676);
nand U5379 (N_5379,N_1350,N_1034);
nor U5380 (N_5380,N_3400,N_4325);
and U5381 (N_5381,N_496,N_4139);
xor U5382 (N_5382,N_1382,N_2168);
or U5383 (N_5383,N_1912,N_2433);
nor U5384 (N_5384,N_478,N_3851);
and U5385 (N_5385,N_2384,N_2173);
nand U5386 (N_5386,N_1038,N_3775);
xnor U5387 (N_5387,N_3252,N_1444);
and U5388 (N_5388,N_4727,N_787);
nand U5389 (N_5389,N_4427,N_596);
and U5390 (N_5390,N_4647,N_2998);
nor U5391 (N_5391,N_529,N_3163);
or U5392 (N_5392,N_3053,N_2000);
nor U5393 (N_5393,N_3912,N_3568);
nand U5394 (N_5394,N_2918,N_1262);
or U5395 (N_5395,N_3026,N_2932);
or U5396 (N_5396,N_3684,N_277);
nand U5397 (N_5397,N_2844,N_1499);
nand U5398 (N_5398,N_1286,N_4022);
nand U5399 (N_5399,N_4755,N_652);
and U5400 (N_5400,N_1913,N_691);
xor U5401 (N_5401,N_2386,N_1588);
and U5402 (N_5402,N_3222,N_3037);
nor U5403 (N_5403,N_4055,N_3564);
and U5404 (N_5404,N_41,N_3722);
or U5405 (N_5405,N_3479,N_1422);
nor U5406 (N_5406,N_971,N_384);
nand U5407 (N_5407,N_4886,N_3239);
or U5408 (N_5408,N_2559,N_1029);
and U5409 (N_5409,N_4970,N_3729);
and U5410 (N_5410,N_3645,N_1699);
and U5411 (N_5411,N_1062,N_2984);
and U5412 (N_5412,N_3418,N_419);
nand U5413 (N_5413,N_3235,N_2274);
nand U5414 (N_5414,N_3866,N_647);
nand U5415 (N_5415,N_211,N_285);
or U5416 (N_5416,N_1121,N_2801);
xnor U5417 (N_5417,N_945,N_2472);
xor U5418 (N_5418,N_127,N_521);
or U5419 (N_5419,N_1325,N_28);
and U5420 (N_5420,N_2715,N_1407);
and U5421 (N_5421,N_1782,N_4815);
nand U5422 (N_5422,N_2322,N_3591);
nor U5423 (N_5423,N_199,N_464);
nand U5424 (N_5424,N_1012,N_1095);
nor U5425 (N_5425,N_2345,N_3779);
and U5426 (N_5426,N_3630,N_438);
and U5427 (N_5427,N_2994,N_352);
nor U5428 (N_5428,N_1993,N_4771);
or U5429 (N_5429,N_4118,N_4218);
nor U5430 (N_5430,N_2143,N_436);
nor U5431 (N_5431,N_4226,N_2746);
nand U5432 (N_5432,N_3060,N_3482);
nand U5433 (N_5433,N_2815,N_134);
nor U5434 (N_5434,N_577,N_3291);
and U5435 (N_5435,N_1688,N_2516);
xor U5436 (N_5436,N_2228,N_2855);
nor U5437 (N_5437,N_1252,N_2391);
or U5438 (N_5438,N_4070,N_974);
nor U5439 (N_5439,N_4391,N_4299);
or U5440 (N_5440,N_4632,N_2643);
or U5441 (N_5441,N_978,N_4207);
nand U5442 (N_5442,N_3093,N_3727);
nand U5443 (N_5443,N_1567,N_3543);
and U5444 (N_5444,N_369,N_1428);
nor U5445 (N_5445,N_2751,N_3546);
or U5446 (N_5446,N_3217,N_604);
nand U5447 (N_5447,N_431,N_4934);
and U5448 (N_5448,N_3784,N_1011);
nand U5449 (N_5449,N_3805,N_1456);
nand U5450 (N_5450,N_2034,N_704);
nand U5451 (N_5451,N_923,N_4262);
and U5452 (N_5452,N_2289,N_2587);
nor U5453 (N_5453,N_3242,N_3430);
nor U5454 (N_5454,N_585,N_2028);
xor U5455 (N_5455,N_144,N_1115);
nor U5456 (N_5456,N_651,N_2253);
nor U5457 (N_5457,N_3539,N_3127);
nand U5458 (N_5458,N_101,N_1498);
nand U5459 (N_5459,N_1777,N_1364);
xnor U5460 (N_5460,N_1344,N_89);
or U5461 (N_5461,N_1885,N_626);
nand U5462 (N_5462,N_4607,N_1847);
and U5463 (N_5463,N_4241,N_4402);
and U5464 (N_5464,N_1808,N_4821);
and U5465 (N_5465,N_4810,N_868);
and U5466 (N_5466,N_2928,N_4919);
nor U5467 (N_5467,N_1278,N_4015);
nand U5468 (N_5468,N_4196,N_2004);
and U5469 (N_5469,N_3160,N_3002);
or U5470 (N_5470,N_1053,N_1473);
and U5471 (N_5471,N_4056,N_4608);
or U5472 (N_5472,N_4927,N_928);
and U5473 (N_5473,N_3861,N_3571);
nor U5474 (N_5474,N_4911,N_2030);
or U5475 (N_5475,N_1807,N_4588);
and U5476 (N_5476,N_2166,N_4164);
xor U5477 (N_5477,N_4140,N_4079);
or U5478 (N_5478,N_4418,N_1901);
and U5479 (N_5479,N_2661,N_4807);
nor U5480 (N_5480,N_1103,N_660);
xnor U5481 (N_5481,N_1403,N_4468);
and U5482 (N_5482,N_3365,N_442);
or U5483 (N_5483,N_2152,N_212);
xnor U5484 (N_5484,N_748,N_2354);
or U5485 (N_5485,N_812,N_4940);
nor U5486 (N_5486,N_4716,N_3959);
or U5487 (N_5487,N_3042,N_1929);
or U5488 (N_5488,N_2668,N_769);
and U5489 (N_5489,N_826,N_30);
or U5490 (N_5490,N_306,N_4923);
xor U5491 (N_5491,N_4265,N_4452);
nor U5492 (N_5492,N_3169,N_3362);
xnor U5493 (N_5493,N_2795,N_2842);
or U5494 (N_5494,N_3059,N_3991);
nand U5495 (N_5495,N_4915,N_108);
xor U5496 (N_5496,N_1900,N_366);
nor U5497 (N_5497,N_1058,N_1552);
or U5498 (N_5498,N_1279,N_2221);
or U5499 (N_5499,N_4984,N_2959);
and U5500 (N_5500,N_4011,N_783);
and U5501 (N_5501,N_110,N_1302);
nor U5502 (N_5502,N_709,N_4032);
xnor U5503 (N_5503,N_1516,N_968);
nor U5504 (N_5504,N_4944,N_4888);
or U5505 (N_5505,N_4869,N_1823);
and U5506 (N_5506,N_4338,N_3574);
nor U5507 (N_5507,N_3384,N_4679);
and U5508 (N_5508,N_4825,N_4394);
nand U5509 (N_5509,N_746,N_4745);
and U5510 (N_5510,N_1826,N_178);
nand U5511 (N_5511,N_1315,N_2797);
xnor U5512 (N_5512,N_1903,N_3994);
nor U5513 (N_5513,N_4072,N_4613);
or U5514 (N_5514,N_2290,N_4366);
nand U5515 (N_5515,N_2364,N_2181);
xor U5516 (N_5516,N_4405,N_2828);
nand U5517 (N_5517,N_2493,N_2799);
or U5518 (N_5518,N_1926,N_3441);
xnor U5519 (N_5519,N_4592,N_394);
nor U5520 (N_5520,N_1145,N_1207);
xnor U5521 (N_5521,N_1768,N_2775);
nor U5522 (N_5522,N_3179,N_3013);
nand U5523 (N_5523,N_258,N_2304);
xnor U5524 (N_5524,N_4758,N_4960);
xor U5525 (N_5525,N_1773,N_333);
or U5526 (N_5526,N_4981,N_4876);
nor U5527 (N_5527,N_1969,N_297);
and U5528 (N_5528,N_136,N_1179);
nor U5529 (N_5529,N_3605,N_1240);
nor U5530 (N_5530,N_1031,N_2388);
nand U5531 (N_5531,N_4779,N_46);
and U5532 (N_5532,N_1701,N_3440);
nand U5533 (N_5533,N_1003,N_1157);
or U5534 (N_5534,N_4310,N_2457);
xor U5535 (N_5535,N_1126,N_1394);
and U5536 (N_5536,N_4776,N_3685);
and U5537 (N_5537,N_1642,N_2449);
nand U5538 (N_5538,N_1525,N_3086);
xnor U5539 (N_5539,N_2276,N_78);
and U5540 (N_5540,N_4378,N_2425);
nand U5541 (N_5541,N_4955,N_2698);
xor U5542 (N_5542,N_3819,N_1544);
nor U5543 (N_5543,N_2496,N_4989);
and U5544 (N_5544,N_1253,N_3933);
or U5545 (N_5545,N_1687,N_4186);
and U5546 (N_5546,N_2203,N_2822);
xor U5547 (N_5547,N_3215,N_2409);
or U5548 (N_5548,N_467,N_3532);
and U5549 (N_5549,N_3317,N_4227);
or U5550 (N_5550,N_2085,N_887);
and U5551 (N_5551,N_1859,N_1843);
and U5552 (N_5552,N_3765,N_707);
and U5553 (N_5553,N_4875,N_483);
nand U5554 (N_5554,N_140,N_1299);
and U5555 (N_5555,N_1512,N_1137);
xnor U5556 (N_5556,N_4544,N_4563);
or U5557 (N_5557,N_4698,N_4748);
nor U5558 (N_5558,N_3073,N_2958);
and U5559 (N_5559,N_2951,N_3454);
and U5560 (N_5560,N_3212,N_2677);
or U5561 (N_5561,N_2820,N_2990);
or U5562 (N_5562,N_2262,N_1650);
or U5563 (N_5563,N_2893,N_3559);
nand U5564 (N_5564,N_3656,N_2072);
nor U5565 (N_5565,N_4658,N_410);
and U5566 (N_5566,N_2089,N_2058);
or U5567 (N_5567,N_1977,N_2962);
or U5568 (N_5568,N_2454,N_197);
nand U5569 (N_5569,N_3954,N_1839);
and U5570 (N_5570,N_311,N_2628);
nand U5571 (N_5571,N_2342,N_4444);
nor U5572 (N_5572,N_1047,N_2137);
or U5573 (N_5573,N_986,N_4696);
nand U5574 (N_5574,N_246,N_3461);
xor U5575 (N_5575,N_3345,N_1232);
or U5576 (N_5576,N_2832,N_3286);
nor U5577 (N_5577,N_3890,N_686);
nor U5578 (N_5578,N_331,N_4559);
xor U5579 (N_5579,N_2907,N_2989);
nand U5580 (N_5580,N_234,N_714);
and U5581 (N_5581,N_2392,N_3371);
or U5582 (N_5582,N_1507,N_2450);
and U5583 (N_5583,N_181,N_3650);
and U5584 (N_5584,N_2403,N_3960);
and U5585 (N_5585,N_3924,N_4621);
and U5586 (N_5586,N_2970,N_927);
xnor U5587 (N_5587,N_360,N_2727);
and U5588 (N_5588,N_4722,N_2295);
nand U5589 (N_5589,N_1792,N_1704);
nor U5590 (N_5590,N_741,N_210);
nand U5591 (N_5591,N_550,N_2674);
nor U5592 (N_5592,N_882,N_3223);
nand U5593 (N_5593,N_2,N_3337);
or U5594 (N_5594,N_3885,N_4850);
or U5595 (N_5595,N_1894,N_1756);
nor U5596 (N_5596,N_4013,N_547);
or U5597 (N_5597,N_4347,N_3817);
or U5598 (N_5598,N_4604,N_32);
and U5599 (N_5599,N_2857,N_2814);
or U5600 (N_5600,N_2639,N_4510);
nand U5601 (N_5601,N_1528,N_3236);
or U5602 (N_5602,N_2941,N_3346);
or U5603 (N_5603,N_1739,N_595);
nor U5604 (N_5604,N_224,N_171);
nor U5605 (N_5605,N_4536,N_316);
nor U5606 (N_5606,N_4272,N_3288);
nand U5607 (N_5607,N_4728,N_1078);
and U5608 (N_5608,N_1746,N_1335);
nand U5609 (N_5609,N_4219,N_2140);
and U5610 (N_5610,N_3968,N_2782);
nor U5611 (N_5611,N_3623,N_972);
nand U5612 (N_5612,N_2358,N_3474);
nor U5613 (N_5613,N_1744,N_4478);
nor U5614 (N_5614,N_3661,N_4205);
nor U5615 (N_5615,N_3392,N_2052);
nand U5616 (N_5616,N_2422,N_2885);
and U5617 (N_5617,N_1891,N_3649);
or U5618 (N_5618,N_2942,N_964);
nor U5619 (N_5619,N_4584,N_3485);
or U5620 (N_5620,N_560,N_1218);
nand U5621 (N_5621,N_1641,N_149);
xnor U5622 (N_5622,N_908,N_2284);
nor U5623 (N_5623,N_4263,N_330);
xor U5624 (N_5624,N_1709,N_4935);
or U5625 (N_5625,N_1889,N_543);
nor U5626 (N_5626,N_3610,N_2243);
nor U5627 (N_5627,N_3436,N_3326);
nor U5628 (N_5628,N_4708,N_4656);
nor U5629 (N_5629,N_4649,N_615);
xnor U5630 (N_5630,N_3871,N_1556);
or U5631 (N_5631,N_3836,N_4639);
or U5632 (N_5632,N_2258,N_791);
or U5633 (N_5633,N_2593,N_3178);
or U5634 (N_5634,N_1573,N_3203);
or U5635 (N_5635,N_2500,N_3975);
or U5636 (N_5636,N_1636,N_97);
or U5637 (N_5637,N_1962,N_4003);
or U5638 (N_5638,N_2474,N_468);
nor U5639 (N_5639,N_3761,N_4519);
and U5640 (N_5640,N_569,N_2678);
nand U5641 (N_5641,N_2275,N_661);
or U5642 (N_5642,N_2710,N_823);
or U5643 (N_5643,N_1442,N_3283);
nand U5644 (N_5644,N_3528,N_3031);
nor U5645 (N_5645,N_4705,N_735);
and U5646 (N_5646,N_1489,N_4052);
nor U5647 (N_5647,N_1369,N_1741);
or U5648 (N_5648,N_3170,N_3606);
or U5649 (N_5649,N_1059,N_3005);
nand U5650 (N_5650,N_1951,N_3428);
nand U5651 (N_5651,N_4000,N_522);
or U5652 (N_5652,N_813,N_2242);
or U5653 (N_5653,N_434,N_4785);
nor U5654 (N_5654,N_1661,N_18);
nand U5655 (N_5655,N_2931,N_2882);
and U5656 (N_5656,N_1201,N_677);
or U5657 (N_5657,N_3385,N_133);
nor U5658 (N_5658,N_2106,N_3374);
nor U5659 (N_5659,N_761,N_4942);
nand U5660 (N_5660,N_2956,N_4926);
or U5661 (N_5661,N_2133,N_473);
nor U5662 (N_5662,N_513,N_1543);
nor U5663 (N_5663,N_3225,N_84);
or U5664 (N_5664,N_3098,N_1645);
nand U5665 (N_5665,N_2625,N_3541);
or U5666 (N_5666,N_94,N_1371);
xnor U5667 (N_5667,N_975,N_3134);
xor U5668 (N_5668,N_717,N_916);
xnor U5669 (N_5669,N_4323,N_3146);
or U5670 (N_5670,N_4027,N_50);
nor U5671 (N_5671,N_310,N_1285);
and U5672 (N_5672,N_3653,N_172);
and U5673 (N_5673,N_3631,N_3055);
or U5674 (N_5674,N_2537,N_4308);
nand U5675 (N_5675,N_2196,N_559);
or U5676 (N_5676,N_3598,N_2389);
or U5677 (N_5677,N_1848,N_481);
or U5678 (N_5678,N_4983,N_1596);
or U5679 (N_5679,N_985,N_1541);
nand U5680 (N_5680,N_4450,N_949);
and U5681 (N_5681,N_951,N_1713);
or U5682 (N_5682,N_1732,N_2895);
nor U5683 (N_5683,N_676,N_4472);
and U5684 (N_5684,N_4163,N_4317);
xnor U5685 (N_5685,N_878,N_4751);
nand U5686 (N_5686,N_1368,N_2344);
and U5687 (N_5687,N_2046,N_3092);
or U5688 (N_5688,N_1549,N_2498);
xnor U5689 (N_5689,N_3749,N_2713);
xor U5690 (N_5690,N_2519,N_3942);
nor U5691 (N_5691,N_2807,N_2843);
nand U5692 (N_5692,N_1384,N_4978);
xnor U5693 (N_5693,N_3529,N_1203);
nand U5694 (N_5694,N_4910,N_70);
xor U5695 (N_5695,N_3159,N_4814);
and U5696 (N_5696,N_151,N_3677);
nand U5697 (N_5697,N_806,N_1606);
nand U5698 (N_5698,N_1707,N_3126);
or U5699 (N_5699,N_2241,N_619);
nand U5700 (N_5700,N_2808,N_2877);
and U5701 (N_5701,N_92,N_22);
nor U5702 (N_5702,N_4388,N_2898);
and U5703 (N_5703,N_3048,N_3231);
xnor U5704 (N_5704,N_1410,N_4179);
or U5705 (N_5705,N_3491,N_1211);
nor U5706 (N_5706,N_2227,N_2528);
nand U5707 (N_5707,N_4088,N_4282);
nor U5708 (N_5708,N_1497,N_1693);
nand U5709 (N_5709,N_1695,N_2742);
or U5710 (N_5710,N_1318,N_611);
and U5711 (N_5711,N_3240,N_4065);
xnor U5712 (N_5712,N_571,N_4849);
nor U5713 (N_5713,N_3421,N_3758);
and U5714 (N_5714,N_1358,N_4293);
nor U5715 (N_5715,N_4528,N_4932);
nand U5716 (N_5716,N_4436,N_4334);
and U5717 (N_5717,N_4147,N_21);
nor U5718 (N_5718,N_976,N_3226);
and U5719 (N_5719,N_3459,N_555);
nor U5720 (N_5720,N_3921,N_320);
or U5721 (N_5721,N_3285,N_3621);
and U5722 (N_5722,N_3054,N_4671);
or U5723 (N_5723,N_1147,N_3593);
nand U5724 (N_5724,N_2303,N_2879);
or U5725 (N_5725,N_1184,N_3167);
or U5726 (N_5726,N_4281,N_2145);
and U5727 (N_5727,N_1820,N_349);
nor U5728 (N_5728,N_33,N_2291);
and U5729 (N_5729,N_1272,N_4353);
and U5730 (N_5730,N_124,N_4178);
and U5731 (N_5731,N_4093,N_1448);
or U5732 (N_5732,N_358,N_2309);
nand U5733 (N_5733,N_3452,N_3567);
or U5734 (N_5734,N_313,N_856);
nor U5735 (N_5735,N_1093,N_1170);
nor U5736 (N_5736,N_4212,N_3221);
or U5737 (N_5737,N_3802,N_145);
and U5738 (N_5738,N_3897,N_240);
nand U5739 (N_5739,N_982,N_3100);
nand U5740 (N_5740,N_1071,N_4652);
xor U5741 (N_5741,N_4576,N_3860);
nand U5742 (N_5742,N_2521,N_1568);
nor U5743 (N_5743,N_3865,N_2355);
and U5744 (N_5744,N_147,N_800);
and U5745 (N_5745,N_1327,N_3820);
and U5746 (N_5746,N_4853,N_524);
nor U5747 (N_5747,N_4835,N_2620);
and U5748 (N_5748,N_612,N_3533);
nand U5749 (N_5749,N_3972,N_1445);
nand U5750 (N_5750,N_844,N_3207);
nand U5751 (N_5751,N_2129,N_1182);
and U5752 (N_5752,N_1055,N_3944);
nand U5753 (N_5753,N_4887,N_4666);
and U5754 (N_5754,N_1441,N_3251);
and U5755 (N_5755,N_4297,N_3030);
nor U5756 (N_5756,N_1319,N_3816);
xor U5757 (N_5757,N_3829,N_2170);
or U5758 (N_5758,N_1172,N_4339);
or U5759 (N_5759,N_2983,N_4798);
nor U5760 (N_5760,N_2213,N_2199);
and U5761 (N_5761,N_1465,N_4949);
or U5762 (N_5762,N_3916,N_872);
or U5763 (N_5763,N_4474,N_36);
nor U5764 (N_5764,N_4531,N_606);
and U5765 (N_5765,N_565,N_3785);
and U5766 (N_5766,N_2405,N_1373);
nand U5767 (N_5767,N_4217,N_3359);
nor U5768 (N_5768,N_3691,N_3121);
or U5769 (N_5769,N_1802,N_4399);
and U5770 (N_5770,N_2878,N_1094);
and U5771 (N_5771,N_2162,N_2119);
nor U5772 (N_5772,N_57,N_2927);
or U5773 (N_5773,N_3183,N_2725);
nand U5774 (N_5774,N_2925,N_4717);
nor U5775 (N_5775,N_2633,N_3039);
and U5776 (N_5776,N_4095,N_3766);
and U5777 (N_5777,N_2552,N_1288);
nand U5778 (N_5778,N_584,N_956);
and U5779 (N_5779,N_3717,N_3277);
nand U5780 (N_5780,N_663,N_2585);
nor U5781 (N_5781,N_2254,N_3149);
nand U5782 (N_5782,N_4837,N_13);
or U5783 (N_5783,N_895,N_300);
and U5784 (N_5784,N_1032,N_2486);
or U5785 (N_5785,N_3464,N_2765);
nand U5786 (N_5786,N_3206,N_512);
or U5787 (N_5787,N_2428,N_2128);
or U5788 (N_5788,N_3185,N_4355);
nand U5789 (N_5789,N_777,N_3864);
and U5790 (N_5790,N_4131,N_2259);
nand U5791 (N_5791,N_4931,N_3551);
and U5792 (N_5792,N_4816,N_495);
and U5793 (N_5793,N_2604,N_1475);
or U5794 (N_5794,N_3136,N_3431);
nand U5795 (N_5795,N_4350,N_3142);
nor U5796 (N_5796,N_4546,N_3494);
nor U5797 (N_5797,N_4285,N_4792);
nand U5798 (N_5798,N_4533,N_1084);
or U5799 (N_5799,N_583,N_2370);
nand U5800 (N_5800,N_1978,N_3561);
and U5801 (N_5801,N_4189,N_1819);
and U5802 (N_5802,N_248,N_1437);
nor U5803 (N_5803,N_3745,N_2271);
and U5804 (N_5804,N_2329,N_910);
xor U5805 (N_5805,N_2982,N_2688);
or U5806 (N_5806,N_3445,N_2502);
and U5807 (N_5807,N_1494,N_3522);
or U5808 (N_5808,N_4879,N_1592);
or U5809 (N_5809,N_3173,N_1671);
or U5810 (N_5810,N_2561,N_4644);
xnor U5811 (N_5811,N_534,N_797);
nand U5812 (N_5812,N_1761,N_2739);
nor U5813 (N_5813,N_237,N_3102);
nand U5814 (N_5814,N_848,N_795);
xor U5815 (N_5815,N_3869,N_2219);
or U5816 (N_5816,N_304,N_3689);
and U5817 (N_5817,N_2331,N_630);
nand U5818 (N_5818,N_8,N_906);
or U5819 (N_5819,N_4401,N_2517);
or U5820 (N_5820,N_2094,N_3137);
nand U5821 (N_5821,N_1142,N_1952);
nand U5822 (N_5822,N_336,N_552);
nand U5823 (N_5823,N_4842,N_3232);
and U5824 (N_5824,N_4165,N_1425);
nand U5825 (N_5825,N_617,N_3058);
nor U5826 (N_5826,N_4290,N_2278);
nor U5827 (N_5827,N_1775,N_4143);
nor U5828 (N_5828,N_261,N_1595);
and U5829 (N_5829,N_4638,N_1947);
nand U5830 (N_5830,N_1138,N_4511);
nand U5831 (N_5831,N_4609,N_857);
xor U5832 (N_5832,N_0,N_4060);
nor U5833 (N_5833,N_805,N_784);
nor U5834 (N_5834,N_523,N_3470);
nor U5835 (N_5835,N_454,N_581);
nand U5836 (N_5836,N_301,N_593);
nor U5837 (N_5837,N_511,N_82);
or U5838 (N_5838,N_1697,N_3003);
and U5839 (N_5839,N_825,N_3334);
or U5840 (N_5840,N_600,N_3329);
xor U5841 (N_5841,N_4881,N_4198);
and U5842 (N_5842,N_909,N_1063);
nand U5843 (N_5843,N_4158,N_1006);
or U5844 (N_5844,N_3636,N_2063);
xor U5845 (N_5845,N_4759,N_2307);
or U5846 (N_5846,N_2507,N_3827);
nor U5847 (N_5847,N_3880,N_3734);
and U5848 (N_5848,N_4710,N_1904);
and U5849 (N_5849,N_1146,N_1664);
and U5850 (N_5850,N_3439,N_120);
and U5851 (N_5851,N_2540,N_2318);
nand U5852 (N_5852,N_1975,N_3151);
or U5853 (N_5853,N_2757,N_3710);
nand U5854 (N_5854,N_3253,N_1037);
nor U5855 (N_5855,N_40,N_1938);
nand U5856 (N_5856,N_2488,N_444);
nand U5857 (N_5857,N_175,N_2789);
nor U5858 (N_5858,N_3742,N_4577);
nand U5859 (N_5859,N_1794,N_2871);
or U5860 (N_5860,N_750,N_4210);
or U5861 (N_5861,N_1457,N_2680);
nor U5862 (N_5862,N_1720,N_2572);
nor U5863 (N_5863,N_2719,N_1559);
nand U5864 (N_5864,N_2475,N_1004);
nand U5865 (N_5865,N_757,N_3467);
and U5866 (N_5866,N_1694,N_4612);
nor U5867 (N_5867,N_287,N_679);
and U5868 (N_5868,N_4796,N_166);
and U5869 (N_5869,N_2641,N_123);
nor U5870 (N_5870,N_973,N_736);
nand U5871 (N_5871,N_2656,N_1956);
xnor U5872 (N_5872,N_2861,N_1090);
or U5873 (N_5873,N_4635,N_222);
or U5874 (N_5874,N_2138,N_4552);
nand U5875 (N_5875,N_3917,N_339);
xnor U5876 (N_5876,N_216,N_1980);
and U5877 (N_5877,N_4103,N_689);
or U5878 (N_5878,N_2382,N_3351);
nor U5879 (N_5879,N_1740,N_4951);
xnor U5880 (N_5880,N_2047,N_4868);
or U5881 (N_5881,N_3502,N_3646);
or U5882 (N_5882,N_3307,N_235);
nand U5883 (N_5883,N_2212,N_1881);
nand U5884 (N_5884,N_1248,N_2399);
and U5885 (N_5885,N_3107,N_413);
nor U5886 (N_5886,N_2401,N_2726);
and U5887 (N_5887,N_426,N_163);
and U5888 (N_5888,N_4569,N_3368);
nor U5889 (N_5889,N_808,N_3809);
nand U5890 (N_5890,N_3083,N_2769);
nand U5891 (N_5891,N_3900,N_685);
or U5892 (N_5892,N_2875,N_2340);
and U5893 (N_5893,N_3904,N_227);
nor U5894 (N_5894,N_1638,N_4598);
nor U5895 (N_5895,N_1000,N_1065);
nand U5896 (N_5896,N_3669,N_1020);
and U5897 (N_5897,N_1131,N_558);
xor U5898 (N_5898,N_4606,N_2135);
nor U5899 (N_5899,N_254,N_3279);
nand U5900 (N_5900,N_4172,N_1096);
nand U5901 (N_5901,N_2460,N_3097);
and U5902 (N_5902,N_4772,N_31);
xor U5903 (N_5903,N_2044,N_2638);
or U5904 (N_5904,N_4345,N_416);
or U5905 (N_5905,N_4709,N_378);
and U5906 (N_5906,N_4368,N_1127);
nor U5907 (N_5907,N_2237,N_616);
nor U5908 (N_5908,N_1459,N_2314);
nand U5909 (N_5909,N_758,N_2139);
nand U5910 (N_5910,N_4973,N_4673);
nor U5911 (N_5911,N_4034,N_1469);
nor U5912 (N_5912,N_774,N_2102);
or U5913 (N_5913,N_2015,N_4848);
or U5914 (N_5914,N_580,N_1391);
nand U5915 (N_5915,N_969,N_3629);
nor U5916 (N_5916,N_391,N_4547);
nand U5917 (N_5917,N_4166,N_3080);
nand U5918 (N_5918,N_913,N_3509);
and U5919 (N_5919,N_262,N_811);
nand U5920 (N_5920,N_2793,N_835);
nand U5921 (N_5921,N_2874,N_1745);
or U5922 (N_5922,N_1072,N_4665);
and U5923 (N_5923,N_2368,N_1353);
or U5924 (N_5924,N_1367,N_4493);
nor U5925 (N_5925,N_2938,N_2174);
and U5926 (N_5926,N_3516,N_2665);
or U5927 (N_5927,N_430,N_1451);
or U5928 (N_5928,N_794,N_4376);
xnor U5929 (N_5929,N_1052,N_3507);
nor U5930 (N_5930,N_4565,N_4626);
nor U5931 (N_5931,N_2518,N_3791);
or U5932 (N_5932,N_2265,N_4894);
xnor U5933 (N_5933,N_4233,N_3712);
or U5934 (N_5934,N_1330,N_3813);
nor U5935 (N_5935,N_1526,N_4556);
nor U5936 (N_5936,N_768,N_182);
xor U5937 (N_5937,N_1605,N_1941);
or U5938 (N_5938,N_3833,N_1979);
or U5939 (N_5939,N_1649,N_3460);
and U5940 (N_5940,N_1290,N_4007);
or U5941 (N_5941,N_3489,N_3750);
nor U5942 (N_5942,N_1765,N_362);
or U5943 (N_5943,N_2306,N_1621);
or U5944 (N_5944,N_1931,N_47);
and U5945 (N_5945,N_589,N_329);
xnor U5946 (N_5946,N_288,N_3850);
or U5947 (N_5947,N_2407,N_1124);
nand U5948 (N_5948,N_305,N_3112);
nor U5949 (N_5949,N_2009,N_4251);
nor U5950 (N_5950,N_1829,N_4587);
nand U5951 (N_5951,N_3124,N_2602);
or U5952 (N_5952,N_1958,N_4763);
xor U5953 (N_5953,N_15,N_4438);
and U5954 (N_5954,N_2236,N_3228);
xor U5955 (N_5955,N_778,N_1303);
and U5956 (N_5956,N_1479,N_1164);
and U5957 (N_5957,N_3918,N_4049);
and U5958 (N_5958,N_860,N_765);
nor U5959 (N_5959,N_3198,N_4254);
and U5960 (N_5960,N_3665,N_4783);
or U5961 (N_5961,N_2900,N_2465);
nand U5962 (N_5962,N_3948,N_716);
and U5963 (N_5963,N_1342,N_3259);
nand U5964 (N_5964,N_665,N_1548);
nor U5965 (N_5965,N_3082,N_3433);
nand U5966 (N_5966,N_3695,N_1064);
or U5967 (N_5967,N_4243,N_4653);
nor U5968 (N_5968,N_1917,N_3472);
nor U5969 (N_5969,N_2936,N_2883);
or U5970 (N_5970,N_2510,N_1089);
nor U5971 (N_5971,N_2095,N_3295);
and U5972 (N_5972,N_4836,N_4864);
or U5973 (N_5973,N_1230,N_4757);
or U5974 (N_5974,N_1458,N_2283);
nand U5975 (N_5975,N_3927,N_1361);
nor U5976 (N_5976,N_3216,N_2461);
and U5977 (N_5977,N_3797,N_3911);
and U5978 (N_5978,N_4026,N_2297);
nor U5979 (N_5979,N_2261,N_1550);
xnor U5980 (N_5980,N_3473,N_527);
and U5981 (N_5981,N_3611,N_2946);
nor U5982 (N_5982,N_2693,N_659);
nand U5983 (N_5983,N_1922,N_4087);
or U5984 (N_5984,N_4130,N_3618);
or U5985 (N_5985,N_3118,N_2109);
or U5986 (N_5986,N_1893,N_4154);
nor U5987 (N_5987,N_2920,N_3999);
nor U5988 (N_5988,N_2864,N_4743);
and U5989 (N_5989,N_3052,N_1023);
nor U5990 (N_5990,N_3402,N_3520);
and U5991 (N_5991,N_3519,N_2599);
or U5992 (N_5992,N_2269,N_2190);
or U5993 (N_5993,N_3238,N_3965);
and U5994 (N_5994,N_4897,N_3642);
nand U5995 (N_5995,N_2352,N_2578);
or U5996 (N_5996,N_1800,N_2557);
and U5997 (N_5997,N_4380,N_634);
nor U5998 (N_5998,N_4903,N_1866);
or U5999 (N_5999,N_4063,N_2022);
nor U6000 (N_6000,N_930,N_2992);
nor U6001 (N_6001,N_2430,N_4128);
nand U6002 (N_6002,N_4898,N_1129);
nor U6003 (N_6003,N_4558,N_3952);
nand U6004 (N_6004,N_3196,N_2790);
nor U6005 (N_6005,N_2120,N_3580);
nand U6006 (N_6006,N_374,N_1887);
xor U6007 (N_6007,N_3697,N_2901);
or U6008 (N_6008,N_3996,N_3280);
or U6009 (N_6009,N_896,N_4489);
and U6010 (N_6010,N_1673,N_2260);
xor U6011 (N_6011,N_213,N_2083);
nor U6012 (N_6012,N_3197,N_3450);
nor U6013 (N_6013,N_4668,N_4941);
xor U6014 (N_6014,N_2631,N_1736);
nor U6015 (N_6015,N_955,N_206);
nand U6016 (N_6016,N_1608,N_2630);
or U6017 (N_6017,N_1577,N_2277);
and U6018 (N_6018,N_4206,N_3114);
or U6019 (N_6019,N_4948,N_1351);
or U6020 (N_6020,N_4331,N_991);
or U6021 (N_6021,N_915,N_1028);
nor U6022 (N_6022,N_2248,N_2134);
or U6023 (N_6023,N_4827,N_2159);
nand U6024 (N_6024,N_2762,N_370);
or U6025 (N_6025,N_867,N_1769);
nor U6026 (N_6026,N_517,N_2570);
nor U6027 (N_6027,N_1875,N_2512);
xor U6028 (N_6028,N_1690,N_3171);
and U6029 (N_6029,N_1271,N_4102);
and U6030 (N_6030,N_2881,N_154);
and U6031 (N_6031,N_3557,N_3780);
xor U6032 (N_6032,N_3190,N_586);
and U6033 (N_6033,N_1156,N_4442);
xor U6034 (N_6034,N_4354,N_4012);
nand U6035 (N_6035,N_720,N_2997);
or U6036 (N_6036,N_2595,N_491);
nor U6037 (N_6037,N_3210,N_693);
nand U6038 (N_6038,N_4393,N_4244);
nand U6039 (N_6039,N_654,N_2600);
or U6040 (N_6040,N_3620,N_2263);
xor U6041 (N_6041,N_4683,N_1150);
xor U6042 (N_6042,N_1824,N_3595);
nand U6043 (N_6043,N_1181,N_1388);
nand U6044 (N_6044,N_1522,N_2036);
or U6045 (N_6045,N_2273,N_1876);
and U6046 (N_6046,N_4371,N_2657);
nor U6047 (N_6047,N_3404,N_940);
and U6048 (N_6048,N_4352,N_4543);
nand U6049 (N_6049,N_4086,N_544);
or U6050 (N_6050,N_533,N_3941);
or U6051 (N_6051,N_2547,N_3859);
nor U6052 (N_6052,N_1542,N_793);
and U6053 (N_6053,N_2543,N_3760);
xor U6054 (N_6054,N_236,N_1198);
or U6055 (N_6055,N_4818,N_4035);
and U6056 (N_6056,N_3325,N_4521);
or U6057 (N_6057,N_1305,N_1725);
or U6058 (N_6058,N_548,N_1069);
or U6059 (N_6059,N_4939,N_3773);
nand U6060 (N_6060,N_95,N_2092);
nand U6061 (N_6061,N_4913,N_105);
or U6062 (N_6062,N_3566,N_4986);
nor U6063 (N_6063,N_3703,N_345);
nand U6064 (N_6064,N_2614,N_3713);
nand U6065 (N_6065,N_506,N_636);
nand U6066 (N_6066,N_4557,N_4633);
and U6067 (N_6067,N_2753,N_1466);
nand U6068 (N_6068,N_4802,N_381);
and U6069 (N_6069,N_498,N_2185);
xor U6070 (N_6070,N_4062,N_4997);
nor U6071 (N_6071,N_3488,N_4952);
nor U6072 (N_6072,N_4204,N_3195);
nand U6073 (N_6073,N_4209,N_3801);
nand U6074 (N_6074,N_537,N_4273);
nand U6075 (N_6075,N_1626,N_421);
nor U6076 (N_6076,N_2390,N_2335);
or U6077 (N_6077,N_4137,N_3662);
and U6078 (N_6078,N_2908,N_2031);
and U6079 (N_6079,N_3893,N_4640);
or U6080 (N_6080,N_950,N_816);
and U6081 (N_6081,N_2202,N_2891);
nand U6082 (N_6082,N_3255,N_3338);
nand U6083 (N_6083,N_715,N_4157);
nand U6084 (N_6084,N_4453,N_1443);
or U6085 (N_6085,N_4170,N_3332);
nand U6086 (N_6086,N_4907,N_3333);
or U6087 (N_6087,N_4617,N_3517);
or U6088 (N_6088,N_1323,N_934);
nor U6089 (N_6089,N_3550,N_2854);
or U6090 (N_6090,N_2452,N_1630);
or U6091 (N_6091,N_3744,N_809);
nand U6092 (N_6092,N_4525,N_4773);
nor U6093 (N_6093,N_1419,N_2484);
and U6094 (N_6094,N_1795,N_1583);
and U6095 (N_6095,N_3828,N_2350);
and U6096 (N_6096,N_3202,N_470);
or U6097 (N_6097,N_1920,N_4107);
nor U6098 (N_6098,N_1886,N_622);
nand U6099 (N_6099,N_2141,N_2887);
nand U6100 (N_6100,N_507,N_879);
and U6101 (N_6101,N_4344,N_2714);
and U6102 (N_6102,N_582,N_1581);
nor U6103 (N_6103,N_4400,N_3391);
or U6104 (N_6104,N_3394,N_2780);
nand U6105 (N_6105,N_4194,N_2148);
or U6106 (N_6106,N_1675,N_1643);
xor U6107 (N_6107,N_2679,N_2471);
nand U6108 (N_6108,N_4713,N_3161);
nor U6109 (N_6109,N_4589,N_4039);
and U6110 (N_6110,N_4690,N_3844);
or U6111 (N_6111,N_3361,N_4720);
nand U6112 (N_6112,N_3320,N_4377);
nand U6113 (N_6113,N_4643,N_1481);
and U6114 (N_6114,N_3457,N_3483);
and U6115 (N_6115,N_4414,N_943);
and U6116 (N_6116,N_2395,N_1515);
and U6117 (N_6117,N_2654,N_202);
nand U6118 (N_6118,N_2131,N_4181);
nor U6119 (N_6119,N_2695,N_4586);
xor U6120 (N_6120,N_810,N_4144);
nand U6121 (N_6121,N_1766,N_1689);
nand U6122 (N_6122,N_1154,N_1426);
nor U6123 (N_6123,N_1128,N_3478);
or U6124 (N_6124,N_1413,N_2017);
and U6125 (N_6125,N_3270,N_3289);
nand U6126 (N_6126,N_3434,N_708);
and U6127 (N_6127,N_2144,N_3926);
and U6128 (N_6128,N_1487,N_3435);
xnor U6129 (N_6129,N_4074,N_3964);
or U6130 (N_6130,N_1803,N_3873);
and U6131 (N_6131,N_4234,N_4634);
or U6132 (N_6132,N_1524,N_1277);
and U6133 (N_6133,N_2740,N_193);
xnor U6134 (N_6134,N_2564,N_2652);
nor U6135 (N_6135,N_1566,N_1669);
xor U6136 (N_6136,N_3363,N_3821);
nand U6137 (N_6137,N_2125,N_3634);
nor U6138 (N_6138,N_4410,N_4654);
and U6139 (N_6139,N_3888,N_1635);
xnor U6140 (N_6140,N_4490,N_2321);
nand U6141 (N_6141,N_1274,N_4092);
or U6142 (N_6142,N_4126,N_3993);
and U6143 (N_6143,N_268,N_3405);
nor U6144 (N_6144,N_321,N_1111);
and U6145 (N_6145,N_3513,N_2731);
nand U6146 (N_6146,N_1212,N_1039);
nor U6147 (N_6147,N_653,N_4311);
nor U6148 (N_6148,N_4482,N_2824);
nand U6149 (N_6149,N_1509,N_2033);
nor U6150 (N_6150,N_1665,N_500);
or U6151 (N_6151,N_4494,N_12);
or U6152 (N_6152,N_3044,N_563);
nand U6153 (N_6153,N_546,N_56);
nand U6154 (N_6154,N_4180,N_2088);
nand U6155 (N_6155,N_1554,N_4406);
and U6156 (N_6156,N_4968,N_1778);
or U6157 (N_6157,N_501,N_2006);
nor U6158 (N_6158,N_3701,N_1224);
nor U6159 (N_6159,N_2495,N_263);
nand U6160 (N_6160,N_60,N_1463);
and U6161 (N_6161,N_3373,N_3581);
and U6162 (N_6162,N_3466,N_1234);
or U6163 (N_6163,N_1346,N_1024);
and U6164 (N_6164,N_2594,N_2624);
and U6165 (N_6165,N_2118,N_727);
or U6166 (N_6166,N_1575,N_2366);
or U6167 (N_6167,N_164,N_2005);
nor U6168 (N_6168,N_781,N_3041);
nand U6169 (N_6169,N_2201,N_2147);
xnor U6170 (N_6170,N_1119,N_2402);
and U6171 (N_6171,N_970,N_1927);
and U6172 (N_6172,N_4793,N_334);
or U6173 (N_6173,N_4426,N_2439);
nor U6174 (N_6174,N_3049,N_278);
and U6175 (N_6175,N_1502,N_1171);
nor U6176 (N_6176,N_4480,N_649);
xor U6177 (N_6177,N_4375,N_2023);
and U6178 (N_6178,N_4109,N_1634);
nand U6179 (N_6179,N_1312,N_1217);
xnor U6180 (N_6180,N_4629,N_624);
nor U6181 (N_6181,N_1565,N_1309);
xor U6182 (N_6182,N_4646,N_2777);
xnor U6183 (N_6183,N_1082,N_2965);
nand U6184 (N_6184,N_2529,N_2632);
nor U6185 (N_6185,N_979,N_1703);
nand U6186 (N_6186,N_1167,N_2785);
xor U6187 (N_6187,N_4826,N_4854);
or U6188 (N_6188,N_2057,N_177);
and U6189 (N_6189,N_3200,N_4947);
and U6190 (N_6190,N_2884,N_2664);
and U6191 (N_6191,N_3110,N_2468);
xor U6192 (N_6192,N_4516,N_1538);
nand U6193 (N_6193,N_2301,N_2986);
or U6194 (N_6194,N_4688,N_4889);
or U6195 (N_6195,N_4694,N_3111);
and U6196 (N_6196,N_3938,N_1002);
nand U6197 (N_6197,N_4780,N_3973);
and U6198 (N_6198,N_3493,N_2343);
and U6199 (N_6199,N_196,N_4208);
nand U6200 (N_6200,N_4136,N_1492);
nor U6201 (N_6201,N_1282,N_2865);
nor U6202 (N_6202,N_1220,N_4754);
or U6203 (N_6203,N_4834,N_933);
or U6204 (N_6204,N_4651,N_1587);
and U6205 (N_6205,N_2365,N_1504);
nand U6206 (N_6206,N_1010,N_1793);
and U6207 (N_6207,N_2481,N_2724);
nor U6208 (N_6208,N_4440,N_2049);
or U6209 (N_6209,N_3552,N_1080);
nor U6210 (N_6210,N_3622,N_4768);
nor U6211 (N_6211,N_870,N_3312);
and U6212 (N_6212,N_106,N_4295);
nor U6213 (N_6213,N_669,N_4085);
nand U6214 (N_6214,N_3298,N_1911);
nand U6215 (N_6215,N_2567,N_719);
or U6216 (N_6216,N_3987,N_551);
and U6217 (N_6217,N_3521,N_2550);
nand U6218 (N_6218,N_3406,N_2107);
nand U6219 (N_6219,N_2852,N_865);
nor U6220 (N_6220,N_3264,N_2442);
and U6221 (N_6221,N_3989,N_3047);
and U6222 (N_6222,N_1805,N_1995);
nor U6223 (N_6223,N_3336,N_77);
xnor U6224 (N_6224,N_286,N_1505);
and U6225 (N_6225,N_1991,N_3909);
nor U6226 (N_6226,N_2821,N_2491);
and U6227 (N_6227,N_2683,N_3408);
and U6228 (N_6228,N_2955,N_4867);
nand U6229 (N_6229,N_2850,N_3162);
or U6230 (N_6230,N_960,N_1946);
or U6231 (N_6231,N_2226,N_732);
or U6232 (N_6232,N_3211,N_2346);
nor U6233 (N_6233,N_2961,N_2776);
xor U6234 (N_6234,N_1133,N_539);
and U6235 (N_6235,N_265,N_292);
nand U6236 (N_6236,N_4291,N_2681);
nand U6237 (N_6237,N_3009,N_967);
or U6238 (N_6238,N_3067,N_3348);
or U6239 (N_6239,N_1226,N_904);
and U6240 (N_6240,N_3823,N_1174);
and U6241 (N_6241,N_655,N_4946);
nor U6242 (N_6242,N_1574,N_3747);
nor U6243 (N_6243,N_183,N_2913);
and U6244 (N_6244,N_668,N_2016);
and U6245 (N_6245,N_4257,N_3379);
or U6246 (N_6246,N_1343,N_3905);
or U6247 (N_6247,N_2398,N_2767);
nand U6248 (N_6248,N_2252,N_2554);
xnor U6249 (N_6249,N_2061,N_168);
and U6250 (N_6250,N_1710,N_3863);
xnor U6251 (N_6251,N_4373,N_3397);
or U6252 (N_6252,N_3908,N_3503);
and U6253 (N_6253,N_3463,N_1195);
nor U6254 (N_6254,N_2445,N_2110);
or U6255 (N_6255,N_1320,N_3984);
or U6256 (N_6256,N_4301,N_1953);
and U6257 (N_6257,N_1604,N_4839);
nor U6258 (N_6258,N_4943,N_725);
nand U6259 (N_6259,N_3297,N_1818);
nor U6260 (N_6260,N_1658,N_2020);
nor U6261 (N_6261,N_1868,N_3832);
or U6262 (N_6262,N_2362,N_2917);
or U6263 (N_6263,N_59,N_840);
and U6264 (N_6264,N_4462,N_2332);
or U6265 (N_6265,N_2257,N_3659);
nor U6266 (N_6266,N_1825,N_3099);
and U6267 (N_6267,N_2949,N_409);
and U6268 (N_6268,N_1132,N_4972);
xnor U6269 (N_6269,N_4247,N_3776);
and U6270 (N_6270,N_2655,N_4537);
and U6271 (N_6271,N_674,N_932);
nand U6272 (N_6272,N_4661,N_130);
and U6273 (N_6273,N_4466,N_3344);
nand U6274 (N_6274,N_3914,N_2077);
xnor U6275 (N_6275,N_829,N_4117);
nor U6276 (N_6276,N_983,N_2292);
and U6277 (N_6277,N_1705,N_4041);
nand U6278 (N_6278,N_1974,N_2161);
nor U6279 (N_6279,N_869,N_682);
nand U6280 (N_6280,N_2218,N_1339);
and U6281 (N_6281,N_422,N_1961);
xnor U6282 (N_6282,N_184,N_1045);
nand U6283 (N_6283,N_2831,N_1940);
xor U6284 (N_6284,N_4238,N_4094);
nor U6285 (N_6285,N_3094,N_2093);
or U6286 (N_6286,N_935,N_113);
nand U6287 (N_6287,N_1706,N_2588);
or U6288 (N_6288,N_4023,N_4676);
or U6289 (N_6289,N_3957,N_4805);
and U6290 (N_6290,N_1022,N_2788);
nor U6291 (N_6291,N_745,N_4362);
xnor U6292 (N_6292,N_2319,N_4384);
and U6293 (N_6293,N_713,N_281);
xor U6294 (N_6294,N_1105,N_1061);
and U6295 (N_6295,N_2079,N_1586);
nand U6296 (N_6296,N_99,N_3934);
nand U6297 (N_6297,N_924,N_4304);
nand U6298 (N_6298,N_4803,N_2193);
or U6299 (N_6299,N_3347,N_2586);
nand U6300 (N_6300,N_4962,N_3308);
or U6301 (N_6301,N_1731,N_4701);
nor U6302 (N_6302,N_1965,N_2569);
or U6303 (N_6303,N_3721,N_2999);
nand U6304 (N_6304,N_4343,N_4162);
nor U6305 (N_6305,N_4515,N_2702);
or U6306 (N_6306,N_4791,N_3199);
xnor U6307 (N_6307,N_233,N_1488);
nand U6308 (N_6308,N_48,N_4250);
xor U6309 (N_6309,N_1719,N_4073);
or U6310 (N_6310,N_1558,N_71);
nor U6311 (N_6311,N_1787,N_204);
nor U6312 (N_6312,N_1539,N_3164);
or U6313 (N_6313,N_656,N_1971);
nor U6314 (N_6314,N_4808,N_1321);
or U6315 (N_6315,N_3318,N_1579);
nor U6316 (N_6316,N_4289,N_568);
nand U6317 (N_6317,N_3849,N_1044);
nor U6318 (N_6318,N_4799,N_3079);
nor U6319 (N_6319,N_4737,N_2380);
nor U6320 (N_6320,N_350,N_2836);
nor U6321 (N_6321,N_1390,N_2818);
or U6322 (N_6322,N_1990,N_2296);
nor U6323 (N_6323,N_2960,N_2966);
nand U6324 (N_6324,N_1804,N_1396);
nand U6325 (N_6325,N_2752,N_1708);
nor U6326 (N_6326,N_3990,N_2098);
nand U6327 (N_6327,N_531,N_3644);
xor U6328 (N_6328,N_1799,N_3799);
or U6329 (N_6329,N_19,N_228);
nand U6330 (N_6330,N_2646,N_1183);
nand U6331 (N_6331,N_3166,N_4124);
and U6332 (N_6332,N_2590,N_424);
nor U6333 (N_6333,N_1607,N_4084);
or U6334 (N_6334,N_2230,N_2381);
xnor U6335 (N_6335,N_509,N_1763);
or U6336 (N_6336,N_4303,N_3061);
nand U6337 (N_6337,N_4058,N_4554);
nand U6338 (N_6338,N_2387,N_705);
or U6339 (N_6339,N_4999,N_1654);
nor U6340 (N_6340,N_2717,N_137);
nand U6341 (N_6341,N_1194,N_3514);
nand U6342 (N_6342,N_4583,N_4730);
nand U6343 (N_6343,N_3723,N_4123);
or U6344 (N_6344,N_4457,N_3000);
or U6345 (N_6345,N_3204,N_3105);
nand U6346 (N_6346,N_1293,N_760);
nor U6347 (N_6347,N_293,N_1041);
and U6348 (N_6348,N_4040,N_4917);
and U6349 (N_6349,N_449,N_4270);
nor U6350 (N_6350,N_3881,N_4505);
nand U6351 (N_6351,N_4677,N_2485);
nor U6352 (N_6352,N_1311,N_3711);
nor U6353 (N_6353,N_3462,N_4267);
xnor U6354 (N_6354,N_1864,N_2195);
or U6355 (N_6355,N_3481,N_1202);
or U6356 (N_6356,N_4851,N_487);
or U6357 (N_6357,N_4264,N_919);
nand U6358 (N_6358,N_4985,N_1888);
nor U6359 (N_6359,N_1967,N_3868);
nand U6360 (N_6360,N_2396,N_1593);
nand U6361 (N_6361,N_2096,N_4631);
or U6362 (N_6362,N_3725,N_3692);
nand U6363 (N_6363,N_2373,N_1810);
and U6364 (N_6364,N_2779,N_4573);
nand U6365 (N_6365,N_4485,N_2845);
nor U6366 (N_6366,N_3057,N_3108);
and U6367 (N_6367,N_1870,N_1714);
or U6368 (N_6368,N_1796,N_2704);
xnor U6369 (N_6369,N_2763,N_4833);
nor U6370 (N_6370,N_3122,N_937);
and U6371 (N_6371,N_4744,N_3271);
nand U6372 (N_6372,N_1854,N_1379);
nand U6373 (N_6373,N_1478,N_4623);
and U6374 (N_6374,N_1790,N_4443);
or U6375 (N_6375,N_4382,N_931);
or U6376 (N_6376,N_308,N_1933);
nand U6377 (N_6377,N_3265,N_4534);
or U6378 (N_6378,N_4549,N_2733);
or U6379 (N_6379,N_3154,N_4561);
and U6380 (N_6380,N_4342,N_1616);
or U6381 (N_6381,N_2837,N_2872);
nand U6382 (N_6382,N_2032,N_3293);
and U6383 (N_6383,N_4648,N_4184);
or U6384 (N_6384,N_3840,N_64);
or U6385 (N_6385,N_1480,N_1221);
or U6386 (N_6386,N_3928,N_2192);
and U6387 (N_6387,N_2003,N_999);
nand U6388 (N_6388,N_3920,N_398);
or U6389 (N_6389,N_4125,N_3024);
nand U6390 (N_6390,N_3287,N_3069);
and U6391 (N_6391,N_3413,N_2423);
and U6392 (N_6392,N_4811,N_4704);
and U6393 (N_6393,N_1599,N_4268);
xor U6394 (N_6394,N_2121,N_1289);
xnor U6395 (N_6395,N_1857,N_4672);
and U6396 (N_6396,N_1114,N_119);
and U6397 (N_6397,N_899,N_833);
nor U6398 (N_6398,N_1506,N_4502);
and U6399 (N_6399,N_3401,N_3590);
nand U6400 (N_6400,N_1546,N_4702);
nand U6401 (N_6401,N_3753,N_1100);
and U6402 (N_6402,N_332,N_954);
and U6403 (N_6403,N_2372,N_1383);
and U6404 (N_6404,N_241,N_490);
or U6405 (N_6405,N_29,N_1186);
and U6406 (N_6406,N_1584,N_3109);
nor U6407 (N_6407,N_3705,N_2756);
and U6408 (N_6408,N_3095,N_3525);
nor U6409 (N_6409,N_23,N_1416);
nor U6410 (N_6410,N_3575,N_1085);
nand U6411 (N_6411,N_1067,N_2694);
and U6412 (N_6412,N_938,N_4900);
and U6413 (N_6413,N_1040,N_3953);
or U6414 (N_6414,N_1098,N_2473);
nand U6415 (N_6415,N_2353,N_1280);
xnor U6416 (N_6416,N_2408,N_1284);
and U6417 (N_6417,N_4545,N_2910);
nand U6418 (N_6418,N_618,N_4969);
xor U6419 (N_6419,N_764,N_613);
or U6420 (N_6420,N_3410,N_4945);
nand U6421 (N_6421,N_4774,N_1249);
nand U6422 (N_6422,N_2435,N_4650);
and U6423 (N_6423,N_363,N_2432);
nand U6424 (N_6424,N_3544,N_3609);
nand U6425 (N_6425,N_389,N_3730);
nor U6426 (N_6426,N_4195,N_1027);
or U6427 (N_6427,N_4929,N_1844);
and U6428 (N_6428,N_2663,N_939);
nor U6429 (N_6429,N_373,N_1334);
nor U6430 (N_6430,N_459,N_667);
xor U6431 (N_6431,N_475,N_3693);
nor U6432 (N_6432,N_1657,N_567);
nor U6433 (N_6433,N_4141,N_2527);
or U6434 (N_6434,N_4461,N_3407);
or U6435 (N_6435,N_2976,N_218);
nand U6436 (N_6436,N_3985,N_2080);
and U6437 (N_6437,N_1270,N_1957);
or U6438 (N_6438,N_2048,N_4067);
xnor U6439 (N_6439,N_525,N_687);
or U6440 (N_6440,N_4675,N_4961);
and U6441 (N_6441,N_2905,N_4950);
or U6442 (N_6442,N_2627,N_1018);
nand U6443 (N_6443,N_3576,N_1845);
or U6444 (N_6444,N_1292,N_3891);
and U6445 (N_6445,N_1837,N_2720);
nand U6446 (N_6446,N_3432,N_290);
or U6447 (N_6447,N_4223,N_2288);
or U6448 (N_6448,N_4498,N_734);
nor U6449 (N_6449,N_3011,N_929);
nand U6450 (N_6450,N_886,N_3438);
or U6451 (N_6451,N_1653,N_256);
or U6452 (N_6452,N_2208,N_3658);
or U6453 (N_6453,N_3923,N_2055);
xnor U6454 (N_6454,N_1365,N_3458);
nor U6455 (N_6455,N_2803,N_4464);
xnor U6456 (N_6456,N_4127,N_3570);
nor U6457 (N_6457,N_1738,N_4912);
or U6458 (N_6458,N_1493,N_2225);
and U6459 (N_6459,N_2555,N_1883);
nand U6460 (N_6460,N_1850,N_2915);
nor U6461 (N_6461,N_1682,N_4707);
xnor U6462 (N_6462,N_325,N_1485);
or U6463 (N_6463,N_4249,N_2768);
or U6464 (N_6464,N_648,N_528);
nand U6465 (N_6465,N_2571,N_3696);
nor U6466 (N_6466,N_4043,N_3560);
nor U6467 (N_6467,N_1033,N_17);
xor U6468 (N_6468,N_2182,N_1404);
nor U6469 (N_6469,N_3853,N_1017);
nor U6470 (N_6470,N_4581,N_3616);
or U6471 (N_6471,N_3141,N_3443);
nand U6472 (N_6472,N_3449,N_3767);
xnor U6473 (N_6473,N_4367,N_1187);
or U6474 (N_6474,N_4038,N_4469);
xor U6475 (N_6475,N_695,N_3841);
nor U6476 (N_6476,N_3599,N_2787);
and U6477 (N_6477,N_2298,N_298);
or U6478 (N_6478,N_3248,N_2607);
and U6479 (N_6479,N_299,N_3001);
xor U6480 (N_6480,N_2066,N_3422);
and U6481 (N_6481,N_671,N_397);
nand U6482 (N_6482,N_1997,N_4404);
nand U6483 (N_6483,N_3355,N_2911);
or U6484 (N_6484,N_128,N_1798);
or U6485 (N_6485,N_4447,N_1160);
nand U6486 (N_6486,N_673,N_3945);
nand U6487 (N_6487,N_1897,N_2863);
nand U6488 (N_6488,N_2076,N_3020);
nor U6489 (N_6489,N_2231,N_3688);
nand U6490 (N_6490,N_2256,N_3021);
and U6491 (N_6491,N_1724,N_4302);
and U6492 (N_6492,N_4214,N_629);
nor U6493 (N_6493,N_445,N_1245);
and U6494 (N_6494,N_4822,N_859);
nor U6495 (N_6495,N_1594,N_646);
or U6496 (N_6496,N_2606,N_1421);
and U6497 (N_6497,N_461,N_3654);
nor U6498 (N_6498,N_1519,N_2605);
and U6499 (N_6499,N_3101,N_640);
nor U6500 (N_6500,N_3922,N_4287);
nor U6501 (N_6501,N_1813,N_2944);
nor U6502 (N_6502,N_232,N_2953);
or U6503 (N_6503,N_4725,N_2008);
or U6504 (N_6504,N_3050,N_773);
nor U6505 (N_6505,N_1935,N_3940);
xor U6506 (N_6506,N_253,N_2892);
nand U6507 (N_6507,N_4954,N_1267);
xor U6508 (N_6508,N_1923,N_3955);
nand U6509 (N_6509,N_2839,N_4574);
or U6510 (N_6510,N_2267,N_1821);
and U6511 (N_6511,N_2754,N_3892);
or U6512 (N_6512,N_2459,N_4899);
nor U6513 (N_6513,N_2097,N_4435);
and U6514 (N_6514,N_4359,N_817);
nand U6515 (N_6515,N_2204,N_4928);
and U6516 (N_6516,N_675,N_4408);
or U6517 (N_6517,N_1833,N_3152);
or U6518 (N_6518,N_3499,N_639);
nand U6519 (N_6519,N_3381,N_2220);
nor U6520 (N_6520,N_3125,N_86);
nand U6521 (N_6521,N_4856,N_2553);
and U6522 (N_6522,N_3495,N_1570);
and U6523 (N_6523,N_4363,N_1057);
or U6524 (N_6524,N_3589,N_3588);
nand U6525 (N_6525,N_3831,N_4370);
and U6526 (N_6526,N_1460,N_1874);
or U6527 (N_6527,N_4369,N_3870);
and U6528 (N_6528,N_766,N_4216);
nand U6529 (N_6529,N_185,N_3950);
nor U6530 (N_6530,N_3746,N_4819);
nand U6531 (N_6531,N_1758,N_2476);
or U6532 (N_6532,N_3878,N_2690);
nand U6533 (N_6533,N_14,N_3754);
or U6534 (N_6534,N_587,N_1257);
and U6535 (N_6535,N_2834,N_3986);
nor U6536 (N_6536,N_3027,N_3790);
nand U6537 (N_6537,N_3417,N_3193);
or U6538 (N_6538,N_2622,N_1265);
nand U6539 (N_6539,N_1973,N_854);
xnor U6540 (N_6540,N_1503,N_701);
and U6541 (N_6541,N_4571,N_4740);
nand U6542 (N_6542,N_3234,N_526);
nand U6543 (N_6543,N_890,N_858);
or U6544 (N_6544,N_4417,N_1791);
nand U6545 (N_6545,N_4451,N_3810);
xor U6546 (N_6546,N_3707,N_3269);
and U6547 (N_6547,N_143,N_1436);
nor U6548 (N_6548,N_1007,N_2513);
and U6549 (N_6549,N_4193,N_3768);
and U6550 (N_6550,N_2406,N_83);
and U6551 (N_6551,N_4721,N_914);
nand U6552 (N_6552,N_1216,N_1472);
nor U6553 (N_6553,N_3103,N_4004);
or U6554 (N_6554,N_90,N_1250);
nor U6555 (N_6555,N_4346,N_4112);
or U6556 (N_6556,N_3607,N_2299);
nand U6557 (N_6557,N_4495,N_4089);
nor U6558 (N_6558,N_4448,N_3569);
nor U6559 (N_6559,N_1223,N_3774);
and U6560 (N_6560,N_3172,N_118);
and U6561 (N_6561,N_2167,N_460);
or U6562 (N_6562,N_2264,N_3446);
or U6563 (N_6563,N_850,N_1880);
nor U6564 (N_6564,N_4882,N_153);
nor U6565 (N_6565,N_3839,N_74);
or U6566 (N_6566,N_1545,N_3411);
or U6567 (N_6567,N_4314,N_3040);
xnor U6568 (N_6568,N_3919,N_4812);
and U6569 (N_6569,N_2708,N_3088);
or U6570 (N_6570,N_2549,N_3104);
or U6571 (N_6571,N_2692,N_4322);
or U6572 (N_6572,N_2305,N_4275);
or U6573 (N_6573,N_2082,N_2711);
nor U6574 (N_6574,N_3943,N_2019);
or U6575 (N_6575,N_818,N_155);
xnor U6576 (N_6576,N_756,N_4902);
nor U6577 (N_6577,N_219,N_1389);
or U6578 (N_6578,N_3419,N_4324);
or U6579 (N_6579,N_726,N_4855);
nor U6580 (N_6580,N_4548,N_1372);
or U6581 (N_6581,N_2116,N_3322);
nor U6582 (N_6582,N_3585,N_4880);
xnor U6583 (N_6583,N_2067,N_1755);
and U6584 (N_6584,N_2478,N_390);
nor U6585 (N_6585,N_1097,N_4059);
nand U6586 (N_6586,N_4691,N_3935);
xnor U6587 (N_6587,N_1942,N_3062);
or U6588 (N_6588,N_2123,N_388);
and U6589 (N_6589,N_4349,N_2833);
nor U6590 (N_6590,N_319,N_4746);
and U6591 (N_6591,N_1527,N_752);
nor U6592 (N_6592,N_176,N_1015);
nor U6593 (N_6593,N_3315,N_4503);
nand U6594 (N_6594,N_4992,N_3530);
and U6595 (N_6595,N_4680,N_4076);
nand U6596 (N_6596,N_1102,N_4356);
xnor U6597 (N_6597,N_407,N_710);
nor U6598 (N_6598,N_2180,N_2351);
nor U6599 (N_6599,N_415,N_3951);
nand U6600 (N_6600,N_1585,N_4817);
nor U6601 (N_6601,N_963,N_4527);
nand U6602 (N_6602,N_4389,N_4159);
nand U6603 (N_6603,N_6,N_488);
xnor U6604 (N_6604,N_4767,N_1337);
nand U6605 (N_6605,N_722,N_1520);
nor U6606 (N_6606,N_4235,N_2729);
xor U6607 (N_6607,N_2246,N_4215);
nand U6608 (N_6608,N_3562,N_2723);
nand U6609 (N_6609,N_1895,N_25);
or U6610 (N_6610,N_4305,N_238);
or U6611 (N_6611,N_1401,N_3331);
nand U6612 (N_6612,N_4042,N_243);
nor U6613 (N_6613,N_203,N_3862);
nand U6614 (N_6614,N_628,N_4695);
and U6615 (N_6615,N_2943,N_2532);
and U6616 (N_6616,N_2541,N_1268);
nand U6617 (N_6617,N_471,N_1691);
nor U6618 (N_6618,N_751,N_2268);
nand U6619 (N_6619,N_338,N_4407);
nor U6620 (N_6620,N_2736,N_2812);
nand U6621 (N_6621,N_2114,N_2985);
nor U6622 (N_6622,N_728,N_1192);
and U6623 (N_6623,N_2451,N_54);
nor U6624 (N_6624,N_251,N_58);
or U6625 (N_6625,N_1771,N_2239);
nand U6626 (N_6626,N_2330,N_451);
nor U6627 (N_6627,N_4008,N_418);
nor U6628 (N_6628,N_2229,N_2216);
nand U6629 (N_6629,N_180,N_260);
xnor U6630 (N_6630,N_632,N_3314);
and U6631 (N_6631,N_918,N_2002);
nand U6632 (N_6632,N_3023,N_3718);
nor U6633 (N_6633,N_542,N_2737);
nand U6634 (N_6634,N_1996,N_1235);
nor U6635 (N_6635,N_884,N_3545);
nor U6636 (N_6636,N_2829,N_1092);
nor U6637 (N_6637,N_2738,N_1836);
or U6638 (N_6638,N_3416,N_1521);
and U6639 (N_6639,N_1684,N_3294);
nor U6640 (N_6640,N_1622,N_3471);
or U6641 (N_6641,N_862,N_4976);
or U6642 (N_6642,N_3309,N_1447);
or U6643 (N_6643,N_4655,N_4590);
xor U6644 (N_6644,N_3651,N_1400);
nand U6645 (N_6645,N_2163,N_3135);
or U6646 (N_6646,N_2972,N_1214);
nand U6647 (N_6647,N_1175,N_1672);
or U6648 (N_6648,N_432,N_141);
xnor U6649 (N_6649,N_2579,N_1964);
and U6650 (N_6650,N_3165,N_4806);
nor U6651 (N_6651,N_2414,N_643);
nor U6652 (N_6652,N_3465,N_3772);
nand U6653 (N_6653,N_189,N_79);
or U6654 (N_6654,N_4146,N_644);
and U6655 (N_6655,N_3276,N_2902);
nor U6656 (N_6656,N_2642,N_98);
nor U6657 (N_6657,N_112,N_462);
nor U6658 (N_6658,N_3427,N_4895);
nand U6659 (N_6659,N_3182,N_3257);
nand U6660 (N_6660,N_2709,N_3078);
nand U6661 (N_6661,N_2503,N_3025);
nor U6662 (N_6662,N_2224,N_138);
and U6663 (N_6663,N_3847,N_4148);
nor U6664 (N_6664,N_2113,N_4765);
xor U6665 (N_6665,N_936,N_4425);
nand U6666 (N_6666,N_690,N_376);
and U6667 (N_6667,N_4732,N_603);
or U6668 (N_6668,N_4009,N_4852);
nor U6669 (N_6669,N_504,N_3628);
nand U6670 (N_6670,N_1986,N_4575);
and U6671 (N_6671,N_3534,N_2580);
or U6672 (N_6672,N_3969,N_3736);
or U6673 (N_6673,N_1153,N_186);
nand U6674 (N_6674,N_1696,N_578);
and U6675 (N_6675,N_1770,N_836);
nand U6676 (N_6676,N_2744,N_150);
nor U6677 (N_6677,N_1733,N_2438);
or U6678 (N_6678,N_3085,N_4922);
nor U6679 (N_6679,N_4151,N_4958);
xor U6680 (N_6680,N_3983,N_1125);
xnor U6681 (N_6681,N_1134,N_3978);
xnor U6682 (N_6682,N_497,N_1939);
and U6683 (N_6683,N_3292,N_4005);
nand U6684 (N_6684,N_414,N_2339);
xnor U6685 (N_6685,N_294,N_2545);
and U6686 (N_6686,N_1169,N_2531);
nand U6687 (N_6687,N_2919,N_2054);
nand U6688 (N_6688,N_4700,N_3096);
nand U6689 (N_6689,N_4628,N_3268);
nand U6690 (N_6690,N_3582,N_1668);
nor U6691 (N_6691,N_1721,N_864);
and U6692 (N_6692,N_4564,N_1363);
and U6693 (N_6693,N_4908,N_4266);
or U6694 (N_6694,N_2800,N_267);
xnor U6695 (N_6695,N_2848,N_4610);
or U6696 (N_6696,N_4823,N_2287);
or U6697 (N_6697,N_4959,N_1101);
or U6698 (N_6698,N_1910,N_3806);
nand U6699 (N_6699,N_2378,N_1591);
nor U6700 (N_6700,N_2431,N_874);
xnor U6701 (N_6701,N_2209,N_162);
nand U6702 (N_6702,N_3015,N_4183);
and U6703 (N_6703,N_1222,N_1760);
nand U6704 (N_6704,N_456,N_3592);
nor U6705 (N_6705,N_400,N_1863);
or U6706 (N_6706,N_3272,N_4104);
or U6707 (N_6707,N_4213,N_4953);
nor U6708 (N_6708,N_2158,N_608);
nand U6709 (N_6709,N_4240,N_958);
or U6710 (N_6710,N_3875,N_3981);
or U6711 (N_6711,N_3837,N_3682);
nand U6712 (N_6712,N_2479,N_341);
and U6713 (N_6713,N_2065,N_1613);
or U6714 (N_6714,N_4108,N_4309);
nand U6715 (N_6715,N_1945,N_962);
and U6716 (N_6716,N_2175,N_4572);
nand U6717 (N_6717,N_1326,N_4507);
or U6718 (N_6718,N_2397,N_3686);
xnor U6719 (N_6719,N_4597,N_888);
or U6720 (N_6720,N_4364,N_2105);
nand U6721 (N_6721,N_3380,N_2419);
and U6722 (N_6722,N_1140,N_3016);
nand U6723 (N_6723,N_776,N_729);
nand U6724 (N_6724,N_4329,N_3281);
xor U6725 (N_6725,N_361,N_4071);
or U6726 (N_6726,N_3655,N_1998);
nor U6727 (N_6727,N_3424,N_3678);
nor U6728 (N_6728,N_4261,N_4053);
or U6729 (N_6729,N_1784,N_4278);
nand U6730 (N_6730,N_3354,N_1849);
and U6731 (N_6731,N_1702,N_4506);
or U6732 (N_6732,N_3907,N_1068);
and U6733 (N_6733,N_1332,N_3176);
nand U6734 (N_6734,N_1716,N_3382);
and U6735 (N_6735,N_3387,N_4603);
or U6736 (N_6736,N_2760,N_489);
or U6737 (N_6737,N_3139,N_3879);
and U6738 (N_6738,N_3506,N_4357);
nand U6739 (N_6739,N_3770,N_4872);
and U6740 (N_6740,N_156,N_1123);
and U6741 (N_6741,N_1036,N_4762);
nor U6742 (N_6742,N_423,N_700);
or U6743 (N_6743,N_2200,N_142);
nor U6744 (N_6744,N_1614,N_2741);
nand U6745 (N_6745,N_2369,N_2750);
nand U6746 (N_6746,N_3739,N_2086);
xor U6747 (N_6747,N_2667,N_3045);
or U6748 (N_6748,N_2492,N_4176);
and U6749 (N_6749,N_4689,N_3258);
or U6750 (N_6750,N_4083,N_2179);
and U6751 (N_6751,N_992,N_3227);
nor U6752 (N_6752,N_4152,N_62);
nor U6753 (N_6753,N_944,N_4481);
or U6754 (N_6754,N_3856,N_1449);
nor U6755 (N_6755,N_4428,N_2659);
xnor U6756 (N_6756,N_952,N_170);
xnor U6757 (N_6757,N_1260,N_3155);
nor U6758 (N_6758,N_2470,N_4741);
and U6759 (N_6759,N_343,N_1338);
nor U6760 (N_6760,N_4030,N_4990);
nor U6761 (N_6761,N_4891,N_1686);
nand U6762 (N_6762,N_2745,N_1717);
and U6763 (N_6763,N_2151,N_2952);
nand U6764 (N_6764,N_815,N_3647);
and U6765 (N_6765,N_2169,N_519);
nor U6766 (N_6766,N_4599,N_3213);
nor U6767 (N_6767,N_3731,N_2245);
or U6768 (N_6768,N_2383,N_2873);
xnor U6769 (N_6769,N_4050,N_706);
nand U6770 (N_6770,N_427,N_2437);
and U6771 (N_6771,N_3624,N_703);
nor U6772 (N_6772,N_3936,N_788);
or U6773 (N_6773,N_3034,N_905);
nor U6774 (N_6774,N_893,N_2400);
or U6775 (N_6775,N_386,N_2534);
nand U6776 (N_6776,N_1106,N_102);
nand U6777 (N_6777,N_2178,N_4201);
and U6778 (N_6778,N_3572,N_4224);
nor U6779 (N_6779,N_396,N_1304);
or U6780 (N_6780,N_4699,N_4484);
or U6781 (N_6781,N_2456,N_3256);
nor U6782 (N_6782,N_1251,N_2313);
nor U6783 (N_6783,N_2619,N_4622);
and U6784 (N_6784,N_605,N_598);
or U6785 (N_6785,N_4091,N_4420);
nor U6786 (N_6786,N_35,N_4432);
or U6787 (N_6787,N_3554,N_3068);
or U6788 (N_6788,N_1259,N_355);
and U6789 (N_6789,N_1204,N_326);
nor U6790 (N_6790,N_1233,N_2059);
nor U6791 (N_6791,N_635,N_55);
xor U6792 (N_6792,N_2111,N_2551);
and U6793 (N_6793,N_1925,N_2205);
or U6794 (N_6794,N_2759,N_4738);
nand U6795 (N_6795,N_1751,N_1905);
nand U6796 (N_6796,N_3876,N_1178);
or U6797 (N_6797,N_4248,N_2858);
nor U6798 (N_6798,N_2069,N_3487);
and U6799 (N_6799,N_200,N_2979);
nand U6800 (N_6800,N_4149,N_995);
nor U6801 (N_6801,N_2802,N_2609);
nor U6802 (N_6802,N_1822,N_824);
and U6803 (N_6803,N_837,N_894);
nor U6804 (N_6804,N_4840,N_4736);
xnor U6805 (N_6805,N_417,N_4734);
nor U6806 (N_6806,N_1648,N_1514);
or U6807 (N_6807,N_7,N_1075);
nor U6808 (N_6808,N_2347,N_2771);
and U6809 (N_6809,N_3743,N_1609);
or U6810 (N_6810,N_2165,N_493);
nand U6811 (N_6811,N_4637,N_3666);
nor U6812 (N_6812,N_2310,N_2360);
nor U6813 (N_6813,N_4341,N_2126);
and U6814 (N_6814,N_1827,N_1331);
and U6815 (N_6815,N_229,N_681);
xnor U6816 (N_6816,N_3420,N_4752);
and U6817 (N_6817,N_2187,N_3072);
or U6818 (N_6818,N_4167,N_903);
nand U6819 (N_6819,N_357,N_3737);
nor U6820 (N_6820,N_1209,N_2480);
nor U6821 (N_6821,N_116,N_2804);
nor U6822 (N_6822,N_4979,N_4351);
nor U6823 (N_6823,N_3614,N_1759);
nor U6824 (N_6824,N_892,N_3150);
nand U6825 (N_6825,N_820,N_188);
or U6826 (N_6826,N_1016,N_3388);
or U6827 (N_6827,N_2860,N_1417);
or U6828 (N_6828,N_67,N_3680);
or U6829 (N_6829,N_4245,N_561);
nand U6830 (N_6830,N_4365,N_3477);
nor U6831 (N_6831,N_1985,N_4509);
or U6832 (N_6832,N_3174,N_1060);
and U6833 (N_6833,N_2675,N_1091);
or U6834 (N_6834,N_3663,N_4423);
and U6835 (N_6835,N_469,N_1659);
or U6836 (N_6836,N_1215,N_291);
nor U6837 (N_6837,N_4993,N_2648);
or U6838 (N_6838,N_3531,N_3339);
or U6839 (N_6839,N_959,N_1517);
nor U6840 (N_6840,N_1611,N_798);
nor U6841 (N_6841,N_2240,N_1440);
or U6842 (N_6842,N_2796,N_87);
nor U6843 (N_6843,N_4750,N_2117);
nor U6844 (N_6844,N_3184,N_4237);
and U6845 (N_6845,N_1789,N_3698);
nor U6846 (N_6846,N_4253,N_819);
and U6847 (N_6847,N_2703,N_2939);
nor U6848 (N_6848,N_3299,N_3455);
and U6849 (N_6849,N_428,N_1430);
nand U6850 (N_6850,N_2749,N_1801);
and U6851 (N_6851,N_4232,N_4458);
nand U6852 (N_6852,N_3635,N_2676);
and U6853 (N_6853,N_3330,N_1283);
and U6854 (N_6854,N_1612,N_807);
or U6855 (N_6855,N_2375,N_264);
or U6856 (N_6856,N_1264,N_3974);
or U6857 (N_6857,N_3615,N_831);
and U6858 (N_6858,N_2525,N_2658);
nand U6859 (N_6859,N_1079,N_4663);
or U6860 (N_6860,N_2894,N_2672);
nor U6861 (N_6861,N_782,N_2045);
or U6862 (N_6862,N_1308,N_2251);
nand U6863 (N_6863,N_2700,N_3261);
or U6864 (N_6864,N_49,N_3266);
or U6865 (N_6865,N_3674,N_4542);
nor U6866 (N_6866,N_453,N_2255);
nand U6867 (N_6867,N_737,N_3748);
nor U6868 (N_6868,N_448,N_3148);
and U6869 (N_6869,N_242,N_65);
or U6870 (N_6870,N_1779,N_4228);
nand U6871 (N_6871,N_2336,N_1374);
or U6872 (N_6872,N_4933,N_3376);
and U6873 (N_6873,N_1772,N_4477);
and U6874 (N_6874,N_1402,N_1812);
and U6875 (N_6875,N_1375,N_3220);
nor U6876 (N_6876,N_518,N_3735);
and U6877 (N_6877,N_4918,N_2421);
nand U6878 (N_6878,N_3186,N_4319);
and U6879 (N_6879,N_4614,N_4786);
nand U6880 (N_6880,N_4906,N_3988);
and U6881 (N_6881,N_1155,N_3882);
nor U6882 (N_6882,N_1930,N_239);
nor U6883 (N_6883,N_2490,N_3667);
nand U6884 (N_6884,N_4090,N_3901);
xnor U6885 (N_6885,N_4562,N_1152);
nand U6886 (N_6886,N_395,N_4361);
nor U6887 (N_6887,N_1219,N_1988);
or U6888 (N_6888,N_564,N_1381);
nand U6889 (N_6889,N_3490,N_566);
nor U6890 (N_6890,N_4017,N_4775);
and U6891 (N_6891,N_3732,N_4051);
nor U6892 (N_6892,N_1921,N_1376);
or U6893 (N_6893,N_2810,N_3751);
nor U6894 (N_6894,N_3505,N_594);
nand U6895 (N_6895,N_1495,N_1561);
nor U6896 (N_6896,N_4258,N_3812);
nor U6897 (N_6897,N_1341,N_2051);
xnor U6898 (N_6898,N_3752,N_3451);
or U6899 (N_6899,N_1423,N_754);
nor U6900 (N_6900,N_3115,N_1872);
or U6901 (N_6901,N_3633,N_738);
xnor U6902 (N_6902,N_4605,N_3895);
nand U6903 (N_6903,N_650,N_2562);
nand U6904 (N_6904,N_2728,N_3657);
nor U6905 (N_6905,N_1345,N_4529);
nand U6906 (N_6906,N_3602,N_2548);
nand U6907 (N_6907,N_2214,N_680);
nor U6908 (N_6908,N_1161,N_4379);
and U6909 (N_6909,N_1135,N_1177);
or U6910 (N_6910,N_573,N_1972);
and U6911 (N_6911,N_516,N_2157);
nand U6912 (N_6912,N_406,N_4994);
and U6913 (N_6913,N_174,N_3811);
and U6914 (N_6914,N_2640,N_1862);
nor U6915 (N_6915,N_3932,N_2282);
nor U6916 (N_6916,N_443,N_2718);
nor U6917 (N_6917,N_1113,N_309);
nor U6918 (N_6918,N_2320,N_3963);
and U6919 (N_6919,N_3930,N_3741);
and U6920 (N_6920,N_457,N_2326);
or U6921 (N_6921,N_2573,N_2914);
and U6922 (N_6922,N_3807,N_2840);
and U6923 (N_6923,N_2957,N_1838);
nand U6924 (N_6924,N_4664,N_1861);
and U6925 (N_6925,N_1722,N_2784);
or U6926 (N_6926,N_4114,N_2969);
xnor U6927 (N_6927,N_2696,N_3883);
or U6928 (N_6928,N_4120,N_4077);
or U6929 (N_6929,N_1700,N_1300);
or U6930 (N_6930,N_3386,N_3762);
or U6931 (N_6931,N_2458,N_599);
or U6932 (N_6932,N_3510,N_4909);
nor U6933 (N_6933,N_803,N_4975);
or U6934 (N_6934,N_2849,N_3757);
nand U6935 (N_6935,N_4991,N_275);
nand U6936 (N_6936,N_4155,N_1685);
nor U6937 (N_6937,N_1130,N_42);
nor U6938 (N_6938,N_3573,N_252);
or U6939 (N_6939,N_2835,N_1398);
nor U6940 (N_6940,N_1578,N_452);
nor U6941 (N_6941,N_2424,N_4645);
or U6942 (N_6942,N_2616,N_4277);
and U6943 (N_6943,N_3738,N_2235);
or U6944 (N_6944,N_4508,N_3316);
nor U6945 (N_6945,N_804,N_4916);
or U6946 (N_6946,N_377,N_2635);
nand U6947 (N_6947,N_3038,N_834);
xnor U6948 (N_6948,N_3553,N_1048);
nand U6949 (N_6949,N_2950,N_3931);
nand U6950 (N_6950,N_3638,N_772);
nand U6951 (N_6951,N_3356,N_2618);
or U6952 (N_6952,N_3129,N_4029);
nor U6953 (N_6953,N_4097,N_402);
and U6954 (N_6954,N_1553,N_4252);
or U6955 (N_6955,N_830,N_1296);
nor U6956 (N_6956,N_2576,N_1406);
nand U6957 (N_6957,N_2426,N_2464);
and U6958 (N_6958,N_508,N_5);
or U6959 (N_6959,N_2010,N_2819);
xnor U6960 (N_6960,N_2722,N_3352);
nand U6961 (N_6961,N_3064,N_3670);
and U6962 (N_6962,N_1269,N_353);
nor U6963 (N_6963,N_2811,N_479);
nor U6964 (N_6964,N_4259,N_4538);
or U6965 (N_6965,N_1647,N_2210);
and U6966 (N_6966,N_1676,N_2712);
xnor U6967 (N_6967,N_3323,N_996);
nor U6968 (N_6968,N_4135,N_2371);
and U6969 (N_6969,N_1043,N_1547);
nand U6970 (N_6970,N_4901,N_2916);
or U6971 (N_6971,N_1200,N_3824);
or U6972 (N_6972,N_1399,N_2316);
or U6973 (N_6973,N_4578,N_1471);
nor U6974 (N_6974,N_3961,N_4315);
nand U6975 (N_6975,N_2716,N_3872);
and U6976 (N_6976,N_4956,N_2584);
or U6977 (N_6977,N_4965,N_3889);
nor U6978 (N_6978,N_2266,N_545);
nand U6979 (N_6979,N_4412,N_3415);
and U6980 (N_6980,N_4028,N_702);
or U6981 (N_6981,N_1513,N_721);
or U6982 (N_6982,N_1049,N_3147);
nor U6983 (N_6983,N_1618,N_3783);
nor U6984 (N_6984,N_4924,N_1467);
nor U6985 (N_6985,N_439,N_792);
and U6986 (N_6986,N_1013,N_1627);
or U6987 (N_6987,N_340,N_763);
nor U6988 (N_6988,N_4385,N_198);
nor U6989 (N_6989,N_1786,N_1619);
nor U6990 (N_6990,N_4937,N_2623);
nand U6991 (N_6991,N_4535,N_2581);
and U6992 (N_6992,N_348,N_4411);
or U6993 (N_6993,N_739,N_2427);
or U6994 (N_6994,N_2270,N_4419);
or U6995 (N_6995,N_2809,N_1551);
nor U6996 (N_6996,N_2963,N_984);
nand U6997 (N_6997,N_135,N_4242);
nand U6998 (N_6998,N_2924,N_52);
and U6999 (N_6999,N_2612,N_2446);
nand U7000 (N_7000,N_2743,N_3205);
nor U7001 (N_7001,N_4075,N_39);
or U7002 (N_7002,N_1108,N_4739);
nand U7003 (N_7003,N_4514,N_3032);
or U7004 (N_7004,N_3180,N_4288);
and U7005 (N_7005,N_4593,N_4134);
and U7006 (N_7006,N_4859,N_2115);
xor U7007 (N_7007,N_2577,N_4517);
nand U7008 (N_7008,N_2223,N_2029);
nand U7009 (N_7009,N_190,N_696);
or U7010 (N_7010,N_3089,N_3652);
and U7011 (N_7011,N_2127,N_4298);
nor U7012 (N_7012,N_2499,N_1743);
nor U7013 (N_7013,N_4328,N_2666);
nand U7014 (N_7014,N_1828,N_3278);
nand U7015 (N_7015,N_881,N_230);
or U7016 (N_7016,N_3577,N_3902);
and U7017 (N_7017,N_2448,N_3641);
xnor U7018 (N_7018,N_2684,N_2453);
and U7019 (N_7019,N_2794,N_2191);
or U7020 (N_7020,N_4486,N_3369);
nor U7021 (N_7021,N_4512,N_4980);
and U7022 (N_7022,N_3612,N_2781);
nor U7023 (N_7023,N_3091,N_1241);
and U7024 (N_7024,N_53,N_103);
nand U7025 (N_7025,N_2758,N_91);
xnor U7026 (N_7026,N_549,N_3596);
and U7027 (N_7027,N_2429,N_891);
nand U7028 (N_7028,N_2899,N_76);
and U7029 (N_7029,N_4831,N_405);
or U7030 (N_7030,N_2766,N_259);
and U7031 (N_7031,N_379,N_3398);
nor U7032 (N_7032,N_4121,N_1557);
and U7033 (N_7033,N_3046,N_3542);
xnor U7034 (N_7034,N_2483,N_2394);
nor U7035 (N_7035,N_179,N_3128);
nor U7036 (N_7036,N_3903,N_3997);
or U7037 (N_7037,N_2280,N_1511);
or U7038 (N_7038,N_3219,N_3008);
nor U7039 (N_7039,N_4192,N_2232);
and U7040 (N_7040,N_1762,N_3769);
and U7041 (N_7041,N_3910,N_2412);
or U7042 (N_7042,N_3740,N_3845);
nand U7043 (N_7043,N_3671,N_514);
or U7044 (N_7044,N_627,N_3429);
nor U7045 (N_7045,N_1433,N_770);
xnor U7046 (N_7046,N_4579,N_3830);
xor U7047 (N_7047,N_1679,N_4111);
or U7048 (N_7048,N_2420,N_2806);
nor U7049 (N_7049,N_4336,N_3887);
nand U7050 (N_7050,N_2817,N_344);
nand U7051 (N_7051,N_1225,N_1454);
xor U7052 (N_7052,N_4966,N_3781);
or U7053 (N_7053,N_1474,N_111);
or U7054 (N_7054,N_4449,N_2041);
nor U7055 (N_7055,N_4316,N_2132);
nor U7056 (N_7056,N_1646,N_2940);
nand U7057 (N_7057,N_441,N_484);
xor U7058 (N_7058,N_161,N_314);
nand U7059 (N_7059,N_749,N_1892);
or U7060 (N_7060,N_1674,N_208);
nand U7061 (N_7061,N_3187,N_1166);
nor U7062 (N_7062,N_4168,N_1981);
and U7063 (N_7063,N_3608,N_1083);
nand U7064 (N_7064,N_2176,N_4904);
or U7065 (N_7065,N_1734,N_2447);
and U7066 (N_7066,N_2411,N_3826);
nor U7067 (N_7067,N_312,N_1362);
nor U7068 (N_7068,N_4866,N_901);
and U7069 (N_7069,N_2886,N_3586);
nand U7070 (N_7070,N_3237,N_3694);
and U7071 (N_7071,N_4693,N_1273);
and U7072 (N_7072,N_4479,N_2770);
nor U7073 (N_7073,N_2597,N_192);
nand U7074 (N_7074,N_1797,N_131);
nor U7075 (N_7075,N_638,N_2466);
and U7076 (N_7076,N_1136,N_125);
or U7077 (N_7077,N_2890,N_4967);
nor U7078 (N_7078,N_3364,N_1879);
and U7079 (N_7079,N_607,N_1173);
nand U7080 (N_7080,N_4570,N_2367);
nand U7081 (N_7081,N_3733,N_2324);
nand U7082 (N_7082,N_1191,N_2026);
and U7083 (N_7083,N_2691,N_2393);
nand U7084 (N_7084,N_3874,N_1533);
nor U7085 (N_7085,N_4463,N_3683);
or U7086 (N_7086,N_2361,N_4843);
nand U7087 (N_7087,N_4016,N_3194);
and U7088 (N_7088,N_1632,N_3855);
and U7089 (N_7089,N_117,N_412);
and U7090 (N_7090,N_2888,N_3143);
or U7091 (N_7091,N_2071,N_1970);
and U7092 (N_7092,N_699,N_2160);
nor U7093 (N_7093,N_3877,N_2040);
or U7094 (N_7094,N_4832,N_1928);
nand U7095 (N_7095,N_1266,N_4312);
and U7096 (N_7096,N_169,N_3224);
or U7097 (N_7097,N_852,N_3679);
nor U7098 (N_7098,N_2434,N_3390);
xor U7099 (N_7099,N_3700,N_3699);
xnor U7100 (N_7100,N_1723,N_4530);
nor U7101 (N_7101,N_2669,N_1229);
and U7102 (N_7102,N_3675,N_3724);
and U7103 (N_7103,N_1227,N_2904);
and U7104 (N_7104,N_429,N_4372);
or U7105 (N_7105,N_3412,N_3526);
and U7106 (N_7106,N_284,N_1088);
nand U7107 (N_7107,N_4129,N_2520);
and U7108 (N_7108,N_505,N_4156);
or U7109 (N_7109,N_4398,N_2981);
xnor U7110 (N_7110,N_4256,N_579);
or U7111 (N_7111,N_2774,N_324);
nand U7112 (N_7112,N_1009,N_1193);
nand U7113 (N_7113,N_1944,N_3825);
nor U7114 (N_7114,N_3423,N_1667);
nor U7115 (N_7115,N_3795,N_4018);
nor U7116 (N_7116,N_664,N_855);
nor U7117 (N_7117,N_1865,N_4667);
or U7118 (N_7118,N_88,N_1898);
or U7119 (N_7119,N_1867,N_2328);
nor U7120 (N_7120,N_3245,N_997);
nor U7121 (N_7121,N_214,N_4636);
or U7122 (N_7122,N_3342,N_4753);
xor U7123 (N_7123,N_3218,N_1180);
or U7124 (N_7124,N_1846,N_1287);
or U7125 (N_7125,N_4010,N_2560);
nand U7126 (N_7126,N_2311,N_1434);
nor U7127 (N_7127,N_762,N_2073);
and U7128 (N_7128,N_4476,N_4024);
and U7129 (N_7129,N_146,N_4396);
and U7130 (N_7130,N_2506,N_1776);
and U7131 (N_7131,N_4568,N_365);
and U7132 (N_7132,N_1934,N_3966);
or U7133 (N_7133,N_2732,N_712);
nor U7134 (N_7134,N_4459,N_2786);
and U7135 (N_7135,N_2194,N_3175);
and U7136 (N_7136,N_2558,N_2416);
xor U7137 (N_7137,N_1356,N_2869);
nand U7138 (N_7138,N_1692,N_3558);
xor U7139 (N_7139,N_953,N_1452);
nand U7140 (N_7140,N_1752,N_2954);
or U7141 (N_7141,N_957,N_4684);
nand U7142 (N_7142,N_225,N_591);
nor U7143 (N_7143,N_1035,N_96);
or U7144 (N_7144,N_3262,N_270);
nand U7145 (N_7145,N_4221,N_37);
nor U7146 (N_7146,N_1729,N_755);
nand U7147 (N_7147,N_3116,N_2592);
and U7148 (N_7148,N_3275,N_1842);
and U7149 (N_7149,N_3138,N_4788);
or U7150 (N_7150,N_2707,N_2996);
or U7151 (N_7151,N_3469,N_3886);
and U7152 (N_7152,N_1001,N_1298);
and U7153 (N_7153,N_2926,N_1831);
and U7154 (N_7154,N_733,N_1307);
and U7155 (N_7155,N_1237,N_1924);
nor U7156 (N_7156,N_1954,N_3583);
or U7157 (N_7157,N_4153,N_3563);
or U7158 (N_7158,N_4555,N_4132);
nand U7159 (N_7159,N_247,N_3214);
nor U7160 (N_7160,N_3244,N_4838);
and U7161 (N_7161,N_68,N_540);
or U7162 (N_7162,N_3962,N_4971);
and U7163 (N_7163,N_4513,N_2826);
xnor U7164 (N_7164,N_3081,N_3033);
or U7165 (N_7165,N_1640,N_4335);
and U7166 (N_7166,N_3804,N_724);
and U7167 (N_7167,N_920,N_3664);
nand U7168 (N_7168,N_2701,N_4106);
and U7169 (N_7169,N_494,N_645);
nand U7170 (N_7170,N_4064,N_597);
and U7171 (N_7171,N_1902,N_1834);
xnor U7172 (N_7172,N_2636,N_743);
nand U7173 (N_7173,N_4439,N_2706);
or U7174 (N_7174,N_1151,N_1397);
or U7175 (N_7175,N_907,N_283);
or U7176 (N_7176,N_2827,N_965);
nand U7177 (N_7177,N_694,N_502);
nor U7178 (N_7178,N_3716,N_3290);
nor U7179 (N_7179,N_576,N_121);
nor U7180 (N_7180,N_3243,N_3854);
nand U7181 (N_7181,N_4467,N_802);
nor U7182 (N_7182,N_3714,N_3777);
or U7183 (N_7183,N_4620,N_2671);
or U7184 (N_7184,N_3535,N_2524);
nor U7185 (N_7185,N_3814,N_226);
and U7186 (N_7186,N_990,N_1385);
nand U7187 (N_7187,N_4697,N_4175);
nor U7188 (N_7188,N_1617,N_4236);
nor U7189 (N_7189,N_404,N_2649);
nand U7190 (N_7190,N_3515,N_2556);
nand U7191 (N_7191,N_1276,N_194);
nand U7192 (N_7192,N_158,N_1754);
xnor U7193 (N_7193,N_1199,N_4320);
nand U7194 (N_7194,N_1066,N_4794);
nor U7195 (N_7195,N_678,N_4231);
and U7196 (N_7196,N_2699,N_866);
nand U7197 (N_7197,N_3357,N_3475);
nand U7198 (N_7198,N_347,N_1242);
or U7199 (N_7199,N_1435,N_3119);
nand U7200 (N_7200,N_3578,N_2934);
nand U7201 (N_7201,N_4174,N_380);
and U7202 (N_7202,N_4321,N_4229);
and U7203 (N_7203,N_3022,N_3613);
and U7204 (N_7204,N_4845,N_1785);
nand U7205 (N_7205,N_2922,N_2608);
or U7206 (N_7206,N_3643,N_4348);
nor U7207 (N_7207,N_356,N_1620);
nand U7208 (N_7208,N_2410,N_2626);
or U7209 (N_7209,N_3192,N_2515);
nor U7210 (N_7210,N_2084,N_1615);
nor U7211 (N_7211,N_2964,N_3842);
or U7212 (N_7212,N_1158,N_4630);
nor U7213 (N_7213,N_1087,N_1431);
and U7214 (N_7214,N_2050,N_4847);
nand U7215 (N_7215,N_411,N_966);
or U7216 (N_7216,N_2870,N_796);
nor U7217 (N_7217,N_4522,N_4115);
nand U7218 (N_7218,N_4977,N_3992);
nand U7219 (N_7219,N_3673,N_2975);
nand U7220 (N_7220,N_2596,N_2538);
or U7221 (N_7221,N_38,N_280);
or U7222 (N_7222,N_1715,N_2868);
nor U7223 (N_7223,N_104,N_3014);
nor U7224 (N_7224,N_1660,N_4497);
xnor U7225 (N_7225,N_3512,N_1120);
nor U7226 (N_7226,N_255,N_4326);
nand U7227 (N_7227,N_3915,N_4686);
or U7228 (N_7228,N_2001,N_303);
nand U7229 (N_7229,N_4360,N_2660);
or U7230 (N_7230,N_863,N_4188);
nor U7231 (N_7231,N_1074,N_1943);
and U7232 (N_7232,N_3168,N_1461);
and U7233 (N_7233,N_403,N_1535);
and U7234 (N_7234,N_4504,N_4374);
xnor U7235 (N_7235,N_2504,N_4279);
nand U7236 (N_7236,N_2250,N_2101);
or U7237 (N_7237,N_1168,N_2281);
or U7238 (N_7238,N_2645,N_1347);
nand U7239 (N_7239,N_4078,N_1860);
or U7240 (N_7240,N_2544,N_2735);
or U7241 (N_7241,N_3018,N_1835);
or U7242 (N_7242,N_1852,N_2315);
nand U7243 (N_7243,N_4333,N_3627);
xor U7244 (N_7244,N_2670,N_80);
nor U7245 (N_7245,N_1529,N_4098);
nand U7246 (N_7246,N_3496,N_2896);
or U7247 (N_7247,N_187,N_2705);
or U7248 (N_7248,N_1976,N_2244);
nor U7249 (N_7249,N_926,N_620);
or U7250 (N_7250,N_3311,N_1104);
nand U7251 (N_7251,N_2482,N_4877);
nand U7252 (N_7252,N_1190,N_4061);
and U7253 (N_7253,N_801,N_2909);
or U7254 (N_7254,N_2075,N_2325);
or U7255 (N_7255,N_4539,N_1246);
nor U7256 (N_7256,N_1148,N_3625);
and U7257 (N_7257,N_642,N_2011);
and U7258 (N_7258,N_4415,N_2921);
and U7259 (N_7259,N_1774,N_3681);
xor U7260 (N_7260,N_1056,N_2441);
or U7261 (N_7261,N_1750,N_1767);
and U7262 (N_7262,N_3852,N_3453);
and U7263 (N_7263,N_2078,N_1254);
xor U7264 (N_7264,N_3273,N_1042);
and U7265 (N_7265,N_1165,N_2249);
or U7266 (N_7266,N_4844,N_4409);
nor U7267 (N_7267,N_2025,N_889);
or U7268 (N_7268,N_4790,N_1915);
nand U7269 (N_7269,N_4169,N_2993);
or U7270 (N_7270,N_3301,N_2477);
nand U7271 (N_7271,N_2164,N_3377);
nand U7272 (N_7272,N_2846,N_109);
or U7273 (N_7273,N_2487,N_3305);
nor U7274 (N_7274,N_4173,N_2530);
nand U7275 (N_7275,N_1840,N_4766);
nand U7276 (N_7276,N_3442,N_3690);
and U7277 (N_7277,N_1256,N_4276);
nor U7278 (N_7278,N_575,N_602);
nor U7279 (N_7279,N_1420,N_4424);
nor U7280 (N_7280,N_3524,N_3956);
or U7281 (N_7281,N_536,N_2935);
nand U7282 (N_7282,N_1666,N_2197);
or U7283 (N_7283,N_2511,N_637);
nor U7284 (N_7284,N_1014,N_3508);
or U7285 (N_7285,N_1239,N_2146);
and U7286 (N_7286,N_2068,N_4182);
nand U7287 (N_7287,N_3632,N_1841);
nand U7288 (N_7288,N_2272,N_1210);
xor U7289 (N_7289,N_4809,N_1295);
xnor U7290 (N_7290,N_2014,N_2108);
or U7291 (N_7291,N_3076,N_1882);
xor U7292 (N_7292,N_3480,N_450);
and U7293 (N_7293,N_44,N_1757);
nor U7294 (N_7294,N_435,N_2042);
or U7295 (N_7295,N_4641,N_4974);
xnor U7296 (N_7296,N_1054,N_503);
nor U7297 (N_7297,N_4110,N_666);
nor U7298 (N_7298,N_1231,N_3640);
or U7299 (N_7299,N_4271,N_3668);
xor U7300 (N_7300,N_4105,N_3708);
xor U7301 (N_7301,N_3906,N_1855);
nand U7302 (N_7302,N_1046,N_2755);
or U7303 (N_7303,N_4203,N_480);
and U7304 (N_7304,N_1255,N_633);
and U7305 (N_7305,N_4925,N_322);
or U7306 (N_7306,N_1352,N_2060);
and U7307 (N_7307,N_4601,N_1907);
nor U7308 (N_7308,N_3070,N_4841);
nor U7309 (N_7309,N_1726,N_4025);
or U7310 (N_7310,N_3818,N_1832);
or U7311 (N_7311,N_3947,N_2761);
nand U7312 (N_7312,N_3764,N_3065);
nor U7313 (N_7313,N_3249,N_4222);
or U7314 (N_7314,N_2357,N_4723);
or U7315 (N_7315,N_1950,N_3004);
or U7316 (N_7316,N_4596,N_4113);
nor U7317 (N_7317,N_3353,N_245);
nor U7318 (N_7318,N_3584,N_3019);
nor U7319 (N_7319,N_4300,N_1118);
xor U7320 (N_7320,N_1959,N_440);
and U7321 (N_7321,N_2563,N_3536);
nand U7322 (N_7322,N_4964,N_775);
nor U7323 (N_7323,N_1531,N_2539);
nor U7324 (N_7324,N_3303,N_1683);
nand U7325 (N_7325,N_2198,N_4957);
or U7326 (N_7326,N_1536,N_4239);
or U7327 (N_7327,N_2816,N_898);
or U7328 (N_7328,N_4199,N_4313);
nor U7329 (N_7329,N_1070,N_173);
nand U7330 (N_7330,N_244,N_148);
nor U7331 (N_7331,N_1937,N_2062);
xor U7332 (N_7332,N_3209,N_4296);
nor U7333 (N_7333,N_4483,N_4187);
nor U7334 (N_7334,N_4002,N_250);
nand U7335 (N_7335,N_570,N_2489);
and U7336 (N_7336,N_4260,N_3720);
and U7337 (N_7337,N_4824,N_4619);
or U7338 (N_7338,N_1392,N_1482);
xor U7339 (N_7339,N_623,N_4747);
or U7340 (N_7340,N_672,N_2334);
nor U7341 (N_7341,N_327,N_4764);
or U7342 (N_7342,N_1360,N_747);
nand U7343 (N_7343,N_4769,N_3782);
xor U7344 (N_7344,N_1484,N_2013);
nand U7345 (N_7345,N_2823,N_4230);
nand U7346 (N_7346,N_4982,N_683);
nor U7347 (N_7347,N_4829,N_3468);
nor U7348 (N_7348,N_1631,N_759);
nand U7349 (N_7349,N_917,N_2973);
and U7350 (N_7350,N_2601,N_1989);
and U7351 (N_7351,N_3383,N_4865);
and U7352 (N_7352,N_987,N_1984);
nand U7353 (N_7353,N_2333,N_2889);
nor U7354 (N_7354,N_26,N_3896);
or U7355 (N_7355,N_2207,N_3939);
and U7356 (N_7356,N_1188,N_3771);
or U7357 (N_7357,N_2748,N_520);
and U7358 (N_7358,N_4998,N_2974);
nand U7359 (N_7359,N_3617,N_2012);
nand U7360 (N_7360,N_1387,N_1073);
and U7361 (N_7361,N_948,N_790);
xor U7362 (N_7362,N_2689,N_4327);
nor U7363 (N_7363,N_3113,N_4487);
and U7364 (N_7364,N_3971,N_4397);
nor U7365 (N_7365,N_1764,N_4733);
xnor U7366 (N_7366,N_3755,N_4054);
and U7367 (N_7367,N_2574,N_2991);
and U7368 (N_7368,N_1349,N_4861);
nor U7369 (N_7369,N_3867,N_2149);
xnor U7370 (N_7370,N_2747,N_3600);
nor U7371 (N_7371,N_1393,N_1340);
nor U7372 (N_7372,N_2279,N_1490);
xor U7373 (N_7373,N_2721,N_3763);
xnor U7374 (N_7374,N_463,N_3074);
and U7375 (N_7375,N_3793,N_372);
nand U7376 (N_7376,N_73,N_1026);
nand U7377 (N_7377,N_1378,N_2912);
nor U7378 (N_7378,N_1412,N_2566);
nor U7379 (N_7379,N_1491,N_1149);
and U7380 (N_7380,N_1455,N_1496);
and U7381 (N_7381,N_307,N_157);
or U7382 (N_7382,N_4211,N_1809);
or U7383 (N_7383,N_2847,N_4518);
or U7384 (N_7384,N_93,N_3350);
nor U7385 (N_7385,N_1322,N_273);
or U7386 (N_7386,N_2348,N_3254);
nor U7387 (N_7387,N_2629,N_4726);
nor U7388 (N_7388,N_4099,N_81);
or U7389 (N_7389,N_4860,N_4532);
nor U7390 (N_7390,N_3898,N_465);
xor U7391 (N_7391,N_2064,N_2099);
or U7392 (N_7392,N_3484,N_2830);
and U7393 (N_7393,N_662,N_3518);
and U7394 (N_7394,N_3360,N_2349);
or U7395 (N_7395,N_2568,N_1747);
nand U7396 (N_7396,N_1727,N_625);
and U7397 (N_7397,N_114,N_1366);
nor U7398 (N_7398,N_3300,N_4430);
nand U7399 (N_7399,N_843,N_342);
nor U7400 (N_7400,N_2104,N_4787);
nor U7401 (N_7401,N_2522,N_4627);
and U7402 (N_7402,N_1918,N_2150);
or U7403 (N_7403,N_821,N_1143);
nor U7404 (N_7404,N_2945,N_1623);
or U7405 (N_7405,N_3028,N_3660);
and U7406 (N_7406,N_2634,N_167);
and U7407 (N_7407,N_1313,N_4191);
nor U7408 (N_7408,N_832,N_3349);
and U7409 (N_7409,N_2565,N_658);
or U7410 (N_7410,N_499,N_1405);
nor U7411 (N_7411,N_3500,N_2100);
nor U7412 (N_7412,N_2686,N_3511);
or U7413 (N_7413,N_535,N_4756);
nand U7414 (N_7414,N_2418,N_2615);
and U7415 (N_7415,N_4033,N_3704);
nand U7416 (N_7416,N_63,N_1562);
xor U7417 (N_7417,N_2112,N_4905);
or U7418 (N_7418,N_425,N_2880);
nor U7419 (N_7419,N_1261,N_3153);
nand U7420 (N_7420,N_2293,N_786);
nand U7421 (N_7421,N_1139,N_2653);
and U7422 (N_7422,N_1316,N_3796);
and U7423 (N_7423,N_4642,N_1117);
and U7424 (N_7424,N_3925,N_1377);
nor U7425 (N_7425,N_2730,N_4777);
and U7426 (N_7426,N_3982,N_126);
nor U7427 (N_7427,N_2156,N_1462);
and U7428 (N_7428,N_72,N_3304);
and U7429 (N_7429,N_4801,N_2613);
nor U7430 (N_7430,N_420,N_4566);
or U7431 (N_7431,N_10,N_3414);
and U7432 (N_7432,N_367,N_1899);
or U7433 (N_7433,N_3036,N_3389);
or U7434 (N_7434,N_3822,N_2673);
nand U7435 (N_7435,N_2463,N_2018);
and U7436 (N_7436,N_742,N_447);
xnor U7437 (N_7437,N_4445,N_318);
or U7438 (N_7438,N_2377,N_4749);
nor U7439 (N_7439,N_4670,N_4283);
and U7440 (N_7440,N_2501,N_4659);
and U7441 (N_7441,N_1510,N_1418);
and U7442 (N_7442,N_3296,N_785);
or U7443 (N_7443,N_532,N_3843);
or U7444 (N_7444,N_4100,N_1534);
or U7445 (N_7445,N_1966,N_4692);
xnor U7446 (N_7446,N_4431,N_3188);
and U7447 (N_7447,N_2217,N_2363);
nand U7448 (N_7448,N_4455,N_2233);
nor U7449 (N_7449,N_4674,N_3130);
nand U7450 (N_7450,N_2142,N_2947);
and U7451 (N_7451,N_1628,N_1081);
nand U7452 (N_7452,N_4611,N_3035);
nand U7453 (N_7453,N_1987,N_554);
and U7454 (N_7454,N_711,N_2644);
or U7455 (N_7455,N_4770,N_1735);
and U7456 (N_7456,N_3639,N_474);
nor U7457 (N_7457,N_1662,N_2825);
and U7458 (N_7458,N_4789,N_4624);
xnor U7459 (N_7459,N_911,N_1159);
nand U7460 (N_7460,N_3084,N_323);
or U7461 (N_7461,N_2153,N_1243);
and U7462 (N_7462,N_922,N_515);
and U7463 (N_7463,N_1427,N_3846);
xnor U7464 (N_7464,N_946,N_2978);
nand U7465 (N_7465,N_3051,N_1468);
xor U7466 (N_7466,N_3426,N_4883);
xnor U7467 (N_7467,N_51,N_3006);
or U7468 (N_7468,N_3456,N_1589);
and U7469 (N_7469,N_3319,N_2583);
and U7470 (N_7470,N_610,N_4122);
and U7471 (N_7471,N_3437,N_2007);
or U7472 (N_7472,N_1890,N_4930);
and U7473 (N_7473,N_2323,N_4921);
xor U7474 (N_7474,N_1753,N_4177);
nor U7475 (N_7475,N_4318,N_4068);
and U7476 (N_7476,N_1602,N_3604);
nor U7477 (N_7477,N_1656,N_4488);
xnor U7478 (N_7478,N_3378,N_4150);
nor U7479 (N_7479,N_2172,N_846);
or U7480 (N_7480,N_4081,N_2772);
or U7481 (N_7481,N_849,N_2087);
and U7482 (N_7482,N_2685,N_1306);
or U7483 (N_7483,N_4540,N_4340);
and U7484 (N_7484,N_2300,N_296);
or U7485 (N_7485,N_1411,N_3370);
nand U7486 (N_7486,N_3786,N_988);
or U7487 (N_7487,N_4987,N_4019);
nand U7488 (N_7488,N_165,N_2376);
nor U7489 (N_7489,N_69,N_3012);
and U7490 (N_7490,N_1681,N_1333);
xnor U7491 (N_7491,N_195,N_1906);
or U7492 (N_7492,N_2056,N_1518);
nand U7493 (N_7493,N_466,N_3324);
or U7494 (N_7494,N_4804,N_3448);
nand U7495 (N_7495,N_1639,N_4551);
nand U7496 (N_7496,N_4171,N_1439);
nand U7497 (N_7497,N_1955,N_4742);
or U7498 (N_7498,N_3444,N_328);
and U7499 (N_7499,N_1359,N_614);
or U7500 (N_7500,N_4887,N_2697);
nor U7501 (N_7501,N_532,N_3505);
and U7502 (N_7502,N_4945,N_713);
nor U7503 (N_7503,N_475,N_4368);
or U7504 (N_7504,N_2032,N_2158);
and U7505 (N_7505,N_4240,N_470);
nor U7506 (N_7506,N_138,N_2086);
nor U7507 (N_7507,N_436,N_4659);
xnor U7508 (N_7508,N_664,N_2773);
nor U7509 (N_7509,N_1745,N_3906);
or U7510 (N_7510,N_563,N_320);
nor U7511 (N_7511,N_4321,N_4185);
xnor U7512 (N_7512,N_919,N_1419);
nand U7513 (N_7513,N_1580,N_4558);
nor U7514 (N_7514,N_3880,N_4808);
nor U7515 (N_7515,N_2462,N_466);
nand U7516 (N_7516,N_4980,N_3921);
and U7517 (N_7517,N_240,N_4294);
or U7518 (N_7518,N_2807,N_2787);
and U7519 (N_7519,N_622,N_1812);
xor U7520 (N_7520,N_4112,N_1982);
nand U7521 (N_7521,N_3898,N_533);
and U7522 (N_7522,N_2628,N_2774);
nand U7523 (N_7523,N_1462,N_4609);
nor U7524 (N_7524,N_999,N_834);
nor U7525 (N_7525,N_924,N_1472);
nand U7526 (N_7526,N_1616,N_388);
nor U7527 (N_7527,N_2085,N_2064);
nand U7528 (N_7528,N_4256,N_2072);
and U7529 (N_7529,N_1254,N_1369);
and U7530 (N_7530,N_1904,N_2739);
nand U7531 (N_7531,N_3627,N_1881);
nor U7532 (N_7532,N_2957,N_2655);
and U7533 (N_7533,N_142,N_730);
nor U7534 (N_7534,N_1522,N_1408);
or U7535 (N_7535,N_3749,N_4405);
and U7536 (N_7536,N_4178,N_4243);
and U7537 (N_7537,N_168,N_2929);
xor U7538 (N_7538,N_1057,N_2811);
nand U7539 (N_7539,N_184,N_3418);
xnor U7540 (N_7540,N_736,N_3432);
or U7541 (N_7541,N_1102,N_236);
nand U7542 (N_7542,N_1915,N_2315);
nand U7543 (N_7543,N_980,N_2848);
and U7544 (N_7544,N_4894,N_1168);
xor U7545 (N_7545,N_4017,N_3472);
or U7546 (N_7546,N_1899,N_4668);
xnor U7547 (N_7547,N_1222,N_746);
or U7548 (N_7548,N_2614,N_3199);
nor U7549 (N_7549,N_2443,N_4876);
xor U7550 (N_7550,N_1607,N_2738);
and U7551 (N_7551,N_291,N_2358);
and U7552 (N_7552,N_18,N_4911);
xor U7553 (N_7553,N_4192,N_2512);
nand U7554 (N_7554,N_4416,N_2746);
or U7555 (N_7555,N_1885,N_4732);
nor U7556 (N_7556,N_4671,N_2387);
nor U7557 (N_7557,N_4889,N_2507);
nor U7558 (N_7558,N_1309,N_3798);
nand U7559 (N_7559,N_3531,N_1666);
and U7560 (N_7560,N_3995,N_2839);
or U7561 (N_7561,N_1741,N_4296);
xnor U7562 (N_7562,N_278,N_4279);
nand U7563 (N_7563,N_1984,N_841);
xor U7564 (N_7564,N_2571,N_4972);
nor U7565 (N_7565,N_3403,N_1403);
and U7566 (N_7566,N_3608,N_1211);
or U7567 (N_7567,N_637,N_3300);
and U7568 (N_7568,N_3650,N_368);
nor U7569 (N_7569,N_3133,N_2047);
nand U7570 (N_7570,N_1675,N_2202);
and U7571 (N_7571,N_4215,N_239);
or U7572 (N_7572,N_1971,N_3737);
or U7573 (N_7573,N_4849,N_941);
nand U7574 (N_7574,N_1169,N_1111);
nor U7575 (N_7575,N_2741,N_196);
xnor U7576 (N_7576,N_4258,N_2375);
or U7577 (N_7577,N_3732,N_2822);
nand U7578 (N_7578,N_682,N_1424);
or U7579 (N_7579,N_2857,N_1319);
or U7580 (N_7580,N_2353,N_3708);
and U7581 (N_7581,N_4691,N_3367);
or U7582 (N_7582,N_110,N_4798);
and U7583 (N_7583,N_1780,N_525);
or U7584 (N_7584,N_3629,N_2638);
and U7585 (N_7585,N_2687,N_2283);
xnor U7586 (N_7586,N_3078,N_2670);
and U7587 (N_7587,N_2164,N_4888);
or U7588 (N_7588,N_1695,N_3251);
nand U7589 (N_7589,N_887,N_4266);
nor U7590 (N_7590,N_982,N_990);
or U7591 (N_7591,N_1721,N_4075);
or U7592 (N_7592,N_50,N_1114);
nand U7593 (N_7593,N_3412,N_4803);
nor U7594 (N_7594,N_1070,N_4097);
nand U7595 (N_7595,N_1401,N_3772);
nor U7596 (N_7596,N_1514,N_2892);
xor U7597 (N_7597,N_2124,N_4309);
xnor U7598 (N_7598,N_3363,N_1295);
and U7599 (N_7599,N_1232,N_4542);
or U7600 (N_7600,N_45,N_731);
or U7601 (N_7601,N_3140,N_2316);
xnor U7602 (N_7602,N_246,N_2460);
or U7603 (N_7603,N_2556,N_2774);
nor U7604 (N_7604,N_3751,N_3660);
and U7605 (N_7605,N_3139,N_3362);
and U7606 (N_7606,N_4053,N_2826);
or U7607 (N_7607,N_4352,N_3708);
and U7608 (N_7608,N_2085,N_3301);
and U7609 (N_7609,N_3167,N_4370);
and U7610 (N_7610,N_3137,N_1988);
and U7611 (N_7611,N_4265,N_1696);
nor U7612 (N_7612,N_1074,N_3917);
or U7613 (N_7613,N_4448,N_4076);
and U7614 (N_7614,N_3217,N_4654);
or U7615 (N_7615,N_1507,N_2326);
xor U7616 (N_7616,N_3182,N_357);
nor U7617 (N_7617,N_4231,N_553);
and U7618 (N_7618,N_2970,N_1413);
or U7619 (N_7619,N_2494,N_4367);
nor U7620 (N_7620,N_4470,N_1345);
nor U7621 (N_7621,N_1816,N_4812);
and U7622 (N_7622,N_1055,N_4505);
xor U7623 (N_7623,N_566,N_1546);
nor U7624 (N_7624,N_577,N_4986);
or U7625 (N_7625,N_1892,N_604);
xnor U7626 (N_7626,N_3844,N_4973);
nand U7627 (N_7627,N_2180,N_4503);
and U7628 (N_7628,N_15,N_2972);
and U7629 (N_7629,N_677,N_1718);
or U7630 (N_7630,N_4153,N_2615);
or U7631 (N_7631,N_3924,N_1790);
nand U7632 (N_7632,N_4580,N_2891);
and U7633 (N_7633,N_4815,N_2715);
xor U7634 (N_7634,N_2878,N_873);
nor U7635 (N_7635,N_4058,N_1659);
or U7636 (N_7636,N_4816,N_2472);
nand U7637 (N_7637,N_4741,N_1778);
xor U7638 (N_7638,N_3250,N_3405);
and U7639 (N_7639,N_2165,N_1627);
and U7640 (N_7640,N_3218,N_4491);
or U7641 (N_7641,N_2162,N_4642);
or U7642 (N_7642,N_2532,N_4540);
or U7643 (N_7643,N_4327,N_1052);
or U7644 (N_7644,N_2879,N_623);
nand U7645 (N_7645,N_3395,N_3772);
nor U7646 (N_7646,N_4279,N_4226);
or U7647 (N_7647,N_4916,N_4879);
nand U7648 (N_7648,N_15,N_4876);
nand U7649 (N_7649,N_4719,N_3269);
nor U7650 (N_7650,N_2161,N_1606);
nand U7651 (N_7651,N_3206,N_2363);
and U7652 (N_7652,N_969,N_4931);
and U7653 (N_7653,N_2922,N_1601);
or U7654 (N_7654,N_2886,N_4142);
and U7655 (N_7655,N_989,N_2423);
and U7656 (N_7656,N_2508,N_3124);
or U7657 (N_7657,N_2982,N_4830);
or U7658 (N_7658,N_2316,N_2034);
nor U7659 (N_7659,N_4482,N_1481);
and U7660 (N_7660,N_771,N_4678);
and U7661 (N_7661,N_4485,N_450);
or U7662 (N_7662,N_4038,N_38);
and U7663 (N_7663,N_2930,N_235);
nand U7664 (N_7664,N_733,N_3022);
or U7665 (N_7665,N_2686,N_4886);
and U7666 (N_7666,N_2961,N_2299);
and U7667 (N_7667,N_3910,N_899);
nor U7668 (N_7668,N_4460,N_4765);
or U7669 (N_7669,N_4273,N_2272);
and U7670 (N_7670,N_1229,N_3269);
and U7671 (N_7671,N_2588,N_4988);
or U7672 (N_7672,N_1687,N_4252);
and U7673 (N_7673,N_3505,N_2588);
nor U7674 (N_7674,N_2503,N_3013);
nand U7675 (N_7675,N_1680,N_3988);
nand U7676 (N_7676,N_506,N_4639);
and U7677 (N_7677,N_1415,N_3801);
and U7678 (N_7678,N_2318,N_2316);
nand U7679 (N_7679,N_2012,N_2825);
nor U7680 (N_7680,N_3751,N_3387);
xor U7681 (N_7681,N_3467,N_2142);
nand U7682 (N_7682,N_2939,N_4472);
and U7683 (N_7683,N_4133,N_4919);
or U7684 (N_7684,N_3,N_1657);
or U7685 (N_7685,N_2240,N_3275);
xor U7686 (N_7686,N_113,N_4887);
nand U7687 (N_7687,N_2250,N_1040);
xnor U7688 (N_7688,N_1007,N_3837);
nand U7689 (N_7689,N_3729,N_1197);
nand U7690 (N_7690,N_640,N_4383);
or U7691 (N_7691,N_1276,N_3617);
xnor U7692 (N_7692,N_4556,N_4853);
nor U7693 (N_7693,N_864,N_4721);
nor U7694 (N_7694,N_2109,N_2729);
nand U7695 (N_7695,N_3646,N_3286);
nor U7696 (N_7696,N_804,N_138);
and U7697 (N_7697,N_1217,N_3169);
nor U7698 (N_7698,N_3146,N_2121);
nand U7699 (N_7699,N_4306,N_4396);
and U7700 (N_7700,N_1832,N_2953);
nand U7701 (N_7701,N_2210,N_2703);
or U7702 (N_7702,N_4617,N_2130);
or U7703 (N_7703,N_2456,N_1459);
and U7704 (N_7704,N_3448,N_4955);
nor U7705 (N_7705,N_1238,N_2786);
nand U7706 (N_7706,N_548,N_3706);
and U7707 (N_7707,N_3680,N_551);
or U7708 (N_7708,N_4483,N_4339);
or U7709 (N_7709,N_1716,N_380);
and U7710 (N_7710,N_2794,N_3386);
nor U7711 (N_7711,N_4105,N_1816);
nand U7712 (N_7712,N_4173,N_1255);
nor U7713 (N_7713,N_1960,N_3445);
or U7714 (N_7714,N_1573,N_3067);
and U7715 (N_7715,N_1089,N_3080);
xnor U7716 (N_7716,N_3012,N_3895);
or U7717 (N_7717,N_4700,N_720);
and U7718 (N_7718,N_1581,N_314);
nand U7719 (N_7719,N_3196,N_2730);
or U7720 (N_7720,N_4567,N_3456);
nand U7721 (N_7721,N_213,N_312);
or U7722 (N_7722,N_2083,N_1737);
xnor U7723 (N_7723,N_1484,N_1631);
and U7724 (N_7724,N_3275,N_4527);
or U7725 (N_7725,N_46,N_483);
nand U7726 (N_7726,N_98,N_740);
nor U7727 (N_7727,N_722,N_3519);
or U7728 (N_7728,N_1579,N_1198);
and U7729 (N_7729,N_4801,N_1642);
nand U7730 (N_7730,N_3279,N_3171);
nand U7731 (N_7731,N_1746,N_447);
or U7732 (N_7732,N_3991,N_1918);
and U7733 (N_7733,N_2067,N_1727);
or U7734 (N_7734,N_4473,N_1681);
nor U7735 (N_7735,N_4835,N_4425);
xor U7736 (N_7736,N_1194,N_4118);
or U7737 (N_7737,N_3001,N_1793);
or U7738 (N_7738,N_4704,N_1635);
nand U7739 (N_7739,N_135,N_1863);
or U7740 (N_7740,N_3593,N_4711);
and U7741 (N_7741,N_2117,N_3186);
or U7742 (N_7742,N_4525,N_2943);
xor U7743 (N_7743,N_1946,N_1336);
or U7744 (N_7744,N_4098,N_2394);
nand U7745 (N_7745,N_849,N_3369);
nand U7746 (N_7746,N_3437,N_1608);
nand U7747 (N_7747,N_3051,N_32);
and U7748 (N_7748,N_4127,N_4395);
and U7749 (N_7749,N_4050,N_101);
or U7750 (N_7750,N_266,N_4936);
nand U7751 (N_7751,N_1442,N_4655);
nand U7752 (N_7752,N_1769,N_3524);
and U7753 (N_7753,N_2109,N_2619);
or U7754 (N_7754,N_3979,N_868);
and U7755 (N_7755,N_2909,N_2043);
xnor U7756 (N_7756,N_4899,N_1300);
nand U7757 (N_7757,N_3424,N_1680);
or U7758 (N_7758,N_4001,N_3647);
xnor U7759 (N_7759,N_509,N_3595);
or U7760 (N_7760,N_559,N_1297);
or U7761 (N_7761,N_3574,N_2892);
nand U7762 (N_7762,N_1386,N_1888);
and U7763 (N_7763,N_4506,N_2879);
nor U7764 (N_7764,N_391,N_917);
nand U7765 (N_7765,N_2684,N_483);
or U7766 (N_7766,N_2806,N_2137);
nand U7767 (N_7767,N_3095,N_601);
nor U7768 (N_7768,N_870,N_2287);
and U7769 (N_7769,N_4682,N_1374);
or U7770 (N_7770,N_821,N_3101);
nor U7771 (N_7771,N_1777,N_744);
nor U7772 (N_7772,N_1951,N_3055);
nor U7773 (N_7773,N_1939,N_4704);
nand U7774 (N_7774,N_4825,N_671);
nor U7775 (N_7775,N_3859,N_1854);
or U7776 (N_7776,N_3365,N_90);
or U7777 (N_7777,N_3672,N_3135);
nand U7778 (N_7778,N_4888,N_206);
nor U7779 (N_7779,N_4714,N_1920);
nand U7780 (N_7780,N_3982,N_612);
nor U7781 (N_7781,N_3483,N_3094);
nor U7782 (N_7782,N_4912,N_2628);
or U7783 (N_7783,N_2096,N_1414);
nor U7784 (N_7784,N_3091,N_1738);
and U7785 (N_7785,N_491,N_943);
nand U7786 (N_7786,N_2324,N_1027);
nor U7787 (N_7787,N_2621,N_4703);
nor U7788 (N_7788,N_2097,N_1807);
or U7789 (N_7789,N_4187,N_3221);
or U7790 (N_7790,N_1078,N_2170);
nor U7791 (N_7791,N_1535,N_2384);
or U7792 (N_7792,N_2440,N_1536);
xnor U7793 (N_7793,N_1197,N_2891);
nor U7794 (N_7794,N_164,N_3420);
xnor U7795 (N_7795,N_4281,N_870);
or U7796 (N_7796,N_1009,N_2481);
or U7797 (N_7797,N_833,N_16);
or U7798 (N_7798,N_4965,N_3943);
and U7799 (N_7799,N_4800,N_4983);
or U7800 (N_7800,N_818,N_675);
and U7801 (N_7801,N_816,N_3974);
nand U7802 (N_7802,N_3152,N_1930);
and U7803 (N_7803,N_4250,N_2701);
nor U7804 (N_7804,N_696,N_3388);
and U7805 (N_7805,N_2616,N_527);
or U7806 (N_7806,N_373,N_4982);
nand U7807 (N_7807,N_3338,N_2897);
and U7808 (N_7808,N_4037,N_3673);
xor U7809 (N_7809,N_2459,N_2147);
xor U7810 (N_7810,N_2912,N_4550);
and U7811 (N_7811,N_3311,N_1607);
and U7812 (N_7812,N_4223,N_4049);
nor U7813 (N_7813,N_551,N_280);
nor U7814 (N_7814,N_1331,N_3624);
nand U7815 (N_7815,N_2146,N_2554);
xnor U7816 (N_7816,N_2750,N_3401);
nand U7817 (N_7817,N_2172,N_4403);
nand U7818 (N_7818,N_3854,N_143);
or U7819 (N_7819,N_2495,N_1859);
nor U7820 (N_7820,N_48,N_4050);
or U7821 (N_7821,N_1307,N_3255);
and U7822 (N_7822,N_2274,N_1508);
nand U7823 (N_7823,N_1297,N_626);
nor U7824 (N_7824,N_1831,N_773);
nor U7825 (N_7825,N_911,N_4783);
or U7826 (N_7826,N_351,N_3151);
and U7827 (N_7827,N_492,N_4764);
or U7828 (N_7828,N_4367,N_1480);
and U7829 (N_7829,N_340,N_2873);
nor U7830 (N_7830,N_1480,N_3663);
and U7831 (N_7831,N_3177,N_2623);
xor U7832 (N_7832,N_572,N_1580);
and U7833 (N_7833,N_3972,N_4848);
or U7834 (N_7834,N_1012,N_912);
and U7835 (N_7835,N_2178,N_2387);
and U7836 (N_7836,N_1445,N_4899);
or U7837 (N_7837,N_4119,N_2347);
or U7838 (N_7838,N_4416,N_2436);
nor U7839 (N_7839,N_2691,N_1019);
and U7840 (N_7840,N_137,N_1440);
or U7841 (N_7841,N_3959,N_1888);
and U7842 (N_7842,N_252,N_644);
or U7843 (N_7843,N_4054,N_2877);
or U7844 (N_7844,N_2044,N_3674);
nand U7845 (N_7845,N_3209,N_4260);
nand U7846 (N_7846,N_3345,N_69);
nor U7847 (N_7847,N_2270,N_4223);
nor U7848 (N_7848,N_3384,N_4720);
nand U7849 (N_7849,N_4176,N_3015);
xnor U7850 (N_7850,N_1877,N_129);
nor U7851 (N_7851,N_2252,N_1592);
xor U7852 (N_7852,N_2244,N_1891);
and U7853 (N_7853,N_3609,N_4303);
nor U7854 (N_7854,N_1419,N_3519);
nor U7855 (N_7855,N_3204,N_197);
xor U7856 (N_7856,N_4123,N_4456);
nor U7857 (N_7857,N_117,N_3642);
and U7858 (N_7858,N_487,N_3123);
or U7859 (N_7859,N_839,N_4082);
and U7860 (N_7860,N_262,N_1169);
or U7861 (N_7861,N_855,N_4048);
nand U7862 (N_7862,N_2074,N_4146);
or U7863 (N_7863,N_2541,N_1768);
and U7864 (N_7864,N_101,N_2040);
nor U7865 (N_7865,N_805,N_1718);
nand U7866 (N_7866,N_480,N_783);
nor U7867 (N_7867,N_390,N_498);
or U7868 (N_7868,N_4184,N_4874);
nand U7869 (N_7869,N_3667,N_3277);
xnor U7870 (N_7870,N_1940,N_4289);
nor U7871 (N_7871,N_2635,N_1214);
nor U7872 (N_7872,N_788,N_3686);
and U7873 (N_7873,N_3152,N_1073);
or U7874 (N_7874,N_417,N_4006);
xor U7875 (N_7875,N_118,N_1841);
nand U7876 (N_7876,N_1562,N_1924);
nor U7877 (N_7877,N_1157,N_4515);
nor U7878 (N_7878,N_2257,N_2927);
nand U7879 (N_7879,N_2647,N_2976);
and U7880 (N_7880,N_2069,N_3964);
nor U7881 (N_7881,N_1207,N_1848);
or U7882 (N_7882,N_2624,N_1768);
nor U7883 (N_7883,N_2350,N_282);
nand U7884 (N_7884,N_3048,N_2825);
or U7885 (N_7885,N_4345,N_1463);
nand U7886 (N_7886,N_731,N_675);
nand U7887 (N_7887,N_691,N_1554);
nor U7888 (N_7888,N_3886,N_2285);
or U7889 (N_7889,N_2852,N_149);
or U7890 (N_7890,N_211,N_1121);
nor U7891 (N_7891,N_3769,N_2492);
xor U7892 (N_7892,N_4266,N_3659);
and U7893 (N_7893,N_2865,N_63);
nand U7894 (N_7894,N_3442,N_2892);
or U7895 (N_7895,N_1869,N_4364);
or U7896 (N_7896,N_3291,N_1343);
nor U7897 (N_7897,N_1990,N_1674);
nor U7898 (N_7898,N_2366,N_2619);
or U7899 (N_7899,N_1291,N_1419);
or U7900 (N_7900,N_3179,N_3734);
nor U7901 (N_7901,N_975,N_2227);
and U7902 (N_7902,N_410,N_3365);
xor U7903 (N_7903,N_507,N_441);
or U7904 (N_7904,N_1812,N_4220);
nand U7905 (N_7905,N_4560,N_1113);
nand U7906 (N_7906,N_2788,N_3813);
nor U7907 (N_7907,N_2891,N_1969);
nor U7908 (N_7908,N_696,N_4221);
and U7909 (N_7909,N_1006,N_2767);
or U7910 (N_7910,N_1147,N_561);
nor U7911 (N_7911,N_101,N_2428);
nand U7912 (N_7912,N_889,N_4643);
nand U7913 (N_7913,N_4746,N_4807);
nand U7914 (N_7914,N_2103,N_1155);
and U7915 (N_7915,N_4863,N_3499);
xnor U7916 (N_7916,N_2672,N_1884);
or U7917 (N_7917,N_1043,N_1359);
nor U7918 (N_7918,N_3376,N_2993);
and U7919 (N_7919,N_2994,N_1921);
xnor U7920 (N_7920,N_1897,N_2832);
nor U7921 (N_7921,N_2393,N_2578);
nand U7922 (N_7922,N_4430,N_4890);
xnor U7923 (N_7923,N_2718,N_1216);
nor U7924 (N_7924,N_4153,N_3177);
or U7925 (N_7925,N_2169,N_3890);
or U7926 (N_7926,N_1254,N_3538);
or U7927 (N_7927,N_1096,N_3042);
or U7928 (N_7928,N_1151,N_586);
and U7929 (N_7929,N_1634,N_3055);
and U7930 (N_7930,N_176,N_510);
xnor U7931 (N_7931,N_592,N_2728);
and U7932 (N_7932,N_463,N_3239);
and U7933 (N_7933,N_3516,N_3499);
and U7934 (N_7934,N_4160,N_2844);
xor U7935 (N_7935,N_1411,N_3062);
and U7936 (N_7936,N_1583,N_2045);
nor U7937 (N_7937,N_2483,N_2291);
nor U7938 (N_7938,N_1727,N_3642);
nor U7939 (N_7939,N_4016,N_1584);
nand U7940 (N_7940,N_3515,N_780);
or U7941 (N_7941,N_3149,N_3320);
nand U7942 (N_7942,N_3434,N_3842);
or U7943 (N_7943,N_2713,N_3671);
nor U7944 (N_7944,N_4727,N_2944);
and U7945 (N_7945,N_1153,N_4070);
and U7946 (N_7946,N_3544,N_2301);
nand U7947 (N_7947,N_4443,N_3472);
xnor U7948 (N_7948,N_2496,N_36);
nand U7949 (N_7949,N_3870,N_1740);
nor U7950 (N_7950,N_4605,N_1334);
or U7951 (N_7951,N_2420,N_578);
nor U7952 (N_7952,N_3211,N_2015);
nor U7953 (N_7953,N_3807,N_2523);
or U7954 (N_7954,N_4316,N_4);
or U7955 (N_7955,N_4011,N_2989);
and U7956 (N_7956,N_509,N_3909);
nor U7957 (N_7957,N_2203,N_2234);
nor U7958 (N_7958,N_4236,N_593);
or U7959 (N_7959,N_1777,N_3529);
or U7960 (N_7960,N_4771,N_3973);
or U7961 (N_7961,N_2597,N_3703);
nor U7962 (N_7962,N_1731,N_708);
or U7963 (N_7963,N_977,N_44);
nand U7964 (N_7964,N_4184,N_4547);
and U7965 (N_7965,N_83,N_4538);
and U7966 (N_7966,N_680,N_3589);
nand U7967 (N_7967,N_1770,N_3634);
xor U7968 (N_7968,N_2941,N_1777);
nor U7969 (N_7969,N_3812,N_2775);
nor U7970 (N_7970,N_3827,N_2820);
and U7971 (N_7971,N_4631,N_4819);
and U7972 (N_7972,N_83,N_1133);
xor U7973 (N_7973,N_3688,N_2392);
nor U7974 (N_7974,N_3851,N_2506);
nand U7975 (N_7975,N_2474,N_964);
xnor U7976 (N_7976,N_3516,N_726);
nor U7977 (N_7977,N_1602,N_3768);
xnor U7978 (N_7978,N_2572,N_412);
or U7979 (N_7979,N_2743,N_4698);
nand U7980 (N_7980,N_3374,N_2345);
nand U7981 (N_7981,N_2259,N_3954);
and U7982 (N_7982,N_3822,N_1051);
nor U7983 (N_7983,N_2486,N_1502);
nand U7984 (N_7984,N_3261,N_937);
and U7985 (N_7985,N_982,N_4874);
nor U7986 (N_7986,N_2433,N_1112);
and U7987 (N_7987,N_3411,N_813);
nor U7988 (N_7988,N_3656,N_3327);
nor U7989 (N_7989,N_4445,N_3086);
nand U7990 (N_7990,N_4346,N_1212);
nand U7991 (N_7991,N_3227,N_4871);
and U7992 (N_7992,N_4871,N_3635);
nand U7993 (N_7993,N_3019,N_407);
or U7994 (N_7994,N_4567,N_1762);
nor U7995 (N_7995,N_3439,N_351);
or U7996 (N_7996,N_1842,N_3192);
nor U7997 (N_7997,N_2512,N_4588);
nand U7998 (N_7998,N_4843,N_3875);
nor U7999 (N_7999,N_3875,N_2024);
xor U8000 (N_8000,N_2789,N_4998);
and U8001 (N_8001,N_353,N_985);
xor U8002 (N_8002,N_4801,N_2818);
or U8003 (N_8003,N_4828,N_2143);
or U8004 (N_8004,N_1222,N_2841);
nand U8005 (N_8005,N_1612,N_101);
or U8006 (N_8006,N_470,N_2322);
nor U8007 (N_8007,N_3139,N_208);
nor U8008 (N_8008,N_2858,N_1552);
or U8009 (N_8009,N_3118,N_14);
xor U8010 (N_8010,N_397,N_3729);
nor U8011 (N_8011,N_1418,N_3428);
and U8012 (N_8012,N_4534,N_4084);
or U8013 (N_8013,N_1427,N_3549);
nand U8014 (N_8014,N_1994,N_3811);
and U8015 (N_8015,N_3884,N_335);
nor U8016 (N_8016,N_94,N_967);
nand U8017 (N_8017,N_230,N_4171);
xor U8018 (N_8018,N_3984,N_2762);
nand U8019 (N_8019,N_3627,N_2830);
nor U8020 (N_8020,N_368,N_4693);
or U8021 (N_8021,N_889,N_4000);
xnor U8022 (N_8022,N_2411,N_2675);
and U8023 (N_8023,N_2195,N_2243);
nor U8024 (N_8024,N_3155,N_4373);
or U8025 (N_8025,N_2708,N_1902);
xor U8026 (N_8026,N_2183,N_124);
and U8027 (N_8027,N_3662,N_4929);
nand U8028 (N_8028,N_1052,N_776);
nand U8029 (N_8029,N_3185,N_12);
and U8030 (N_8030,N_1780,N_2447);
nand U8031 (N_8031,N_4497,N_474);
nor U8032 (N_8032,N_4749,N_1816);
nor U8033 (N_8033,N_2016,N_2333);
nor U8034 (N_8034,N_4424,N_441);
or U8035 (N_8035,N_4619,N_3693);
nand U8036 (N_8036,N_1417,N_412);
nor U8037 (N_8037,N_2552,N_3557);
and U8038 (N_8038,N_4931,N_4686);
nor U8039 (N_8039,N_1501,N_2196);
and U8040 (N_8040,N_263,N_1572);
or U8041 (N_8041,N_2083,N_1460);
and U8042 (N_8042,N_2056,N_3338);
nor U8043 (N_8043,N_2421,N_1068);
or U8044 (N_8044,N_894,N_483);
nand U8045 (N_8045,N_1247,N_1812);
and U8046 (N_8046,N_1138,N_1217);
nand U8047 (N_8047,N_321,N_3921);
and U8048 (N_8048,N_4257,N_1393);
and U8049 (N_8049,N_2351,N_3664);
nor U8050 (N_8050,N_4717,N_2595);
nor U8051 (N_8051,N_1091,N_1872);
xor U8052 (N_8052,N_3647,N_62);
or U8053 (N_8053,N_2010,N_347);
and U8054 (N_8054,N_157,N_3292);
xor U8055 (N_8055,N_4620,N_4170);
xor U8056 (N_8056,N_3020,N_315);
nor U8057 (N_8057,N_2146,N_1155);
nor U8058 (N_8058,N_1962,N_2512);
nand U8059 (N_8059,N_592,N_3926);
nor U8060 (N_8060,N_1567,N_2623);
nor U8061 (N_8061,N_999,N_4566);
nand U8062 (N_8062,N_1423,N_3695);
or U8063 (N_8063,N_1169,N_2530);
nand U8064 (N_8064,N_873,N_335);
xor U8065 (N_8065,N_2890,N_3593);
xnor U8066 (N_8066,N_891,N_2320);
nand U8067 (N_8067,N_213,N_2538);
and U8068 (N_8068,N_4805,N_4756);
and U8069 (N_8069,N_1762,N_3519);
or U8070 (N_8070,N_3830,N_2224);
nor U8071 (N_8071,N_2267,N_141);
or U8072 (N_8072,N_1028,N_4574);
and U8073 (N_8073,N_1647,N_1063);
and U8074 (N_8074,N_1573,N_1805);
nor U8075 (N_8075,N_3889,N_251);
nand U8076 (N_8076,N_2607,N_2754);
and U8077 (N_8077,N_3770,N_839);
xnor U8078 (N_8078,N_3476,N_2322);
nand U8079 (N_8079,N_2106,N_1476);
xnor U8080 (N_8080,N_2173,N_63);
and U8081 (N_8081,N_1708,N_4564);
or U8082 (N_8082,N_4732,N_4685);
and U8083 (N_8083,N_384,N_2559);
nor U8084 (N_8084,N_3077,N_4866);
and U8085 (N_8085,N_1499,N_2299);
xor U8086 (N_8086,N_3536,N_1818);
or U8087 (N_8087,N_226,N_3351);
xor U8088 (N_8088,N_3141,N_3739);
and U8089 (N_8089,N_810,N_2685);
xor U8090 (N_8090,N_1475,N_1831);
nor U8091 (N_8091,N_3094,N_4711);
and U8092 (N_8092,N_4029,N_3667);
and U8093 (N_8093,N_2848,N_441);
nor U8094 (N_8094,N_2630,N_2112);
nor U8095 (N_8095,N_2040,N_3851);
nand U8096 (N_8096,N_998,N_3591);
or U8097 (N_8097,N_3502,N_3901);
and U8098 (N_8098,N_4602,N_3687);
or U8099 (N_8099,N_1174,N_2393);
nand U8100 (N_8100,N_1933,N_1555);
nor U8101 (N_8101,N_531,N_1688);
and U8102 (N_8102,N_1755,N_1942);
and U8103 (N_8103,N_4635,N_4855);
xor U8104 (N_8104,N_1600,N_4252);
or U8105 (N_8105,N_3396,N_247);
or U8106 (N_8106,N_2071,N_1599);
nor U8107 (N_8107,N_3282,N_1739);
nor U8108 (N_8108,N_4101,N_1788);
nor U8109 (N_8109,N_838,N_869);
or U8110 (N_8110,N_3311,N_4940);
nand U8111 (N_8111,N_3641,N_4719);
nor U8112 (N_8112,N_1852,N_3381);
nand U8113 (N_8113,N_1602,N_4327);
nor U8114 (N_8114,N_4289,N_2208);
nand U8115 (N_8115,N_1087,N_1633);
nand U8116 (N_8116,N_4078,N_766);
or U8117 (N_8117,N_3861,N_4884);
and U8118 (N_8118,N_4601,N_1594);
nor U8119 (N_8119,N_4984,N_2502);
xnor U8120 (N_8120,N_542,N_4885);
nand U8121 (N_8121,N_1194,N_833);
or U8122 (N_8122,N_3552,N_521);
and U8123 (N_8123,N_3092,N_3629);
xnor U8124 (N_8124,N_1479,N_4347);
or U8125 (N_8125,N_171,N_1739);
nand U8126 (N_8126,N_1532,N_799);
or U8127 (N_8127,N_1923,N_1595);
and U8128 (N_8128,N_3258,N_2858);
xor U8129 (N_8129,N_2544,N_232);
and U8130 (N_8130,N_3156,N_1803);
and U8131 (N_8131,N_2127,N_2852);
nor U8132 (N_8132,N_4667,N_4552);
nor U8133 (N_8133,N_4041,N_2957);
or U8134 (N_8134,N_3208,N_3884);
or U8135 (N_8135,N_675,N_4586);
nor U8136 (N_8136,N_1586,N_2972);
or U8137 (N_8137,N_5,N_3252);
xor U8138 (N_8138,N_1338,N_1368);
nand U8139 (N_8139,N_2397,N_4772);
nor U8140 (N_8140,N_2963,N_4785);
nand U8141 (N_8141,N_4202,N_38);
nor U8142 (N_8142,N_3945,N_352);
or U8143 (N_8143,N_4436,N_3721);
nand U8144 (N_8144,N_722,N_27);
nand U8145 (N_8145,N_4500,N_210);
or U8146 (N_8146,N_2010,N_2155);
nand U8147 (N_8147,N_3225,N_263);
or U8148 (N_8148,N_897,N_4179);
nor U8149 (N_8149,N_113,N_3549);
nand U8150 (N_8150,N_182,N_3115);
xor U8151 (N_8151,N_793,N_1390);
and U8152 (N_8152,N_4275,N_2745);
nor U8153 (N_8153,N_2000,N_1721);
and U8154 (N_8154,N_958,N_434);
nor U8155 (N_8155,N_4571,N_2690);
nand U8156 (N_8156,N_2693,N_3519);
and U8157 (N_8157,N_3594,N_1198);
and U8158 (N_8158,N_1828,N_2518);
or U8159 (N_8159,N_2469,N_2617);
xor U8160 (N_8160,N_2800,N_2737);
nor U8161 (N_8161,N_417,N_1247);
xnor U8162 (N_8162,N_1751,N_4100);
nor U8163 (N_8163,N_4495,N_2058);
xor U8164 (N_8164,N_1557,N_3221);
xor U8165 (N_8165,N_2558,N_3083);
xor U8166 (N_8166,N_3527,N_4556);
or U8167 (N_8167,N_2719,N_985);
nand U8168 (N_8168,N_2024,N_210);
or U8169 (N_8169,N_4084,N_3752);
nor U8170 (N_8170,N_3503,N_3223);
nor U8171 (N_8171,N_2221,N_4585);
xnor U8172 (N_8172,N_2352,N_4991);
or U8173 (N_8173,N_1071,N_3616);
nand U8174 (N_8174,N_962,N_3024);
or U8175 (N_8175,N_2321,N_2100);
and U8176 (N_8176,N_4349,N_368);
or U8177 (N_8177,N_2906,N_4562);
nor U8178 (N_8178,N_1623,N_2594);
nor U8179 (N_8179,N_1724,N_1947);
nand U8180 (N_8180,N_3007,N_1680);
nand U8181 (N_8181,N_4879,N_794);
nand U8182 (N_8182,N_2184,N_4948);
nand U8183 (N_8183,N_411,N_2131);
and U8184 (N_8184,N_3800,N_4980);
nor U8185 (N_8185,N_2043,N_4827);
xor U8186 (N_8186,N_2457,N_615);
or U8187 (N_8187,N_4858,N_1009);
nand U8188 (N_8188,N_4224,N_1668);
nand U8189 (N_8189,N_2186,N_4161);
nor U8190 (N_8190,N_2134,N_4748);
or U8191 (N_8191,N_3919,N_2379);
and U8192 (N_8192,N_2570,N_4900);
and U8193 (N_8193,N_706,N_2267);
nand U8194 (N_8194,N_2305,N_1363);
and U8195 (N_8195,N_3587,N_967);
and U8196 (N_8196,N_4113,N_3204);
nor U8197 (N_8197,N_2123,N_2803);
xnor U8198 (N_8198,N_1871,N_1709);
or U8199 (N_8199,N_1964,N_764);
or U8200 (N_8200,N_186,N_3567);
nor U8201 (N_8201,N_2024,N_2480);
or U8202 (N_8202,N_145,N_2593);
or U8203 (N_8203,N_4862,N_400);
nor U8204 (N_8204,N_2052,N_2307);
nand U8205 (N_8205,N_579,N_2269);
and U8206 (N_8206,N_2409,N_313);
xnor U8207 (N_8207,N_2450,N_4696);
xnor U8208 (N_8208,N_1662,N_3251);
nand U8209 (N_8209,N_3222,N_967);
nand U8210 (N_8210,N_2037,N_3737);
nand U8211 (N_8211,N_4030,N_4354);
nor U8212 (N_8212,N_2478,N_4758);
and U8213 (N_8213,N_3254,N_1309);
nor U8214 (N_8214,N_3981,N_2574);
or U8215 (N_8215,N_4118,N_4191);
nand U8216 (N_8216,N_914,N_513);
or U8217 (N_8217,N_3198,N_2234);
nand U8218 (N_8218,N_1201,N_4941);
and U8219 (N_8219,N_4867,N_4041);
nand U8220 (N_8220,N_3521,N_2087);
nand U8221 (N_8221,N_1281,N_4205);
or U8222 (N_8222,N_2644,N_1818);
nor U8223 (N_8223,N_2852,N_4584);
and U8224 (N_8224,N_208,N_3785);
or U8225 (N_8225,N_3532,N_1261);
and U8226 (N_8226,N_1592,N_4396);
xnor U8227 (N_8227,N_4188,N_136);
nand U8228 (N_8228,N_2620,N_3409);
xnor U8229 (N_8229,N_1641,N_4946);
xor U8230 (N_8230,N_1024,N_2840);
or U8231 (N_8231,N_1849,N_92);
nand U8232 (N_8232,N_769,N_2704);
or U8233 (N_8233,N_361,N_110);
nor U8234 (N_8234,N_233,N_4469);
nor U8235 (N_8235,N_47,N_2605);
nor U8236 (N_8236,N_1123,N_4477);
nand U8237 (N_8237,N_3906,N_4714);
and U8238 (N_8238,N_995,N_3125);
nor U8239 (N_8239,N_947,N_4477);
and U8240 (N_8240,N_3061,N_1017);
nor U8241 (N_8241,N_4021,N_158);
or U8242 (N_8242,N_3788,N_4834);
nand U8243 (N_8243,N_190,N_856);
and U8244 (N_8244,N_586,N_134);
and U8245 (N_8245,N_3031,N_1131);
nand U8246 (N_8246,N_1936,N_1550);
or U8247 (N_8247,N_4549,N_3564);
nor U8248 (N_8248,N_3710,N_2944);
or U8249 (N_8249,N_2909,N_3770);
or U8250 (N_8250,N_4294,N_4645);
xor U8251 (N_8251,N_4688,N_2801);
nor U8252 (N_8252,N_3872,N_705);
nor U8253 (N_8253,N_4000,N_1833);
nor U8254 (N_8254,N_1421,N_3939);
or U8255 (N_8255,N_2399,N_1348);
nor U8256 (N_8256,N_4817,N_2316);
nand U8257 (N_8257,N_4922,N_379);
nand U8258 (N_8258,N_1400,N_2872);
and U8259 (N_8259,N_2147,N_3663);
nand U8260 (N_8260,N_3278,N_3860);
nand U8261 (N_8261,N_593,N_4526);
or U8262 (N_8262,N_634,N_2680);
and U8263 (N_8263,N_4064,N_3347);
and U8264 (N_8264,N_2975,N_2816);
nand U8265 (N_8265,N_4973,N_3241);
or U8266 (N_8266,N_3705,N_3967);
and U8267 (N_8267,N_569,N_2800);
nand U8268 (N_8268,N_4565,N_2399);
nand U8269 (N_8269,N_4467,N_4154);
xor U8270 (N_8270,N_1248,N_498);
or U8271 (N_8271,N_4717,N_2297);
and U8272 (N_8272,N_3431,N_405);
or U8273 (N_8273,N_824,N_636);
or U8274 (N_8274,N_950,N_630);
nand U8275 (N_8275,N_861,N_1884);
xnor U8276 (N_8276,N_1392,N_2170);
nor U8277 (N_8277,N_354,N_2297);
nand U8278 (N_8278,N_1150,N_2584);
xor U8279 (N_8279,N_4092,N_4742);
and U8280 (N_8280,N_4609,N_2184);
and U8281 (N_8281,N_2151,N_1403);
or U8282 (N_8282,N_3618,N_2186);
nand U8283 (N_8283,N_2188,N_1589);
and U8284 (N_8284,N_387,N_1980);
or U8285 (N_8285,N_3681,N_4987);
nand U8286 (N_8286,N_1700,N_2835);
and U8287 (N_8287,N_172,N_2276);
nor U8288 (N_8288,N_751,N_4757);
nand U8289 (N_8289,N_1438,N_712);
nand U8290 (N_8290,N_2091,N_881);
nor U8291 (N_8291,N_512,N_2871);
nand U8292 (N_8292,N_2635,N_1360);
nor U8293 (N_8293,N_460,N_4608);
nor U8294 (N_8294,N_2063,N_4565);
nand U8295 (N_8295,N_4297,N_3905);
nor U8296 (N_8296,N_2432,N_4179);
nor U8297 (N_8297,N_2499,N_2334);
nor U8298 (N_8298,N_643,N_3731);
and U8299 (N_8299,N_4413,N_1829);
or U8300 (N_8300,N_351,N_2712);
nor U8301 (N_8301,N_1481,N_1620);
or U8302 (N_8302,N_3993,N_4483);
xnor U8303 (N_8303,N_2008,N_3323);
nor U8304 (N_8304,N_4401,N_4146);
nand U8305 (N_8305,N_1897,N_2796);
nand U8306 (N_8306,N_2887,N_4565);
or U8307 (N_8307,N_2492,N_630);
nand U8308 (N_8308,N_3782,N_246);
nor U8309 (N_8309,N_3136,N_1987);
nand U8310 (N_8310,N_4646,N_793);
nor U8311 (N_8311,N_1931,N_2799);
xor U8312 (N_8312,N_1479,N_4878);
nand U8313 (N_8313,N_787,N_3472);
xor U8314 (N_8314,N_1309,N_3177);
and U8315 (N_8315,N_492,N_395);
xnor U8316 (N_8316,N_4589,N_1956);
or U8317 (N_8317,N_4520,N_2743);
and U8318 (N_8318,N_3061,N_280);
nor U8319 (N_8319,N_2752,N_1861);
xor U8320 (N_8320,N_2993,N_1685);
nor U8321 (N_8321,N_1204,N_1711);
nand U8322 (N_8322,N_3065,N_2978);
or U8323 (N_8323,N_40,N_549);
nand U8324 (N_8324,N_4825,N_1764);
xnor U8325 (N_8325,N_2402,N_1126);
and U8326 (N_8326,N_4075,N_1794);
nand U8327 (N_8327,N_3651,N_4667);
and U8328 (N_8328,N_3331,N_3734);
xnor U8329 (N_8329,N_1263,N_1113);
and U8330 (N_8330,N_1560,N_2738);
nor U8331 (N_8331,N_3872,N_528);
nor U8332 (N_8332,N_2595,N_2211);
xnor U8333 (N_8333,N_2860,N_562);
and U8334 (N_8334,N_967,N_1125);
nand U8335 (N_8335,N_621,N_4180);
or U8336 (N_8336,N_1948,N_3355);
or U8337 (N_8337,N_620,N_3249);
and U8338 (N_8338,N_2683,N_1922);
or U8339 (N_8339,N_1811,N_2235);
and U8340 (N_8340,N_4744,N_2190);
xnor U8341 (N_8341,N_4545,N_3637);
or U8342 (N_8342,N_4978,N_2650);
or U8343 (N_8343,N_3176,N_1412);
or U8344 (N_8344,N_2424,N_1001);
nand U8345 (N_8345,N_3614,N_1450);
nor U8346 (N_8346,N_3494,N_2902);
nand U8347 (N_8347,N_1526,N_1360);
nor U8348 (N_8348,N_4129,N_57);
and U8349 (N_8349,N_3316,N_2975);
and U8350 (N_8350,N_3942,N_2431);
or U8351 (N_8351,N_898,N_384);
nand U8352 (N_8352,N_245,N_3789);
and U8353 (N_8353,N_3376,N_313);
and U8354 (N_8354,N_437,N_3904);
nor U8355 (N_8355,N_4879,N_1764);
and U8356 (N_8356,N_269,N_1176);
and U8357 (N_8357,N_3196,N_4795);
and U8358 (N_8358,N_719,N_2987);
nor U8359 (N_8359,N_807,N_3154);
or U8360 (N_8360,N_3001,N_3721);
or U8361 (N_8361,N_2696,N_438);
and U8362 (N_8362,N_68,N_3575);
nand U8363 (N_8363,N_3254,N_1044);
or U8364 (N_8364,N_1675,N_3594);
and U8365 (N_8365,N_2328,N_4227);
xor U8366 (N_8366,N_4530,N_2204);
and U8367 (N_8367,N_3698,N_4953);
and U8368 (N_8368,N_3070,N_2655);
and U8369 (N_8369,N_2802,N_4767);
xnor U8370 (N_8370,N_3366,N_4430);
and U8371 (N_8371,N_4998,N_1339);
or U8372 (N_8372,N_613,N_1561);
nor U8373 (N_8373,N_1714,N_399);
or U8374 (N_8374,N_1519,N_3566);
or U8375 (N_8375,N_660,N_883);
xnor U8376 (N_8376,N_31,N_2653);
or U8377 (N_8377,N_4998,N_2839);
nand U8378 (N_8378,N_3319,N_1933);
or U8379 (N_8379,N_3361,N_1467);
or U8380 (N_8380,N_11,N_4241);
and U8381 (N_8381,N_2551,N_4520);
nand U8382 (N_8382,N_2424,N_2252);
nand U8383 (N_8383,N_1037,N_2549);
xor U8384 (N_8384,N_4419,N_289);
nor U8385 (N_8385,N_3154,N_2366);
xnor U8386 (N_8386,N_1428,N_1200);
nor U8387 (N_8387,N_4530,N_398);
nor U8388 (N_8388,N_302,N_215);
nand U8389 (N_8389,N_4670,N_4586);
and U8390 (N_8390,N_2616,N_656);
or U8391 (N_8391,N_1230,N_4458);
and U8392 (N_8392,N_2012,N_1976);
or U8393 (N_8393,N_2942,N_3794);
or U8394 (N_8394,N_2965,N_1937);
nand U8395 (N_8395,N_798,N_4644);
or U8396 (N_8396,N_3905,N_2917);
or U8397 (N_8397,N_4760,N_34);
xor U8398 (N_8398,N_800,N_4450);
nor U8399 (N_8399,N_2097,N_3149);
and U8400 (N_8400,N_2636,N_1816);
nor U8401 (N_8401,N_3115,N_4285);
and U8402 (N_8402,N_417,N_4090);
nor U8403 (N_8403,N_4310,N_1100);
or U8404 (N_8404,N_1670,N_3482);
and U8405 (N_8405,N_4800,N_665);
nor U8406 (N_8406,N_1398,N_4458);
nor U8407 (N_8407,N_4342,N_4138);
and U8408 (N_8408,N_4010,N_1922);
and U8409 (N_8409,N_3413,N_1932);
or U8410 (N_8410,N_4617,N_4515);
and U8411 (N_8411,N_1108,N_2982);
nand U8412 (N_8412,N_2175,N_3319);
and U8413 (N_8413,N_1457,N_1427);
nand U8414 (N_8414,N_698,N_1121);
nor U8415 (N_8415,N_3639,N_281);
nand U8416 (N_8416,N_1918,N_1579);
or U8417 (N_8417,N_3872,N_2290);
nand U8418 (N_8418,N_4483,N_2823);
nand U8419 (N_8419,N_2843,N_2432);
or U8420 (N_8420,N_4937,N_4005);
nor U8421 (N_8421,N_1832,N_426);
and U8422 (N_8422,N_259,N_914);
nor U8423 (N_8423,N_1795,N_3335);
xor U8424 (N_8424,N_3987,N_982);
nand U8425 (N_8425,N_4797,N_2036);
and U8426 (N_8426,N_4970,N_1653);
nor U8427 (N_8427,N_4921,N_3565);
or U8428 (N_8428,N_3181,N_2016);
or U8429 (N_8429,N_3094,N_2834);
nor U8430 (N_8430,N_2310,N_4015);
or U8431 (N_8431,N_2251,N_395);
xnor U8432 (N_8432,N_2353,N_4374);
nand U8433 (N_8433,N_2131,N_3668);
or U8434 (N_8434,N_4725,N_2340);
nand U8435 (N_8435,N_4901,N_3598);
nor U8436 (N_8436,N_2227,N_1643);
and U8437 (N_8437,N_3604,N_2405);
nor U8438 (N_8438,N_2127,N_187);
or U8439 (N_8439,N_379,N_4670);
nand U8440 (N_8440,N_2297,N_3332);
nand U8441 (N_8441,N_2797,N_684);
xor U8442 (N_8442,N_1190,N_1684);
and U8443 (N_8443,N_697,N_1105);
or U8444 (N_8444,N_1075,N_313);
nor U8445 (N_8445,N_2970,N_3561);
and U8446 (N_8446,N_3685,N_20);
nand U8447 (N_8447,N_2999,N_376);
and U8448 (N_8448,N_695,N_3730);
nor U8449 (N_8449,N_3817,N_934);
nand U8450 (N_8450,N_4608,N_4249);
and U8451 (N_8451,N_2144,N_589);
nand U8452 (N_8452,N_1603,N_1994);
and U8453 (N_8453,N_1435,N_1203);
nor U8454 (N_8454,N_3530,N_2986);
nand U8455 (N_8455,N_910,N_907);
nor U8456 (N_8456,N_1765,N_4410);
nor U8457 (N_8457,N_3317,N_2791);
nor U8458 (N_8458,N_2742,N_2579);
nor U8459 (N_8459,N_4890,N_305);
nor U8460 (N_8460,N_2808,N_938);
nand U8461 (N_8461,N_2017,N_2347);
or U8462 (N_8462,N_1580,N_4293);
nor U8463 (N_8463,N_4603,N_2564);
nor U8464 (N_8464,N_3986,N_4909);
xor U8465 (N_8465,N_2890,N_3812);
nor U8466 (N_8466,N_1624,N_2578);
xnor U8467 (N_8467,N_4571,N_717);
nor U8468 (N_8468,N_4159,N_450);
xnor U8469 (N_8469,N_4586,N_1512);
nor U8470 (N_8470,N_2640,N_4219);
nand U8471 (N_8471,N_3039,N_1443);
nor U8472 (N_8472,N_899,N_2258);
nor U8473 (N_8473,N_2671,N_138);
nand U8474 (N_8474,N_94,N_1547);
nand U8475 (N_8475,N_661,N_4209);
nand U8476 (N_8476,N_2828,N_1113);
and U8477 (N_8477,N_3345,N_2976);
and U8478 (N_8478,N_3486,N_3576);
or U8479 (N_8479,N_2696,N_3492);
nand U8480 (N_8480,N_212,N_3873);
nor U8481 (N_8481,N_532,N_4765);
nand U8482 (N_8482,N_2637,N_3330);
nor U8483 (N_8483,N_4867,N_4751);
nand U8484 (N_8484,N_2987,N_1495);
and U8485 (N_8485,N_4245,N_4399);
or U8486 (N_8486,N_4538,N_4903);
or U8487 (N_8487,N_300,N_4302);
xor U8488 (N_8488,N_4508,N_1039);
or U8489 (N_8489,N_2769,N_3521);
or U8490 (N_8490,N_1346,N_3382);
or U8491 (N_8491,N_1230,N_4724);
nand U8492 (N_8492,N_1683,N_2183);
or U8493 (N_8493,N_2711,N_1626);
nor U8494 (N_8494,N_2261,N_3316);
nand U8495 (N_8495,N_4070,N_4437);
or U8496 (N_8496,N_4514,N_4626);
or U8497 (N_8497,N_3214,N_4091);
and U8498 (N_8498,N_4640,N_68);
or U8499 (N_8499,N_621,N_2854);
or U8500 (N_8500,N_903,N_2957);
or U8501 (N_8501,N_1011,N_3165);
nand U8502 (N_8502,N_2331,N_485);
or U8503 (N_8503,N_2296,N_1163);
or U8504 (N_8504,N_3598,N_922);
or U8505 (N_8505,N_622,N_4921);
and U8506 (N_8506,N_570,N_1375);
xor U8507 (N_8507,N_419,N_4334);
nor U8508 (N_8508,N_4817,N_1882);
or U8509 (N_8509,N_1288,N_3400);
and U8510 (N_8510,N_4928,N_4508);
nor U8511 (N_8511,N_4685,N_41);
nor U8512 (N_8512,N_1302,N_3990);
or U8513 (N_8513,N_2667,N_423);
nor U8514 (N_8514,N_2037,N_1028);
or U8515 (N_8515,N_3754,N_1682);
and U8516 (N_8516,N_568,N_2797);
or U8517 (N_8517,N_3774,N_2888);
or U8518 (N_8518,N_4863,N_1795);
or U8519 (N_8519,N_3006,N_1106);
nor U8520 (N_8520,N_4959,N_4319);
or U8521 (N_8521,N_4963,N_297);
nor U8522 (N_8522,N_273,N_31);
or U8523 (N_8523,N_2964,N_1759);
or U8524 (N_8524,N_1072,N_3054);
xor U8525 (N_8525,N_1279,N_481);
and U8526 (N_8526,N_990,N_2928);
nor U8527 (N_8527,N_572,N_1356);
xor U8528 (N_8528,N_1661,N_51);
or U8529 (N_8529,N_1711,N_2787);
nor U8530 (N_8530,N_4071,N_1892);
nand U8531 (N_8531,N_1284,N_4117);
or U8532 (N_8532,N_1183,N_4145);
or U8533 (N_8533,N_2967,N_850);
nor U8534 (N_8534,N_3230,N_1994);
or U8535 (N_8535,N_1563,N_1507);
and U8536 (N_8536,N_3710,N_4717);
nor U8537 (N_8537,N_3039,N_4539);
nor U8538 (N_8538,N_4224,N_1513);
nand U8539 (N_8539,N_1468,N_931);
nor U8540 (N_8540,N_4482,N_1602);
and U8541 (N_8541,N_4863,N_4088);
and U8542 (N_8542,N_100,N_2512);
nand U8543 (N_8543,N_1393,N_3035);
and U8544 (N_8544,N_4815,N_4511);
nand U8545 (N_8545,N_6,N_2724);
or U8546 (N_8546,N_1113,N_2303);
nor U8547 (N_8547,N_3104,N_4053);
nand U8548 (N_8548,N_4552,N_4527);
xor U8549 (N_8549,N_2826,N_505);
xnor U8550 (N_8550,N_1878,N_356);
xnor U8551 (N_8551,N_3056,N_4599);
and U8552 (N_8552,N_613,N_3133);
nand U8553 (N_8553,N_1136,N_2685);
or U8554 (N_8554,N_3453,N_4884);
nor U8555 (N_8555,N_1853,N_4615);
or U8556 (N_8556,N_3843,N_205);
xor U8557 (N_8557,N_4,N_4906);
or U8558 (N_8558,N_1582,N_2574);
nand U8559 (N_8559,N_1810,N_1755);
or U8560 (N_8560,N_4382,N_1210);
or U8561 (N_8561,N_2187,N_2726);
xnor U8562 (N_8562,N_2610,N_1416);
nand U8563 (N_8563,N_4067,N_737);
and U8564 (N_8564,N_821,N_2991);
nand U8565 (N_8565,N_3131,N_2633);
xnor U8566 (N_8566,N_1744,N_1481);
nand U8567 (N_8567,N_83,N_4658);
or U8568 (N_8568,N_2148,N_3462);
or U8569 (N_8569,N_3540,N_370);
or U8570 (N_8570,N_3474,N_217);
nor U8571 (N_8571,N_3423,N_93);
and U8572 (N_8572,N_4895,N_1240);
nand U8573 (N_8573,N_3375,N_3262);
nor U8574 (N_8574,N_1627,N_540);
and U8575 (N_8575,N_2086,N_1038);
and U8576 (N_8576,N_1517,N_2056);
or U8577 (N_8577,N_2538,N_2335);
nor U8578 (N_8578,N_1877,N_1826);
and U8579 (N_8579,N_3791,N_951);
or U8580 (N_8580,N_1106,N_210);
nand U8581 (N_8581,N_4705,N_2839);
nand U8582 (N_8582,N_4370,N_1139);
nor U8583 (N_8583,N_1254,N_2926);
nand U8584 (N_8584,N_636,N_2306);
nand U8585 (N_8585,N_848,N_2183);
or U8586 (N_8586,N_2461,N_1944);
nor U8587 (N_8587,N_969,N_2478);
and U8588 (N_8588,N_1119,N_3867);
and U8589 (N_8589,N_59,N_2718);
nand U8590 (N_8590,N_1534,N_4558);
nor U8591 (N_8591,N_1395,N_4051);
or U8592 (N_8592,N_4247,N_3326);
nor U8593 (N_8593,N_3809,N_3511);
nand U8594 (N_8594,N_2422,N_3355);
or U8595 (N_8595,N_2316,N_3533);
nand U8596 (N_8596,N_160,N_2926);
nor U8597 (N_8597,N_4236,N_1491);
nor U8598 (N_8598,N_2183,N_1585);
and U8599 (N_8599,N_3342,N_2322);
nand U8600 (N_8600,N_605,N_2549);
nand U8601 (N_8601,N_2350,N_3067);
and U8602 (N_8602,N_3132,N_4873);
nand U8603 (N_8603,N_1011,N_2033);
xor U8604 (N_8604,N_115,N_1672);
xnor U8605 (N_8605,N_161,N_3065);
nand U8606 (N_8606,N_1506,N_1618);
and U8607 (N_8607,N_2908,N_564);
or U8608 (N_8608,N_4300,N_1298);
nor U8609 (N_8609,N_4005,N_326);
nand U8610 (N_8610,N_968,N_543);
and U8611 (N_8611,N_1070,N_4671);
and U8612 (N_8612,N_67,N_4795);
or U8613 (N_8613,N_1538,N_3747);
nand U8614 (N_8614,N_431,N_4389);
xor U8615 (N_8615,N_2320,N_3163);
nand U8616 (N_8616,N_2121,N_1275);
nand U8617 (N_8617,N_857,N_61);
nand U8618 (N_8618,N_2557,N_1755);
nand U8619 (N_8619,N_1548,N_2200);
and U8620 (N_8620,N_2071,N_935);
xnor U8621 (N_8621,N_2280,N_2055);
xor U8622 (N_8622,N_3653,N_4357);
nand U8623 (N_8623,N_2967,N_2997);
nand U8624 (N_8624,N_709,N_470);
and U8625 (N_8625,N_3244,N_1633);
nand U8626 (N_8626,N_2607,N_326);
nor U8627 (N_8627,N_225,N_219);
or U8628 (N_8628,N_58,N_2222);
nor U8629 (N_8629,N_1095,N_3998);
or U8630 (N_8630,N_2086,N_2857);
and U8631 (N_8631,N_3655,N_786);
xor U8632 (N_8632,N_4786,N_4787);
xnor U8633 (N_8633,N_469,N_4132);
and U8634 (N_8634,N_2198,N_4246);
or U8635 (N_8635,N_2892,N_2237);
nand U8636 (N_8636,N_4922,N_1661);
nand U8637 (N_8637,N_451,N_2961);
or U8638 (N_8638,N_1055,N_106);
or U8639 (N_8639,N_3125,N_904);
and U8640 (N_8640,N_684,N_3358);
or U8641 (N_8641,N_4742,N_2201);
nand U8642 (N_8642,N_3515,N_2214);
nor U8643 (N_8643,N_4244,N_1920);
and U8644 (N_8644,N_2542,N_1225);
or U8645 (N_8645,N_2551,N_891);
nor U8646 (N_8646,N_1764,N_2570);
and U8647 (N_8647,N_457,N_3780);
or U8648 (N_8648,N_173,N_4527);
nor U8649 (N_8649,N_64,N_373);
and U8650 (N_8650,N_2681,N_1988);
nand U8651 (N_8651,N_3653,N_1282);
or U8652 (N_8652,N_2843,N_1213);
or U8653 (N_8653,N_2668,N_1413);
nand U8654 (N_8654,N_37,N_4424);
and U8655 (N_8655,N_2691,N_2011);
nand U8656 (N_8656,N_4271,N_4085);
and U8657 (N_8657,N_2518,N_67);
nor U8658 (N_8658,N_4308,N_530);
and U8659 (N_8659,N_3113,N_3047);
and U8660 (N_8660,N_4378,N_911);
or U8661 (N_8661,N_409,N_4594);
or U8662 (N_8662,N_3403,N_485);
nand U8663 (N_8663,N_2742,N_4736);
nand U8664 (N_8664,N_4606,N_2853);
nor U8665 (N_8665,N_2555,N_1761);
nor U8666 (N_8666,N_3550,N_3572);
nor U8667 (N_8667,N_876,N_1354);
nor U8668 (N_8668,N_4340,N_4438);
or U8669 (N_8669,N_2885,N_496);
nor U8670 (N_8670,N_1603,N_2054);
nand U8671 (N_8671,N_3836,N_4124);
nor U8672 (N_8672,N_3739,N_1599);
or U8673 (N_8673,N_4516,N_2047);
xor U8674 (N_8674,N_650,N_3610);
and U8675 (N_8675,N_2890,N_224);
nor U8676 (N_8676,N_2101,N_1870);
or U8677 (N_8677,N_3784,N_233);
and U8678 (N_8678,N_1589,N_516);
nand U8679 (N_8679,N_2719,N_3026);
or U8680 (N_8680,N_4591,N_3486);
xor U8681 (N_8681,N_1190,N_4782);
and U8682 (N_8682,N_1576,N_4137);
and U8683 (N_8683,N_610,N_4995);
and U8684 (N_8684,N_1405,N_4602);
nand U8685 (N_8685,N_2844,N_1206);
nand U8686 (N_8686,N_400,N_1441);
xor U8687 (N_8687,N_3891,N_3492);
or U8688 (N_8688,N_4590,N_3439);
and U8689 (N_8689,N_3051,N_348);
or U8690 (N_8690,N_444,N_2049);
or U8691 (N_8691,N_443,N_3462);
nand U8692 (N_8692,N_4244,N_800);
and U8693 (N_8693,N_418,N_1059);
nand U8694 (N_8694,N_2406,N_3017);
or U8695 (N_8695,N_2636,N_2050);
nand U8696 (N_8696,N_3957,N_306);
nor U8697 (N_8697,N_3612,N_884);
and U8698 (N_8698,N_4027,N_1286);
nor U8699 (N_8699,N_2434,N_51);
nand U8700 (N_8700,N_2593,N_2703);
or U8701 (N_8701,N_347,N_1078);
and U8702 (N_8702,N_1172,N_2038);
nor U8703 (N_8703,N_3891,N_605);
xnor U8704 (N_8704,N_1653,N_3309);
nand U8705 (N_8705,N_228,N_2646);
nor U8706 (N_8706,N_3858,N_2981);
and U8707 (N_8707,N_2130,N_2689);
and U8708 (N_8708,N_2952,N_2731);
nand U8709 (N_8709,N_514,N_2892);
xor U8710 (N_8710,N_2618,N_4079);
nand U8711 (N_8711,N_4699,N_3536);
nand U8712 (N_8712,N_3929,N_2890);
or U8713 (N_8713,N_81,N_4545);
and U8714 (N_8714,N_2813,N_4092);
nor U8715 (N_8715,N_2883,N_3826);
or U8716 (N_8716,N_2000,N_3999);
or U8717 (N_8717,N_3768,N_3228);
nand U8718 (N_8718,N_1756,N_3043);
and U8719 (N_8719,N_2674,N_2769);
nor U8720 (N_8720,N_2845,N_3776);
xnor U8721 (N_8721,N_4000,N_55);
and U8722 (N_8722,N_1357,N_3464);
or U8723 (N_8723,N_82,N_577);
or U8724 (N_8724,N_1419,N_2921);
nand U8725 (N_8725,N_1459,N_217);
nor U8726 (N_8726,N_2921,N_515);
or U8727 (N_8727,N_2687,N_4269);
nand U8728 (N_8728,N_1293,N_40);
and U8729 (N_8729,N_4195,N_2250);
and U8730 (N_8730,N_1091,N_2240);
nor U8731 (N_8731,N_1440,N_170);
nand U8732 (N_8732,N_2505,N_1497);
nand U8733 (N_8733,N_3525,N_4629);
and U8734 (N_8734,N_4559,N_3874);
or U8735 (N_8735,N_4712,N_4406);
and U8736 (N_8736,N_1305,N_2355);
nor U8737 (N_8737,N_4457,N_4072);
or U8738 (N_8738,N_2716,N_1617);
or U8739 (N_8739,N_1289,N_1454);
or U8740 (N_8740,N_772,N_3731);
or U8741 (N_8741,N_601,N_1749);
xor U8742 (N_8742,N_2029,N_2073);
xor U8743 (N_8743,N_1674,N_4346);
or U8744 (N_8744,N_2806,N_4899);
nand U8745 (N_8745,N_454,N_1934);
and U8746 (N_8746,N_2117,N_660);
or U8747 (N_8747,N_3531,N_2059);
and U8748 (N_8748,N_2509,N_3865);
nand U8749 (N_8749,N_3118,N_2921);
nor U8750 (N_8750,N_1041,N_3721);
nand U8751 (N_8751,N_732,N_2403);
or U8752 (N_8752,N_4584,N_2658);
or U8753 (N_8753,N_2993,N_2061);
nand U8754 (N_8754,N_1609,N_2356);
xnor U8755 (N_8755,N_4802,N_1250);
or U8756 (N_8756,N_3934,N_2632);
or U8757 (N_8757,N_1107,N_2891);
or U8758 (N_8758,N_2050,N_1502);
nor U8759 (N_8759,N_1541,N_2431);
and U8760 (N_8760,N_2177,N_4140);
and U8761 (N_8761,N_1072,N_4169);
and U8762 (N_8762,N_509,N_633);
xnor U8763 (N_8763,N_4228,N_1475);
and U8764 (N_8764,N_3157,N_1877);
nor U8765 (N_8765,N_3010,N_3577);
nor U8766 (N_8766,N_1840,N_347);
and U8767 (N_8767,N_787,N_4407);
and U8768 (N_8768,N_2201,N_2996);
and U8769 (N_8769,N_3446,N_3719);
or U8770 (N_8770,N_3598,N_32);
or U8771 (N_8771,N_3403,N_1333);
nand U8772 (N_8772,N_3614,N_1112);
and U8773 (N_8773,N_1800,N_2207);
nor U8774 (N_8774,N_3211,N_1391);
nand U8775 (N_8775,N_233,N_1431);
and U8776 (N_8776,N_2634,N_1845);
nand U8777 (N_8777,N_2812,N_3181);
or U8778 (N_8778,N_3242,N_1267);
nor U8779 (N_8779,N_2510,N_2840);
nor U8780 (N_8780,N_4374,N_1494);
and U8781 (N_8781,N_4181,N_4619);
nor U8782 (N_8782,N_1546,N_2652);
and U8783 (N_8783,N_1710,N_492);
or U8784 (N_8784,N_1740,N_581);
nor U8785 (N_8785,N_2072,N_4834);
and U8786 (N_8786,N_3744,N_3435);
xnor U8787 (N_8787,N_2586,N_3802);
or U8788 (N_8788,N_3988,N_2126);
nor U8789 (N_8789,N_1401,N_2950);
or U8790 (N_8790,N_841,N_398);
nor U8791 (N_8791,N_426,N_1980);
xor U8792 (N_8792,N_2665,N_3603);
nand U8793 (N_8793,N_2119,N_4574);
nand U8794 (N_8794,N_3128,N_2878);
nand U8795 (N_8795,N_2949,N_4848);
or U8796 (N_8796,N_2836,N_235);
or U8797 (N_8797,N_3304,N_430);
or U8798 (N_8798,N_3821,N_555);
nor U8799 (N_8799,N_1405,N_3185);
and U8800 (N_8800,N_4335,N_4504);
and U8801 (N_8801,N_3698,N_1443);
nor U8802 (N_8802,N_3021,N_1996);
nand U8803 (N_8803,N_4825,N_1954);
and U8804 (N_8804,N_3696,N_705);
nor U8805 (N_8805,N_86,N_721);
nor U8806 (N_8806,N_4116,N_4436);
or U8807 (N_8807,N_3325,N_1118);
xor U8808 (N_8808,N_662,N_4183);
and U8809 (N_8809,N_4862,N_4186);
nor U8810 (N_8810,N_4739,N_2408);
or U8811 (N_8811,N_2486,N_126);
and U8812 (N_8812,N_499,N_4788);
nor U8813 (N_8813,N_619,N_2862);
nor U8814 (N_8814,N_1142,N_1308);
nor U8815 (N_8815,N_2513,N_413);
and U8816 (N_8816,N_3136,N_1672);
or U8817 (N_8817,N_1564,N_2082);
nand U8818 (N_8818,N_1634,N_2689);
xor U8819 (N_8819,N_4778,N_1623);
and U8820 (N_8820,N_1781,N_3654);
or U8821 (N_8821,N_1804,N_3933);
xor U8822 (N_8822,N_382,N_3670);
and U8823 (N_8823,N_2165,N_3818);
nand U8824 (N_8824,N_27,N_598);
xor U8825 (N_8825,N_4391,N_4125);
nor U8826 (N_8826,N_2778,N_51);
nand U8827 (N_8827,N_3648,N_2714);
and U8828 (N_8828,N_3715,N_2592);
and U8829 (N_8829,N_2881,N_2117);
xor U8830 (N_8830,N_503,N_932);
nand U8831 (N_8831,N_200,N_1651);
nand U8832 (N_8832,N_298,N_1286);
xor U8833 (N_8833,N_682,N_3241);
or U8834 (N_8834,N_207,N_1102);
nor U8835 (N_8835,N_2443,N_4576);
and U8836 (N_8836,N_3754,N_1586);
nor U8837 (N_8837,N_3506,N_4782);
nand U8838 (N_8838,N_4523,N_567);
nor U8839 (N_8839,N_4742,N_1501);
nor U8840 (N_8840,N_2116,N_4271);
nand U8841 (N_8841,N_4955,N_2090);
nor U8842 (N_8842,N_21,N_715);
nand U8843 (N_8843,N_4208,N_4096);
nor U8844 (N_8844,N_1812,N_1617);
nor U8845 (N_8845,N_48,N_4759);
xnor U8846 (N_8846,N_1328,N_4644);
nor U8847 (N_8847,N_773,N_313);
nand U8848 (N_8848,N_4078,N_4631);
xnor U8849 (N_8849,N_4312,N_1652);
nand U8850 (N_8850,N_3782,N_3665);
and U8851 (N_8851,N_4995,N_2237);
nand U8852 (N_8852,N_4569,N_983);
nor U8853 (N_8853,N_3254,N_2637);
nor U8854 (N_8854,N_1863,N_1582);
xnor U8855 (N_8855,N_1518,N_3832);
or U8856 (N_8856,N_2714,N_2295);
and U8857 (N_8857,N_4971,N_4926);
nand U8858 (N_8858,N_3669,N_1987);
or U8859 (N_8859,N_3867,N_4540);
and U8860 (N_8860,N_586,N_1604);
nor U8861 (N_8861,N_2372,N_1510);
or U8862 (N_8862,N_139,N_778);
or U8863 (N_8863,N_697,N_4571);
or U8864 (N_8864,N_1092,N_3842);
and U8865 (N_8865,N_4740,N_3286);
or U8866 (N_8866,N_4322,N_353);
nor U8867 (N_8867,N_1537,N_3419);
or U8868 (N_8868,N_3731,N_4436);
or U8869 (N_8869,N_741,N_2293);
xor U8870 (N_8870,N_2059,N_393);
nor U8871 (N_8871,N_1132,N_338);
and U8872 (N_8872,N_1665,N_3971);
xor U8873 (N_8873,N_2070,N_2314);
nor U8874 (N_8874,N_225,N_2962);
or U8875 (N_8875,N_2489,N_2343);
and U8876 (N_8876,N_513,N_668);
nor U8877 (N_8877,N_566,N_3467);
or U8878 (N_8878,N_536,N_4331);
and U8879 (N_8879,N_4079,N_2506);
xor U8880 (N_8880,N_4316,N_4225);
nor U8881 (N_8881,N_1624,N_3036);
or U8882 (N_8882,N_1977,N_2485);
nor U8883 (N_8883,N_2133,N_2191);
nand U8884 (N_8884,N_372,N_168);
or U8885 (N_8885,N_1683,N_2409);
and U8886 (N_8886,N_2232,N_1251);
or U8887 (N_8887,N_2129,N_4411);
or U8888 (N_8888,N_1957,N_1953);
nor U8889 (N_8889,N_4539,N_2445);
or U8890 (N_8890,N_2027,N_1370);
or U8891 (N_8891,N_3100,N_4889);
xor U8892 (N_8892,N_819,N_4031);
nor U8893 (N_8893,N_774,N_2354);
nor U8894 (N_8894,N_733,N_3287);
nor U8895 (N_8895,N_4150,N_1000);
and U8896 (N_8896,N_1940,N_4419);
nand U8897 (N_8897,N_266,N_2600);
xnor U8898 (N_8898,N_4494,N_3979);
or U8899 (N_8899,N_4503,N_1908);
or U8900 (N_8900,N_279,N_473);
and U8901 (N_8901,N_1962,N_1331);
or U8902 (N_8902,N_688,N_4232);
nand U8903 (N_8903,N_4443,N_4118);
xnor U8904 (N_8904,N_2768,N_4496);
or U8905 (N_8905,N_368,N_1383);
nor U8906 (N_8906,N_4704,N_328);
nand U8907 (N_8907,N_3764,N_4993);
and U8908 (N_8908,N_3916,N_2818);
nand U8909 (N_8909,N_4656,N_4537);
nor U8910 (N_8910,N_4169,N_2361);
nand U8911 (N_8911,N_2653,N_1764);
nand U8912 (N_8912,N_3927,N_262);
xnor U8913 (N_8913,N_2839,N_532);
or U8914 (N_8914,N_3014,N_4408);
or U8915 (N_8915,N_2720,N_3799);
and U8916 (N_8916,N_3663,N_2440);
and U8917 (N_8917,N_4202,N_2333);
or U8918 (N_8918,N_1134,N_4933);
nor U8919 (N_8919,N_442,N_3336);
nor U8920 (N_8920,N_994,N_1944);
or U8921 (N_8921,N_17,N_4123);
or U8922 (N_8922,N_4516,N_1288);
nand U8923 (N_8923,N_4441,N_2200);
nand U8924 (N_8924,N_2976,N_1246);
nor U8925 (N_8925,N_2088,N_1036);
xnor U8926 (N_8926,N_2065,N_4147);
nand U8927 (N_8927,N_2753,N_752);
and U8928 (N_8928,N_3414,N_2589);
and U8929 (N_8929,N_3988,N_3197);
or U8930 (N_8930,N_2488,N_2650);
and U8931 (N_8931,N_3008,N_3985);
or U8932 (N_8932,N_1232,N_269);
and U8933 (N_8933,N_2036,N_1920);
and U8934 (N_8934,N_2471,N_391);
nor U8935 (N_8935,N_3273,N_4362);
nor U8936 (N_8936,N_2892,N_2042);
xor U8937 (N_8937,N_4111,N_3225);
nor U8938 (N_8938,N_2204,N_1379);
nor U8939 (N_8939,N_1896,N_627);
nand U8940 (N_8940,N_1147,N_4506);
nor U8941 (N_8941,N_1887,N_3783);
or U8942 (N_8942,N_2028,N_3374);
and U8943 (N_8943,N_1491,N_1773);
or U8944 (N_8944,N_2186,N_2320);
and U8945 (N_8945,N_495,N_2126);
nand U8946 (N_8946,N_1829,N_2363);
nor U8947 (N_8947,N_3680,N_4852);
nor U8948 (N_8948,N_1894,N_346);
nand U8949 (N_8949,N_3974,N_56);
and U8950 (N_8950,N_358,N_3025);
and U8951 (N_8951,N_1225,N_3403);
nand U8952 (N_8952,N_4086,N_2150);
and U8953 (N_8953,N_2687,N_716);
nor U8954 (N_8954,N_4386,N_830);
or U8955 (N_8955,N_3181,N_191);
nand U8956 (N_8956,N_2444,N_3120);
xnor U8957 (N_8957,N_4094,N_4851);
nor U8958 (N_8958,N_2342,N_1558);
xor U8959 (N_8959,N_922,N_4647);
nand U8960 (N_8960,N_1579,N_431);
or U8961 (N_8961,N_2994,N_1070);
xnor U8962 (N_8962,N_276,N_3924);
xnor U8963 (N_8963,N_959,N_3858);
and U8964 (N_8964,N_2127,N_2963);
nor U8965 (N_8965,N_4064,N_4470);
nor U8966 (N_8966,N_280,N_1897);
xor U8967 (N_8967,N_1726,N_3923);
nor U8968 (N_8968,N_257,N_1129);
nand U8969 (N_8969,N_4368,N_1260);
and U8970 (N_8970,N_311,N_4521);
nor U8971 (N_8971,N_103,N_4459);
or U8972 (N_8972,N_1591,N_960);
or U8973 (N_8973,N_2176,N_139);
xnor U8974 (N_8974,N_2932,N_4868);
nand U8975 (N_8975,N_4799,N_3985);
nand U8976 (N_8976,N_2516,N_1501);
or U8977 (N_8977,N_3348,N_23);
xnor U8978 (N_8978,N_3426,N_4114);
or U8979 (N_8979,N_3487,N_1777);
or U8980 (N_8980,N_785,N_3402);
and U8981 (N_8981,N_4254,N_3389);
or U8982 (N_8982,N_3930,N_4144);
and U8983 (N_8983,N_3074,N_1533);
and U8984 (N_8984,N_172,N_3130);
xor U8985 (N_8985,N_1469,N_2783);
nor U8986 (N_8986,N_2055,N_1734);
xnor U8987 (N_8987,N_1855,N_4557);
nand U8988 (N_8988,N_643,N_772);
or U8989 (N_8989,N_1163,N_672);
xor U8990 (N_8990,N_2412,N_2340);
or U8991 (N_8991,N_4210,N_1986);
and U8992 (N_8992,N_606,N_475);
nand U8993 (N_8993,N_3546,N_2715);
or U8994 (N_8994,N_4657,N_1842);
nor U8995 (N_8995,N_3873,N_360);
and U8996 (N_8996,N_60,N_3067);
xor U8997 (N_8997,N_885,N_1637);
nand U8998 (N_8998,N_4839,N_310);
nor U8999 (N_8999,N_3578,N_2702);
nor U9000 (N_9000,N_4179,N_326);
and U9001 (N_9001,N_3761,N_946);
or U9002 (N_9002,N_498,N_2614);
nor U9003 (N_9003,N_773,N_3221);
or U9004 (N_9004,N_2865,N_4496);
nand U9005 (N_9005,N_407,N_4401);
nor U9006 (N_9006,N_4698,N_1694);
xor U9007 (N_9007,N_375,N_4640);
nand U9008 (N_9008,N_4956,N_3763);
nand U9009 (N_9009,N_3519,N_1942);
nor U9010 (N_9010,N_1524,N_2964);
nor U9011 (N_9011,N_4965,N_1813);
and U9012 (N_9012,N_2858,N_1000);
xnor U9013 (N_9013,N_4124,N_3317);
and U9014 (N_9014,N_1516,N_3314);
xor U9015 (N_9015,N_524,N_3790);
and U9016 (N_9016,N_2041,N_936);
nand U9017 (N_9017,N_4681,N_4169);
and U9018 (N_9018,N_901,N_2113);
and U9019 (N_9019,N_4493,N_1489);
xnor U9020 (N_9020,N_336,N_3318);
nor U9021 (N_9021,N_2225,N_1351);
nor U9022 (N_9022,N_2101,N_543);
nand U9023 (N_9023,N_3926,N_4147);
nor U9024 (N_9024,N_2402,N_3665);
or U9025 (N_9025,N_1644,N_4419);
nand U9026 (N_9026,N_3959,N_2623);
xnor U9027 (N_9027,N_3704,N_915);
or U9028 (N_9028,N_3810,N_4857);
nand U9029 (N_9029,N_1821,N_4275);
nand U9030 (N_9030,N_71,N_4840);
or U9031 (N_9031,N_1930,N_1452);
nor U9032 (N_9032,N_3452,N_4773);
nand U9033 (N_9033,N_1197,N_4640);
nor U9034 (N_9034,N_684,N_4033);
and U9035 (N_9035,N_806,N_4649);
nand U9036 (N_9036,N_2371,N_325);
nand U9037 (N_9037,N_4737,N_3178);
or U9038 (N_9038,N_683,N_4591);
and U9039 (N_9039,N_218,N_1429);
nand U9040 (N_9040,N_741,N_4698);
nand U9041 (N_9041,N_512,N_4318);
and U9042 (N_9042,N_4547,N_3176);
and U9043 (N_9043,N_2306,N_2572);
nand U9044 (N_9044,N_402,N_688);
xnor U9045 (N_9045,N_1190,N_3606);
nand U9046 (N_9046,N_579,N_1193);
and U9047 (N_9047,N_492,N_1528);
nand U9048 (N_9048,N_4538,N_1418);
nand U9049 (N_9049,N_2159,N_3062);
or U9050 (N_9050,N_4432,N_3720);
nor U9051 (N_9051,N_3087,N_2733);
nand U9052 (N_9052,N_1197,N_2089);
xor U9053 (N_9053,N_3457,N_278);
nor U9054 (N_9054,N_750,N_1202);
nor U9055 (N_9055,N_3679,N_4135);
nor U9056 (N_9056,N_1435,N_3133);
and U9057 (N_9057,N_156,N_3826);
or U9058 (N_9058,N_1120,N_4384);
nor U9059 (N_9059,N_1846,N_2790);
nand U9060 (N_9060,N_987,N_4795);
or U9061 (N_9061,N_2581,N_2386);
and U9062 (N_9062,N_4378,N_3732);
and U9063 (N_9063,N_4029,N_3695);
or U9064 (N_9064,N_2885,N_2866);
nor U9065 (N_9065,N_1302,N_3791);
nor U9066 (N_9066,N_4403,N_1580);
or U9067 (N_9067,N_277,N_4585);
or U9068 (N_9068,N_674,N_2351);
or U9069 (N_9069,N_1017,N_4327);
or U9070 (N_9070,N_448,N_3419);
and U9071 (N_9071,N_1589,N_3380);
nand U9072 (N_9072,N_4577,N_3521);
or U9073 (N_9073,N_3627,N_2710);
and U9074 (N_9074,N_1161,N_4208);
or U9075 (N_9075,N_1507,N_2815);
nor U9076 (N_9076,N_3156,N_2831);
and U9077 (N_9077,N_3768,N_74);
and U9078 (N_9078,N_1383,N_1370);
xnor U9079 (N_9079,N_2427,N_1596);
and U9080 (N_9080,N_1602,N_2595);
nor U9081 (N_9081,N_2987,N_3253);
or U9082 (N_9082,N_878,N_2854);
or U9083 (N_9083,N_2707,N_4723);
or U9084 (N_9084,N_3242,N_2900);
nor U9085 (N_9085,N_3667,N_3237);
xnor U9086 (N_9086,N_4700,N_2504);
nor U9087 (N_9087,N_1907,N_1643);
nor U9088 (N_9088,N_2465,N_2359);
and U9089 (N_9089,N_492,N_2965);
nand U9090 (N_9090,N_491,N_3472);
or U9091 (N_9091,N_4691,N_3485);
and U9092 (N_9092,N_1462,N_3030);
xor U9093 (N_9093,N_902,N_1626);
nand U9094 (N_9094,N_519,N_1232);
nor U9095 (N_9095,N_3071,N_581);
nor U9096 (N_9096,N_3136,N_4429);
nand U9097 (N_9097,N_1962,N_4802);
and U9098 (N_9098,N_4401,N_1675);
and U9099 (N_9099,N_2747,N_2533);
nor U9100 (N_9100,N_4979,N_2939);
nand U9101 (N_9101,N_2891,N_577);
and U9102 (N_9102,N_280,N_3796);
nand U9103 (N_9103,N_1442,N_783);
or U9104 (N_9104,N_4052,N_1137);
or U9105 (N_9105,N_2866,N_2183);
nor U9106 (N_9106,N_2978,N_4892);
or U9107 (N_9107,N_4729,N_3602);
and U9108 (N_9108,N_817,N_2726);
and U9109 (N_9109,N_3634,N_2011);
nand U9110 (N_9110,N_1658,N_2956);
nor U9111 (N_9111,N_717,N_192);
and U9112 (N_9112,N_1317,N_1462);
xor U9113 (N_9113,N_872,N_4303);
nor U9114 (N_9114,N_1474,N_120);
or U9115 (N_9115,N_3935,N_3620);
nand U9116 (N_9116,N_4118,N_2998);
nor U9117 (N_9117,N_3638,N_1780);
and U9118 (N_9118,N_3597,N_2479);
xnor U9119 (N_9119,N_4722,N_2259);
xor U9120 (N_9120,N_1165,N_1562);
or U9121 (N_9121,N_1933,N_214);
or U9122 (N_9122,N_3118,N_2322);
or U9123 (N_9123,N_1098,N_914);
nor U9124 (N_9124,N_1571,N_187);
xnor U9125 (N_9125,N_4552,N_1430);
and U9126 (N_9126,N_1452,N_4711);
nor U9127 (N_9127,N_4881,N_1970);
nor U9128 (N_9128,N_4388,N_1418);
nand U9129 (N_9129,N_3349,N_2242);
nor U9130 (N_9130,N_4728,N_4740);
nor U9131 (N_9131,N_3280,N_1453);
nand U9132 (N_9132,N_1497,N_445);
nand U9133 (N_9133,N_956,N_3693);
nor U9134 (N_9134,N_4763,N_216);
nand U9135 (N_9135,N_63,N_2479);
or U9136 (N_9136,N_3065,N_1912);
nor U9137 (N_9137,N_195,N_1805);
or U9138 (N_9138,N_550,N_2435);
nand U9139 (N_9139,N_4463,N_1293);
and U9140 (N_9140,N_454,N_3214);
and U9141 (N_9141,N_42,N_2955);
and U9142 (N_9142,N_4762,N_3027);
nand U9143 (N_9143,N_176,N_3567);
or U9144 (N_9144,N_1685,N_4188);
nand U9145 (N_9145,N_3815,N_2205);
nor U9146 (N_9146,N_4838,N_606);
or U9147 (N_9147,N_4348,N_723);
nor U9148 (N_9148,N_2678,N_30);
nand U9149 (N_9149,N_4732,N_2416);
and U9150 (N_9150,N_3436,N_837);
and U9151 (N_9151,N_891,N_3442);
and U9152 (N_9152,N_268,N_477);
nand U9153 (N_9153,N_3278,N_2853);
or U9154 (N_9154,N_857,N_4089);
nand U9155 (N_9155,N_255,N_14);
nor U9156 (N_9156,N_1954,N_3682);
nand U9157 (N_9157,N_1242,N_4951);
xor U9158 (N_9158,N_4927,N_3028);
or U9159 (N_9159,N_3364,N_3303);
or U9160 (N_9160,N_4171,N_381);
and U9161 (N_9161,N_1356,N_1322);
nand U9162 (N_9162,N_2008,N_1674);
and U9163 (N_9163,N_4460,N_1413);
and U9164 (N_9164,N_2153,N_2653);
and U9165 (N_9165,N_4202,N_1849);
nand U9166 (N_9166,N_3847,N_3555);
and U9167 (N_9167,N_1788,N_3545);
nor U9168 (N_9168,N_898,N_429);
or U9169 (N_9169,N_3022,N_3079);
and U9170 (N_9170,N_1843,N_2134);
or U9171 (N_9171,N_1278,N_2433);
and U9172 (N_9172,N_3237,N_1971);
or U9173 (N_9173,N_121,N_670);
and U9174 (N_9174,N_2740,N_2645);
nand U9175 (N_9175,N_1097,N_1216);
nand U9176 (N_9176,N_1493,N_888);
and U9177 (N_9177,N_4985,N_4946);
or U9178 (N_9178,N_3987,N_2633);
or U9179 (N_9179,N_381,N_4775);
or U9180 (N_9180,N_3164,N_3721);
or U9181 (N_9181,N_854,N_3480);
or U9182 (N_9182,N_4019,N_3150);
or U9183 (N_9183,N_2094,N_3599);
nor U9184 (N_9184,N_2736,N_1812);
or U9185 (N_9185,N_3423,N_525);
or U9186 (N_9186,N_2942,N_695);
xnor U9187 (N_9187,N_2908,N_3533);
and U9188 (N_9188,N_877,N_1615);
xnor U9189 (N_9189,N_4863,N_1541);
nand U9190 (N_9190,N_1148,N_409);
or U9191 (N_9191,N_103,N_2417);
and U9192 (N_9192,N_2733,N_3669);
or U9193 (N_9193,N_896,N_3563);
nor U9194 (N_9194,N_28,N_520);
or U9195 (N_9195,N_180,N_3777);
nand U9196 (N_9196,N_1697,N_4069);
or U9197 (N_9197,N_1364,N_4135);
and U9198 (N_9198,N_3656,N_1430);
or U9199 (N_9199,N_2344,N_3298);
nor U9200 (N_9200,N_4480,N_1519);
nand U9201 (N_9201,N_2989,N_4639);
or U9202 (N_9202,N_770,N_2114);
or U9203 (N_9203,N_3485,N_3853);
xnor U9204 (N_9204,N_2567,N_4235);
nor U9205 (N_9205,N_2684,N_4174);
nor U9206 (N_9206,N_364,N_2817);
and U9207 (N_9207,N_4221,N_4789);
or U9208 (N_9208,N_4558,N_3773);
nor U9209 (N_9209,N_1947,N_1685);
or U9210 (N_9210,N_3395,N_1204);
nor U9211 (N_9211,N_1010,N_887);
nand U9212 (N_9212,N_2992,N_4303);
or U9213 (N_9213,N_4086,N_1455);
nor U9214 (N_9214,N_814,N_201);
or U9215 (N_9215,N_1602,N_1237);
nor U9216 (N_9216,N_4027,N_1937);
nor U9217 (N_9217,N_1167,N_1439);
and U9218 (N_9218,N_3559,N_3317);
nor U9219 (N_9219,N_4606,N_253);
and U9220 (N_9220,N_2222,N_2597);
or U9221 (N_9221,N_4147,N_3414);
xnor U9222 (N_9222,N_1256,N_2050);
nand U9223 (N_9223,N_3055,N_501);
nand U9224 (N_9224,N_175,N_3823);
or U9225 (N_9225,N_1931,N_3860);
nand U9226 (N_9226,N_4278,N_210);
nand U9227 (N_9227,N_4041,N_3883);
or U9228 (N_9228,N_2771,N_3796);
and U9229 (N_9229,N_1160,N_4049);
nand U9230 (N_9230,N_3704,N_2538);
nand U9231 (N_9231,N_3288,N_4438);
nor U9232 (N_9232,N_450,N_1038);
or U9233 (N_9233,N_578,N_4467);
or U9234 (N_9234,N_4087,N_4651);
nand U9235 (N_9235,N_4905,N_113);
or U9236 (N_9236,N_2815,N_757);
nand U9237 (N_9237,N_4622,N_3971);
or U9238 (N_9238,N_2888,N_3902);
nand U9239 (N_9239,N_434,N_1306);
nand U9240 (N_9240,N_238,N_2367);
nand U9241 (N_9241,N_1393,N_52);
nand U9242 (N_9242,N_3489,N_1542);
or U9243 (N_9243,N_874,N_3816);
or U9244 (N_9244,N_886,N_2641);
xor U9245 (N_9245,N_739,N_3223);
nor U9246 (N_9246,N_4949,N_4887);
nand U9247 (N_9247,N_4133,N_2345);
nor U9248 (N_9248,N_2633,N_3201);
nor U9249 (N_9249,N_904,N_4656);
or U9250 (N_9250,N_1338,N_1274);
or U9251 (N_9251,N_2593,N_3818);
nor U9252 (N_9252,N_1383,N_2208);
or U9253 (N_9253,N_70,N_1239);
or U9254 (N_9254,N_1822,N_4504);
or U9255 (N_9255,N_244,N_10);
or U9256 (N_9256,N_3915,N_584);
or U9257 (N_9257,N_4760,N_4375);
and U9258 (N_9258,N_1901,N_2256);
xnor U9259 (N_9259,N_1002,N_3946);
nand U9260 (N_9260,N_3556,N_1082);
or U9261 (N_9261,N_3693,N_4353);
and U9262 (N_9262,N_3172,N_4644);
nor U9263 (N_9263,N_3694,N_3785);
nand U9264 (N_9264,N_1585,N_1376);
xnor U9265 (N_9265,N_2236,N_1706);
and U9266 (N_9266,N_3386,N_4549);
nor U9267 (N_9267,N_761,N_1599);
nand U9268 (N_9268,N_1064,N_2596);
and U9269 (N_9269,N_390,N_1021);
nand U9270 (N_9270,N_610,N_3790);
and U9271 (N_9271,N_4695,N_2740);
and U9272 (N_9272,N_3320,N_1807);
nor U9273 (N_9273,N_4112,N_4866);
and U9274 (N_9274,N_4992,N_836);
nor U9275 (N_9275,N_4995,N_882);
nand U9276 (N_9276,N_983,N_2910);
nor U9277 (N_9277,N_3768,N_390);
or U9278 (N_9278,N_284,N_1941);
or U9279 (N_9279,N_3604,N_1276);
nor U9280 (N_9280,N_1137,N_3642);
nand U9281 (N_9281,N_4062,N_4334);
and U9282 (N_9282,N_1135,N_2060);
xnor U9283 (N_9283,N_660,N_375);
nand U9284 (N_9284,N_3066,N_315);
or U9285 (N_9285,N_2450,N_629);
or U9286 (N_9286,N_1458,N_997);
nor U9287 (N_9287,N_2889,N_4040);
nor U9288 (N_9288,N_2725,N_439);
nand U9289 (N_9289,N_3238,N_2904);
and U9290 (N_9290,N_2414,N_3452);
nor U9291 (N_9291,N_4958,N_1916);
and U9292 (N_9292,N_4746,N_3634);
and U9293 (N_9293,N_3728,N_2362);
nor U9294 (N_9294,N_2272,N_4158);
or U9295 (N_9295,N_638,N_2892);
nand U9296 (N_9296,N_4200,N_506);
nor U9297 (N_9297,N_2872,N_3458);
and U9298 (N_9298,N_1143,N_3096);
and U9299 (N_9299,N_4792,N_4462);
nor U9300 (N_9300,N_4209,N_4643);
nor U9301 (N_9301,N_2938,N_4807);
or U9302 (N_9302,N_3363,N_1676);
and U9303 (N_9303,N_4987,N_1627);
and U9304 (N_9304,N_4678,N_156);
or U9305 (N_9305,N_306,N_1073);
xnor U9306 (N_9306,N_3333,N_3379);
nor U9307 (N_9307,N_1932,N_47);
nor U9308 (N_9308,N_4588,N_719);
nand U9309 (N_9309,N_1009,N_690);
nor U9310 (N_9310,N_26,N_3490);
nor U9311 (N_9311,N_603,N_2222);
nor U9312 (N_9312,N_4087,N_3473);
or U9313 (N_9313,N_2667,N_1274);
or U9314 (N_9314,N_1446,N_2799);
or U9315 (N_9315,N_4351,N_2259);
and U9316 (N_9316,N_67,N_411);
xnor U9317 (N_9317,N_1000,N_4310);
nand U9318 (N_9318,N_4964,N_4667);
xor U9319 (N_9319,N_390,N_2659);
nor U9320 (N_9320,N_3169,N_3565);
or U9321 (N_9321,N_3440,N_3680);
nor U9322 (N_9322,N_4742,N_4865);
nand U9323 (N_9323,N_1454,N_1239);
or U9324 (N_9324,N_4889,N_1530);
and U9325 (N_9325,N_1953,N_1309);
or U9326 (N_9326,N_3897,N_2589);
nand U9327 (N_9327,N_291,N_3574);
or U9328 (N_9328,N_2583,N_1623);
nor U9329 (N_9329,N_1831,N_4998);
xnor U9330 (N_9330,N_357,N_1210);
or U9331 (N_9331,N_3996,N_2828);
and U9332 (N_9332,N_2506,N_4055);
nor U9333 (N_9333,N_1653,N_2587);
nor U9334 (N_9334,N_4449,N_4774);
nand U9335 (N_9335,N_3565,N_2460);
xor U9336 (N_9336,N_3951,N_3822);
or U9337 (N_9337,N_4651,N_900);
xor U9338 (N_9338,N_4099,N_4477);
nor U9339 (N_9339,N_653,N_643);
or U9340 (N_9340,N_2716,N_484);
and U9341 (N_9341,N_341,N_3416);
and U9342 (N_9342,N_4503,N_4247);
or U9343 (N_9343,N_580,N_2023);
or U9344 (N_9344,N_2942,N_1976);
or U9345 (N_9345,N_4886,N_2610);
or U9346 (N_9346,N_172,N_2805);
or U9347 (N_9347,N_4068,N_1185);
nor U9348 (N_9348,N_4788,N_2487);
nor U9349 (N_9349,N_1060,N_808);
or U9350 (N_9350,N_4819,N_2359);
nor U9351 (N_9351,N_4037,N_2240);
and U9352 (N_9352,N_3246,N_4396);
nor U9353 (N_9353,N_2743,N_1303);
or U9354 (N_9354,N_4912,N_2906);
nor U9355 (N_9355,N_1971,N_3426);
nand U9356 (N_9356,N_3197,N_2768);
and U9357 (N_9357,N_639,N_4864);
xnor U9358 (N_9358,N_2491,N_4239);
or U9359 (N_9359,N_573,N_650);
nor U9360 (N_9360,N_694,N_3028);
nor U9361 (N_9361,N_1425,N_604);
and U9362 (N_9362,N_3557,N_378);
nor U9363 (N_9363,N_4706,N_4641);
nor U9364 (N_9364,N_4178,N_1546);
nor U9365 (N_9365,N_3021,N_2316);
xor U9366 (N_9366,N_1087,N_1147);
and U9367 (N_9367,N_4986,N_2615);
and U9368 (N_9368,N_876,N_999);
nand U9369 (N_9369,N_1859,N_4227);
nor U9370 (N_9370,N_3225,N_2361);
nor U9371 (N_9371,N_3179,N_325);
nand U9372 (N_9372,N_428,N_4711);
or U9373 (N_9373,N_1482,N_1478);
nor U9374 (N_9374,N_3646,N_4601);
or U9375 (N_9375,N_2009,N_2125);
or U9376 (N_9376,N_4813,N_2237);
nand U9377 (N_9377,N_4579,N_4207);
or U9378 (N_9378,N_958,N_103);
nand U9379 (N_9379,N_2980,N_2762);
nand U9380 (N_9380,N_2106,N_989);
nor U9381 (N_9381,N_3821,N_2921);
and U9382 (N_9382,N_3456,N_3642);
and U9383 (N_9383,N_1250,N_2079);
nor U9384 (N_9384,N_854,N_4203);
nor U9385 (N_9385,N_605,N_3425);
nor U9386 (N_9386,N_623,N_2647);
nand U9387 (N_9387,N_828,N_2100);
xnor U9388 (N_9388,N_2537,N_4141);
or U9389 (N_9389,N_4229,N_4199);
nand U9390 (N_9390,N_545,N_363);
xnor U9391 (N_9391,N_521,N_593);
xnor U9392 (N_9392,N_4967,N_2959);
or U9393 (N_9393,N_1905,N_47);
or U9394 (N_9394,N_4077,N_4894);
or U9395 (N_9395,N_2857,N_410);
or U9396 (N_9396,N_457,N_4393);
or U9397 (N_9397,N_3118,N_2121);
nor U9398 (N_9398,N_3765,N_3879);
or U9399 (N_9399,N_2611,N_4254);
nor U9400 (N_9400,N_849,N_1146);
or U9401 (N_9401,N_314,N_966);
and U9402 (N_9402,N_2835,N_4885);
nor U9403 (N_9403,N_949,N_4279);
and U9404 (N_9404,N_4141,N_3159);
nand U9405 (N_9405,N_979,N_3615);
and U9406 (N_9406,N_1235,N_3684);
nand U9407 (N_9407,N_2918,N_3759);
or U9408 (N_9408,N_2136,N_2256);
nand U9409 (N_9409,N_2389,N_3150);
nand U9410 (N_9410,N_1542,N_2078);
and U9411 (N_9411,N_715,N_4865);
and U9412 (N_9412,N_1264,N_1767);
xor U9413 (N_9413,N_1231,N_234);
nor U9414 (N_9414,N_1280,N_4539);
and U9415 (N_9415,N_2700,N_2190);
or U9416 (N_9416,N_2407,N_4577);
nor U9417 (N_9417,N_3835,N_2780);
or U9418 (N_9418,N_4315,N_1397);
nor U9419 (N_9419,N_2549,N_342);
nand U9420 (N_9420,N_2884,N_1409);
xnor U9421 (N_9421,N_4953,N_1373);
or U9422 (N_9422,N_894,N_2015);
nand U9423 (N_9423,N_2436,N_1825);
and U9424 (N_9424,N_1116,N_730);
nand U9425 (N_9425,N_2391,N_2588);
or U9426 (N_9426,N_426,N_2519);
or U9427 (N_9427,N_3081,N_1779);
or U9428 (N_9428,N_1346,N_2038);
nand U9429 (N_9429,N_1762,N_1634);
or U9430 (N_9430,N_2842,N_2888);
nor U9431 (N_9431,N_1010,N_4124);
nand U9432 (N_9432,N_2313,N_3171);
or U9433 (N_9433,N_3948,N_2265);
and U9434 (N_9434,N_2501,N_4893);
nand U9435 (N_9435,N_3346,N_1952);
and U9436 (N_9436,N_3119,N_2403);
nor U9437 (N_9437,N_2784,N_49);
nand U9438 (N_9438,N_1731,N_3320);
nand U9439 (N_9439,N_1567,N_4378);
nand U9440 (N_9440,N_4198,N_2522);
nand U9441 (N_9441,N_4110,N_2080);
xnor U9442 (N_9442,N_501,N_4489);
or U9443 (N_9443,N_2611,N_4851);
and U9444 (N_9444,N_154,N_2086);
and U9445 (N_9445,N_1270,N_2092);
or U9446 (N_9446,N_4944,N_2458);
nor U9447 (N_9447,N_4402,N_2910);
nor U9448 (N_9448,N_478,N_3434);
nand U9449 (N_9449,N_2086,N_4191);
nor U9450 (N_9450,N_3095,N_2355);
nand U9451 (N_9451,N_4584,N_3993);
and U9452 (N_9452,N_1357,N_3753);
nor U9453 (N_9453,N_4820,N_1960);
xnor U9454 (N_9454,N_2787,N_4849);
or U9455 (N_9455,N_1970,N_3055);
and U9456 (N_9456,N_917,N_2222);
nor U9457 (N_9457,N_1119,N_4067);
nor U9458 (N_9458,N_2843,N_1939);
and U9459 (N_9459,N_409,N_3386);
nor U9460 (N_9460,N_1535,N_1071);
or U9461 (N_9461,N_4106,N_2692);
nor U9462 (N_9462,N_3492,N_1443);
or U9463 (N_9463,N_2319,N_1047);
xnor U9464 (N_9464,N_1063,N_273);
nor U9465 (N_9465,N_2897,N_4478);
nor U9466 (N_9466,N_631,N_4498);
and U9467 (N_9467,N_2412,N_2682);
and U9468 (N_9468,N_4101,N_434);
nor U9469 (N_9469,N_319,N_3751);
nor U9470 (N_9470,N_1287,N_459);
xor U9471 (N_9471,N_4347,N_4248);
nand U9472 (N_9472,N_422,N_3880);
nor U9473 (N_9473,N_4072,N_1450);
nand U9474 (N_9474,N_1240,N_1162);
nor U9475 (N_9475,N_127,N_3110);
or U9476 (N_9476,N_4076,N_4396);
nor U9477 (N_9477,N_1899,N_530);
and U9478 (N_9478,N_4274,N_4812);
xnor U9479 (N_9479,N_3115,N_694);
nor U9480 (N_9480,N_4647,N_3753);
nor U9481 (N_9481,N_3907,N_3779);
nor U9482 (N_9482,N_893,N_570);
xor U9483 (N_9483,N_4146,N_3530);
or U9484 (N_9484,N_4075,N_4011);
nand U9485 (N_9485,N_2744,N_512);
nand U9486 (N_9486,N_3088,N_91);
nand U9487 (N_9487,N_4528,N_322);
nor U9488 (N_9488,N_411,N_612);
or U9489 (N_9489,N_1590,N_2232);
or U9490 (N_9490,N_3658,N_2665);
nor U9491 (N_9491,N_4390,N_3806);
nor U9492 (N_9492,N_3851,N_1942);
or U9493 (N_9493,N_4331,N_4260);
xnor U9494 (N_9494,N_593,N_1550);
or U9495 (N_9495,N_3937,N_753);
nor U9496 (N_9496,N_3481,N_2170);
nor U9497 (N_9497,N_2807,N_393);
xor U9498 (N_9498,N_4170,N_4235);
and U9499 (N_9499,N_3047,N_1501);
nand U9500 (N_9500,N_229,N_3865);
or U9501 (N_9501,N_3413,N_1957);
and U9502 (N_9502,N_2250,N_4352);
or U9503 (N_9503,N_2512,N_4330);
nor U9504 (N_9504,N_875,N_2469);
and U9505 (N_9505,N_567,N_54);
nor U9506 (N_9506,N_262,N_1970);
or U9507 (N_9507,N_1142,N_4222);
or U9508 (N_9508,N_213,N_4618);
nand U9509 (N_9509,N_2408,N_796);
nor U9510 (N_9510,N_457,N_4796);
nand U9511 (N_9511,N_2877,N_30);
nand U9512 (N_9512,N_479,N_3503);
and U9513 (N_9513,N_4554,N_3424);
and U9514 (N_9514,N_2921,N_3112);
xor U9515 (N_9515,N_544,N_1329);
nor U9516 (N_9516,N_1840,N_664);
nand U9517 (N_9517,N_4684,N_2787);
nor U9518 (N_9518,N_2746,N_3244);
and U9519 (N_9519,N_4681,N_4821);
nor U9520 (N_9520,N_2208,N_180);
nor U9521 (N_9521,N_1838,N_2830);
and U9522 (N_9522,N_4934,N_3780);
or U9523 (N_9523,N_2080,N_3320);
and U9524 (N_9524,N_3844,N_4908);
nand U9525 (N_9525,N_3288,N_1743);
nand U9526 (N_9526,N_2898,N_2464);
nor U9527 (N_9527,N_1940,N_1646);
nor U9528 (N_9528,N_1760,N_3885);
or U9529 (N_9529,N_1162,N_4203);
and U9530 (N_9530,N_257,N_479);
nor U9531 (N_9531,N_545,N_4513);
or U9532 (N_9532,N_475,N_485);
nand U9533 (N_9533,N_1114,N_2451);
or U9534 (N_9534,N_3566,N_590);
nand U9535 (N_9535,N_1644,N_677);
nand U9536 (N_9536,N_1703,N_4606);
nor U9537 (N_9537,N_3271,N_450);
or U9538 (N_9538,N_2573,N_1524);
and U9539 (N_9539,N_4817,N_1743);
and U9540 (N_9540,N_2579,N_2113);
nor U9541 (N_9541,N_3943,N_4846);
nand U9542 (N_9542,N_1728,N_2670);
nor U9543 (N_9543,N_976,N_2806);
xor U9544 (N_9544,N_3198,N_3439);
nor U9545 (N_9545,N_3990,N_270);
nand U9546 (N_9546,N_2760,N_2629);
nor U9547 (N_9547,N_4094,N_1155);
or U9548 (N_9548,N_3991,N_2253);
nand U9549 (N_9549,N_3451,N_1042);
nand U9550 (N_9550,N_1090,N_2886);
and U9551 (N_9551,N_2392,N_1019);
nand U9552 (N_9552,N_2678,N_488);
nor U9553 (N_9553,N_3267,N_85);
nand U9554 (N_9554,N_1234,N_2194);
nand U9555 (N_9555,N_1952,N_357);
nand U9556 (N_9556,N_2772,N_703);
xnor U9557 (N_9557,N_1399,N_186);
or U9558 (N_9558,N_3752,N_3235);
nand U9559 (N_9559,N_3763,N_1843);
or U9560 (N_9560,N_4689,N_1238);
or U9561 (N_9561,N_2246,N_3986);
and U9562 (N_9562,N_610,N_1739);
nor U9563 (N_9563,N_1492,N_378);
nand U9564 (N_9564,N_3233,N_2694);
xnor U9565 (N_9565,N_1846,N_2324);
nor U9566 (N_9566,N_860,N_2080);
nand U9567 (N_9567,N_3773,N_785);
or U9568 (N_9568,N_4897,N_1630);
or U9569 (N_9569,N_2723,N_1475);
and U9570 (N_9570,N_197,N_1398);
and U9571 (N_9571,N_2589,N_3424);
xor U9572 (N_9572,N_986,N_452);
and U9573 (N_9573,N_1655,N_3981);
xnor U9574 (N_9574,N_4495,N_3425);
nand U9575 (N_9575,N_4766,N_982);
xnor U9576 (N_9576,N_385,N_2417);
or U9577 (N_9577,N_1418,N_2136);
nor U9578 (N_9578,N_1095,N_1239);
nor U9579 (N_9579,N_2231,N_622);
nand U9580 (N_9580,N_3412,N_3955);
nand U9581 (N_9581,N_1248,N_2833);
or U9582 (N_9582,N_2742,N_1931);
and U9583 (N_9583,N_2106,N_108);
nor U9584 (N_9584,N_4802,N_45);
nor U9585 (N_9585,N_1208,N_3205);
or U9586 (N_9586,N_21,N_2310);
nor U9587 (N_9587,N_4613,N_4197);
nand U9588 (N_9588,N_2933,N_4127);
nand U9589 (N_9589,N_266,N_1424);
or U9590 (N_9590,N_3744,N_689);
or U9591 (N_9591,N_1165,N_4602);
and U9592 (N_9592,N_2981,N_3866);
nor U9593 (N_9593,N_4888,N_87);
nand U9594 (N_9594,N_2259,N_4532);
and U9595 (N_9595,N_339,N_73);
and U9596 (N_9596,N_3545,N_951);
xnor U9597 (N_9597,N_783,N_1953);
or U9598 (N_9598,N_1783,N_4243);
and U9599 (N_9599,N_1104,N_1027);
nor U9600 (N_9600,N_638,N_1301);
or U9601 (N_9601,N_3806,N_3966);
nand U9602 (N_9602,N_4896,N_3538);
nor U9603 (N_9603,N_2590,N_3765);
xnor U9604 (N_9604,N_1799,N_3829);
and U9605 (N_9605,N_1143,N_4389);
xor U9606 (N_9606,N_3495,N_1049);
nand U9607 (N_9607,N_2322,N_3294);
nand U9608 (N_9608,N_623,N_3760);
or U9609 (N_9609,N_1714,N_3678);
and U9610 (N_9610,N_3906,N_1674);
nor U9611 (N_9611,N_3067,N_3867);
and U9612 (N_9612,N_4349,N_2030);
and U9613 (N_9613,N_3953,N_4139);
nand U9614 (N_9614,N_1272,N_420);
and U9615 (N_9615,N_2516,N_3799);
and U9616 (N_9616,N_260,N_339);
nor U9617 (N_9617,N_4266,N_2562);
nor U9618 (N_9618,N_651,N_1125);
or U9619 (N_9619,N_4005,N_847);
and U9620 (N_9620,N_4012,N_4422);
and U9621 (N_9621,N_1799,N_3005);
nand U9622 (N_9622,N_4359,N_49);
xnor U9623 (N_9623,N_3164,N_3360);
nand U9624 (N_9624,N_80,N_1924);
nor U9625 (N_9625,N_4208,N_1380);
nand U9626 (N_9626,N_628,N_1596);
nor U9627 (N_9627,N_3800,N_1520);
xor U9628 (N_9628,N_4453,N_3894);
nor U9629 (N_9629,N_483,N_653);
nor U9630 (N_9630,N_1557,N_4382);
and U9631 (N_9631,N_2804,N_1504);
xnor U9632 (N_9632,N_4026,N_3993);
nand U9633 (N_9633,N_1108,N_4307);
nor U9634 (N_9634,N_860,N_2254);
or U9635 (N_9635,N_3248,N_2985);
nand U9636 (N_9636,N_4388,N_1978);
nand U9637 (N_9637,N_3186,N_1477);
nand U9638 (N_9638,N_1238,N_507);
nor U9639 (N_9639,N_366,N_1764);
xor U9640 (N_9640,N_1932,N_1300);
and U9641 (N_9641,N_531,N_231);
nand U9642 (N_9642,N_2838,N_2806);
nand U9643 (N_9643,N_389,N_1957);
nand U9644 (N_9644,N_2158,N_26);
nand U9645 (N_9645,N_343,N_4123);
and U9646 (N_9646,N_668,N_304);
or U9647 (N_9647,N_2519,N_3924);
nor U9648 (N_9648,N_24,N_2861);
or U9649 (N_9649,N_1503,N_4995);
nand U9650 (N_9650,N_2446,N_503);
xnor U9651 (N_9651,N_3264,N_4225);
nand U9652 (N_9652,N_3067,N_3835);
and U9653 (N_9653,N_652,N_2354);
or U9654 (N_9654,N_4547,N_334);
nor U9655 (N_9655,N_4383,N_4870);
xor U9656 (N_9656,N_2223,N_940);
or U9657 (N_9657,N_645,N_4539);
or U9658 (N_9658,N_1287,N_4776);
and U9659 (N_9659,N_830,N_1961);
nand U9660 (N_9660,N_672,N_368);
nand U9661 (N_9661,N_199,N_782);
xnor U9662 (N_9662,N_3452,N_2447);
nor U9663 (N_9663,N_1496,N_3043);
xor U9664 (N_9664,N_431,N_1503);
nor U9665 (N_9665,N_544,N_1223);
or U9666 (N_9666,N_6,N_1318);
and U9667 (N_9667,N_2412,N_3487);
nor U9668 (N_9668,N_473,N_1740);
or U9669 (N_9669,N_4974,N_4170);
nor U9670 (N_9670,N_2983,N_1835);
or U9671 (N_9671,N_704,N_2448);
or U9672 (N_9672,N_341,N_1376);
nand U9673 (N_9673,N_4966,N_3336);
nand U9674 (N_9674,N_980,N_661);
or U9675 (N_9675,N_2128,N_607);
or U9676 (N_9676,N_4601,N_4551);
nor U9677 (N_9677,N_2613,N_1667);
or U9678 (N_9678,N_1044,N_3807);
xor U9679 (N_9679,N_175,N_3441);
or U9680 (N_9680,N_3607,N_2412);
or U9681 (N_9681,N_4281,N_2128);
nor U9682 (N_9682,N_3102,N_3357);
xnor U9683 (N_9683,N_329,N_644);
nor U9684 (N_9684,N_2812,N_1047);
nand U9685 (N_9685,N_4547,N_4244);
or U9686 (N_9686,N_2808,N_201);
nand U9687 (N_9687,N_245,N_257);
nor U9688 (N_9688,N_1488,N_2995);
or U9689 (N_9689,N_346,N_230);
nand U9690 (N_9690,N_3444,N_4871);
or U9691 (N_9691,N_4428,N_1977);
and U9692 (N_9692,N_388,N_4908);
nor U9693 (N_9693,N_1558,N_1939);
nor U9694 (N_9694,N_2949,N_1075);
or U9695 (N_9695,N_4395,N_398);
nor U9696 (N_9696,N_1257,N_2062);
and U9697 (N_9697,N_4938,N_4679);
and U9698 (N_9698,N_677,N_1457);
or U9699 (N_9699,N_389,N_2707);
nand U9700 (N_9700,N_3003,N_2957);
nor U9701 (N_9701,N_4000,N_1750);
nor U9702 (N_9702,N_2184,N_1911);
xnor U9703 (N_9703,N_4807,N_198);
xor U9704 (N_9704,N_268,N_1575);
and U9705 (N_9705,N_2294,N_2439);
nor U9706 (N_9706,N_2096,N_521);
or U9707 (N_9707,N_4615,N_4863);
or U9708 (N_9708,N_3312,N_1971);
and U9709 (N_9709,N_4055,N_3627);
nand U9710 (N_9710,N_1959,N_3102);
nor U9711 (N_9711,N_3579,N_3026);
or U9712 (N_9712,N_2363,N_2795);
nand U9713 (N_9713,N_4033,N_3244);
and U9714 (N_9714,N_1976,N_4924);
nand U9715 (N_9715,N_4776,N_2089);
or U9716 (N_9716,N_1507,N_3271);
or U9717 (N_9717,N_4408,N_15);
and U9718 (N_9718,N_248,N_4650);
nor U9719 (N_9719,N_271,N_708);
and U9720 (N_9720,N_780,N_1632);
nand U9721 (N_9721,N_4211,N_2712);
or U9722 (N_9722,N_1753,N_1640);
nand U9723 (N_9723,N_988,N_4123);
nor U9724 (N_9724,N_883,N_506);
and U9725 (N_9725,N_1459,N_2443);
nor U9726 (N_9726,N_1926,N_3561);
and U9727 (N_9727,N_1960,N_579);
nand U9728 (N_9728,N_2625,N_89);
nand U9729 (N_9729,N_1592,N_3140);
or U9730 (N_9730,N_851,N_1596);
and U9731 (N_9731,N_3510,N_4115);
nor U9732 (N_9732,N_2758,N_641);
and U9733 (N_9733,N_2998,N_645);
or U9734 (N_9734,N_4581,N_3419);
nor U9735 (N_9735,N_304,N_2348);
or U9736 (N_9736,N_2316,N_830);
nand U9737 (N_9737,N_2028,N_3732);
and U9738 (N_9738,N_3528,N_3495);
nor U9739 (N_9739,N_3468,N_2723);
or U9740 (N_9740,N_1670,N_1729);
nand U9741 (N_9741,N_509,N_1269);
and U9742 (N_9742,N_3749,N_1309);
xor U9743 (N_9743,N_3892,N_2699);
or U9744 (N_9744,N_3477,N_1166);
or U9745 (N_9745,N_612,N_3394);
or U9746 (N_9746,N_481,N_1058);
and U9747 (N_9747,N_3878,N_4434);
nor U9748 (N_9748,N_195,N_3862);
nand U9749 (N_9749,N_160,N_2080);
or U9750 (N_9750,N_4389,N_2145);
and U9751 (N_9751,N_3462,N_3200);
nor U9752 (N_9752,N_2330,N_4479);
and U9753 (N_9753,N_1129,N_1179);
xor U9754 (N_9754,N_3243,N_359);
xnor U9755 (N_9755,N_3552,N_423);
or U9756 (N_9756,N_4513,N_2034);
nand U9757 (N_9757,N_637,N_4377);
or U9758 (N_9758,N_2372,N_2038);
nand U9759 (N_9759,N_2163,N_4086);
nor U9760 (N_9760,N_2444,N_4004);
nand U9761 (N_9761,N_3470,N_4409);
nor U9762 (N_9762,N_456,N_4634);
or U9763 (N_9763,N_3120,N_1267);
nor U9764 (N_9764,N_3212,N_4648);
or U9765 (N_9765,N_1620,N_2725);
or U9766 (N_9766,N_1969,N_2569);
nand U9767 (N_9767,N_3967,N_2191);
nand U9768 (N_9768,N_522,N_2803);
and U9769 (N_9769,N_4759,N_4224);
nor U9770 (N_9770,N_1187,N_2418);
nor U9771 (N_9771,N_1704,N_2398);
nor U9772 (N_9772,N_3281,N_1913);
or U9773 (N_9773,N_1219,N_3450);
nor U9774 (N_9774,N_2998,N_478);
or U9775 (N_9775,N_1427,N_4442);
nor U9776 (N_9776,N_1865,N_1710);
nand U9777 (N_9777,N_3900,N_1437);
and U9778 (N_9778,N_2165,N_2657);
and U9779 (N_9779,N_739,N_516);
nor U9780 (N_9780,N_3785,N_1600);
or U9781 (N_9781,N_855,N_668);
and U9782 (N_9782,N_4732,N_2069);
or U9783 (N_9783,N_2174,N_1055);
nand U9784 (N_9784,N_4209,N_4638);
nor U9785 (N_9785,N_1907,N_1947);
xnor U9786 (N_9786,N_4571,N_603);
or U9787 (N_9787,N_859,N_792);
nor U9788 (N_9788,N_3225,N_1774);
nand U9789 (N_9789,N_1869,N_755);
and U9790 (N_9790,N_3233,N_65);
xnor U9791 (N_9791,N_1797,N_2876);
nand U9792 (N_9792,N_3599,N_308);
or U9793 (N_9793,N_4782,N_1470);
nor U9794 (N_9794,N_3018,N_376);
or U9795 (N_9795,N_2478,N_1333);
or U9796 (N_9796,N_4048,N_2555);
or U9797 (N_9797,N_882,N_4994);
nor U9798 (N_9798,N_2720,N_1696);
or U9799 (N_9799,N_3915,N_1802);
nand U9800 (N_9800,N_85,N_983);
and U9801 (N_9801,N_3198,N_161);
nand U9802 (N_9802,N_2180,N_630);
and U9803 (N_9803,N_647,N_409);
xor U9804 (N_9804,N_3466,N_3132);
xor U9805 (N_9805,N_3008,N_298);
or U9806 (N_9806,N_4571,N_2824);
nor U9807 (N_9807,N_3984,N_4527);
or U9808 (N_9808,N_299,N_425);
nand U9809 (N_9809,N_4185,N_3737);
nand U9810 (N_9810,N_2782,N_659);
nor U9811 (N_9811,N_4815,N_604);
and U9812 (N_9812,N_2046,N_2823);
nand U9813 (N_9813,N_3811,N_2603);
and U9814 (N_9814,N_2532,N_979);
xnor U9815 (N_9815,N_3702,N_1248);
xnor U9816 (N_9816,N_1379,N_2191);
nand U9817 (N_9817,N_2955,N_4642);
nor U9818 (N_9818,N_1940,N_3487);
nand U9819 (N_9819,N_3012,N_1784);
nor U9820 (N_9820,N_3991,N_2869);
xor U9821 (N_9821,N_2382,N_248);
nor U9822 (N_9822,N_1592,N_4147);
or U9823 (N_9823,N_2665,N_1765);
nor U9824 (N_9824,N_1155,N_4273);
nor U9825 (N_9825,N_4456,N_2947);
and U9826 (N_9826,N_2252,N_342);
nand U9827 (N_9827,N_1407,N_4983);
or U9828 (N_9828,N_2420,N_2979);
and U9829 (N_9829,N_3474,N_3596);
nand U9830 (N_9830,N_3152,N_2980);
or U9831 (N_9831,N_1942,N_2783);
and U9832 (N_9832,N_3667,N_3640);
and U9833 (N_9833,N_3765,N_3050);
or U9834 (N_9834,N_610,N_3517);
or U9835 (N_9835,N_4267,N_2269);
and U9836 (N_9836,N_93,N_934);
nand U9837 (N_9837,N_1588,N_3198);
nor U9838 (N_9838,N_2840,N_168);
nand U9839 (N_9839,N_1153,N_49);
or U9840 (N_9840,N_1038,N_1923);
and U9841 (N_9841,N_3258,N_1942);
and U9842 (N_9842,N_727,N_3780);
nor U9843 (N_9843,N_1414,N_4382);
or U9844 (N_9844,N_3783,N_1466);
xor U9845 (N_9845,N_2208,N_975);
or U9846 (N_9846,N_1809,N_2929);
nor U9847 (N_9847,N_1976,N_3812);
and U9848 (N_9848,N_2690,N_4530);
or U9849 (N_9849,N_4714,N_4321);
or U9850 (N_9850,N_1894,N_4063);
and U9851 (N_9851,N_1922,N_3274);
or U9852 (N_9852,N_4926,N_4159);
nand U9853 (N_9853,N_4610,N_1752);
nand U9854 (N_9854,N_2369,N_4668);
or U9855 (N_9855,N_910,N_1715);
nor U9856 (N_9856,N_4751,N_279);
nor U9857 (N_9857,N_4638,N_2139);
or U9858 (N_9858,N_2283,N_853);
nor U9859 (N_9859,N_3128,N_38);
and U9860 (N_9860,N_3064,N_4681);
or U9861 (N_9861,N_2151,N_4882);
nand U9862 (N_9862,N_3962,N_1674);
nand U9863 (N_9863,N_1188,N_1623);
and U9864 (N_9864,N_2825,N_1414);
or U9865 (N_9865,N_4120,N_4658);
nor U9866 (N_9866,N_466,N_3019);
nand U9867 (N_9867,N_1419,N_528);
and U9868 (N_9868,N_3500,N_3774);
or U9869 (N_9869,N_1356,N_1443);
nand U9870 (N_9870,N_2003,N_4891);
and U9871 (N_9871,N_3283,N_3926);
or U9872 (N_9872,N_4708,N_1638);
and U9873 (N_9873,N_2053,N_356);
nand U9874 (N_9874,N_1608,N_2404);
nand U9875 (N_9875,N_4599,N_423);
or U9876 (N_9876,N_1564,N_1160);
nor U9877 (N_9877,N_4763,N_4896);
or U9878 (N_9878,N_4367,N_4351);
and U9879 (N_9879,N_3408,N_2200);
nand U9880 (N_9880,N_1698,N_1413);
nor U9881 (N_9881,N_3866,N_3178);
and U9882 (N_9882,N_4616,N_2451);
and U9883 (N_9883,N_465,N_3029);
nor U9884 (N_9884,N_812,N_236);
nor U9885 (N_9885,N_1017,N_2989);
nand U9886 (N_9886,N_4232,N_2959);
and U9887 (N_9887,N_2227,N_1579);
xnor U9888 (N_9888,N_969,N_2595);
nand U9889 (N_9889,N_318,N_1404);
and U9890 (N_9890,N_677,N_4529);
or U9891 (N_9891,N_1321,N_4521);
xnor U9892 (N_9892,N_4702,N_1810);
and U9893 (N_9893,N_3549,N_3747);
nand U9894 (N_9894,N_2203,N_975);
or U9895 (N_9895,N_4678,N_2754);
or U9896 (N_9896,N_4843,N_288);
and U9897 (N_9897,N_2523,N_4424);
nand U9898 (N_9898,N_988,N_3662);
and U9899 (N_9899,N_2208,N_4018);
or U9900 (N_9900,N_2690,N_4698);
nor U9901 (N_9901,N_3282,N_1817);
or U9902 (N_9902,N_3156,N_4843);
nand U9903 (N_9903,N_4350,N_4068);
nand U9904 (N_9904,N_3878,N_844);
nor U9905 (N_9905,N_2256,N_2139);
or U9906 (N_9906,N_1465,N_773);
or U9907 (N_9907,N_203,N_2922);
and U9908 (N_9908,N_1278,N_4407);
or U9909 (N_9909,N_4781,N_4510);
nand U9910 (N_9910,N_1935,N_2556);
and U9911 (N_9911,N_3035,N_2325);
and U9912 (N_9912,N_966,N_2397);
or U9913 (N_9913,N_538,N_320);
xnor U9914 (N_9914,N_1653,N_3415);
or U9915 (N_9915,N_4360,N_1596);
and U9916 (N_9916,N_1857,N_3112);
nor U9917 (N_9917,N_3969,N_2611);
nand U9918 (N_9918,N_1731,N_3058);
or U9919 (N_9919,N_3283,N_561);
and U9920 (N_9920,N_4044,N_4005);
nor U9921 (N_9921,N_4047,N_3803);
or U9922 (N_9922,N_413,N_3569);
nand U9923 (N_9923,N_3319,N_3459);
and U9924 (N_9924,N_3771,N_25);
nor U9925 (N_9925,N_1336,N_4799);
nor U9926 (N_9926,N_1937,N_1289);
xnor U9927 (N_9927,N_2237,N_4776);
and U9928 (N_9928,N_3656,N_4678);
and U9929 (N_9929,N_678,N_1511);
and U9930 (N_9930,N_1089,N_4117);
and U9931 (N_9931,N_3800,N_4615);
and U9932 (N_9932,N_1487,N_1634);
nand U9933 (N_9933,N_3303,N_4899);
or U9934 (N_9934,N_3934,N_134);
and U9935 (N_9935,N_4155,N_4013);
nand U9936 (N_9936,N_4143,N_1471);
or U9937 (N_9937,N_4003,N_3232);
and U9938 (N_9938,N_4337,N_4391);
and U9939 (N_9939,N_2209,N_4305);
and U9940 (N_9940,N_1439,N_4139);
or U9941 (N_9941,N_3216,N_2619);
or U9942 (N_9942,N_1756,N_4675);
nand U9943 (N_9943,N_865,N_3322);
or U9944 (N_9944,N_117,N_3305);
xnor U9945 (N_9945,N_1770,N_3774);
nor U9946 (N_9946,N_2472,N_3788);
or U9947 (N_9947,N_4766,N_2799);
xor U9948 (N_9948,N_3966,N_3519);
nand U9949 (N_9949,N_2945,N_1128);
nand U9950 (N_9950,N_2011,N_1543);
or U9951 (N_9951,N_4794,N_4163);
xor U9952 (N_9952,N_3871,N_3412);
nor U9953 (N_9953,N_3093,N_3894);
nand U9954 (N_9954,N_1022,N_128);
nand U9955 (N_9955,N_4216,N_510);
nor U9956 (N_9956,N_2878,N_1539);
and U9957 (N_9957,N_576,N_291);
and U9958 (N_9958,N_4630,N_4140);
nor U9959 (N_9959,N_3298,N_414);
nor U9960 (N_9960,N_2124,N_4871);
nand U9961 (N_9961,N_2343,N_3557);
or U9962 (N_9962,N_3578,N_159);
nand U9963 (N_9963,N_4465,N_3166);
nand U9964 (N_9964,N_386,N_2851);
nand U9965 (N_9965,N_3430,N_3470);
and U9966 (N_9966,N_2555,N_2676);
nor U9967 (N_9967,N_2025,N_57);
and U9968 (N_9968,N_3782,N_918);
and U9969 (N_9969,N_49,N_2830);
or U9970 (N_9970,N_1409,N_1180);
nor U9971 (N_9971,N_800,N_525);
or U9972 (N_9972,N_3247,N_2097);
and U9973 (N_9973,N_37,N_4748);
nor U9974 (N_9974,N_2900,N_2722);
and U9975 (N_9975,N_2756,N_212);
nor U9976 (N_9976,N_1603,N_3012);
and U9977 (N_9977,N_2227,N_3804);
nor U9978 (N_9978,N_632,N_1931);
nor U9979 (N_9979,N_1303,N_3562);
or U9980 (N_9980,N_3426,N_3632);
or U9981 (N_9981,N_8,N_4947);
xnor U9982 (N_9982,N_2090,N_4446);
nand U9983 (N_9983,N_2504,N_328);
and U9984 (N_9984,N_3602,N_169);
nor U9985 (N_9985,N_3070,N_4583);
or U9986 (N_9986,N_646,N_320);
and U9987 (N_9987,N_4144,N_1043);
nand U9988 (N_9988,N_1202,N_4540);
nand U9989 (N_9989,N_10,N_521);
nor U9990 (N_9990,N_4548,N_1048);
xor U9991 (N_9991,N_3919,N_1171);
or U9992 (N_9992,N_1885,N_599);
and U9993 (N_9993,N_1903,N_1681);
nand U9994 (N_9994,N_4262,N_535);
or U9995 (N_9995,N_3758,N_4270);
and U9996 (N_9996,N_22,N_820);
nand U9997 (N_9997,N_1875,N_3847);
or U9998 (N_9998,N_3688,N_2623);
nand U9999 (N_9999,N_1725,N_1108);
or UO_0 (O_0,N_5013,N_9546);
or UO_1 (O_1,N_8289,N_7070);
nor UO_2 (O_2,N_8370,N_7613);
or UO_3 (O_3,N_8387,N_7114);
nand UO_4 (O_4,N_5698,N_7253);
nor UO_5 (O_5,N_8534,N_7961);
and UO_6 (O_6,N_6354,N_6092);
nand UO_7 (O_7,N_9825,N_5281);
nand UO_8 (O_8,N_5196,N_8514);
or UO_9 (O_9,N_6721,N_8186);
and UO_10 (O_10,N_9902,N_7716);
nand UO_11 (O_11,N_7315,N_5528);
xnor UO_12 (O_12,N_5119,N_7875);
or UO_13 (O_13,N_8709,N_8160);
nor UO_14 (O_14,N_6466,N_9551);
or UO_15 (O_15,N_7828,N_8141);
nand UO_16 (O_16,N_7068,N_8298);
and UO_17 (O_17,N_9203,N_8461);
nand UO_18 (O_18,N_7703,N_6235);
or UO_19 (O_19,N_6425,N_8663);
nand UO_20 (O_20,N_6545,N_7037);
or UO_21 (O_21,N_6278,N_6516);
nor UO_22 (O_22,N_6826,N_8815);
or UO_23 (O_23,N_7733,N_5045);
and UO_24 (O_24,N_7481,N_9453);
and UO_25 (O_25,N_8979,N_6269);
and UO_26 (O_26,N_5527,N_8446);
or UO_27 (O_27,N_5733,N_8331);
and UO_28 (O_28,N_6757,N_9225);
nor UO_29 (O_29,N_8517,N_5006);
nor UO_30 (O_30,N_5850,N_6376);
nand UO_31 (O_31,N_5942,N_5994);
nand UO_32 (O_32,N_5678,N_5416);
and UO_33 (O_33,N_5621,N_7029);
nor UO_34 (O_34,N_5054,N_6271);
or UO_35 (O_35,N_9596,N_9013);
or UO_36 (O_36,N_6836,N_8126);
nand UO_37 (O_37,N_8895,N_6020);
nor UO_38 (O_38,N_7311,N_5271);
or UO_39 (O_39,N_6620,N_9310);
nor UO_40 (O_40,N_7897,N_8661);
nand UO_41 (O_41,N_9305,N_6406);
nand UO_42 (O_42,N_6776,N_8422);
or UO_43 (O_43,N_5614,N_7260);
nand UO_44 (O_44,N_5635,N_6230);
nor UO_45 (O_45,N_9866,N_8632);
or UO_46 (O_46,N_9835,N_6614);
and UO_47 (O_47,N_5682,N_8834);
and UO_48 (O_48,N_7922,N_8396);
nor UO_49 (O_49,N_8500,N_8305);
nor UO_50 (O_50,N_6774,N_5376);
xnor UO_51 (O_51,N_9830,N_5947);
and UO_52 (O_52,N_9528,N_9821);
or UO_53 (O_53,N_9151,N_6844);
and UO_54 (O_54,N_9800,N_9387);
or UO_55 (O_55,N_8220,N_9253);
nand UO_56 (O_56,N_5267,N_5774);
and UO_57 (O_57,N_5563,N_8248);
nand UO_58 (O_58,N_7985,N_6482);
and UO_59 (O_59,N_6348,N_5868);
or UO_60 (O_60,N_7034,N_8616);
nand UO_61 (O_61,N_8109,N_8269);
nand UO_62 (O_62,N_6310,N_9642);
or UO_63 (O_63,N_5131,N_5508);
nor UO_64 (O_64,N_7378,N_9009);
or UO_65 (O_65,N_7097,N_9176);
nor UO_66 (O_66,N_9805,N_5005);
xor UO_67 (O_67,N_5448,N_5787);
nor UO_68 (O_68,N_9402,N_7633);
or UO_69 (O_69,N_9038,N_6123);
nand UO_70 (O_70,N_7067,N_9125);
nand UO_71 (O_71,N_7040,N_5676);
or UO_72 (O_72,N_5568,N_7126);
nand UO_73 (O_73,N_8841,N_9918);
or UO_74 (O_74,N_6041,N_9892);
xor UO_75 (O_75,N_5529,N_8839);
xor UO_76 (O_76,N_9264,N_7510);
or UO_77 (O_77,N_7280,N_8243);
or UO_78 (O_78,N_9313,N_9332);
or UO_79 (O_79,N_7491,N_9245);
and UO_80 (O_80,N_9717,N_9719);
nand UO_81 (O_81,N_6962,N_7272);
nand UO_82 (O_82,N_7972,N_8166);
nand UO_83 (O_83,N_8956,N_6222);
and UO_84 (O_84,N_6115,N_9165);
and UO_85 (O_85,N_9148,N_6445);
nand UO_86 (O_86,N_7222,N_7150);
nor UO_87 (O_87,N_8902,N_8785);
nor UO_88 (O_88,N_6402,N_7538);
or UO_89 (O_89,N_9083,N_5195);
and UO_90 (O_90,N_7359,N_8254);
nand UO_91 (O_91,N_5512,N_7012);
and UO_92 (O_92,N_9811,N_8252);
nor UO_93 (O_93,N_7653,N_7172);
nand UO_94 (O_94,N_6733,N_5216);
or UO_95 (O_95,N_6394,N_5366);
and UO_96 (O_96,N_9451,N_8949);
nand UO_97 (O_97,N_8747,N_5422);
xor UO_98 (O_98,N_6810,N_9256);
or UO_99 (O_99,N_6190,N_6508);
xnor UO_100 (O_100,N_9887,N_7738);
nand UO_101 (O_101,N_8637,N_6752);
and UO_102 (O_102,N_9163,N_7783);
or UO_103 (O_103,N_6048,N_6573);
and UO_104 (O_104,N_8607,N_6586);
nand UO_105 (O_105,N_8447,N_6108);
and UO_106 (O_106,N_9628,N_6770);
nand UO_107 (O_107,N_9792,N_9485);
and UO_108 (O_108,N_8284,N_9577);
nor UO_109 (O_109,N_5155,N_5017);
and UO_110 (O_110,N_9932,N_5011);
or UO_111 (O_111,N_7024,N_9737);
and UO_112 (O_112,N_7986,N_6887);
or UO_113 (O_113,N_7519,N_5824);
xnor UO_114 (O_114,N_6154,N_9959);
nand UO_115 (O_115,N_7808,N_8643);
nand UO_116 (O_116,N_7680,N_8065);
nor UO_117 (O_117,N_5975,N_5709);
nand UO_118 (O_118,N_9957,N_5526);
or UO_119 (O_119,N_8750,N_5143);
nand UO_120 (O_120,N_8678,N_5773);
and UO_121 (O_121,N_7841,N_8568);
xnor UO_122 (O_122,N_9634,N_7873);
nor UO_123 (O_123,N_7837,N_5796);
xnor UO_124 (O_124,N_9073,N_9353);
and UO_125 (O_125,N_9519,N_7347);
nor UO_126 (O_126,N_8941,N_7054);
nor UO_127 (O_127,N_8569,N_5900);
xor UO_128 (O_128,N_8348,N_6529);
or UO_129 (O_129,N_5415,N_5133);
or UO_130 (O_130,N_8480,N_9820);
and UO_131 (O_131,N_9321,N_8170);
or UO_132 (O_132,N_6572,N_9948);
xor UO_133 (O_133,N_6399,N_8960);
nor UO_134 (O_134,N_7902,N_6241);
or UO_135 (O_135,N_5488,N_5918);
nand UO_136 (O_136,N_5021,N_6579);
nor UO_137 (O_137,N_7404,N_8017);
or UO_138 (O_138,N_8946,N_8394);
nand UO_139 (O_139,N_9075,N_7982);
or UO_140 (O_140,N_9605,N_6935);
nor UO_141 (O_141,N_5081,N_8216);
and UO_142 (O_142,N_8911,N_8420);
nor UO_143 (O_143,N_8307,N_6499);
nand UO_144 (O_144,N_6063,N_8688);
nor UO_145 (O_145,N_7848,N_9895);
nand UO_146 (O_146,N_5615,N_8177);
or UO_147 (O_147,N_5727,N_9541);
xnor UO_148 (O_148,N_5842,N_9096);
and UO_149 (O_149,N_6143,N_7386);
and UO_150 (O_150,N_7598,N_5327);
or UO_151 (O_151,N_8824,N_9891);
or UO_152 (O_152,N_6022,N_8219);
or UO_153 (O_153,N_5714,N_6148);
and UO_154 (O_154,N_6793,N_6449);
nor UO_155 (O_155,N_6907,N_7515);
or UO_156 (O_156,N_6863,N_7130);
nand UO_157 (O_157,N_8585,N_6486);
or UO_158 (O_158,N_8975,N_7977);
and UO_159 (O_159,N_6293,N_5108);
nand UO_160 (O_160,N_5840,N_9319);
nand UO_161 (O_161,N_5163,N_5295);
and UO_162 (O_162,N_9104,N_6309);
nand UO_163 (O_163,N_7597,N_6555);
nand UO_164 (O_164,N_5539,N_5022);
and UO_165 (O_165,N_7241,N_7697);
or UO_166 (O_166,N_8261,N_6038);
and UO_167 (O_167,N_7630,N_5479);
xnor UO_168 (O_168,N_5540,N_7340);
nor UO_169 (O_169,N_9436,N_6012);
and UO_170 (O_170,N_8826,N_5386);
or UO_171 (O_171,N_9662,N_6035);
nor UO_172 (O_172,N_9708,N_7686);
nor UO_173 (O_173,N_9135,N_7433);
nor UO_174 (O_174,N_6943,N_5016);
and UO_175 (O_175,N_5089,N_9316);
or UO_176 (O_176,N_9512,N_5972);
and UO_177 (O_177,N_7930,N_6578);
nand UO_178 (O_178,N_8801,N_9268);
nand UO_179 (O_179,N_7147,N_7537);
and UO_180 (O_180,N_5681,N_5565);
or UO_181 (O_181,N_6231,N_6939);
nor UO_182 (O_182,N_9962,N_7533);
or UO_183 (O_183,N_7942,N_7732);
nand UO_184 (O_184,N_7674,N_8711);
nor UO_185 (O_185,N_5241,N_7066);
or UO_186 (O_186,N_5489,N_8345);
nor UO_187 (O_187,N_5307,N_5482);
or UO_188 (O_188,N_5930,N_6695);
or UO_189 (O_189,N_7285,N_9914);
nand UO_190 (O_190,N_9289,N_6053);
nor UO_191 (O_191,N_6911,N_8463);
and UO_192 (O_192,N_5335,N_6172);
and UO_193 (O_193,N_7736,N_6921);
and UO_194 (O_194,N_8303,N_7335);
nand UO_195 (O_195,N_7127,N_9014);
nor UO_196 (O_196,N_5057,N_6392);
or UO_197 (O_197,N_7775,N_9753);
xnor UO_198 (O_198,N_8809,N_6133);
and UO_199 (O_199,N_9702,N_5076);
nand UO_200 (O_200,N_8677,N_5828);
and UO_201 (O_201,N_9364,N_8584);
xnor UO_202 (O_202,N_8428,N_8885);
or UO_203 (O_203,N_7685,N_5889);
and UO_204 (O_204,N_8513,N_9182);
or UO_205 (O_205,N_9735,N_7091);
nand UO_206 (O_206,N_8840,N_5538);
and UO_207 (O_207,N_9864,N_9495);
and UO_208 (O_208,N_5302,N_8057);
and UO_209 (O_209,N_7795,N_8433);
nand UO_210 (O_210,N_9214,N_5244);
nand UO_211 (O_211,N_9237,N_6030);
xnor UO_212 (O_212,N_7678,N_5860);
and UO_213 (O_213,N_8007,N_5050);
and UO_214 (O_214,N_9466,N_7008);
or UO_215 (O_215,N_5124,N_8787);
and UO_216 (O_216,N_6896,N_7745);
nand UO_217 (O_217,N_6446,N_7714);
xnor UO_218 (O_218,N_5931,N_5537);
xor UO_219 (O_219,N_9184,N_6481);
nor UO_220 (O_220,N_9993,N_6125);
nor UO_221 (O_221,N_6386,N_6709);
and UO_222 (O_222,N_9697,N_8628);
nand UO_223 (O_223,N_5484,N_9026);
or UO_224 (O_224,N_8759,N_6430);
nor UO_225 (O_225,N_9623,N_8635);
nor UO_226 (O_226,N_8951,N_7208);
or UO_227 (O_227,N_9973,N_5659);
and UO_228 (O_228,N_8820,N_9745);
nor UO_229 (O_229,N_8575,N_8606);
xor UO_230 (O_230,N_6355,N_8594);
xor UO_231 (O_231,N_8444,N_5243);
nand UO_232 (O_232,N_9802,N_9930);
xnor UO_233 (O_233,N_6951,N_8054);
nor UO_234 (O_234,N_9718,N_6680);
xnor UO_235 (O_235,N_5815,N_7954);
nand UO_236 (O_236,N_9205,N_5401);
nand UO_237 (O_237,N_9826,N_7125);
xor UO_238 (O_238,N_5801,N_8184);
or UO_239 (O_239,N_7266,N_7996);
xnor UO_240 (O_240,N_5719,N_9257);
nand UO_241 (O_241,N_6812,N_9230);
and UO_242 (O_242,N_9040,N_6996);
or UO_243 (O_243,N_9335,N_5495);
nor UO_244 (O_244,N_5798,N_8919);
nor UO_245 (O_245,N_8933,N_9143);
and UO_246 (O_246,N_7947,N_6847);
and UO_247 (O_247,N_5861,N_6729);
nand UO_248 (O_248,N_7143,N_7536);
nand UO_249 (O_249,N_7225,N_6510);
nand UO_250 (O_250,N_7402,N_6672);
nor UO_251 (O_251,N_6541,N_6470);
nor UO_252 (O_252,N_8765,N_6275);
or UO_253 (O_253,N_8980,N_5166);
nor UO_254 (O_254,N_8909,N_5349);
nand UO_255 (O_255,N_7850,N_7909);
nor UO_256 (O_256,N_6912,N_9124);
or UO_257 (O_257,N_5957,N_8664);
nor UO_258 (O_258,N_5873,N_7577);
and UO_259 (O_259,N_9549,N_8786);
and UO_260 (O_260,N_9691,N_5321);
nor UO_261 (O_261,N_7554,N_8851);
nand UO_262 (O_262,N_6626,N_8278);
nor UO_263 (O_263,N_6450,N_5939);
or UO_264 (O_264,N_8324,N_7473);
nor UO_265 (O_265,N_6040,N_8070);
nand UO_266 (O_266,N_6152,N_9033);
or UO_267 (O_267,N_6690,N_9782);
nand UO_268 (O_268,N_7463,N_5616);
or UO_269 (O_269,N_8409,N_5036);
and UO_270 (O_270,N_6627,N_7606);
and UO_271 (O_271,N_5266,N_5212);
nand UO_272 (O_272,N_6571,N_9952);
xnor UO_273 (O_273,N_7937,N_5726);
or UO_274 (O_274,N_5988,N_5684);
and UO_275 (O_275,N_6232,N_6807);
nor UO_276 (O_276,N_5769,N_5954);
and UO_277 (O_277,N_8772,N_7590);
and UO_278 (O_278,N_5091,N_6057);
xnor UO_279 (O_279,N_7403,N_8091);
xor UO_280 (O_280,N_7166,N_9990);
nand UO_281 (O_281,N_5569,N_8648);
and UO_282 (O_282,N_9599,N_8322);
xor UO_283 (O_283,N_7492,N_6089);
and UO_284 (O_284,N_7165,N_6443);
xor UO_285 (O_285,N_6609,N_6352);
nand UO_286 (O_286,N_5835,N_8614);
and UO_287 (O_287,N_8958,N_5193);
nor UO_288 (O_288,N_6795,N_7220);
nand UO_289 (O_289,N_5012,N_8586);
nor UO_290 (O_290,N_7093,N_9638);
nand UO_291 (O_291,N_9566,N_6305);
nand UO_292 (O_292,N_9833,N_5309);
nand UO_293 (O_293,N_6639,N_5269);
nand UO_294 (O_294,N_9232,N_5984);
nor UO_295 (O_295,N_9141,N_5973);
and UO_296 (O_296,N_8764,N_9224);
or UO_297 (O_297,N_5661,N_7702);
nand UO_298 (O_298,N_8489,N_6936);
and UO_299 (O_299,N_9363,N_7596);
nor UO_300 (O_300,N_8268,N_9018);
nor UO_301 (O_301,N_8150,N_5812);
nor UO_302 (O_302,N_8942,N_9196);
and UO_303 (O_303,N_7277,N_9654);
and UO_304 (O_304,N_9243,N_6250);
nor UO_305 (O_305,N_5795,N_5142);
or UO_306 (O_306,N_7073,N_9049);
and UO_307 (O_307,N_8692,N_9815);
and UO_308 (O_308,N_7973,N_8889);
or UO_309 (O_309,N_5120,N_6464);
nor UO_310 (O_310,N_8768,N_7207);
nand UO_311 (O_311,N_8213,N_5061);
nor UO_312 (O_312,N_9710,N_8224);
or UO_313 (O_313,N_8351,N_5202);
and UO_314 (O_314,N_6905,N_8888);
and UO_315 (O_315,N_6457,N_5003);
and UO_316 (O_316,N_5403,N_5179);
nor UO_317 (O_317,N_9780,N_8506);
or UO_318 (O_318,N_5296,N_8292);
nor UO_319 (O_319,N_5458,N_8967);
xnor UO_320 (O_320,N_7584,N_5953);
or UO_321 (O_321,N_7323,N_6461);
nor UO_322 (O_322,N_6483,N_5707);
and UO_323 (O_323,N_9444,N_6773);
xor UO_324 (O_324,N_9777,N_8246);
nand UO_325 (O_325,N_8122,N_9425);
nand UO_326 (O_326,N_9762,N_5999);
or UO_327 (O_327,N_6332,N_6409);
and UO_328 (O_328,N_8326,N_6408);
nor UO_329 (O_329,N_5360,N_7699);
or UO_330 (O_330,N_6494,N_9056);
nor UO_331 (O_331,N_5749,N_5979);
xor UO_332 (O_332,N_5697,N_8432);
and UO_333 (O_333,N_9352,N_6149);
or UO_334 (O_334,N_9482,N_7546);
nor UO_335 (O_335,N_5759,N_9211);
or UO_336 (O_336,N_9396,N_7022);
or UO_337 (O_337,N_7957,N_6944);
or UO_338 (O_338,N_6712,N_9302);
xnor UO_339 (O_339,N_8483,N_7761);
or UO_340 (O_340,N_8465,N_9161);
and UO_341 (O_341,N_6834,N_7965);
nor UO_342 (O_342,N_9273,N_7968);
and UO_343 (O_343,N_9481,N_5917);
xor UO_344 (O_344,N_6313,N_6279);
and UO_345 (O_345,N_6363,N_6244);
or UO_346 (O_346,N_8358,N_6135);
nand UO_347 (O_347,N_5444,N_7128);
nor UO_348 (O_348,N_8223,N_9137);
and UO_349 (O_349,N_8095,N_6946);
nor UO_350 (O_350,N_9729,N_7031);
nor UO_351 (O_351,N_5059,N_5075);
or UO_352 (O_352,N_8469,N_6373);
or UO_353 (O_353,N_7483,N_7926);
nand UO_354 (O_354,N_6223,N_7906);
and UO_355 (O_355,N_5080,N_6985);
or UO_356 (O_356,N_8864,N_8683);
xnor UO_357 (O_357,N_8317,N_9950);
or UO_358 (O_358,N_9395,N_6766);
and UO_359 (O_359,N_7729,N_6168);
xnor UO_360 (O_360,N_6248,N_9544);
xnor UO_361 (O_361,N_5078,N_6359);
nor UO_362 (O_362,N_6633,N_9852);
or UO_363 (O_363,N_6934,N_7429);
or UO_364 (O_364,N_6480,N_7593);
and UO_365 (O_365,N_9924,N_6253);
nand UO_366 (O_366,N_8380,N_6725);
and UO_367 (O_367,N_7441,N_8442);
or UO_368 (O_368,N_7489,N_8069);
or UO_369 (O_369,N_5753,N_7294);
and UO_370 (O_370,N_8312,N_8361);
and UO_371 (O_371,N_9410,N_5729);
nand UO_372 (O_372,N_6666,N_9876);
or UO_373 (O_373,N_5786,N_7490);
or UO_374 (O_374,N_8222,N_8060);
xor UO_375 (O_375,N_6920,N_6740);
nor UO_376 (O_376,N_6800,N_7883);
nor UO_377 (O_377,N_6853,N_7187);
and UO_378 (O_378,N_8127,N_7364);
and UO_379 (O_379,N_5126,N_9457);
or UO_380 (O_380,N_6517,N_8587);
nand UO_381 (O_381,N_8753,N_9011);
or UO_382 (O_382,N_9626,N_9497);
nand UO_383 (O_383,N_5268,N_9149);
or UO_384 (O_384,N_7047,N_7956);
nand UO_385 (O_385,N_9508,N_6025);
nor UO_386 (O_386,N_9756,N_9912);
xnor UO_387 (O_387,N_6438,N_9198);
nor UO_388 (O_388,N_7249,N_6631);
nor UO_389 (O_389,N_9744,N_8399);
and UO_390 (O_390,N_5418,N_8424);
nor UO_391 (O_391,N_9447,N_7813);
or UO_392 (O_392,N_9167,N_7343);
nand UO_393 (O_393,N_7310,N_9020);
nor UO_394 (O_394,N_9153,N_6021);
nor UO_395 (O_395,N_7728,N_5328);
and UO_396 (O_396,N_8953,N_9849);
xor UO_397 (O_397,N_8563,N_8842);
and UO_398 (O_398,N_6525,N_9515);
xor UO_399 (O_399,N_5001,N_7531);
and UO_400 (O_400,N_9538,N_6391);
or UO_401 (O_401,N_5863,N_7677);
or UO_402 (O_402,N_5689,N_7035);
and UO_403 (O_403,N_8571,N_9565);
nor UO_404 (O_404,N_5663,N_9720);
or UO_405 (O_405,N_9222,N_9129);
and UO_406 (O_406,N_9078,N_8674);
nor UO_407 (O_407,N_9272,N_7052);
and UO_408 (O_408,N_9282,N_7111);
or UO_409 (O_409,N_8940,N_8462);
xor UO_410 (O_410,N_8962,N_5948);
nor UO_411 (O_411,N_7069,N_8472);
nor UO_412 (O_412,N_8829,N_7217);
and UO_413 (O_413,N_7970,N_9956);
nand UO_414 (O_414,N_6447,N_8320);
nor UO_415 (O_415,N_8932,N_5134);
nand UO_416 (O_416,N_5921,N_8187);
xor UO_417 (O_417,N_9883,N_8573);
or UO_418 (O_418,N_7915,N_5841);
and UO_419 (O_419,N_9320,N_5555);
and UO_420 (O_420,N_5221,N_7013);
nor UO_421 (O_421,N_9068,N_9769);
nand UO_422 (O_422,N_5329,N_6903);
or UO_423 (O_423,N_5852,N_7363);
or UO_424 (O_424,N_5901,N_8917);
nor UO_425 (O_425,N_6113,N_9084);
nor UO_426 (O_426,N_9323,N_7624);
or UO_427 (O_427,N_9998,N_5570);
and UO_428 (O_428,N_6849,N_7565);
and UO_429 (O_429,N_7796,N_8006);
or UO_430 (O_430,N_5218,N_8011);
nor UO_431 (O_431,N_9598,N_5279);
nor UO_432 (O_432,N_7818,N_8198);
or UO_433 (O_433,N_6220,N_5490);
and UO_434 (O_434,N_6867,N_9855);
nand UO_435 (O_435,N_5138,N_7948);
or UO_436 (O_436,N_9683,N_9180);
nand UO_437 (O_437,N_9029,N_7842);
nor UO_438 (O_438,N_9187,N_8355);
or UO_439 (O_439,N_7271,N_7375);
nor UO_440 (O_440,N_5652,N_9270);
or UO_441 (O_441,N_6745,N_5331);
xnor UO_442 (O_442,N_9250,N_9897);
or UO_443 (O_443,N_7623,N_7969);
nor UO_444 (O_444,N_5043,N_9770);
nor UO_445 (O_445,N_8578,N_7507);
and UO_446 (O_446,N_6894,N_5367);
and UO_447 (O_447,N_6610,N_7450);
nor UO_448 (O_448,N_9365,N_8649);
or UO_449 (O_449,N_5365,N_5789);
and UO_450 (O_450,N_9974,N_9381);
or UO_451 (O_451,N_5591,N_7050);
and UO_452 (O_452,N_6882,N_7064);
nor UO_453 (O_453,N_5424,N_6665);
nand UO_454 (O_454,N_6557,N_8113);
or UO_455 (O_455,N_8724,N_6109);
xor UO_456 (O_456,N_6284,N_6054);
xor UO_457 (O_457,N_7251,N_8918);
and UO_458 (O_458,N_9220,N_7238);
xor UO_459 (O_459,N_5153,N_7667);
nand UO_460 (O_460,N_5671,N_6224);
nor UO_461 (O_461,N_8987,N_8959);
nand UO_462 (O_462,N_5886,N_8402);
or UO_463 (O_463,N_8245,N_6563);
or UO_464 (O_464,N_9767,N_6346);
and UO_465 (O_465,N_6604,N_8638);
and UO_466 (O_466,N_6380,N_8474);
nand UO_467 (O_467,N_8549,N_7135);
nor UO_468 (O_468,N_9529,N_5653);
nor UO_469 (O_469,N_5230,N_6013);
nor UO_470 (O_470,N_5412,N_7105);
nand UO_471 (O_471,N_7301,N_5870);
and UO_472 (O_472,N_5602,N_6839);
nand UO_473 (O_473,N_8673,N_6865);
and UO_474 (O_474,N_8236,N_9870);
and UO_475 (O_475,N_5536,N_8035);
nand UO_476 (O_476,N_8334,N_8715);
or UO_477 (O_477,N_7239,N_8372);
nand UO_478 (O_478,N_5601,N_9379);
xor UO_479 (O_479,N_9567,N_6804);
or UO_480 (O_480,N_8650,N_5587);
or UO_481 (O_481,N_7326,N_6898);
and UO_482 (O_482,N_6821,N_6657);
nand UO_483 (O_483,N_6426,N_9590);
xor UO_484 (O_484,N_6838,N_5720);
and UO_485 (O_485,N_8619,N_8374);
nor UO_486 (O_486,N_5592,N_5950);
or UO_487 (O_487,N_8155,N_7821);
xnor UO_488 (O_488,N_7788,N_7479);
nor UO_489 (O_489,N_5969,N_5702);
nor UO_490 (O_490,N_6216,N_6442);
nand UO_491 (O_491,N_8300,N_7539);
or UO_492 (O_492,N_8906,N_5946);
or UO_493 (O_493,N_8403,N_8737);
and UO_494 (O_494,N_6061,N_8590);
or UO_495 (O_495,N_5696,N_9439);
and UO_496 (O_496,N_7435,N_9281);
nand UO_497 (O_497,N_5916,N_7063);
nand UO_498 (O_498,N_5157,N_9061);
nor UO_499 (O_499,N_8912,N_9002);
and UO_500 (O_500,N_9488,N_8542);
nand UO_501 (O_501,N_8330,N_6588);
nand UO_502 (O_502,N_7185,N_7269);
and UO_503 (O_503,N_6974,N_8565);
or UO_504 (O_504,N_7765,N_7505);
nand UO_505 (O_505,N_7711,N_9936);
and UO_506 (O_506,N_8235,N_9809);
or UO_507 (O_507,N_5648,N_8891);
or UO_508 (O_508,N_6338,N_9255);
and UO_509 (O_509,N_8207,N_9489);
or UO_510 (O_510,N_6412,N_9563);
or UO_511 (O_511,N_6972,N_8294);
and UO_512 (O_512,N_5438,N_9446);
nor UO_513 (O_513,N_6062,N_6146);
nand UO_514 (O_514,N_7572,N_8032);
or UO_515 (O_515,N_6876,N_7025);
and UO_516 (O_516,N_5983,N_8013);
and UO_517 (O_517,N_5522,N_6213);
xor UO_518 (O_518,N_6377,N_7303);
and UO_519 (O_519,N_7390,N_6045);
nand UO_520 (O_520,N_6005,N_9942);
and UO_521 (O_521,N_6490,N_9456);
and UO_522 (O_522,N_9470,N_6368);
and UO_523 (O_523,N_9139,N_6723);
nor UO_524 (O_524,N_8316,N_5521);
or UO_525 (O_525,N_6085,N_8996);
and UO_526 (O_526,N_8232,N_7626);
nand UO_527 (O_527,N_6407,N_6067);
and UO_528 (O_528,N_6937,N_7474);
nor UO_529 (O_529,N_8407,N_5315);
nand UO_530 (O_530,N_5265,N_9636);
nand UO_531 (O_531,N_9053,N_7346);
nand UO_532 (O_532,N_8288,N_7910);
and UO_533 (O_533,N_9525,N_5836);
and UO_534 (O_534,N_6121,N_9492);
and UO_535 (O_535,N_7261,N_6414);
and UO_536 (O_536,N_9520,N_6065);
nand UO_537 (O_537,N_9929,N_7555);
and UO_538 (O_538,N_9127,N_9343);
nor UO_539 (O_539,N_7576,N_6949);
nand UO_540 (O_540,N_6993,N_7950);
nor UO_541 (O_541,N_9955,N_5262);
xor UO_542 (O_542,N_9960,N_6966);
nand UO_543 (O_543,N_7424,N_8210);
and UO_544 (O_544,N_7092,N_8344);
xor UO_545 (O_545,N_8784,N_5477);
or UO_546 (O_546,N_8148,N_6634);
xnor UO_547 (O_547,N_9449,N_7924);
nor UO_548 (O_548,N_8093,N_8272);
or UO_549 (O_549,N_9045,N_7551);
and UO_550 (O_550,N_8831,N_6315);
or UO_551 (O_551,N_9975,N_7080);
and UO_552 (O_552,N_9653,N_7202);
and UO_553 (O_553,N_6307,N_5629);
nand UO_554 (O_554,N_7570,N_9964);
or UO_555 (O_555,N_6249,N_7825);
and UO_556 (O_556,N_6183,N_9012);
xnor UO_557 (O_557,N_5363,N_9862);
nand UO_558 (O_558,N_8666,N_5459);
and UO_559 (O_559,N_9724,N_6845);
and UO_560 (O_560,N_9824,N_6817);
and UO_561 (O_561,N_5177,N_9415);
or UO_562 (O_562,N_8205,N_8162);
nor UO_563 (O_563,N_6330,N_8634);
nand UO_564 (O_564,N_9067,N_9686);
nor UO_565 (O_565,N_5274,N_8779);
or UO_566 (O_566,N_9941,N_9617);
and UO_567 (O_567,N_5405,N_7290);
and UO_568 (O_568,N_9411,N_8583);
or UO_569 (O_569,N_9841,N_5442);
nor UO_570 (O_570,N_9832,N_8208);
nor UO_571 (O_571,N_7055,N_9089);
and UO_572 (O_572,N_5923,N_5169);
and UO_573 (O_573,N_9663,N_5117);
or UO_574 (O_574,N_6160,N_6983);
xnor UO_575 (O_575,N_5156,N_9838);
or UO_576 (O_576,N_5217,N_7218);
and UO_577 (O_577,N_8313,N_9610);
nand UO_578 (O_578,N_5710,N_8277);
nand UO_579 (O_579,N_9716,N_8020);
nand UO_580 (O_580,N_8192,N_8998);
and UO_581 (O_581,N_5088,N_6214);
or UO_582 (O_582,N_5576,N_9513);
xor UO_583 (O_583,N_8740,N_6091);
nand UO_584 (O_584,N_8044,N_9659);
nor UO_585 (O_585,N_9179,N_6869);
nand UO_586 (O_586,N_7840,N_9399);
nor UO_587 (O_587,N_8875,N_6033);
or UO_588 (O_588,N_6678,N_5097);
or UO_589 (O_589,N_8612,N_7221);
or UO_590 (O_590,N_8486,N_6551);
nand UO_591 (O_591,N_5330,N_7643);
and UO_592 (O_592,N_8789,N_9758);
and UO_593 (O_593,N_7388,N_6628);
or UO_594 (O_594,N_6217,N_6743);
nand UO_595 (O_595,N_6922,N_8830);
nand UO_596 (O_596,N_7940,N_9306);
and UO_597 (O_597,N_8337,N_9150);
nand UO_598 (O_598,N_6792,N_8026);
or UO_599 (O_599,N_5435,N_8066);
nor UO_600 (O_600,N_9641,N_8053);
or UO_601 (O_601,N_6110,N_7094);
nand UO_602 (O_602,N_6353,N_6268);
nand UO_603 (O_603,N_6398,N_8237);
nand UO_604 (O_604,N_7543,N_7535);
and UO_605 (O_605,N_6750,N_6708);
xnor UO_606 (O_606,N_9842,N_8360);
nor UO_607 (O_607,N_8748,N_7406);
nor UO_608 (O_608,N_9839,N_7866);
nand UO_609 (O_609,N_9213,N_8338);
or UO_610 (O_610,N_7568,N_6077);
nor UO_611 (O_611,N_7465,N_6989);
nor UO_612 (O_612,N_8546,N_6429);
or UO_613 (O_613,N_5892,N_9120);
or UO_614 (O_614,N_9799,N_8808);
and UO_615 (O_615,N_6370,N_7312);
xnor UO_616 (O_616,N_6512,N_9774);
and UO_617 (O_617,N_6724,N_9556);
or UO_618 (O_618,N_9793,N_8792);
or UO_619 (O_619,N_7668,N_8818);
nor UO_620 (O_620,N_6396,N_8072);
and UO_621 (O_621,N_8392,N_7717);
nor UO_622 (O_622,N_5312,N_6906);
and UO_623 (O_623,N_8952,N_8504);
xor UO_624 (O_624,N_9021,N_8279);
xnor UO_625 (O_625,N_5718,N_9637);
xnor UO_626 (O_626,N_5190,N_9235);
nor UO_627 (O_627,N_8588,N_7102);
or UO_628 (O_628,N_5603,N_5270);
xor UO_629 (O_629,N_8105,N_7928);
nor UO_630 (O_630,N_6668,N_8973);
nor UO_631 (O_631,N_9888,N_7661);
or UO_632 (O_632,N_8657,N_5249);
nand UO_633 (O_633,N_8544,N_5949);
nor UO_634 (O_634,N_9742,N_8812);
and UO_635 (O_635,N_8828,N_6748);
nor UO_636 (O_636,N_5589,N_9298);
nand UO_637 (O_637,N_6629,N_8507);
nor UO_638 (O_638,N_6423,N_5783);
or UO_639 (O_639,N_5192,N_5518);
nand UO_640 (O_640,N_7891,N_6987);
nor UO_641 (O_641,N_7787,N_9764);
and UO_642 (O_642,N_9276,N_8640);
nor UO_643 (O_643,N_8074,N_5278);
nand UO_644 (O_644,N_5204,N_5818);
nor UO_645 (O_645,N_8846,N_7430);
nand UO_646 (O_646,N_9069,N_6421);
or UO_647 (O_647,N_9370,N_6952);
and UO_648 (O_648,N_9715,N_5171);
nor UO_649 (O_649,N_6929,N_8676);
nand UO_650 (O_650,N_6116,N_7811);
or UO_651 (O_651,N_8641,N_7530);
nand UO_652 (O_652,N_8089,N_9407);
nor UO_653 (O_653,N_8943,N_9091);
xnor UO_654 (O_654,N_8671,N_5445);
xnor UO_655 (O_655,N_8297,N_6463);
nor UO_656 (O_656,N_8097,N_7123);
nand UO_657 (O_657,N_7806,N_5334);
nor UO_658 (O_658,N_9795,N_7145);
or UO_659 (O_659,N_8804,N_9345);
or UO_660 (O_660,N_8495,N_9904);
or UO_661 (O_661,N_7857,N_9722);
nand UO_662 (O_662,N_5007,N_9658);
nand UO_663 (O_663,N_6397,N_7189);
nor UO_664 (O_664,N_8061,N_8622);
and UO_665 (O_665,N_6539,N_7345);
nand UO_666 (O_666,N_6915,N_6607);
xor UO_667 (O_667,N_8561,N_6856);
nor UO_668 (O_668,N_7669,N_8249);
or UO_669 (O_669,N_7334,N_9156);
nor UO_670 (O_670,N_7781,N_9145);
xnor UO_671 (O_671,N_8581,N_7754);
nor UO_672 (O_672,N_6765,N_5041);
or UO_673 (O_673,N_9126,N_8477);
xnor UO_674 (O_674,N_5144,N_6714);
and UO_675 (O_675,N_9560,N_5552);
or UO_676 (O_676,N_8368,N_5880);
nand UO_677 (O_677,N_5251,N_5756);
and UO_678 (O_678,N_9386,N_7720);
and UO_679 (O_679,N_5324,N_9966);
and UO_680 (O_680,N_6675,N_7204);
and UO_681 (O_681,N_5819,N_8525);
nor UO_682 (O_682,N_5377,N_7200);
nand UO_683 (O_683,N_5214,N_5636);
or UO_684 (O_684,N_5044,N_5300);
and UO_685 (O_685,N_6060,N_5731);
or UO_686 (O_686,N_8976,N_7722);
or UO_687 (O_687,N_9093,N_8848);
xor UO_688 (O_688,N_7405,N_7892);
nor UO_689 (O_689,N_8385,N_7000);
xor UO_690 (O_690,N_7057,N_7959);
nand UO_691 (O_691,N_6647,N_8774);
nand UO_692 (O_692,N_9215,N_9342);
and UO_693 (O_693,N_7646,N_5582);
and UO_694 (O_694,N_5807,N_8161);
or UO_695 (O_695,N_9236,N_5340);
nor UO_696 (O_696,N_8111,N_6468);
and UO_697 (O_697,N_5686,N_9186);
nand UO_698 (O_698,N_5910,N_6643);
nand UO_699 (O_699,N_8886,N_6488);
nand UO_700 (O_700,N_5201,N_9279);
and UO_701 (O_701,N_7336,N_6895);
or UO_702 (O_702,N_5253,N_6126);
and UO_703 (O_703,N_5932,N_9578);
or UO_704 (O_704,N_5936,N_5154);
xor UO_705 (O_705,N_5754,N_7882);
nand UO_706 (O_706,N_9183,N_7357);
xor UO_707 (O_707,N_5139,N_8466);
nand UO_708 (O_708,N_9431,N_8541);
nand UO_709 (O_709,N_9763,N_8098);
or UO_710 (O_710,N_9269,N_5721);
nor UO_711 (O_711,N_6401,N_5297);
nor UO_712 (O_712,N_5666,N_9639);
and UO_713 (O_713,N_9574,N_5639);
nand UO_714 (O_714,N_7023,N_7112);
and UO_715 (O_715,N_9158,N_6436);
or UO_716 (O_716,N_9652,N_5486);
nor UO_717 (O_717,N_9747,N_8413);
nor UO_718 (O_718,N_8094,N_6877);
nor UO_719 (O_719,N_8859,N_9733);
and UO_720 (O_720,N_9755,N_8773);
xnor UO_721 (O_721,N_6208,N_5110);
or UO_722 (O_722,N_6498,N_9972);
nor UO_723 (O_723,N_5895,N_7077);
nand UO_724 (O_724,N_5817,N_8080);
or UO_725 (O_725,N_5121,N_6564);
and UO_726 (O_726,N_6493,N_6802);
nand UO_727 (O_727,N_9893,N_8048);
or UO_728 (O_728,N_7760,N_8104);
or UO_729 (O_729,N_8171,N_5668);
or UO_730 (O_730,N_8103,N_7296);
nor UO_731 (O_731,N_6662,N_9375);
nor UO_732 (O_732,N_6753,N_8130);
nand UO_733 (O_733,N_5752,N_9570);
nor UO_734 (O_734,N_8897,N_8690);
nor UO_735 (O_735,N_6384,N_9024);
or UO_736 (O_736,N_5956,N_7934);
nor UO_737 (O_737,N_7300,N_5531);
nand UO_738 (O_738,N_9871,N_5800);
and UO_739 (O_739,N_7943,N_6768);
nand UO_740 (O_740,N_8712,N_9757);
and UO_741 (O_741,N_5716,N_6659);
or UO_742 (O_742,N_8263,N_6870);
or UO_743 (O_743,N_6129,N_9057);
nor UO_744 (O_744,N_6207,N_9297);
and UO_745 (O_745,N_6884,N_7095);
nor UO_746 (O_746,N_8636,N_8869);
nand UO_747 (O_747,N_7427,N_5883);
and UO_748 (O_748,N_8377,N_9309);
nor UO_749 (O_749,N_6472,N_6159);
or UO_750 (O_750,N_9065,N_8539);
and UO_751 (O_751,N_7867,N_6964);
nor UO_752 (O_752,N_8231,N_7488);
and UO_753 (O_753,N_9423,N_7801);
and UO_754 (O_754,N_5175,N_8833);
nand UO_755 (O_755,N_7861,N_9015);
or UO_756 (O_756,N_7592,N_8763);
xor UO_757 (O_757,N_5205,N_7524);
or UO_758 (O_758,N_9576,N_8416);
nand UO_759 (O_759,N_8359,N_9499);
or UO_760 (O_760,N_6328,N_5712);
nor UO_761 (O_761,N_7142,N_8642);
or UO_762 (O_762,N_8821,N_8611);
and UO_763 (O_763,N_6018,N_5597);
nor UO_764 (O_764,N_8689,N_9649);
and UO_765 (O_765,N_8555,N_8647);
xnor UO_766 (O_766,N_6866,N_5113);
and UO_767 (O_767,N_7665,N_5455);
and UO_768 (O_768,N_8382,N_6536);
and UO_769 (O_769,N_7901,N_8770);
nand UO_770 (O_770,N_8795,N_9039);
nand UO_771 (O_771,N_7153,N_7654);
nor UO_772 (O_772,N_5035,N_6081);
xor UO_773 (O_773,N_8620,N_6164);
and UO_774 (O_774,N_5766,N_7101);
and UO_775 (O_775,N_6540,N_7152);
nand UO_776 (O_776,N_6674,N_8937);
xnor UO_777 (O_777,N_8075,N_7368);
or UO_778 (O_778,N_9464,N_9290);
nand UO_779 (O_779,N_8476,N_9383);
nand UO_780 (O_780,N_9430,N_6205);
nor UO_781 (O_781,N_5993,N_9532);
nor UO_782 (O_782,N_6615,N_7352);
and UO_783 (O_783,N_5015,N_9404);
nor UO_784 (O_784,N_6756,N_7800);
xnor UO_785 (O_785,N_5394,N_8376);
nor UO_786 (O_786,N_7734,N_7567);
or UO_787 (O_787,N_7499,N_7860);
and UO_788 (O_788,N_8438,N_5468);
and UO_789 (O_789,N_7575,N_9537);
and UO_790 (O_790,N_9635,N_6526);
nand UO_791 (O_791,N_6625,N_5768);
nand UO_792 (O_792,N_9479,N_8551);
nor UO_793 (O_793,N_8308,N_9886);
or UO_794 (O_794,N_7003,N_6100);
nor UO_795 (O_795,N_7513,N_8807);
nand UO_796 (O_796,N_7476,N_8491);
or UO_797 (O_797,N_6916,N_5701);
nor UO_798 (O_798,N_8000,N_7620);
xor UO_799 (O_799,N_9687,N_9315);
xnor UO_800 (O_800,N_7385,N_9978);
and UO_801 (O_801,N_9884,N_5705);
nor UO_802 (O_802,N_7360,N_6799);
or UO_803 (O_803,N_9746,N_5853);
nand UO_804 (O_804,N_6677,N_7446);
nand UO_805 (O_805,N_9668,N_5160);
and UO_806 (O_806,N_6043,N_8096);
nand UO_807 (O_807,N_9217,N_8115);
and UO_808 (O_808,N_8140,N_7638);
and UO_809 (O_809,N_6069,N_9422);
nand UO_810 (O_810,N_5610,N_7553);
or UO_811 (O_811,N_7079,N_6296);
and UO_812 (O_812,N_7018,N_8214);
and UO_813 (O_813,N_7282,N_8435);
and UO_814 (O_814,N_9614,N_5092);
nor UO_815 (O_815,N_7214,N_7466);
and UO_816 (O_816,N_9133,N_6097);
nand UO_817 (O_817,N_7502,N_6506);
xnor UO_818 (O_818,N_7322,N_6132);
and UO_819 (O_819,N_6042,N_6519);
or UO_820 (O_820,N_7026,N_7652);
or UO_821 (O_821,N_8796,N_5894);
nand UO_822 (O_822,N_6051,N_5254);
nand UO_823 (O_823,N_9317,N_8723);
nor UO_824 (O_824,N_6681,N_8468);
nand UO_825 (O_825,N_9818,N_9648);
nand UO_826 (O_826,N_9007,N_8615);
nand UO_827 (O_827,N_7475,N_8920);
nor UO_828 (O_828,N_8603,N_7588);
nor UO_829 (O_829,N_5926,N_8945);
nand UO_830 (O_830,N_7199,N_8287);
nand UO_831 (O_831,N_5290,N_9027);
nor UO_832 (O_832,N_7289,N_8473);
nand UO_833 (O_833,N_6685,N_7240);
nand UO_834 (O_834,N_9607,N_7019);
or UO_835 (O_835,N_9690,N_8537);
nand UO_836 (O_836,N_5925,N_5679);
xnor UO_837 (O_837,N_7137,N_5220);
xor UO_838 (O_838,N_8354,N_8580);
nor UO_839 (O_839,N_7213,N_5240);
xor UO_840 (O_840,N_8769,N_5982);
nor UO_841 (O_841,N_6948,N_6297);
and UO_842 (O_842,N_6434,N_7723);
and UO_843 (O_843,N_8055,N_8684);
or UO_844 (O_844,N_6927,N_5385);
nand UO_845 (O_845,N_7673,N_9730);
nand UO_846 (O_846,N_9700,N_5319);
or UO_847 (O_847,N_5887,N_5090);
or UO_848 (O_848,N_5888,N_9968);
nor UO_849 (O_849,N_6975,N_9487);
nor UO_850 (O_850,N_7319,N_9958);
nand UO_851 (O_851,N_8414,N_7992);
and UO_852 (O_852,N_7131,N_9174);
nand UO_853 (O_853,N_6221,N_7791);
and UO_854 (O_854,N_9494,N_6521);
xnor UO_855 (O_855,N_8972,N_5493);
and UO_856 (O_856,N_5532,N_8022);
nor UO_857 (O_857,N_6094,N_6967);
nor UO_858 (O_858,N_7864,N_8116);
and UO_859 (O_859,N_9362,N_7084);
xnor UO_860 (O_860,N_8042,N_7698);
nor UO_861 (O_861,N_9743,N_9459);
xor UO_862 (O_862,N_5343,N_7608);
nor UO_863 (O_863,N_7912,N_8211);
or UO_864 (O_864,N_7274,N_5772);
and UO_865 (O_865,N_7556,N_9784);
or UO_866 (O_866,N_7297,N_6875);
or UO_867 (O_867,N_6292,N_8086);
nand UO_868 (O_868,N_6302,N_6161);
nand UO_869 (O_869,N_8882,N_9003);
and UO_870 (O_870,N_8131,N_9630);
nand UO_871 (O_871,N_8730,N_8343);
and UO_872 (O_872,N_9969,N_7459);
and UO_873 (O_873,N_8698,N_5261);
nor UO_874 (O_874,N_8434,N_9670);
or UO_875 (O_875,N_7509,N_8591);
and UO_876 (O_876,N_6676,N_9553);
nand UO_877 (O_877,N_7320,N_6320);
and UO_878 (O_878,N_6237,N_7500);
nor UO_879 (O_879,N_6758,N_7980);
xor UO_880 (O_880,N_9765,N_8134);
nor UO_881 (O_881,N_9377,N_7332);
or UO_882 (O_882,N_8128,N_7594);
xor UO_883 (O_883,N_5830,N_5130);
nand UO_884 (O_884,N_8421,N_7027);
nand UO_885 (O_885,N_9354,N_7362);
or UO_886 (O_886,N_5778,N_6535);
and UO_887 (O_887,N_8974,N_6027);
nor UO_888 (O_888,N_6600,N_8872);
and UO_889 (O_889,N_5325,N_8713);
or UO_890 (O_890,N_9771,N_7009);
nor UO_891 (O_891,N_7932,N_9921);
nor UO_892 (O_892,N_8225,N_5129);
and UO_893 (O_893,N_8030,N_9689);
or UO_894 (O_894,N_8056,N_9667);
nor UO_895 (O_895,N_9080,N_8206);
and UO_896 (O_896,N_5181,N_8129);
xnor UO_897 (O_897,N_8318,N_8101);
nand UO_898 (O_898,N_6111,N_9885);
nand UO_899 (O_899,N_9548,N_5170);
and UO_900 (O_900,N_8655,N_8700);
nand UO_901 (O_901,N_7042,N_6638);
nor UO_902 (O_902,N_9094,N_9695);
nand UO_903 (O_903,N_9502,N_7411);
xnor UO_904 (O_904,N_9227,N_7755);
and UO_905 (O_905,N_6958,N_5105);
nand UO_906 (O_906,N_7232,N_9602);
and UO_907 (O_907,N_8703,N_7087);
nand UO_908 (O_908,N_8078,N_7284);
xor UO_909 (O_909,N_8255,N_8512);
nor UO_910 (O_910,N_5945,N_5148);
nor UO_911 (O_911,N_9189,N_6385);
nor UO_912 (O_912,N_9336,N_5937);
nor UO_913 (O_913,N_5374,N_7835);
nand UO_914 (O_914,N_9391,N_5111);
nor UO_915 (O_915,N_7807,N_9727);
and UO_916 (O_916,N_7888,N_6605);
and UO_917 (O_917,N_8806,N_9263);
nand UO_918 (O_918,N_6715,N_9822);
nand UO_919 (O_919,N_6028,N_8488);
nand UO_920 (O_920,N_8244,N_7743);
and UO_921 (O_921,N_5802,N_5417);
xnor UO_922 (O_922,N_9169,N_6961);
nand UO_923 (O_923,N_7350,N_7122);
nor UO_924 (O_924,N_7921,N_8400);
and UO_925 (O_925,N_7181,N_9527);
and UO_926 (O_926,N_9646,N_6050);
or UO_927 (O_927,N_5959,N_9712);
or UO_928 (O_928,N_9675,N_9274);
and UO_929 (O_929,N_8280,N_5940);
or UO_930 (O_930,N_6347,N_9935);
and UO_931 (O_931,N_6788,N_7398);
or UO_932 (O_932,N_7895,N_6011);
and UO_933 (O_933,N_7295,N_5371);
and UO_934 (O_934,N_6679,N_6416);
nand UO_935 (O_935,N_6259,N_5382);
and UO_936 (O_936,N_7418,N_6167);
nand UO_937 (O_937,N_7038,N_6886);
or UO_938 (O_938,N_9041,N_5875);
and UO_939 (O_939,N_9997,N_6592);
xor UO_940 (O_940,N_8005,N_8265);
and UO_941 (O_941,N_9660,N_6010);
and UO_942 (O_942,N_7955,N_5619);
nor UO_943 (O_943,N_9249,N_8274);
or UO_944 (O_944,N_8605,N_5431);
nor UO_945 (O_945,N_5577,N_9076);
nand UO_946 (O_946,N_7560,N_9545);
and UO_947 (O_947,N_6378,N_9144);
and UO_948 (O_948,N_8721,N_9922);
nor UO_949 (O_949,N_9152,N_5893);
nor UO_950 (O_950,N_5039,N_7817);
nand UO_951 (O_951,N_8241,N_6760);
nand UO_952 (O_952,N_9943,N_9725);
or UO_953 (O_953,N_6688,N_9846);
xor UO_954 (O_954,N_9171,N_9147);
nor UO_955 (O_955,N_7750,N_6965);
xor UO_956 (O_956,N_9330,N_9059);
xor UO_957 (O_957,N_7104,N_9445);
nand UO_958 (O_958,N_7585,N_7508);
or UO_959 (O_959,N_9010,N_5372);
and UO_960 (O_960,N_8375,N_5485);
xor UO_961 (O_961,N_6543,N_9834);
nor UO_962 (O_962,N_8532,N_7764);
or UO_963 (O_963,N_8485,N_5093);
or UO_964 (O_964,N_7419,N_9122);
or UO_965 (O_965,N_5058,N_7276);
and UO_966 (O_966,N_6885,N_6441);
or UO_967 (O_967,N_5974,N_9437);
and UO_968 (O_968,N_7062,N_8281);
nand UO_969 (O_969,N_9803,N_5285);
and UO_970 (O_970,N_6435,N_5680);
nand UO_971 (O_971,N_6816,N_6264);
xor UO_972 (O_972,N_9741,N_7461);
xnor UO_973 (O_973,N_5782,N_5391);
xor UO_974 (O_974,N_5611,N_8566);
nor UO_975 (O_975,N_8197,N_9530);
nand UO_976 (O_976,N_7971,N_8853);
xnor UO_977 (O_977,N_8600,N_7642);
nor UO_978 (O_978,N_5728,N_8340);
nor UO_979 (O_979,N_5534,N_6369);
nor UO_980 (O_980,N_6454,N_6140);
or UO_981 (O_981,N_8260,N_9679);
nor UO_982 (O_982,N_7695,N_7721);
and UO_983 (O_983,N_6741,N_7559);
xor UO_984 (O_984,N_7414,N_9814);
and UO_985 (O_985,N_6938,N_9098);
nor UO_986 (O_986,N_5524,N_9095);
and UO_987 (O_987,N_7451,N_6495);
or UO_988 (O_988,N_8720,N_9325);
or UO_989 (O_989,N_8123,N_7967);
nand UO_990 (O_990,N_9995,N_8589);
or UO_991 (O_991,N_5810,N_9218);
and UO_992 (O_992,N_8227,N_9714);
nand UO_993 (O_993,N_9994,N_8879);
xnor UO_994 (O_994,N_6601,N_7273);
xnor UO_995 (O_995,N_5223,N_9484);
and UO_996 (O_996,N_7082,N_6784);
nand UO_997 (O_997,N_6988,N_9229);
or UO_998 (O_998,N_9099,N_6641);
nor UO_999 (O_999,N_6861,N_5976);
nor UO_1000 (O_1000,N_5462,N_5906);
nor UO_1001 (O_1001,N_7262,N_7923);
xnor UO_1002 (O_1002,N_9109,N_6763);
nor UO_1003 (O_1003,N_7752,N_9123);
nor UO_1004 (O_1004,N_9414,N_9376);
and UO_1005 (O_1005,N_6749,N_6603);
and UO_1006 (O_1006,N_8938,N_5470);
or UO_1007 (O_1007,N_7635,N_5439);
and UO_1008 (O_1008,N_7233,N_9254);
and UO_1009 (O_1009,N_9164,N_9155);
nor UO_1010 (O_1010,N_9341,N_5425);
or UO_1011 (O_1011,N_5072,N_9087);
or UO_1012 (O_1012,N_6174,N_7735);
or UO_1013 (O_1013,N_7283,N_9808);
and UO_1014 (O_1014,N_9564,N_8063);
or UO_1015 (O_1015,N_6880,N_9597);
and UO_1016 (O_1016,N_7958,N_6890);
nand UO_1017 (O_1017,N_8068,N_5657);
and UO_1018 (O_1018,N_5258,N_5839);
and UO_1019 (O_1019,N_8680,N_9329);
and UO_1020 (O_1020,N_7945,N_7704);
or UO_1021 (O_1021,N_8301,N_5226);
and UO_1022 (O_1022,N_8363,N_9951);
and UO_1023 (O_1023,N_7964,N_7367);
nand UO_1024 (O_1024,N_5320,N_8991);
or UO_1025 (O_1025,N_6698,N_8884);
nor UO_1026 (O_1026,N_8610,N_9588);
or UO_1027 (O_1027,N_6507,N_7211);
or UO_1028 (O_1028,N_5432,N_6699);
nand UO_1029 (O_1029,N_7603,N_9294);
nand UO_1030 (O_1030,N_6547,N_6640);
or UO_1031 (O_1031,N_9314,N_8717);
nand UO_1032 (O_1032,N_6086,N_8738);
or UO_1033 (O_1033,N_5890,N_5188);
and UO_1034 (O_1034,N_9490,N_5159);
and UO_1035 (O_1035,N_8405,N_8847);
or UO_1036 (O_1036,N_5102,N_5402);
nor UO_1037 (O_1037,N_5443,N_9810);
nand UO_1038 (O_1038,N_7587,N_6854);
or UO_1039 (O_1039,N_7522,N_6194);
or UO_1040 (O_1040,N_8404,N_6561);
or UO_1041 (O_1041,N_7827,N_7884);
or UO_1042 (O_1042,N_7160,N_6968);
and UO_1043 (O_1043,N_5487,N_5164);
xor UO_1044 (O_1044,N_5345,N_6803);
xor UO_1045 (O_1045,N_9170,N_8810);
nand UO_1046 (O_1046,N_7329,N_6462);
xnor UO_1047 (O_1047,N_5546,N_9406);
or UO_1048 (O_1048,N_6188,N_5627);
nor UO_1049 (O_1049,N_7753,N_7183);
nor UO_1050 (O_1050,N_6182,N_6868);
nand UO_1051 (O_1051,N_7146,N_7829);
or UO_1052 (O_1052,N_7700,N_9036);
and UO_1053 (O_1053,N_8914,N_5775);
xnor UO_1054 (O_1054,N_7615,N_6088);
xnor UO_1055 (O_1055,N_6797,N_8613);
and UO_1056 (O_1056,N_6093,N_7339);
or UO_1057 (O_1057,N_9766,N_7184);
xnor UO_1058 (O_1058,N_7178,N_7440);
and UO_1059 (O_1059,N_5291,N_7212);
nand UO_1060 (O_1060,N_6783,N_9971);
xnor UO_1061 (O_1061,N_8850,N_6405);
nor UO_1062 (O_1062,N_5743,N_9583);
nand UO_1063 (O_1063,N_6589,N_7812);
and UO_1064 (O_1064,N_5741,N_7705);
or UO_1065 (O_1065,N_5420,N_5934);
xor UO_1066 (O_1066,N_7248,N_9208);
xnor UO_1067 (O_1067,N_5299,N_7756);
and UO_1068 (O_1068,N_6263,N_5519);
xor UO_1069 (O_1069,N_5547,N_8907);
nand UO_1070 (O_1070,N_5128,N_5687);
or UO_1071 (O_1071,N_7636,N_9547);
nor UO_1072 (O_1072,N_8201,N_6331);
nand UO_1073 (O_1073,N_6560,N_5797);
nand UO_1074 (O_1074,N_7933,N_7383);
nand UO_1075 (O_1075,N_8656,N_7803);
and UO_1076 (O_1076,N_6645,N_7438);
and UO_1077 (O_1077,N_5053,N_9160);
and UO_1078 (O_1078,N_8644,N_9856);
and UO_1079 (O_1079,N_8880,N_9312);
and UO_1080 (O_1080,N_9072,N_9680);
nor UO_1081 (O_1081,N_7229,N_8456);
xor UO_1082 (O_1082,N_7192,N_6139);
nand UO_1083 (O_1083,N_8459,N_6819);
or UO_1084 (O_1084,N_8861,N_5933);
nand UO_1085 (O_1085,N_9051,N_6580);
and UO_1086 (O_1086,N_7528,N_8038);
nor UO_1087 (O_1087,N_7434,N_5467);
nand UO_1088 (O_1088,N_5541,N_7890);
nand UO_1089 (O_1089,N_5289,N_8487);
and UO_1090 (O_1090,N_8088,N_7979);
nand UO_1091 (O_1091,N_9246,N_6787);
and UO_1092 (O_1092,N_9603,N_5390);
and UO_1093 (O_1093,N_6177,N_5542);
xnor UO_1094 (O_1094,N_6452,N_9202);
nor UO_1095 (O_1095,N_6095,N_9693);
and UO_1096 (O_1096,N_5502,N_6785);
or UO_1097 (O_1097,N_7448,N_8373);
nor UO_1098 (O_1098,N_7637,N_8118);
nor UO_1099 (O_1099,N_5625,N_9736);
nor UO_1100 (O_1100,N_8475,N_7709);
nand UO_1101 (O_1101,N_9452,N_8827);
xor UO_1102 (O_1102,N_7810,N_9328);
and UO_1103 (O_1103,N_6879,N_7086);
nor UO_1104 (O_1104,N_8865,N_5986);
nor UO_1105 (O_1105,N_8948,N_8599);
and UO_1106 (O_1106,N_6118,N_6562);
nand UO_1107 (O_1107,N_8350,N_5392);
and UO_1108 (O_1108,N_7978,N_7408);
and UO_1109 (O_1109,N_8825,N_6782);
and UO_1110 (O_1110,N_6960,N_6813);
nand UO_1111 (O_1111,N_6970,N_9536);
xnor UO_1112 (O_1112,N_5622,N_5135);
or UO_1113 (O_1113,N_9207,N_8482);
or UO_1114 (O_1114,N_8173,N_9678);
or UO_1115 (O_1115,N_5550,N_6361);
nor UO_1116 (O_1116,N_5028,N_6335);
and UO_1117 (O_1117,N_6180,N_7304);
nor UO_1118 (O_1118,N_5284,N_5399);
or UO_1119 (O_1119,N_8560,N_5008);
or UO_1120 (O_1120,N_8411,N_5107);
or UO_1121 (O_1121,N_5700,N_9234);
and UO_1122 (O_1122,N_5361,N_8027);
and UO_1123 (O_1123,N_5647,N_5967);
nor UO_1124 (O_1124,N_7136,N_6686);
nand UO_1125 (O_1125,N_9666,N_6176);
nand UO_1126 (O_1126,N_5876,N_5746);
nor UO_1127 (O_1127,N_7372,N_9773);
nand UO_1128 (O_1128,N_8993,N_7908);
xnor UO_1129 (O_1129,N_5638,N_7885);
xor UO_1130 (O_1130,N_6052,N_5688);
xnor UO_1131 (O_1131,N_8726,N_8047);
and UO_1132 (O_1132,N_7072,N_9542);
xor UO_1133 (O_1133,N_6017,N_8509);
nor UO_1134 (O_1134,N_6204,N_5997);
nand UO_1135 (O_1135,N_8230,N_5504);
nor UO_1136 (O_1136,N_7512,N_9682);
nand UO_1137 (O_1137,N_5239,N_5585);
nand UO_1138 (O_1138,N_9079,N_7089);
or UO_1139 (O_1139,N_5821,N_8921);
or UO_1140 (O_1140,N_7759,N_9327);
nor UO_1141 (O_1141,N_5685,N_7707);
nand UO_1142 (O_1142,N_7206,N_6156);
nor UO_1143 (O_1143,N_7657,N_8204);
nand UO_1144 (O_1144,N_8735,N_8369);
or UO_1145 (O_1145,N_6940,N_6599);
and UO_1146 (O_1146,N_5397,N_7975);
nor UO_1147 (O_1147,N_8633,N_8143);
nor UO_1148 (O_1148,N_7544,N_7658);
xnor UO_1149 (O_1149,N_9114,N_5903);
nor UO_1150 (O_1150,N_7120,N_8783);
and UO_1151 (O_1151,N_7619,N_8947);
and UO_1152 (O_1152,N_5071,N_6808);
nand UO_1153 (O_1153,N_6671,N_8151);
or UO_1154 (O_1154,N_5583,N_9671);
nor UO_1155 (O_1155,N_7454,N_6102);
and UO_1156 (O_1156,N_7993,N_7371);
nand UO_1157 (O_1157,N_5834,N_5255);
and UO_1158 (O_1158,N_7098,N_8970);
or UO_1159 (O_1159,N_5593,N_5306);
and UO_1160 (O_1160,N_9301,N_8749);
nand UO_1161 (O_1161,N_8349,N_6707);
nand UO_1162 (O_1162,N_8714,N_8253);
and UO_1163 (O_1163,N_5004,N_7518);
nand UO_1164 (O_1164,N_7264,N_6336);
and UO_1165 (O_1165,N_8771,N_9019);
xnor UO_1166 (O_1166,N_8332,N_6422);
and UO_1167 (O_1167,N_8866,N_6789);
nand UO_1168 (O_1168,N_9580,N_5571);
or UO_1169 (O_1169,N_6185,N_6984);
and UO_1170 (O_1170,N_6120,N_7046);
nor UO_1171 (O_1171,N_8559,N_5935);
or UO_1172 (O_1172,N_7863,N_8479);
and UO_1173 (O_1173,N_6673,N_9371);
and UO_1174 (O_1174,N_8944,N_5358);
or UO_1175 (O_1175,N_8502,N_8777);
xnor UO_1176 (O_1176,N_7843,N_9776);
or UO_1177 (O_1177,N_8290,N_7349);
nand UO_1178 (O_1178,N_5806,N_6319);
and UO_1179 (O_1179,N_9115,N_8729);
or UO_1180 (O_1180,N_9976,N_5747);
and UO_1181 (O_1181,N_6574,N_5065);
or UO_1182 (O_1182,N_9260,N_6192);
and UO_1183 (O_1183,N_6585,N_9275);
nor UO_1184 (O_1184,N_8024,N_9761);
nand UO_1185 (O_1185,N_5375,N_6718);
or UO_1186 (O_1186,N_5237,N_9338);
xnor UO_1187 (O_1187,N_9121,N_5829);
and UO_1188 (O_1188,N_7586,N_6227);
nand UO_1189 (O_1189,N_5640,N_7726);
and UO_1190 (O_1190,N_6606,N_6294);
nand UO_1191 (O_1191,N_8905,N_7030);
or UO_1192 (O_1192,N_7157,N_8406);
and UO_1193 (O_1193,N_8572,N_8696);
xor UO_1194 (O_1194,N_6947,N_5557);
and UO_1195 (O_1195,N_7498,N_5250);
nor UO_1196 (O_1196,N_8496,N_8395);
and UO_1197 (O_1197,N_8685,N_6304);
nor UO_1198 (O_1198,N_6285,N_8267);
and UO_1199 (O_1199,N_9424,N_7925);
xnor UO_1200 (O_1200,N_8968,N_8133);
nor UO_1201 (O_1201,N_7358,N_5777);
and UO_1202 (O_1202,N_7313,N_6702);
nand UO_1203 (O_1203,N_9172,N_8417);
nand UO_1204 (O_1204,N_7472,N_5715);
and UO_1205 (O_1205,N_8481,N_8702);
nand UO_1206 (O_1206,N_8533,N_9711);
nor UO_1207 (O_1207,N_8926,N_5150);
nor UO_1208 (O_1208,N_8218,N_7852);
and UO_1209 (O_1209,N_9008,N_6329);
nand UO_1210 (O_1210,N_5147,N_7681);
xnor UO_1211 (O_1211,N_7059,N_7182);
or UO_1212 (O_1212,N_8217,N_9555);
nand UO_1213 (O_1213,N_8706,N_9698);
or UO_1214 (O_1214,N_9349,N_9473);
and UO_1215 (O_1215,N_7872,N_7324);
xnor UO_1216 (O_1216,N_5145,N_8107);
and UO_1217 (O_1217,N_8986,N_7495);
nor UO_1218 (O_1218,N_6862,N_6410);
xor UO_1219 (O_1219,N_5469,N_9367);
nand UO_1220 (O_1220,N_7784,N_9066);
and UO_1221 (O_1221,N_9581,N_8592);
nor UO_1222 (O_1222,N_6492,N_8904);
and UO_1223 (O_1223,N_5276,N_8073);
or UO_1224 (O_1224,N_8333,N_5225);
nor UO_1225 (O_1225,N_8790,N_9110);
or UO_1226 (O_1226,N_5617,N_5457);
or UO_1227 (O_1227,N_6917,N_8992);
or UO_1228 (O_1228,N_5056,N_8758);
nor UO_1229 (O_1229,N_7672,N_6262);
nor UO_1230 (O_1230,N_6274,N_7645);
or UO_1231 (O_1231,N_6367,N_8138);
nor UO_1232 (O_1232,N_7896,N_6658);
and UO_1233 (O_1233,N_9552,N_8518);
xnor UO_1234 (O_1234,N_5180,N_9428);
and UO_1235 (O_1235,N_8295,N_9390);
nor UO_1236 (O_1236,N_8780,N_7452);
and UO_1237 (O_1237,N_6058,N_6233);
and UO_1238 (O_1238,N_5736,N_7412);
and UO_1239 (O_1239,N_8543,N_9288);
and UO_1240 (O_1240,N_6340,N_6134);
nand UO_1241 (O_1241,N_8707,N_9347);
nand UO_1242 (O_1242,N_9028,N_8181);
and UO_1243 (O_1243,N_7799,N_7355);
or UO_1244 (O_1244,N_7670,N_9827);
nand UO_1245 (O_1245,N_7916,N_8077);
nor UO_1246 (O_1246,N_9775,N_5847);
nor UO_1247 (O_1247,N_8860,N_6691);
or UO_1248 (O_1248,N_6841,N_5409);
nor UO_1249 (O_1249,N_5362,N_7342);
nor UO_1250 (O_1250,N_9086,N_7293);
nor UO_1251 (O_1251,N_6290,N_7016);
or UO_1252 (O_1252,N_8966,N_8234);
nand UO_1253 (O_1253,N_8654,N_5423);
or UO_1254 (O_1254,N_8383,N_6534);
nor UO_1255 (O_1255,N_7380,N_9783);
nor UO_1256 (O_1256,N_8202,N_9326);
nor UO_1257 (O_1257,N_8900,N_8233);
or UO_1258 (O_1258,N_9461,N_7690);
nor UO_1259 (O_1259,N_9468,N_7090);
nand UO_1260 (O_1260,N_7991,N_5030);
nor UO_1261 (O_1261,N_6272,N_5843);
nor UO_1262 (O_1262,N_9360,N_8498);
xnor UO_1263 (O_1263,N_9285,N_8817);
and UO_1264 (O_1264,N_7718,N_5427);
nand UO_1265 (O_1265,N_5898,N_7946);
nand UO_1266 (O_1266,N_6910,N_9804);
or UO_1267 (O_1267,N_6145,N_9162);
nor UO_1268 (O_1268,N_8084,N_5907);
or UO_1269 (O_1269,N_8137,N_6980);
and UO_1270 (O_1270,N_7651,N_8802);
and UO_1271 (O_1271,N_7230,N_8325);
and UO_1272 (O_1272,N_6528,N_5317);
nor UO_1273 (O_1273,N_7844,N_9606);
xnor UO_1274 (O_1274,N_9136,N_9847);
or UO_1275 (O_1275,N_9867,N_7666);
and UO_1276 (O_1276,N_8467,N_8371);
and UO_1277 (O_1277,N_6345,N_7314);
nor UO_1278 (O_1278,N_5844,N_6287);
nand UO_1279 (O_1279,N_6076,N_8757);
nor UO_1280 (O_1280,N_6872,N_8535);
or UO_1281 (O_1281,N_9295,N_9627);
and UO_1282 (O_1282,N_8125,N_8309);
and UO_1283 (O_1283,N_5724,N_6151);
nand UO_1284 (O_1284,N_5544,N_9209);
or UO_1285 (O_1285,N_9277,N_9882);
and UO_1286 (O_1286,N_6538,N_5556);
or UO_1287 (O_1287,N_5242,N_6963);
nand UO_1288 (O_1288,N_7002,N_8916);
or UO_1289 (O_1289,N_9665,N_5025);
xnor UO_1290 (O_1290,N_7607,N_8854);
or UO_1291 (O_1291,N_9177,N_5472);
nor UO_1292 (O_1292,N_6106,N_7049);
or UO_1293 (O_1293,N_8193,N_5885);
and UO_1294 (O_1294,N_5838,N_6850);
nand UO_1295 (O_1295,N_9643,N_8189);
nor UO_1296 (O_1296,N_8283,N_6226);
or UO_1297 (O_1297,N_5618,N_5286);
and UO_1298 (O_1298,N_8928,N_9477);
or UO_1299 (O_1299,N_5173,N_9781);
or UO_1300 (O_1300,N_6730,N_8310);
nor UO_1301 (O_1301,N_5019,N_5811);
nand UO_1302 (O_1302,N_8110,N_9516);
nor UO_1303 (O_1303,N_5594,N_5920);
nor UO_1304 (O_1304,N_6871,N_9193);
xnor UO_1305 (O_1305,N_7919,N_6427);
nor UO_1306 (O_1306,N_8282,N_9382);
nor UO_1307 (O_1307,N_6491,N_9097);
or UO_1308 (O_1308,N_6479,N_8898);
nand UO_1309 (O_1309,N_9522,N_6169);
nand UO_1310 (O_1310,N_6362,N_9088);
and UO_1311 (O_1311,N_8838,N_5304);
nor UO_1312 (O_1312,N_6165,N_8357);
and UO_1313 (O_1313,N_9674,N_6608);
nand UO_1314 (O_1314,N_9419,N_5646);
and UO_1315 (O_1315,N_5637,N_9509);
nand UO_1316 (O_1316,N_7226,N_8667);
and UO_1317 (O_1317,N_7647,N_6388);
and UO_1318 (O_1318,N_9427,N_5559);
or UO_1319 (O_1319,N_6316,N_5184);
or UO_1320 (O_1320,N_7918,N_7250);
or UO_1321 (O_1321,N_5014,N_6694);
nor UO_1322 (O_1322,N_8971,N_6298);
nand UO_1323 (O_1323,N_5357,N_5670);
nor UO_1324 (O_1324,N_5246,N_9923);
nor UO_1325 (O_1325,N_7790,N_5046);
nor UO_1326 (O_1326,N_7561,N_6128);
or UO_1327 (O_1327,N_6781,N_5106);
nor UO_1328 (O_1328,N_5200,N_8609);
nand UO_1329 (O_1329,N_8031,N_7786);
or UO_1330 (O_1330,N_7384,N_6074);
or UO_1331 (O_1331,N_9655,N_9632);
and UO_1332 (O_1332,N_6245,N_9429);
and UO_1333 (O_1333,N_6777,N_9361);
or UO_1334 (O_1334,N_9772,N_7614);
or UO_1335 (O_1335,N_5437,N_6083);
and UO_1336 (O_1336,N_8687,N_8321);
nand UO_1337 (O_1337,N_6238,N_9899);
or UO_1338 (O_1338,N_8978,N_6899);
nor UO_1339 (O_1339,N_8868,N_7421);
and UO_1340 (O_1340,N_6624,N_5554);
and UO_1341 (O_1341,N_7337,N_8427);
or UO_1342 (O_1342,N_6349,N_7288);
nor UO_1343 (O_1343,N_6489,N_6591);
and UO_1344 (O_1344,N_5859,N_5506);
nor UO_1345 (O_1345,N_8455,N_7566);
nor UO_1346 (O_1346,N_7321,N_7395);
or UO_1347 (O_1347,N_9573,N_6451);
xnor UO_1348 (O_1348,N_7715,N_9624);
or UO_1349 (O_1349,N_6822,N_7862);
nor UO_1350 (O_1350,N_7158,N_7044);
or UO_1351 (O_1351,N_9608,N_5558);
nor UO_1352 (O_1352,N_9618,N_7851);
nand UO_1353 (O_1353,N_7748,N_8803);
and UO_1354 (O_1354,N_8950,N_5905);
or UO_1355 (O_1355,N_9460,N_6209);
xor UO_1356 (O_1356,N_5136,N_5808);
and UO_1357 (O_1357,N_5067,N_6537);
and UO_1358 (O_1358,N_6170,N_9589);
and UO_1359 (O_1359,N_6448,N_7683);
or UO_1360 (O_1360,N_9118,N_5314);
and UO_1361 (O_1361,N_9178,N_6684);
nor UO_1362 (O_1362,N_6267,N_5505);
or UO_1363 (O_1363,N_8927,N_9107);
or UO_1364 (O_1364,N_8625,N_7571);
xnor UO_1365 (O_1365,N_7331,N_9190);
or UO_1366 (O_1366,N_6131,N_8939);
nor UO_1367 (O_1367,N_6029,N_9223);
and UO_1368 (O_1368,N_5118,N_9759);
or UO_1369 (O_1369,N_8327,N_7692);
or UO_1370 (O_1370,N_6798,N_6326);
or UO_1371 (O_1371,N_7516,N_7076);
nand UO_1372 (O_1372,N_9794,N_5421);
nand UO_1373 (O_1373,N_5855,N_5573);
nor UO_1374 (O_1374,N_6764,N_9318);
nor UO_1375 (O_1375,N_7532,N_9523);
nor UO_1376 (O_1376,N_6909,N_6554);
nor UO_1377 (O_1377,N_7278,N_8190);
or UO_1378 (O_1378,N_8159,N_7847);
nand UO_1379 (O_1379,N_8936,N_8388);
nand UO_1380 (O_1380,N_7869,N_5779);
or UO_1381 (O_1381,N_7629,N_7215);
and UO_1382 (O_1382,N_5804,N_8577);
and UO_1383 (O_1383,N_6550,N_5690);
or UO_1384 (O_1384,N_8652,N_6036);
or UO_1385 (O_1385,N_6602,N_6210);
nor UO_1386 (O_1386,N_6558,N_8856);
and UO_1387 (O_1387,N_6700,N_5856);
and UO_1388 (O_1388,N_8493,N_6374);
xor UO_1389 (O_1389,N_5140,N_6073);
and UO_1390 (O_1390,N_5207,N_5515);
nor UO_1391 (O_1391,N_9514,N_8167);
nor UO_1392 (O_1392,N_5055,N_5125);
nor UO_1393 (O_1393,N_5348,N_8156);
or UO_1394 (O_1394,N_9919,N_5549);
and UO_1395 (O_1395,N_6286,N_9754);
or UO_1396 (O_1396,N_5672,N_8855);
nor UO_1397 (O_1397,N_9261,N_7768);
nand UO_1398 (O_1398,N_7231,N_7941);
or UO_1399 (O_1399,N_9601,N_9192);
and UO_1400 (O_1400,N_9154,N_7121);
and UO_1401 (O_1401,N_8695,N_5293);
xnor UO_1402 (O_1402,N_7078,N_6475);
or UO_1403 (O_1403,N_8440,N_8999);
or UO_1404 (O_1404,N_7006,N_6203);
nor UO_1405 (O_1405,N_5062,N_7898);
and UO_1406 (O_1406,N_7767,N_6945);
nor UO_1407 (O_1407,N_9412,N_8727);
nor UO_1408 (O_1408,N_6533,N_6002);
and UO_1409 (O_1409,N_7797,N_8490);
and UO_1410 (O_1410,N_7361,N_8651);
and UO_1411 (O_1411,N_6542,N_6453);
and UO_1412 (O_1412,N_9369,N_7564);
nand UO_1413 (O_1413,N_9906,N_8452);
and UO_1414 (O_1414,N_5466,N_6809);
or UO_1415 (O_1415,N_7219,N_6667);
nor UO_1416 (O_1416,N_5198,N_8183);
and UO_1417 (O_1417,N_5735,N_5112);
nand UO_1418 (O_1418,N_8681,N_5996);
xnor UO_1419 (O_1419,N_8969,N_6381);
nand UO_1420 (O_1420,N_9945,N_6990);
xnor UO_1421 (O_1421,N_5641,N_5545);
nand UO_1422 (O_1422,N_8558,N_9988);
and UO_1423 (O_1423,N_6395,N_6956);
or UO_1424 (O_1424,N_5624,N_5600);
nor UO_1425 (O_1425,N_5581,N_5379);
xnor UO_1426 (O_1426,N_8697,N_9130);
nand UO_1427 (O_1427,N_7804,N_6257);
nor UO_1428 (O_1428,N_9510,N_6727);
or UO_1429 (O_1429,N_5252,N_7832);
and UO_1430 (O_1430,N_5123,N_9881);
nand UO_1431 (O_1431,N_9197,N_8863);
and UO_1432 (O_1432,N_5874,N_7562);
or UO_1433 (O_1433,N_9940,N_9688);
or UO_1434 (O_1434,N_6341,N_7392);
nand UO_1435 (O_1435,N_7511,N_8762);
and UO_1436 (O_1436,N_6883,N_6300);
nor UO_1437 (O_1437,N_6023,N_5400);
nor UO_1438 (O_1438,N_9503,N_9465);
or UO_1439 (O_1439,N_5691,N_6520);
and UO_1440 (O_1440,N_6037,N_8389);
nand UO_1441 (O_1441,N_5094,N_5395);
nand UO_1442 (O_1442,N_7527,N_9030);
or UO_1443 (O_1443,N_7880,N_9194);
nor UO_1444 (O_1444,N_6372,N_5051);
nand UO_1445 (O_1445,N_6570,N_5231);
or UO_1446 (O_1446,N_6583,N_8849);
and UO_1447 (O_1447,N_9593,N_6923);
xor UO_1448 (O_1448,N_6251,N_8002);
or UO_1449 (O_1449,N_9348,N_6742);
nand UO_1450 (O_1450,N_9507,N_5683);
and UO_1451 (O_1451,N_8291,N_6105);
nor UO_1452 (O_1452,N_9685,N_8315);
and UO_1453 (O_1453,N_6584,N_6382);
xor UO_1454 (O_1454,N_9791,N_6327);
xor UO_1455 (O_1455,N_5943,N_7730);
or UO_1456 (O_1456,N_6342,N_8034);
nor UO_1457 (O_1457,N_9248,N_8453);
nand UO_1458 (O_1458,N_8100,N_6713);
or UO_1459 (O_1459,N_5608,N_6080);
and UO_1460 (O_1460,N_7468,N_6200);
or UO_1461 (O_1461,N_5222,N_5992);
and UO_1462 (O_1462,N_6755,N_9111);
nor UO_1463 (O_1463,N_6393,N_8798);
nand UO_1464 (O_1464,N_7247,N_8384);
nand UO_1465 (O_1465,N_9621,N_9228);
xor UO_1466 (O_1466,N_7148,N_7550);
and UO_1467 (O_1467,N_5256,N_7774);
nand UO_1468 (O_1468,N_5127,N_8415);
or UO_1469 (O_1469,N_5699,N_7088);
xor UO_1470 (O_1470,N_5354,N_5634);
or UO_1471 (O_1471,N_7485,N_5561);
nand UO_1472 (O_1472,N_6459,N_9113);
or UO_1473 (O_1473,N_5454,N_5187);
or UO_1474 (O_1474,N_9368,N_7344);
nand UO_1475 (O_1475,N_7581,N_8311);
nor UO_1476 (O_1476,N_7254,N_7494);
and UO_1477 (O_1477,N_9787,N_9657);
and UO_1478 (O_1478,N_9905,N_7696);
and UO_1479 (O_1479,N_6098,N_9392);
xnor UO_1480 (O_1480,N_5152,N_6814);
and UO_1481 (O_1481,N_8076,N_6432);
xnor UO_1482 (O_1482,N_7747,N_7151);
and UO_1483 (O_1483,N_7417,N_9241);
or UO_1484 (O_1484,N_6471,N_5070);
nand UO_1485 (O_1485,N_8018,N_8645);
or UO_1486 (O_1486,N_6513,N_8679);
and UO_1487 (O_1487,N_7021,N_8314);
and UO_1488 (O_1488,N_9865,N_8050);
and UO_1489 (O_1489,N_8988,N_5430);
xnor UO_1490 (O_1490,N_5476,N_6219);
nand UO_1491 (O_1491,N_8025,N_8732);
or UO_1492 (O_1492,N_7831,N_6419);
nand UO_1493 (O_1493,N_7416,N_8367);
and UO_1494 (O_1494,N_5816,N_5132);
or UO_1495 (O_1495,N_6215,N_8124);
nor UO_1496 (O_1496,N_6087,N_5799);
nor UO_1497 (O_1497,N_7655,N_9963);
nand UO_1498 (O_1498,N_7439,N_9504);
nor UO_1499 (O_1499,N_6504,N_5332);
endmodule