module basic_1500_15000_2000_60_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_1045,In_1307);
xor U1 (N_1,In_658,In_536);
and U2 (N_2,In_571,In_674);
and U3 (N_3,In_653,In_1497);
or U4 (N_4,In_1492,In_1140);
and U5 (N_5,In_226,In_1336);
nor U6 (N_6,In_169,In_1299);
or U7 (N_7,In_1192,In_187);
nor U8 (N_8,In_1365,In_796);
nor U9 (N_9,In_1031,In_834);
or U10 (N_10,In_515,In_1340);
nand U11 (N_11,In_681,In_716);
nand U12 (N_12,In_1369,In_998);
nor U13 (N_13,In_512,In_1062);
and U14 (N_14,In_670,In_1129);
xor U15 (N_15,In_1003,In_853);
nand U16 (N_16,In_167,In_1450);
nand U17 (N_17,In_1073,In_983);
or U18 (N_18,In_559,In_560);
or U19 (N_19,In_881,In_1154);
xnor U20 (N_20,In_67,In_908);
or U21 (N_21,In_686,In_1110);
and U22 (N_22,In_1412,In_683);
xnor U23 (N_23,In_1390,In_1020);
nor U24 (N_24,In_427,In_337);
and U25 (N_25,In_1309,In_832);
and U26 (N_26,In_583,In_1370);
nand U27 (N_27,In_112,In_646);
nor U28 (N_28,In_966,In_673);
nand U29 (N_29,In_434,In_847);
or U30 (N_30,In_550,In_1130);
or U31 (N_31,In_1253,In_609);
nand U32 (N_32,In_51,In_772);
nand U33 (N_33,In_189,In_878);
and U34 (N_34,In_861,In_305);
nor U35 (N_35,In_1418,In_655);
xor U36 (N_36,In_216,In_184);
xnor U37 (N_37,In_1105,In_720);
nor U38 (N_38,In_761,In_730);
xnor U39 (N_39,In_445,In_736);
nand U40 (N_40,In_126,In_1178);
and U41 (N_41,In_1074,In_895);
nand U42 (N_42,In_397,In_221);
and U43 (N_43,In_188,In_32);
nor U44 (N_44,In_709,In_178);
nand U45 (N_45,In_977,In_432);
and U46 (N_46,In_152,In_933);
or U47 (N_47,In_680,In_1421);
or U48 (N_48,In_902,In_920);
nand U49 (N_49,In_464,In_639);
and U50 (N_50,In_1126,In_575);
or U51 (N_51,In_1375,In_972);
and U52 (N_52,In_1368,In_1173);
or U53 (N_53,In_992,In_484);
nand U54 (N_54,In_119,In_2);
and U55 (N_55,In_153,In_462);
or U56 (N_56,In_558,In_1422);
and U57 (N_57,In_260,In_669);
xnor U58 (N_58,In_961,In_668);
or U59 (N_59,In_628,In_1437);
nand U60 (N_60,In_986,In_504);
xor U61 (N_61,In_369,In_461);
and U62 (N_62,In_648,In_726);
nand U63 (N_63,In_1429,In_848);
nand U64 (N_64,In_243,In_1224);
nor U65 (N_65,In_1040,In_1168);
nand U66 (N_66,In_146,In_752);
or U67 (N_67,In_223,In_723);
xnor U68 (N_68,In_236,In_1187);
xnor U69 (N_69,In_980,In_812);
or U70 (N_70,In_879,In_778);
nand U71 (N_71,In_917,In_1015);
and U72 (N_72,In_302,In_1352);
xnor U73 (N_73,In_725,In_603);
nor U74 (N_74,In_962,In_54);
and U75 (N_75,In_165,In_754);
and U76 (N_76,In_727,In_1278);
or U77 (N_77,In_508,In_921);
and U78 (N_78,In_1066,In_1282);
nand U79 (N_79,In_311,In_1294);
and U80 (N_80,In_963,In_134);
nand U81 (N_81,In_222,In_995);
xnor U82 (N_82,In_25,In_940);
nand U83 (N_83,In_261,In_210);
xor U84 (N_84,In_1327,In_1259);
and U85 (N_85,In_106,In_617);
xnor U86 (N_86,In_964,In_328);
xnor U87 (N_87,In_836,In_802);
xnor U88 (N_88,In_783,In_85);
xor U89 (N_89,In_935,In_565);
or U90 (N_90,In_627,In_593);
xor U91 (N_91,In_1402,In_1213);
or U92 (N_92,In_396,In_419);
or U93 (N_93,In_450,In_1247);
nor U94 (N_94,In_1498,In_1306);
and U95 (N_95,In_1443,In_949);
and U96 (N_96,In_1258,In_551);
xor U97 (N_97,In_356,In_359);
or U98 (N_98,In_459,In_74);
xnor U99 (N_99,In_372,In_102);
or U100 (N_100,In_68,In_477);
or U101 (N_101,In_4,In_734);
nand U102 (N_102,In_1001,In_1332);
or U103 (N_103,In_1433,In_466);
nand U104 (N_104,In_637,In_497);
or U105 (N_105,In_804,In_290);
nor U106 (N_106,In_1069,In_109);
xor U107 (N_107,In_854,In_561);
or U108 (N_108,In_1133,In_1287);
xnor U109 (N_109,In_330,In_1029);
nor U110 (N_110,In_181,In_1403);
nand U111 (N_111,In_1022,In_1397);
nand U112 (N_112,In_267,In_1139);
xnor U113 (N_113,In_448,In_914);
nor U114 (N_114,In_621,In_326);
and U115 (N_115,In_244,In_1083);
nand U116 (N_116,In_624,In_1354);
xnor U117 (N_117,In_1274,In_846);
and U118 (N_118,In_1209,In_491);
nor U119 (N_119,In_810,In_288);
xor U120 (N_120,In_1423,In_1010);
nor U121 (N_121,In_403,In_241);
nand U122 (N_122,In_1084,In_1158);
and U123 (N_123,In_1042,In_387);
nand U124 (N_124,In_546,In_443);
and U125 (N_125,In_5,In_517);
and U126 (N_126,In_422,In_1101);
or U127 (N_127,In_912,In_13);
xor U128 (N_128,In_896,In_1373);
or U129 (N_129,In_227,In_488);
nand U130 (N_130,In_95,In_629);
or U131 (N_131,In_873,In_163);
and U132 (N_132,In_755,In_430);
nand U133 (N_133,In_785,In_46);
and U134 (N_134,In_883,In_80);
nor U135 (N_135,In_346,In_1115);
nor U136 (N_136,In_1326,In_538);
nor U137 (N_137,In_361,In_811);
xor U138 (N_138,In_179,In_1440);
xor U139 (N_139,In_1358,In_943);
or U140 (N_140,In_421,In_1302);
xor U141 (N_141,In_1479,In_235);
and U142 (N_142,In_1261,In_132);
nand U143 (N_143,In_1220,In_332);
nand U144 (N_144,In_160,In_280);
and U145 (N_145,In_1273,In_925);
xnor U146 (N_146,In_1350,In_121);
and U147 (N_147,In_981,In_656);
xnor U148 (N_148,In_1449,In_254);
xnor U149 (N_149,In_148,In_1068);
nor U150 (N_150,In_1235,In_566);
and U151 (N_151,In_945,In_1219);
and U152 (N_152,In_388,In_350);
xor U153 (N_153,In_510,In_1036);
nand U154 (N_154,In_1,In_1266);
nand U155 (N_155,In_1198,In_97);
or U156 (N_156,In_620,In_1246);
nand U157 (N_157,In_718,In_447);
xor U158 (N_158,In_867,In_742);
xor U159 (N_159,In_1314,In_602);
xor U160 (N_160,In_82,In_301);
or U161 (N_161,In_947,In_1098);
and U162 (N_162,In_65,In_706);
nand U163 (N_163,In_1455,In_1233);
and U164 (N_164,In_283,In_1148);
or U165 (N_165,In_1468,In_395);
and U166 (N_166,In_835,In_1216);
and U167 (N_167,In_1017,In_199);
xor U168 (N_168,In_207,In_56);
xnor U169 (N_169,In_692,In_663);
or U170 (N_170,In_699,In_996);
or U171 (N_171,In_92,In_939);
xnor U172 (N_172,In_1499,In_118);
or U173 (N_173,In_341,In_161);
xnor U174 (N_174,In_1271,In_292);
and U175 (N_175,In_798,In_822);
or U176 (N_176,In_768,In_1431);
nor U177 (N_177,In_310,In_764);
or U178 (N_178,In_379,In_580);
or U179 (N_179,In_500,In_1156);
and U180 (N_180,In_313,In_1337);
nand U181 (N_181,In_779,In_606);
or U182 (N_182,In_463,In_1063);
or U183 (N_183,In_1002,In_1035);
nor U184 (N_184,In_1109,In_1049);
or U185 (N_185,In_1471,In_431);
or U186 (N_186,In_277,In_38);
nand U187 (N_187,In_1495,In_868);
or U188 (N_188,In_414,In_58);
nand U189 (N_189,In_322,In_759);
or U190 (N_190,In_619,In_122);
xnor U191 (N_191,In_127,In_149);
or U192 (N_192,In_271,In_1131);
xor U193 (N_193,In_631,In_1033);
and U194 (N_194,In_885,In_1195);
or U195 (N_195,In_1215,In_1023);
or U196 (N_196,In_308,In_824);
xor U197 (N_197,In_480,In_1467);
nor U198 (N_198,In_735,In_470);
nand U199 (N_199,In_731,In_1362);
or U200 (N_200,In_857,In_492);
xnor U201 (N_201,In_479,In_76);
or U202 (N_202,In_159,In_978);
or U203 (N_203,In_625,In_863);
or U204 (N_204,In_1071,In_423);
nor U205 (N_205,In_893,In_245);
and U206 (N_206,In_927,In_139);
and U207 (N_207,In_1312,In_1413);
nor U208 (N_208,In_1276,In_1102);
nand U209 (N_209,In_1268,In_608);
or U210 (N_210,In_1311,In_1018);
xor U211 (N_211,In_887,In_398);
nand U212 (N_212,In_553,In_540);
or U213 (N_213,In_931,In_647);
xnor U214 (N_214,In_378,In_532);
xnor U215 (N_215,In_1136,In_386);
and U216 (N_216,In_1396,In_1447);
and U217 (N_217,In_1118,In_390);
nor U218 (N_218,In_1292,In_840);
nor U219 (N_219,In_460,In_710);
xnor U220 (N_220,In_700,In_79);
nor U221 (N_221,In_150,In_708);
nor U222 (N_222,In_592,In_733);
nand U223 (N_223,In_909,In_702);
nor U224 (N_224,In_1037,In_123);
and U225 (N_225,In_1197,In_130);
or U226 (N_226,In_894,In_472);
and U227 (N_227,In_1088,In_852);
and U228 (N_228,In_220,In_1225);
or U229 (N_229,In_1211,In_1272);
nand U230 (N_230,In_1163,In_1123);
xor U231 (N_231,In_829,In_166);
nand U232 (N_232,In_93,In_89);
xnor U233 (N_233,In_1316,In_974);
and U234 (N_234,In_1174,In_452);
nor U235 (N_235,In_630,In_86);
and U236 (N_236,In_475,In_103);
or U237 (N_237,In_780,In_594);
and U238 (N_238,In_1053,In_1108);
or U239 (N_239,In_850,In_324);
nand U240 (N_240,In_1059,In_108);
xnor U241 (N_241,In_1021,In_664);
or U242 (N_242,In_1103,In_749);
nor U243 (N_243,In_192,In_340);
or U244 (N_244,In_1189,In_882);
nor U245 (N_245,In_272,In_530);
xnor U246 (N_246,In_1466,In_458);
nor U247 (N_247,In_316,In_1322);
or U248 (N_248,In_1205,In_24);
or U249 (N_249,In_688,In_531);
nor U250 (N_250,N_105,In_839);
nor U251 (N_251,In_751,In_273);
nand U252 (N_252,In_1411,In_349);
or U253 (N_253,In_249,In_1406);
nor U254 (N_254,In_418,N_5);
xnor U255 (N_255,In_384,In_1161);
xnor U256 (N_256,In_293,In_440);
nor U257 (N_257,In_923,N_106);
or U258 (N_258,In_219,In_794);
and U259 (N_259,In_217,In_872);
xor U260 (N_260,In_1484,In_634);
xnor U261 (N_261,In_537,In_513);
nor U262 (N_262,In_1043,N_39);
xnor U263 (N_263,In_255,In_1222);
xor U264 (N_264,In_1313,N_141);
nor U265 (N_265,In_793,In_131);
nor U266 (N_266,In_1207,In_672);
or U267 (N_267,In_952,In_856);
and U268 (N_268,In_469,N_151);
nand U269 (N_269,In_1416,In_493);
and U270 (N_270,N_80,In_564);
or U271 (N_271,In_1398,In_490);
and U272 (N_272,In_202,In_521);
nand U273 (N_273,N_130,In_898);
xor U274 (N_274,N_241,In_111);
nor U275 (N_275,N_53,In_1414);
or U276 (N_276,In_474,In_684);
xnor U277 (N_277,In_377,In_1104);
nand U278 (N_278,In_1204,In_170);
nand U279 (N_279,In_717,In_544);
nor U280 (N_280,In_1289,In_1277);
xnor U281 (N_281,In_238,In_555);
nor U282 (N_282,In_632,N_32);
nor U283 (N_283,In_1330,N_173);
or U284 (N_284,In_285,In_1107);
or U285 (N_285,In_693,In_194);
xnor U286 (N_286,In_1394,In_997);
and U287 (N_287,In_87,In_1335);
nand U288 (N_288,In_1128,In_1463);
nor U289 (N_289,In_214,In_666);
nand U290 (N_290,N_209,In_1376);
and U291 (N_291,N_204,N_116);
xnor U292 (N_292,In_107,In_34);
nand U293 (N_293,N_232,In_234);
nand U294 (N_294,In_204,In_66);
nor U295 (N_295,In_904,In_158);
and U296 (N_296,In_270,N_215);
or U297 (N_297,In_366,In_1093);
nand U298 (N_298,In_274,In_1342);
nor U299 (N_299,In_406,In_1080);
and U300 (N_300,In_411,In_282);
and U301 (N_301,In_91,In_233);
nor U302 (N_302,In_884,In_1328);
and U303 (N_303,In_1087,N_175);
nor U304 (N_304,In_1363,N_56);
xnor U305 (N_305,In_968,N_206);
nand U306 (N_306,N_244,In_610);
nor U307 (N_307,In_1435,In_1349);
xnor U308 (N_308,In_1480,In_1119);
or U309 (N_309,In_27,In_748);
nor U310 (N_310,In_101,N_94);
or U311 (N_311,In_180,In_1125);
and U312 (N_312,In_1190,N_192);
nor U313 (N_313,N_55,In_781);
nor U314 (N_314,In_1157,In_1208);
and U315 (N_315,In_1478,In_251);
nor U316 (N_316,In_690,N_207);
nor U317 (N_317,In_859,In_548);
nand U318 (N_318,N_82,In_352);
and U319 (N_319,In_1228,In_975);
and U320 (N_320,In_394,In_1099);
or U321 (N_321,In_622,In_1252);
and U322 (N_322,In_110,In_671);
nand U323 (N_323,N_140,In_816);
or U324 (N_324,In_1283,In_821);
or U325 (N_325,N_134,In_1286);
or U326 (N_326,In_1120,In_286);
and U327 (N_327,In_1210,In_104);
nand U328 (N_328,In_612,In_843);
and U329 (N_329,N_179,In_1072);
nor U330 (N_330,In_1318,In_645);
xor U331 (N_331,In_1399,In_412);
xor U332 (N_332,In_616,In_505);
nor U333 (N_333,In_1308,In_105);
nor U334 (N_334,N_34,N_20);
and U335 (N_335,In_971,N_104);
nand U336 (N_336,In_1485,In_516);
or U337 (N_337,In_215,N_228);
xnor U338 (N_338,In_374,In_1193);
nor U339 (N_339,In_1470,N_200);
nand U340 (N_340,In_888,In_642);
nor U341 (N_341,In_711,In_263);
xor U342 (N_342,In_957,N_211);
nand U343 (N_343,In_1381,In_239);
and U344 (N_344,In_495,N_59);
xor U345 (N_345,In_831,In_1025);
or U346 (N_346,N_15,In_232);
xor U347 (N_347,In_154,In_665);
and U348 (N_348,In_237,In_1171);
or U349 (N_349,In_30,In_573);
nand U350 (N_350,In_42,In_314);
xor U351 (N_351,N_248,N_147);
and U352 (N_352,In_597,In_1013);
nand U353 (N_353,In_1295,In_14);
xnor U354 (N_354,N_139,In_362);
xor U355 (N_355,In_318,In_231);
nor U356 (N_356,In_409,In_415);
nand U357 (N_357,In_333,In_529);
nor U358 (N_358,In_1428,In_381);
or U359 (N_359,In_18,In_1092);
xnor U360 (N_360,N_218,In_502);
nor U361 (N_361,In_6,N_152);
nand U362 (N_362,In_578,In_1444);
nor U363 (N_363,N_237,N_148);
or U364 (N_364,In_509,In_654);
nor U365 (N_365,In_115,In_1434);
and U366 (N_366,In_864,In_813);
nor U367 (N_367,In_958,In_814);
nand U368 (N_368,In_1196,In_696);
xor U369 (N_369,In_763,In_762);
or U370 (N_370,In_449,In_1378);
nand U371 (N_371,In_203,In_1483);
and U372 (N_372,In_1027,In_1245);
and U373 (N_373,N_89,In_874);
nor U374 (N_374,In_1079,N_238);
nand U375 (N_375,In_23,N_26);
nor U376 (N_376,In_1305,In_444);
or U377 (N_377,In_549,In_1032);
xnor U378 (N_378,In_331,In_468);
nor U379 (N_379,In_789,N_67);
and U380 (N_380,In_801,In_1395);
nand U381 (N_381,N_122,In_402);
nor U382 (N_382,In_1388,N_62);
and U383 (N_383,In_809,In_941);
nor U384 (N_384,In_1095,N_114);
or U385 (N_385,In_1386,In_1430);
xnor U386 (N_386,N_75,In_62);
nor U387 (N_387,In_1425,In_1293);
xnor U388 (N_388,In_830,In_607);
and U389 (N_389,In_1475,In_1357);
nor U390 (N_390,In_496,In_31);
or U391 (N_391,In_899,N_191);
and U392 (N_392,In_584,In_704);
or U393 (N_393,In_499,In_162);
nand U394 (N_394,In_77,In_511);
nor U395 (N_395,In_689,N_117);
nand U396 (N_396,In_55,In_334);
nor U397 (N_397,In_776,In_737);
nor U398 (N_398,In_416,N_71);
nor U399 (N_399,N_47,N_81);
or U400 (N_400,In_435,In_201);
nor U401 (N_401,In_1076,N_90);
nor U402 (N_402,In_28,N_85);
and U403 (N_403,In_309,In_436);
nor U404 (N_404,In_640,In_745);
nand U405 (N_405,In_53,N_186);
or U406 (N_406,N_61,N_203);
nand U407 (N_407,In_928,In_1009);
nor U408 (N_408,In_527,In_960);
or U409 (N_409,In_442,In_1251);
or U410 (N_410,In_456,In_1400);
xnor U411 (N_411,In_451,In_1367);
xnor U412 (N_412,N_18,In_638);
nand U413 (N_413,In_269,N_109);
xor U414 (N_414,N_108,N_28);
xnor U415 (N_415,In_965,In_1124);
nand U416 (N_416,In_862,In_389);
nor U417 (N_417,In_1325,In_858);
or U418 (N_418,N_180,In_787);
xor U419 (N_419,In_1364,In_224);
nor U420 (N_420,In_345,In_155);
xnor U421 (N_421,In_147,In_740);
and U422 (N_422,In_1151,N_205);
or U423 (N_423,In_1232,In_1476);
and U424 (N_424,In_1182,In_1355);
nand U425 (N_425,In_335,In_347);
and U426 (N_426,In_1201,In_252);
nor U427 (N_427,In_1382,In_52);
nor U428 (N_428,In_315,In_317);
xor U429 (N_429,N_36,In_876);
and U430 (N_430,In_946,In_542);
nor U431 (N_431,In_1097,In_1481);
and U432 (N_432,In_1046,In_919);
nand U433 (N_433,In_247,In_1446);
nor U434 (N_434,In_803,In_1324);
xor U435 (N_435,N_95,In_1380);
or U436 (N_436,In_401,In_886);
and U437 (N_437,In_1490,In_765);
nor U438 (N_438,In_405,In_124);
nand U439 (N_439,In_1242,N_14);
xor U440 (N_440,N_70,In_1114);
nor U441 (N_441,In_63,In_339);
nand U442 (N_442,In_643,N_166);
and U443 (N_443,In_891,In_633);
or U444 (N_444,In_1417,In_694);
xor U445 (N_445,In_498,In_1138);
nor U446 (N_446,In_1451,In_1441);
nand U447 (N_447,In_1177,In_39);
xor U448 (N_448,In_1345,In_545);
xnor U449 (N_449,In_41,N_99);
nand U450 (N_450,In_1344,In_1038);
and U451 (N_451,N_226,N_160);
or U452 (N_452,N_96,N_169);
and U453 (N_453,In_636,In_1269);
nor U454 (N_454,In_1214,In_136);
and U455 (N_455,N_66,In_1061);
or U456 (N_456,In_905,In_1472);
nor U457 (N_457,In_1482,In_1353);
or U458 (N_458,In_1144,In_855);
nand U459 (N_459,In_44,N_154);
xnor U460 (N_460,N_38,In_924);
xor U461 (N_461,In_790,In_1048);
or U462 (N_462,In_1134,N_31);
or U463 (N_463,In_382,N_236);
nor U464 (N_464,In_1385,In_144);
or U465 (N_465,In_753,In_1212);
nor U466 (N_466,In_1067,In_370);
xnor U467 (N_467,N_74,N_164);
nor U468 (N_468,N_35,In_64);
nor U469 (N_469,In_129,N_143);
or U470 (N_470,In_808,In_782);
or U471 (N_471,In_767,In_870);
and U472 (N_472,In_662,N_194);
or U473 (N_473,N_142,In_156);
and U474 (N_474,N_128,N_231);
and U475 (N_475,In_732,In_937);
nor U476 (N_476,In_534,In_1077);
xnor U477 (N_477,In_1052,In_951);
nand U478 (N_478,In_441,In_133);
nand U479 (N_479,In_926,N_42);
xnor U480 (N_480,In_907,In_959);
nand U481 (N_481,N_92,In_209);
or U482 (N_482,In_969,In_626);
nand U483 (N_483,In_1487,In_256);
or U484 (N_484,N_60,In_543);
nand U485 (N_485,In_266,In_1113);
nor U486 (N_486,In_47,In_1166);
nand U487 (N_487,N_16,N_23);
and U488 (N_488,In_1329,N_46);
or U489 (N_489,In_729,In_426);
or U490 (N_490,In_797,N_219);
xor U491 (N_491,In_1094,In_1223);
nor U492 (N_492,In_182,N_17);
or U493 (N_493,In_1089,In_1256);
nor U494 (N_494,In_503,In_999);
or U495 (N_495,In_1203,In_900);
nand U496 (N_496,In_33,In_1300);
and U497 (N_497,N_223,N_233);
nand U498 (N_498,In_1202,In_113);
or U499 (N_499,In_930,In_114);
nand U500 (N_500,N_217,In_817);
nand U501 (N_501,In_211,In_1270);
and U502 (N_502,In_218,In_84);
nand U503 (N_503,N_454,N_407);
nand U504 (N_504,In_596,In_598);
or U505 (N_505,N_83,In_72);
and U506 (N_506,In_1255,In_677);
xor U507 (N_507,N_414,In_0);
nand U508 (N_508,N_301,In_922);
nor U509 (N_509,In_618,In_875);
nor U510 (N_510,N_159,In_1415);
and U511 (N_511,In_576,In_183);
or U512 (N_512,In_81,In_1284);
and U513 (N_513,In_83,N_37);
xnor U514 (N_514,N_267,N_181);
nand U515 (N_515,In_1112,N_457);
xor U516 (N_516,N_275,In_1457);
xnor U517 (N_517,N_328,N_258);
xnor U518 (N_518,In_1194,In_1383);
or U519 (N_519,N_297,In_659);
or U520 (N_520,N_224,N_201);
xor U521 (N_521,N_277,N_363);
and U522 (N_522,N_392,In_392);
and U523 (N_523,N_292,In_1047);
xnor U524 (N_524,In_721,N_421);
nor U525 (N_525,N_335,In_932);
and U526 (N_526,N_121,N_489);
or U527 (N_527,In_438,In_319);
or U528 (N_528,N_426,In_1405);
xnor U529 (N_529,N_375,N_284);
nor U530 (N_530,In_248,N_458);
and U531 (N_531,In_1149,In_719);
and U532 (N_532,In_1008,N_372);
and U533 (N_533,N_468,In_75);
xor U534 (N_534,N_54,In_19);
xor U535 (N_535,N_350,N_86);
and U536 (N_536,N_494,In_1169);
or U537 (N_537,In_455,In_523);
and U538 (N_538,N_401,In_481);
nor U539 (N_539,In_407,In_1279);
nand U540 (N_540,N_385,N_429);
nand U541 (N_541,N_486,In_644);
xor U542 (N_542,N_93,In_116);
xnor U543 (N_543,N_354,In_775);
and U544 (N_544,N_460,N_126);
xnor U545 (N_545,N_161,N_176);
nand U546 (N_546,N_131,N_91);
nor U547 (N_547,In_206,N_252);
nand U548 (N_548,N_187,N_321);
and U549 (N_549,In_554,N_381);
or U550 (N_550,In_1408,In_649);
xor U551 (N_551,In_652,N_153);
or U552 (N_552,In_871,In_1339);
xor U553 (N_553,In_1410,In_667);
and U554 (N_554,In_1267,N_311);
xnor U555 (N_555,N_303,In_198);
nand U556 (N_556,In_259,In_845);
xnor U557 (N_557,In_228,In_911);
and U558 (N_558,In_57,In_1488);
xor U559 (N_559,In_1234,N_296);
nand U560 (N_560,N_485,N_52);
nor U561 (N_561,In_1351,In_577);
and U562 (N_562,In_383,N_402);
or U563 (N_563,In_143,N_113);
and U564 (N_564,N_2,N_21);
or U565 (N_565,In_1041,In_471);
nand U566 (N_566,In_229,N_387);
nor U567 (N_567,In_242,N_355);
xor U568 (N_568,In_525,In_1121);
xnor U569 (N_569,In_1419,In_777);
nand U570 (N_570,N_488,In_1474);
or U571 (N_571,In_760,N_110);
and U572 (N_572,In_1333,In_1150);
nand U573 (N_573,In_623,In_357);
nand U574 (N_574,N_393,N_425);
and U575 (N_575,N_382,In_485);
nor U576 (N_576,In_714,In_71);
or U577 (N_577,N_172,In_1461);
and U578 (N_578,In_164,N_380);
or U579 (N_579,In_1391,In_743);
xnor U580 (N_580,In_1427,In_1265);
nor U581 (N_581,In_604,N_496);
or U582 (N_582,N_273,N_341);
or U583 (N_583,In_424,In_901);
and U584 (N_584,N_476,N_119);
xnor U585 (N_585,In_373,N_222);
nor U586 (N_586,N_327,In_329);
and U587 (N_587,N_449,In_1304);
or U588 (N_588,N_12,N_102);
nor U589 (N_589,In_1469,In_1051);
and U590 (N_590,In_520,In_993);
xnor U591 (N_591,In_94,N_293);
nand U592 (N_592,N_49,In_849);
or U593 (N_593,N_250,In_979);
nor U594 (N_594,In_120,In_800);
or U595 (N_595,In_1462,N_450);
nand U596 (N_596,In_1028,In_138);
nand U597 (N_597,In_994,N_45);
or U598 (N_598,In_90,N_115);
nor U599 (N_599,In_1496,N_491);
xnor U600 (N_600,In_174,In_1019);
and U601 (N_601,N_58,N_334);
nor U602 (N_602,In_413,In_581);
xnor U603 (N_603,N_279,N_325);
or U604 (N_604,N_445,N_394);
nor U605 (N_605,In_691,N_497);
nor U606 (N_606,In_1347,In_323);
or U607 (N_607,In_371,In_246);
nand U608 (N_608,In_11,In_1206);
nand U609 (N_609,N_492,In_99);
nand U610 (N_610,In_1226,In_1016);
nand U611 (N_611,In_1145,In_991);
nand U612 (N_612,In_1426,N_170);
nand U613 (N_613,In_1146,In_641);
or U614 (N_614,N_251,N_234);
or U615 (N_615,In_695,In_806);
nand U616 (N_616,In_157,In_866);
or U617 (N_617,In_1106,In_750);
nor U618 (N_618,N_475,In_1082);
or U619 (N_619,In_984,N_349);
nor U620 (N_620,In_567,N_274);
or U621 (N_621,In_205,N_9);
xnor U622 (N_622,N_400,N_373);
nor U623 (N_623,N_225,In_657);
nor U624 (N_624,In_599,In_844);
nand U625 (N_625,N_462,In_815);
or U626 (N_626,N_359,In_195);
nor U627 (N_627,N_220,N_403);
nand U628 (N_628,In_841,In_1452);
xnor U629 (N_629,N_287,In_1160);
nand U630 (N_630,N_269,In_375);
or U631 (N_631,In_1236,In_284);
or U632 (N_632,N_469,N_319);
and U633 (N_633,N_427,N_177);
xor U634 (N_634,N_408,In_906);
xnor U635 (N_635,In_50,N_132);
or U636 (N_636,N_27,In_1439);
nand U637 (N_637,N_345,N_315);
xnor U638 (N_638,In_944,In_385);
nand U639 (N_639,In_1264,In_1039);
or U640 (N_640,In_1135,N_322);
nor U641 (N_641,N_298,In_877);
or U642 (N_642,In_1165,N_73);
nand U643 (N_643,N_336,In_1346);
or U644 (N_644,N_165,In_1142);
xnor U645 (N_645,In_890,In_1243);
nor U646 (N_646,N_137,N_123);
xnor U647 (N_647,In_1379,In_828);
nand U648 (N_648,N_443,In_651);
nand U649 (N_649,N_316,N_331);
nand U650 (N_650,In_391,N_444);
or U651 (N_651,In_1116,N_434);
xor U652 (N_652,In_60,In_1360);
and U653 (N_653,In_1155,N_302);
nand U654 (N_654,In_348,N_410);
nand U655 (N_655,In_950,In_1230);
and U656 (N_656,N_391,In_1011);
or U657 (N_657,N_495,N_299);
xor U658 (N_658,N_356,In_1473);
nand U659 (N_659,In_225,In_1085);
or U660 (N_660,In_1409,N_470);
xnor U661 (N_661,In_805,In_1331);
and U662 (N_662,In_819,In_454);
nand U663 (N_663,In_1359,In_1070);
and U664 (N_664,In_482,N_371);
and U665 (N_665,N_419,N_259);
nor U666 (N_666,N_30,In_1275);
nor U667 (N_667,In_1241,In_78);
and U668 (N_668,In_1323,N_4);
or U669 (N_669,In_1006,In_738);
and U670 (N_670,N_196,In_196);
xor U671 (N_671,In_660,N_490);
and U672 (N_672,In_408,In_49);
and U673 (N_673,N_452,In_21);
or U674 (N_674,N_430,In_1239);
xor U675 (N_675,N_361,In_1064);
or U676 (N_676,In_368,In_514);
nand U677 (N_677,In_177,In_29);
nand U678 (N_678,In_1054,In_1221);
and U679 (N_679,N_111,In_268);
and U680 (N_680,N_227,In_1248);
nand U681 (N_681,N_308,In_1170);
xor U682 (N_682,In_1217,N_50);
xor U683 (N_683,In_1091,In_903);
xor U684 (N_684,In_1024,In_1338);
nand U685 (N_685,N_411,In_1404);
or U686 (N_686,In_1262,In_137);
or U687 (N_687,In_8,In_574);
nor U688 (N_688,N_210,In_942);
xor U689 (N_689,N_249,N_351);
xnor U690 (N_690,N_72,N_286);
nand U691 (N_691,In_483,N_309);
nand U692 (N_692,In_851,In_417);
xor U693 (N_693,In_701,N_79);
or U694 (N_694,In_1387,In_1438);
or U695 (N_695,In_48,In_298);
or U696 (N_696,N_57,In_685);
nand U697 (N_697,N_455,In_36);
nand U698 (N_698,In_823,N_171);
or U699 (N_699,In_519,In_172);
nand U700 (N_700,In_1056,N_283);
nand U701 (N_701,In_586,In_45);
xor U702 (N_702,In_1057,In_1458);
nor U703 (N_703,In_552,N_33);
xnor U704 (N_704,N_483,In_703);
nor U705 (N_705,In_303,N_482);
or U706 (N_706,In_722,In_257);
and U707 (N_707,In_141,N_229);
nand U708 (N_708,In_354,N_432);
nand U709 (N_709,N_367,N_247);
or U710 (N_710,In_1320,N_479);
or U711 (N_711,In_687,In_275);
or U712 (N_712,N_420,N_25);
nor U713 (N_713,In_990,In_250);
nand U714 (N_714,N_162,In_476);
nand U715 (N_715,In_12,In_213);
and U716 (N_716,N_480,N_463);
xor U717 (N_717,In_562,In_428);
xnor U718 (N_718,N_498,N_310);
and U719 (N_719,In_336,In_1432);
xnor U720 (N_720,In_1420,In_773);
and U721 (N_721,In_568,In_707);
or U722 (N_722,N_183,In_1372);
xor U723 (N_723,In_10,In_1238);
or U724 (N_724,N_270,N_431);
or U725 (N_725,In_7,In_747);
nand U726 (N_726,In_1180,In_591);
nor U727 (N_727,In_151,N_193);
nand U728 (N_728,N_97,In_1249);
nor U729 (N_729,In_1181,In_1465);
xnor U730 (N_730,N_481,In_1147);
or U731 (N_731,In_96,N_243);
nor U732 (N_732,In_807,In_117);
nor U733 (N_733,In_1371,N_88);
or U734 (N_734,N_406,N_399);
nand U735 (N_735,In_9,In_784);
nand U736 (N_736,In_40,In_1254);
nor U737 (N_737,N_40,In_1240);
and U738 (N_738,In_473,In_457);
xor U739 (N_739,N_461,In_929);
or U740 (N_740,In_1030,N_239);
nor U741 (N_741,In_563,In_953);
xnor U742 (N_742,In_300,In_613);
and U743 (N_743,In_833,N_197);
or U744 (N_744,N_433,In_579);
xnor U745 (N_745,In_1227,N_253);
or U746 (N_746,N_124,In_769);
or U747 (N_747,N_8,In_291);
xor U748 (N_748,N_374,N_435);
or U749 (N_749,In_1007,N_135);
and U750 (N_750,In_973,N_174);
or U751 (N_751,N_343,N_735);
nand U752 (N_752,In_1164,N_709);
nor U753 (N_753,In_988,N_519);
xnor U754 (N_754,In_37,N_398);
xnor U755 (N_755,N_586,In_279);
xor U756 (N_756,In_774,N_506);
xnor U757 (N_757,N_572,In_363);
or U758 (N_758,In_507,N_510);
or U759 (N_759,N_43,N_68);
nor U760 (N_760,In_1000,In_358);
nand U761 (N_761,N_609,N_651);
nand U762 (N_762,N_29,N_384);
nor U763 (N_763,N_746,N_418);
and U764 (N_764,N_304,N_24);
xor U765 (N_765,In_425,N_337);
xnor U766 (N_766,In_433,In_758);
nor U767 (N_767,In_278,N_569);
nand U768 (N_768,N_673,In_59);
nand U769 (N_769,In_661,In_698);
and U770 (N_770,In_171,In_682);
and U771 (N_771,In_556,N_667);
nor U772 (N_772,In_61,In_1152);
or U773 (N_773,N_600,In_1491);
or U774 (N_774,In_1162,In_827);
xor U775 (N_775,N_145,N_294);
xnor U776 (N_776,N_723,N_671);
nand U777 (N_777,In_880,In_678);
or U778 (N_778,N_362,In_3);
and U779 (N_779,In_1218,In_1341);
nand U780 (N_780,In_1186,In_916);
nand U781 (N_781,N_738,N_745);
nand U782 (N_782,N_136,N_540);
nand U783 (N_783,In_1184,N_714);
xnor U784 (N_784,N_416,In_478);
nor U785 (N_785,N_446,N_724);
or U786 (N_786,N_221,N_138);
and U787 (N_787,N_694,In_915);
or U788 (N_788,N_439,N_693);
nand U789 (N_789,N_377,N_306);
or U790 (N_790,N_404,N_559);
or U791 (N_791,N_665,In_1179);
nor U792 (N_792,N_635,N_566);
xor U793 (N_793,N_474,N_574);
nor U794 (N_794,In_826,In_1111);
nor U795 (N_795,N_593,N_307);
or U796 (N_796,N_348,N_438);
nor U797 (N_797,In_1172,N_254);
nor U798 (N_798,N_630,N_670);
xnor U799 (N_799,N_530,N_202);
or U800 (N_800,N_710,N_645);
or U801 (N_801,N_289,N_639);
nand U802 (N_802,In_547,N_590);
xor U803 (N_803,In_611,In_1290);
and U804 (N_804,N_397,In_1263);
nor U805 (N_805,N_702,N_594);
xnor U806 (N_806,In_766,N_508);
xor U807 (N_807,N_704,In_1392);
xnor U808 (N_808,In_193,N_619);
xor U809 (N_809,In_200,N_317);
or U810 (N_810,N_338,In_675);
and U811 (N_811,In_1348,In_1442);
nand U812 (N_812,N_255,In_1096);
xnor U813 (N_813,N_41,In_1456);
nor U814 (N_814,In_535,N_653);
and U815 (N_815,N_507,N_451);
nand U816 (N_816,In_1384,In_601);
xor U817 (N_817,In_792,N_580);
nand U818 (N_818,N_168,N_733);
nor U819 (N_819,N_515,N_669);
and U820 (N_820,N_625,N_558);
xor U821 (N_821,In_296,In_838);
nand U822 (N_822,N_376,N_686);
xnor U823 (N_823,In_1389,In_967);
or U824 (N_824,In_1143,N_538);
nor U825 (N_825,In_344,N_685);
or U826 (N_826,N_358,N_747);
xnor U827 (N_827,N_295,N_532);
and U828 (N_828,N_396,N_19);
nor U829 (N_829,N_727,N_663);
xor U830 (N_830,N_466,In_325);
nand U831 (N_831,N_370,N_634);
and U832 (N_832,N_395,In_1486);
nand U833 (N_833,In_304,In_1237);
xor U834 (N_834,N_643,N_741);
and U835 (N_835,In_771,N_329);
nor U836 (N_836,N_245,N_272);
nand U837 (N_837,In_1285,N_208);
or U838 (N_838,N_87,N_291);
nand U839 (N_839,N_649,In_712);
and U840 (N_840,N_617,N_412);
or U841 (N_841,N_212,N_612);
and U842 (N_842,N_555,N_549);
and U843 (N_843,In_1321,N_553);
or U844 (N_844,In_1078,In_1291);
nor U845 (N_845,N_683,N_260);
nand U846 (N_846,In_35,N_263);
xnor U847 (N_847,In_724,N_365);
xor U848 (N_848,In_570,In_892);
and U849 (N_849,N_0,N_533);
nor U850 (N_850,In_1303,In_321);
xnor U851 (N_851,In_1014,N_146);
xor U852 (N_852,N_697,N_195);
or U853 (N_853,In_795,N_749);
xor U854 (N_854,In_1229,In_173);
and U855 (N_855,In_355,N_13);
and U856 (N_856,In_865,In_1356);
and U857 (N_857,In_489,N_51);
and U858 (N_858,In_265,N_616);
xor U859 (N_859,In_1494,N_560);
nor U860 (N_860,N_703,In_770);
xor U861 (N_861,N_632,N_712);
nand U862 (N_862,In_589,In_1401);
nand U863 (N_863,In_820,In_145);
nand U864 (N_864,In_1489,In_1034);
or U865 (N_865,In_1050,N_717);
and U866 (N_866,In_88,In_1132);
xnor U867 (N_867,N_120,N_539);
nand U868 (N_868,In_467,In_1374);
and U869 (N_869,In_791,N_129);
nor U870 (N_870,N_503,In_956);
nand U871 (N_871,N_214,N_677);
nand U872 (N_872,In_605,N_150);
nand U873 (N_873,N_579,In_746);
and U874 (N_874,N_516,N_280);
xnor U875 (N_875,In_26,In_1185);
nor U876 (N_876,N_84,N_568);
xnor U877 (N_877,N_282,N_518);
or U878 (N_878,N_366,N_672);
and U879 (N_879,In_1153,In_588);
xor U880 (N_880,N_198,N_342);
and U881 (N_881,In_786,In_989);
nor U882 (N_882,N_711,In_1244);
and U883 (N_883,N_369,N_534);
and U884 (N_884,N_524,In_429);
nand U885 (N_885,N_567,In_1288);
and U886 (N_886,N_708,In_1060);
or U887 (N_887,In_1191,In_1393);
nor U888 (N_888,N_737,In_910);
nor U889 (N_889,N_611,N_563);
nor U890 (N_890,In_1257,In_705);
nand U891 (N_891,N_675,In_399);
or U892 (N_892,In_1297,N_437);
nand U893 (N_893,N_647,N_514);
nand U894 (N_894,N_107,N_378);
or U895 (N_895,N_535,In_1250);
nor U896 (N_896,N_601,N_472);
nand U897 (N_897,N_290,N_544);
nor U898 (N_898,In_17,N_78);
xnor U899 (N_899,N_606,In_518);
xor U900 (N_900,N_163,In_494);
nand U901 (N_901,In_20,N_464);
and U902 (N_902,N_627,N_722);
nand U903 (N_903,In_22,N_687);
nand U904 (N_904,N_256,N_517);
nand U905 (N_905,N_577,In_788);
nor U906 (N_906,In_1100,In_600);
and U907 (N_907,N_64,In_524);
and U908 (N_908,N_10,N_676);
xor U909 (N_909,In_1493,N_320);
nor U910 (N_910,N_487,N_644);
nor U911 (N_911,N_587,In_1004);
or U912 (N_912,N_633,N_386);
and U913 (N_913,In_897,N_556);
and U914 (N_914,N_261,In_1464);
nand U915 (N_915,In_486,N_608);
or U916 (N_916,N_628,In_140);
nand U917 (N_917,In_1281,N_629);
xnor U918 (N_918,N_720,In_1081);
and U919 (N_919,In_168,In_1167);
or U920 (N_920,N_631,N_442);
nor U921 (N_921,N_554,In_954);
nand U922 (N_922,N_422,In_70);
or U923 (N_923,N_564,In_1459);
nor U924 (N_924,In_289,In_506);
and U925 (N_925,In_175,N_719);
xor U926 (N_926,N_357,N_453);
xnor U927 (N_927,In_1445,N_595);
or U928 (N_928,N_240,In_741);
and U929 (N_929,N_618,N_526);
nand U930 (N_930,In_1260,N_100);
nor U931 (N_931,In_15,N_312);
or U932 (N_932,In_351,N_447);
xnor U933 (N_933,In_1366,N_692);
and U934 (N_934,N_257,N_571);
and U935 (N_935,In_1317,In_918);
nand U936 (N_936,N_748,In_1183);
nor U937 (N_937,N_613,N_281);
nand U938 (N_938,N_330,N_678);
nand U939 (N_939,In_297,N_188);
nor U940 (N_940,N_661,In_1296);
xnor U941 (N_941,In_343,In_364);
nand U942 (N_942,N_591,In_1175);
or U943 (N_943,In_1310,N_499);
and U944 (N_944,In_614,In_208);
or U945 (N_945,N_278,N_185);
or U946 (N_946,N_103,N_734);
and U947 (N_947,N_413,N_565);
xor U948 (N_948,N_592,In_404);
nand U949 (N_949,N_189,N_265);
nor U950 (N_950,N_323,N_696);
nor U951 (N_951,N_484,N_548);
or U952 (N_952,N_557,N_583);
nand U953 (N_953,N_230,N_379);
xor U954 (N_954,N_614,N_184);
xnor U955 (N_955,N_642,N_648);
or U956 (N_956,N_268,N_716);
nand U957 (N_957,N_666,N_144);
and U958 (N_958,N_155,N_715);
and U959 (N_959,In_197,In_757);
and U960 (N_960,In_1141,N_417);
or U961 (N_961,N_660,N_581);
and U962 (N_962,N_536,N_657);
nand U963 (N_963,N_428,N_127);
or U964 (N_964,In_365,N_300);
nand U965 (N_965,N_473,N_383);
nand U966 (N_966,N_602,N_588);
or U967 (N_967,In_125,In_913);
xor U968 (N_968,In_1448,N_264);
xnor U969 (N_969,N_388,In_676);
or U970 (N_970,N_101,N_705);
nand U971 (N_971,N_347,N_596);
or U972 (N_972,N_699,In_697);
xnor U973 (N_973,In_569,In_1188);
and U974 (N_974,N_77,In_1460);
nand U975 (N_975,In_635,N_728);
nor U976 (N_976,In_679,In_1454);
nor U977 (N_977,N_326,N_646);
xor U978 (N_978,N_156,In_987);
or U979 (N_979,In_281,In_934);
nand U980 (N_980,N_679,In_541);
nand U981 (N_981,In_360,In_453);
nand U982 (N_982,N_477,N_680);
nor U983 (N_983,In_650,N_542);
xor U984 (N_984,N_707,N_511);
nor U985 (N_985,In_420,N_537);
nor U986 (N_986,N_743,N_65);
and U987 (N_987,N_324,In_1477);
or U988 (N_988,N_48,N_691);
nor U989 (N_989,In_437,In_982);
nand U990 (N_990,N_465,N_543);
and U991 (N_991,N_3,N_235);
nor U992 (N_992,In_799,In_1407);
nand U993 (N_993,N_528,N_112);
or U994 (N_994,N_216,N_659);
xor U995 (N_995,N_684,N_664);
and U996 (N_996,In_587,N_69);
nor U997 (N_997,N_353,N_314);
xnor U998 (N_998,In_295,In_842);
xnor U999 (N_999,N_681,In_585);
and U1000 (N_1000,N_833,N_522);
or U1001 (N_1001,N_980,N_796);
and U1002 (N_1002,N_866,In_264);
nor U1003 (N_1003,N_801,In_294);
nand U1004 (N_1004,In_258,N_63);
nand U1005 (N_1005,N_509,N_774);
or U1006 (N_1006,N_368,N_809);
and U1007 (N_1007,N_897,N_605);
and U1008 (N_1008,In_73,N_792);
and U1009 (N_1009,N_620,N_785);
or U1010 (N_1010,N_621,N_862);
xor U1011 (N_1011,N_964,N_758);
nor U1012 (N_1012,N_902,N_641);
xnor U1013 (N_1013,N_984,N_932);
or U1014 (N_1014,N_640,N_941);
xor U1015 (N_1015,N_318,N_940);
nor U1016 (N_1016,N_662,N_931);
or U1017 (N_1017,N_847,N_893);
xor U1018 (N_1018,N_7,N_780);
nor U1019 (N_1019,N_979,N_158);
and U1020 (N_1020,N_860,In_728);
nor U1021 (N_1021,N_655,N_882);
xnor U1022 (N_1022,N_892,N_652);
nor U1023 (N_1023,N_907,N_527);
nand U1024 (N_1024,N_901,N_914);
nor U1025 (N_1025,N_190,N_547);
or U1026 (N_1026,N_467,N_726);
xnor U1027 (N_1027,N_871,N_958);
nand U1028 (N_1028,N_636,N_840);
or U1029 (N_1029,N_459,N_551);
or U1030 (N_1030,In_1005,N_529);
or U1031 (N_1031,N_584,N_928);
nand U1032 (N_1032,N_935,In_287);
or U1033 (N_1033,N_763,N_167);
xnor U1034 (N_1034,N_262,In_320);
nor U1035 (N_1035,N_986,N_793);
nor U1036 (N_1036,In_307,N_149);
nor U1037 (N_1037,In_400,N_779);
nand U1038 (N_1038,N_828,N_858);
and U1039 (N_1039,N_761,N_523);
or U1040 (N_1040,N_963,N_423);
nor U1041 (N_1041,N_11,N_757);
nand U1042 (N_1042,In_1176,In_572);
or U1043 (N_1043,N_813,N_844);
xnor U1044 (N_1044,N_390,N_759);
and U1045 (N_1045,In_1065,N_784);
and U1046 (N_1046,In_185,N_890);
or U1047 (N_1047,N_898,N_967);
nor U1048 (N_1048,N_895,N_943);
nand U1049 (N_1049,N_831,In_533);
xnor U1050 (N_1050,N_700,N_525);
nand U1051 (N_1051,N_851,N_807);
and U1052 (N_1052,In_98,N_313);
xor U1053 (N_1053,In_186,N_585);
xor U1054 (N_1054,In_393,N_841);
xor U1055 (N_1055,In_1231,N_997);
or U1056 (N_1056,In_69,In_312);
xor U1057 (N_1057,N_471,In_970);
xor U1058 (N_1058,In_1075,N_576);
nor U1059 (N_1059,N_546,N_995);
nand U1060 (N_1060,In_1315,N_769);
or U1061 (N_1061,In_615,N_919);
nor U1062 (N_1062,In_1298,N_827);
nand U1063 (N_1063,N_604,N_961);
nor U1064 (N_1064,N_731,N_810);
nand U1065 (N_1065,N_730,N_903);
or U1066 (N_1066,N_750,N_781);
nor U1067 (N_1067,In_100,N_953);
nand U1068 (N_1068,N_912,N_624);
or U1069 (N_1069,N_977,N_910);
or U1070 (N_1070,N_288,N_656);
xor U1071 (N_1071,N_440,In_16);
xor U1072 (N_1072,N_22,N_900);
or U1073 (N_1073,N_884,N_883);
xnor U1074 (N_1074,N_765,N_946);
xnor U1075 (N_1075,N_835,N_982);
or U1076 (N_1076,N_531,In_1199);
nand U1077 (N_1077,N_870,N_894);
nor U1078 (N_1078,N_340,N_550);
nor U1079 (N_1079,N_856,N_623);
xor U1080 (N_1080,N_874,N_346);
and U1081 (N_1081,N_775,N_713);
and U1082 (N_1082,N_972,N_821);
or U1083 (N_1083,N_513,N_436);
nand U1084 (N_1084,N_808,N_843);
nor U1085 (N_1085,N_917,N_865);
nor U1086 (N_1086,N_285,N_819);
nor U1087 (N_1087,In_1453,N_415);
xnor U1088 (N_1088,N_545,N_959);
nand U1089 (N_1089,In_253,N_915);
and U1090 (N_1090,N_857,N_832);
xor U1091 (N_1091,In_353,N_921);
nand U1092 (N_1092,N_424,N_133);
nand U1093 (N_1093,In_1122,N_456);
and U1094 (N_1094,N_876,N_861);
and U1095 (N_1095,N_770,N_911);
xnor U1096 (N_1096,N_782,N_983);
xnor U1097 (N_1097,N_790,N_803);
xnor U1098 (N_1098,N_966,N_626);
and U1099 (N_1099,N_913,N_949);
or U1100 (N_1100,In_410,N_881);
xor U1101 (N_1101,In_487,N_930);
and U1102 (N_1102,N_839,N_603);
nor U1103 (N_1103,N_922,N_637);
or U1104 (N_1104,N_850,N_815);
or U1105 (N_1105,N_934,N_981);
nor U1106 (N_1106,N_991,N_674);
nand U1107 (N_1107,N_923,N_875);
nor U1108 (N_1108,In_1117,N_778);
nor U1109 (N_1109,In_299,In_825);
xnor U1110 (N_1110,N_504,N_607);
and U1111 (N_1111,N_962,N_777);
xnor U1112 (N_1112,N_182,N_952);
and U1113 (N_1113,N_501,N_849);
nor U1114 (N_1114,N_753,In_528);
nor U1115 (N_1115,N_806,N_76);
xnor U1116 (N_1116,N_561,N_389);
xnor U1117 (N_1117,In_860,In_465);
nor U1118 (N_1118,In_262,N_948);
nand U1119 (N_1119,N_965,In_1137);
and U1120 (N_1120,N_570,N_246);
nor U1121 (N_1121,N_899,N_879);
nand U1122 (N_1122,In_1334,N_721);
xor U1123 (N_1123,In_240,N_578);
xnor U1124 (N_1124,N_927,In_744);
nor U1125 (N_1125,N_752,N_799);
nand U1126 (N_1126,In_869,In_1280);
xor U1127 (N_1127,N_904,N_970);
nor U1128 (N_1128,N_736,N_824);
nor U1129 (N_1129,N_823,N_994);
nor U1130 (N_1130,N_754,In_595);
nand U1131 (N_1131,In_327,N_725);
and U1132 (N_1132,N_689,In_526);
nand U1133 (N_1133,N_500,In_191);
nand U1134 (N_1134,In_557,N_1);
nand U1135 (N_1135,N_788,N_794);
xor U1136 (N_1136,N_950,N_178);
and U1137 (N_1137,N_762,N_993);
and U1138 (N_1138,N_521,N_125);
nor U1139 (N_1139,N_638,N_744);
nand U1140 (N_1140,In_142,N_957);
xor U1141 (N_1141,N_955,N_772);
nand U1142 (N_1142,N_760,In_936);
and U1143 (N_1143,N_886,N_756);
or U1144 (N_1144,In_190,In_539);
or U1145 (N_1145,N_985,N_951);
nand U1146 (N_1146,N_956,N_742);
and U1147 (N_1147,N_969,N_848);
and U1148 (N_1148,N_266,N_573);
xnor U1149 (N_1149,N_118,N_541);
xnor U1150 (N_1150,In_582,N_854);
or U1151 (N_1151,N_992,N_942);
nand U1152 (N_1152,N_597,In_135);
nor U1153 (N_1153,In_1319,N_802);
nor U1154 (N_1154,N_975,N_493);
or U1155 (N_1155,N_838,N_896);
xnor U1156 (N_1156,N_6,N_925);
nand U1157 (N_1157,In_43,In_739);
nand U1158 (N_1158,N_920,N_817);
xor U1159 (N_1159,N_786,N_695);
nor U1160 (N_1160,In_1377,N_816);
nand U1161 (N_1161,N_333,N_947);
and U1162 (N_1162,N_938,N_974);
xnor U1163 (N_1163,In_306,N_582);
nand U1164 (N_1164,In_1127,N_797);
or U1165 (N_1165,N_199,N_768);
xor U1166 (N_1166,N_939,In_1159);
nand U1167 (N_1167,N_971,N_751);
xor U1168 (N_1168,N_718,N_905);
and U1169 (N_1169,N_906,N_877);
xnor U1170 (N_1170,In_985,N_867);
nand U1171 (N_1171,N_945,N_213);
nor U1172 (N_1172,N_859,N_599);
nand U1173 (N_1173,In_446,N_853);
and U1174 (N_1174,In_938,N_739);
or U1175 (N_1175,N_987,N_864);
nor U1176 (N_1176,In_590,N_916);
nor U1177 (N_1177,N_891,N_783);
xor U1178 (N_1178,In_1026,In_1424);
nand U1179 (N_1179,N_740,In_212);
nor U1180 (N_1180,N_650,N_845);
nand U1181 (N_1181,N_944,N_830);
nand U1182 (N_1182,N_598,N_988);
nor U1183 (N_1183,N_755,In_818);
and U1184 (N_1184,N_688,N_787);
or U1185 (N_1185,N_575,In_439);
or U1186 (N_1186,N_829,N_936);
nand U1187 (N_1187,N_767,In_837);
xor U1188 (N_1188,N_872,In_1436);
and U1189 (N_1189,In_128,N_998);
nand U1190 (N_1190,N_520,N_441);
and U1191 (N_1191,N_771,N_502);
xnor U1192 (N_1192,N_690,N_773);
xor U1193 (N_1193,N_615,N_658);
xnor U1194 (N_1194,N_814,N_873);
xor U1195 (N_1195,In_376,In_1301);
nand U1196 (N_1196,N_846,In_1090);
nor U1197 (N_1197,N_339,N_999);
xnor U1198 (N_1198,N_701,N_834);
nand U1199 (N_1199,In_1012,In_713);
or U1200 (N_1200,N_805,N_800);
or U1201 (N_1201,N_918,In_1044);
or U1202 (N_1202,N_976,N_776);
xor U1203 (N_1203,N_332,N_610);
xor U1204 (N_1204,N_909,N_954);
or U1205 (N_1205,N_552,N_562);
or U1206 (N_1206,N_789,N_305);
nand U1207 (N_1207,N_842,N_622);
nand U1208 (N_1208,N_820,In_176);
xnor U1209 (N_1209,N_360,N_929);
xnor U1210 (N_1210,N_764,N_978);
and U1211 (N_1211,N_880,N_732);
or U1212 (N_1212,N_791,N_812);
nor U1213 (N_1213,In_955,N_826);
nor U1214 (N_1214,N_822,In_501);
or U1215 (N_1215,In_1343,In_342);
or U1216 (N_1216,In_1200,N_589);
and U1217 (N_1217,In_230,N_937);
and U1218 (N_1218,N_512,N_706);
nor U1219 (N_1219,N_448,N_729);
or U1220 (N_1220,N_276,N_885);
or U1221 (N_1221,N_990,N_271);
or U1222 (N_1222,N_352,In_380);
and U1223 (N_1223,N_344,N_863);
xor U1224 (N_1224,N_405,N_98);
or U1225 (N_1225,N_795,N_924);
nor U1226 (N_1226,N_878,N_505);
or U1227 (N_1227,In_1361,N_888);
xnor U1228 (N_1228,N_852,N_668);
xnor U1229 (N_1229,N_409,N_478);
nand U1230 (N_1230,In_976,N_682);
or U1231 (N_1231,N_157,N_968);
and U1232 (N_1232,N_798,In_276);
xor U1233 (N_1233,N_989,N_868);
or U1234 (N_1234,N_837,N_933);
nor U1235 (N_1235,N_960,N_855);
nor U1236 (N_1236,N_889,N_825);
and U1237 (N_1237,In_1086,N_364);
nor U1238 (N_1238,In_1055,N_887);
and U1239 (N_1239,In_889,N_869);
nand U1240 (N_1240,In_1058,N_926);
and U1241 (N_1241,N_44,N_654);
nand U1242 (N_1242,N_818,In_715);
or U1243 (N_1243,N_996,N_973);
and U1244 (N_1244,N_908,N_811);
nor U1245 (N_1245,In_338,In_522);
nand U1246 (N_1246,In_367,N_766);
xor U1247 (N_1247,N_242,In_756);
or U1248 (N_1248,In_948,N_804);
nor U1249 (N_1249,N_836,N_698);
nand U1250 (N_1250,N_1065,N_1008);
or U1251 (N_1251,N_1153,N_1126);
xor U1252 (N_1252,N_1034,N_1172);
or U1253 (N_1253,N_1243,N_1030);
xor U1254 (N_1254,N_1085,N_1188);
xnor U1255 (N_1255,N_1209,N_1148);
or U1256 (N_1256,N_1011,N_1158);
and U1257 (N_1257,N_1194,N_1131);
or U1258 (N_1258,N_1138,N_1039);
nand U1259 (N_1259,N_1101,N_1185);
or U1260 (N_1260,N_1244,N_1060);
xor U1261 (N_1261,N_1087,N_1140);
and U1262 (N_1262,N_1130,N_1088);
nor U1263 (N_1263,N_1061,N_1068);
xnor U1264 (N_1264,N_1227,N_1203);
nor U1265 (N_1265,N_1136,N_1178);
xor U1266 (N_1266,N_1013,N_1116);
or U1267 (N_1267,N_1122,N_1142);
xnor U1268 (N_1268,N_1047,N_1173);
nand U1269 (N_1269,N_1231,N_1204);
xor U1270 (N_1270,N_1189,N_1151);
nand U1271 (N_1271,N_1191,N_1001);
and U1272 (N_1272,N_1134,N_1081);
nand U1273 (N_1273,N_1141,N_1053);
xor U1274 (N_1274,N_1024,N_1006);
nand U1275 (N_1275,N_1202,N_1145);
xnor U1276 (N_1276,N_1124,N_1089);
and U1277 (N_1277,N_1070,N_1223);
and U1278 (N_1278,N_1029,N_1078);
nand U1279 (N_1279,N_1105,N_1082);
xor U1280 (N_1280,N_1120,N_1071);
and U1281 (N_1281,N_1051,N_1248);
xnor U1282 (N_1282,N_1009,N_1111);
xnor U1283 (N_1283,N_1055,N_1159);
nor U1284 (N_1284,N_1230,N_1043);
and U1285 (N_1285,N_1176,N_1035);
nand U1286 (N_1286,N_1000,N_1002);
or U1287 (N_1287,N_1196,N_1219);
and U1288 (N_1288,N_1031,N_1090);
or U1289 (N_1289,N_1193,N_1183);
nand U1290 (N_1290,N_1229,N_1072);
or U1291 (N_1291,N_1163,N_1137);
nand U1292 (N_1292,N_1160,N_1226);
or U1293 (N_1293,N_1046,N_1113);
nand U1294 (N_1294,N_1077,N_1074);
nor U1295 (N_1295,N_1169,N_1170);
or U1296 (N_1296,N_1125,N_1014);
or U1297 (N_1297,N_1118,N_1215);
and U1298 (N_1298,N_1040,N_1063);
nor U1299 (N_1299,N_1218,N_1239);
xor U1300 (N_1300,N_1012,N_1049);
xnor U1301 (N_1301,N_1207,N_1144);
and U1302 (N_1302,N_1018,N_1042);
and U1303 (N_1303,N_1073,N_1208);
nand U1304 (N_1304,N_1161,N_1044);
nor U1305 (N_1305,N_1057,N_1224);
nand U1306 (N_1306,N_1247,N_1076);
xnor U1307 (N_1307,N_1119,N_1147);
nand U1308 (N_1308,N_1184,N_1020);
or U1309 (N_1309,N_1109,N_1028);
and U1310 (N_1310,N_1036,N_1143);
and U1311 (N_1311,N_1180,N_1033);
or U1312 (N_1312,N_1080,N_1240);
nand U1313 (N_1313,N_1054,N_1106);
xor U1314 (N_1314,N_1093,N_1171);
xor U1315 (N_1315,N_1015,N_1238);
nor U1316 (N_1316,N_1017,N_1110);
and U1317 (N_1317,N_1233,N_1175);
and U1318 (N_1318,N_1146,N_1177);
nand U1319 (N_1319,N_1075,N_1064);
or U1320 (N_1320,N_1007,N_1195);
nor U1321 (N_1321,N_1149,N_1100);
xor U1322 (N_1322,N_1212,N_1132);
nor U1323 (N_1323,N_1222,N_1025);
and U1324 (N_1324,N_1135,N_1199);
nand U1325 (N_1325,N_1150,N_1117);
nand U1326 (N_1326,N_1198,N_1127);
nand U1327 (N_1327,N_1058,N_1200);
nor U1328 (N_1328,N_1108,N_1104);
nor U1329 (N_1329,N_1133,N_1050);
xor U1330 (N_1330,N_1016,N_1112);
or U1331 (N_1331,N_1056,N_1242);
or U1332 (N_1332,N_1181,N_1022);
xor U1333 (N_1333,N_1048,N_1084);
nor U1334 (N_1334,N_1079,N_1246);
or U1335 (N_1335,N_1190,N_1155);
and U1336 (N_1336,N_1096,N_1211);
xor U1337 (N_1337,N_1164,N_1026);
and U1338 (N_1338,N_1004,N_1167);
nor U1339 (N_1339,N_1027,N_1019);
nand U1340 (N_1340,N_1192,N_1201);
nor U1341 (N_1341,N_1156,N_1095);
nor U1342 (N_1342,N_1069,N_1232);
and U1343 (N_1343,N_1052,N_1066);
nand U1344 (N_1344,N_1216,N_1092);
xor U1345 (N_1345,N_1234,N_1228);
nor U1346 (N_1346,N_1086,N_1123);
xnor U1347 (N_1347,N_1091,N_1010);
and U1348 (N_1348,N_1237,N_1179);
and U1349 (N_1349,N_1062,N_1221);
and U1350 (N_1350,N_1083,N_1186);
xnor U1351 (N_1351,N_1129,N_1162);
xor U1352 (N_1352,N_1235,N_1103);
nor U1353 (N_1353,N_1213,N_1128);
or U1354 (N_1354,N_1182,N_1107);
nor U1355 (N_1355,N_1005,N_1139);
xor U1356 (N_1356,N_1121,N_1097);
nor U1357 (N_1357,N_1045,N_1210);
or U1358 (N_1358,N_1099,N_1041);
or U1359 (N_1359,N_1220,N_1098);
and U1360 (N_1360,N_1157,N_1152);
nand U1361 (N_1361,N_1037,N_1197);
or U1362 (N_1362,N_1245,N_1023);
xnor U1363 (N_1363,N_1114,N_1094);
nand U1364 (N_1364,N_1166,N_1067);
nor U1365 (N_1365,N_1217,N_1059);
and U1366 (N_1366,N_1187,N_1236);
nand U1367 (N_1367,N_1168,N_1102);
xor U1368 (N_1368,N_1038,N_1032);
nand U1369 (N_1369,N_1214,N_1206);
nor U1370 (N_1370,N_1249,N_1205);
or U1371 (N_1371,N_1241,N_1154);
nand U1372 (N_1372,N_1115,N_1174);
nor U1373 (N_1373,N_1021,N_1165);
or U1374 (N_1374,N_1003,N_1225);
and U1375 (N_1375,N_1120,N_1037);
nand U1376 (N_1376,N_1045,N_1151);
nor U1377 (N_1377,N_1083,N_1192);
nand U1378 (N_1378,N_1037,N_1073);
xnor U1379 (N_1379,N_1215,N_1090);
or U1380 (N_1380,N_1121,N_1215);
nand U1381 (N_1381,N_1078,N_1229);
or U1382 (N_1382,N_1024,N_1124);
or U1383 (N_1383,N_1159,N_1197);
or U1384 (N_1384,N_1096,N_1124);
xor U1385 (N_1385,N_1169,N_1056);
nor U1386 (N_1386,N_1002,N_1247);
or U1387 (N_1387,N_1031,N_1071);
nand U1388 (N_1388,N_1045,N_1241);
and U1389 (N_1389,N_1037,N_1045);
nand U1390 (N_1390,N_1228,N_1239);
nor U1391 (N_1391,N_1080,N_1199);
nor U1392 (N_1392,N_1100,N_1194);
xor U1393 (N_1393,N_1057,N_1159);
xor U1394 (N_1394,N_1153,N_1183);
nand U1395 (N_1395,N_1132,N_1023);
nor U1396 (N_1396,N_1221,N_1184);
xor U1397 (N_1397,N_1032,N_1108);
or U1398 (N_1398,N_1180,N_1039);
nor U1399 (N_1399,N_1193,N_1151);
and U1400 (N_1400,N_1116,N_1212);
or U1401 (N_1401,N_1213,N_1122);
or U1402 (N_1402,N_1034,N_1010);
and U1403 (N_1403,N_1192,N_1123);
or U1404 (N_1404,N_1045,N_1152);
or U1405 (N_1405,N_1075,N_1097);
nor U1406 (N_1406,N_1243,N_1209);
and U1407 (N_1407,N_1037,N_1000);
nand U1408 (N_1408,N_1204,N_1029);
nor U1409 (N_1409,N_1223,N_1129);
or U1410 (N_1410,N_1227,N_1092);
nand U1411 (N_1411,N_1157,N_1010);
and U1412 (N_1412,N_1083,N_1051);
nand U1413 (N_1413,N_1101,N_1152);
or U1414 (N_1414,N_1167,N_1136);
nand U1415 (N_1415,N_1212,N_1204);
nor U1416 (N_1416,N_1026,N_1114);
or U1417 (N_1417,N_1000,N_1070);
xnor U1418 (N_1418,N_1066,N_1031);
and U1419 (N_1419,N_1208,N_1019);
or U1420 (N_1420,N_1054,N_1058);
nor U1421 (N_1421,N_1113,N_1168);
and U1422 (N_1422,N_1039,N_1028);
or U1423 (N_1423,N_1187,N_1233);
nor U1424 (N_1424,N_1138,N_1246);
nor U1425 (N_1425,N_1149,N_1134);
nand U1426 (N_1426,N_1083,N_1208);
and U1427 (N_1427,N_1091,N_1073);
nor U1428 (N_1428,N_1177,N_1204);
nand U1429 (N_1429,N_1248,N_1081);
or U1430 (N_1430,N_1199,N_1046);
nand U1431 (N_1431,N_1130,N_1128);
nand U1432 (N_1432,N_1195,N_1117);
xor U1433 (N_1433,N_1182,N_1112);
nor U1434 (N_1434,N_1014,N_1230);
and U1435 (N_1435,N_1122,N_1096);
and U1436 (N_1436,N_1221,N_1006);
or U1437 (N_1437,N_1074,N_1239);
nand U1438 (N_1438,N_1178,N_1123);
or U1439 (N_1439,N_1017,N_1197);
xnor U1440 (N_1440,N_1117,N_1101);
xnor U1441 (N_1441,N_1191,N_1185);
xnor U1442 (N_1442,N_1152,N_1172);
nor U1443 (N_1443,N_1212,N_1020);
xor U1444 (N_1444,N_1152,N_1184);
or U1445 (N_1445,N_1108,N_1245);
nand U1446 (N_1446,N_1015,N_1060);
xnor U1447 (N_1447,N_1233,N_1077);
or U1448 (N_1448,N_1163,N_1064);
xnor U1449 (N_1449,N_1063,N_1092);
nor U1450 (N_1450,N_1225,N_1131);
xnor U1451 (N_1451,N_1171,N_1074);
or U1452 (N_1452,N_1144,N_1044);
xnor U1453 (N_1453,N_1001,N_1246);
nor U1454 (N_1454,N_1232,N_1173);
nor U1455 (N_1455,N_1245,N_1183);
nor U1456 (N_1456,N_1216,N_1090);
or U1457 (N_1457,N_1169,N_1246);
nor U1458 (N_1458,N_1169,N_1106);
and U1459 (N_1459,N_1205,N_1109);
and U1460 (N_1460,N_1138,N_1122);
xor U1461 (N_1461,N_1035,N_1187);
and U1462 (N_1462,N_1054,N_1086);
xor U1463 (N_1463,N_1179,N_1110);
and U1464 (N_1464,N_1092,N_1001);
xor U1465 (N_1465,N_1029,N_1161);
and U1466 (N_1466,N_1144,N_1082);
and U1467 (N_1467,N_1108,N_1095);
nand U1468 (N_1468,N_1078,N_1190);
or U1469 (N_1469,N_1195,N_1160);
xnor U1470 (N_1470,N_1060,N_1137);
nand U1471 (N_1471,N_1248,N_1195);
nand U1472 (N_1472,N_1186,N_1047);
nor U1473 (N_1473,N_1176,N_1078);
and U1474 (N_1474,N_1178,N_1175);
or U1475 (N_1475,N_1076,N_1130);
and U1476 (N_1476,N_1234,N_1079);
or U1477 (N_1477,N_1239,N_1069);
and U1478 (N_1478,N_1127,N_1124);
nor U1479 (N_1479,N_1143,N_1043);
xor U1480 (N_1480,N_1125,N_1204);
nor U1481 (N_1481,N_1125,N_1249);
xnor U1482 (N_1482,N_1175,N_1227);
nand U1483 (N_1483,N_1180,N_1232);
xnor U1484 (N_1484,N_1095,N_1015);
nand U1485 (N_1485,N_1174,N_1076);
xor U1486 (N_1486,N_1241,N_1022);
nor U1487 (N_1487,N_1092,N_1234);
or U1488 (N_1488,N_1013,N_1023);
and U1489 (N_1489,N_1054,N_1074);
or U1490 (N_1490,N_1170,N_1051);
or U1491 (N_1491,N_1203,N_1032);
and U1492 (N_1492,N_1048,N_1226);
xnor U1493 (N_1493,N_1165,N_1190);
or U1494 (N_1494,N_1051,N_1011);
and U1495 (N_1495,N_1082,N_1003);
nand U1496 (N_1496,N_1130,N_1133);
or U1497 (N_1497,N_1024,N_1154);
nand U1498 (N_1498,N_1120,N_1140);
nor U1499 (N_1499,N_1240,N_1183);
xnor U1500 (N_1500,N_1427,N_1326);
xnor U1501 (N_1501,N_1478,N_1464);
nand U1502 (N_1502,N_1444,N_1308);
nand U1503 (N_1503,N_1268,N_1447);
and U1504 (N_1504,N_1455,N_1417);
xnor U1505 (N_1505,N_1275,N_1419);
and U1506 (N_1506,N_1484,N_1305);
nand U1507 (N_1507,N_1259,N_1420);
nand U1508 (N_1508,N_1365,N_1441);
or U1509 (N_1509,N_1440,N_1396);
or U1510 (N_1510,N_1258,N_1357);
xnor U1511 (N_1511,N_1261,N_1466);
xnor U1512 (N_1512,N_1352,N_1250);
nor U1513 (N_1513,N_1371,N_1462);
nor U1514 (N_1514,N_1297,N_1376);
nand U1515 (N_1515,N_1392,N_1412);
nor U1516 (N_1516,N_1318,N_1313);
or U1517 (N_1517,N_1360,N_1349);
nor U1518 (N_1518,N_1348,N_1272);
nor U1519 (N_1519,N_1322,N_1362);
xnor U1520 (N_1520,N_1351,N_1446);
nor U1521 (N_1521,N_1283,N_1435);
xor U1522 (N_1522,N_1428,N_1255);
nor U1523 (N_1523,N_1418,N_1271);
or U1524 (N_1524,N_1468,N_1398);
xor U1525 (N_1525,N_1451,N_1469);
nand U1526 (N_1526,N_1498,N_1397);
nand U1527 (N_1527,N_1356,N_1491);
and U1528 (N_1528,N_1363,N_1285);
and U1529 (N_1529,N_1452,N_1324);
or U1530 (N_1530,N_1408,N_1264);
xor U1531 (N_1531,N_1463,N_1299);
or U1532 (N_1532,N_1343,N_1485);
nor U1533 (N_1533,N_1367,N_1339);
and U1534 (N_1534,N_1415,N_1267);
xnor U1535 (N_1535,N_1496,N_1253);
or U1536 (N_1536,N_1486,N_1375);
nand U1537 (N_1537,N_1424,N_1390);
xnor U1538 (N_1538,N_1430,N_1393);
nand U1539 (N_1539,N_1345,N_1474);
nand U1540 (N_1540,N_1379,N_1301);
or U1541 (N_1541,N_1481,N_1429);
and U1542 (N_1542,N_1361,N_1304);
xor U1543 (N_1543,N_1274,N_1369);
and U1544 (N_1544,N_1286,N_1309);
nor U1545 (N_1545,N_1494,N_1328);
and U1546 (N_1546,N_1273,N_1437);
or U1547 (N_1547,N_1374,N_1456);
nand U1548 (N_1548,N_1350,N_1317);
or U1549 (N_1549,N_1282,N_1316);
nand U1550 (N_1550,N_1329,N_1284);
and U1551 (N_1551,N_1459,N_1262);
or U1552 (N_1552,N_1405,N_1497);
nor U1553 (N_1553,N_1490,N_1473);
nor U1554 (N_1554,N_1394,N_1277);
and U1555 (N_1555,N_1260,N_1439);
and U1556 (N_1556,N_1487,N_1460);
or U1557 (N_1557,N_1383,N_1354);
nor U1558 (N_1558,N_1499,N_1296);
nand U1559 (N_1559,N_1436,N_1421);
xnor U1560 (N_1560,N_1332,N_1422);
or U1561 (N_1561,N_1377,N_1409);
and U1562 (N_1562,N_1450,N_1489);
xor U1563 (N_1563,N_1334,N_1406);
xnor U1564 (N_1564,N_1461,N_1381);
nand U1565 (N_1565,N_1280,N_1373);
nand U1566 (N_1566,N_1287,N_1288);
and U1567 (N_1567,N_1300,N_1384);
and U1568 (N_1568,N_1327,N_1294);
nor U1569 (N_1569,N_1411,N_1290);
xnor U1570 (N_1570,N_1404,N_1298);
nand U1571 (N_1571,N_1279,N_1303);
xor U1572 (N_1572,N_1346,N_1302);
nand U1573 (N_1573,N_1458,N_1425);
and U1574 (N_1574,N_1488,N_1414);
xnor U1575 (N_1575,N_1465,N_1330);
nor U1576 (N_1576,N_1493,N_1403);
nand U1577 (N_1577,N_1331,N_1407);
and U1578 (N_1578,N_1442,N_1292);
nor U1579 (N_1579,N_1378,N_1470);
xor U1580 (N_1580,N_1320,N_1480);
nand U1581 (N_1581,N_1380,N_1257);
nand U1582 (N_1582,N_1479,N_1289);
nand U1583 (N_1583,N_1337,N_1389);
nor U1584 (N_1584,N_1431,N_1395);
and U1585 (N_1585,N_1453,N_1336);
nor U1586 (N_1586,N_1342,N_1310);
xnor U1587 (N_1587,N_1410,N_1454);
nor U1588 (N_1588,N_1385,N_1370);
nor U1589 (N_1589,N_1266,N_1457);
and U1590 (N_1590,N_1483,N_1340);
and U1591 (N_1591,N_1423,N_1311);
nand U1592 (N_1592,N_1438,N_1387);
nor U1593 (N_1593,N_1335,N_1416);
or U1594 (N_1594,N_1449,N_1359);
and U1595 (N_1595,N_1319,N_1281);
nor U1596 (N_1596,N_1386,N_1291);
nor U1597 (N_1597,N_1364,N_1426);
and U1598 (N_1598,N_1443,N_1471);
nor U1599 (N_1599,N_1321,N_1269);
nor U1600 (N_1600,N_1323,N_1445);
or U1601 (N_1601,N_1399,N_1353);
nand U1602 (N_1602,N_1413,N_1344);
and U1603 (N_1603,N_1358,N_1400);
and U1604 (N_1604,N_1256,N_1293);
xnor U1605 (N_1605,N_1448,N_1315);
nand U1606 (N_1606,N_1402,N_1475);
and U1607 (N_1607,N_1355,N_1270);
xnor U1608 (N_1608,N_1333,N_1314);
and U1609 (N_1609,N_1276,N_1492);
xnor U1610 (N_1610,N_1251,N_1312);
and U1611 (N_1611,N_1368,N_1265);
xor U1612 (N_1612,N_1347,N_1254);
or U1613 (N_1613,N_1476,N_1366);
xnor U1614 (N_1614,N_1382,N_1434);
and U1615 (N_1615,N_1372,N_1388);
nor U1616 (N_1616,N_1482,N_1391);
nor U1617 (N_1617,N_1467,N_1495);
and U1618 (N_1618,N_1433,N_1306);
and U1619 (N_1619,N_1252,N_1325);
nor U1620 (N_1620,N_1432,N_1263);
xnor U1621 (N_1621,N_1278,N_1295);
or U1622 (N_1622,N_1338,N_1477);
or U1623 (N_1623,N_1401,N_1472);
nor U1624 (N_1624,N_1341,N_1307);
and U1625 (N_1625,N_1250,N_1445);
and U1626 (N_1626,N_1269,N_1268);
and U1627 (N_1627,N_1262,N_1364);
xor U1628 (N_1628,N_1350,N_1412);
nor U1629 (N_1629,N_1444,N_1273);
and U1630 (N_1630,N_1403,N_1446);
and U1631 (N_1631,N_1294,N_1304);
nor U1632 (N_1632,N_1253,N_1448);
or U1633 (N_1633,N_1291,N_1412);
or U1634 (N_1634,N_1407,N_1312);
nor U1635 (N_1635,N_1256,N_1476);
xnor U1636 (N_1636,N_1471,N_1395);
and U1637 (N_1637,N_1419,N_1432);
and U1638 (N_1638,N_1276,N_1358);
nand U1639 (N_1639,N_1273,N_1439);
nand U1640 (N_1640,N_1258,N_1333);
or U1641 (N_1641,N_1282,N_1481);
nor U1642 (N_1642,N_1364,N_1438);
or U1643 (N_1643,N_1425,N_1472);
xor U1644 (N_1644,N_1347,N_1280);
xnor U1645 (N_1645,N_1258,N_1389);
nor U1646 (N_1646,N_1296,N_1334);
xnor U1647 (N_1647,N_1488,N_1384);
and U1648 (N_1648,N_1377,N_1347);
nor U1649 (N_1649,N_1367,N_1453);
nor U1650 (N_1650,N_1379,N_1384);
or U1651 (N_1651,N_1343,N_1278);
or U1652 (N_1652,N_1387,N_1334);
or U1653 (N_1653,N_1301,N_1453);
nor U1654 (N_1654,N_1256,N_1301);
xor U1655 (N_1655,N_1428,N_1273);
nor U1656 (N_1656,N_1429,N_1369);
or U1657 (N_1657,N_1387,N_1271);
nand U1658 (N_1658,N_1271,N_1281);
nor U1659 (N_1659,N_1444,N_1400);
and U1660 (N_1660,N_1461,N_1437);
nor U1661 (N_1661,N_1447,N_1424);
nor U1662 (N_1662,N_1374,N_1412);
xor U1663 (N_1663,N_1339,N_1385);
and U1664 (N_1664,N_1425,N_1334);
nand U1665 (N_1665,N_1491,N_1291);
xnor U1666 (N_1666,N_1449,N_1274);
xor U1667 (N_1667,N_1489,N_1498);
and U1668 (N_1668,N_1281,N_1431);
or U1669 (N_1669,N_1296,N_1493);
xnor U1670 (N_1670,N_1373,N_1346);
and U1671 (N_1671,N_1494,N_1413);
or U1672 (N_1672,N_1267,N_1479);
or U1673 (N_1673,N_1388,N_1488);
xnor U1674 (N_1674,N_1370,N_1330);
nor U1675 (N_1675,N_1294,N_1313);
xor U1676 (N_1676,N_1258,N_1250);
and U1677 (N_1677,N_1425,N_1362);
or U1678 (N_1678,N_1398,N_1445);
or U1679 (N_1679,N_1478,N_1309);
and U1680 (N_1680,N_1313,N_1365);
nor U1681 (N_1681,N_1441,N_1358);
or U1682 (N_1682,N_1443,N_1307);
and U1683 (N_1683,N_1408,N_1290);
or U1684 (N_1684,N_1473,N_1364);
and U1685 (N_1685,N_1490,N_1353);
and U1686 (N_1686,N_1268,N_1486);
nand U1687 (N_1687,N_1458,N_1264);
nand U1688 (N_1688,N_1288,N_1325);
nand U1689 (N_1689,N_1338,N_1368);
nand U1690 (N_1690,N_1492,N_1432);
xor U1691 (N_1691,N_1371,N_1476);
xor U1692 (N_1692,N_1475,N_1286);
xor U1693 (N_1693,N_1291,N_1297);
nand U1694 (N_1694,N_1403,N_1378);
nor U1695 (N_1695,N_1404,N_1395);
nor U1696 (N_1696,N_1492,N_1280);
nand U1697 (N_1697,N_1435,N_1415);
nand U1698 (N_1698,N_1437,N_1279);
xor U1699 (N_1699,N_1276,N_1326);
xor U1700 (N_1700,N_1349,N_1277);
xor U1701 (N_1701,N_1324,N_1326);
or U1702 (N_1702,N_1435,N_1421);
xnor U1703 (N_1703,N_1495,N_1454);
xnor U1704 (N_1704,N_1432,N_1423);
and U1705 (N_1705,N_1432,N_1294);
nand U1706 (N_1706,N_1372,N_1448);
xnor U1707 (N_1707,N_1260,N_1402);
nor U1708 (N_1708,N_1451,N_1305);
or U1709 (N_1709,N_1295,N_1495);
nor U1710 (N_1710,N_1355,N_1352);
or U1711 (N_1711,N_1270,N_1442);
nor U1712 (N_1712,N_1305,N_1474);
or U1713 (N_1713,N_1333,N_1463);
nand U1714 (N_1714,N_1290,N_1259);
nor U1715 (N_1715,N_1420,N_1353);
nor U1716 (N_1716,N_1480,N_1422);
and U1717 (N_1717,N_1411,N_1320);
xnor U1718 (N_1718,N_1251,N_1373);
nand U1719 (N_1719,N_1425,N_1358);
and U1720 (N_1720,N_1383,N_1392);
xnor U1721 (N_1721,N_1465,N_1285);
xor U1722 (N_1722,N_1321,N_1366);
xnor U1723 (N_1723,N_1289,N_1497);
nand U1724 (N_1724,N_1263,N_1255);
nand U1725 (N_1725,N_1393,N_1327);
or U1726 (N_1726,N_1280,N_1489);
nor U1727 (N_1727,N_1384,N_1310);
xor U1728 (N_1728,N_1443,N_1473);
and U1729 (N_1729,N_1293,N_1487);
and U1730 (N_1730,N_1384,N_1421);
or U1731 (N_1731,N_1368,N_1305);
and U1732 (N_1732,N_1497,N_1444);
and U1733 (N_1733,N_1427,N_1438);
and U1734 (N_1734,N_1341,N_1434);
xor U1735 (N_1735,N_1421,N_1337);
nand U1736 (N_1736,N_1421,N_1336);
or U1737 (N_1737,N_1458,N_1379);
nor U1738 (N_1738,N_1351,N_1441);
or U1739 (N_1739,N_1456,N_1413);
nand U1740 (N_1740,N_1396,N_1366);
nand U1741 (N_1741,N_1473,N_1272);
or U1742 (N_1742,N_1361,N_1287);
and U1743 (N_1743,N_1496,N_1333);
xor U1744 (N_1744,N_1489,N_1392);
xnor U1745 (N_1745,N_1392,N_1395);
and U1746 (N_1746,N_1466,N_1286);
nand U1747 (N_1747,N_1347,N_1266);
xor U1748 (N_1748,N_1328,N_1308);
xnor U1749 (N_1749,N_1352,N_1402);
or U1750 (N_1750,N_1647,N_1506);
nor U1751 (N_1751,N_1604,N_1714);
and U1752 (N_1752,N_1706,N_1503);
xnor U1753 (N_1753,N_1513,N_1615);
nor U1754 (N_1754,N_1687,N_1578);
xor U1755 (N_1755,N_1605,N_1542);
xnor U1756 (N_1756,N_1616,N_1569);
and U1757 (N_1757,N_1568,N_1594);
and U1758 (N_1758,N_1638,N_1626);
xnor U1759 (N_1759,N_1514,N_1662);
or U1760 (N_1760,N_1587,N_1732);
nand U1761 (N_1761,N_1510,N_1711);
nor U1762 (N_1762,N_1674,N_1689);
nor U1763 (N_1763,N_1541,N_1606);
nand U1764 (N_1764,N_1637,N_1565);
or U1765 (N_1765,N_1535,N_1737);
nor U1766 (N_1766,N_1658,N_1553);
xnor U1767 (N_1767,N_1531,N_1611);
xor U1768 (N_1768,N_1505,N_1559);
xnor U1769 (N_1769,N_1718,N_1533);
or U1770 (N_1770,N_1666,N_1555);
or U1771 (N_1771,N_1585,N_1546);
or U1772 (N_1772,N_1598,N_1523);
xnor U1773 (N_1773,N_1702,N_1614);
nand U1774 (N_1774,N_1726,N_1599);
nor U1775 (N_1775,N_1654,N_1511);
or U1776 (N_1776,N_1592,N_1691);
or U1777 (N_1777,N_1669,N_1620);
nor U1778 (N_1778,N_1504,N_1566);
and U1779 (N_1779,N_1748,N_1704);
xor U1780 (N_1780,N_1622,N_1636);
nand U1781 (N_1781,N_1625,N_1683);
nor U1782 (N_1782,N_1558,N_1619);
nand U1783 (N_1783,N_1629,N_1652);
nand U1784 (N_1784,N_1593,N_1602);
nor U1785 (N_1785,N_1573,N_1534);
or U1786 (N_1786,N_1586,N_1618);
xor U1787 (N_1787,N_1589,N_1627);
nand U1788 (N_1788,N_1730,N_1590);
or U1789 (N_1789,N_1639,N_1635);
nor U1790 (N_1790,N_1547,N_1676);
nand U1791 (N_1791,N_1610,N_1608);
nor U1792 (N_1792,N_1551,N_1725);
nand U1793 (N_1793,N_1717,N_1507);
nand U1794 (N_1794,N_1684,N_1664);
or U1795 (N_1795,N_1663,N_1747);
nand U1796 (N_1796,N_1649,N_1650);
and U1797 (N_1797,N_1502,N_1716);
and U1798 (N_1798,N_1544,N_1562);
or U1799 (N_1799,N_1520,N_1517);
xnor U1800 (N_1800,N_1521,N_1540);
nand U1801 (N_1801,N_1576,N_1681);
or U1802 (N_1802,N_1697,N_1731);
nand U1803 (N_1803,N_1537,N_1550);
and U1804 (N_1804,N_1656,N_1524);
and U1805 (N_1805,N_1686,N_1612);
xnor U1806 (N_1806,N_1575,N_1528);
nor U1807 (N_1807,N_1539,N_1709);
or U1808 (N_1808,N_1713,N_1582);
or U1809 (N_1809,N_1668,N_1660);
nand U1810 (N_1810,N_1705,N_1560);
or U1811 (N_1811,N_1563,N_1557);
xnor U1812 (N_1812,N_1742,N_1740);
nand U1813 (N_1813,N_1538,N_1549);
or U1814 (N_1814,N_1543,N_1679);
and U1815 (N_1815,N_1579,N_1518);
nor U1816 (N_1816,N_1703,N_1548);
or U1817 (N_1817,N_1500,N_1675);
nor U1818 (N_1818,N_1532,N_1600);
or U1819 (N_1819,N_1634,N_1692);
and U1820 (N_1820,N_1583,N_1745);
or U1821 (N_1821,N_1688,N_1596);
or U1822 (N_1822,N_1655,N_1741);
or U1823 (N_1823,N_1722,N_1595);
nor U1824 (N_1824,N_1671,N_1597);
or U1825 (N_1825,N_1685,N_1603);
or U1826 (N_1826,N_1530,N_1670);
xor U1827 (N_1827,N_1640,N_1651);
or U1828 (N_1828,N_1693,N_1719);
and U1829 (N_1829,N_1648,N_1633);
nand U1830 (N_1830,N_1574,N_1645);
xnor U1831 (N_1831,N_1723,N_1581);
nor U1832 (N_1832,N_1545,N_1571);
xnor U1833 (N_1833,N_1708,N_1749);
nor U1834 (N_1834,N_1694,N_1617);
nor U1835 (N_1835,N_1501,N_1728);
or U1836 (N_1836,N_1712,N_1727);
or U1837 (N_1837,N_1623,N_1659);
xnor U1838 (N_1838,N_1721,N_1509);
xnor U1839 (N_1839,N_1696,N_1536);
xnor U1840 (N_1840,N_1621,N_1577);
and U1841 (N_1841,N_1665,N_1552);
and U1842 (N_1842,N_1522,N_1529);
or U1843 (N_1843,N_1734,N_1729);
nand U1844 (N_1844,N_1690,N_1653);
xor U1845 (N_1845,N_1746,N_1570);
xnor U1846 (N_1846,N_1630,N_1743);
or U1847 (N_1847,N_1601,N_1588);
or U1848 (N_1848,N_1739,N_1682);
or U1849 (N_1849,N_1519,N_1515);
or U1850 (N_1850,N_1698,N_1673);
nor U1851 (N_1851,N_1657,N_1672);
nor U1852 (N_1852,N_1632,N_1642);
or U1853 (N_1853,N_1516,N_1607);
and U1854 (N_1854,N_1580,N_1609);
and U1855 (N_1855,N_1744,N_1564);
nor U1856 (N_1856,N_1526,N_1613);
or U1857 (N_1857,N_1707,N_1591);
nand U1858 (N_1858,N_1715,N_1661);
nor U1859 (N_1859,N_1720,N_1677);
xor U1860 (N_1860,N_1646,N_1628);
nand U1861 (N_1861,N_1508,N_1724);
and U1862 (N_1862,N_1701,N_1643);
nor U1863 (N_1863,N_1700,N_1584);
xnor U1864 (N_1864,N_1554,N_1738);
or U1865 (N_1865,N_1699,N_1710);
and U1866 (N_1866,N_1512,N_1631);
or U1867 (N_1867,N_1561,N_1736);
or U1868 (N_1868,N_1527,N_1678);
nand U1869 (N_1869,N_1556,N_1624);
xnor U1870 (N_1870,N_1567,N_1733);
xor U1871 (N_1871,N_1572,N_1680);
xor U1872 (N_1872,N_1667,N_1735);
nand U1873 (N_1873,N_1644,N_1525);
nor U1874 (N_1874,N_1695,N_1641);
nor U1875 (N_1875,N_1709,N_1708);
xor U1876 (N_1876,N_1520,N_1510);
nand U1877 (N_1877,N_1569,N_1643);
or U1878 (N_1878,N_1702,N_1745);
nor U1879 (N_1879,N_1631,N_1655);
xnor U1880 (N_1880,N_1524,N_1647);
xor U1881 (N_1881,N_1651,N_1577);
or U1882 (N_1882,N_1731,N_1561);
nor U1883 (N_1883,N_1706,N_1703);
nand U1884 (N_1884,N_1501,N_1637);
nand U1885 (N_1885,N_1531,N_1744);
xnor U1886 (N_1886,N_1620,N_1586);
nand U1887 (N_1887,N_1525,N_1579);
nand U1888 (N_1888,N_1597,N_1560);
nand U1889 (N_1889,N_1534,N_1725);
nand U1890 (N_1890,N_1743,N_1646);
nor U1891 (N_1891,N_1562,N_1534);
or U1892 (N_1892,N_1609,N_1744);
or U1893 (N_1893,N_1623,N_1670);
and U1894 (N_1894,N_1630,N_1677);
nand U1895 (N_1895,N_1513,N_1545);
nor U1896 (N_1896,N_1637,N_1589);
and U1897 (N_1897,N_1696,N_1693);
or U1898 (N_1898,N_1720,N_1699);
nand U1899 (N_1899,N_1633,N_1714);
xnor U1900 (N_1900,N_1688,N_1585);
xnor U1901 (N_1901,N_1630,N_1594);
nand U1902 (N_1902,N_1606,N_1589);
xnor U1903 (N_1903,N_1607,N_1714);
xnor U1904 (N_1904,N_1515,N_1720);
or U1905 (N_1905,N_1590,N_1607);
nand U1906 (N_1906,N_1739,N_1721);
nor U1907 (N_1907,N_1500,N_1735);
xnor U1908 (N_1908,N_1554,N_1500);
nand U1909 (N_1909,N_1501,N_1568);
xnor U1910 (N_1910,N_1718,N_1609);
xnor U1911 (N_1911,N_1542,N_1546);
nor U1912 (N_1912,N_1664,N_1603);
or U1913 (N_1913,N_1679,N_1744);
nand U1914 (N_1914,N_1635,N_1688);
xnor U1915 (N_1915,N_1621,N_1553);
nand U1916 (N_1916,N_1605,N_1643);
nand U1917 (N_1917,N_1532,N_1652);
nor U1918 (N_1918,N_1630,N_1732);
nand U1919 (N_1919,N_1610,N_1580);
nand U1920 (N_1920,N_1613,N_1516);
and U1921 (N_1921,N_1735,N_1682);
and U1922 (N_1922,N_1650,N_1695);
xnor U1923 (N_1923,N_1545,N_1554);
nand U1924 (N_1924,N_1559,N_1644);
or U1925 (N_1925,N_1532,N_1668);
or U1926 (N_1926,N_1690,N_1669);
nand U1927 (N_1927,N_1705,N_1594);
nand U1928 (N_1928,N_1595,N_1609);
nor U1929 (N_1929,N_1562,N_1530);
and U1930 (N_1930,N_1613,N_1733);
or U1931 (N_1931,N_1679,N_1533);
or U1932 (N_1932,N_1688,N_1701);
xor U1933 (N_1933,N_1558,N_1685);
or U1934 (N_1934,N_1593,N_1540);
xor U1935 (N_1935,N_1620,N_1642);
or U1936 (N_1936,N_1740,N_1561);
or U1937 (N_1937,N_1710,N_1655);
nand U1938 (N_1938,N_1637,N_1584);
nand U1939 (N_1939,N_1551,N_1565);
or U1940 (N_1940,N_1552,N_1725);
nand U1941 (N_1941,N_1680,N_1595);
or U1942 (N_1942,N_1580,N_1677);
nor U1943 (N_1943,N_1597,N_1735);
or U1944 (N_1944,N_1572,N_1726);
xnor U1945 (N_1945,N_1645,N_1592);
nor U1946 (N_1946,N_1680,N_1594);
nand U1947 (N_1947,N_1691,N_1575);
nor U1948 (N_1948,N_1636,N_1598);
nor U1949 (N_1949,N_1719,N_1695);
xnor U1950 (N_1950,N_1643,N_1665);
or U1951 (N_1951,N_1713,N_1697);
and U1952 (N_1952,N_1675,N_1724);
nor U1953 (N_1953,N_1721,N_1579);
or U1954 (N_1954,N_1646,N_1732);
and U1955 (N_1955,N_1738,N_1555);
or U1956 (N_1956,N_1605,N_1633);
nand U1957 (N_1957,N_1645,N_1619);
nor U1958 (N_1958,N_1612,N_1670);
or U1959 (N_1959,N_1633,N_1621);
nand U1960 (N_1960,N_1719,N_1743);
nor U1961 (N_1961,N_1615,N_1660);
and U1962 (N_1962,N_1555,N_1634);
or U1963 (N_1963,N_1584,N_1517);
and U1964 (N_1964,N_1619,N_1739);
or U1965 (N_1965,N_1720,N_1670);
or U1966 (N_1966,N_1708,N_1587);
nor U1967 (N_1967,N_1675,N_1615);
nand U1968 (N_1968,N_1550,N_1534);
nor U1969 (N_1969,N_1749,N_1602);
or U1970 (N_1970,N_1590,N_1683);
or U1971 (N_1971,N_1745,N_1602);
and U1972 (N_1972,N_1683,N_1665);
nor U1973 (N_1973,N_1658,N_1618);
nand U1974 (N_1974,N_1615,N_1642);
xor U1975 (N_1975,N_1511,N_1508);
nor U1976 (N_1976,N_1620,N_1693);
nor U1977 (N_1977,N_1565,N_1558);
nand U1978 (N_1978,N_1545,N_1666);
nand U1979 (N_1979,N_1747,N_1672);
or U1980 (N_1980,N_1735,N_1700);
or U1981 (N_1981,N_1610,N_1516);
or U1982 (N_1982,N_1598,N_1647);
xnor U1983 (N_1983,N_1608,N_1526);
nor U1984 (N_1984,N_1602,N_1537);
nor U1985 (N_1985,N_1599,N_1507);
or U1986 (N_1986,N_1667,N_1540);
nor U1987 (N_1987,N_1548,N_1512);
nor U1988 (N_1988,N_1747,N_1575);
xnor U1989 (N_1989,N_1504,N_1573);
nand U1990 (N_1990,N_1643,N_1593);
or U1991 (N_1991,N_1556,N_1582);
or U1992 (N_1992,N_1536,N_1640);
and U1993 (N_1993,N_1576,N_1708);
nor U1994 (N_1994,N_1538,N_1542);
nand U1995 (N_1995,N_1694,N_1523);
and U1996 (N_1996,N_1568,N_1634);
nor U1997 (N_1997,N_1593,N_1648);
nor U1998 (N_1998,N_1735,N_1702);
and U1999 (N_1999,N_1570,N_1637);
nor U2000 (N_2000,N_1951,N_1800);
nor U2001 (N_2001,N_1910,N_1887);
nand U2002 (N_2002,N_1945,N_1790);
nand U2003 (N_2003,N_1834,N_1863);
or U2004 (N_2004,N_1971,N_1832);
and U2005 (N_2005,N_1801,N_1983);
or U2006 (N_2006,N_1860,N_1818);
xor U2007 (N_2007,N_1908,N_1862);
or U2008 (N_2008,N_1967,N_1905);
or U2009 (N_2009,N_1822,N_1962);
xor U2010 (N_2010,N_1859,N_1872);
xor U2011 (N_2011,N_1789,N_1806);
or U2012 (N_2012,N_1886,N_1949);
nor U2013 (N_2013,N_1935,N_1838);
nor U2014 (N_2014,N_1825,N_1830);
nor U2015 (N_2015,N_1885,N_1954);
xnor U2016 (N_2016,N_1869,N_1900);
nor U2017 (N_2017,N_1952,N_1810);
nor U2018 (N_2018,N_1858,N_1928);
and U2019 (N_2019,N_1996,N_1940);
and U2020 (N_2020,N_1955,N_1839);
or U2021 (N_2021,N_1836,N_1811);
xnor U2022 (N_2022,N_1965,N_1751);
xnor U2023 (N_2023,N_1849,N_1823);
and U2024 (N_2024,N_1929,N_1914);
or U2025 (N_2025,N_1754,N_1911);
nor U2026 (N_2026,N_1817,N_1840);
and U2027 (N_2027,N_1968,N_1786);
nand U2028 (N_2028,N_1852,N_1969);
or U2029 (N_2029,N_1960,N_1813);
xor U2030 (N_2030,N_1854,N_1927);
or U2031 (N_2031,N_1936,N_1847);
or U2032 (N_2032,N_1979,N_1775);
nor U2033 (N_2033,N_1850,N_1913);
nand U2034 (N_2034,N_1959,N_1763);
nand U2035 (N_2035,N_1779,N_1774);
nand U2036 (N_2036,N_1805,N_1851);
and U2037 (N_2037,N_1844,N_1938);
nand U2038 (N_2038,N_1988,N_1808);
nand U2039 (N_2039,N_1899,N_1815);
nand U2040 (N_2040,N_1941,N_1989);
xnor U2041 (N_2041,N_1820,N_1895);
xor U2042 (N_2042,N_1835,N_1921);
nand U2043 (N_2043,N_1843,N_1865);
or U2044 (N_2044,N_1819,N_1776);
xnor U2045 (N_2045,N_1963,N_1981);
xnor U2046 (N_2046,N_1904,N_1975);
nor U2047 (N_2047,N_1829,N_1757);
nand U2048 (N_2048,N_1897,N_1966);
nor U2049 (N_2049,N_1809,N_1853);
xnor U2050 (N_2050,N_1957,N_1958);
xor U2051 (N_2051,N_1974,N_1842);
and U2052 (N_2052,N_1793,N_1920);
or U2053 (N_2053,N_1791,N_1993);
and U2054 (N_2054,N_1856,N_1934);
xnor U2055 (N_2055,N_1784,N_1752);
xnor U2056 (N_2056,N_1907,N_1942);
or U2057 (N_2057,N_1964,N_1803);
and U2058 (N_2058,N_1773,N_1902);
nor U2059 (N_2059,N_1777,N_1990);
and U2060 (N_2060,N_1939,N_1937);
nand U2061 (N_2061,N_1956,N_1798);
nor U2062 (N_2062,N_1876,N_1785);
xor U2063 (N_2063,N_1980,N_1778);
xnor U2064 (N_2064,N_1892,N_1873);
xnor U2065 (N_2065,N_1894,N_1781);
and U2066 (N_2066,N_1901,N_1946);
and U2067 (N_2067,N_1909,N_1917);
nand U2068 (N_2068,N_1769,N_1992);
nand U2069 (N_2069,N_1864,N_1787);
nor U2070 (N_2070,N_1976,N_1759);
and U2071 (N_2071,N_1932,N_1953);
or U2072 (N_2072,N_1877,N_1881);
and U2073 (N_2073,N_1889,N_1772);
nand U2074 (N_2074,N_1994,N_1797);
or U2075 (N_2075,N_1987,N_1995);
or U2076 (N_2076,N_1788,N_1771);
nor U2077 (N_2077,N_1896,N_1978);
nor U2078 (N_2078,N_1767,N_1879);
nand U2079 (N_2079,N_1926,N_1875);
or U2080 (N_2080,N_1756,N_1985);
nor U2081 (N_2081,N_1977,N_1828);
or U2082 (N_2082,N_1972,N_1874);
nand U2083 (N_2083,N_1750,N_1986);
and U2084 (N_2084,N_1821,N_1761);
xnor U2085 (N_2085,N_1944,N_1826);
xor U2086 (N_2086,N_1916,N_1884);
nand U2087 (N_2087,N_1984,N_1794);
nor U2088 (N_2088,N_1883,N_1912);
or U2089 (N_2089,N_1861,N_1882);
nor U2090 (N_2090,N_1868,N_1857);
xnor U2091 (N_2091,N_1991,N_1925);
and U2092 (N_2092,N_1766,N_1947);
nand U2093 (N_2093,N_1802,N_1845);
nand U2094 (N_2094,N_1970,N_1933);
and U2095 (N_2095,N_1762,N_1755);
nand U2096 (N_2096,N_1918,N_1837);
nand U2097 (N_2097,N_1783,N_1931);
and U2098 (N_2098,N_1915,N_1782);
xor U2099 (N_2099,N_1824,N_1870);
or U2100 (N_2100,N_1888,N_1982);
or U2101 (N_2101,N_1796,N_1799);
and U2102 (N_2102,N_1961,N_1760);
or U2103 (N_2103,N_1841,N_1922);
nor U2104 (N_2104,N_1878,N_1753);
nor U2105 (N_2105,N_1846,N_1923);
nor U2106 (N_2106,N_1930,N_1866);
and U2107 (N_2107,N_1999,N_1997);
xor U2108 (N_2108,N_1848,N_1867);
nor U2109 (N_2109,N_1924,N_1973);
and U2110 (N_2110,N_1795,N_1758);
or U2111 (N_2111,N_1807,N_1770);
and U2112 (N_2112,N_1816,N_1871);
or U2113 (N_2113,N_1943,N_1919);
or U2114 (N_2114,N_1890,N_1898);
and U2115 (N_2115,N_1814,N_1792);
nor U2116 (N_2116,N_1764,N_1891);
or U2117 (N_2117,N_1893,N_1831);
xnor U2118 (N_2118,N_1998,N_1903);
nand U2119 (N_2119,N_1948,N_1765);
xnor U2120 (N_2120,N_1827,N_1833);
or U2121 (N_2121,N_1950,N_1768);
nor U2122 (N_2122,N_1804,N_1906);
or U2123 (N_2123,N_1780,N_1812);
xnor U2124 (N_2124,N_1880,N_1855);
xor U2125 (N_2125,N_1862,N_1930);
and U2126 (N_2126,N_1957,N_1841);
or U2127 (N_2127,N_1907,N_1806);
or U2128 (N_2128,N_1785,N_1945);
or U2129 (N_2129,N_1874,N_1938);
or U2130 (N_2130,N_1885,N_1872);
nand U2131 (N_2131,N_1833,N_1798);
or U2132 (N_2132,N_1960,N_1789);
and U2133 (N_2133,N_1803,N_1860);
nor U2134 (N_2134,N_1786,N_1908);
xor U2135 (N_2135,N_1762,N_1992);
xor U2136 (N_2136,N_1775,N_1760);
and U2137 (N_2137,N_1841,N_1851);
or U2138 (N_2138,N_1810,N_1804);
xor U2139 (N_2139,N_1976,N_1879);
or U2140 (N_2140,N_1790,N_1865);
xnor U2141 (N_2141,N_1811,N_1772);
xnor U2142 (N_2142,N_1989,N_1831);
and U2143 (N_2143,N_1837,N_1916);
nor U2144 (N_2144,N_1785,N_1925);
nor U2145 (N_2145,N_1815,N_1905);
nor U2146 (N_2146,N_1958,N_1798);
nor U2147 (N_2147,N_1868,N_1836);
and U2148 (N_2148,N_1917,N_1801);
nor U2149 (N_2149,N_1795,N_1847);
nor U2150 (N_2150,N_1879,N_1924);
xnor U2151 (N_2151,N_1757,N_1918);
xnor U2152 (N_2152,N_1829,N_1975);
xor U2153 (N_2153,N_1855,N_1982);
nor U2154 (N_2154,N_1847,N_1801);
nand U2155 (N_2155,N_1824,N_1780);
xor U2156 (N_2156,N_1926,N_1974);
and U2157 (N_2157,N_1983,N_1750);
and U2158 (N_2158,N_1872,N_1989);
nor U2159 (N_2159,N_1838,N_1934);
nor U2160 (N_2160,N_1976,N_1849);
nor U2161 (N_2161,N_1905,N_1839);
and U2162 (N_2162,N_1891,N_1953);
nand U2163 (N_2163,N_1862,N_1937);
or U2164 (N_2164,N_1754,N_1873);
nand U2165 (N_2165,N_1995,N_1979);
and U2166 (N_2166,N_1895,N_1936);
xnor U2167 (N_2167,N_1997,N_1821);
xor U2168 (N_2168,N_1978,N_1975);
or U2169 (N_2169,N_1909,N_1943);
nor U2170 (N_2170,N_1902,N_1889);
nor U2171 (N_2171,N_1870,N_1971);
nand U2172 (N_2172,N_1808,N_1792);
or U2173 (N_2173,N_1865,N_1825);
nor U2174 (N_2174,N_1758,N_1965);
nand U2175 (N_2175,N_1797,N_1897);
nand U2176 (N_2176,N_1915,N_1997);
nand U2177 (N_2177,N_1877,N_1814);
or U2178 (N_2178,N_1867,N_1833);
xor U2179 (N_2179,N_1823,N_1998);
nor U2180 (N_2180,N_1960,N_1875);
nand U2181 (N_2181,N_1866,N_1814);
or U2182 (N_2182,N_1804,N_1923);
and U2183 (N_2183,N_1769,N_1823);
nand U2184 (N_2184,N_1928,N_1832);
and U2185 (N_2185,N_1877,N_1764);
xor U2186 (N_2186,N_1816,N_1821);
or U2187 (N_2187,N_1975,N_1819);
nand U2188 (N_2188,N_1839,N_1819);
and U2189 (N_2189,N_1803,N_1829);
xnor U2190 (N_2190,N_1776,N_1906);
nor U2191 (N_2191,N_1899,N_1801);
xor U2192 (N_2192,N_1969,N_1976);
nand U2193 (N_2193,N_1823,N_1937);
and U2194 (N_2194,N_1950,N_1827);
xor U2195 (N_2195,N_1935,N_1912);
or U2196 (N_2196,N_1807,N_1870);
or U2197 (N_2197,N_1804,N_1929);
xor U2198 (N_2198,N_1983,N_1810);
or U2199 (N_2199,N_1928,N_1763);
nor U2200 (N_2200,N_1810,N_1980);
nand U2201 (N_2201,N_1840,N_1940);
xnor U2202 (N_2202,N_1796,N_1912);
nor U2203 (N_2203,N_1787,N_1849);
xor U2204 (N_2204,N_1879,N_1913);
xor U2205 (N_2205,N_1788,N_1810);
xor U2206 (N_2206,N_1782,N_1847);
or U2207 (N_2207,N_1908,N_1890);
xnor U2208 (N_2208,N_1989,N_1877);
nand U2209 (N_2209,N_1911,N_1833);
nor U2210 (N_2210,N_1953,N_1851);
nand U2211 (N_2211,N_1754,N_1792);
and U2212 (N_2212,N_1968,N_1854);
nor U2213 (N_2213,N_1854,N_1837);
nand U2214 (N_2214,N_1841,N_1949);
xor U2215 (N_2215,N_1797,N_1855);
nor U2216 (N_2216,N_1772,N_1809);
nor U2217 (N_2217,N_1757,N_1824);
nand U2218 (N_2218,N_1790,N_1892);
or U2219 (N_2219,N_1951,N_1818);
and U2220 (N_2220,N_1767,N_1806);
nor U2221 (N_2221,N_1755,N_1883);
or U2222 (N_2222,N_1995,N_1834);
nand U2223 (N_2223,N_1970,N_1963);
xor U2224 (N_2224,N_1971,N_1799);
and U2225 (N_2225,N_1973,N_1916);
xor U2226 (N_2226,N_1869,N_1882);
nand U2227 (N_2227,N_1985,N_1940);
or U2228 (N_2228,N_1850,N_1967);
nand U2229 (N_2229,N_1959,N_1869);
and U2230 (N_2230,N_1930,N_1944);
nand U2231 (N_2231,N_1858,N_1809);
and U2232 (N_2232,N_1824,N_1809);
xnor U2233 (N_2233,N_1760,N_1997);
xor U2234 (N_2234,N_1824,N_1947);
or U2235 (N_2235,N_1801,N_1819);
or U2236 (N_2236,N_1916,N_1819);
nand U2237 (N_2237,N_1878,N_1861);
nor U2238 (N_2238,N_1977,N_1998);
nor U2239 (N_2239,N_1768,N_1988);
and U2240 (N_2240,N_1902,N_1948);
and U2241 (N_2241,N_1766,N_1914);
nor U2242 (N_2242,N_1828,N_1766);
nor U2243 (N_2243,N_1767,N_1952);
or U2244 (N_2244,N_1779,N_1796);
nor U2245 (N_2245,N_1794,N_1951);
nand U2246 (N_2246,N_1792,N_1930);
or U2247 (N_2247,N_1956,N_1936);
nor U2248 (N_2248,N_1776,N_1817);
or U2249 (N_2249,N_1916,N_1928);
or U2250 (N_2250,N_2079,N_2071);
and U2251 (N_2251,N_2223,N_2149);
and U2252 (N_2252,N_2221,N_2207);
and U2253 (N_2253,N_2039,N_2067);
or U2254 (N_2254,N_2162,N_2174);
nand U2255 (N_2255,N_2157,N_2072);
xnor U2256 (N_2256,N_2141,N_2108);
nor U2257 (N_2257,N_2089,N_2109);
and U2258 (N_2258,N_2004,N_2211);
xor U2259 (N_2259,N_2025,N_2020);
nor U2260 (N_2260,N_2138,N_2115);
nand U2261 (N_2261,N_2200,N_2126);
nand U2262 (N_2262,N_2027,N_2076);
and U2263 (N_2263,N_2229,N_2209);
nor U2264 (N_2264,N_2058,N_2159);
nor U2265 (N_2265,N_2180,N_2172);
nand U2266 (N_2266,N_2236,N_2217);
nand U2267 (N_2267,N_2206,N_2069);
nor U2268 (N_2268,N_2068,N_2083);
or U2269 (N_2269,N_2199,N_2167);
and U2270 (N_2270,N_2234,N_2015);
or U2271 (N_2271,N_2054,N_2008);
and U2272 (N_2272,N_2118,N_2010);
nand U2273 (N_2273,N_2124,N_2210);
and U2274 (N_2274,N_2001,N_2006);
and U2275 (N_2275,N_2034,N_2193);
and U2276 (N_2276,N_2014,N_2232);
xnor U2277 (N_2277,N_2030,N_2235);
nor U2278 (N_2278,N_2100,N_2048);
nand U2279 (N_2279,N_2065,N_2133);
nor U2280 (N_2280,N_2037,N_2135);
nor U2281 (N_2281,N_2191,N_2005);
xnor U2282 (N_2282,N_2085,N_2201);
and U2283 (N_2283,N_2213,N_2044);
and U2284 (N_2284,N_2168,N_2063);
and U2285 (N_2285,N_2050,N_2190);
nand U2286 (N_2286,N_2074,N_2224);
xor U2287 (N_2287,N_2032,N_2024);
and U2288 (N_2288,N_2097,N_2233);
xnor U2289 (N_2289,N_2040,N_2158);
xnor U2290 (N_2290,N_2123,N_2111);
and U2291 (N_2291,N_2002,N_2171);
nor U2292 (N_2292,N_2066,N_2205);
nand U2293 (N_2293,N_2018,N_2077);
xor U2294 (N_2294,N_2237,N_2246);
or U2295 (N_2295,N_2227,N_2219);
nor U2296 (N_2296,N_2196,N_2122);
nor U2297 (N_2297,N_2041,N_2120);
and U2298 (N_2298,N_2183,N_2086);
nor U2299 (N_2299,N_2084,N_2218);
and U2300 (N_2300,N_2243,N_2075);
nand U2301 (N_2301,N_2179,N_2178);
nand U2302 (N_2302,N_2105,N_2245);
nor U2303 (N_2303,N_2240,N_2078);
or U2304 (N_2304,N_2038,N_2012);
xor U2305 (N_2305,N_2082,N_2177);
or U2306 (N_2306,N_2103,N_2112);
and U2307 (N_2307,N_2194,N_2017);
or U2308 (N_2308,N_2139,N_2182);
or U2309 (N_2309,N_2137,N_2101);
xnor U2310 (N_2310,N_2053,N_2073);
nand U2311 (N_2311,N_2049,N_2204);
nor U2312 (N_2312,N_2147,N_2247);
xnor U2313 (N_2313,N_2092,N_2175);
nor U2314 (N_2314,N_2152,N_2029);
and U2315 (N_2315,N_2131,N_2031);
or U2316 (N_2316,N_2143,N_2114);
nor U2317 (N_2317,N_2125,N_2203);
nand U2318 (N_2318,N_2028,N_2148);
xor U2319 (N_2319,N_2136,N_2062);
and U2320 (N_2320,N_2104,N_2144);
xnor U2321 (N_2321,N_2127,N_2156);
nor U2322 (N_2322,N_2192,N_2061);
nand U2323 (N_2323,N_2214,N_2176);
xor U2324 (N_2324,N_2093,N_2166);
or U2325 (N_2325,N_2216,N_2153);
and U2326 (N_2326,N_2225,N_2164);
and U2327 (N_2327,N_2116,N_2188);
nand U2328 (N_2328,N_2021,N_2249);
nand U2329 (N_2329,N_2099,N_2026);
nor U2330 (N_2330,N_2181,N_2119);
nor U2331 (N_2331,N_2134,N_2186);
and U2332 (N_2332,N_2107,N_2242);
and U2333 (N_2333,N_2239,N_2163);
and U2334 (N_2334,N_2052,N_2110);
and U2335 (N_2335,N_2132,N_2060);
nand U2336 (N_2336,N_2244,N_2189);
nand U2337 (N_2337,N_2238,N_2043);
nand U2338 (N_2338,N_2051,N_2230);
or U2339 (N_2339,N_2212,N_2173);
and U2340 (N_2340,N_2187,N_2091);
or U2341 (N_2341,N_2011,N_2220);
nand U2342 (N_2342,N_2113,N_2129);
nand U2343 (N_2343,N_2121,N_2198);
nor U2344 (N_2344,N_2140,N_2184);
nor U2345 (N_2345,N_2007,N_2161);
or U2346 (N_2346,N_2036,N_2208);
xor U2347 (N_2347,N_2064,N_2056);
nand U2348 (N_2348,N_2095,N_2185);
and U2349 (N_2349,N_2098,N_2009);
and U2350 (N_2350,N_2096,N_2013);
and U2351 (N_2351,N_2117,N_2146);
or U2352 (N_2352,N_2154,N_2150);
nor U2353 (N_2353,N_2046,N_2022);
xnor U2354 (N_2354,N_2228,N_2165);
and U2355 (N_2355,N_2033,N_2195);
nor U2356 (N_2356,N_2130,N_2106);
nor U2357 (N_2357,N_2045,N_2016);
nand U2358 (N_2358,N_2019,N_2197);
and U2359 (N_2359,N_2248,N_2087);
xor U2360 (N_2360,N_2151,N_2215);
and U2361 (N_2361,N_2102,N_2070);
nor U2362 (N_2362,N_2142,N_2080);
xnor U2363 (N_2363,N_2090,N_2169);
xnor U2364 (N_2364,N_2145,N_2088);
and U2365 (N_2365,N_2055,N_2241);
nor U2366 (N_2366,N_2081,N_2042);
nor U2367 (N_2367,N_2000,N_2094);
nor U2368 (N_2368,N_2057,N_2059);
xor U2369 (N_2369,N_2170,N_2035);
and U2370 (N_2370,N_2155,N_2128);
xnor U2371 (N_2371,N_2003,N_2047);
nand U2372 (N_2372,N_2226,N_2160);
and U2373 (N_2373,N_2222,N_2023);
nand U2374 (N_2374,N_2202,N_2231);
nor U2375 (N_2375,N_2044,N_2175);
and U2376 (N_2376,N_2164,N_2204);
or U2377 (N_2377,N_2092,N_2054);
and U2378 (N_2378,N_2081,N_2125);
and U2379 (N_2379,N_2043,N_2009);
or U2380 (N_2380,N_2187,N_2238);
nand U2381 (N_2381,N_2136,N_2238);
and U2382 (N_2382,N_2127,N_2169);
nor U2383 (N_2383,N_2159,N_2047);
nand U2384 (N_2384,N_2147,N_2005);
nor U2385 (N_2385,N_2052,N_2199);
or U2386 (N_2386,N_2246,N_2182);
or U2387 (N_2387,N_2224,N_2176);
xor U2388 (N_2388,N_2100,N_2147);
xnor U2389 (N_2389,N_2197,N_2113);
xor U2390 (N_2390,N_2142,N_2123);
nor U2391 (N_2391,N_2229,N_2081);
nand U2392 (N_2392,N_2041,N_2204);
or U2393 (N_2393,N_2144,N_2221);
and U2394 (N_2394,N_2117,N_2089);
nor U2395 (N_2395,N_2159,N_2064);
nand U2396 (N_2396,N_2161,N_2090);
xnor U2397 (N_2397,N_2118,N_2207);
and U2398 (N_2398,N_2107,N_2223);
xnor U2399 (N_2399,N_2067,N_2026);
nor U2400 (N_2400,N_2136,N_2109);
and U2401 (N_2401,N_2233,N_2108);
and U2402 (N_2402,N_2205,N_2001);
nand U2403 (N_2403,N_2171,N_2243);
and U2404 (N_2404,N_2119,N_2040);
xnor U2405 (N_2405,N_2249,N_2119);
nand U2406 (N_2406,N_2149,N_2063);
nand U2407 (N_2407,N_2217,N_2149);
nor U2408 (N_2408,N_2016,N_2046);
or U2409 (N_2409,N_2059,N_2121);
or U2410 (N_2410,N_2056,N_2016);
nand U2411 (N_2411,N_2086,N_2126);
xnor U2412 (N_2412,N_2196,N_2203);
nor U2413 (N_2413,N_2027,N_2216);
nand U2414 (N_2414,N_2053,N_2249);
and U2415 (N_2415,N_2013,N_2234);
xnor U2416 (N_2416,N_2226,N_2052);
and U2417 (N_2417,N_2082,N_2156);
nand U2418 (N_2418,N_2139,N_2243);
nor U2419 (N_2419,N_2157,N_2124);
nand U2420 (N_2420,N_2007,N_2086);
nor U2421 (N_2421,N_2090,N_2002);
nand U2422 (N_2422,N_2123,N_2116);
nand U2423 (N_2423,N_2060,N_2101);
or U2424 (N_2424,N_2174,N_2088);
and U2425 (N_2425,N_2172,N_2078);
nand U2426 (N_2426,N_2142,N_2084);
or U2427 (N_2427,N_2122,N_2202);
nor U2428 (N_2428,N_2066,N_2225);
or U2429 (N_2429,N_2192,N_2245);
xnor U2430 (N_2430,N_2131,N_2220);
and U2431 (N_2431,N_2125,N_2065);
or U2432 (N_2432,N_2116,N_2173);
or U2433 (N_2433,N_2016,N_2163);
or U2434 (N_2434,N_2165,N_2017);
and U2435 (N_2435,N_2119,N_2172);
nor U2436 (N_2436,N_2112,N_2201);
and U2437 (N_2437,N_2110,N_2139);
nor U2438 (N_2438,N_2124,N_2027);
or U2439 (N_2439,N_2056,N_2086);
and U2440 (N_2440,N_2007,N_2192);
nor U2441 (N_2441,N_2058,N_2124);
xor U2442 (N_2442,N_2068,N_2215);
or U2443 (N_2443,N_2080,N_2037);
and U2444 (N_2444,N_2093,N_2120);
nor U2445 (N_2445,N_2107,N_2221);
nor U2446 (N_2446,N_2096,N_2048);
and U2447 (N_2447,N_2049,N_2030);
nor U2448 (N_2448,N_2022,N_2111);
nor U2449 (N_2449,N_2186,N_2160);
nor U2450 (N_2450,N_2048,N_2042);
nand U2451 (N_2451,N_2100,N_2145);
xnor U2452 (N_2452,N_2095,N_2043);
nand U2453 (N_2453,N_2125,N_2160);
nor U2454 (N_2454,N_2112,N_2144);
xnor U2455 (N_2455,N_2102,N_2227);
nor U2456 (N_2456,N_2172,N_2152);
xnor U2457 (N_2457,N_2178,N_2111);
or U2458 (N_2458,N_2212,N_2162);
and U2459 (N_2459,N_2062,N_2187);
and U2460 (N_2460,N_2096,N_2046);
nor U2461 (N_2461,N_2162,N_2223);
xnor U2462 (N_2462,N_2214,N_2188);
nand U2463 (N_2463,N_2080,N_2093);
or U2464 (N_2464,N_2155,N_2037);
xor U2465 (N_2465,N_2141,N_2197);
or U2466 (N_2466,N_2239,N_2107);
xnor U2467 (N_2467,N_2172,N_2165);
nand U2468 (N_2468,N_2235,N_2139);
xor U2469 (N_2469,N_2185,N_2104);
nand U2470 (N_2470,N_2120,N_2238);
and U2471 (N_2471,N_2218,N_2040);
and U2472 (N_2472,N_2100,N_2125);
nor U2473 (N_2473,N_2050,N_2162);
or U2474 (N_2474,N_2181,N_2245);
nor U2475 (N_2475,N_2066,N_2112);
nand U2476 (N_2476,N_2058,N_2099);
xnor U2477 (N_2477,N_2249,N_2098);
xor U2478 (N_2478,N_2213,N_2032);
nor U2479 (N_2479,N_2083,N_2247);
nor U2480 (N_2480,N_2169,N_2094);
or U2481 (N_2481,N_2110,N_2121);
nand U2482 (N_2482,N_2208,N_2092);
or U2483 (N_2483,N_2057,N_2011);
nor U2484 (N_2484,N_2151,N_2226);
nor U2485 (N_2485,N_2186,N_2081);
and U2486 (N_2486,N_2085,N_2210);
xnor U2487 (N_2487,N_2118,N_2003);
xor U2488 (N_2488,N_2239,N_2198);
or U2489 (N_2489,N_2039,N_2004);
nor U2490 (N_2490,N_2132,N_2194);
and U2491 (N_2491,N_2108,N_2230);
or U2492 (N_2492,N_2104,N_2062);
xor U2493 (N_2493,N_2119,N_2237);
or U2494 (N_2494,N_2127,N_2008);
nand U2495 (N_2495,N_2117,N_2208);
and U2496 (N_2496,N_2018,N_2175);
xnor U2497 (N_2497,N_2030,N_2087);
or U2498 (N_2498,N_2053,N_2013);
nor U2499 (N_2499,N_2022,N_2173);
nor U2500 (N_2500,N_2460,N_2422);
xor U2501 (N_2501,N_2350,N_2409);
nor U2502 (N_2502,N_2353,N_2465);
and U2503 (N_2503,N_2297,N_2450);
xor U2504 (N_2504,N_2440,N_2300);
nor U2505 (N_2505,N_2340,N_2462);
and U2506 (N_2506,N_2360,N_2301);
xnor U2507 (N_2507,N_2310,N_2278);
and U2508 (N_2508,N_2293,N_2386);
or U2509 (N_2509,N_2378,N_2364);
and U2510 (N_2510,N_2493,N_2388);
nand U2511 (N_2511,N_2483,N_2427);
or U2512 (N_2512,N_2257,N_2289);
and U2513 (N_2513,N_2255,N_2403);
nand U2514 (N_2514,N_2410,N_2327);
nand U2515 (N_2515,N_2441,N_2391);
nand U2516 (N_2516,N_2251,N_2338);
or U2517 (N_2517,N_2472,N_2296);
nand U2518 (N_2518,N_2426,N_2343);
nand U2519 (N_2519,N_2497,N_2254);
and U2520 (N_2520,N_2405,N_2298);
and U2521 (N_2521,N_2366,N_2412);
xnor U2522 (N_2522,N_2288,N_2341);
nand U2523 (N_2523,N_2373,N_2307);
or U2524 (N_2524,N_2276,N_2316);
and U2525 (N_2525,N_2397,N_2357);
nor U2526 (N_2526,N_2362,N_2287);
and U2527 (N_2527,N_2491,N_2279);
nor U2528 (N_2528,N_2286,N_2385);
and U2529 (N_2529,N_2349,N_2262);
nor U2530 (N_2530,N_2393,N_2354);
xor U2531 (N_2531,N_2376,N_2281);
xnor U2532 (N_2532,N_2265,N_2344);
xor U2533 (N_2533,N_2408,N_2299);
nand U2534 (N_2534,N_2335,N_2291);
nor U2535 (N_2535,N_2496,N_2459);
and U2536 (N_2536,N_2448,N_2458);
xor U2537 (N_2537,N_2481,N_2345);
and U2538 (N_2538,N_2277,N_2361);
and U2539 (N_2539,N_2404,N_2271);
or U2540 (N_2540,N_2417,N_2489);
xnor U2541 (N_2541,N_2444,N_2267);
nand U2542 (N_2542,N_2419,N_2273);
nor U2543 (N_2543,N_2348,N_2428);
and U2544 (N_2544,N_2321,N_2442);
nand U2545 (N_2545,N_2443,N_2423);
or U2546 (N_2546,N_2379,N_2309);
xor U2547 (N_2547,N_2250,N_2326);
xor U2548 (N_2548,N_2433,N_2424);
nand U2549 (N_2549,N_2467,N_2274);
xor U2550 (N_2550,N_2461,N_2306);
xnor U2551 (N_2551,N_2328,N_2375);
or U2552 (N_2552,N_2434,N_2383);
nor U2553 (N_2553,N_2372,N_2312);
nor U2554 (N_2554,N_2454,N_2401);
or U2555 (N_2555,N_2320,N_2333);
and U2556 (N_2556,N_2394,N_2272);
and U2557 (N_2557,N_2305,N_2499);
and U2558 (N_2558,N_2421,N_2471);
xor U2559 (N_2559,N_2359,N_2449);
nand U2560 (N_2560,N_2407,N_2494);
nand U2561 (N_2561,N_2304,N_2399);
nand U2562 (N_2562,N_2352,N_2395);
nor U2563 (N_2563,N_2445,N_2464);
nor U2564 (N_2564,N_2392,N_2264);
or U2565 (N_2565,N_2363,N_2325);
nor U2566 (N_2566,N_2389,N_2406);
nand U2567 (N_2567,N_2377,N_2457);
nand U2568 (N_2568,N_2371,N_2477);
xnor U2569 (N_2569,N_2336,N_2480);
nor U2570 (N_2570,N_2329,N_2285);
or U2571 (N_2571,N_2475,N_2263);
and U2572 (N_2572,N_2490,N_2339);
nand U2573 (N_2573,N_2319,N_2484);
and U2574 (N_2574,N_2318,N_2252);
or U2575 (N_2575,N_2351,N_2469);
and U2576 (N_2576,N_2369,N_2429);
and U2577 (N_2577,N_2314,N_2294);
nor U2578 (N_2578,N_2368,N_2398);
xor U2579 (N_2579,N_2258,N_2436);
nand U2580 (N_2580,N_2413,N_2492);
xor U2581 (N_2581,N_2446,N_2414);
nor U2582 (N_2582,N_2400,N_2367);
xor U2583 (N_2583,N_2468,N_2275);
or U2584 (N_2584,N_2487,N_2485);
xor U2585 (N_2585,N_2290,N_2380);
and U2586 (N_2586,N_2420,N_2315);
xnor U2587 (N_2587,N_2259,N_2456);
nor U2588 (N_2588,N_2280,N_2313);
nor U2589 (N_2589,N_2431,N_2466);
or U2590 (N_2590,N_2358,N_2455);
nand U2591 (N_2591,N_2430,N_2283);
nand U2592 (N_2592,N_2476,N_2253);
or U2593 (N_2593,N_2473,N_2303);
nor U2594 (N_2594,N_2346,N_2308);
xnor U2595 (N_2595,N_2268,N_2384);
nand U2596 (N_2596,N_2432,N_2387);
or U2597 (N_2597,N_2261,N_2330);
nand U2598 (N_2598,N_2411,N_2334);
xnor U2599 (N_2599,N_2415,N_2292);
nand U2600 (N_2600,N_2317,N_2322);
and U2601 (N_2601,N_2470,N_2365);
and U2602 (N_2602,N_2266,N_2295);
or U2603 (N_2603,N_2382,N_2324);
or U2604 (N_2604,N_2374,N_2495);
xnor U2605 (N_2605,N_2337,N_2355);
nor U2606 (N_2606,N_2381,N_2435);
and U2607 (N_2607,N_2282,N_2451);
xor U2608 (N_2608,N_2270,N_2486);
xor U2609 (N_2609,N_2463,N_2474);
nor U2610 (N_2610,N_2478,N_2347);
and U2611 (N_2611,N_2439,N_2302);
xor U2612 (N_2612,N_2331,N_2453);
nand U2613 (N_2613,N_2256,N_2356);
or U2614 (N_2614,N_2482,N_2447);
nand U2615 (N_2615,N_2416,N_2370);
and U2616 (N_2616,N_2396,N_2498);
xor U2617 (N_2617,N_2260,N_2311);
and U2618 (N_2618,N_2452,N_2323);
and U2619 (N_2619,N_2390,N_2269);
nand U2620 (N_2620,N_2418,N_2332);
or U2621 (N_2621,N_2402,N_2479);
nand U2622 (N_2622,N_2438,N_2425);
xnor U2623 (N_2623,N_2437,N_2488);
and U2624 (N_2624,N_2284,N_2342);
nand U2625 (N_2625,N_2397,N_2464);
nand U2626 (N_2626,N_2369,N_2413);
nor U2627 (N_2627,N_2335,N_2430);
nor U2628 (N_2628,N_2437,N_2280);
nand U2629 (N_2629,N_2408,N_2478);
or U2630 (N_2630,N_2498,N_2460);
and U2631 (N_2631,N_2371,N_2466);
nor U2632 (N_2632,N_2287,N_2256);
or U2633 (N_2633,N_2490,N_2320);
nor U2634 (N_2634,N_2261,N_2353);
or U2635 (N_2635,N_2259,N_2271);
or U2636 (N_2636,N_2329,N_2343);
or U2637 (N_2637,N_2338,N_2323);
xor U2638 (N_2638,N_2340,N_2255);
and U2639 (N_2639,N_2407,N_2295);
xnor U2640 (N_2640,N_2481,N_2341);
and U2641 (N_2641,N_2404,N_2372);
nor U2642 (N_2642,N_2273,N_2378);
nand U2643 (N_2643,N_2439,N_2301);
and U2644 (N_2644,N_2421,N_2374);
nand U2645 (N_2645,N_2412,N_2443);
xor U2646 (N_2646,N_2386,N_2332);
nand U2647 (N_2647,N_2297,N_2434);
and U2648 (N_2648,N_2457,N_2460);
nand U2649 (N_2649,N_2315,N_2341);
nand U2650 (N_2650,N_2413,N_2308);
or U2651 (N_2651,N_2280,N_2293);
xnor U2652 (N_2652,N_2272,N_2373);
xor U2653 (N_2653,N_2446,N_2322);
nand U2654 (N_2654,N_2391,N_2389);
nand U2655 (N_2655,N_2315,N_2492);
nor U2656 (N_2656,N_2365,N_2401);
xnor U2657 (N_2657,N_2364,N_2286);
nand U2658 (N_2658,N_2444,N_2414);
or U2659 (N_2659,N_2339,N_2379);
nor U2660 (N_2660,N_2283,N_2328);
and U2661 (N_2661,N_2318,N_2412);
nor U2662 (N_2662,N_2357,N_2266);
nand U2663 (N_2663,N_2352,N_2456);
nor U2664 (N_2664,N_2303,N_2498);
nand U2665 (N_2665,N_2434,N_2268);
nand U2666 (N_2666,N_2392,N_2468);
or U2667 (N_2667,N_2430,N_2417);
nand U2668 (N_2668,N_2270,N_2327);
nand U2669 (N_2669,N_2492,N_2287);
nand U2670 (N_2670,N_2325,N_2288);
or U2671 (N_2671,N_2272,N_2468);
or U2672 (N_2672,N_2264,N_2467);
xnor U2673 (N_2673,N_2386,N_2307);
and U2674 (N_2674,N_2418,N_2313);
nand U2675 (N_2675,N_2304,N_2351);
nand U2676 (N_2676,N_2318,N_2470);
and U2677 (N_2677,N_2480,N_2272);
nor U2678 (N_2678,N_2402,N_2268);
and U2679 (N_2679,N_2340,N_2455);
nand U2680 (N_2680,N_2489,N_2362);
and U2681 (N_2681,N_2263,N_2422);
nor U2682 (N_2682,N_2426,N_2260);
and U2683 (N_2683,N_2415,N_2409);
nor U2684 (N_2684,N_2260,N_2435);
nand U2685 (N_2685,N_2413,N_2441);
nand U2686 (N_2686,N_2403,N_2447);
nor U2687 (N_2687,N_2309,N_2398);
and U2688 (N_2688,N_2271,N_2439);
and U2689 (N_2689,N_2444,N_2317);
and U2690 (N_2690,N_2372,N_2374);
and U2691 (N_2691,N_2370,N_2389);
nor U2692 (N_2692,N_2457,N_2432);
xnor U2693 (N_2693,N_2474,N_2363);
nor U2694 (N_2694,N_2307,N_2391);
nor U2695 (N_2695,N_2435,N_2282);
nor U2696 (N_2696,N_2408,N_2284);
nor U2697 (N_2697,N_2325,N_2293);
and U2698 (N_2698,N_2328,N_2264);
and U2699 (N_2699,N_2269,N_2327);
xor U2700 (N_2700,N_2399,N_2328);
nor U2701 (N_2701,N_2306,N_2404);
or U2702 (N_2702,N_2284,N_2293);
and U2703 (N_2703,N_2348,N_2455);
and U2704 (N_2704,N_2322,N_2351);
or U2705 (N_2705,N_2412,N_2338);
xor U2706 (N_2706,N_2263,N_2469);
and U2707 (N_2707,N_2325,N_2361);
and U2708 (N_2708,N_2281,N_2468);
nor U2709 (N_2709,N_2329,N_2310);
nor U2710 (N_2710,N_2342,N_2369);
nand U2711 (N_2711,N_2263,N_2324);
or U2712 (N_2712,N_2422,N_2255);
and U2713 (N_2713,N_2318,N_2254);
nor U2714 (N_2714,N_2438,N_2480);
or U2715 (N_2715,N_2458,N_2340);
xor U2716 (N_2716,N_2278,N_2436);
nand U2717 (N_2717,N_2379,N_2475);
or U2718 (N_2718,N_2355,N_2396);
xnor U2719 (N_2719,N_2401,N_2261);
or U2720 (N_2720,N_2447,N_2434);
or U2721 (N_2721,N_2464,N_2250);
nand U2722 (N_2722,N_2426,N_2428);
nand U2723 (N_2723,N_2299,N_2421);
nand U2724 (N_2724,N_2451,N_2428);
and U2725 (N_2725,N_2341,N_2312);
or U2726 (N_2726,N_2365,N_2314);
and U2727 (N_2727,N_2263,N_2412);
or U2728 (N_2728,N_2268,N_2273);
nand U2729 (N_2729,N_2282,N_2424);
and U2730 (N_2730,N_2403,N_2499);
and U2731 (N_2731,N_2483,N_2423);
nor U2732 (N_2732,N_2251,N_2351);
xnor U2733 (N_2733,N_2410,N_2421);
or U2734 (N_2734,N_2494,N_2347);
nor U2735 (N_2735,N_2499,N_2409);
xnor U2736 (N_2736,N_2300,N_2452);
or U2737 (N_2737,N_2437,N_2264);
and U2738 (N_2738,N_2320,N_2482);
xnor U2739 (N_2739,N_2427,N_2438);
or U2740 (N_2740,N_2485,N_2266);
and U2741 (N_2741,N_2449,N_2429);
nand U2742 (N_2742,N_2353,N_2389);
nand U2743 (N_2743,N_2316,N_2357);
or U2744 (N_2744,N_2432,N_2277);
xor U2745 (N_2745,N_2313,N_2499);
xor U2746 (N_2746,N_2285,N_2266);
or U2747 (N_2747,N_2366,N_2262);
nand U2748 (N_2748,N_2448,N_2339);
and U2749 (N_2749,N_2351,N_2342);
nand U2750 (N_2750,N_2507,N_2721);
and U2751 (N_2751,N_2610,N_2708);
and U2752 (N_2752,N_2618,N_2725);
nand U2753 (N_2753,N_2642,N_2624);
xor U2754 (N_2754,N_2713,N_2746);
nor U2755 (N_2755,N_2560,N_2651);
and U2756 (N_2756,N_2653,N_2536);
nand U2757 (N_2757,N_2644,N_2579);
and U2758 (N_2758,N_2611,N_2600);
and U2759 (N_2759,N_2679,N_2513);
or U2760 (N_2760,N_2733,N_2662);
and U2761 (N_2761,N_2565,N_2646);
nor U2762 (N_2762,N_2620,N_2722);
or U2763 (N_2763,N_2745,N_2728);
nand U2764 (N_2764,N_2572,N_2629);
and U2765 (N_2765,N_2524,N_2730);
nand U2766 (N_2766,N_2682,N_2688);
nand U2767 (N_2767,N_2580,N_2686);
and U2768 (N_2768,N_2720,N_2741);
nand U2769 (N_2769,N_2650,N_2661);
and U2770 (N_2770,N_2526,N_2707);
and U2771 (N_2771,N_2717,N_2607);
or U2772 (N_2772,N_2576,N_2568);
and U2773 (N_2773,N_2530,N_2598);
xor U2774 (N_2774,N_2664,N_2675);
and U2775 (N_2775,N_2564,N_2599);
xnor U2776 (N_2776,N_2515,N_2633);
and U2777 (N_2777,N_2590,N_2609);
and U2778 (N_2778,N_2547,N_2587);
nor U2779 (N_2779,N_2652,N_2692);
nand U2780 (N_2780,N_2593,N_2550);
nor U2781 (N_2781,N_2561,N_2663);
and U2782 (N_2782,N_2632,N_2527);
xor U2783 (N_2783,N_2696,N_2676);
xor U2784 (N_2784,N_2724,N_2578);
nand U2785 (N_2785,N_2567,N_2591);
and U2786 (N_2786,N_2539,N_2509);
and U2787 (N_2787,N_2573,N_2612);
and U2788 (N_2788,N_2672,N_2608);
xor U2789 (N_2789,N_2712,N_2525);
and U2790 (N_2790,N_2582,N_2678);
nor U2791 (N_2791,N_2709,N_2729);
xnor U2792 (N_2792,N_2695,N_2674);
nor U2793 (N_2793,N_2699,N_2702);
or U2794 (N_2794,N_2585,N_2641);
xnor U2795 (N_2795,N_2531,N_2583);
nor U2796 (N_2796,N_2541,N_2669);
nand U2797 (N_2797,N_2516,N_2706);
nor U2798 (N_2798,N_2630,N_2704);
or U2799 (N_2799,N_2700,N_2698);
or U2800 (N_2800,N_2691,N_2718);
or U2801 (N_2801,N_2736,N_2680);
xnor U2802 (N_2802,N_2606,N_2594);
or U2803 (N_2803,N_2654,N_2634);
or U2804 (N_2804,N_2538,N_2640);
nand U2805 (N_2805,N_2545,N_2559);
and U2806 (N_2806,N_2537,N_2555);
or U2807 (N_2807,N_2595,N_2657);
nand U2808 (N_2808,N_2687,N_2658);
nand U2809 (N_2809,N_2738,N_2744);
or U2810 (N_2810,N_2617,N_2747);
and U2811 (N_2811,N_2649,N_2512);
and U2812 (N_2812,N_2726,N_2740);
and U2813 (N_2813,N_2703,N_2616);
nand U2814 (N_2814,N_2500,N_2619);
or U2815 (N_2815,N_2570,N_2731);
nand U2816 (N_2816,N_2518,N_2643);
or U2817 (N_2817,N_2626,N_2532);
and U2818 (N_2818,N_2689,N_2670);
nor U2819 (N_2819,N_2571,N_2749);
xnor U2820 (N_2820,N_2519,N_2628);
nor U2821 (N_2821,N_2627,N_2723);
nor U2822 (N_2822,N_2522,N_2529);
and U2823 (N_2823,N_2521,N_2714);
and U2824 (N_2824,N_2710,N_2737);
nand U2825 (N_2825,N_2665,N_2533);
nor U2826 (N_2826,N_2558,N_2681);
xor U2827 (N_2827,N_2631,N_2563);
xor U2828 (N_2828,N_2562,N_2542);
nand U2829 (N_2829,N_2732,N_2656);
and U2830 (N_2830,N_2544,N_2711);
nand U2831 (N_2831,N_2543,N_2623);
or U2832 (N_2832,N_2546,N_2506);
nor U2833 (N_2833,N_2739,N_2734);
or U2834 (N_2834,N_2554,N_2715);
xor U2835 (N_2835,N_2666,N_2719);
xor U2836 (N_2836,N_2556,N_2647);
nor U2837 (N_2837,N_2552,N_2705);
or U2838 (N_2838,N_2508,N_2589);
or U2839 (N_2839,N_2684,N_2645);
xor U2840 (N_2840,N_2727,N_2637);
and U2841 (N_2841,N_2639,N_2671);
xor U2842 (N_2842,N_2569,N_2586);
or U2843 (N_2843,N_2735,N_2523);
nor U2844 (N_2844,N_2601,N_2502);
nor U2845 (N_2845,N_2605,N_2553);
nor U2846 (N_2846,N_2636,N_2520);
or U2847 (N_2847,N_2615,N_2551);
nand U2848 (N_2848,N_2505,N_2575);
nor U2849 (N_2849,N_2574,N_2549);
nand U2850 (N_2850,N_2602,N_2603);
and U2851 (N_2851,N_2504,N_2511);
nand U2852 (N_2852,N_2597,N_2668);
xnor U2853 (N_2853,N_2514,N_2604);
nor U2854 (N_2854,N_2638,N_2667);
xor U2855 (N_2855,N_2701,N_2697);
and U2856 (N_2856,N_2548,N_2621);
and U2857 (N_2857,N_2517,N_2584);
nand U2858 (N_2858,N_2528,N_2742);
or U2859 (N_2859,N_2535,N_2716);
xnor U2860 (N_2860,N_2748,N_2648);
or U2861 (N_2861,N_2577,N_2501);
nor U2862 (N_2862,N_2694,N_2557);
xnor U2863 (N_2863,N_2622,N_2659);
and U2864 (N_2864,N_2534,N_2503);
xor U2865 (N_2865,N_2510,N_2677);
and U2866 (N_2866,N_2596,N_2614);
and U2867 (N_2867,N_2635,N_2690);
nor U2868 (N_2868,N_2685,N_2655);
and U2869 (N_2869,N_2625,N_2673);
nor U2870 (N_2870,N_2566,N_2693);
xor U2871 (N_2871,N_2683,N_2588);
and U2872 (N_2872,N_2743,N_2540);
xnor U2873 (N_2873,N_2660,N_2592);
or U2874 (N_2874,N_2581,N_2613);
or U2875 (N_2875,N_2582,N_2595);
and U2876 (N_2876,N_2653,N_2644);
and U2877 (N_2877,N_2550,N_2516);
or U2878 (N_2878,N_2512,N_2628);
or U2879 (N_2879,N_2633,N_2577);
nand U2880 (N_2880,N_2617,N_2629);
nand U2881 (N_2881,N_2670,N_2723);
xor U2882 (N_2882,N_2730,N_2527);
nor U2883 (N_2883,N_2589,N_2697);
and U2884 (N_2884,N_2736,N_2607);
and U2885 (N_2885,N_2584,N_2625);
or U2886 (N_2886,N_2686,N_2542);
nor U2887 (N_2887,N_2670,N_2660);
nor U2888 (N_2888,N_2581,N_2622);
xor U2889 (N_2889,N_2672,N_2607);
nor U2890 (N_2890,N_2675,N_2553);
xnor U2891 (N_2891,N_2646,N_2710);
or U2892 (N_2892,N_2610,N_2706);
or U2893 (N_2893,N_2743,N_2575);
and U2894 (N_2894,N_2744,N_2549);
or U2895 (N_2895,N_2572,N_2583);
and U2896 (N_2896,N_2641,N_2574);
and U2897 (N_2897,N_2691,N_2654);
nor U2898 (N_2898,N_2545,N_2638);
and U2899 (N_2899,N_2668,N_2525);
and U2900 (N_2900,N_2592,N_2513);
xor U2901 (N_2901,N_2641,N_2618);
nor U2902 (N_2902,N_2560,N_2631);
and U2903 (N_2903,N_2675,N_2652);
nor U2904 (N_2904,N_2642,N_2585);
and U2905 (N_2905,N_2524,N_2533);
and U2906 (N_2906,N_2626,N_2663);
nor U2907 (N_2907,N_2524,N_2680);
xnor U2908 (N_2908,N_2641,N_2591);
and U2909 (N_2909,N_2683,N_2716);
nand U2910 (N_2910,N_2555,N_2595);
and U2911 (N_2911,N_2588,N_2673);
and U2912 (N_2912,N_2547,N_2606);
nand U2913 (N_2913,N_2501,N_2597);
nor U2914 (N_2914,N_2530,N_2748);
or U2915 (N_2915,N_2633,N_2538);
nand U2916 (N_2916,N_2542,N_2682);
xor U2917 (N_2917,N_2565,N_2667);
or U2918 (N_2918,N_2572,N_2717);
and U2919 (N_2919,N_2631,N_2726);
xnor U2920 (N_2920,N_2687,N_2535);
xor U2921 (N_2921,N_2731,N_2579);
xnor U2922 (N_2922,N_2719,N_2520);
nand U2923 (N_2923,N_2605,N_2620);
xor U2924 (N_2924,N_2555,N_2653);
nor U2925 (N_2925,N_2539,N_2558);
and U2926 (N_2926,N_2524,N_2557);
nor U2927 (N_2927,N_2506,N_2741);
nor U2928 (N_2928,N_2695,N_2566);
xor U2929 (N_2929,N_2608,N_2710);
nor U2930 (N_2930,N_2712,N_2744);
and U2931 (N_2931,N_2633,N_2718);
or U2932 (N_2932,N_2570,N_2726);
xor U2933 (N_2933,N_2690,N_2652);
nor U2934 (N_2934,N_2691,N_2529);
xor U2935 (N_2935,N_2646,N_2506);
xor U2936 (N_2936,N_2719,N_2693);
and U2937 (N_2937,N_2573,N_2692);
and U2938 (N_2938,N_2587,N_2563);
xnor U2939 (N_2939,N_2525,N_2612);
nor U2940 (N_2940,N_2574,N_2602);
or U2941 (N_2941,N_2540,N_2746);
or U2942 (N_2942,N_2570,N_2527);
nor U2943 (N_2943,N_2566,N_2732);
xnor U2944 (N_2944,N_2597,N_2559);
nand U2945 (N_2945,N_2603,N_2567);
or U2946 (N_2946,N_2627,N_2710);
and U2947 (N_2947,N_2723,N_2676);
nor U2948 (N_2948,N_2720,N_2746);
or U2949 (N_2949,N_2736,N_2540);
or U2950 (N_2950,N_2692,N_2544);
and U2951 (N_2951,N_2634,N_2529);
xnor U2952 (N_2952,N_2735,N_2692);
and U2953 (N_2953,N_2615,N_2729);
xor U2954 (N_2954,N_2653,N_2542);
xnor U2955 (N_2955,N_2649,N_2506);
or U2956 (N_2956,N_2648,N_2708);
xnor U2957 (N_2957,N_2567,N_2734);
nand U2958 (N_2958,N_2539,N_2681);
and U2959 (N_2959,N_2678,N_2709);
nor U2960 (N_2960,N_2584,N_2700);
nand U2961 (N_2961,N_2687,N_2725);
nand U2962 (N_2962,N_2587,N_2595);
nand U2963 (N_2963,N_2552,N_2666);
or U2964 (N_2964,N_2681,N_2676);
xor U2965 (N_2965,N_2635,N_2712);
and U2966 (N_2966,N_2707,N_2712);
nor U2967 (N_2967,N_2624,N_2654);
nor U2968 (N_2968,N_2703,N_2525);
xor U2969 (N_2969,N_2703,N_2732);
or U2970 (N_2970,N_2515,N_2594);
nor U2971 (N_2971,N_2640,N_2614);
or U2972 (N_2972,N_2609,N_2550);
or U2973 (N_2973,N_2620,N_2547);
xnor U2974 (N_2974,N_2523,N_2624);
nor U2975 (N_2975,N_2542,N_2738);
and U2976 (N_2976,N_2656,N_2654);
nor U2977 (N_2977,N_2509,N_2707);
nor U2978 (N_2978,N_2669,N_2516);
nor U2979 (N_2979,N_2746,N_2739);
xor U2980 (N_2980,N_2578,N_2659);
and U2981 (N_2981,N_2522,N_2664);
and U2982 (N_2982,N_2615,N_2741);
nor U2983 (N_2983,N_2671,N_2527);
nor U2984 (N_2984,N_2507,N_2523);
xor U2985 (N_2985,N_2554,N_2536);
xnor U2986 (N_2986,N_2741,N_2694);
nand U2987 (N_2987,N_2586,N_2683);
xnor U2988 (N_2988,N_2683,N_2545);
and U2989 (N_2989,N_2543,N_2539);
nand U2990 (N_2990,N_2690,N_2642);
nand U2991 (N_2991,N_2689,N_2505);
nand U2992 (N_2992,N_2669,N_2744);
and U2993 (N_2993,N_2654,N_2611);
and U2994 (N_2994,N_2580,N_2572);
nor U2995 (N_2995,N_2686,N_2653);
and U2996 (N_2996,N_2664,N_2551);
xnor U2997 (N_2997,N_2695,N_2715);
nor U2998 (N_2998,N_2604,N_2702);
nor U2999 (N_2999,N_2722,N_2616);
nand U3000 (N_3000,N_2937,N_2909);
nor U3001 (N_3001,N_2807,N_2808);
and U3002 (N_3002,N_2759,N_2900);
or U3003 (N_3003,N_2978,N_2813);
or U3004 (N_3004,N_2964,N_2819);
nor U3005 (N_3005,N_2907,N_2851);
nor U3006 (N_3006,N_2848,N_2893);
xnor U3007 (N_3007,N_2864,N_2873);
nand U3008 (N_3008,N_2932,N_2857);
nor U3009 (N_3009,N_2891,N_2753);
xor U3010 (N_3010,N_2804,N_2858);
nand U3011 (N_3011,N_2809,N_2999);
xor U3012 (N_3012,N_2773,N_2788);
or U3013 (N_3013,N_2765,N_2866);
xnor U3014 (N_3014,N_2822,N_2918);
and U3015 (N_3015,N_2885,N_2842);
nand U3016 (N_3016,N_2993,N_2958);
nand U3017 (N_3017,N_2985,N_2942);
nand U3018 (N_3018,N_2938,N_2935);
nand U3019 (N_3019,N_2766,N_2856);
nor U3020 (N_3020,N_2929,N_2795);
and U3021 (N_3021,N_2820,N_2855);
nand U3022 (N_3022,N_2976,N_2781);
and U3023 (N_3023,N_2810,N_2859);
or U3024 (N_3024,N_2934,N_2940);
and U3025 (N_3025,N_2923,N_2965);
xnor U3026 (N_3026,N_2862,N_2984);
or U3027 (N_3027,N_2975,N_2756);
or U3028 (N_3028,N_2752,N_2877);
nor U3029 (N_3029,N_2917,N_2959);
nand U3030 (N_3030,N_2950,N_2802);
nor U3031 (N_3031,N_2869,N_2779);
nand U3032 (N_3032,N_2751,N_2780);
or U3033 (N_3033,N_2894,N_2931);
nand U3034 (N_3034,N_2990,N_2953);
nand U3035 (N_3035,N_2829,N_2969);
and U3036 (N_3036,N_2811,N_2995);
nand U3037 (N_3037,N_2833,N_2835);
and U3038 (N_3038,N_2831,N_2761);
or U3039 (N_3039,N_2889,N_2824);
nand U3040 (N_3040,N_2988,N_2956);
and U3041 (N_3041,N_2830,N_2878);
and U3042 (N_3042,N_2767,N_2800);
and U3043 (N_3043,N_2832,N_2883);
nor U3044 (N_3044,N_2963,N_2881);
or U3045 (N_3045,N_2794,N_2774);
nor U3046 (N_3046,N_2943,N_2998);
or U3047 (N_3047,N_2768,N_2754);
or U3048 (N_3048,N_2861,N_2896);
and U3049 (N_3049,N_2933,N_2930);
or U3050 (N_3050,N_2845,N_2871);
xnor U3051 (N_3051,N_2758,N_2901);
nor U3052 (N_3052,N_2805,N_2836);
or U3053 (N_3053,N_2903,N_2874);
xnor U3054 (N_3054,N_2983,N_2916);
or U3055 (N_3055,N_2875,N_2823);
and U3056 (N_3056,N_2818,N_2913);
nor U3057 (N_3057,N_2952,N_2868);
or U3058 (N_3058,N_2910,N_2801);
nand U3059 (N_3059,N_2936,N_2921);
xnor U3060 (N_3060,N_2815,N_2991);
nand U3061 (N_3061,N_2782,N_2927);
and U3062 (N_3062,N_2949,N_2772);
xnor U3063 (N_3063,N_2899,N_2863);
or U3064 (N_3064,N_2787,N_2939);
nand U3065 (N_3065,N_2895,N_2890);
or U3066 (N_3066,N_2853,N_2989);
nand U3067 (N_3067,N_2986,N_2840);
xnor U3068 (N_3068,N_2915,N_2926);
or U3069 (N_3069,N_2816,N_2902);
nor U3070 (N_3070,N_2783,N_2797);
nor U3071 (N_3071,N_2971,N_2867);
xnor U3072 (N_3072,N_2945,N_2860);
xnor U3073 (N_3073,N_2947,N_2821);
and U3074 (N_3074,N_2888,N_2996);
xor U3075 (N_3075,N_2799,N_2914);
xnor U3076 (N_3076,N_2898,N_2960);
xnor U3077 (N_3077,N_2849,N_2967);
and U3078 (N_3078,N_2944,N_2786);
nand U3079 (N_3079,N_2948,N_2897);
nor U3080 (N_3080,N_2957,N_2973);
or U3081 (N_3081,N_2928,N_2962);
nand U3082 (N_3082,N_2852,N_2979);
nand U3083 (N_3083,N_2972,N_2760);
nand U3084 (N_3084,N_2763,N_2884);
nor U3085 (N_3085,N_2762,N_2784);
and U3086 (N_3086,N_2846,N_2764);
nor U3087 (N_3087,N_2755,N_2887);
nor U3088 (N_3088,N_2980,N_2865);
nand U3089 (N_3089,N_2825,N_2798);
or U3090 (N_3090,N_2771,N_2776);
and U3091 (N_3091,N_2843,N_2997);
xor U3092 (N_3092,N_2922,N_2977);
nand U3093 (N_3093,N_2812,N_2775);
nand U3094 (N_3094,N_2777,N_2912);
or U3095 (N_3095,N_2924,N_2828);
nand U3096 (N_3096,N_2908,N_2880);
or U3097 (N_3097,N_2837,N_2941);
xnor U3098 (N_3098,N_2981,N_2904);
nor U3099 (N_3099,N_2968,N_2982);
nand U3100 (N_3100,N_2882,N_2974);
and U3101 (N_3101,N_2886,N_2920);
nor U3102 (N_3102,N_2789,N_2757);
nor U3103 (N_3103,N_2872,N_2992);
nor U3104 (N_3104,N_2750,N_2906);
nor U3105 (N_3105,N_2791,N_2827);
nand U3106 (N_3106,N_2870,N_2796);
nand U3107 (N_3107,N_2769,N_2778);
nand U3108 (N_3108,N_2925,N_2841);
nand U3109 (N_3109,N_2919,N_2951);
or U3110 (N_3110,N_2838,N_2879);
or U3111 (N_3111,N_2955,N_2905);
and U3112 (N_3112,N_2770,N_2785);
and U3113 (N_3113,N_2844,N_2839);
or U3114 (N_3114,N_2987,N_2850);
nor U3115 (N_3115,N_2854,N_2970);
nor U3116 (N_3116,N_2817,N_2793);
nor U3117 (N_3117,N_2946,N_2847);
nand U3118 (N_3118,N_2792,N_2954);
nand U3119 (N_3119,N_2966,N_2803);
or U3120 (N_3120,N_2892,N_2806);
nand U3121 (N_3121,N_2790,N_2834);
nor U3122 (N_3122,N_2961,N_2994);
nor U3123 (N_3123,N_2876,N_2814);
or U3124 (N_3124,N_2911,N_2826);
or U3125 (N_3125,N_2931,N_2850);
xnor U3126 (N_3126,N_2799,N_2804);
and U3127 (N_3127,N_2778,N_2918);
or U3128 (N_3128,N_2750,N_2837);
nand U3129 (N_3129,N_2768,N_2807);
or U3130 (N_3130,N_2852,N_2860);
nand U3131 (N_3131,N_2937,N_2942);
or U3132 (N_3132,N_2932,N_2750);
and U3133 (N_3133,N_2773,N_2750);
nand U3134 (N_3134,N_2895,N_2827);
nor U3135 (N_3135,N_2772,N_2779);
or U3136 (N_3136,N_2867,N_2779);
or U3137 (N_3137,N_2935,N_2939);
and U3138 (N_3138,N_2931,N_2935);
nand U3139 (N_3139,N_2934,N_2989);
and U3140 (N_3140,N_2783,N_2943);
xor U3141 (N_3141,N_2977,N_2949);
xor U3142 (N_3142,N_2846,N_2834);
xnor U3143 (N_3143,N_2879,N_2963);
xnor U3144 (N_3144,N_2763,N_2890);
and U3145 (N_3145,N_2755,N_2800);
or U3146 (N_3146,N_2881,N_2993);
nand U3147 (N_3147,N_2869,N_2937);
xor U3148 (N_3148,N_2905,N_2776);
nand U3149 (N_3149,N_2913,N_2920);
and U3150 (N_3150,N_2814,N_2815);
xnor U3151 (N_3151,N_2795,N_2900);
nand U3152 (N_3152,N_2986,N_2767);
or U3153 (N_3153,N_2805,N_2781);
and U3154 (N_3154,N_2809,N_2934);
nor U3155 (N_3155,N_2931,N_2753);
and U3156 (N_3156,N_2792,N_2866);
or U3157 (N_3157,N_2963,N_2893);
nor U3158 (N_3158,N_2805,N_2822);
or U3159 (N_3159,N_2795,N_2854);
xnor U3160 (N_3160,N_2777,N_2852);
xor U3161 (N_3161,N_2812,N_2965);
and U3162 (N_3162,N_2953,N_2842);
nor U3163 (N_3163,N_2994,N_2917);
nand U3164 (N_3164,N_2945,N_2845);
and U3165 (N_3165,N_2897,N_2966);
nand U3166 (N_3166,N_2812,N_2825);
xor U3167 (N_3167,N_2894,N_2979);
nor U3168 (N_3168,N_2999,N_2995);
and U3169 (N_3169,N_2866,N_2927);
xor U3170 (N_3170,N_2968,N_2752);
nand U3171 (N_3171,N_2961,N_2893);
nor U3172 (N_3172,N_2898,N_2776);
nand U3173 (N_3173,N_2832,N_2890);
and U3174 (N_3174,N_2798,N_2890);
xnor U3175 (N_3175,N_2853,N_2908);
xnor U3176 (N_3176,N_2984,N_2948);
xor U3177 (N_3177,N_2754,N_2816);
nand U3178 (N_3178,N_2763,N_2815);
nor U3179 (N_3179,N_2788,N_2751);
xnor U3180 (N_3180,N_2963,N_2760);
or U3181 (N_3181,N_2946,N_2943);
or U3182 (N_3182,N_2758,N_2944);
xor U3183 (N_3183,N_2915,N_2761);
nor U3184 (N_3184,N_2765,N_2956);
xnor U3185 (N_3185,N_2835,N_2917);
nand U3186 (N_3186,N_2767,N_2916);
nand U3187 (N_3187,N_2946,N_2834);
and U3188 (N_3188,N_2935,N_2862);
nor U3189 (N_3189,N_2974,N_2866);
and U3190 (N_3190,N_2769,N_2753);
xor U3191 (N_3191,N_2827,N_2963);
and U3192 (N_3192,N_2781,N_2836);
nor U3193 (N_3193,N_2896,N_2972);
or U3194 (N_3194,N_2804,N_2915);
nor U3195 (N_3195,N_2887,N_2800);
or U3196 (N_3196,N_2928,N_2875);
or U3197 (N_3197,N_2750,N_2916);
nor U3198 (N_3198,N_2844,N_2952);
nand U3199 (N_3199,N_2755,N_2975);
xnor U3200 (N_3200,N_2769,N_2784);
or U3201 (N_3201,N_2831,N_2959);
nor U3202 (N_3202,N_2839,N_2915);
or U3203 (N_3203,N_2876,N_2859);
and U3204 (N_3204,N_2810,N_2987);
xor U3205 (N_3205,N_2844,N_2905);
nand U3206 (N_3206,N_2842,N_2887);
and U3207 (N_3207,N_2805,N_2759);
and U3208 (N_3208,N_2760,N_2807);
and U3209 (N_3209,N_2807,N_2983);
nor U3210 (N_3210,N_2767,N_2995);
nand U3211 (N_3211,N_2792,N_2801);
and U3212 (N_3212,N_2782,N_2770);
nor U3213 (N_3213,N_2806,N_2846);
nor U3214 (N_3214,N_2824,N_2964);
nor U3215 (N_3215,N_2811,N_2899);
and U3216 (N_3216,N_2940,N_2798);
xnor U3217 (N_3217,N_2946,N_2783);
nor U3218 (N_3218,N_2773,N_2939);
xnor U3219 (N_3219,N_2839,N_2919);
nand U3220 (N_3220,N_2849,N_2880);
nor U3221 (N_3221,N_2892,N_2988);
or U3222 (N_3222,N_2819,N_2751);
nor U3223 (N_3223,N_2969,N_2941);
xor U3224 (N_3224,N_2868,N_2964);
nand U3225 (N_3225,N_2979,N_2840);
or U3226 (N_3226,N_2801,N_2806);
and U3227 (N_3227,N_2819,N_2908);
or U3228 (N_3228,N_2837,N_2876);
nand U3229 (N_3229,N_2857,N_2847);
nand U3230 (N_3230,N_2930,N_2839);
and U3231 (N_3231,N_2767,N_2811);
xnor U3232 (N_3232,N_2862,N_2871);
xor U3233 (N_3233,N_2756,N_2896);
xor U3234 (N_3234,N_2762,N_2886);
nor U3235 (N_3235,N_2769,N_2751);
xnor U3236 (N_3236,N_2946,N_2786);
nor U3237 (N_3237,N_2971,N_2959);
xnor U3238 (N_3238,N_2804,N_2960);
nand U3239 (N_3239,N_2973,N_2954);
or U3240 (N_3240,N_2931,N_2973);
nor U3241 (N_3241,N_2971,N_2776);
and U3242 (N_3242,N_2882,N_2766);
nor U3243 (N_3243,N_2893,N_2773);
nand U3244 (N_3244,N_2788,N_2973);
and U3245 (N_3245,N_2869,N_2901);
nor U3246 (N_3246,N_2819,N_2867);
nor U3247 (N_3247,N_2773,N_2948);
nor U3248 (N_3248,N_2754,N_2961);
and U3249 (N_3249,N_2887,N_2949);
nor U3250 (N_3250,N_3027,N_3093);
nand U3251 (N_3251,N_3085,N_3072);
nor U3252 (N_3252,N_3003,N_3062);
xor U3253 (N_3253,N_3104,N_3133);
and U3254 (N_3254,N_3078,N_3198);
nor U3255 (N_3255,N_3102,N_3241);
and U3256 (N_3256,N_3197,N_3022);
or U3257 (N_3257,N_3118,N_3081);
xnor U3258 (N_3258,N_3245,N_3044);
nand U3259 (N_3259,N_3225,N_3184);
xnor U3260 (N_3260,N_3105,N_3191);
nor U3261 (N_3261,N_3060,N_3006);
nor U3262 (N_3262,N_3100,N_3247);
or U3263 (N_3263,N_3106,N_3140);
nor U3264 (N_3264,N_3094,N_3188);
nor U3265 (N_3265,N_3190,N_3182);
or U3266 (N_3266,N_3178,N_3200);
xnor U3267 (N_3267,N_3013,N_3199);
xnor U3268 (N_3268,N_3208,N_3015);
nor U3269 (N_3269,N_3186,N_3171);
xor U3270 (N_3270,N_3244,N_3090);
nand U3271 (N_3271,N_3172,N_3150);
xnor U3272 (N_3272,N_3210,N_3214);
nor U3273 (N_3273,N_3152,N_3056);
and U3274 (N_3274,N_3074,N_3234);
xnor U3275 (N_3275,N_3219,N_3235);
xor U3276 (N_3276,N_3157,N_3032);
or U3277 (N_3277,N_3057,N_3046);
nor U3278 (N_3278,N_3114,N_3024);
nor U3279 (N_3279,N_3069,N_3142);
and U3280 (N_3280,N_3159,N_3227);
xor U3281 (N_3281,N_3113,N_3066);
nor U3282 (N_3282,N_3124,N_3127);
xor U3283 (N_3283,N_3092,N_3224);
or U3284 (N_3284,N_3165,N_3000);
nor U3285 (N_3285,N_3248,N_3033);
nand U3286 (N_3286,N_3231,N_3230);
xnor U3287 (N_3287,N_3059,N_3193);
nor U3288 (N_3288,N_3161,N_3091);
nor U3289 (N_3289,N_3026,N_3229);
and U3290 (N_3290,N_3131,N_3134);
nor U3291 (N_3291,N_3132,N_3052);
xnor U3292 (N_3292,N_3109,N_3168);
or U3293 (N_3293,N_3023,N_3147);
xnor U3294 (N_3294,N_3146,N_3122);
and U3295 (N_3295,N_3045,N_3086);
nor U3296 (N_3296,N_3116,N_3179);
nand U3297 (N_3297,N_3129,N_3055);
xnor U3298 (N_3298,N_3183,N_3149);
nand U3299 (N_3299,N_3119,N_3038);
nand U3300 (N_3300,N_3110,N_3007);
or U3301 (N_3301,N_3151,N_3148);
and U3302 (N_3302,N_3195,N_3061);
and U3303 (N_3303,N_3173,N_3115);
and U3304 (N_3304,N_3240,N_3189);
or U3305 (N_3305,N_3097,N_3123);
nand U3306 (N_3306,N_3121,N_3242);
xor U3307 (N_3307,N_3192,N_3065);
nor U3308 (N_3308,N_3163,N_3169);
and U3309 (N_3309,N_3226,N_3028);
nand U3310 (N_3310,N_3220,N_3041);
xor U3311 (N_3311,N_3036,N_3130);
xnor U3312 (N_3312,N_3137,N_3181);
or U3313 (N_3313,N_3040,N_3099);
nor U3314 (N_3314,N_3243,N_3143);
nor U3315 (N_3315,N_3216,N_3030);
and U3316 (N_3316,N_3098,N_3180);
and U3317 (N_3317,N_3237,N_3201);
and U3318 (N_3318,N_3016,N_3073);
or U3319 (N_3319,N_3096,N_3010);
nor U3320 (N_3320,N_3095,N_3012);
nor U3321 (N_3321,N_3205,N_3031);
and U3322 (N_3322,N_3138,N_3029);
and U3323 (N_3323,N_3017,N_3203);
xnor U3324 (N_3324,N_3037,N_3067);
nand U3325 (N_3325,N_3042,N_3054);
nand U3326 (N_3326,N_3177,N_3202);
xnor U3327 (N_3327,N_3153,N_3047);
and U3328 (N_3328,N_3246,N_3126);
xnor U3329 (N_3329,N_3077,N_3136);
and U3330 (N_3330,N_3020,N_3079);
and U3331 (N_3331,N_3228,N_3004);
nand U3332 (N_3332,N_3160,N_3107);
nand U3333 (N_3333,N_3058,N_3048);
and U3334 (N_3334,N_3011,N_3164);
xnor U3335 (N_3335,N_3014,N_3236);
and U3336 (N_3336,N_3158,N_3112);
nor U3337 (N_3337,N_3043,N_3128);
or U3338 (N_3338,N_3084,N_3209);
xnor U3339 (N_3339,N_3144,N_3141);
nand U3340 (N_3340,N_3162,N_3238);
and U3341 (N_3341,N_3005,N_3194);
or U3342 (N_3342,N_3232,N_3021);
nand U3343 (N_3343,N_3111,N_3049);
and U3344 (N_3344,N_3204,N_3117);
and U3345 (N_3345,N_3239,N_3145);
and U3346 (N_3346,N_3002,N_3070);
nand U3347 (N_3347,N_3215,N_3185);
nand U3348 (N_3348,N_3139,N_3125);
and U3349 (N_3349,N_3089,N_3222);
nor U3350 (N_3350,N_3156,N_3068);
and U3351 (N_3351,N_3218,N_3249);
or U3352 (N_3352,N_3050,N_3064);
nand U3353 (N_3353,N_3087,N_3108);
or U3354 (N_3354,N_3076,N_3167);
xor U3355 (N_3355,N_3082,N_3008);
nor U3356 (N_3356,N_3213,N_3083);
nor U3357 (N_3357,N_3154,N_3039);
and U3358 (N_3358,N_3166,N_3075);
or U3359 (N_3359,N_3174,N_3018);
or U3360 (N_3360,N_3009,N_3120);
nand U3361 (N_3361,N_3001,N_3103);
nor U3362 (N_3362,N_3207,N_3212);
xor U3363 (N_3363,N_3035,N_3080);
nor U3364 (N_3364,N_3217,N_3175);
and U3365 (N_3365,N_3088,N_3223);
and U3366 (N_3366,N_3019,N_3051);
nand U3367 (N_3367,N_3221,N_3211);
or U3368 (N_3368,N_3135,N_3025);
and U3369 (N_3369,N_3187,N_3053);
xnor U3370 (N_3370,N_3155,N_3206);
xor U3371 (N_3371,N_3170,N_3063);
xnor U3372 (N_3372,N_3233,N_3176);
xor U3373 (N_3373,N_3071,N_3196);
nand U3374 (N_3374,N_3101,N_3034);
nor U3375 (N_3375,N_3212,N_3169);
xnor U3376 (N_3376,N_3240,N_3162);
nor U3377 (N_3377,N_3181,N_3000);
or U3378 (N_3378,N_3162,N_3074);
or U3379 (N_3379,N_3019,N_3140);
or U3380 (N_3380,N_3096,N_3041);
nand U3381 (N_3381,N_3147,N_3062);
nand U3382 (N_3382,N_3008,N_3077);
or U3383 (N_3383,N_3155,N_3067);
nand U3384 (N_3384,N_3117,N_3240);
nand U3385 (N_3385,N_3125,N_3145);
or U3386 (N_3386,N_3222,N_3171);
nor U3387 (N_3387,N_3073,N_3105);
xor U3388 (N_3388,N_3178,N_3246);
and U3389 (N_3389,N_3110,N_3156);
or U3390 (N_3390,N_3213,N_3013);
or U3391 (N_3391,N_3032,N_3128);
and U3392 (N_3392,N_3087,N_3155);
and U3393 (N_3393,N_3038,N_3077);
and U3394 (N_3394,N_3185,N_3030);
nor U3395 (N_3395,N_3071,N_3230);
nand U3396 (N_3396,N_3191,N_3234);
xor U3397 (N_3397,N_3237,N_3117);
or U3398 (N_3398,N_3185,N_3207);
nand U3399 (N_3399,N_3065,N_3115);
nand U3400 (N_3400,N_3068,N_3047);
or U3401 (N_3401,N_3129,N_3240);
and U3402 (N_3402,N_3016,N_3237);
nand U3403 (N_3403,N_3102,N_3076);
or U3404 (N_3404,N_3218,N_3112);
and U3405 (N_3405,N_3215,N_3179);
and U3406 (N_3406,N_3138,N_3099);
xnor U3407 (N_3407,N_3242,N_3110);
nor U3408 (N_3408,N_3141,N_3193);
or U3409 (N_3409,N_3158,N_3048);
and U3410 (N_3410,N_3228,N_3141);
or U3411 (N_3411,N_3063,N_3026);
nor U3412 (N_3412,N_3029,N_3203);
or U3413 (N_3413,N_3077,N_3200);
and U3414 (N_3414,N_3046,N_3087);
xnor U3415 (N_3415,N_3049,N_3004);
or U3416 (N_3416,N_3040,N_3192);
nand U3417 (N_3417,N_3056,N_3100);
or U3418 (N_3418,N_3034,N_3243);
and U3419 (N_3419,N_3238,N_3215);
nor U3420 (N_3420,N_3045,N_3211);
or U3421 (N_3421,N_3078,N_3103);
or U3422 (N_3422,N_3191,N_3206);
nand U3423 (N_3423,N_3068,N_3171);
and U3424 (N_3424,N_3192,N_3140);
or U3425 (N_3425,N_3206,N_3170);
nand U3426 (N_3426,N_3128,N_3105);
and U3427 (N_3427,N_3085,N_3036);
and U3428 (N_3428,N_3232,N_3027);
xor U3429 (N_3429,N_3226,N_3064);
or U3430 (N_3430,N_3145,N_3022);
or U3431 (N_3431,N_3192,N_3058);
nand U3432 (N_3432,N_3102,N_3163);
and U3433 (N_3433,N_3226,N_3133);
xor U3434 (N_3434,N_3145,N_3192);
xnor U3435 (N_3435,N_3089,N_3212);
nor U3436 (N_3436,N_3073,N_3111);
xor U3437 (N_3437,N_3075,N_3152);
xor U3438 (N_3438,N_3119,N_3011);
xnor U3439 (N_3439,N_3174,N_3164);
nor U3440 (N_3440,N_3108,N_3214);
xor U3441 (N_3441,N_3139,N_3012);
or U3442 (N_3442,N_3001,N_3070);
or U3443 (N_3443,N_3018,N_3026);
xnor U3444 (N_3444,N_3034,N_3119);
and U3445 (N_3445,N_3034,N_3031);
and U3446 (N_3446,N_3185,N_3096);
xor U3447 (N_3447,N_3152,N_3130);
xnor U3448 (N_3448,N_3013,N_3077);
nor U3449 (N_3449,N_3162,N_3191);
or U3450 (N_3450,N_3140,N_3208);
nor U3451 (N_3451,N_3006,N_3174);
xnor U3452 (N_3452,N_3198,N_3157);
nor U3453 (N_3453,N_3134,N_3000);
and U3454 (N_3454,N_3055,N_3209);
and U3455 (N_3455,N_3156,N_3028);
nand U3456 (N_3456,N_3024,N_3165);
nand U3457 (N_3457,N_3217,N_3191);
nor U3458 (N_3458,N_3220,N_3154);
or U3459 (N_3459,N_3132,N_3241);
xor U3460 (N_3460,N_3051,N_3023);
xor U3461 (N_3461,N_3235,N_3037);
nand U3462 (N_3462,N_3212,N_3092);
nand U3463 (N_3463,N_3050,N_3126);
nand U3464 (N_3464,N_3070,N_3055);
or U3465 (N_3465,N_3233,N_3137);
nor U3466 (N_3466,N_3154,N_3102);
or U3467 (N_3467,N_3146,N_3233);
xor U3468 (N_3468,N_3009,N_3036);
xnor U3469 (N_3469,N_3003,N_3079);
or U3470 (N_3470,N_3181,N_3224);
or U3471 (N_3471,N_3018,N_3156);
xor U3472 (N_3472,N_3201,N_3173);
or U3473 (N_3473,N_3083,N_3032);
xor U3474 (N_3474,N_3224,N_3015);
nor U3475 (N_3475,N_3245,N_3114);
or U3476 (N_3476,N_3192,N_3109);
and U3477 (N_3477,N_3108,N_3153);
and U3478 (N_3478,N_3073,N_3035);
xor U3479 (N_3479,N_3131,N_3020);
and U3480 (N_3480,N_3096,N_3042);
and U3481 (N_3481,N_3173,N_3000);
nand U3482 (N_3482,N_3236,N_3091);
nor U3483 (N_3483,N_3059,N_3140);
xor U3484 (N_3484,N_3020,N_3096);
xnor U3485 (N_3485,N_3114,N_3002);
or U3486 (N_3486,N_3124,N_3248);
or U3487 (N_3487,N_3030,N_3215);
and U3488 (N_3488,N_3108,N_3047);
and U3489 (N_3489,N_3209,N_3178);
xnor U3490 (N_3490,N_3023,N_3219);
or U3491 (N_3491,N_3226,N_3212);
or U3492 (N_3492,N_3216,N_3006);
xnor U3493 (N_3493,N_3234,N_3134);
nor U3494 (N_3494,N_3009,N_3240);
nand U3495 (N_3495,N_3040,N_3190);
and U3496 (N_3496,N_3124,N_3140);
nand U3497 (N_3497,N_3122,N_3031);
nand U3498 (N_3498,N_3228,N_3163);
xnor U3499 (N_3499,N_3095,N_3004);
xor U3500 (N_3500,N_3487,N_3445);
and U3501 (N_3501,N_3422,N_3464);
nand U3502 (N_3502,N_3428,N_3307);
or U3503 (N_3503,N_3356,N_3410);
or U3504 (N_3504,N_3308,N_3296);
xor U3505 (N_3505,N_3455,N_3411);
or U3506 (N_3506,N_3279,N_3477);
nand U3507 (N_3507,N_3355,N_3453);
or U3508 (N_3508,N_3479,N_3350);
nor U3509 (N_3509,N_3274,N_3393);
xnor U3510 (N_3510,N_3302,N_3435);
xnor U3511 (N_3511,N_3348,N_3374);
and U3512 (N_3512,N_3354,N_3475);
xnor U3513 (N_3513,N_3347,N_3363);
nand U3514 (N_3514,N_3346,N_3291);
xnor U3515 (N_3515,N_3367,N_3266);
nand U3516 (N_3516,N_3462,N_3421);
xnor U3517 (N_3517,N_3285,N_3376);
xor U3518 (N_3518,N_3265,N_3353);
xnor U3519 (N_3519,N_3398,N_3481);
xnor U3520 (N_3520,N_3454,N_3264);
nor U3521 (N_3521,N_3322,N_3489);
and U3522 (N_3522,N_3324,N_3309);
or U3523 (N_3523,N_3345,N_3305);
and U3524 (N_3524,N_3333,N_3391);
nor U3525 (N_3525,N_3463,N_3427);
nand U3526 (N_3526,N_3271,N_3289);
nand U3527 (N_3527,N_3405,N_3250);
or U3528 (N_3528,N_3277,N_3303);
xnor U3529 (N_3529,N_3442,N_3377);
nor U3530 (N_3530,N_3495,N_3280);
xnor U3531 (N_3531,N_3425,N_3297);
nand U3532 (N_3532,N_3287,N_3384);
xor U3533 (N_3533,N_3432,N_3357);
and U3534 (N_3534,N_3358,N_3491);
or U3535 (N_3535,N_3300,N_3449);
nand U3536 (N_3536,N_3434,N_3292);
nor U3537 (N_3537,N_3318,N_3360);
or U3538 (N_3538,N_3373,N_3419);
nand U3539 (N_3539,N_3320,N_3493);
and U3540 (N_3540,N_3415,N_3440);
or U3541 (N_3541,N_3254,N_3331);
and U3542 (N_3542,N_3402,N_3337);
xnor U3543 (N_3543,N_3334,N_3286);
and U3544 (N_3544,N_3490,N_3283);
xnor U3545 (N_3545,N_3329,N_3446);
xor U3546 (N_3546,N_3466,N_3459);
or U3547 (N_3547,N_3443,N_3400);
and U3548 (N_3548,N_3387,N_3263);
nor U3549 (N_3549,N_3335,N_3315);
and U3550 (N_3550,N_3252,N_3364);
xnor U3551 (N_3551,N_3260,N_3257);
nand U3552 (N_3552,N_3258,N_3496);
or U3553 (N_3553,N_3304,N_3371);
nor U3554 (N_3554,N_3394,N_3430);
nand U3555 (N_3555,N_3494,N_3328);
xnor U3556 (N_3556,N_3412,N_3276);
nor U3557 (N_3557,N_3407,N_3436);
nor U3558 (N_3558,N_3255,N_3311);
and U3559 (N_3559,N_3467,N_3259);
and U3560 (N_3560,N_3429,N_3444);
xnor U3561 (N_3561,N_3299,N_3416);
and U3562 (N_3562,N_3361,N_3456);
xnor U3563 (N_3563,N_3409,N_3439);
nand U3564 (N_3564,N_3482,N_3272);
or U3565 (N_3565,N_3288,N_3423);
xnor U3566 (N_3566,N_3386,N_3473);
nand U3567 (N_3567,N_3267,N_3441);
and U3568 (N_3568,N_3294,N_3368);
or U3569 (N_3569,N_3389,N_3270);
xnor U3570 (N_3570,N_3485,N_3484);
nor U3571 (N_3571,N_3301,N_3471);
and U3572 (N_3572,N_3379,N_3392);
xor U3573 (N_3573,N_3396,N_3472);
nand U3574 (N_3574,N_3349,N_3492);
nor U3575 (N_3575,N_3497,N_3408);
nor U3576 (N_3576,N_3327,N_3268);
nor U3577 (N_3577,N_3284,N_3480);
xnor U3578 (N_3578,N_3381,N_3380);
nand U3579 (N_3579,N_3293,N_3290);
or U3580 (N_3580,N_3262,N_3424);
and U3581 (N_3581,N_3298,N_3447);
nand U3582 (N_3582,N_3306,N_3498);
nand U3583 (N_3583,N_3321,N_3316);
nand U3584 (N_3584,N_3366,N_3278);
and U3585 (N_3585,N_3338,N_3406);
and U3586 (N_3586,N_3403,N_3251);
nand U3587 (N_3587,N_3341,N_3332);
nand U3588 (N_3588,N_3351,N_3476);
nand U3589 (N_3589,N_3343,N_3344);
xnor U3590 (N_3590,N_3438,N_3488);
xnor U3591 (N_3591,N_3388,N_3486);
nor U3592 (N_3592,N_3282,N_3418);
and U3593 (N_3593,N_3426,N_3457);
or U3594 (N_3594,N_3399,N_3310);
and U3595 (N_3595,N_3420,N_3401);
nand U3596 (N_3596,N_3372,N_3256);
xnor U3597 (N_3597,N_3352,N_3468);
or U3598 (N_3598,N_3397,N_3253);
and U3599 (N_3599,N_3336,N_3261);
nor U3600 (N_3600,N_3451,N_3295);
nor U3601 (N_3601,N_3269,N_3339);
or U3602 (N_3602,N_3474,N_3314);
xor U3603 (N_3603,N_3369,N_3450);
or U3604 (N_3604,N_3281,N_3323);
xor U3605 (N_3605,N_3469,N_3362);
or U3606 (N_3606,N_3452,N_3385);
or U3607 (N_3607,N_3273,N_3413);
or U3608 (N_3608,N_3483,N_3375);
and U3609 (N_3609,N_3275,N_3448);
nand U3610 (N_3610,N_3342,N_3382);
or U3611 (N_3611,N_3395,N_3390);
nor U3612 (N_3612,N_3431,N_3359);
nand U3613 (N_3613,N_3319,N_3365);
nand U3614 (N_3614,N_3414,N_3378);
and U3615 (N_3615,N_3325,N_3404);
or U3616 (N_3616,N_3370,N_3478);
and U3617 (N_3617,N_3312,N_3460);
or U3618 (N_3618,N_3499,N_3461);
or U3619 (N_3619,N_3465,N_3326);
and U3620 (N_3620,N_3417,N_3340);
and U3621 (N_3621,N_3317,N_3458);
nor U3622 (N_3622,N_3383,N_3470);
and U3623 (N_3623,N_3437,N_3313);
xor U3624 (N_3624,N_3330,N_3433);
xor U3625 (N_3625,N_3351,N_3462);
xnor U3626 (N_3626,N_3433,N_3378);
xnor U3627 (N_3627,N_3448,N_3359);
xnor U3628 (N_3628,N_3320,N_3433);
nand U3629 (N_3629,N_3438,N_3443);
or U3630 (N_3630,N_3274,N_3331);
xnor U3631 (N_3631,N_3307,N_3446);
nor U3632 (N_3632,N_3268,N_3497);
xnor U3633 (N_3633,N_3451,N_3433);
or U3634 (N_3634,N_3382,N_3420);
or U3635 (N_3635,N_3386,N_3272);
nor U3636 (N_3636,N_3383,N_3278);
or U3637 (N_3637,N_3317,N_3275);
xor U3638 (N_3638,N_3431,N_3486);
nand U3639 (N_3639,N_3350,N_3442);
nand U3640 (N_3640,N_3317,N_3478);
and U3641 (N_3641,N_3383,N_3368);
xor U3642 (N_3642,N_3364,N_3411);
nor U3643 (N_3643,N_3312,N_3339);
nor U3644 (N_3644,N_3295,N_3362);
nand U3645 (N_3645,N_3486,N_3255);
or U3646 (N_3646,N_3327,N_3424);
and U3647 (N_3647,N_3376,N_3312);
and U3648 (N_3648,N_3391,N_3435);
nor U3649 (N_3649,N_3467,N_3422);
and U3650 (N_3650,N_3341,N_3364);
or U3651 (N_3651,N_3318,N_3379);
and U3652 (N_3652,N_3438,N_3468);
nor U3653 (N_3653,N_3343,N_3289);
nor U3654 (N_3654,N_3379,N_3430);
xor U3655 (N_3655,N_3467,N_3460);
nand U3656 (N_3656,N_3397,N_3295);
and U3657 (N_3657,N_3427,N_3351);
xnor U3658 (N_3658,N_3303,N_3373);
xor U3659 (N_3659,N_3332,N_3300);
or U3660 (N_3660,N_3372,N_3415);
and U3661 (N_3661,N_3489,N_3262);
or U3662 (N_3662,N_3362,N_3391);
and U3663 (N_3663,N_3308,N_3473);
and U3664 (N_3664,N_3304,N_3328);
or U3665 (N_3665,N_3279,N_3430);
nor U3666 (N_3666,N_3436,N_3424);
nor U3667 (N_3667,N_3286,N_3253);
and U3668 (N_3668,N_3304,N_3394);
nand U3669 (N_3669,N_3431,N_3305);
and U3670 (N_3670,N_3353,N_3264);
or U3671 (N_3671,N_3289,N_3344);
and U3672 (N_3672,N_3325,N_3343);
or U3673 (N_3673,N_3386,N_3356);
or U3674 (N_3674,N_3310,N_3451);
nand U3675 (N_3675,N_3412,N_3297);
xor U3676 (N_3676,N_3320,N_3452);
or U3677 (N_3677,N_3413,N_3261);
nor U3678 (N_3678,N_3492,N_3365);
nor U3679 (N_3679,N_3336,N_3257);
xnor U3680 (N_3680,N_3447,N_3336);
xor U3681 (N_3681,N_3453,N_3429);
and U3682 (N_3682,N_3291,N_3321);
nand U3683 (N_3683,N_3363,N_3302);
or U3684 (N_3684,N_3323,N_3292);
and U3685 (N_3685,N_3490,N_3459);
or U3686 (N_3686,N_3370,N_3303);
nand U3687 (N_3687,N_3479,N_3251);
or U3688 (N_3688,N_3488,N_3305);
nor U3689 (N_3689,N_3276,N_3431);
or U3690 (N_3690,N_3466,N_3433);
xor U3691 (N_3691,N_3341,N_3425);
nor U3692 (N_3692,N_3459,N_3434);
nand U3693 (N_3693,N_3363,N_3494);
and U3694 (N_3694,N_3498,N_3291);
nor U3695 (N_3695,N_3285,N_3318);
xor U3696 (N_3696,N_3366,N_3307);
nor U3697 (N_3697,N_3398,N_3483);
and U3698 (N_3698,N_3419,N_3342);
nand U3699 (N_3699,N_3458,N_3483);
and U3700 (N_3700,N_3397,N_3258);
nand U3701 (N_3701,N_3370,N_3277);
or U3702 (N_3702,N_3422,N_3323);
nand U3703 (N_3703,N_3261,N_3293);
nand U3704 (N_3704,N_3453,N_3421);
and U3705 (N_3705,N_3466,N_3444);
nand U3706 (N_3706,N_3311,N_3395);
or U3707 (N_3707,N_3464,N_3384);
nor U3708 (N_3708,N_3441,N_3350);
nand U3709 (N_3709,N_3419,N_3404);
and U3710 (N_3710,N_3356,N_3498);
xnor U3711 (N_3711,N_3262,N_3471);
and U3712 (N_3712,N_3380,N_3497);
xor U3713 (N_3713,N_3324,N_3361);
nand U3714 (N_3714,N_3417,N_3299);
nand U3715 (N_3715,N_3292,N_3400);
xor U3716 (N_3716,N_3369,N_3372);
and U3717 (N_3717,N_3348,N_3306);
or U3718 (N_3718,N_3402,N_3333);
and U3719 (N_3719,N_3457,N_3262);
and U3720 (N_3720,N_3349,N_3498);
xnor U3721 (N_3721,N_3472,N_3330);
and U3722 (N_3722,N_3438,N_3465);
xnor U3723 (N_3723,N_3440,N_3340);
xnor U3724 (N_3724,N_3336,N_3357);
and U3725 (N_3725,N_3289,N_3356);
and U3726 (N_3726,N_3342,N_3336);
xnor U3727 (N_3727,N_3452,N_3498);
or U3728 (N_3728,N_3331,N_3412);
or U3729 (N_3729,N_3276,N_3266);
and U3730 (N_3730,N_3429,N_3477);
and U3731 (N_3731,N_3268,N_3376);
xnor U3732 (N_3732,N_3304,N_3494);
xnor U3733 (N_3733,N_3353,N_3476);
xor U3734 (N_3734,N_3262,N_3452);
and U3735 (N_3735,N_3394,N_3416);
nor U3736 (N_3736,N_3445,N_3275);
xor U3737 (N_3737,N_3358,N_3426);
xnor U3738 (N_3738,N_3273,N_3488);
nand U3739 (N_3739,N_3456,N_3296);
and U3740 (N_3740,N_3299,N_3348);
nand U3741 (N_3741,N_3357,N_3383);
xor U3742 (N_3742,N_3271,N_3338);
xor U3743 (N_3743,N_3337,N_3465);
nor U3744 (N_3744,N_3421,N_3319);
xnor U3745 (N_3745,N_3333,N_3288);
nand U3746 (N_3746,N_3452,N_3451);
or U3747 (N_3747,N_3335,N_3484);
xor U3748 (N_3748,N_3469,N_3496);
or U3749 (N_3749,N_3427,N_3289);
xor U3750 (N_3750,N_3542,N_3587);
or U3751 (N_3751,N_3661,N_3696);
nand U3752 (N_3752,N_3613,N_3599);
or U3753 (N_3753,N_3703,N_3510);
xor U3754 (N_3754,N_3736,N_3645);
or U3755 (N_3755,N_3611,N_3697);
or U3756 (N_3756,N_3671,N_3530);
and U3757 (N_3757,N_3676,N_3614);
or U3758 (N_3758,N_3602,N_3648);
nand U3759 (N_3759,N_3529,N_3742);
xor U3760 (N_3760,N_3543,N_3695);
and U3761 (N_3761,N_3655,N_3709);
xor U3762 (N_3762,N_3501,N_3535);
or U3763 (N_3763,N_3739,N_3679);
nand U3764 (N_3764,N_3660,N_3749);
or U3765 (N_3765,N_3719,N_3634);
nand U3766 (N_3766,N_3615,N_3647);
nand U3767 (N_3767,N_3629,N_3511);
and U3768 (N_3768,N_3564,N_3650);
nand U3769 (N_3769,N_3522,N_3507);
and U3770 (N_3770,N_3681,N_3637);
or U3771 (N_3771,N_3576,N_3536);
xor U3772 (N_3772,N_3571,N_3577);
xnor U3773 (N_3773,N_3603,N_3627);
and U3774 (N_3774,N_3624,N_3531);
and U3775 (N_3775,N_3512,N_3705);
nor U3776 (N_3776,N_3714,N_3636);
nor U3777 (N_3777,N_3688,N_3666);
nor U3778 (N_3778,N_3517,N_3509);
xor U3779 (N_3779,N_3644,N_3580);
xor U3780 (N_3780,N_3523,N_3560);
xnor U3781 (N_3781,N_3566,N_3622);
nand U3782 (N_3782,N_3534,N_3693);
xnor U3783 (N_3783,N_3584,N_3539);
nand U3784 (N_3784,N_3582,N_3735);
nor U3785 (N_3785,N_3589,N_3658);
xnor U3786 (N_3786,N_3659,N_3569);
xor U3787 (N_3787,N_3585,N_3649);
or U3788 (N_3788,N_3716,N_3675);
nor U3789 (N_3789,N_3712,N_3729);
nor U3790 (N_3790,N_3557,N_3654);
and U3791 (N_3791,N_3707,N_3575);
or U3792 (N_3792,N_3640,N_3626);
nand U3793 (N_3793,N_3653,N_3711);
xor U3794 (N_3794,N_3718,N_3593);
xnor U3795 (N_3795,N_3521,N_3673);
and U3796 (N_3796,N_3638,N_3746);
nor U3797 (N_3797,N_3672,N_3607);
nand U3798 (N_3798,N_3595,N_3568);
nand U3799 (N_3799,N_3664,N_3702);
xnor U3800 (N_3800,N_3533,N_3694);
xor U3801 (N_3801,N_3528,N_3670);
and U3802 (N_3802,N_3631,N_3601);
nand U3803 (N_3803,N_3706,N_3741);
nor U3804 (N_3804,N_3724,N_3728);
and U3805 (N_3805,N_3594,N_3731);
or U3806 (N_3806,N_3565,N_3526);
or U3807 (N_3807,N_3605,N_3617);
nand U3808 (N_3808,N_3723,N_3691);
or U3809 (N_3809,N_3633,N_3646);
nand U3810 (N_3810,N_3684,N_3727);
nand U3811 (N_3811,N_3733,N_3537);
xor U3812 (N_3812,N_3540,N_3532);
or U3813 (N_3813,N_3516,N_3726);
nor U3814 (N_3814,N_3692,N_3685);
and U3815 (N_3815,N_3596,N_3620);
nor U3816 (N_3816,N_3721,N_3725);
nor U3817 (N_3817,N_3553,N_3519);
nor U3818 (N_3818,N_3588,N_3551);
nor U3819 (N_3819,N_3583,N_3518);
nor U3820 (N_3820,N_3738,N_3630);
or U3821 (N_3821,N_3687,N_3698);
xnor U3822 (N_3822,N_3642,N_3690);
nor U3823 (N_3823,N_3545,N_3722);
xor U3824 (N_3824,N_3546,N_3515);
or U3825 (N_3825,N_3668,N_3682);
xnor U3826 (N_3826,N_3561,N_3678);
nand U3827 (N_3827,N_3683,N_3541);
nor U3828 (N_3828,N_3552,N_3555);
nand U3829 (N_3829,N_3639,N_3563);
nand U3830 (N_3830,N_3700,N_3732);
nor U3831 (N_3831,N_3740,N_3701);
or U3832 (N_3832,N_3667,N_3548);
xnor U3833 (N_3833,N_3503,N_3710);
or U3834 (N_3834,N_3635,N_3610);
xnor U3835 (N_3835,N_3651,N_3656);
and U3836 (N_3836,N_3674,N_3665);
nand U3837 (N_3837,N_3504,N_3717);
xnor U3838 (N_3838,N_3554,N_3598);
xnor U3839 (N_3839,N_3556,N_3748);
and U3840 (N_3840,N_3559,N_3558);
and U3841 (N_3841,N_3500,N_3715);
xor U3842 (N_3842,N_3520,N_3618);
or U3843 (N_3843,N_3708,N_3669);
nor U3844 (N_3844,N_3689,N_3734);
and U3845 (N_3845,N_3527,N_3621);
nor U3846 (N_3846,N_3704,N_3567);
or U3847 (N_3847,N_3525,N_3606);
or U3848 (N_3848,N_3609,N_3597);
nor U3849 (N_3849,N_3513,N_3506);
or U3850 (N_3850,N_3744,N_3590);
xnor U3851 (N_3851,N_3604,N_3573);
or U3852 (N_3852,N_3547,N_3544);
nor U3853 (N_3853,N_3608,N_3619);
xnor U3854 (N_3854,N_3502,N_3730);
or U3855 (N_3855,N_3680,N_3737);
and U3856 (N_3856,N_3745,N_3549);
nand U3857 (N_3857,N_3628,N_3586);
or U3858 (N_3858,N_3747,N_3643);
xor U3859 (N_3859,N_3600,N_3538);
xor U3860 (N_3860,N_3578,N_3612);
nor U3861 (N_3861,N_3625,N_3657);
nor U3862 (N_3862,N_3699,N_3570);
and U3863 (N_3863,N_3572,N_3508);
nor U3864 (N_3864,N_3686,N_3505);
nor U3865 (N_3865,N_3514,N_3743);
nand U3866 (N_3866,N_3623,N_3592);
nor U3867 (N_3867,N_3581,N_3652);
nor U3868 (N_3868,N_3677,N_3641);
or U3869 (N_3869,N_3562,N_3713);
or U3870 (N_3870,N_3663,N_3579);
and U3871 (N_3871,N_3524,N_3591);
and U3872 (N_3872,N_3720,N_3550);
nand U3873 (N_3873,N_3574,N_3632);
or U3874 (N_3874,N_3662,N_3616);
xnor U3875 (N_3875,N_3734,N_3507);
nor U3876 (N_3876,N_3694,N_3743);
and U3877 (N_3877,N_3606,N_3679);
or U3878 (N_3878,N_3600,N_3730);
nor U3879 (N_3879,N_3707,N_3515);
nand U3880 (N_3880,N_3665,N_3515);
and U3881 (N_3881,N_3575,N_3565);
xnor U3882 (N_3882,N_3685,N_3739);
or U3883 (N_3883,N_3509,N_3626);
nor U3884 (N_3884,N_3530,N_3564);
or U3885 (N_3885,N_3548,N_3553);
and U3886 (N_3886,N_3546,N_3738);
nand U3887 (N_3887,N_3612,N_3531);
nand U3888 (N_3888,N_3624,N_3622);
and U3889 (N_3889,N_3621,N_3548);
xor U3890 (N_3890,N_3511,N_3555);
or U3891 (N_3891,N_3596,N_3567);
or U3892 (N_3892,N_3507,N_3662);
and U3893 (N_3893,N_3694,N_3741);
or U3894 (N_3894,N_3512,N_3572);
or U3895 (N_3895,N_3613,N_3501);
or U3896 (N_3896,N_3572,N_3621);
xor U3897 (N_3897,N_3582,N_3741);
nor U3898 (N_3898,N_3557,N_3640);
or U3899 (N_3899,N_3615,N_3668);
and U3900 (N_3900,N_3676,N_3707);
nand U3901 (N_3901,N_3569,N_3574);
and U3902 (N_3902,N_3622,N_3541);
nor U3903 (N_3903,N_3717,N_3513);
nand U3904 (N_3904,N_3562,N_3538);
xnor U3905 (N_3905,N_3652,N_3714);
or U3906 (N_3906,N_3546,N_3540);
and U3907 (N_3907,N_3687,N_3529);
nor U3908 (N_3908,N_3690,N_3520);
or U3909 (N_3909,N_3671,N_3545);
nor U3910 (N_3910,N_3735,N_3586);
or U3911 (N_3911,N_3655,N_3725);
xor U3912 (N_3912,N_3602,N_3732);
or U3913 (N_3913,N_3701,N_3598);
nor U3914 (N_3914,N_3578,N_3744);
nor U3915 (N_3915,N_3550,N_3608);
xor U3916 (N_3916,N_3672,N_3557);
xor U3917 (N_3917,N_3616,N_3501);
nand U3918 (N_3918,N_3519,N_3563);
xnor U3919 (N_3919,N_3713,N_3749);
nand U3920 (N_3920,N_3728,N_3602);
or U3921 (N_3921,N_3660,N_3614);
xor U3922 (N_3922,N_3560,N_3592);
nand U3923 (N_3923,N_3549,N_3576);
nor U3924 (N_3924,N_3695,N_3618);
nor U3925 (N_3925,N_3547,N_3643);
or U3926 (N_3926,N_3691,N_3635);
and U3927 (N_3927,N_3630,N_3523);
nand U3928 (N_3928,N_3508,N_3571);
nor U3929 (N_3929,N_3649,N_3620);
xor U3930 (N_3930,N_3739,N_3527);
and U3931 (N_3931,N_3693,N_3578);
xor U3932 (N_3932,N_3545,N_3527);
or U3933 (N_3933,N_3717,N_3575);
or U3934 (N_3934,N_3733,N_3569);
nor U3935 (N_3935,N_3552,N_3734);
or U3936 (N_3936,N_3533,N_3674);
or U3937 (N_3937,N_3668,N_3613);
nand U3938 (N_3938,N_3550,N_3669);
or U3939 (N_3939,N_3514,N_3500);
nand U3940 (N_3940,N_3665,N_3673);
nor U3941 (N_3941,N_3668,N_3585);
or U3942 (N_3942,N_3674,N_3737);
or U3943 (N_3943,N_3617,N_3660);
nand U3944 (N_3944,N_3652,N_3531);
xor U3945 (N_3945,N_3592,N_3635);
nor U3946 (N_3946,N_3516,N_3547);
and U3947 (N_3947,N_3526,N_3635);
or U3948 (N_3948,N_3616,N_3695);
or U3949 (N_3949,N_3696,N_3616);
xor U3950 (N_3950,N_3608,N_3591);
nand U3951 (N_3951,N_3590,N_3692);
nand U3952 (N_3952,N_3704,N_3561);
or U3953 (N_3953,N_3661,N_3676);
or U3954 (N_3954,N_3526,N_3569);
or U3955 (N_3955,N_3517,N_3722);
nor U3956 (N_3956,N_3513,N_3522);
nor U3957 (N_3957,N_3506,N_3594);
nand U3958 (N_3958,N_3599,N_3521);
and U3959 (N_3959,N_3617,N_3667);
and U3960 (N_3960,N_3541,N_3728);
and U3961 (N_3961,N_3736,N_3738);
xnor U3962 (N_3962,N_3744,N_3602);
nand U3963 (N_3963,N_3680,N_3608);
nor U3964 (N_3964,N_3693,N_3722);
nor U3965 (N_3965,N_3626,N_3737);
nand U3966 (N_3966,N_3536,N_3515);
xnor U3967 (N_3967,N_3665,N_3716);
xor U3968 (N_3968,N_3559,N_3576);
nor U3969 (N_3969,N_3651,N_3502);
and U3970 (N_3970,N_3645,N_3699);
or U3971 (N_3971,N_3543,N_3722);
nor U3972 (N_3972,N_3584,N_3536);
and U3973 (N_3973,N_3721,N_3618);
nor U3974 (N_3974,N_3695,N_3620);
nor U3975 (N_3975,N_3688,N_3534);
nand U3976 (N_3976,N_3746,N_3525);
nand U3977 (N_3977,N_3740,N_3680);
and U3978 (N_3978,N_3658,N_3619);
and U3979 (N_3979,N_3555,N_3594);
xnor U3980 (N_3980,N_3573,N_3744);
nor U3981 (N_3981,N_3578,N_3548);
or U3982 (N_3982,N_3741,N_3730);
nor U3983 (N_3983,N_3701,N_3514);
or U3984 (N_3984,N_3536,N_3645);
or U3985 (N_3985,N_3599,N_3522);
nand U3986 (N_3986,N_3637,N_3590);
xor U3987 (N_3987,N_3725,N_3575);
or U3988 (N_3988,N_3525,N_3716);
nand U3989 (N_3989,N_3606,N_3624);
nor U3990 (N_3990,N_3650,N_3511);
and U3991 (N_3991,N_3546,N_3712);
xor U3992 (N_3992,N_3707,N_3614);
nor U3993 (N_3993,N_3504,N_3644);
and U3994 (N_3994,N_3739,N_3601);
xnor U3995 (N_3995,N_3661,N_3720);
or U3996 (N_3996,N_3643,N_3657);
nand U3997 (N_3997,N_3652,N_3738);
or U3998 (N_3998,N_3546,N_3656);
xor U3999 (N_3999,N_3740,N_3500);
xnor U4000 (N_4000,N_3944,N_3975);
xnor U4001 (N_4001,N_3750,N_3957);
and U4002 (N_4002,N_3946,N_3877);
and U4003 (N_4003,N_3780,N_3829);
nor U4004 (N_4004,N_3866,N_3755);
nand U4005 (N_4005,N_3800,N_3852);
nand U4006 (N_4006,N_3831,N_3867);
xnor U4007 (N_4007,N_3931,N_3835);
and U4008 (N_4008,N_3954,N_3865);
nor U4009 (N_4009,N_3897,N_3970);
and U4010 (N_4010,N_3887,N_3815);
xor U4011 (N_4011,N_3996,N_3777);
nor U4012 (N_4012,N_3804,N_3870);
and U4013 (N_4013,N_3979,N_3905);
nand U4014 (N_4014,N_3952,N_3994);
nor U4015 (N_4015,N_3774,N_3768);
nor U4016 (N_4016,N_3837,N_3767);
nand U4017 (N_4017,N_3834,N_3909);
or U4018 (N_4018,N_3825,N_3960);
nor U4019 (N_4019,N_3933,N_3809);
xor U4020 (N_4020,N_3964,N_3941);
xnor U4021 (N_4021,N_3935,N_3902);
xnor U4022 (N_4022,N_3971,N_3851);
or U4023 (N_4023,N_3788,N_3930);
nor U4024 (N_4024,N_3812,N_3885);
nor U4025 (N_4025,N_3886,N_3983);
xor U4026 (N_4026,N_3982,N_3875);
nor U4027 (N_4027,N_3816,N_3791);
xor U4028 (N_4028,N_3758,N_3951);
nand U4029 (N_4029,N_3969,N_3919);
nor U4030 (N_4030,N_3890,N_3936);
xor U4031 (N_4031,N_3943,N_3832);
and U4032 (N_4032,N_3784,N_3923);
and U4033 (N_4033,N_3911,N_3989);
or U4034 (N_4034,N_3843,N_3786);
xor U4035 (N_4035,N_3908,N_3904);
nand U4036 (N_4036,N_3918,N_3797);
nand U4037 (N_4037,N_3949,N_3836);
or U4038 (N_4038,N_3795,N_3962);
and U4039 (N_4039,N_3891,N_3848);
nand U4040 (N_4040,N_3820,N_3956);
and U4041 (N_4041,N_3880,N_3775);
nand U4042 (N_4042,N_3789,N_3817);
xnor U4043 (N_4043,N_3916,N_3929);
nor U4044 (N_4044,N_3760,N_3999);
nor U4045 (N_4045,N_3871,N_3756);
xnor U4046 (N_4046,N_3798,N_3819);
or U4047 (N_4047,N_3861,N_3910);
nand U4048 (N_4048,N_3781,N_3850);
nor U4049 (N_4049,N_3934,N_3938);
nand U4050 (N_4050,N_3882,N_3922);
nor U4051 (N_4051,N_3892,N_3813);
nand U4052 (N_4052,N_3940,N_3811);
or U4053 (N_4053,N_3828,N_3972);
or U4054 (N_4054,N_3839,N_3876);
xor U4055 (N_4055,N_3894,N_3937);
xor U4056 (N_4056,N_3821,N_3921);
nor U4057 (N_4057,N_3898,N_3939);
nor U4058 (N_4058,N_3782,N_3808);
nand U4059 (N_4059,N_3805,N_3776);
and U4060 (N_4060,N_3846,N_3984);
and U4061 (N_4061,N_3823,N_3783);
or U4062 (N_4062,N_3754,N_3874);
and U4063 (N_4063,N_3751,N_3945);
or U4064 (N_4064,N_3925,N_3796);
and U4065 (N_4065,N_3790,N_3822);
and U4066 (N_4066,N_3947,N_3833);
or U4067 (N_4067,N_3906,N_3967);
xor U4068 (N_4068,N_3872,N_3857);
nor U4069 (N_4069,N_3824,N_3987);
nand U4070 (N_4070,N_3860,N_3966);
nand U4071 (N_4071,N_3985,N_3842);
and U4072 (N_4072,N_3993,N_3927);
or U4073 (N_4073,N_3968,N_3903);
nand U4074 (N_4074,N_3988,N_3838);
nand U4075 (N_4075,N_3879,N_3849);
nand U4076 (N_4076,N_3978,N_3818);
nor U4077 (N_4077,N_3868,N_3873);
or U4078 (N_4078,N_3765,N_3763);
or U4079 (N_4079,N_3884,N_3974);
xor U4080 (N_4080,N_3965,N_3840);
nor U4081 (N_4081,N_3853,N_3787);
and U4082 (N_4082,N_3963,N_3883);
xnor U4083 (N_4083,N_3948,N_3900);
nand U4084 (N_4084,N_3864,N_3863);
or U4085 (N_4085,N_3926,N_3955);
and U4086 (N_4086,N_3771,N_3830);
nand U4087 (N_4087,N_3973,N_3827);
nand U4088 (N_4088,N_3757,N_3913);
or U4089 (N_4089,N_3761,N_3907);
nand U4090 (N_4090,N_3990,N_3998);
nor U4091 (N_4091,N_3770,N_3924);
nor U4092 (N_4092,N_3893,N_3792);
or U4093 (N_4093,N_3901,N_3814);
nand U4094 (N_4094,N_3992,N_3766);
nor U4095 (N_4095,N_3912,N_3959);
xnor U4096 (N_4096,N_3881,N_3802);
and U4097 (N_4097,N_3810,N_3844);
or U4098 (N_4098,N_3759,N_3845);
xor U4099 (N_4099,N_3855,N_3961);
or U4100 (N_4100,N_3779,N_3801);
xnor U4101 (N_4101,N_3793,N_3799);
and U4102 (N_4102,N_3878,N_3914);
nor U4103 (N_4103,N_3895,N_3807);
nand U4104 (N_4104,N_3991,N_3856);
or U4105 (N_4105,N_3826,N_3862);
nor U4106 (N_4106,N_3806,N_3977);
xnor U4107 (N_4107,N_3803,N_3764);
nor U4108 (N_4108,N_3847,N_3942);
and U4109 (N_4109,N_3976,N_3995);
or U4110 (N_4110,N_3888,N_3772);
xor U4111 (N_4111,N_3986,N_3785);
nand U4112 (N_4112,N_3752,N_3981);
or U4113 (N_4113,N_3896,N_3932);
nand U4114 (N_4114,N_3778,N_3915);
xnor U4115 (N_4115,N_3950,N_3928);
and U4116 (N_4116,N_3997,N_3917);
nor U4117 (N_4117,N_3889,N_3869);
or U4118 (N_4118,N_3773,N_3920);
or U4119 (N_4119,N_3858,N_3762);
and U4120 (N_4120,N_3841,N_3753);
nor U4121 (N_4121,N_3958,N_3794);
xor U4122 (N_4122,N_3899,N_3854);
xor U4123 (N_4123,N_3980,N_3769);
and U4124 (N_4124,N_3953,N_3859);
nand U4125 (N_4125,N_3811,N_3873);
xnor U4126 (N_4126,N_3943,N_3912);
xnor U4127 (N_4127,N_3919,N_3928);
nand U4128 (N_4128,N_3767,N_3829);
nor U4129 (N_4129,N_3918,N_3858);
nand U4130 (N_4130,N_3886,N_3993);
nor U4131 (N_4131,N_3998,N_3908);
or U4132 (N_4132,N_3956,N_3761);
nand U4133 (N_4133,N_3791,N_3981);
xor U4134 (N_4134,N_3987,N_3945);
nand U4135 (N_4135,N_3839,N_3798);
xnor U4136 (N_4136,N_3949,N_3975);
xor U4137 (N_4137,N_3785,N_3881);
and U4138 (N_4138,N_3777,N_3920);
nand U4139 (N_4139,N_3943,N_3858);
xor U4140 (N_4140,N_3825,N_3979);
and U4141 (N_4141,N_3798,N_3939);
xnor U4142 (N_4142,N_3784,N_3762);
and U4143 (N_4143,N_3835,N_3853);
xnor U4144 (N_4144,N_3774,N_3927);
and U4145 (N_4145,N_3890,N_3873);
nand U4146 (N_4146,N_3880,N_3789);
and U4147 (N_4147,N_3881,N_3843);
and U4148 (N_4148,N_3888,N_3947);
or U4149 (N_4149,N_3917,N_3927);
or U4150 (N_4150,N_3778,N_3994);
or U4151 (N_4151,N_3765,N_3986);
nand U4152 (N_4152,N_3910,N_3996);
and U4153 (N_4153,N_3814,N_3866);
nand U4154 (N_4154,N_3841,N_3889);
nor U4155 (N_4155,N_3998,N_3979);
nand U4156 (N_4156,N_3801,N_3777);
nand U4157 (N_4157,N_3999,N_3931);
nor U4158 (N_4158,N_3907,N_3814);
xnor U4159 (N_4159,N_3958,N_3912);
nor U4160 (N_4160,N_3837,N_3954);
xnor U4161 (N_4161,N_3806,N_3905);
and U4162 (N_4162,N_3776,N_3886);
nand U4163 (N_4163,N_3840,N_3851);
xor U4164 (N_4164,N_3941,N_3922);
and U4165 (N_4165,N_3843,N_3768);
and U4166 (N_4166,N_3760,N_3974);
nand U4167 (N_4167,N_3914,N_3999);
nor U4168 (N_4168,N_3823,N_3787);
or U4169 (N_4169,N_3867,N_3995);
and U4170 (N_4170,N_3951,N_3801);
or U4171 (N_4171,N_3988,N_3828);
xnor U4172 (N_4172,N_3991,N_3899);
nand U4173 (N_4173,N_3887,N_3866);
nand U4174 (N_4174,N_3940,N_3920);
nor U4175 (N_4175,N_3830,N_3766);
nand U4176 (N_4176,N_3907,N_3781);
or U4177 (N_4177,N_3951,N_3765);
nor U4178 (N_4178,N_3878,N_3761);
nand U4179 (N_4179,N_3868,N_3818);
xor U4180 (N_4180,N_3815,N_3751);
xnor U4181 (N_4181,N_3998,N_3835);
nor U4182 (N_4182,N_3774,N_3946);
xnor U4183 (N_4183,N_3751,N_3870);
or U4184 (N_4184,N_3790,N_3936);
or U4185 (N_4185,N_3751,N_3795);
nand U4186 (N_4186,N_3943,N_3907);
xor U4187 (N_4187,N_3845,N_3890);
nand U4188 (N_4188,N_3754,N_3826);
or U4189 (N_4189,N_3883,N_3971);
nand U4190 (N_4190,N_3791,N_3762);
nand U4191 (N_4191,N_3916,N_3827);
nand U4192 (N_4192,N_3976,N_3884);
nor U4193 (N_4193,N_3856,N_3802);
or U4194 (N_4194,N_3768,N_3793);
nand U4195 (N_4195,N_3863,N_3998);
and U4196 (N_4196,N_3873,N_3895);
xnor U4197 (N_4197,N_3975,N_3977);
nand U4198 (N_4198,N_3901,N_3831);
or U4199 (N_4199,N_3820,N_3874);
nor U4200 (N_4200,N_3877,N_3937);
xor U4201 (N_4201,N_3982,N_3766);
nor U4202 (N_4202,N_3802,N_3765);
or U4203 (N_4203,N_3829,N_3956);
nor U4204 (N_4204,N_3965,N_3996);
nand U4205 (N_4205,N_3824,N_3986);
or U4206 (N_4206,N_3828,N_3803);
or U4207 (N_4207,N_3929,N_3788);
nor U4208 (N_4208,N_3958,N_3875);
or U4209 (N_4209,N_3942,N_3990);
nor U4210 (N_4210,N_3813,N_3910);
nor U4211 (N_4211,N_3777,N_3823);
nor U4212 (N_4212,N_3880,N_3930);
and U4213 (N_4213,N_3756,N_3774);
nor U4214 (N_4214,N_3809,N_3934);
or U4215 (N_4215,N_3846,N_3835);
and U4216 (N_4216,N_3768,N_3876);
or U4217 (N_4217,N_3846,N_3865);
or U4218 (N_4218,N_3788,N_3947);
nand U4219 (N_4219,N_3751,N_3975);
or U4220 (N_4220,N_3901,N_3836);
nand U4221 (N_4221,N_3981,N_3991);
xnor U4222 (N_4222,N_3975,N_3971);
nand U4223 (N_4223,N_3804,N_3905);
and U4224 (N_4224,N_3881,N_3782);
xor U4225 (N_4225,N_3810,N_3922);
nand U4226 (N_4226,N_3972,N_3974);
and U4227 (N_4227,N_3942,N_3844);
nor U4228 (N_4228,N_3934,N_3811);
nor U4229 (N_4229,N_3989,N_3820);
and U4230 (N_4230,N_3953,N_3833);
nand U4231 (N_4231,N_3976,N_3867);
and U4232 (N_4232,N_3783,N_3759);
nor U4233 (N_4233,N_3835,N_3868);
or U4234 (N_4234,N_3972,N_3801);
nor U4235 (N_4235,N_3770,N_3781);
xnor U4236 (N_4236,N_3844,N_3979);
nor U4237 (N_4237,N_3901,N_3963);
nand U4238 (N_4238,N_3810,N_3936);
xnor U4239 (N_4239,N_3855,N_3816);
nor U4240 (N_4240,N_3754,N_3890);
or U4241 (N_4241,N_3916,N_3944);
nand U4242 (N_4242,N_3840,N_3787);
nand U4243 (N_4243,N_3918,N_3757);
xnor U4244 (N_4244,N_3925,N_3960);
xnor U4245 (N_4245,N_3973,N_3947);
or U4246 (N_4246,N_3788,N_3851);
or U4247 (N_4247,N_3765,N_3798);
nand U4248 (N_4248,N_3772,N_3877);
nand U4249 (N_4249,N_3808,N_3935);
or U4250 (N_4250,N_4003,N_4153);
and U4251 (N_4251,N_4127,N_4006);
and U4252 (N_4252,N_4130,N_4134);
or U4253 (N_4253,N_4037,N_4043);
xnor U4254 (N_4254,N_4107,N_4116);
xor U4255 (N_4255,N_4243,N_4149);
nand U4256 (N_4256,N_4102,N_4217);
or U4257 (N_4257,N_4060,N_4146);
nand U4258 (N_4258,N_4161,N_4052);
or U4259 (N_4259,N_4123,N_4084);
xnor U4260 (N_4260,N_4183,N_4030);
xnor U4261 (N_4261,N_4168,N_4198);
nand U4262 (N_4262,N_4209,N_4128);
or U4263 (N_4263,N_4109,N_4223);
and U4264 (N_4264,N_4176,N_4119);
or U4265 (N_4265,N_4141,N_4036);
nand U4266 (N_4266,N_4182,N_4186);
xnor U4267 (N_4267,N_4103,N_4154);
or U4268 (N_4268,N_4048,N_4051);
and U4269 (N_4269,N_4234,N_4246);
or U4270 (N_4270,N_4118,N_4108);
nor U4271 (N_4271,N_4025,N_4180);
nand U4272 (N_4272,N_4171,N_4053);
nand U4273 (N_4273,N_4095,N_4063);
or U4274 (N_4274,N_4150,N_4225);
nor U4275 (N_4275,N_4111,N_4142);
xor U4276 (N_4276,N_4078,N_4069);
nand U4277 (N_4277,N_4211,N_4214);
or U4278 (N_4278,N_4086,N_4055);
and U4279 (N_4279,N_4148,N_4206);
and U4280 (N_4280,N_4028,N_4241);
nor U4281 (N_4281,N_4244,N_4188);
nand U4282 (N_4282,N_4210,N_4104);
nand U4283 (N_4283,N_4079,N_4233);
nor U4284 (N_4284,N_4236,N_4085);
or U4285 (N_4285,N_4229,N_4017);
nand U4286 (N_4286,N_4039,N_4219);
nand U4287 (N_4287,N_4100,N_4035);
or U4288 (N_4288,N_4106,N_4167);
nand U4289 (N_4289,N_4073,N_4212);
xnor U4290 (N_4290,N_4092,N_4090);
nor U4291 (N_4291,N_4228,N_4059);
or U4292 (N_4292,N_4170,N_4139);
xor U4293 (N_4293,N_4178,N_4248);
and U4294 (N_4294,N_4164,N_4247);
xnor U4295 (N_4295,N_4125,N_4091);
xor U4296 (N_4296,N_4066,N_4020);
nor U4297 (N_4297,N_4001,N_4213);
xnor U4298 (N_4298,N_4072,N_4221);
and U4299 (N_4299,N_4019,N_4007);
xor U4300 (N_4300,N_4195,N_4207);
and U4301 (N_4301,N_4169,N_4172);
or U4302 (N_4302,N_4094,N_4245);
and U4303 (N_4303,N_4239,N_4013);
nor U4304 (N_4304,N_4181,N_4187);
or U4305 (N_4305,N_4012,N_4158);
and U4306 (N_4306,N_4046,N_4038);
nand U4307 (N_4307,N_4068,N_4041);
nor U4308 (N_4308,N_4065,N_4205);
nand U4309 (N_4309,N_4208,N_4122);
nor U4310 (N_4310,N_4224,N_4157);
and U4311 (N_4311,N_4126,N_4121);
xor U4312 (N_4312,N_4101,N_4216);
nand U4313 (N_4313,N_4004,N_4184);
xor U4314 (N_4314,N_4061,N_4200);
and U4315 (N_4315,N_4238,N_4202);
nor U4316 (N_4316,N_4230,N_4194);
xor U4317 (N_4317,N_4014,N_4031);
xnor U4318 (N_4318,N_4129,N_4049);
or U4319 (N_4319,N_4156,N_4018);
or U4320 (N_4320,N_4016,N_4227);
nand U4321 (N_4321,N_4144,N_4115);
nor U4322 (N_4322,N_4192,N_4147);
and U4323 (N_4323,N_4218,N_4110);
or U4324 (N_4324,N_4005,N_4138);
nor U4325 (N_4325,N_4249,N_4074);
or U4326 (N_4326,N_4056,N_4163);
and U4327 (N_4327,N_4196,N_4026);
nor U4328 (N_4328,N_4098,N_4058);
xor U4329 (N_4329,N_4137,N_4190);
nand U4330 (N_4330,N_4027,N_4050);
xnor U4331 (N_4331,N_4160,N_4132);
and U4332 (N_4332,N_4203,N_4177);
nand U4333 (N_4333,N_4240,N_4226);
nand U4334 (N_4334,N_4075,N_4062);
xnor U4335 (N_4335,N_4159,N_4097);
and U4336 (N_4336,N_4145,N_4002);
and U4337 (N_4337,N_4047,N_4215);
xnor U4338 (N_4338,N_4076,N_4204);
xor U4339 (N_4339,N_4201,N_4189);
nor U4340 (N_4340,N_4023,N_4057);
nor U4341 (N_4341,N_4173,N_4011);
nand U4342 (N_4342,N_4185,N_4193);
and U4343 (N_4343,N_4008,N_4151);
nor U4344 (N_4344,N_4220,N_4237);
xor U4345 (N_4345,N_4174,N_4033);
nor U4346 (N_4346,N_4045,N_4232);
xnor U4347 (N_4347,N_4152,N_4235);
xor U4348 (N_4348,N_4087,N_4136);
or U4349 (N_4349,N_4093,N_4131);
nand U4350 (N_4350,N_4112,N_4175);
nand U4351 (N_4351,N_4222,N_4022);
and U4352 (N_4352,N_4114,N_4088);
nand U4353 (N_4353,N_4140,N_4191);
nor U4354 (N_4354,N_4117,N_4096);
nand U4355 (N_4355,N_4071,N_4162);
and U4356 (N_4356,N_4120,N_4080);
or U4357 (N_4357,N_4099,N_4143);
or U4358 (N_4358,N_4067,N_4044);
and U4359 (N_4359,N_4197,N_4064);
nand U4360 (N_4360,N_4021,N_4070);
nand U4361 (N_4361,N_4089,N_4032);
nand U4362 (N_4362,N_4083,N_4179);
and U4363 (N_4363,N_4166,N_4133);
nand U4364 (N_4364,N_4040,N_4034);
xnor U4365 (N_4365,N_4082,N_4009);
nor U4366 (N_4366,N_4135,N_4042);
nand U4367 (N_4367,N_4024,N_4199);
and U4368 (N_4368,N_4124,N_4165);
and U4369 (N_4369,N_4155,N_4105);
and U4370 (N_4370,N_4000,N_4010);
or U4371 (N_4371,N_4077,N_4015);
nor U4372 (N_4372,N_4081,N_4231);
nor U4373 (N_4373,N_4054,N_4242);
nand U4374 (N_4374,N_4113,N_4029);
nor U4375 (N_4375,N_4016,N_4003);
and U4376 (N_4376,N_4035,N_4161);
nand U4377 (N_4377,N_4211,N_4139);
and U4378 (N_4378,N_4047,N_4010);
or U4379 (N_4379,N_4146,N_4043);
or U4380 (N_4380,N_4231,N_4079);
xor U4381 (N_4381,N_4177,N_4130);
or U4382 (N_4382,N_4018,N_4230);
xor U4383 (N_4383,N_4091,N_4018);
nor U4384 (N_4384,N_4154,N_4024);
and U4385 (N_4385,N_4229,N_4147);
or U4386 (N_4386,N_4040,N_4058);
nand U4387 (N_4387,N_4154,N_4097);
nor U4388 (N_4388,N_4114,N_4068);
nor U4389 (N_4389,N_4044,N_4246);
or U4390 (N_4390,N_4067,N_4235);
nor U4391 (N_4391,N_4191,N_4055);
nand U4392 (N_4392,N_4068,N_4066);
or U4393 (N_4393,N_4138,N_4083);
nand U4394 (N_4394,N_4039,N_4236);
or U4395 (N_4395,N_4021,N_4100);
nand U4396 (N_4396,N_4233,N_4005);
and U4397 (N_4397,N_4121,N_4063);
xor U4398 (N_4398,N_4103,N_4205);
nand U4399 (N_4399,N_4133,N_4242);
and U4400 (N_4400,N_4171,N_4127);
and U4401 (N_4401,N_4194,N_4065);
nor U4402 (N_4402,N_4214,N_4069);
nand U4403 (N_4403,N_4101,N_4228);
and U4404 (N_4404,N_4115,N_4077);
nor U4405 (N_4405,N_4219,N_4062);
or U4406 (N_4406,N_4085,N_4239);
or U4407 (N_4407,N_4232,N_4214);
xor U4408 (N_4408,N_4018,N_4157);
and U4409 (N_4409,N_4078,N_4180);
nor U4410 (N_4410,N_4089,N_4137);
or U4411 (N_4411,N_4178,N_4223);
xor U4412 (N_4412,N_4035,N_4160);
xor U4413 (N_4413,N_4163,N_4239);
or U4414 (N_4414,N_4045,N_4187);
nor U4415 (N_4415,N_4147,N_4176);
xor U4416 (N_4416,N_4144,N_4149);
nand U4417 (N_4417,N_4030,N_4244);
or U4418 (N_4418,N_4186,N_4066);
and U4419 (N_4419,N_4152,N_4075);
nand U4420 (N_4420,N_4214,N_4023);
nand U4421 (N_4421,N_4040,N_4144);
nor U4422 (N_4422,N_4243,N_4136);
nand U4423 (N_4423,N_4123,N_4012);
nand U4424 (N_4424,N_4026,N_4179);
nand U4425 (N_4425,N_4068,N_4073);
and U4426 (N_4426,N_4150,N_4223);
nand U4427 (N_4427,N_4126,N_4245);
xor U4428 (N_4428,N_4059,N_4023);
or U4429 (N_4429,N_4132,N_4081);
or U4430 (N_4430,N_4138,N_4214);
nand U4431 (N_4431,N_4065,N_4032);
or U4432 (N_4432,N_4223,N_4211);
nand U4433 (N_4433,N_4177,N_4009);
and U4434 (N_4434,N_4216,N_4099);
xnor U4435 (N_4435,N_4026,N_4202);
xor U4436 (N_4436,N_4056,N_4033);
nor U4437 (N_4437,N_4138,N_4147);
nor U4438 (N_4438,N_4204,N_4024);
nor U4439 (N_4439,N_4067,N_4228);
xnor U4440 (N_4440,N_4144,N_4212);
nor U4441 (N_4441,N_4159,N_4023);
or U4442 (N_4442,N_4174,N_4125);
nand U4443 (N_4443,N_4116,N_4133);
and U4444 (N_4444,N_4248,N_4213);
nand U4445 (N_4445,N_4071,N_4159);
nand U4446 (N_4446,N_4048,N_4147);
xnor U4447 (N_4447,N_4172,N_4151);
nand U4448 (N_4448,N_4051,N_4019);
xnor U4449 (N_4449,N_4207,N_4185);
nor U4450 (N_4450,N_4146,N_4016);
and U4451 (N_4451,N_4003,N_4071);
or U4452 (N_4452,N_4199,N_4143);
and U4453 (N_4453,N_4030,N_4037);
nor U4454 (N_4454,N_4152,N_4163);
xnor U4455 (N_4455,N_4021,N_4169);
xnor U4456 (N_4456,N_4135,N_4062);
nor U4457 (N_4457,N_4184,N_4089);
xnor U4458 (N_4458,N_4223,N_4004);
xnor U4459 (N_4459,N_4121,N_4057);
xnor U4460 (N_4460,N_4209,N_4239);
and U4461 (N_4461,N_4064,N_4046);
and U4462 (N_4462,N_4020,N_4169);
xnor U4463 (N_4463,N_4153,N_4045);
or U4464 (N_4464,N_4109,N_4073);
and U4465 (N_4465,N_4058,N_4222);
and U4466 (N_4466,N_4032,N_4028);
nand U4467 (N_4467,N_4205,N_4197);
nand U4468 (N_4468,N_4220,N_4188);
and U4469 (N_4469,N_4092,N_4194);
or U4470 (N_4470,N_4069,N_4158);
nand U4471 (N_4471,N_4081,N_4192);
nor U4472 (N_4472,N_4078,N_4087);
nand U4473 (N_4473,N_4126,N_4217);
nand U4474 (N_4474,N_4023,N_4206);
and U4475 (N_4475,N_4019,N_4079);
nand U4476 (N_4476,N_4035,N_4216);
xnor U4477 (N_4477,N_4031,N_4050);
nor U4478 (N_4478,N_4101,N_4010);
or U4479 (N_4479,N_4228,N_4005);
and U4480 (N_4480,N_4196,N_4240);
and U4481 (N_4481,N_4019,N_4168);
nor U4482 (N_4482,N_4077,N_4242);
and U4483 (N_4483,N_4028,N_4177);
nor U4484 (N_4484,N_4162,N_4057);
or U4485 (N_4485,N_4078,N_4113);
xor U4486 (N_4486,N_4158,N_4219);
xnor U4487 (N_4487,N_4009,N_4101);
xnor U4488 (N_4488,N_4020,N_4228);
nor U4489 (N_4489,N_4023,N_4236);
xnor U4490 (N_4490,N_4246,N_4122);
nand U4491 (N_4491,N_4229,N_4129);
and U4492 (N_4492,N_4088,N_4096);
nor U4493 (N_4493,N_4078,N_4215);
nor U4494 (N_4494,N_4016,N_4236);
and U4495 (N_4495,N_4096,N_4113);
or U4496 (N_4496,N_4093,N_4027);
and U4497 (N_4497,N_4027,N_4074);
and U4498 (N_4498,N_4169,N_4236);
nor U4499 (N_4499,N_4087,N_4196);
nor U4500 (N_4500,N_4340,N_4384);
and U4501 (N_4501,N_4469,N_4462);
nand U4502 (N_4502,N_4457,N_4405);
nor U4503 (N_4503,N_4365,N_4320);
nor U4504 (N_4504,N_4290,N_4287);
and U4505 (N_4505,N_4482,N_4266);
nand U4506 (N_4506,N_4388,N_4443);
and U4507 (N_4507,N_4464,N_4252);
xor U4508 (N_4508,N_4428,N_4262);
and U4509 (N_4509,N_4352,N_4300);
or U4510 (N_4510,N_4339,N_4331);
or U4511 (N_4511,N_4424,N_4474);
nor U4512 (N_4512,N_4460,N_4281);
xnor U4513 (N_4513,N_4465,N_4477);
nor U4514 (N_4514,N_4323,N_4383);
or U4515 (N_4515,N_4393,N_4497);
or U4516 (N_4516,N_4408,N_4347);
nor U4517 (N_4517,N_4298,N_4329);
or U4518 (N_4518,N_4414,N_4299);
xnor U4519 (N_4519,N_4260,N_4434);
and U4520 (N_4520,N_4385,N_4472);
xor U4521 (N_4521,N_4371,N_4445);
nor U4522 (N_4522,N_4412,N_4325);
xnor U4523 (N_4523,N_4406,N_4256);
and U4524 (N_4524,N_4440,N_4452);
or U4525 (N_4525,N_4416,N_4369);
and U4526 (N_4526,N_4448,N_4302);
and U4527 (N_4527,N_4419,N_4476);
and U4528 (N_4528,N_4410,N_4399);
nor U4529 (N_4529,N_4390,N_4335);
nand U4530 (N_4530,N_4484,N_4435);
nand U4531 (N_4531,N_4431,N_4350);
or U4532 (N_4532,N_4489,N_4386);
nor U4533 (N_4533,N_4278,N_4346);
and U4534 (N_4534,N_4473,N_4432);
nand U4535 (N_4535,N_4306,N_4475);
nand U4536 (N_4536,N_4355,N_4328);
xor U4537 (N_4537,N_4312,N_4427);
xor U4538 (N_4538,N_4470,N_4313);
nand U4539 (N_4539,N_4254,N_4495);
and U4540 (N_4540,N_4283,N_4433);
nor U4541 (N_4541,N_4295,N_4370);
or U4542 (N_4542,N_4444,N_4311);
or U4543 (N_4543,N_4269,N_4250);
nor U4544 (N_4544,N_4351,N_4353);
or U4545 (N_4545,N_4317,N_4285);
or U4546 (N_4546,N_4326,N_4275);
nor U4547 (N_4547,N_4467,N_4334);
nand U4548 (N_4548,N_4341,N_4272);
xor U4549 (N_4549,N_4292,N_4490);
nand U4550 (N_4550,N_4322,N_4439);
nand U4551 (N_4551,N_4319,N_4332);
nand U4552 (N_4552,N_4310,N_4389);
and U4553 (N_4553,N_4491,N_4263);
and U4554 (N_4554,N_4418,N_4348);
xor U4555 (N_4555,N_4358,N_4437);
or U4556 (N_4556,N_4461,N_4401);
nor U4557 (N_4557,N_4451,N_4360);
xor U4558 (N_4558,N_4466,N_4493);
xnor U4559 (N_4559,N_4421,N_4430);
or U4560 (N_4560,N_4316,N_4446);
nand U4561 (N_4561,N_4337,N_4463);
or U4562 (N_4562,N_4487,N_4381);
or U4563 (N_4563,N_4314,N_4288);
nand U4564 (N_4564,N_4425,N_4382);
and U4565 (N_4565,N_4293,N_4296);
xnor U4566 (N_4566,N_4488,N_4376);
xnor U4567 (N_4567,N_4361,N_4447);
and U4568 (N_4568,N_4392,N_4307);
or U4569 (N_4569,N_4494,N_4282);
or U4570 (N_4570,N_4366,N_4327);
xor U4571 (N_4571,N_4407,N_4276);
nand U4572 (N_4572,N_4413,N_4258);
nand U4573 (N_4573,N_4284,N_4397);
xor U4574 (N_4574,N_4455,N_4318);
xnor U4575 (N_4575,N_4496,N_4442);
nor U4576 (N_4576,N_4264,N_4261);
or U4577 (N_4577,N_4342,N_4459);
nor U4578 (N_4578,N_4257,N_4404);
or U4579 (N_4579,N_4273,N_4279);
nor U4580 (N_4580,N_4400,N_4301);
xor U4581 (N_4581,N_4357,N_4330);
nand U4582 (N_4582,N_4486,N_4423);
and U4583 (N_4583,N_4315,N_4394);
nand U4584 (N_4584,N_4409,N_4387);
xor U4585 (N_4585,N_4344,N_4415);
nand U4586 (N_4586,N_4305,N_4255);
nor U4587 (N_4587,N_4368,N_4259);
xor U4588 (N_4588,N_4359,N_4426);
nor U4589 (N_4589,N_4471,N_4308);
nand U4590 (N_4590,N_4429,N_4267);
xnor U4591 (N_4591,N_4345,N_4372);
xnor U4592 (N_4592,N_4289,N_4492);
or U4593 (N_4593,N_4349,N_4333);
and U4594 (N_4594,N_4417,N_4377);
and U4595 (N_4595,N_4270,N_4441);
xnor U4596 (N_4596,N_4291,N_4324);
and U4597 (N_4597,N_4294,N_4378);
or U4598 (N_4598,N_4379,N_4303);
nand U4599 (N_4599,N_4396,N_4253);
xor U4600 (N_4600,N_4251,N_4374);
nor U4601 (N_4601,N_4356,N_4456);
nand U4602 (N_4602,N_4380,N_4280);
xor U4603 (N_4603,N_4277,N_4411);
or U4604 (N_4604,N_4321,N_4395);
or U4605 (N_4605,N_4265,N_4478);
or U4606 (N_4606,N_4364,N_4373);
xor U4607 (N_4607,N_4375,N_4271);
nand U4608 (N_4608,N_4422,N_4398);
nand U4609 (N_4609,N_4268,N_4468);
nor U4610 (N_4610,N_4338,N_4286);
xor U4611 (N_4611,N_4453,N_4354);
nor U4612 (N_4612,N_4402,N_4481);
nor U4613 (N_4613,N_4480,N_4297);
nand U4614 (N_4614,N_4391,N_4449);
nand U4615 (N_4615,N_4483,N_4498);
nor U4616 (N_4616,N_4343,N_4274);
xor U4617 (N_4617,N_4367,N_4436);
xnor U4618 (N_4618,N_4450,N_4458);
or U4619 (N_4619,N_4479,N_4336);
nor U4620 (N_4620,N_4363,N_4438);
nand U4621 (N_4621,N_4403,N_4362);
nand U4622 (N_4622,N_4309,N_4420);
or U4623 (N_4623,N_4499,N_4304);
nand U4624 (N_4624,N_4485,N_4454);
nand U4625 (N_4625,N_4335,N_4349);
xnor U4626 (N_4626,N_4337,N_4355);
and U4627 (N_4627,N_4454,N_4458);
or U4628 (N_4628,N_4276,N_4398);
nor U4629 (N_4629,N_4467,N_4357);
nand U4630 (N_4630,N_4466,N_4306);
nor U4631 (N_4631,N_4409,N_4430);
nor U4632 (N_4632,N_4492,N_4330);
xor U4633 (N_4633,N_4499,N_4343);
and U4634 (N_4634,N_4499,N_4296);
and U4635 (N_4635,N_4273,N_4256);
xnor U4636 (N_4636,N_4463,N_4417);
xor U4637 (N_4637,N_4315,N_4306);
nand U4638 (N_4638,N_4312,N_4393);
nand U4639 (N_4639,N_4294,N_4340);
or U4640 (N_4640,N_4428,N_4427);
and U4641 (N_4641,N_4446,N_4292);
nor U4642 (N_4642,N_4301,N_4478);
and U4643 (N_4643,N_4317,N_4395);
xnor U4644 (N_4644,N_4474,N_4350);
nand U4645 (N_4645,N_4478,N_4472);
or U4646 (N_4646,N_4380,N_4465);
nor U4647 (N_4647,N_4429,N_4436);
nor U4648 (N_4648,N_4382,N_4301);
nand U4649 (N_4649,N_4390,N_4475);
nor U4650 (N_4650,N_4453,N_4334);
and U4651 (N_4651,N_4361,N_4257);
xnor U4652 (N_4652,N_4387,N_4331);
and U4653 (N_4653,N_4332,N_4390);
nor U4654 (N_4654,N_4428,N_4398);
xnor U4655 (N_4655,N_4383,N_4336);
or U4656 (N_4656,N_4373,N_4393);
nor U4657 (N_4657,N_4456,N_4289);
and U4658 (N_4658,N_4318,N_4487);
nand U4659 (N_4659,N_4277,N_4268);
and U4660 (N_4660,N_4304,N_4440);
or U4661 (N_4661,N_4451,N_4452);
or U4662 (N_4662,N_4457,N_4296);
and U4663 (N_4663,N_4448,N_4458);
nor U4664 (N_4664,N_4413,N_4331);
nor U4665 (N_4665,N_4345,N_4388);
nor U4666 (N_4666,N_4313,N_4334);
nor U4667 (N_4667,N_4498,N_4487);
nand U4668 (N_4668,N_4410,N_4382);
or U4669 (N_4669,N_4445,N_4490);
or U4670 (N_4670,N_4478,N_4450);
or U4671 (N_4671,N_4334,N_4310);
and U4672 (N_4672,N_4393,N_4269);
xor U4673 (N_4673,N_4487,N_4371);
and U4674 (N_4674,N_4380,N_4288);
nor U4675 (N_4675,N_4428,N_4495);
and U4676 (N_4676,N_4296,N_4254);
nand U4677 (N_4677,N_4291,N_4434);
nor U4678 (N_4678,N_4285,N_4298);
and U4679 (N_4679,N_4467,N_4315);
or U4680 (N_4680,N_4417,N_4454);
xor U4681 (N_4681,N_4356,N_4322);
and U4682 (N_4682,N_4298,N_4477);
and U4683 (N_4683,N_4406,N_4332);
and U4684 (N_4684,N_4266,N_4259);
xor U4685 (N_4685,N_4430,N_4351);
xnor U4686 (N_4686,N_4484,N_4284);
nor U4687 (N_4687,N_4439,N_4416);
or U4688 (N_4688,N_4350,N_4337);
xor U4689 (N_4689,N_4344,N_4363);
xor U4690 (N_4690,N_4459,N_4430);
nor U4691 (N_4691,N_4328,N_4336);
and U4692 (N_4692,N_4280,N_4293);
xnor U4693 (N_4693,N_4286,N_4390);
nor U4694 (N_4694,N_4399,N_4452);
nor U4695 (N_4695,N_4305,N_4377);
nand U4696 (N_4696,N_4421,N_4273);
xor U4697 (N_4697,N_4272,N_4321);
nor U4698 (N_4698,N_4269,N_4437);
xor U4699 (N_4699,N_4472,N_4388);
or U4700 (N_4700,N_4480,N_4260);
nor U4701 (N_4701,N_4415,N_4466);
nor U4702 (N_4702,N_4390,N_4494);
xor U4703 (N_4703,N_4412,N_4351);
nor U4704 (N_4704,N_4449,N_4397);
xnor U4705 (N_4705,N_4341,N_4473);
xnor U4706 (N_4706,N_4381,N_4480);
xor U4707 (N_4707,N_4395,N_4418);
or U4708 (N_4708,N_4288,N_4452);
and U4709 (N_4709,N_4361,N_4251);
nor U4710 (N_4710,N_4485,N_4295);
or U4711 (N_4711,N_4493,N_4340);
nand U4712 (N_4712,N_4417,N_4328);
or U4713 (N_4713,N_4285,N_4485);
and U4714 (N_4714,N_4435,N_4377);
and U4715 (N_4715,N_4450,N_4360);
xor U4716 (N_4716,N_4289,N_4352);
or U4717 (N_4717,N_4449,N_4258);
and U4718 (N_4718,N_4339,N_4343);
nor U4719 (N_4719,N_4394,N_4475);
or U4720 (N_4720,N_4276,N_4349);
xor U4721 (N_4721,N_4370,N_4345);
or U4722 (N_4722,N_4350,N_4382);
and U4723 (N_4723,N_4250,N_4458);
or U4724 (N_4724,N_4426,N_4416);
or U4725 (N_4725,N_4497,N_4460);
and U4726 (N_4726,N_4428,N_4459);
xnor U4727 (N_4727,N_4296,N_4361);
or U4728 (N_4728,N_4262,N_4427);
and U4729 (N_4729,N_4262,N_4310);
and U4730 (N_4730,N_4440,N_4269);
and U4731 (N_4731,N_4280,N_4397);
nand U4732 (N_4732,N_4439,N_4449);
and U4733 (N_4733,N_4476,N_4448);
nand U4734 (N_4734,N_4488,N_4277);
and U4735 (N_4735,N_4396,N_4405);
or U4736 (N_4736,N_4276,N_4347);
and U4737 (N_4737,N_4316,N_4408);
nand U4738 (N_4738,N_4365,N_4448);
or U4739 (N_4739,N_4273,N_4315);
or U4740 (N_4740,N_4430,N_4498);
and U4741 (N_4741,N_4309,N_4349);
xnor U4742 (N_4742,N_4469,N_4268);
or U4743 (N_4743,N_4494,N_4445);
xor U4744 (N_4744,N_4311,N_4366);
xor U4745 (N_4745,N_4257,N_4283);
or U4746 (N_4746,N_4467,N_4270);
xor U4747 (N_4747,N_4299,N_4383);
nor U4748 (N_4748,N_4444,N_4286);
and U4749 (N_4749,N_4307,N_4441);
and U4750 (N_4750,N_4555,N_4643);
and U4751 (N_4751,N_4638,N_4749);
xnor U4752 (N_4752,N_4669,N_4628);
or U4753 (N_4753,N_4514,N_4704);
or U4754 (N_4754,N_4713,N_4561);
nand U4755 (N_4755,N_4513,N_4591);
nor U4756 (N_4756,N_4539,N_4613);
nand U4757 (N_4757,N_4564,N_4578);
nor U4758 (N_4758,N_4590,N_4720);
xor U4759 (N_4759,N_4505,N_4573);
or U4760 (N_4760,N_4667,N_4640);
nor U4761 (N_4761,N_4579,N_4503);
nor U4762 (N_4762,N_4666,N_4646);
nand U4763 (N_4763,N_4575,N_4728);
or U4764 (N_4764,N_4615,N_4595);
nor U4765 (N_4765,N_4625,N_4620);
nor U4766 (N_4766,N_4527,N_4512);
or U4767 (N_4767,N_4501,N_4629);
xor U4768 (N_4768,N_4518,N_4616);
nand U4769 (N_4769,N_4529,N_4682);
xnor U4770 (N_4770,N_4663,N_4535);
nor U4771 (N_4771,N_4627,N_4739);
nand U4772 (N_4772,N_4708,N_4692);
xnor U4773 (N_4773,N_4710,N_4695);
nor U4774 (N_4774,N_4607,N_4596);
xor U4775 (N_4775,N_4737,N_4538);
or U4776 (N_4776,N_4520,N_4626);
xnor U4777 (N_4777,N_4624,N_4617);
nand U4778 (N_4778,N_4515,N_4719);
nor U4779 (N_4779,N_4565,N_4655);
nor U4780 (N_4780,N_4690,N_4588);
nand U4781 (N_4781,N_4597,N_4724);
nand U4782 (N_4782,N_4605,N_4521);
and U4783 (N_4783,N_4697,N_4542);
nor U4784 (N_4784,N_4696,N_4693);
xnor U4785 (N_4785,N_4689,N_4623);
xnor U4786 (N_4786,N_4664,N_4691);
xnor U4787 (N_4787,N_4592,N_4545);
or U4788 (N_4788,N_4712,N_4621);
nand U4789 (N_4789,N_4594,N_4651);
nor U4790 (N_4790,N_4662,N_4653);
or U4791 (N_4791,N_4504,N_4654);
nor U4792 (N_4792,N_4601,N_4531);
nand U4793 (N_4793,N_4570,N_4526);
nor U4794 (N_4794,N_4675,N_4726);
and U4795 (N_4795,N_4510,N_4733);
nor U4796 (N_4796,N_4560,N_4644);
nand U4797 (N_4797,N_4676,N_4530);
nand U4798 (N_4798,N_4547,N_4516);
and U4799 (N_4799,N_4686,N_4583);
xor U4800 (N_4800,N_4577,N_4725);
xnor U4801 (N_4801,N_4706,N_4648);
and U4802 (N_4802,N_4658,N_4727);
or U4803 (N_4803,N_4522,N_4670);
nor U4804 (N_4804,N_4523,N_4748);
or U4805 (N_4805,N_4568,N_4685);
nand U4806 (N_4806,N_4649,N_4723);
xor U4807 (N_4807,N_4582,N_4618);
or U4808 (N_4808,N_4534,N_4536);
nor U4809 (N_4809,N_4735,N_4645);
nor U4810 (N_4810,N_4742,N_4598);
and U4811 (N_4811,N_4673,N_4745);
and U4812 (N_4812,N_4525,N_4507);
and U4813 (N_4813,N_4684,N_4567);
or U4814 (N_4814,N_4674,N_4734);
xnor U4815 (N_4815,N_4587,N_4537);
or U4816 (N_4816,N_4672,N_4548);
and U4817 (N_4817,N_4715,N_4540);
nand U4818 (N_4818,N_4702,N_4608);
nand U4819 (N_4819,N_4677,N_4604);
xnor U4820 (N_4820,N_4569,N_4688);
nand U4821 (N_4821,N_4705,N_4718);
and U4822 (N_4822,N_4559,N_4659);
and U4823 (N_4823,N_4665,N_4701);
xnor U4824 (N_4824,N_4610,N_4687);
or U4825 (N_4825,N_4586,N_4611);
nand U4826 (N_4826,N_4668,N_4500);
nor U4827 (N_4827,N_4679,N_4511);
nand U4828 (N_4828,N_4707,N_4632);
or U4829 (N_4829,N_4619,N_4699);
or U4830 (N_4830,N_4639,N_4543);
or U4831 (N_4831,N_4711,N_4546);
xnor U4832 (N_4832,N_4614,N_4642);
and U4833 (N_4833,N_4647,N_4622);
and U4834 (N_4834,N_4576,N_4631);
xor U4835 (N_4835,N_4671,N_4636);
nor U4836 (N_4836,N_4716,N_4572);
or U4837 (N_4837,N_4731,N_4656);
nand U4838 (N_4838,N_4747,N_4599);
xnor U4839 (N_4839,N_4732,N_4660);
and U4840 (N_4840,N_4729,N_4549);
and U4841 (N_4841,N_4517,N_4574);
or U4842 (N_4842,N_4585,N_4506);
nor U4843 (N_4843,N_4528,N_4633);
and U4844 (N_4844,N_4612,N_4556);
or U4845 (N_4845,N_4600,N_4571);
nor U4846 (N_4846,N_4550,N_4741);
or U4847 (N_4847,N_4709,N_4714);
and U4848 (N_4848,N_4589,N_4722);
nor U4849 (N_4849,N_4551,N_4593);
or U4850 (N_4850,N_4609,N_4524);
nand U4851 (N_4851,N_4721,N_4603);
and U4852 (N_4852,N_4637,N_4657);
and U4853 (N_4853,N_4681,N_4508);
xor U4854 (N_4854,N_4738,N_4740);
and U4855 (N_4855,N_4730,N_4703);
or U4856 (N_4856,N_4630,N_4678);
nand U4857 (N_4857,N_4554,N_4634);
nor U4858 (N_4858,N_4680,N_4683);
xnor U4859 (N_4859,N_4584,N_4566);
xor U4860 (N_4860,N_4558,N_4519);
and U4861 (N_4861,N_4541,N_4553);
nand U4862 (N_4862,N_4641,N_4650);
nor U4863 (N_4863,N_4602,N_4652);
or U4864 (N_4864,N_4581,N_4700);
nor U4865 (N_4865,N_4744,N_4635);
nor U4866 (N_4866,N_4509,N_4694);
or U4867 (N_4867,N_4502,N_4743);
nand U4868 (N_4868,N_4580,N_4532);
xor U4869 (N_4869,N_4544,N_4563);
xnor U4870 (N_4870,N_4606,N_4661);
xor U4871 (N_4871,N_4562,N_4736);
and U4872 (N_4872,N_4552,N_4698);
and U4873 (N_4873,N_4557,N_4717);
xor U4874 (N_4874,N_4746,N_4533);
nand U4875 (N_4875,N_4568,N_4564);
xnor U4876 (N_4876,N_4706,N_4590);
nand U4877 (N_4877,N_4536,N_4721);
nor U4878 (N_4878,N_4589,N_4683);
nor U4879 (N_4879,N_4710,N_4642);
and U4880 (N_4880,N_4554,N_4560);
nand U4881 (N_4881,N_4737,N_4531);
or U4882 (N_4882,N_4520,N_4734);
and U4883 (N_4883,N_4681,N_4546);
nor U4884 (N_4884,N_4652,N_4715);
nor U4885 (N_4885,N_4699,N_4648);
and U4886 (N_4886,N_4611,N_4637);
nand U4887 (N_4887,N_4532,N_4500);
and U4888 (N_4888,N_4516,N_4689);
nor U4889 (N_4889,N_4633,N_4584);
or U4890 (N_4890,N_4627,N_4540);
nand U4891 (N_4891,N_4715,N_4628);
xnor U4892 (N_4892,N_4552,N_4519);
and U4893 (N_4893,N_4666,N_4563);
xor U4894 (N_4894,N_4746,N_4653);
or U4895 (N_4895,N_4550,N_4599);
nand U4896 (N_4896,N_4642,N_4519);
or U4897 (N_4897,N_4692,N_4640);
nand U4898 (N_4898,N_4520,N_4547);
xnor U4899 (N_4899,N_4742,N_4632);
and U4900 (N_4900,N_4513,N_4529);
xnor U4901 (N_4901,N_4660,N_4548);
and U4902 (N_4902,N_4683,N_4642);
nor U4903 (N_4903,N_4567,N_4534);
nand U4904 (N_4904,N_4696,N_4681);
or U4905 (N_4905,N_4745,N_4707);
nand U4906 (N_4906,N_4505,N_4553);
nor U4907 (N_4907,N_4742,N_4518);
nor U4908 (N_4908,N_4594,N_4655);
nor U4909 (N_4909,N_4518,N_4697);
nand U4910 (N_4910,N_4595,N_4658);
nor U4911 (N_4911,N_4575,N_4569);
xor U4912 (N_4912,N_4625,N_4522);
or U4913 (N_4913,N_4687,N_4515);
nand U4914 (N_4914,N_4591,N_4555);
nor U4915 (N_4915,N_4620,N_4529);
nand U4916 (N_4916,N_4572,N_4571);
or U4917 (N_4917,N_4564,N_4699);
and U4918 (N_4918,N_4703,N_4558);
and U4919 (N_4919,N_4621,N_4530);
nand U4920 (N_4920,N_4628,N_4568);
and U4921 (N_4921,N_4681,N_4683);
xnor U4922 (N_4922,N_4663,N_4502);
or U4923 (N_4923,N_4624,N_4665);
and U4924 (N_4924,N_4583,N_4658);
or U4925 (N_4925,N_4720,N_4744);
or U4926 (N_4926,N_4678,N_4679);
xnor U4927 (N_4927,N_4644,N_4638);
or U4928 (N_4928,N_4571,N_4664);
xor U4929 (N_4929,N_4551,N_4700);
xor U4930 (N_4930,N_4683,N_4611);
and U4931 (N_4931,N_4744,N_4709);
or U4932 (N_4932,N_4526,N_4692);
nor U4933 (N_4933,N_4712,N_4640);
xnor U4934 (N_4934,N_4558,N_4635);
nor U4935 (N_4935,N_4749,N_4731);
nand U4936 (N_4936,N_4602,N_4517);
nor U4937 (N_4937,N_4521,N_4693);
or U4938 (N_4938,N_4622,N_4677);
nand U4939 (N_4939,N_4592,N_4622);
or U4940 (N_4940,N_4557,N_4648);
nand U4941 (N_4941,N_4706,N_4526);
nor U4942 (N_4942,N_4556,N_4712);
nand U4943 (N_4943,N_4623,N_4505);
or U4944 (N_4944,N_4715,N_4668);
and U4945 (N_4945,N_4547,N_4562);
or U4946 (N_4946,N_4688,N_4673);
and U4947 (N_4947,N_4548,N_4626);
and U4948 (N_4948,N_4645,N_4546);
or U4949 (N_4949,N_4607,N_4739);
nor U4950 (N_4950,N_4560,N_4636);
nor U4951 (N_4951,N_4519,N_4733);
and U4952 (N_4952,N_4525,N_4518);
nor U4953 (N_4953,N_4507,N_4601);
xnor U4954 (N_4954,N_4654,N_4572);
or U4955 (N_4955,N_4688,N_4531);
and U4956 (N_4956,N_4644,N_4666);
and U4957 (N_4957,N_4722,N_4649);
or U4958 (N_4958,N_4745,N_4663);
nor U4959 (N_4959,N_4530,N_4618);
or U4960 (N_4960,N_4709,N_4728);
or U4961 (N_4961,N_4503,N_4560);
nand U4962 (N_4962,N_4623,N_4509);
or U4963 (N_4963,N_4721,N_4599);
nand U4964 (N_4964,N_4566,N_4643);
or U4965 (N_4965,N_4628,N_4552);
nand U4966 (N_4966,N_4573,N_4586);
xor U4967 (N_4967,N_4650,N_4710);
nor U4968 (N_4968,N_4588,N_4506);
nand U4969 (N_4969,N_4616,N_4575);
nand U4970 (N_4970,N_4575,N_4658);
xnor U4971 (N_4971,N_4642,N_4744);
xor U4972 (N_4972,N_4584,N_4712);
nor U4973 (N_4973,N_4696,N_4745);
and U4974 (N_4974,N_4563,N_4694);
xnor U4975 (N_4975,N_4559,N_4626);
nand U4976 (N_4976,N_4703,N_4505);
nand U4977 (N_4977,N_4636,N_4577);
nand U4978 (N_4978,N_4503,N_4646);
nor U4979 (N_4979,N_4538,N_4501);
xnor U4980 (N_4980,N_4619,N_4638);
nor U4981 (N_4981,N_4585,N_4714);
nor U4982 (N_4982,N_4594,N_4550);
or U4983 (N_4983,N_4692,N_4703);
nor U4984 (N_4984,N_4684,N_4558);
nand U4985 (N_4985,N_4716,N_4652);
nand U4986 (N_4986,N_4504,N_4677);
nand U4987 (N_4987,N_4551,N_4674);
xor U4988 (N_4988,N_4529,N_4665);
or U4989 (N_4989,N_4653,N_4594);
or U4990 (N_4990,N_4736,N_4518);
or U4991 (N_4991,N_4637,N_4544);
or U4992 (N_4992,N_4590,N_4513);
nor U4993 (N_4993,N_4617,N_4734);
nor U4994 (N_4994,N_4749,N_4595);
xnor U4995 (N_4995,N_4574,N_4508);
nor U4996 (N_4996,N_4648,N_4613);
nand U4997 (N_4997,N_4644,N_4546);
nand U4998 (N_4998,N_4557,N_4615);
and U4999 (N_4999,N_4647,N_4683);
nand U5000 (N_5000,N_4834,N_4772);
nor U5001 (N_5001,N_4956,N_4985);
nand U5002 (N_5002,N_4983,N_4911);
nand U5003 (N_5003,N_4895,N_4998);
nand U5004 (N_5004,N_4984,N_4768);
xor U5005 (N_5005,N_4946,N_4972);
nand U5006 (N_5006,N_4824,N_4879);
nor U5007 (N_5007,N_4961,N_4893);
nor U5008 (N_5008,N_4812,N_4819);
nand U5009 (N_5009,N_4842,N_4873);
nand U5010 (N_5010,N_4838,N_4865);
nor U5011 (N_5011,N_4871,N_4943);
or U5012 (N_5012,N_4992,N_4951);
or U5013 (N_5013,N_4790,N_4885);
nand U5014 (N_5014,N_4816,N_4804);
xnor U5015 (N_5015,N_4821,N_4909);
xnor U5016 (N_5016,N_4907,N_4887);
or U5017 (N_5017,N_4839,N_4960);
or U5018 (N_5018,N_4898,N_4773);
nor U5019 (N_5019,N_4903,N_4784);
or U5020 (N_5020,N_4797,N_4916);
or U5021 (N_5021,N_4979,N_4932);
nand U5022 (N_5022,N_4837,N_4771);
or U5023 (N_5023,N_4931,N_4817);
xor U5024 (N_5024,N_4905,N_4766);
nand U5025 (N_5025,N_4802,N_4823);
xor U5026 (N_5026,N_4763,N_4954);
nor U5027 (N_5027,N_4798,N_4910);
nand U5028 (N_5028,N_4927,N_4929);
and U5029 (N_5029,N_4936,N_4840);
and U5030 (N_5030,N_4755,N_4825);
and U5031 (N_5031,N_4974,N_4852);
or U5032 (N_5032,N_4814,N_4869);
and U5033 (N_5033,N_4944,N_4897);
or U5034 (N_5034,N_4891,N_4882);
or U5035 (N_5035,N_4775,N_4789);
or U5036 (N_5036,N_4901,N_4783);
xnor U5037 (N_5037,N_4937,N_4836);
and U5038 (N_5038,N_4762,N_4966);
nand U5039 (N_5039,N_4877,N_4958);
or U5040 (N_5040,N_4963,N_4853);
xor U5041 (N_5041,N_4926,N_4851);
nand U5042 (N_5042,N_4919,N_4870);
nor U5043 (N_5043,N_4808,N_4805);
or U5044 (N_5044,N_4862,N_4922);
or U5045 (N_5045,N_4997,N_4953);
xor U5046 (N_5046,N_4938,N_4968);
and U5047 (N_5047,N_4883,N_4861);
xor U5048 (N_5048,N_4999,N_4978);
nand U5049 (N_5049,N_4913,N_4781);
or U5050 (N_5050,N_4795,N_4982);
and U5051 (N_5051,N_4874,N_4925);
xnor U5052 (N_5052,N_4856,N_4930);
xnor U5053 (N_5053,N_4902,N_4769);
or U5054 (N_5054,N_4900,N_4947);
or U5055 (N_5055,N_4977,N_4878);
nand U5056 (N_5056,N_4987,N_4796);
or U5057 (N_5057,N_4765,N_4807);
nand U5058 (N_5058,N_4787,N_4886);
nand U5059 (N_5059,N_4906,N_4940);
nor U5060 (N_5060,N_4815,N_4845);
nand U5061 (N_5061,N_4971,N_4924);
or U5062 (N_5062,N_4764,N_4778);
nand U5063 (N_5063,N_4993,N_4801);
or U5064 (N_5064,N_4829,N_4875);
xor U5065 (N_5065,N_4849,N_4908);
xor U5066 (N_5066,N_4912,N_4793);
or U5067 (N_5067,N_4975,N_4872);
nor U5068 (N_5068,N_4969,N_4761);
nand U5069 (N_5069,N_4918,N_4976);
or U5070 (N_5070,N_4970,N_4818);
nand U5071 (N_5071,N_4994,N_4811);
nand U5072 (N_5072,N_4884,N_4986);
nand U5073 (N_5073,N_4841,N_4806);
or U5074 (N_5074,N_4915,N_4751);
nand U5075 (N_5075,N_4803,N_4813);
xnor U5076 (N_5076,N_4880,N_4995);
nand U5077 (N_5077,N_4760,N_4866);
or U5078 (N_5078,N_4933,N_4859);
nand U5079 (N_5079,N_4962,N_4830);
xor U5080 (N_5080,N_4832,N_4914);
nand U5081 (N_5081,N_4864,N_4881);
xnor U5082 (N_5082,N_4923,N_4809);
or U5083 (N_5083,N_4920,N_4867);
and U5084 (N_5084,N_4799,N_4935);
xnor U5085 (N_5085,N_4770,N_4820);
and U5086 (N_5086,N_4843,N_4868);
xor U5087 (N_5087,N_4948,N_4756);
and U5088 (N_5088,N_4827,N_4896);
nand U5089 (N_5089,N_4828,N_4752);
nor U5090 (N_5090,N_4889,N_4890);
nor U5091 (N_5091,N_4894,N_4757);
and U5092 (N_5092,N_4964,N_4965);
and U5093 (N_5093,N_4928,N_4800);
xnor U5094 (N_5094,N_4782,N_4750);
nor U5095 (N_5095,N_4950,N_4774);
nor U5096 (N_5096,N_4846,N_4791);
nand U5097 (N_5097,N_4899,N_4955);
nand U5098 (N_5098,N_4876,N_4860);
or U5099 (N_5099,N_4952,N_4904);
nand U5100 (N_5100,N_4981,N_4959);
nor U5101 (N_5101,N_4957,N_4996);
xnor U5102 (N_5102,N_4759,N_4939);
nand U5103 (N_5103,N_4921,N_4942);
nand U5104 (N_5104,N_4831,N_4826);
xnor U5105 (N_5105,N_4854,N_4835);
nor U5106 (N_5106,N_4858,N_4888);
xor U5107 (N_5107,N_4917,N_4792);
or U5108 (N_5108,N_4758,N_4967);
nor U5109 (N_5109,N_4855,N_4780);
or U5110 (N_5110,N_4989,N_4980);
nand U5111 (N_5111,N_4753,N_4945);
or U5112 (N_5112,N_4777,N_4844);
nand U5113 (N_5113,N_4857,N_4892);
and U5114 (N_5114,N_4810,N_4847);
and U5115 (N_5115,N_4848,N_4788);
and U5116 (N_5116,N_4850,N_4833);
nor U5117 (N_5117,N_4776,N_4786);
nand U5118 (N_5118,N_4973,N_4991);
or U5119 (N_5119,N_4949,N_4988);
or U5120 (N_5120,N_4754,N_4779);
xnor U5121 (N_5121,N_4863,N_4785);
and U5122 (N_5122,N_4822,N_4767);
xor U5123 (N_5123,N_4934,N_4794);
or U5124 (N_5124,N_4941,N_4990);
xnor U5125 (N_5125,N_4906,N_4926);
nor U5126 (N_5126,N_4949,N_4848);
xnor U5127 (N_5127,N_4960,N_4986);
or U5128 (N_5128,N_4938,N_4896);
or U5129 (N_5129,N_4989,N_4975);
xor U5130 (N_5130,N_4985,N_4930);
nor U5131 (N_5131,N_4859,N_4772);
nor U5132 (N_5132,N_4962,N_4976);
xor U5133 (N_5133,N_4894,N_4850);
nor U5134 (N_5134,N_4876,N_4992);
nor U5135 (N_5135,N_4795,N_4902);
nor U5136 (N_5136,N_4954,N_4989);
nor U5137 (N_5137,N_4929,N_4875);
nand U5138 (N_5138,N_4921,N_4775);
or U5139 (N_5139,N_4804,N_4817);
nand U5140 (N_5140,N_4761,N_4970);
or U5141 (N_5141,N_4782,N_4851);
nand U5142 (N_5142,N_4824,N_4793);
xnor U5143 (N_5143,N_4813,N_4870);
or U5144 (N_5144,N_4850,N_4769);
nand U5145 (N_5145,N_4863,N_4867);
nor U5146 (N_5146,N_4887,N_4987);
or U5147 (N_5147,N_4922,N_4921);
and U5148 (N_5148,N_4976,N_4865);
and U5149 (N_5149,N_4794,N_4804);
nor U5150 (N_5150,N_4775,N_4871);
and U5151 (N_5151,N_4976,N_4834);
nand U5152 (N_5152,N_4854,N_4821);
nand U5153 (N_5153,N_4827,N_4751);
or U5154 (N_5154,N_4753,N_4999);
nand U5155 (N_5155,N_4954,N_4810);
nor U5156 (N_5156,N_4772,N_4876);
nor U5157 (N_5157,N_4909,N_4975);
or U5158 (N_5158,N_4971,N_4875);
or U5159 (N_5159,N_4942,N_4944);
xnor U5160 (N_5160,N_4837,N_4861);
and U5161 (N_5161,N_4751,N_4875);
and U5162 (N_5162,N_4830,N_4833);
nand U5163 (N_5163,N_4917,N_4751);
or U5164 (N_5164,N_4955,N_4962);
and U5165 (N_5165,N_4877,N_4998);
or U5166 (N_5166,N_4845,N_4941);
nor U5167 (N_5167,N_4934,N_4873);
and U5168 (N_5168,N_4950,N_4837);
nand U5169 (N_5169,N_4932,N_4758);
xor U5170 (N_5170,N_4973,N_4853);
and U5171 (N_5171,N_4973,N_4924);
or U5172 (N_5172,N_4827,N_4887);
xor U5173 (N_5173,N_4929,N_4863);
nor U5174 (N_5174,N_4965,N_4788);
or U5175 (N_5175,N_4798,N_4943);
nor U5176 (N_5176,N_4806,N_4857);
xnor U5177 (N_5177,N_4823,N_4908);
xnor U5178 (N_5178,N_4776,N_4780);
and U5179 (N_5179,N_4953,N_4760);
or U5180 (N_5180,N_4799,N_4772);
and U5181 (N_5181,N_4958,N_4768);
and U5182 (N_5182,N_4775,N_4868);
and U5183 (N_5183,N_4993,N_4983);
nand U5184 (N_5184,N_4794,N_4805);
or U5185 (N_5185,N_4791,N_4837);
xor U5186 (N_5186,N_4939,N_4959);
nand U5187 (N_5187,N_4794,N_4771);
and U5188 (N_5188,N_4975,N_4863);
xnor U5189 (N_5189,N_4778,N_4763);
nor U5190 (N_5190,N_4821,N_4750);
nor U5191 (N_5191,N_4885,N_4778);
or U5192 (N_5192,N_4816,N_4873);
nand U5193 (N_5193,N_4969,N_4792);
xnor U5194 (N_5194,N_4799,N_4817);
xor U5195 (N_5195,N_4960,N_4806);
nor U5196 (N_5196,N_4865,N_4843);
nor U5197 (N_5197,N_4889,N_4871);
nand U5198 (N_5198,N_4875,N_4861);
or U5199 (N_5199,N_4826,N_4896);
nand U5200 (N_5200,N_4906,N_4786);
nand U5201 (N_5201,N_4909,N_4965);
or U5202 (N_5202,N_4750,N_4783);
xnor U5203 (N_5203,N_4817,N_4801);
xnor U5204 (N_5204,N_4996,N_4934);
and U5205 (N_5205,N_4958,N_4863);
and U5206 (N_5206,N_4965,N_4890);
and U5207 (N_5207,N_4854,N_4849);
xnor U5208 (N_5208,N_4947,N_4809);
and U5209 (N_5209,N_4805,N_4918);
or U5210 (N_5210,N_4962,N_4773);
nor U5211 (N_5211,N_4960,N_4804);
xor U5212 (N_5212,N_4757,N_4948);
nor U5213 (N_5213,N_4884,N_4787);
or U5214 (N_5214,N_4947,N_4757);
xor U5215 (N_5215,N_4862,N_4975);
and U5216 (N_5216,N_4847,N_4831);
and U5217 (N_5217,N_4871,N_4970);
and U5218 (N_5218,N_4912,N_4860);
and U5219 (N_5219,N_4858,N_4764);
xor U5220 (N_5220,N_4835,N_4858);
nor U5221 (N_5221,N_4831,N_4988);
nand U5222 (N_5222,N_4854,N_4850);
xnor U5223 (N_5223,N_4835,N_4833);
nor U5224 (N_5224,N_4779,N_4837);
xor U5225 (N_5225,N_4784,N_4773);
or U5226 (N_5226,N_4754,N_4911);
or U5227 (N_5227,N_4978,N_4758);
and U5228 (N_5228,N_4921,N_4797);
xnor U5229 (N_5229,N_4862,N_4960);
and U5230 (N_5230,N_4846,N_4986);
nor U5231 (N_5231,N_4947,N_4760);
nor U5232 (N_5232,N_4959,N_4845);
nor U5233 (N_5233,N_4982,N_4781);
xor U5234 (N_5234,N_4856,N_4754);
nand U5235 (N_5235,N_4809,N_4981);
and U5236 (N_5236,N_4812,N_4966);
xnor U5237 (N_5237,N_4756,N_4899);
nand U5238 (N_5238,N_4904,N_4767);
xnor U5239 (N_5239,N_4752,N_4818);
xor U5240 (N_5240,N_4914,N_4902);
xnor U5241 (N_5241,N_4920,N_4763);
or U5242 (N_5242,N_4846,N_4803);
or U5243 (N_5243,N_4910,N_4823);
nand U5244 (N_5244,N_4924,N_4984);
nand U5245 (N_5245,N_4903,N_4759);
and U5246 (N_5246,N_4937,N_4852);
xor U5247 (N_5247,N_4817,N_4875);
nor U5248 (N_5248,N_4974,N_4883);
xor U5249 (N_5249,N_4909,N_4820);
nand U5250 (N_5250,N_5074,N_5056);
xnor U5251 (N_5251,N_5198,N_5188);
and U5252 (N_5252,N_5190,N_5119);
xor U5253 (N_5253,N_5153,N_5233);
nor U5254 (N_5254,N_5027,N_5066);
or U5255 (N_5255,N_5081,N_5051);
nor U5256 (N_5256,N_5015,N_5013);
or U5257 (N_5257,N_5036,N_5006);
xor U5258 (N_5258,N_5236,N_5131);
xnor U5259 (N_5259,N_5050,N_5052);
nand U5260 (N_5260,N_5109,N_5213);
and U5261 (N_5261,N_5086,N_5162);
and U5262 (N_5262,N_5063,N_5230);
and U5263 (N_5263,N_5249,N_5201);
nor U5264 (N_5264,N_5009,N_5176);
or U5265 (N_5265,N_5165,N_5134);
xnor U5266 (N_5266,N_5208,N_5221);
xor U5267 (N_5267,N_5019,N_5102);
or U5268 (N_5268,N_5042,N_5085);
and U5269 (N_5269,N_5016,N_5135);
or U5270 (N_5270,N_5089,N_5090);
and U5271 (N_5271,N_5128,N_5067);
nand U5272 (N_5272,N_5229,N_5200);
and U5273 (N_5273,N_5043,N_5002);
nor U5274 (N_5274,N_5114,N_5186);
nor U5275 (N_5275,N_5100,N_5166);
or U5276 (N_5276,N_5083,N_5206);
nand U5277 (N_5277,N_5143,N_5111);
nand U5278 (N_5278,N_5168,N_5017);
and U5279 (N_5279,N_5011,N_5193);
and U5280 (N_5280,N_5029,N_5088);
nor U5281 (N_5281,N_5149,N_5199);
or U5282 (N_5282,N_5101,N_5142);
or U5283 (N_5283,N_5174,N_5078);
xnor U5284 (N_5284,N_5008,N_5095);
nand U5285 (N_5285,N_5044,N_5021);
xnor U5286 (N_5286,N_5156,N_5048);
xnor U5287 (N_5287,N_5154,N_5205);
xnor U5288 (N_5288,N_5061,N_5133);
nor U5289 (N_5289,N_5039,N_5218);
or U5290 (N_5290,N_5239,N_5150);
and U5291 (N_5291,N_5004,N_5080);
and U5292 (N_5292,N_5010,N_5209);
or U5293 (N_5293,N_5072,N_5112);
xor U5294 (N_5294,N_5045,N_5227);
or U5295 (N_5295,N_5238,N_5082);
nor U5296 (N_5296,N_5038,N_5245);
xnor U5297 (N_5297,N_5189,N_5196);
or U5298 (N_5298,N_5173,N_5187);
or U5299 (N_5299,N_5022,N_5023);
nor U5300 (N_5300,N_5172,N_5057);
nand U5301 (N_5301,N_5181,N_5248);
nand U5302 (N_5302,N_5025,N_5182);
nand U5303 (N_5303,N_5237,N_5223);
xor U5304 (N_5304,N_5159,N_5026);
nand U5305 (N_5305,N_5120,N_5103);
and U5306 (N_5306,N_5152,N_5091);
and U5307 (N_5307,N_5179,N_5065);
nand U5308 (N_5308,N_5184,N_5139);
or U5309 (N_5309,N_5234,N_5069);
nand U5310 (N_5310,N_5145,N_5059);
and U5311 (N_5311,N_5098,N_5195);
nand U5312 (N_5312,N_5126,N_5020);
and U5313 (N_5313,N_5137,N_5216);
xor U5314 (N_5314,N_5064,N_5243);
and U5315 (N_5315,N_5110,N_5028);
nor U5316 (N_5316,N_5175,N_5092);
nand U5317 (N_5317,N_5107,N_5164);
or U5318 (N_5318,N_5210,N_5183);
nand U5319 (N_5319,N_5024,N_5058);
nand U5320 (N_5320,N_5192,N_5157);
xor U5321 (N_5321,N_5041,N_5005);
nand U5322 (N_5322,N_5144,N_5105);
and U5323 (N_5323,N_5070,N_5084);
xor U5324 (N_5324,N_5123,N_5141);
nor U5325 (N_5325,N_5241,N_5108);
xor U5326 (N_5326,N_5093,N_5033);
nand U5327 (N_5327,N_5117,N_5207);
and U5328 (N_5328,N_5202,N_5071);
xnor U5329 (N_5329,N_5034,N_5099);
nor U5330 (N_5330,N_5185,N_5125);
nand U5331 (N_5331,N_5160,N_5136);
nor U5332 (N_5332,N_5054,N_5014);
nand U5333 (N_5333,N_5155,N_5161);
and U5334 (N_5334,N_5177,N_5106);
xnor U5335 (N_5335,N_5204,N_5232);
nand U5336 (N_5336,N_5235,N_5076);
or U5337 (N_5337,N_5169,N_5104);
nor U5338 (N_5338,N_5032,N_5151);
xor U5339 (N_5339,N_5118,N_5130);
nor U5340 (N_5340,N_5222,N_5115);
nor U5341 (N_5341,N_5079,N_5148);
nor U5342 (N_5342,N_5124,N_5127);
and U5343 (N_5343,N_5018,N_5197);
xor U5344 (N_5344,N_5240,N_5217);
nand U5345 (N_5345,N_5191,N_5113);
or U5346 (N_5346,N_5226,N_5247);
xor U5347 (N_5347,N_5073,N_5140);
or U5348 (N_5348,N_5228,N_5116);
nor U5349 (N_5349,N_5035,N_5138);
and U5350 (N_5350,N_5129,N_5075);
nor U5351 (N_5351,N_5214,N_5047);
xor U5352 (N_5352,N_5003,N_5147);
nand U5353 (N_5353,N_5132,N_5040);
nand U5354 (N_5354,N_5171,N_5231);
or U5355 (N_5355,N_5077,N_5007);
or U5356 (N_5356,N_5030,N_5087);
or U5357 (N_5357,N_5001,N_5121);
nor U5358 (N_5358,N_5244,N_5037);
nand U5359 (N_5359,N_5060,N_5220);
nand U5360 (N_5360,N_5246,N_5096);
nand U5361 (N_5361,N_5224,N_5158);
xor U5362 (N_5362,N_5046,N_5122);
nor U5363 (N_5363,N_5170,N_5194);
and U5364 (N_5364,N_5055,N_5225);
xor U5365 (N_5365,N_5000,N_5012);
nand U5366 (N_5366,N_5167,N_5212);
and U5367 (N_5367,N_5242,N_5211);
nand U5368 (N_5368,N_5031,N_5178);
and U5369 (N_5369,N_5097,N_5094);
and U5370 (N_5370,N_5146,N_5053);
nor U5371 (N_5371,N_5068,N_5163);
or U5372 (N_5372,N_5219,N_5203);
xor U5373 (N_5373,N_5049,N_5215);
and U5374 (N_5374,N_5062,N_5180);
xnor U5375 (N_5375,N_5015,N_5205);
nand U5376 (N_5376,N_5206,N_5123);
xnor U5377 (N_5377,N_5187,N_5051);
or U5378 (N_5378,N_5091,N_5141);
or U5379 (N_5379,N_5231,N_5192);
nor U5380 (N_5380,N_5204,N_5191);
nand U5381 (N_5381,N_5148,N_5195);
and U5382 (N_5382,N_5099,N_5230);
nor U5383 (N_5383,N_5144,N_5181);
nor U5384 (N_5384,N_5206,N_5082);
nand U5385 (N_5385,N_5129,N_5222);
xor U5386 (N_5386,N_5219,N_5105);
nor U5387 (N_5387,N_5128,N_5027);
or U5388 (N_5388,N_5160,N_5131);
and U5389 (N_5389,N_5005,N_5138);
xor U5390 (N_5390,N_5107,N_5237);
xnor U5391 (N_5391,N_5164,N_5037);
nand U5392 (N_5392,N_5227,N_5088);
nand U5393 (N_5393,N_5193,N_5203);
nand U5394 (N_5394,N_5016,N_5236);
xor U5395 (N_5395,N_5235,N_5050);
or U5396 (N_5396,N_5182,N_5115);
nor U5397 (N_5397,N_5162,N_5055);
and U5398 (N_5398,N_5101,N_5111);
or U5399 (N_5399,N_5211,N_5165);
xor U5400 (N_5400,N_5135,N_5245);
or U5401 (N_5401,N_5002,N_5178);
or U5402 (N_5402,N_5207,N_5150);
or U5403 (N_5403,N_5057,N_5163);
nand U5404 (N_5404,N_5227,N_5108);
and U5405 (N_5405,N_5110,N_5088);
nand U5406 (N_5406,N_5123,N_5154);
and U5407 (N_5407,N_5066,N_5062);
nor U5408 (N_5408,N_5217,N_5144);
nor U5409 (N_5409,N_5066,N_5191);
and U5410 (N_5410,N_5105,N_5233);
and U5411 (N_5411,N_5073,N_5079);
nor U5412 (N_5412,N_5071,N_5159);
nor U5413 (N_5413,N_5201,N_5030);
or U5414 (N_5414,N_5143,N_5189);
nor U5415 (N_5415,N_5109,N_5172);
nand U5416 (N_5416,N_5027,N_5249);
xnor U5417 (N_5417,N_5222,N_5151);
xnor U5418 (N_5418,N_5144,N_5036);
or U5419 (N_5419,N_5086,N_5246);
nor U5420 (N_5420,N_5113,N_5207);
nor U5421 (N_5421,N_5116,N_5043);
or U5422 (N_5422,N_5205,N_5026);
nor U5423 (N_5423,N_5233,N_5094);
nor U5424 (N_5424,N_5001,N_5246);
and U5425 (N_5425,N_5052,N_5167);
xor U5426 (N_5426,N_5178,N_5124);
nand U5427 (N_5427,N_5120,N_5128);
and U5428 (N_5428,N_5165,N_5089);
and U5429 (N_5429,N_5068,N_5032);
nand U5430 (N_5430,N_5242,N_5110);
or U5431 (N_5431,N_5238,N_5205);
nand U5432 (N_5432,N_5014,N_5147);
or U5433 (N_5433,N_5173,N_5073);
and U5434 (N_5434,N_5107,N_5210);
and U5435 (N_5435,N_5098,N_5211);
or U5436 (N_5436,N_5095,N_5116);
nor U5437 (N_5437,N_5206,N_5215);
and U5438 (N_5438,N_5017,N_5053);
nand U5439 (N_5439,N_5211,N_5184);
and U5440 (N_5440,N_5009,N_5022);
nor U5441 (N_5441,N_5038,N_5053);
nor U5442 (N_5442,N_5010,N_5246);
nor U5443 (N_5443,N_5189,N_5186);
nand U5444 (N_5444,N_5065,N_5237);
and U5445 (N_5445,N_5029,N_5099);
nor U5446 (N_5446,N_5150,N_5035);
and U5447 (N_5447,N_5145,N_5054);
nor U5448 (N_5448,N_5227,N_5113);
nor U5449 (N_5449,N_5125,N_5108);
nand U5450 (N_5450,N_5039,N_5183);
nand U5451 (N_5451,N_5052,N_5168);
nand U5452 (N_5452,N_5137,N_5176);
nand U5453 (N_5453,N_5074,N_5239);
or U5454 (N_5454,N_5089,N_5040);
and U5455 (N_5455,N_5046,N_5169);
nor U5456 (N_5456,N_5093,N_5199);
nor U5457 (N_5457,N_5170,N_5235);
or U5458 (N_5458,N_5044,N_5079);
xnor U5459 (N_5459,N_5036,N_5021);
and U5460 (N_5460,N_5157,N_5068);
and U5461 (N_5461,N_5000,N_5191);
and U5462 (N_5462,N_5191,N_5098);
or U5463 (N_5463,N_5130,N_5192);
or U5464 (N_5464,N_5184,N_5210);
and U5465 (N_5465,N_5067,N_5144);
nor U5466 (N_5466,N_5073,N_5228);
xnor U5467 (N_5467,N_5132,N_5192);
or U5468 (N_5468,N_5154,N_5069);
nor U5469 (N_5469,N_5062,N_5178);
nand U5470 (N_5470,N_5080,N_5128);
and U5471 (N_5471,N_5210,N_5204);
or U5472 (N_5472,N_5154,N_5028);
nand U5473 (N_5473,N_5053,N_5208);
nand U5474 (N_5474,N_5025,N_5016);
or U5475 (N_5475,N_5124,N_5099);
and U5476 (N_5476,N_5018,N_5233);
and U5477 (N_5477,N_5117,N_5145);
xnor U5478 (N_5478,N_5117,N_5021);
and U5479 (N_5479,N_5212,N_5001);
or U5480 (N_5480,N_5239,N_5169);
xor U5481 (N_5481,N_5016,N_5193);
nand U5482 (N_5482,N_5061,N_5178);
or U5483 (N_5483,N_5190,N_5127);
and U5484 (N_5484,N_5202,N_5086);
xnor U5485 (N_5485,N_5005,N_5124);
nand U5486 (N_5486,N_5174,N_5013);
and U5487 (N_5487,N_5088,N_5215);
nand U5488 (N_5488,N_5010,N_5014);
and U5489 (N_5489,N_5189,N_5135);
nor U5490 (N_5490,N_5120,N_5101);
xnor U5491 (N_5491,N_5073,N_5048);
nor U5492 (N_5492,N_5202,N_5023);
xor U5493 (N_5493,N_5144,N_5053);
or U5494 (N_5494,N_5189,N_5214);
and U5495 (N_5495,N_5228,N_5130);
nand U5496 (N_5496,N_5231,N_5002);
nor U5497 (N_5497,N_5197,N_5238);
and U5498 (N_5498,N_5021,N_5004);
or U5499 (N_5499,N_5186,N_5009);
nand U5500 (N_5500,N_5409,N_5255);
and U5501 (N_5501,N_5489,N_5261);
nand U5502 (N_5502,N_5289,N_5358);
or U5503 (N_5503,N_5473,N_5268);
or U5504 (N_5504,N_5362,N_5460);
nor U5505 (N_5505,N_5407,N_5287);
and U5506 (N_5506,N_5361,N_5399);
or U5507 (N_5507,N_5343,N_5253);
nand U5508 (N_5508,N_5422,N_5281);
nor U5509 (N_5509,N_5423,N_5368);
xor U5510 (N_5510,N_5321,N_5424);
nand U5511 (N_5511,N_5372,N_5332);
nor U5512 (N_5512,N_5316,N_5292);
xnor U5513 (N_5513,N_5263,N_5415);
and U5514 (N_5514,N_5412,N_5339);
and U5515 (N_5515,N_5480,N_5326);
or U5516 (N_5516,N_5301,N_5357);
and U5517 (N_5517,N_5296,N_5383);
and U5518 (N_5518,N_5318,N_5468);
or U5519 (N_5519,N_5366,N_5319);
nand U5520 (N_5520,N_5302,N_5446);
xnor U5521 (N_5521,N_5359,N_5498);
xor U5522 (N_5522,N_5309,N_5496);
nand U5523 (N_5523,N_5450,N_5433);
nor U5524 (N_5524,N_5499,N_5440);
xor U5525 (N_5525,N_5351,N_5384);
nor U5526 (N_5526,N_5444,N_5322);
nand U5527 (N_5527,N_5260,N_5336);
or U5528 (N_5528,N_5454,N_5259);
or U5529 (N_5529,N_5284,N_5390);
or U5530 (N_5530,N_5386,N_5405);
nand U5531 (N_5531,N_5429,N_5467);
or U5532 (N_5532,N_5491,N_5314);
or U5533 (N_5533,N_5411,N_5436);
and U5534 (N_5534,N_5290,N_5455);
nor U5535 (N_5535,N_5312,N_5459);
or U5536 (N_5536,N_5493,N_5396);
nand U5537 (N_5537,N_5387,N_5254);
nand U5538 (N_5538,N_5347,N_5305);
nor U5539 (N_5539,N_5298,N_5435);
or U5540 (N_5540,N_5418,N_5427);
and U5541 (N_5541,N_5282,N_5331);
xnor U5542 (N_5542,N_5341,N_5295);
or U5543 (N_5543,N_5335,N_5342);
and U5544 (N_5544,N_5421,N_5494);
xnor U5545 (N_5545,N_5252,N_5442);
nor U5546 (N_5546,N_5272,N_5367);
xor U5547 (N_5547,N_5293,N_5337);
nor U5548 (N_5548,N_5420,N_5325);
nand U5549 (N_5549,N_5299,N_5307);
and U5550 (N_5550,N_5285,N_5274);
or U5551 (N_5551,N_5381,N_5398);
or U5552 (N_5552,N_5393,N_5266);
nand U5553 (N_5553,N_5371,N_5346);
and U5554 (N_5554,N_5324,N_5392);
nor U5555 (N_5555,N_5291,N_5317);
nand U5556 (N_5556,N_5417,N_5456);
nand U5557 (N_5557,N_5438,N_5490);
or U5558 (N_5558,N_5273,N_5401);
or U5559 (N_5559,N_5300,N_5469);
nand U5560 (N_5560,N_5470,N_5397);
xnor U5561 (N_5561,N_5414,N_5360);
nand U5562 (N_5562,N_5251,N_5445);
nor U5563 (N_5563,N_5431,N_5265);
nor U5564 (N_5564,N_5497,N_5425);
nor U5565 (N_5565,N_5495,N_5308);
and U5566 (N_5566,N_5408,N_5340);
nor U5567 (N_5567,N_5443,N_5416);
or U5568 (N_5568,N_5452,N_5382);
nand U5569 (N_5569,N_5391,N_5356);
nand U5570 (N_5570,N_5471,N_5428);
nand U5571 (N_5571,N_5303,N_5294);
nand U5572 (N_5572,N_5350,N_5388);
nor U5573 (N_5573,N_5441,N_5258);
or U5574 (N_5574,N_5373,N_5395);
nor U5575 (N_5575,N_5365,N_5306);
nand U5576 (N_5576,N_5377,N_5352);
xor U5577 (N_5577,N_5276,N_5482);
or U5578 (N_5578,N_5256,N_5410);
and U5579 (N_5579,N_5457,N_5353);
or U5580 (N_5580,N_5375,N_5463);
and U5581 (N_5581,N_5323,N_5279);
and U5582 (N_5582,N_5462,N_5330);
nand U5583 (N_5583,N_5328,N_5344);
nor U5584 (N_5584,N_5406,N_5264);
or U5585 (N_5585,N_5338,N_5278);
nand U5586 (N_5586,N_5447,N_5354);
xnor U5587 (N_5587,N_5486,N_5376);
or U5588 (N_5588,N_5449,N_5283);
or U5589 (N_5589,N_5439,N_5400);
and U5590 (N_5590,N_5315,N_5370);
xnor U5591 (N_5591,N_5404,N_5413);
xnor U5592 (N_5592,N_5363,N_5434);
nand U5593 (N_5593,N_5257,N_5333);
or U5594 (N_5594,N_5430,N_5481);
xnor U5595 (N_5595,N_5374,N_5355);
or U5596 (N_5596,N_5488,N_5432);
and U5597 (N_5597,N_5364,N_5458);
and U5598 (N_5598,N_5465,N_5310);
nor U5599 (N_5599,N_5286,N_5483);
and U5600 (N_5600,N_5329,N_5271);
nand U5601 (N_5601,N_5478,N_5437);
xnor U5602 (N_5602,N_5348,N_5313);
nand U5603 (N_5603,N_5385,N_5250);
or U5604 (N_5604,N_5476,N_5485);
xor U5605 (N_5605,N_5304,N_5269);
and U5606 (N_5606,N_5402,N_5320);
or U5607 (N_5607,N_5277,N_5267);
nand U5608 (N_5608,N_5378,N_5345);
nand U5609 (N_5609,N_5451,N_5270);
nand U5610 (N_5610,N_5474,N_5475);
xor U5611 (N_5611,N_5311,N_5394);
xnor U5612 (N_5612,N_5369,N_5487);
nor U5613 (N_5613,N_5466,N_5280);
nand U5614 (N_5614,N_5419,N_5403);
nand U5615 (N_5615,N_5453,N_5334);
or U5616 (N_5616,N_5484,N_5479);
and U5617 (N_5617,N_5448,N_5349);
and U5618 (N_5618,N_5461,N_5297);
xnor U5619 (N_5619,N_5492,N_5327);
nor U5620 (N_5620,N_5275,N_5262);
and U5621 (N_5621,N_5288,N_5426);
or U5622 (N_5622,N_5389,N_5464);
nand U5623 (N_5623,N_5379,N_5472);
or U5624 (N_5624,N_5380,N_5477);
nor U5625 (N_5625,N_5361,N_5367);
or U5626 (N_5626,N_5407,N_5254);
nand U5627 (N_5627,N_5333,N_5254);
nand U5628 (N_5628,N_5317,N_5381);
xor U5629 (N_5629,N_5329,N_5251);
nor U5630 (N_5630,N_5391,N_5351);
xnor U5631 (N_5631,N_5350,N_5468);
and U5632 (N_5632,N_5358,N_5306);
nand U5633 (N_5633,N_5470,N_5373);
and U5634 (N_5634,N_5441,N_5279);
nor U5635 (N_5635,N_5462,N_5309);
and U5636 (N_5636,N_5389,N_5436);
nor U5637 (N_5637,N_5428,N_5464);
nand U5638 (N_5638,N_5329,N_5444);
nor U5639 (N_5639,N_5436,N_5304);
nand U5640 (N_5640,N_5395,N_5499);
nand U5641 (N_5641,N_5338,N_5360);
and U5642 (N_5642,N_5354,N_5471);
nand U5643 (N_5643,N_5459,N_5380);
or U5644 (N_5644,N_5481,N_5489);
or U5645 (N_5645,N_5492,N_5287);
or U5646 (N_5646,N_5479,N_5431);
and U5647 (N_5647,N_5353,N_5463);
xnor U5648 (N_5648,N_5362,N_5459);
and U5649 (N_5649,N_5488,N_5483);
or U5650 (N_5650,N_5491,N_5329);
or U5651 (N_5651,N_5419,N_5444);
and U5652 (N_5652,N_5454,N_5494);
xor U5653 (N_5653,N_5393,N_5444);
or U5654 (N_5654,N_5274,N_5485);
nand U5655 (N_5655,N_5276,N_5368);
or U5656 (N_5656,N_5343,N_5418);
or U5657 (N_5657,N_5475,N_5330);
and U5658 (N_5658,N_5428,N_5278);
nand U5659 (N_5659,N_5388,N_5361);
nor U5660 (N_5660,N_5425,N_5281);
or U5661 (N_5661,N_5283,N_5410);
or U5662 (N_5662,N_5257,N_5385);
nand U5663 (N_5663,N_5287,N_5437);
xnor U5664 (N_5664,N_5304,N_5480);
or U5665 (N_5665,N_5327,N_5386);
xnor U5666 (N_5666,N_5300,N_5414);
or U5667 (N_5667,N_5396,N_5361);
xnor U5668 (N_5668,N_5458,N_5372);
nand U5669 (N_5669,N_5309,N_5264);
or U5670 (N_5670,N_5312,N_5423);
nor U5671 (N_5671,N_5291,N_5475);
or U5672 (N_5672,N_5464,N_5369);
nand U5673 (N_5673,N_5334,N_5282);
and U5674 (N_5674,N_5452,N_5380);
and U5675 (N_5675,N_5369,N_5317);
and U5676 (N_5676,N_5269,N_5316);
and U5677 (N_5677,N_5301,N_5253);
nor U5678 (N_5678,N_5340,N_5265);
xnor U5679 (N_5679,N_5329,N_5250);
or U5680 (N_5680,N_5310,N_5474);
and U5681 (N_5681,N_5362,N_5483);
nor U5682 (N_5682,N_5442,N_5335);
nor U5683 (N_5683,N_5282,N_5494);
nor U5684 (N_5684,N_5319,N_5459);
nor U5685 (N_5685,N_5332,N_5254);
nand U5686 (N_5686,N_5291,N_5463);
xnor U5687 (N_5687,N_5260,N_5251);
nand U5688 (N_5688,N_5348,N_5335);
nor U5689 (N_5689,N_5364,N_5443);
nand U5690 (N_5690,N_5330,N_5384);
and U5691 (N_5691,N_5425,N_5411);
nand U5692 (N_5692,N_5374,N_5272);
or U5693 (N_5693,N_5257,N_5452);
or U5694 (N_5694,N_5364,N_5383);
or U5695 (N_5695,N_5495,N_5397);
nand U5696 (N_5696,N_5288,N_5420);
xnor U5697 (N_5697,N_5309,N_5396);
nand U5698 (N_5698,N_5327,N_5402);
nand U5699 (N_5699,N_5359,N_5403);
nand U5700 (N_5700,N_5466,N_5298);
and U5701 (N_5701,N_5277,N_5308);
and U5702 (N_5702,N_5358,N_5489);
nor U5703 (N_5703,N_5466,N_5452);
nor U5704 (N_5704,N_5283,N_5287);
nor U5705 (N_5705,N_5460,N_5350);
xor U5706 (N_5706,N_5317,N_5303);
and U5707 (N_5707,N_5351,N_5286);
or U5708 (N_5708,N_5465,N_5455);
xor U5709 (N_5709,N_5497,N_5276);
nand U5710 (N_5710,N_5347,N_5310);
and U5711 (N_5711,N_5365,N_5267);
nor U5712 (N_5712,N_5424,N_5384);
nand U5713 (N_5713,N_5257,N_5494);
nand U5714 (N_5714,N_5415,N_5483);
nand U5715 (N_5715,N_5349,N_5322);
or U5716 (N_5716,N_5470,N_5454);
or U5717 (N_5717,N_5392,N_5412);
xnor U5718 (N_5718,N_5352,N_5341);
and U5719 (N_5719,N_5263,N_5416);
nor U5720 (N_5720,N_5286,N_5385);
nand U5721 (N_5721,N_5294,N_5299);
nand U5722 (N_5722,N_5259,N_5261);
and U5723 (N_5723,N_5257,N_5263);
nand U5724 (N_5724,N_5432,N_5397);
nand U5725 (N_5725,N_5483,N_5255);
xor U5726 (N_5726,N_5442,N_5355);
and U5727 (N_5727,N_5325,N_5411);
or U5728 (N_5728,N_5257,N_5329);
xor U5729 (N_5729,N_5384,N_5327);
nor U5730 (N_5730,N_5338,N_5420);
or U5731 (N_5731,N_5444,N_5404);
nand U5732 (N_5732,N_5386,N_5265);
nor U5733 (N_5733,N_5283,N_5419);
nand U5734 (N_5734,N_5253,N_5499);
xnor U5735 (N_5735,N_5463,N_5449);
or U5736 (N_5736,N_5458,N_5395);
and U5737 (N_5737,N_5370,N_5491);
nand U5738 (N_5738,N_5367,N_5365);
nor U5739 (N_5739,N_5277,N_5485);
xor U5740 (N_5740,N_5450,N_5261);
nand U5741 (N_5741,N_5451,N_5297);
nand U5742 (N_5742,N_5313,N_5335);
nand U5743 (N_5743,N_5487,N_5320);
or U5744 (N_5744,N_5272,N_5365);
xor U5745 (N_5745,N_5370,N_5272);
xnor U5746 (N_5746,N_5488,N_5260);
nor U5747 (N_5747,N_5283,N_5406);
xor U5748 (N_5748,N_5396,N_5380);
and U5749 (N_5749,N_5257,N_5254);
xnor U5750 (N_5750,N_5649,N_5629);
and U5751 (N_5751,N_5657,N_5637);
xnor U5752 (N_5752,N_5672,N_5506);
nor U5753 (N_5753,N_5538,N_5693);
xnor U5754 (N_5754,N_5699,N_5548);
or U5755 (N_5755,N_5733,N_5728);
nor U5756 (N_5756,N_5616,N_5668);
xor U5757 (N_5757,N_5560,N_5687);
xor U5758 (N_5758,N_5710,N_5692);
and U5759 (N_5759,N_5516,N_5583);
or U5760 (N_5760,N_5582,N_5695);
xor U5761 (N_5761,N_5594,N_5645);
or U5762 (N_5762,N_5540,N_5531);
xnor U5763 (N_5763,N_5606,N_5586);
and U5764 (N_5764,N_5669,N_5577);
xnor U5765 (N_5765,N_5743,N_5740);
nand U5766 (N_5766,N_5720,N_5737);
nor U5767 (N_5767,N_5660,N_5537);
and U5768 (N_5768,N_5524,N_5590);
and U5769 (N_5769,N_5704,N_5562);
or U5770 (N_5770,N_5559,N_5646);
nand U5771 (N_5771,N_5545,N_5510);
or U5772 (N_5772,N_5572,N_5707);
nand U5773 (N_5773,N_5689,N_5734);
and U5774 (N_5774,N_5677,N_5726);
xnor U5775 (N_5775,N_5676,N_5665);
xor U5776 (N_5776,N_5721,N_5638);
nor U5777 (N_5777,N_5662,N_5718);
nand U5778 (N_5778,N_5650,N_5534);
xor U5779 (N_5779,N_5655,N_5610);
and U5780 (N_5780,N_5744,N_5653);
nor U5781 (N_5781,N_5571,N_5711);
nor U5782 (N_5782,N_5643,N_5747);
xor U5783 (N_5783,N_5595,N_5636);
or U5784 (N_5784,N_5748,N_5741);
nor U5785 (N_5785,N_5696,N_5639);
and U5786 (N_5786,N_5719,N_5742);
or U5787 (N_5787,N_5614,N_5659);
nor U5788 (N_5788,N_5640,N_5631);
or U5789 (N_5789,N_5505,N_5714);
or U5790 (N_5790,N_5681,N_5503);
or U5791 (N_5791,N_5634,N_5680);
xnor U5792 (N_5792,N_5683,N_5561);
nand U5793 (N_5793,N_5526,N_5628);
and U5794 (N_5794,N_5557,N_5688);
and U5795 (N_5795,N_5604,N_5729);
and U5796 (N_5796,N_5591,N_5549);
nor U5797 (N_5797,N_5566,N_5554);
nor U5798 (N_5798,N_5609,N_5732);
nand U5799 (N_5799,N_5536,N_5521);
nand U5800 (N_5800,N_5602,N_5541);
or U5801 (N_5801,N_5717,N_5527);
nand U5802 (N_5802,N_5542,N_5520);
or U5803 (N_5803,N_5715,N_5546);
nand U5804 (N_5804,N_5647,N_5567);
xnor U5805 (N_5805,N_5652,N_5623);
and U5806 (N_5806,N_5556,N_5517);
nand U5807 (N_5807,N_5605,N_5598);
nand U5808 (N_5808,N_5635,N_5626);
and U5809 (N_5809,N_5608,N_5550);
and U5810 (N_5810,N_5581,N_5601);
xnor U5811 (N_5811,N_5724,N_5555);
and U5812 (N_5812,N_5619,N_5722);
and U5813 (N_5813,N_5738,N_5575);
nand U5814 (N_5814,N_5679,N_5644);
nand U5815 (N_5815,N_5745,N_5596);
and U5816 (N_5816,N_5535,N_5641);
or U5817 (N_5817,N_5576,N_5523);
xor U5818 (N_5818,N_5611,N_5731);
and U5819 (N_5819,N_5501,N_5713);
xor U5820 (N_5820,N_5735,N_5654);
nand U5821 (N_5821,N_5642,N_5603);
and U5822 (N_5822,N_5518,N_5706);
nand U5823 (N_5823,N_5727,N_5500);
or U5824 (N_5824,N_5633,N_5525);
or U5825 (N_5825,N_5589,N_5587);
or U5826 (N_5826,N_5661,N_5664);
xor U5827 (N_5827,N_5558,N_5599);
nand U5828 (N_5828,N_5612,N_5667);
xnor U5829 (N_5829,N_5564,N_5539);
and U5830 (N_5830,N_5708,N_5632);
nand U5831 (N_5831,N_5697,N_5579);
or U5832 (N_5832,N_5502,N_5716);
and U5833 (N_5833,N_5528,N_5600);
nand U5834 (N_5834,N_5585,N_5725);
nand U5835 (N_5835,N_5515,N_5673);
nand U5836 (N_5836,N_5547,N_5507);
and U5837 (N_5837,N_5705,N_5593);
and U5838 (N_5838,N_5627,N_5622);
and U5839 (N_5839,N_5618,N_5723);
nand U5840 (N_5840,N_5615,N_5573);
nor U5841 (N_5841,N_5685,N_5630);
nand U5842 (N_5842,N_5749,N_5580);
nor U5843 (N_5843,N_5511,N_5519);
or U5844 (N_5844,N_5551,N_5700);
and U5845 (N_5845,N_5621,N_5698);
and U5846 (N_5846,N_5666,N_5656);
nand U5847 (N_5847,N_5568,N_5739);
xnor U5848 (N_5848,N_5691,N_5690);
or U5849 (N_5849,N_5648,N_5709);
or U5850 (N_5850,N_5613,N_5686);
nor U5851 (N_5851,N_5684,N_5592);
or U5852 (N_5852,N_5730,N_5529);
nand U5853 (N_5853,N_5512,N_5620);
and U5854 (N_5854,N_5508,N_5565);
nand U5855 (N_5855,N_5532,N_5588);
and U5856 (N_5856,N_5682,N_5569);
xor U5857 (N_5857,N_5570,N_5509);
nand U5858 (N_5858,N_5678,N_5746);
and U5859 (N_5859,N_5504,N_5543);
and U5860 (N_5860,N_5663,N_5651);
and U5861 (N_5861,N_5530,N_5607);
or U5862 (N_5862,N_5671,N_5597);
xnor U5863 (N_5863,N_5533,N_5670);
nor U5864 (N_5864,N_5553,N_5522);
and U5865 (N_5865,N_5674,N_5578);
nor U5866 (N_5866,N_5702,N_5584);
nor U5867 (N_5867,N_5513,N_5703);
nand U5868 (N_5868,N_5624,N_5514);
and U5869 (N_5869,N_5712,N_5544);
nor U5870 (N_5870,N_5694,N_5736);
nor U5871 (N_5871,N_5617,N_5675);
or U5872 (N_5872,N_5574,N_5563);
xor U5873 (N_5873,N_5552,N_5701);
nor U5874 (N_5874,N_5658,N_5625);
nor U5875 (N_5875,N_5731,N_5721);
nand U5876 (N_5876,N_5565,N_5668);
xor U5877 (N_5877,N_5660,N_5725);
nand U5878 (N_5878,N_5529,N_5638);
xnor U5879 (N_5879,N_5701,N_5708);
or U5880 (N_5880,N_5649,N_5589);
or U5881 (N_5881,N_5579,N_5622);
xnor U5882 (N_5882,N_5581,N_5744);
or U5883 (N_5883,N_5725,N_5532);
and U5884 (N_5884,N_5694,N_5514);
nand U5885 (N_5885,N_5524,N_5729);
xnor U5886 (N_5886,N_5507,N_5743);
or U5887 (N_5887,N_5590,N_5658);
or U5888 (N_5888,N_5547,N_5572);
nand U5889 (N_5889,N_5615,N_5651);
and U5890 (N_5890,N_5678,N_5700);
and U5891 (N_5891,N_5554,N_5519);
or U5892 (N_5892,N_5549,N_5610);
nand U5893 (N_5893,N_5553,N_5605);
xnor U5894 (N_5894,N_5507,N_5573);
or U5895 (N_5895,N_5572,N_5576);
and U5896 (N_5896,N_5746,N_5581);
and U5897 (N_5897,N_5570,N_5668);
and U5898 (N_5898,N_5567,N_5717);
nor U5899 (N_5899,N_5608,N_5613);
or U5900 (N_5900,N_5564,N_5635);
nor U5901 (N_5901,N_5627,N_5541);
and U5902 (N_5902,N_5627,N_5619);
nor U5903 (N_5903,N_5699,N_5544);
xor U5904 (N_5904,N_5513,N_5681);
nand U5905 (N_5905,N_5509,N_5601);
nor U5906 (N_5906,N_5646,N_5639);
nand U5907 (N_5907,N_5625,N_5526);
nand U5908 (N_5908,N_5588,N_5525);
nand U5909 (N_5909,N_5702,N_5632);
or U5910 (N_5910,N_5571,N_5541);
or U5911 (N_5911,N_5671,N_5631);
and U5912 (N_5912,N_5623,N_5586);
xnor U5913 (N_5913,N_5703,N_5661);
and U5914 (N_5914,N_5716,N_5519);
xnor U5915 (N_5915,N_5746,N_5749);
nand U5916 (N_5916,N_5587,N_5748);
nor U5917 (N_5917,N_5525,N_5629);
or U5918 (N_5918,N_5552,N_5620);
or U5919 (N_5919,N_5628,N_5508);
xor U5920 (N_5920,N_5576,N_5559);
xor U5921 (N_5921,N_5686,N_5586);
nor U5922 (N_5922,N_5586,N_5501);
xor U5923 (N_5923,N_5572,N_5519);
nand U5924 (N_5924,N_5535,N_5682);
xor U5925 (N_5925,N_5602,N_5686);
or U5926 (N_5926,N_5570,N_5522);
xor U5927 (N_5927,N_5622,N_5724);
xnor U5928 (N_5928,N_5569,N_5611);
or U5929 (N_5929,N_5734,N_5664);
xnor U5930 (N_5930,N_5600,N_5660);
or U5931 (N_5931,N_5537,N_5595);
nand U5932 (N_5932,N_5669,N_5685);
nor U5933 (N_5933,N_5578,N_5553);
and U5934 (N_5934,N_5618,N_5667);
or U5935 (N_5935,N_5613,N_5591);
or U5936 (N_5936,N_5682,N_5503);
xnor U5937 (N_5937,N_5661,N_5611);
nand U5938 (N_5938,N_5681,N_5668);
and U5939 (N_5939,N_5627,N_5654);
or U5940 (N_5940,N_5572,N_5579);
and U5941 (N_5941,N_5675,N_5740);
nor U5942 (N_5942,N_5671,N_5540);
and U5943 (N_5943,N_5687,N_5747);
nor U5944 (N_5944,N_5689,N_5748);
nor U5945 (N_5945,N_5500,N_5618);
nor U5946 (N_5946,N_5666,N_5563);
nor U5947 (N_5947,N_5632,N_5608);
and U5948 (N_5948,N_5696,N_5607);
nand U5949 (N_5949,N_5698,N_5745);
nand U5950 (N_5950,N_5674,N_5552);
xnor U5951 (N_5951,N_5525,N_5655);
or U5952 (N_5952,N_5639,N_5678);
nand U5953 (N_5953,N_5688,N_5735);
and U5954 (N_5954,N_5614,N_5643);
or U5955 (N_5955,N_5538,N_5539);
xor U5956 (N_5956,N_5672,N_5708);
nand U5957 (N_5957,N_5557,N_5617);
xor U5958 (N_5958,N_5592,N_5742);
nand U5959 (N_5959,N_5694,N_5500);
nor U5960 (N_5960,N_5702,N_5643);
and U5961 (N_5961,N_5536,N_5740);
or U5962 (N_5962,N_5539,N_5669);
nand U5963 (N_5963,N_5717,N_5696);
xnor U5964 (N_5964,N_5681,N_5600);
and U5965 (N_5965,N_5588,N_5712);
nor U5966 (N_5966,N_5719,N_5568);
xor U5967 (N_5967,N_5587,N_5687);
and U5968 (N_5968,N_5718,N_5570);
nand U5969 (N_5969,N_5656,N_5612);
nor U5970 (N_5970,N_5506,N_5579);
or U5971 (N_5971,N_5645,N_5725);
xor U5972 (N_5972,N_5621,N_5548);
or U5973 (N_5973,N_5659,N_5639);
nor U5974 (N_5974,N_5618,N_5571);
or U5975 (N_5975,N_5632,N_5513);
nand U5976 (N_5976,N_5675,N_5574);
or U5977 (N_5977,N_5644,N_5625);
nor U5978 (N_5978,N_5656,N_5741);
and U5979 (N_5979,N_5520,N_5726);
and U5980 (N_5980,N_5742,N_5642);
and U5981 (N_5981,N_5584,N_5565);
or U5982 (N_5982,N_5574,N_5664);
nor U5983 (N_5983,N_5511,N_5740);
nor U5984 (N_5984,N_5569,N_5709);
nand U5985 (N_5985,N_5726,N_5525);
nor U5986 (N_5986,N_5682,N_5661);
or U5987 (N_5987,N_5555,N_5744);
nand U5988 (N_5988,N_5610,N_5588);
or U5989 (N_5989,N_5633,N_5531);
nand U5990 (N_5990,N_5588,N_5559);
nand U5991 (N_5991,N_5519,N_5729);
xor U5992 (N_5992,N_5654,N_5631);
and U5993 (N_5993,N_5727,N_5649);
nor U5994 (N_5994,N_5600,N_5631);
nor U5995 (N_5995,N_5677,N_5601);
and U5996 (N_5996,N_5630,N_5615);
nor U5997 (N_5997,N_5585,N_5640);
nand U5998 (N_5998,N_5552,N_5536);
and U5999 (N_5999,N_5745,N_5682);
or U6000 (N_6000,N_5750,N_5886);
or U6001 (N_6001,N_5773,N_5932);
or U6002 (N_6002,N_5978,N_5839);
xnor U6003 (N_6003,N_5926,N_5766);
nor U6004 (N_6004,N_5816,N_5825);
and U6005 (N_6005,N_5836,N_5865);
nor U6006 (N_6006,N_5866,N_5795);
xnor U6007 (N_6007,N_5972,N_5986);
xnor U6008 (N_6008,N_5798,N_5939);
nand U6009 (N_6009,N_5899,N_5950);
xnor U6010 (N_6010,N_5873,N_5820);
nor U6011 (N_6011,N_5810,N_5760);
xor U6012 (N_6012,N_5813,N_5955);
or U6013 (N_6013,N_5883,N_5753);
nand U6014 (N_6014,N_5974,N_5888);
or U6015 (N_6015,N_5912,N_5847);
or U6016 (N_6016,N_5826,N_5982);
or U6017 (N_6017,N_5992,N_5880);
xnor U6018 (N_6018,N_5889,N_5918);
nand U6019 (N_6019,N_5917,N_5896);
or U6020 (N_6020,N_5925,N_5962);
nand U6021 (N_6021,N_5764,N_5990);
or U6022 (N_6022,N_5811,N_5854);
nand U6023 (N_6023,N_5954,N_5775);
xor U6024 (N_6024,N_5940,N_5969);
nand U6025 (N_6025,N_5961,N_5770);
nor U6026 (N_6026,N_5752,N_5882);
nor U6027 (N_6027,N_5759,N_5995);
xnor U6028 (N_6028,N_5834,N_5861);
or U6029 (N_6029,N_5762,N_5853);
xor U6030 (N_6030,N_5920,N_5944);
xnor U6031 (N_6031,N_5797,N_5876);
nand U6032 (N_6032,N_5779,N_5862);
and U6033 (N_6033,N_5817,N_5870);
nor U6034 (N_6034,N_5914,N_5821);
nand U6035 (N_6035,N_5989,N_5943);
nor U6036 (N_6036,N_5791,N_5987);
or U6037 (N_6037,N_5942,N_5868);
xnor U6038 (N_6038,N_5806,N_5966);
nor U6039 (N_6039,N_5808,N_5963);
xnor U6040 (N_6040,N_5900,N_5823);
or U6041 (N_6041,N_5938,N_5941);
nand U6042 (N_6042,N_5780,N_5828);
nand U6043 (N_6043,N_5934,N_5754);
or U6044 (N_6044,N_5848,N_5913);
or U6045 (N_6045,N_5971,N_5879);
nor U6046 (N_6046,N_5787,N_5875);
nor U6047 (N_6047,N_5906,N_5796);
xor U6048 (N_6048,N_5909,N_5884);
nand U6049 (N_6049,N_5860,N_5818);
or U6050 (N_6050,N_5793,N_5977);
or U6051 (N_6051,N_5758,N_5965);
or U6052 (N_6052,N_5790,N_5778);
nand U6053 (N_6053,N_5960,N_5985);
and U6054 (N_6054,N_5857,N_5894);
or U6055 (N_6055,N_5785,N_5864);
nor U6056 (N_6056,N_5949,N_5973);
or U6057 (N_6057,N_5908,N_5933);
and U6058 (N_6058,N_5794,N_5975);
and U6059 (N_6059,N_5831,N_5792);
nand U6060 (N_6060,N_5997,N_5991);
nor U6061 (N_6061,N_5801,N_5807);
nand U6062 (N_6062,N_5755,N_5852);
nand U6063 (N_6063,N_5980,N_5893);
and U6064 (N_6064,N_5936,N_5910);
xor U6065 (N_6065,N_5769,N_5911);
nor U6066 (N_6066,N_5763,N_5885);
and U6067 (N_6067,N_5895,N_5903);
or U6068 (N_6068,N_5871,N_5907);
nand U6069 (N_6069,N_5856,N_5843);
nand U6070 (N_6070,N_5835,N_5803);
and U6071 (N_6071,N_5959,N_5859);
nand U6072 (N_6072,N_5776,N_5984);
and U6073 (N_6073,N_5953,N_5771);
or U6074 (N_6074,N_5999,N_5858);
nor U6075 (N_6075,N_5842,N_5877);
nor U6076 (N_6076,N_5849,N_5872);
xnor U6077 (N_6077,N_5976,N_5761);
or U6078 (N_6078,N_5952,N_5830);
nand U6079 (N_6079,N_5838,N_5822);
nand U6080 (N_6080,N_5892,N_5781);
or U6081 (N_6081,N_5947,N_5994);
nand U6082 (N_6082,N_5767,N_5874);
and U6083 (N_6083,N_5833,N_5996);
nor U6084 (N_6084,N_5802,N_5964);
and U6085 (N_6085,N_5805,N_5891);
nand U6086 (N_6086,N_5841,N_5921);
nor U6087 (N_6087,N_5829,N_5897);
nand U6088 (N_6088,N_5824,N_5869);
and U6089 (N_6089,N_5804,N_5931);
and U6090 (N_6090,N_5840,N_5774);
and U6091 (N_6091,N_5956,N_5902);
xor U6092 (N_6092,N_5898,N_5846);
nand U6093 (N_6093,N_5772,N_5878);
or U6094 (N_6094,N_5786,N_5788);
nor U6095 (N_6095,N_5887,N_5916);
nor U6096 (N_6096,N_5901,N_5845);
nand U6097 (N_6097,N_5957,N_5777);
nor U6098 (N_6098,N_5945,N_5765);
nand U6099 (N_6099,N_5812,N_5930);
nor U6100 (N_6100,N_5890,N_5783);
nor U6101 (N_6101,N_5979,N_5948);
nand U6102 (N_6102,N_5850,N_5928);
and U6103 (N_6103,N_5867,N_5915);
nor U6104 (N_6104,N_5951,N_5981);
nor U6105 (N_6105,N_5929,N_5968);
and U6106 (N_6106,N_5855,N_5827);
and U6107 (N_6107,N_5782,N_5881);
nand U6108 (N_6108,N_5844,N_5993);
xnor U6109 (N_6109,N_5927,N_5751);
nand U6110 (N_6110,N_5768,N_5757);
nor U6111 (N_6111,N_5919,N_5799);
nor U6112 (N_6112,N_5988,N_5904);
and U6113 (N_6113,N_5922,N_5935);
nor U6114 (N_6114,N_5784,N_5837);
and U6115 (N_6115,N_5998,N_5789);
nand U6116 (N_6116,N_5923,N_5814);
nor U6117 (N_6117,N_5970,N_5937);
or U6118 (N_6118,N_5924,N_5863);
and U6119 (N_6119,N_5832,N_5851);
nand U6120 (N_6120,N_5809,N_5756);
xnor U6121 (N_6121,N_5819,N_5800);
nand U6122 (N_6122,N_5967,N_5946);
xor U6123 (N_6123,N_5815,N_5983);
nor U6124 (N_6124,N_5905,N_5958);
nand U6125 (N_6125,N_5946,N_5876);
nand U6126 (N_6126,N_5838,N_5764);
nand U6127 (N_6127,N_5959,N_5905);
xor U6128 (N_6128,N_5839,N_5949);
nor U6129 (N_6129,N_5986,N_5845);
nor U6130 (N_6130,N_5990,N_5974);
and U6131 (N_6131,N_5978,N_5764);
nand U6132 (N_6132,N_5980,N_5990);
nand U6133 (N_6133,N_5870,N_5781);
xor U6134 (N_6134,N_5812,N_5919);
xnor U6135 (N_6135,N_5999,N_5846);
and U6136 (N_6136,N_5989,N_5964);
nor U6137 (N_6137,N_5870,N_5990);
nand U6138 (N_6138,N_5860,N_5973);
xnor U6139 (N_6139,N_5787,N_5926);
or U6140 (N_6140,N_5907,N_5903);
nand U6141 (N_6141,N_5923,N_5845);
xnor U6142 (N_6142,N_5765,N_5891);
xnor U6143 (N_6143,N_5938,N_5848);
or U6144 (N_6144,N_5930,N_5958);
nor U6145 (N_6145,N_5972,N_5765);
and U6146 (N_6146,N_5969,N_5818);
nand U6147 (N_6147,N_5832,N_5915);
xnor U6148 (N_6148,N_5939,N_5829);
or U6149 (N_6149,N_5777,N_5986);
xor U6150 (N_6150,N_5771,N_5937);
and U6151 (N_6151,N_5970,N_5802);
or U6152 (N_6152,N_5846,N_5883);
or U6153 (N_6153,N_5931,N_5932);
nand U6154 (N_6154,N_5756,N_5827);
xor U6155 (N_6155,N_5891,N_5961);
nand U6156 (N_6156,N_5826,N_5757);
xor U6157 (N_6157,N_5963,N_5905);
and U6158 (N_6158,N_5781,N_5945);
nand U6159 (N_6159,N_5988,N_5790);
nor U6160 (N_6160,N_5801,N_5825);
nand U6161 (N_6161,N_5854,N_5766);
or U6162 (N_6162,N_5973,N_5862);
and U6163 (N_6163,N_5826,N_5890);
nand U6164 (N_6164,N_5835,N_5799);
and U6165 (N_6165,N_5879,N_5794);
or U6166 (N_6166,N_5764,N_5996);
nor U6167 (N_6167,N_5914,N_5789);
and U6168 (N_6168,N_5953,N_5885);
and U6169 (N_6169,N_5922,N_5796);
xor U6170 (N_6170,N_5887,N_5787);
nand U6171 (N_6171,N_5826,N_5842);
nor U6172 (N_6172,N_5915,N_5784);
nand U6173 (N_6173,N_5781,N_5826);
xnor U6174 (N_6174,N_5967,N_5933);
xor U6175 (N_6175,N_5817,N_5959);
nand U6176 (N_6176,N_5753,N_5875);
nor U6177 (N_6177,N_5988,N_5797);
xor U6178 (N_6178,N_5989,N_5907);
and U6179 (N_6179,N_5985,N_5778);
xnor U6180 (N_6180,N_5939,N_5934);
nor U6181 (N_6181,N_5812,N_5960);
and U6182 (N_6182,N_5911,N_5898);
nand U6183 (N_6183,N_5805,N_5857);
nand U6184 (N_6184,N_5784,N_5820);
xnor U6185 (N_6185,N_5761,N_5909);
nand U6186 (N_6186,N_5849,N_5901);
and U6187 (N_6187,N_5771,N_5922);
nor U6188 (N_6188,N_5871,N_5878);
nor U6189 (N_6189,N_5997,N_5928);
xor U6190 (N_6190,N_5895,N_5842);
xnor U6191 (N_6191,N_5779,N_5826);
nor U6192 (N_6192,N_5824,N_5975);
and U6193 (N_6193,N_5872,N_5892);
and U6194 (N_6194,N_5909,N_5842);
and U6195 (N_6195,N_5861,N_5935);
nand U6196 (N_6196,N_5778,N_5776);
nor U6197 (N_6197,N_5978,N_5953);
or U6198 (N_6198,N_5837,N_5850);
and U6199 (N_6199,N_5846,N_5796);
nor U6200 (N_6200,N_5810,N_5946);
xor U6201 (N_6201,N_5919,N_5878);
or U6202 (N_6202,N_5891,N_5771);
nor U6203 (N_6203,N_5983,N_5942);
or U6204 (N_6204,N_5989,N_5769);
and U6205 (N_6205,N_5984,N_5891);
xnor U6206 (N_6206,N_5955,N_5866);
or U6207 (N_6207,N_5750,N_5997);
nor U6208 (N_6208,N_5894,N_5905);
xnor U6209 (N_6209,N_5952,N_5856);
xor U6210 (N_6210,N_5876,N_5828);
nand U6211 (N_6211,N_5779,N_5903);
xor U6212 (N_6212,N_5848,N_5957);
xor U6213 (N_6213,N_5892,N_5956);
or U6214 (N_6214,N_5985,N_5879);
nand U6215 (N_6215,N_5858,N_5853);
and U6216 (N_6216,N_5975,N_5895);
nor U6217 (N_6217,N_5948,N_5982);
and U6218 (N_6218,N_5760,N_5921);
or U6219 (N_6219,N_5891,N_5811);
or U6220 (N_6220,N_5990,N_5883);
nor U6221 (N_6221,N_5792,N_5946);
and U6222 (N_6222,N_5778,N_5770);
nand U6223 (N_6223,N_5840,N_5833);
and U6224 (N_6224,N_5984,N_5854);
or U6225 (N_6225,N_5937,N_5825);
or U6226 (N_6226,N_5756,N_5819);
or U6227 (N_6227,N_5913,N_5917);
nor U6228 (N_6228,N_5788,N_5805);
or U6229 (N_6229,N_5764,N_5788);
nand U6230 (N_6230,N_5783,N_5826);
and U6231 (N_6231,N_5838,N_5863);
nand U6232 (N_6232,N_5776,N_5756);
nand U6233 (N_6233,N_5838,N_5888);
nor U6234 (N_6234,N_5789,N_5969);
nor U6235 (N_6235,N_5991,N_5779);
nor U6236 (N_6236,N_5936,N_5973);
or U6237 (N_6237,N_5926,N_5884);
nor U6238 (N_6238,N_5921,N_5909);
nor U6239 (N_6239,N_5840,N_5771);
and U6240 (N_6240,N_5997,N_5752);
and U6241 (N_6241,N_5929,N_5874);
and U6242 (N_6242,N_5766,N_5871);
nor U6243 (N_6243,N_5938,N_5821);
nor U6244 (N_6244,N_5795,N_5820);
or U6245 (N_6245,N_5894,N_5914);
or U6246 (N_6246,N_5962,N_5814);
nand U6247 (N_6247,N_5926,N_5898);
and U6248 (N_6248,N_5983,N_5840);
nor U6249 (N_6249,N_5914,N_5961);
or U6250 (N_6250,N_6230,N_6078);
or U6251 (N_6251,N_6243,N_6119);
nand U6252 (N_6252,N_6169,N_6132);
xnor U6253 (N_6253,N_6166,N_6070);
and U6254 (N_6254,N_6120,N_6084);
nor U6255 (N_6255,N_6223,N_6147);
and U6256 (N_6256,N_6200,N_6106);
nor U6257 (N_6257,N_6046,N_6179);
nor U6258 (N_6258,N_6074,N_6193);
or U6259 (N_6259,N_6091,N_6064);
nand U6260 (N_6260,N_6054,N_6210);
nor U6261 (N_6261,N_6159,N_6066);
and U6262 (N_6262,N_6211,N_6118);
nand U6263 (N_6263,N_6206,N_6012);
nand U6264 (N_6264,N_6142,N_6201);
nor U6265 (N_6265,N_6103,N_6027);
nand U6266 (N_6266,N_6010,N_6226);
and U6267 (N_6267,N_6059,N_6144);
xnor U6268 (N_6268,N_6067,N_6031);
nor U6269 (N_6269,N_6021,N_6129);
or U6270 (N_6270,N_6182,N_6140);
xor U6271 (N_6271,N_6073,N_6008);
and U6272 (N_6272,N_6057,N_6022);
xnor U6273 (N_6273,N_6168,N_6137);
and U6274 (N_6274,N_6128,N_6075);
nor U6275 (N_6275,N_6247,N_6018);
nor U6276 (N_6276,N_6245,N_6062);
nand U6277 (N_6277,N_6162,N_6056);
and U6278 (N_6278,N_6122,N_6149);
nor U6279 (N_6279,N_6160,N_6170);
nand U6280 (N_6280,N_6101,N_6096);
nor U6281 (N_6281,N_6152,N_6072);
xor U6282 (N_6282,N_6024,N_6034);
and U6283 (N_6283,N_6171,N_6089);
xnor U6284 (N_6284,N_6131,N_6231);
or U6285 (N_6285,N_6048,N_6183);
xnor U6286 (N_6286,N_6248,N_6215);
and U6287 (N_6287,N_6081,N_6164);
or U6288 (N_6288,N_6055,N_6115);
and U6289 (N_6289,N_6172,N_6069);
nand U6290 (N_6290,N_6232,N_6205);
or U6291 (N_6291,N_6195,N_6090);
xor U6292 (N_6292,N_6176,N_6203);
and U6293 (N_6293,N_6039,N_6020);
nor U6294 (N_6294,N_6228,N_6117);
nor U6295 (N_6295,N_6102,N_6240);
nor U6296 (N_6296,N_6212,N_6030);
xnor U6297 (N_6297,N_6001,N_6032);
xor U6298 (N_6298,N_6098,N_6040);
nor U6299 (N_6299,N_6038,N_6107);
nor U6300 (N_6300,N_6173,N_6130);
or U6301 (N_6301,N_6229,N_6016);
and U6302 (N_6302,N_6246,N_6007);
or U6303 (N_6303,N_6043,N_6121);
nor U6304 (N_6304,N_6002,N_6224);
and U6305 (N_6305,N_6242,N_6004);
nor U6306 (N_6306,N_6216,N_6109);
and U6307 (N_6307,N_6123,N_6041);
xnor U6308 (N_6308,N_6196,N_6003);
xnor U6309 (N_6309,N_6023,N_6093);
nand U6310 (N_6310,N_6187,N_6092);
nand U6311 (N_6311,N_6134,N_6053);
and U6312 (N_6312,N_6127,N_6026);
or U6313 (N_6313,N_6049,N_6214);
or U6314 (N_6314,N_6197,N_6204);
nor U6315 (N_6315,N_6082,N_6151);
and U6316 (N_6316,N_6085,N_6236);
nor U6317 (N_6317,N_6194,N_6114);
or U6318 (N_6318,N_6153,N_6156);
nor U6319 (N_6319,N_6241,N_6225);
or U6320 (N_6320,N_6088,N_6178);
xnor U6321 (N_6321,N_6037,N_6198);
xor U6322 (N_6322,N_6108,N_6163);
nand U6323 (N_6323,N_6219,N_6086);
and U6324 (N_6324,N_6113,N_6079);
and U6325 (N_6325,N_6011,N_6150);
xor U6326 (N_6326,N_6235,N_6063);
or U6327 (N_6327,N_6139,N_6009);
nand U6328 (N_6328,N_6174,N_6244);
and U6329 (N_6329,N_6000,N_6154);
nor U6330 (N_6330,N_6076,N_6110);
nand U6331 (N_6331,N_6035,N_6047);
nor U6332 (N_6332,N_6014,N_6133);
xnor U6333 (N_6333,N_6185,N_6068);
nand U6334 (N_6334,N_6017,N_6180);
and U6335 (N_6335,N_6061,N_6050);
or U6336 (N_6336,N_6165,N_6015);
xor U6337 (N_6337,N_6238,N_6029);
xnor U6338 (N_6338,N_6124,N_6157);
nor U6339 (N_6339,N_6135,N_6148);
or U6340 (N_6340,N_6143,N_6005);
xnor U6341 (N_6341,N_6071,N_6138);
and U6342 (N_6342,N_6104,N_6141);
xor U6343 (N_6343,N_6190,N_6094);
nor U6344 (N_6344,N_6249,N_6186);
nand U6345 (N_6345,N_6234,N_6207);
xnor U6346 (N_6346,N_6060,N_6233);
nand U6347 (N_6347,N_6051,N_6100);
or U6348 (N_6348,N_6202,N_6136);
nor U6349 (N_6349,N_6237,N_6036);
xnor U6350 (N_6350,N_6158,N_6227);
and U6351 (N_6351,N_6217,N_6112);
nand U6352 (N_6352,N_6083,N_6145);
nand U6353 (N_6353,N_6058,N_6191);
nand U6354 (N_6354,N_6044,N_6006);
nor U6355 (N_6355,N_6189,N_6221);
nand U6356 (N_6356,N_6013,N_6218);
or U6357 (N_6357,N_6019,N_6188);
and U6358 (N_6358,N_6220,N_6146);
or U6359 (N_6359,N_6167,N_6116);
nor U6360 (N_6360,N_6045,N_6239);
xor U6361 (N_6361,N_6080,N_6161);
nand U6362 (N_6362,N_6095,N_6097);
and U6363 (N_6363,N_6105,N_6177);
and U6364 (N_6364,N_6199,N_6052);
nand U6365 (N_6365,N_6181,N_6099);
and U6366 (N_6366,N_6125,N_6077);
nor U6367 (N_6367,N_6033,N_6209);
and U6368 (N_6368,N_6126,N_6192);
nor U6369 (N_6369,N_6175,N_6065);
nand U6370 (N_6370,N_6213,N_6155);
nand U6371 (N_6371,N_6042,N_6184);
nor U6372 (N_6372,N_6208,N_6222);
nand U6373 (N_6373,N_6111,N_6025);
xnor U6374 (N_6374,N_6087,N_6028);
and U6375 (N_6375,N_6111,N_6108);
or U6376 (N_6376,N_6223,N_6148);
xnor U6377 (N_6377,N_6114,N_6032);
and U6378 (N_6378,N_6226,N_6216);
nor U6379 (N_6379,N_6083,N_6208);
nand U6380 (N_6380,N_6189,N_6004);
or U6381 (N_6381,N_6063,N_6218);
and U6382 (N_6382,N_6220,N_6111);
xor U6383 (N_6383,N_6092,N_6234);
xor U6384 (N_6384,N_6154,N_6224);
nand U6385 (N_6385,N_6078,N_6113);
nand U6386 (N_6386,N_6139,N_6088);
nand U6387 (N_6387,N_6220,N_6095);
and U6388 (N_6388,N_6022,N_6228);
and U6389 (N_6389,N_6106,N_6022);
xnor U6390 (N_6390,N_6232,N_6144);
nand U6391 (N_6391,N_6202,N_6106);
xor U6392 (N_6392,N_6022,N_6027);
nor U6393 (N_6393,N_6145,N_6238);
xnor U6394 (N_6394,N_6242,N_6129);
nand U6395 (N_6395,N_6216,N_6053);
and U6396 (N_6396,N_6064,N_6196);
and U6397 (N_6397,N_6104,N_6197);
or U6398 (N_6398,N_6219,N_6173);
or U6399 (N_6399,N_6112,N_6155);
and U6400 (N_6400,N_6108,N_6222);
and U6401 (N_6401,N_6125,N_6055);
xnor U6402 (N_6402,N_6022,N_6070);
and U6403 (N_6403,N_6228,N_6220);
nor U6404 (N_6404,N_6042,N_6098);
nor U6405 (N_6405,N_6243,N_6114);
nor U6406 (N_6406,N_6207,N_6142);
and U6407 (N_6407,N_6215,N_6011);
or U6408 (N_6408,N_6019,N_6245);
and U6409 (N_6409,N_6036,N_6180);
and U6410 (N_6410,N_6157,N_6229);
and U6411 (N_6411,N_6157,N_6210);
or U6412 (N_6412,N_6161,N_6091);
xnor U6413 (N_6413,N_6040,N_6136);
and U6414 (N_6414,N_6093,N_6081);
and U6415 (N_6415,N_6024,N_6022);
or U6416 (N_6416,N_6216,N_6242);
or U6417 (N_6417,N_6056,N_6051);
nor U6418 (N_6418,N_6082,N_6200);
xor U6419 (N_6419,N_6116,N_6213);
and U6420 (N_6420,N_6050,N_6132);
and U6421 (N_6421,N_6041,N_6181);
or U6422 (N_6422,N_6158,N_6109);
xnor U6423 (N_6423,N_6054,N_6115);
nor U6424 (N_6424,N_6127,N_6039);
or U6425 (N_6425,N_6083,N_6020);
nand U6426 (N_6426,N_6087,N_6080);
nand U6427 (N_6427,N_6203,N_6168);
xnor U6428 (N_6428,N_6187,N_6229);
and U6429 (N_6429,N_6235,N_6101);
xor U6430 (N_6430,N_6238,N_6001);
xnor U6431 (N_6431,N_6029,N_6242);
and U6432 (N_6432,N_6198,N_6233);
nand U6433 (N_6433,N_6238,N_6178);
xor U6434 (N_6434,N_6074,N_6136);
nand U6435 (N_6435,N_6172,N_6203);
and U6436 (N_6436,N_6047,N_6012);
and U6437 (N_6437,N_6214,N_6098);
xor U6438 (N_6438,N_6221,N_6213);
xor U6439 (N_6439,N_6216,N_6061);
or U6440 (N_6440,N_6071,N_6065);
nand U6441 (N_6441,N_6203,N_6059);
nor U6442 (N_6442,N_6056,N_6101);
xnor U6443 (N_6443,N_6223,N_6189);
nor U6444 (N_6444,N_6249,N_6167);
nand U6445 (N_6445,N_6077,N_6144);
and U6446 (N_6446,N_6049,N_6238);
and U6447 (N_6447,N_6082,N_6110);
xor U6448 (N_6448,N_6154,N_6094);
xnor U6449 (N_6449,N_6014,N_6105);
nor U6450 (N_6450,N_6181,N_6093);
or U6451 (N_6451,N_6227,N_6144);
nor U6452 (N_6452,N_6228,N_6024);
xnor U6453 (N_6453,N_6093,N_6242);
nor U6454 (N_6454,N_6095,N_6033);
or U6455 (N_6455,N_6116,N_6124);
xnor U6456 (N_6456,N_6058,N_6053);
xor U6457 (N_6457,N_6023,N_6016);
xnor U6458 (N_6458,N_6034,N_6204);
or U6459 (N_6459,N_6106,N_6026);
nand U6460 (N_6460,N_6077,N_6212);
or U6461 (N_6461,N_6003,N_6139);
or U6462 (N_6462,N_6074,N_6210);
and U6463 (N_6463,N_6127,N_6234);
and U6464 (N_6464,N_6057,N_6085);
xor U6465 (N_6465,N_6209,N_6095);
or U6466 (N_6466,N_6197,N_6054);
and U6467 (N_6467,N_6015,N_6049);
xnor U6468 (N_6468,N_6060,N_6021);
xor U6469 (N_6469,N_6013,N_6130);
and U6470 (N_6470,N_6077,N_6105);
xor U6471 (N_6471,N_6042,N_6030);
and U6472 (N_6472,N_6148,N_6053);
and U6473 (N_6473,N_6051,N_6172);
and U6474 (N_6474,N_6187,N_6131);
or U6475 (N_6475,N_6006,N_6202);
nor U6476 (N_6476,N_6227,N_6089);
or U6477 (N_6477,N_6194,N_6119);
nand U6478 (N_6478,N_6032,N_6103);
and U6479 (N_6479,N_6127,N_6036);
and U6480 (N_6480,N_6051,N_6037);
nor U6481 (N_6481,N_6152,N_6043);
nand U6482 (N_6482,N_6030,N_6092);
and U6483 (N_6483,N_6057,N_6002);
nand U6484 (N_6484,N_6090,N_6086);
nor U6485 (N_6485,N_6031,N_6151);
nor U6486 (N_6486,N_6020,N_6172);
or U6487 (N_6487,N_6024,N_6178);
or U6488 (N_6488,N_6025,N_6090);
nand U6489 (N_6489,N_6074,N_6060);
nand U6490 (N_6490,N_6059,N_6036);
nor U6491 (N_6491,N_6235,N_6105);
and U6492 (N_6492,N_6116,N_6054);
nand U6493 (N_6493,N_6063,N_6009);
and U6494 (N_6494,N_6034,N_6239);
or U6495 (N_6495,N_6223,N_6153);
nand U6496 (N_6496,N_6101,N_6219);
nand U6497 (N_6497,N_6101,N_6015);
nand U6498 (N_6498,N_6092,N_6080);
and U6499 (N_6499,N_6014,N_6145);
nand U6500 (N_6500,N_6353,N_6319);
nand U6501 (N_6501,N_6451,N_6474);
nand U6502 (N_6502,N_6328,N_6271);
and U6503 (N_6503,N_6481,N_6396);
nand U6504 (N_6504,N_6416,N_6358);
nand U6505 (N_6505,N_6432,N_6305);
nor U6506 (N_6506,N_6356,N_6361);
nand U6507 (N_6507,N_6255,N_6311);
or U6508 (N_6508,N_6286,N_6307);
and U6509 (N_6509,N_6440,N_6395);
nor U6510 (N_6510,N_6326,N_6420);
xnor U6511 (N_6511,N_6265,N_6346);
nor U6512 (N_6512,N_6300,N_6471);
xor U6513 (N_6513,N_6386,N_6428);
or U6514 (N_6514,N_6270,N_6272);
nand U6515 (N_6515,N_6350,N_6450);
nor U6516 (N_6516,N_6308,N_6366);
xor U6517 (N_6517,N_6302,N_6339);
xor U6518 (N_6518,N_6313,N_6377);
nor U6519 (N_6519,N_6466,N_6261);
or U6520 (N_6520,N_6490,N_6390);
nor U6521 (N_6521,N_6409,N_6289);
xnor U6522 (N_6522,N_6306,N_6441);
nand U6523 (N_6523,N_6483,N_6403);
nor U6524 (N_6524,N_6340,N_6381);
nand U6525 (N_6525,N_6426,N_6299);
and U6526 (N_6526,N_6318,N_6359);
and U6527 (N_6527,N_6349,N_6292);
or U6528 (N_6528,N_6448,N_6297);
or U6529 (N_6529,N_6452,N_6369);
xnor U6530 (N_6530,N_6257,N_6430);
or U6531 (N_6531,N_6410,N_6417);
or U6532 (N_6532,N_6316,N_6472);
nand U6533 (N_6533,N_6400,N_6365);
nand U6534 (N_6534,N_6315,N_6388);
or U6535 (N_6535,N_6424,N_6415);
nor U6536 (N_6536,N_6372,N_6293);
xnor U6537 (N_6537,N_6476,N_6348);
xor U6538 (N_6538,N_6274,N_6276);
nor U6539 (N_6539,N_6263,N_6370);
xnor U6540 (N_6540,N_6277,N_6254);
xnor U6541 (N_6541,N_6378,N_6433);
nor U6542 (N_6542,N_6488,N_6492);
nor U6543 (N_6543,N_6320,N_6465);
or U6544 (N_6544,N_6491,N_6477);
or U6545 (N_6545,N_6458,N_6411);
or U6546 (N_6546,N_6312,N_6499);
nor U6547 (N_6547,N_6327,N_6489);
nor U6548 (N_6548,N_6285,N_6262);
nor U6549 (N_6549,N_6427,N_6473);
and U6550 (N_6550,N_6280,N_6434);
xor U6551 (N_6551,N_6342,N_6368);
or U6552 (N_6552,N_6383,N_6329);
and U6553 (N_6553,N_6495,N_6301);
or U6554 (N_6554,N_6414,N_6494);
nor U6555 (N_6555,N_6418,N_6475);
xnor U6556 (N_6556,N_6384,N_6407);
xor U6557 (N_6557,N_6404,N_6406);
and U6558 (N_6558,N_6429,N_6455);
nand U6559 (N_6559,N_6282,N_6290);
xor U6560 (N_6560,N_6486,N_6324);
nor U6561 (N_6561,N_6298,N_6291);
or U6562 (N_6562,N_6253,N_6281);
or U6563 (N_6563,N_6493,N_6460);
or U6564 (N_6564,N_6457,N_6397);
or U6565 (N_6565,N_6408,N_6338);
and U6566 (N_6566,N_6337,N_6480);
xor U6567 (N_6567,N_6273,N_6449);
nand U6568 (N_6568,N_6445,N_6421);
and U6569 (N_6569,N_6374,N_6347);
nand U6570 (N_6570,N_6487,N_6354);
nor U6571 (N_6571,N_6321,N_6322);
or U6572 (N_6572,N_6341,N_6278);
xor U6573 (N_6573,N_6267,N_6352);
nor U6574 (N_6574,N_6325,N_6398);
and U6575 (N_6575,N_6367,N_6317);
xor U6576 (N_6576,N_6351,N_6334);
xnor U6577 (N_6577,N_6382,N_6453);
xnor U6578 (N_6578,N_6463,N_6444);
or U6579 (N_6579,N_6288,N_6331);
and U6580 (N_6580,N_6484,N_6284);
and U6581 (N_6581,N_6363,N_6387);
and U6582 (N_6582,N_6443,N_6468);
nand U6583 (N_6583,N_6375,N_6345);
nor U6584 (N_6584,N_6268,N_6258);
or U6585 (N_6585,N_6462,N_6467);
or U6586 (N_6586,N_6309,N_6412);
and U6587 (N_6587,N_6287,N_6402);
nand U6588 (N_6588,N_6413,N_6330);
nor U6589 (N_6589,N_6269,N_6360);
or U6590 (N_6590,N_6436,N_6393);
xnor U6591 (N_6591,N_6454,N_6431);
xnor U6592 (N_6592,N_6379,N_6335);
or U6593 (N_6593,N_6438,N_6394);
and U6594 (N_6594,N_6362,N_6470);
nand U6595 (N_6595,N_6279,N_6251);
or U6596 (N_6596,N_6422,N_6447);
or U6597 (N_6597,N_6295,N_6399);
nor U6598 (N_6598,N_6391,N_6283);
nor U6599 (N_6599,N_6498,N_6419);
nor U6600 (N_6600,N_6380,N_6266);
or U6601 (N_6601,N_6343,N_6435);
nor U6602 (N_6602,N_6459,N_6344);
nor U6603 (N_6603,N_6259,N_6425);
or U6604 (N_6604,N_6478,N_6442);
xnor U6605 (N_6605,N_6264,N_6439);
and U6606 (N_6606,N_6355,N_6485);
nand U6607 (N_6607,N_6275,N_6250);
or U6608 (N_6608,N_6310,N_6336);
and U6609 (N_6609,N_6437,N_6461);
or U6610 (N_6610,N_6479,N_6497);
and U6611 (N_6611,N_6252,N_6373);
nand U6612 (N_6612,N_6323,N_6296);
xor U6613 (N_6613,N_6256,N_6496);
and U6614 (N_6614,N_6385,N_6401);
nand U6615 (N_6615,N_6446,N_6333);
or U6616 (N_6616,N_6456,N_6389);
nor U6617 (N_6617,N_6357,N_6423);
nand U6618 (N_6618,N_6405,N_6464);
nor U6619 (N_6619,N_6376,N_6304);
nand U6620 (N_6620,N_6469,N_6371);
or U6621 (N_6621,N_6482,N_6332);
nand U6622 (N_6622,N_6314,N_6392);
and U6623 (N_6623,N_6364,N_6294);
nor U6624 (N_6624,N_6260,N_6303);
and U6625 (N_6625,N_6455,N_6258);
or U6626 (N_6626,N_6323,N_6391);
nor U6627 (N_6627,N_6309,N_6413);
nor U6628 (N_6628,N_6455,N_6413);
or U6629 (N_6629,N_6369,N_6425);
and U6630 (N_6630,N_6400,N_6492);
and U6631 (N_6631,N_6271,N_6429);
nor U6632 (N_6632,N_6250,N_6489);
nor U6633 (N_6633,N_6259,N_6352);
nand U6634 (N_6634,N_6329,N_6483);
and U6635 (N_6635,N_6320,N_6346);
nand U6636 (N_6636,N_6323,N_6439);
nor U6637 (N_6637,N_6371,N_6313);
nand U6638 (N_6638,N_6399,N_6457);
nand U6639 (N_6639,N_6387,N_6291);
xnor U6640 (N_6640,N_6303,N_6326);
or U6641 (N_6641,N_6287,N_6385);
and U6642 (N_6642,N_6305,N_6412);
and U6643 (N_6643,N_6314,N_6356);
xor U6644 (N_6644,N_6454,N_6262);
xnor U6645 (N_6645,N_6486,N_6314);
nand U6646 (N_6646,N_6487,N_6472);
xnor U6647 (N_6647,N_6349,N_6314);
and U6648 (N_6648,N_6431,N_6288);
nor U6649 (N_6649,N_6326,N_6252);
or U6650 (N_6650,N_6354,N_6260);
or U6651 (N_6651,N_6315,N_6497);
nand U6652 (N_6652,N_6439,N_6332);
and U6653 (N_6653,N_6407,N_6252);
or U6654 (N_6654,N_6329,N_6349);
xnor U6655 (N_6655,N_6482,N_6357);
nor U6656 (N_6656,N_6388,N_6301);
and U6657 (N_6657,N_6331,N_6430);
and U6658 (N_6658,N_6284,N_6331);
and U6659 (N_6659,N_6478,N_6416);
and U6660 (N_6660,N_6294,N_6269);
xnor U6661 (N_6661,N_6306,N_6374);
or U6662 (N_6662,N_6255,N_6284);
and U6663 (N_6663,N_6287,N_6474);
or U6664 (N_6664,N_6396,N_6267);
nor U6665 (N_6665,N_6374,N_6468);
nand U6666 (N_6666,N_6264,N_6408);
xnor U6667 (N_6667,N_6308,N_6401);
nand U6668 (N_6668,N_6461,N_6444);
xor U6669 (N_6669,N_6265,N_6494);
or U6670 (N_6670,N_6340,N_6368);
nand U6671 (N_6671,N_6441,N_6423);
or U6672 (N_6672,N_6437,N_6464);
and U6673 (N_6673,N_6368,N_6262);
and U6674 (N_6674,N_6305,N_6339);
or U6675 (N_6675,N_6415,N_6414);
and U6676 (N_6676,N_6397,N_6315);
nor U6677 (N_6677,N_6322,N_6425);
nor U6678 (N_6678,N_6489,N_6432);
nor U6679 (N_6679,N_6410,N_6393);
xnor U6680 (N_6680,N_6255,N_6398);
nor U6681 (N_6681,N_6495,N_6334);
and U6682 (N_6682,N_6250,N_6273);
or U6683 (N_6683,N_6388,N_6342);
nand U6684 (N_6684,N_6381,N_6373);
and U6685 (N_6685,N_6428,N_6395);
and U6686 (N_6686,N_6333,N_6433);
or U6687 (N_6687,N_6351,N_6366);
xor U6688 (N_6688,N_6376,N_6422);
and U6689 (N_6689,N_6307,N_6402);
nand U6690 (N_6690,N_6469,N_6424);
nor U6691 (N_6691,N_6319,N_6297);
and U6692 (N_6692,N_6329,N_6498);
nand U6693 (N_6693,N_6432,N_6410);
and U6694 (N_6694,N_6345,N_6327);
and U6695 (N_6695,N_6302,N_6288);
nor U6696 (N_6696,N_6362,N_6489);
nand U6697 (N_6697,N_6409,N_6391);
or U6698 (N_6698,N_6256,N_6351);
and U6699 (N_6699,N_6350,N_6444);
nor U6700 (N_6700,N_6276,N_6422);
and U6701 (N_6701,N_6351,N_6343);
nor U6702 (N_6702,N_6402,N_6277);
nor U6703 (N_6703,N_6255,N_6345);
or U6704 (N_6704,N_6464,N_6338);
or U6705 (N_6705,N_6250,N_6408);
nand U6706 (N_6706,N_6285,N_6468);
xnor U6707 (N_6707,N_6361,N_6320);
nand U6708 (N_6708,N_6406,N_6415);
nor U6709 (N_6709,N_6355,N_6332);
and U6710 (N_6710,N_6364,N_6360);
nand U6711 (N_6711,N_6391,N_6392);
nand U6712 (N_6712,N_6323,N_6260);
xor U6713 (N_6713,N_6491,N_6485);
nand U6714 (N_6714,N_6359,N_6351);
xor U6715 (N_6715,N_6473,N_6255);
or U6716 (N_6716,N_6257,N_6397);
or U6717 (N_6717,N_6429,N_6296);
and U6718 (N_6718,N_6479,N_6324);
nor U6719 (N_6719,N_6315,N_6327);
nor U6720 (N_6720,N_6458,N_6417);
nand U6721 (N_6721,N_6291,N_6321);
and U6722 (N_6722,N_6430,N_6283);
nor U6723 (N_6723,N_6405,N_6466);
or U6724 (N_6724,N_6437,N_6256);
nor U6725 (N_6725,N_6344,N_6274);
nand U6726 (N_6726,N_6419,N_6484);
xnor U6727 (N_6727,N_6328,N_6295);
and U6728 (N_6728,N_6451,N_6392);
and U6729 (N_6729,N_6316,N_6335);
xor U6730 (N_6730,N_6277,N_6437);
and U6731 (N_6731,N_6278,N_6496);
nor U6732 (N_6732,N_6253,N_6372);
xnor U6733 (N_6733,N_6337,N_6320);
or U6734 (N_6734,N_6282,N_6423);
xor U6735 (N_6735,N_6363,N_6379);
or U6736 (N_6736,N_6454,N_6296);
and U6737 (N_6737,N_6264,N_6346);
xnor U6738 (N_6738,N_6377,N_6347);
and U6739 (N_6739,N_6468,N_6495);
and U6740 (N_6740,N_6312,N_6414);
or U6741 (N_6741,N_6387,N_6401);
nor U6742 (N_6742,N_6368,N_6358);
nand U6743 (N_6743,N_6365,N_6411);
and U6744 (N_6744,N_6487,N_6347);
nand U6745 (N_6745,N_6421,N_6304);
nor U6746 (N_6746,N_6443,N_6453);
or U6747 (N_6747,N_6311,N_6495);
nor U6748 (N_6748,N_6412,N_6480);
and U6749 (N_6749,N_6314,N_6350);
or U6750 (N_6750,N_6743,N_6650);
and U6751 (N_6751,N_6604,N_6656);
or U6752 (N_6752,N_6553,N_6523);
or U6753 (N_6753,N_6564,N_6692);
nand U6754 (N_6754,N_6521,N_6735);
and U6755 (N_6755,N_6681,N_6688);
and U6756 (N_6756,N_6653,N_6651);
nand U6757 (N_6757,N_6715,N_6520);
nor U6758 (N_6758,N_6675,N_6578);
nor U6759 (N_6759,N_6720,N_6600);
nor U6760 (N_6760,N_6663,N_6555);
xor U6761 (N_6761,N_6562,N_6558);
nor U6762 (N_6762,N_6654,N_6561);
nand U6763 (N_6763,N_6580,N_6566);
nand U6764 (N_6764,N_6565,N_6577);
and U6765 (N_6765,N_6573,N_6507);
xnor U6766 (N_6766,N_6538,N_6599);
xnor U6767 (N_6767,N_6716,N_6543);
nor U6768 (N_6768,N_6524,N_6547);
or U6769 (N_6769,N_6655,N_6643);
or U6770 (N_6770,N_6700,N_6560);
nor U6771 (N_6771,N_6619,N_6626);
or U6772 (N_6772,N_6544,N_6514);
and U6773 (N_6773,N_6625,N_6585);
and U6774 (N_6774,N_6698,N_6724);
nor U6775 (N_6775,N_6574,N_6645);
nor U6776 (N_6776,N_6690,N_6549);
nand U6777 (N_6777,N_6639,N_6737);
nor U6778 (N_6778,N_6537,N_6517);
or U6779 (N_6779,N_6701,N_6622);
and U6780 (N_6780,N_6640,N_6616);
xor U6781 (N_6781,N_6664,N_6508);
xnor U6782 (N_6782,N_6532,N_6670);
xor U6783 (N_6783,N_6552,N_6713);
and U6784 (N_6784,N_6586,N_6527);
nor U6785 (N_6785,N_6595,N_6530);
nor U6786 (N_6786,N_6501,N_6614);
and U6787 (N_6787,N_6541,N_6687);
and U6788 (N_6788,N_6605,N_6534);
and U6789 (N_6789,N_6519,N_6718);
nor U6790 (N_6790,N_6590,N_6647);
nor U6791 (N_6791,N_6696,N_6551);
nor U6792 (N_6792,N_6732,N_6691);
or U6793 (N_6793,N_6730,N_6668);
xnor U6794 (N_6794,N_6748,N_6711);
xor U6795 (N_6795,N_6621,N_6588);
and U6796 (N_6796,N_6575,N_6593);
xor U6797 (N_6797,N_6697,N_6745);
nor U6798 (N_6798,N_6630,N_6506);
nor U6799 (N_6799,N_6661,N_6749);
or U6800 (N_6800,N_6546,N_6740);
nand U6801 (N_6801,N_6576,N_6615);
or U6802 (N_6802,N_6603,N_6602);
or U6803 (N_6803,N_6704,N_6550);
or U6804 (N_6804,N_6567,N_6502);
nor U6805 (N_6805,N_6601,N_6512);
or U6806 (N_6806,N_6708,N_6522);
and U6807 (N_6807,N_6515,N_6738);
or U6808 (N_6808,N_6559,N_6548);
xor U6809 (N_6809,N_6570,N_6678);
or U6810 (N_6810,N_6556,N_6633);
xnor U6811 (N_6811,N_6611,N_6667);
or U6812 (N_6812,N_6648,N_6686);
xnor U6813 (N_6813,N_6657,N_6557);
nand U6814 (N_6814,N_6587,N_6511);
nor U6815 (N_6815,N_6710,N_6747);
nand U6816 (N_6816,N_6609,N_6563);
and U6817 (N_6817,N_6741,N_6510);
and U6818 (N_6818,N_6644,N_6535);
nand U6819 (N_6819,N_6624,N_6528);
or U6820 (N_6820,N_6693,N_6500);
nand U6821 (N_6821,N_6516,N_6568);
nor U6822 (N_6822,N_6707,N_6594);
xor U6823 (N_6823,N_6513,N_6642);
or U6824 (N_6824,N_6682,N_6666);
nor U6825 (N_6825,N_6649,N_6637);
and U6826 (N_6826,N_6542,N_6714);
nand U6827 (N_6827,N_6676,N_6623);
nor U6828 (N_6828,N_6723,N_6536);
nor U6829 (N_6829,N_6736,N_6539);
or U6830 (N_6830,N_6597,N_6646);
nor U6831 (N_6831,N_6733,N_6662);
or U6832 (N_6832,N_6636,N_6734);
nor U6833 (N_6833,N_6652,N_6695);
xor U6834 (N_6834,N_6717,N_6504);
and U6835 (N_6835,N_6607,N_6703);
nand U6836 (N_6836,N_6509,N_6583);
nand U6837 (N_6837,N_6631,N_6683);
xnor U6838 (N_6838,N_6658,N_6627);
and U6839 (N_6839,N_6727,N_6659);
xnor U6840 (N_6840,N_6660,N_6591);
or U6841 (N_6841,N_6746,N_6629);
and U6842 (N_6842,N_6742,N_6608);
nand U6843 (N_6843,N_6729,N_6617);
nor U6844 (N_6844,N_6632,N_6684);
or U6845 (N_6845,N_6721,N_6634);
nand U6846 (N_6846,N_6505,N_6592);
or U6847 (N_6847,N_6589,N_6672);
nand U6848 (N_6848,N_6545,N_6702);
and U6849 (N_6849,N_6598,N_6613);
and U6850 (N_6850,N_6726,N_6706);
nor U6851 (N_6851,N_6739,N_6525);
xnor U6852 (N_6852,N_6610,N_6638);
nor U6853 (N_6853,N_6744,N_6680);
nand U6854 (N_6854,N_6584,N_6606);
and U6855 (N_6855,N_6719,N_6709);
and U6856 (N_6856,N_6531,N_6673);
xnor U6857 (N_6857,N_6679,N_6677);
nand U6858 (N_6858,N_6582,N_6699);
xor U6859 (N_6859,N_6529,N_6596);
or U6860 (N_6860,N_6620,N_6671);
and U6861 (N_6861,N_6669,N_6554);
xnor U6862 (N_6862,N_6685,N_6518);
or U6863 (N_6863,N_6728,N_6712);
nor U6864 (N_6864,N_6540,N_6725);
xnor U6865 (N_6865,N_6581,N_6503);
nand U6866 (N_6866,N_6612,N_6731);
or U6867 (N_6867,N_6569,N_6571);
nor U6868 (N_6868,N_6689,N_6694);
and U6869 (N_6869,N_6635,N_6628);
xnor U6870 (N_6870,N_6579,N_6533);
or U6871 (N_6871,N_6665,N_6705);
xnor U6872 (N_6872,N_6674,N_6641);
nand U6873 (N_6873,N_6722,N_6572);
xnor U6874 (N_6874,N_6526,N_6618);
and U6875 (N_6875,N_6718,N_6683);
nor U6876 (N_6876,N_6627,N_6639);
nand U6877 (N_6877,N_6643,N_6571);
and U6878 (N_6878,N_6608,N_6720);
or U6879 (N_6879,N_6548,N_6679);
nand U6880 (N_6880,N_6670,N_6604);
nand U6881 (N_6881,N_6748,N_6670);
xor U6882 (N_6882,N_6632,N_6639);
and U6883 (N_6883,N_6533,N_6723);
and U6884 (N_6884,N_6616,N_6570);
or U6885 (N_6885,N_6642,N_6675);
and U6886 (N_6886,N_6618,N_6510);
or U6887 (N_6887,N_6532,N_6525);
xnor U6888 (N_6888,N_6739,N_6634);
and U6889 (N_6889,N_6632,N_6571);
nor U6890 (N_6890,N_6556,N_6717);
nand U6891 (N_6891,N_6564,N_6630);
xor U6892 (N_6892,N_6638,N_6554);
xnor U6893 (N_6893,N_6547,N_6726);
or U6894 (N_6894,N_6567,N_6731);
nand U6895 (N_6895,N_6665,N_6728);
nor U6896 (N_6896,N_6541,N_6682);
or U6897 (N_6897,N_6510,N_6517);
xor U6898 (N_6898,N_6705,N_6666);
nand U6899 (N_6899,N_6712,N_6575);
xnor U6900 (N_6900,N_6611,N_6737);
or U6901 (N_6901,N_6693,N_6700);
and U6902 (N_6902,N_6726,N_6743);
xor U6903 (N_6903,N_6744,N_6720);
and U6904 (N_6904,N_6587,N_6654);
or U6905 (N_6905,N_6603,N_6500);
nand U6906 (N_6906,N_6685,N_6571);
and U6907 (N_6907,N_6608,N_6638);
and U6908 (N_6908,N_6611,N_6534);
and U6909 (N_6909,N_6574,N_6604);
and U6910 (N_6910,N_6728,N_6614);
nand U6911 (N_6911,N_6610,N_6534);
nand U6912 (N_6912,N_6571,N_6512);
or U6913 (N_6913,N_6627,N_6538);
nand U6914 (N_6914,N_6742,N_6610);
and U6915 (N_6915,N_6573,N_6506);
or U6916 (N_6916,N_6673,N_6503);
and U6917 (N_6917,N_6664,N_6554);
nor U6918 (N_6918,N_6593,N_6745);
nor U6919 (N_6919,N_6680,N_6690);
and U6920 (N_6920,N_6508,N_6643);
nor U6921 (N_6921,N_6736,N_6537);
nand U6922 (N_6922,N_6637,N_6559);
or U6923 (N_6923,N_6546,N_6682);
nor U6924 (N_6924,N_6519,N_6625);
or U6925 (N_6925,N_6618,N_6550);
and U6926 (N_6926,N_6501,N_6696);
xnor U6927 (N_6927,N_6711,N_6610);
nand U6928 (N_6928,N_6624,N_6610);
nor U6929 (N_6929,N_6592,N_6663);
or U6930 (N_6930,N_6724,N_6579);
nor U6931 (N_6931,N_6670,N_6546);
nor U6932 (N_6932,N_6645,N_6594);
and U6933 (N_6933,N_6547,N_6652);
nor U6934 (N_6934,N_6580,N_6747);
nor U6935 (N_6935,N_6581,N_6649);
nor U6936 (N_6936,N_6648,N_6619);
or U6937 (N_6937,N_6549,N_6687);
nand U6938 (N_6938,N_6730,N_6673);
nand U6939 (N_6939,N_6660,N_6686);
nand U6940 (N_6940,N_6609,N_6589);
xor U6941 (N_6941,N_6648,N_6546);
or U6942 (N_6942,N_6612,N_6645);
nand U6943 (N_6943,N_6663,N_6607);
xnor U6944 (N_6944,N_6705,N_6544);
nand U6945 (N_6945,N_6647,N_6705);
or U6946 (N_6946,N_6577,N_6666);
xnor U6947 (N_6947,N_6724,N_6522);
and U6948 (N_6948,N_6500,N_6596);
nand U6949 (N_6949,N_6586,N_6560);
and U6950 (N_6950,N_6503,N_6660);
nand U6951 (N_6951,N_6749,N_6718);
nor U6952 (N_6952,N_6597,N_6620);
nand U6953 (N_6953,N_6583,N_6603);
and U6954 (N_6954,N_6552,N_6638);
or U6955 (N_6955,N_6573,N_6620);
and U6956 (N_6956,N_6678,N_6598);
nor U6957 (N_6957,N_6512,N_6645);
and U6958 (N_6958,N_6548,N_6681);
and U6959 (N_6959,N_6663,N_6614);
xnor U6960 (N_6960,N_6653,N_6709);
nor U6961 (N_6961,N_6567,N_6662);
or U6962 (N_6962,N_6712,N_6540);
xor U6963 (N_6963,N_6669,N_6676);
xnor U6964 (N_6964,N_6654,N_6541);
or U6965 (N_6965,N_6657,N_6658);
nor U6966 (N_6966,N_6508,N_6667);
and U6967 (N_6967,N_6533,N_6574);
nor U6968 (N_6968,N_6748,N_6659);
xor U6969 (N_6969,N_6631,N_6701);
and U6970 (N_6970,N_6534,N_6616);
xor U6971 (N_6971,N_6728,N_6658);
and U6972 (N_6972,N_6663,N_6669);
nand U6973 (N_6973,N_6549,N_6558);
xnor U6974 (N_6974,N_6562,N_6584);
nand U6975 (N_6975,N_6682,N_6519);
nand U6976 (N_6976,N_6600,N_6646);
xnor U6977 (N_6977,N_6627,N_6501);
nor U6978 (N_6978,N_6705,N_6584);
nand U6979 (N_6979,N_6703,N_6611);
or U6980 (N_6980,N_6521,N_6586);
nand U6981 (N_6981,N_6637,N_6718);
nand U6982 (N_6982,N_6529,N_6650);
nand U6983 (N_6983,N_6655,N_6504);
nor U6984 (N_6984,N_6719,N_6693);
nor U6985 (N_6985,N_6550,N_6588);
or U6986 (N_6986,N_6722,N_6711);
nand U6987 (N_6987,N_6554,N_6534);
and U6988 (N_6988,N_6545,N_6510);
xnor U6989 (N_6989,N_6745,N_6728);
or U6990 (N_6990,N_6724,N_6508);
nor U6991 (N_6991,N_6546,N_6525);
xnor U6992 (N_6992,N_6730,N_6691);
xor U6993 (N_6993,N_6714,N_6550);
nor U6994 (N_6994,N_6519,N_6644);
nor U6995 (N_6995,N_6617,N_6568);
xor U6996 (N_6996,N_6628,N_6551);
nor U6997 (N_6997,N_6640,N_6712);
nor U6998 (N_6998,N_6602,N_6741);
or U6999 (N_6999,N_6546,N_6703);
and U7000 (N_7000,N_6893,N_6955);
and U7001 (N_7001,N_6815,N_6833);
and U7002 (N_7002,N_6896,N_6932);
and U7003 (N_7003,N_6827,N_6768);
xnor U7004 (N_7004,N_6914,N_6843);
and U7005 (N_7005,N_6890,N_6952);
nor U7006 (N_7006,N_6977,N_6899);
nor U7007 (N_7007,N_6796,N_6813);
nand U7008 (N_7008,N_6921,N_6946);
and U7009 (N_7009,N_6781,N_6930);
nand U7010 (N_7010,N_6941,N_6821);
xor U7011 (N_7011,N_6872,N_6972);
nand U7012 (N_7012,N_6857,N_6774);
or U7013 (N_7013,N_6826,N_6775);
nand U7014 (N_7014,N_6840,N_6881);
nand U7015 (N_7015,N_6883,N_6858);
and U7016 (N_7016,N_6853,N_6866);
xor U7017 (N_7017,N_6789,N_6897);
xnor U7018 (N_7018,N_6904,N_6888);
and U7019 (N_7019,N_6874,N_6828);
xor U7020 (N_7020,N_6860,N_6803);
and U7021 (N_7021,N_6825,N_6939);
nor U7022 (N_7022,N_6980,N_6978);
nor U7023 (N_7023,N_6776,N_6937);
xor U7024 (N_7024,N_6832,N_6812);
or U7025 (N_7025,N_6792,N_6993);
or U7026 (N_7026,N_6918,N_6863);
nor U7027 (N_7027,N_6779,N_6973);
or U7028 (N_7028,N_6871,N_6983);
or U7029 (N_7029,N_6911,N_6766);
or U7030 (N_7030,N_6991,N_6926);
or U7031 (N_7031,N_6880,N_6755);
or U7032 (N_7032,N_6777,N_6814);
nor U7033 (N_7033,N_6969,N_6761);
and U7034 (N_7034,N_6886,N_6961);
nand U7035 (N_7035,N_6954,N_6922);
nand U7036 (N_7036,N_6903,N_6979);
or U7037 (N_7037,N_6901,N_6956);
xor U7038 (N_7038,N_6802,N_6895);
nor U7039 (N_7039,N_6758,N_6849);
and U7040 (N_7040,N_6910,N_6982);
nand U7041 (N_7041,N_6794,N_6999);
nand U7042 (N_7042,N_6785,N_6820);
xor U7043 (N_7043,N_6970,N_6879);
or U7044 (N_7044,N_6935,N_6800);
nand U7045 (N_7045,N_6929,N_6753);
xnor U7046 (N_7046,N_6848,N_6798);
nand U7047 (N_7047,N_6942,N_6861);
nand U7048 (N_7048,N_6975,N_6882);
and U7049 (N_7049,N_6894,N_6839);
or U7050 (N_7050,N_6958,N_6898);
and U7051 (N_7051,N_6998,N_6878);
or U7052 (N_7052,N_6810,N_6841);
and U7053 (N_7053,N_6784,N_6864);
nand U7054 (N_7054,N_6960,N_6806);
xnor U7055 (N_7055,N_6995,N_6778);
or U7056 (N_7056,N_6846,N_6764);
or U7057 (N_7057,N_6965,N_6771);
nand U7058 (N_7058,N_6943,N_6763);
and U7059 (N_7059,N_6997,N_6804);
and U7060 (N_7060,N_6767,N_6854);
nor U7061 (N_7061,N_6819,N_6950);
or U7062 (N_7062,N_6752,N_6862);
nor U7063 (N_7063,N_6962,N_6967);
nor U7064 (N_7064,N_6887,N_6934);
and U7065 (N_7065,N_6769,N_6809);
or U7066 (N_7066,N_6944,N_6948);
and U7067 (N_7067,N_6971,N_6940);
and U7068 (N_7068,N_6852,N_6867);
nand U7069 (N_7069,N_6805,N_6987);
and U7070 (N_7070,N_6836,N_6902);
xor U7071 (N_7071,N_6829,N_6868);
nand U7072 (N_7072,N_6762,N_6889);
or U7073 (N_7073,N_6927,N_6985);
xnor U7074 (N_7074,N_6968,N_6884);
nand U7075 (N_7075,N_6877,N_6856);
xnor U7076 (N_7076,N_6850,N_6772);
or U7077 (N_7077,N_6936,N_6757);
nor U7078 (N_7078,N_6783,N_6759);
and U7079 (N_7079,N_6928,N_6844);
and U7080 (N_7080,N_6760,N_6851);
or U7081 (N_7081,N_6966,N_6823);
xor U7082 (N_7082,N_6824,N_6876);
nor U7083 (N_7083,N_6947,N_6992);
or U7084 (N_7084,N_6873,N_6920);
nor U7085 (N_7085,N_6988,N_6986);
nand U7086 (N_7086,N_6831,N_6945);
and U7087 (N_7087,N_6923,N_6782);
nand U7088 (N_7088,N_6917,N_6859);
and U7089 (N_7089,N_6924,N_6816);
nand U7090 (N_7090,N_6976,N_6787);
or U7091 (N_7091,N_6799,N_6913);
xnor U7092 (N_7092,N_6773,N_6830);
xnor U7093 (N_7093,N_6765,N_6750);
and U7094 (N_7094,N_6959,N_6907);
xor U7095 (N_7095,N_6891,N_6984);
xnor U7096 (N_7096,N_6909,N_6786);
nand U7097 (N_7097,N_6885,N_6869);
and U7098 (N_7098,N_6870,N_6808);
and U7099 (N_7099,N_6811,N_6837);
and U7100 (N_7100,N_6905,N_6791);
nor U7101 (N_7101,N_6925,N_6835);
or U7102 (N_7102,N_6933,N_6912);
or U7103 (N_7103,N_6754,N_6915);
nor U7104 (N_7104,N_6989,N_6949);
nor U7105 (N_7105,N_6953,N_6801);
xnor U7106 (N_7106,N_6916,N_6990);
nor U7107 (N_7107,N_6892,N_6807);
or U7108 (N_7108,N_6818,N_6900);
xor U7109 (N_7109,N_6790,N_6756);
and U7110 (N_7110,N_6865,N_6788);
and U7111 (N_7111,N_6780,N_6906);
or U7112 (N_7112,N_6981,N_6797);
nand U7113 (N_7113,N_6855,N_6875);
and U7114 (N_7114,N_6957,N_6751);
and U7115 (N_7115,N_6931,N_6974);
or U7116 (N_7116,N_6919,N_6963);
or U7117 (N_7117,N_6938,N_6996);
nor U7118 (N_7118,N_6795,N_6770);
nor U7119 (N_7119,N_6964,N_6845);
xnor U7120 (N_7120,N_6834,N_6908);
and U7121 (N_7121,N_6842,N_6822);
nand U7122 (N_7122,N_6951,N_6994);
xor U7123 (N_7123,N_6838,N_6847);
xor U7124 (N_7124,N_6793,N_6817);
xnor U7125 (N_7125,N_6895,N_6758);
nand U7126 (N_7126,N_6892,N_6757);
nor U7127 (N_7127,N_6813,N_6970);
or U7128 (N_7128,N_6982,N_6815);
and U7129 (N_7129,N_6946,N_6897);
xnor U7130 (N_7130,N_6861,N_6836);
nand U7131 (N_7131,N_6890,N_6980);
and U7132 (N_7132,N_6964,N_6884);
nand U7133 (N_7133,N_6998,N_6907);
xnor U7134 (N_7134,N_6826,N_6825);
or U7135 (N_7135,N_6917,N_6933);
and U7136 (N_7136,N_6803,N_6811);
xnor U7137 (N_7137,N_6751,N_6852);
or U7138 (N_7138,N_6981,N_6922);
nand U7139 (N_7139,N_6882,N_6750);
nor U7140 (N_7140,N_6840,N_6997);
xor U7141 (N_7141,N_6971,N_6877);
nand U7142 (N_7142,N_6796,N_6844);
or U7143 (N_7143,N_6796,N_6945);
nor U7144 (N_7144,N_6840,N_6896);
and U7145 (N_7145,N_6805,N_6990);
nor U7146 (N_7146,N_6886,N_6967);
and U7147 (N_7147,N_6923,N_6914);
xor U7148 (N_7148,N_6876,N_6899);
and U7149 (N_7149,N_6968,N_6932);
nor U7150 (N_7150,N_6927,N_6764);
nor U7151 (N_7151,N_6816,N_6771);
xnor U7152 (N_7152,N_6912,N_6790);
and U7153 (N_7153,N_6801,N_6815);
and U7154 (N_7154,N_6998,N_6808);
nand U7155 (N_7155,N_6832,N_6926);
and U7156 (N_7156,N_6963,N_6841);
or U7157 (N_7157,N_6877,N_6916);
and U7158 (N_7158,N_6887,N_6971);
nor U7159 (N_7159,N_6860,N_6834);
nor U7160 (N_7160,N_6812,N_6986);
nand U7161 (N_7161,N_6865,N_6849);
nor U7162 (N_7162,N_6989,N_6871);
or U7163 (N_7163,N_6993,N_6832);
nand U7164 (N_7164,N_6890,N_6985);
or U7165 (N_7165,N_6900,N_6843);
and U7166 (N_7166,N_6996,N_6769);
nor U7167 (N_7167,N_6861,N_6853);
nand U7168 (N_7168,N_6799,N_6948);
xnor U7169 (N_7169,N_6818,N_6926);
and U7170 (N_7170,N_6860,N_6778);
nor U7171 (N_7171,N_6834,N_6873);
or U7172 (N_7172,N_6774,N_6869);
xnor U7173 (N_7173,N_6898,N_6789);
and U7174 (N_7174,N_6965,N_6849);
nand U7175 (N_7175,N_6885,N_6969);
xor U7176 (N_7176,N_6791,N_6887);
nor U7177 (N_7177,N_6924,N_6913);
nor U7178 (N_7178,N_6849,N_6810);
or U7179 (N_7179,N_6820,N_6841);
nand U7180 (N_7180,N_6834,N_6800);
nand U7181 (N_7181,N_6973,N_6975);
nand U7182 (N_7182,N_6952,N_6878);
xnor U7183 (N_7183,N_6938,N_6962);
xor U7184 (N_7184,N_6782,N_6769);
nand U7185 (N_7185,N_6837,N_6918);
or U7186 (N_7186,N_6878,N_6949);
nor U7187 (N_7187,N_6885,N_6829);
or U7188 (N_7188,N_6755,N_6795);
nor U7189 (N_7189,N_6765,N_6887);
nor U7190 (N_7190,N_6968,N_6791);
xnor U7191 (N_7191,N_6803,N_6806);
nor U7192 (N_7192,N_6938,N_6824);
xnor U7193 (N_7193,N_6782,N_6862);
nand U7194 (N_7194,N_6951,N_6913);
nand U7195 (N_7195,N_6957,N_6845);
and U7196 (N_7196,N_6869,N_6758);
nand U7197 (N_7197,N_6972,N_6864);
or U7198 (N_7198,N_6881,N_6961);
nand U7199 (N_7199,N_6771,N_6906);
or U7200 (N_7200,N_6863,N_6979);
nor U7201 (N_7201,N_6969,N_6864);
nor U7202 (N_7202,N_6847,N_6855);
xnor U7203 (N_7203,N_6772,N_6880);
xor U7204 (N_7204,N_6864,N_6971);
xnor U7205 (N_7205,N_6758,N_6936);
and U7206 (N_7206,N_6883,N_6895);
xor U7207 (N_7207,N_6769,N_6828);
or U7208 (N_7208,N_6927,N_6897);
or U7209 (N_7209,N_6866,N_6768);
nor U7210 (N_7210,N_6947,N_6896);
xnor U7211 (N_7211,N_6780,N_6977);
xnor U7212 (N_7212,N_6969,N_6862);
or U7213 (N_7213,N_6770,N_6815);
and U7214 (N_7214,N_6999,N_6847);
and U7215 (N_7215,N_6836,N_6888);
or U7216 (N_7216,N_6782,N_6978);
and U7217 (N_7217,N_6959,N_6810);
nor U7218 (N_7218,N_6915,N_6833);
nor U7219 (N_7219,N_6909,N_6953);
xnor U7220 (N_7220,N_6858,N_6800);
nor U7221 (N_7221,N_6859,N_6946);
xnor U7222 (N_7222,N_6844,N_6799);
xnor U7223 (N_7223,N_6858,N_6855);
nand U7224 (N_7224,N_6850,N_6949);
or U7225 (N_7225,N_6858,N_6981);
nand U7226 (N_7226,N_6999,N_6996);
xor U7227 (N_7227,N_6898,N_6972);
xor U7228 (N_7228,N_6952,N_6880);
nor U7229 (N_7229,N_6966,N_6916);
and U7230 (N_7230,N_6761,N_6867);
or U7231 (N_7231,N_6794,N_6875);
xor U7232 (N_7232,N_6823,N_6926);
xor U7233 (N_7233,N_6976,N_6981);
or U7234 (N_7234,N_6995,N_6969);
and U7235 (N_7235,N_6996,N_6908);
xnor U7236 (N_7236,N_6986,N_6755);
nand U7237 (N_7237,N_6872,N_6958);
nand U7238 (N_7238,N_6969,N_6954);
and U7239 (N_7239,N_6932,N_6906);
xnor U7240 (N_7240,N_6832,N_6984);
xnor U7241 (N_7241,N_6813,N_6850);
and U7242 (N_7242,N_6981,N_6819);
or U7243 (N_7243,N_6992,N_6978);
and U7244 (N_7244,N_6824,N_6949);
nor U7245 (N_7245,N_6887,N_6824);
and U7246 (N_7246,N_6893,N_6907);
and U7247 (N_7247,N_6907,N_6857);
xor U7248 (N_7248,N_6929,N_6969);
nand U7249 (N_7249,N_6964,N_6818);
or U7250 (N_7250,N_7120,N_7003);
nand U7251 (N_7251,N_7195,N_7012);
and U7252 (N_7252,N_7167,N_7171);
nand U7253 (N_7253,N_7114,N_7149);
xor U7254 (N_7254,N_7088,N_7204);
nand U7255 (N_7255,N_7113,N_7227);
or U7256 (N_7256,N_7109,N_7168);
nor U7257 (N_7257,N_7131,N_7047);
nor U7258 (N_7258,N_7121,N_7176);
nor U7259 (N_7259,N_7089,N_7102);
nor U7260 (N_7260,N_7134,N_7217);
and U7261 (N_7261,N_7203,N_7162);
xor U7262 (N_7262,N_7188,N_7105);
and U7263 (N_7263,N_7097,N_7142);
nand U7264 (N_7264,N_7035,N_7191);
xnor U7265 (N_7265,N_7236,N_7146);
nor U7266 (N_7266,N_7010,N_7023);
and U7267 (N_7267,N_7243,N_7199);
nor U7268 (N_7268,N_7068,N_7186);
and U7269 (N_7269,N_7185,N_7228);
or U7270 (N_7270,N_7233,N_7237);
nand U7271 (N_7271,N_7169,N_7209);
xnor U7272 (N_7272,N_7156,N_7071);
and U7273 (N_7273,N_7028,N_7235);
nor U7274 (N_7274,N_7231,N_7226);
nor U7275 (N_7275,N_7210,N_7218);
xor U7276 (N_7276,N_7104,N_7213);
or U7277 (N_7277,N_7110,N_7182);
nor U7278 (N_7278,N_7249,N_7192);
xor U7279 (N_7279,N_7174,N_7133);
and U7280 (N_7280,N_7147,N_7202);
and U7281 (N_7281,N_7177,N_7242);
or U7282 (N_7282,N_7041,N_7016);
nand U7283 (N_7283,N_7013,N_7076);
or U7284 (N_7284,N_7241,N_7222);
xor U7285 (N_7285,N_7056,N_7000);
and U7286 (N_7286,N_7164,N_7207);
xor U7287 (N_7287,N_7208,N_7136);
and U7288 (N_7288,N_7206,N_7018);
xnor U7289 (N_7289,N_7048,N_7247);
nand U7290 (N_7290,N_7065,N_7022);
xor U7291 (N_7291,N_7248,N_7154);
xor U7292 (N_7292,N_7062,N_7161);
nand U7293 (N_7293,N_7194,N_7224);
and U7294 (N_7294,N_7152,N_7115);
or U7295 (N_7295,N_7141,N_7096);
nand U7296 (N_7296,N_7126,N_7198);
nor U7297 (N_7297,N_7106,N_7074);
xnor U7298 (N_7298,N_7029,N_7019);
xor U7299 (N_7299,N_7044,N_7196);
or U7300 (N_7300,N_7066,N_7042);
and U7301 (N_7301,N_7092,N_7001);
xor U7302 (N_7302,N_7173,N_7059);
or U7303 (N_7303,N_7043,N_7132);
nor U7304 (N_7304,N_7008,N_7170);
nor U7305 (N_7305,N_7049,N_7038);
or U7306 (N_7306,N_7122,N_7183);
or U7307 (N_7307,N_7034,N_7025);
or U7308 (N_7308,N_7117,N_7094);
nor U7309 (N_7309,N_7212,N_7024);
nand U7310 (N_7310,N_7091,N_7151);
nor U7311 (N_7311,N_7127,N_7053);
nor U7312 (N_7312,N_7211,N_7014);
nand U7313 (N_7313,N_7178,N_7221);
xnor U7314 (N_7314,N_7219,N_7137);
xor U7315 (N_7315,N_7020,N_7086);
nor U7316 (N_7316,N_7036,N_7021);
or U7317 (N_7317,N_7103,N_7118);
and U7318 (N_7318,N_7160,N_7125);
nand U7319 (N_7319,N_7073,N_7039);
nor U7320 (N_7320,N_7232,N_7017);
xor U7321 (N_7321,N_7051,N_7225);
nor U7322 (N_7322,N_7244,N_7119);
nor U7323 (N_7323,N_7033,N_7215);
nor U7324 (N_7324,N_7135,N_7081);
and U7325 (N_7325,N_7004,N_7099);
nand U7326 (N_7326,N_7189,N_7032);
or U7327 (N_7327,N_7148,N_7240);
or U7328 (N_7328,N_7128,N_7138);
nor U7329 (N_7329,N_7112,N_7129);
or U7330 (N_7330,N_7002,N_7229);
nor U7331 (N_7331,N_7158,N_7165);
or U7332 (N_7332,N_7027,N_7163);
xor U7333 (N_7333,N_7246,N_7234);
and U7334 (N_7334,N_7045,N_7187);
nand U7335 (N_7335,N_7087,N_7197);
nor U7336 (N_7336,N_7026,N_7058);
nand U7337 (N_7337,N_7159,N_7030);
nor U7338 (N_7338,N_7072,N_7205);
nor U7339 (N_7339,N_7090,N_7201);
nor U7340 (N_7340,N_7172,N_7220);
and U7341 (N_7341,N_7040,N_7124);
xnor U7342 (N_7342,N_7116,N_7067);
nand U7343 (N_7343,N_7075,N_7184);
xnor U7344 (N_7344,N_7052,N_7238);
and U7345 (N_7345,N_7085,N_7175);
nor U7346 (N_7346,N_7093,N_7084);
xnor U7347 (N_7347,N_7007,N_7111);
xor U7348 (N_7348,N_7123,N_7064);
and U7349 (N_7349,N_7069,N_7079);
nand U7350 (N_7350,N_7130,N_7101);
nor U7351 (N_7351,N_7239,N_7150);
or U7352 (N_7352,N_7006,N_7063);
nor U7353 (N_7353,N_7070,N_7083);
xor U7354 (N_7354,N_7200,N_7179);
nor U7355 (N_7355,N_7078,N_7245);
and U7356 (N_7356,N_7144,N_7193);
or U7357 (N_7357,N_7031,N_7005);
xnor U7358 (N_7358,N_7216,N_7060);
nand U7359 (N_7359,N_7155,N_7057);
or U7360 (N_7360,N_7054,N_7214);
nand U7361 (N_7361,N_7180,N_7046);
nor U7362 (N_7362,N_7015,N_7166);
nor U7363 (N_7363,N_7153,N_7157);
and U7364 (N_7364,N_7011,N_7050);
xor U7365 (N_7365,N_7095,N_7108);
and U7366 (N_7366,N_7037,N_7061);
nor U7367 (N_7367,N_7190,N_7107);
nand U7368 (N_7368,N_7009,N_7143);
or U7369 (N_7369,N_7055,N_7139);
and U7370 (N_7370,N_7181,N_7140);
or U7371 (N_7371,N_7223,N_7080);
or U7372 (N_7372,N_7082,N_7077);
xnor U7373 (N_7373,N_7098,N_7100);
and U7374 (N_7374,N_7145,N_7230);
or U7375 (N_7375,N_7229,N_7090);
nand U7376 (N_7376,N_7006,N_7106);
and U7377 (N_7377,N_7142,N_7047);
and U7378 (N_7378,N_7233,N_7083);
or U7379 (N_7379,N_7163,N_7165);
nand U7380 (N_7380,N_7157,N_7037);
nand U7381 (N_7381,N_7099,N_7102);
nand U7382 (N_7382,N_7105,N_7046);
nand U7383 (N_7383,N_7137,N_7050);
and U7384 (N_7384,N_7113,N_7142);
nor U7385 (N_7385,N_7074,N_7141);
nand U7386 (N_7386,N_7064,N_7072);
or U7387 (N_7387,N_7235,N_7074);
nand U7388 (N_7388,N_7121,N_7157);
nor U7389 (N_7389,N_7044,N_7197);
nor U7390 (N_7390,N_7069,N_7006);
xor U7391 (N_7391,N_7100,N_7153);
nor U7392 (N_7392,N_7062,N_7230);
xor U7393 (N_7393,N_7232,N_7116);
nand U7394 (N_7394,N_7239,N_7166);
or U7395 (N_7395,N_7060,N_7200);
xor U7396 (N_7396,N_7163,N_7048);
or U7397 (N_7397,N_7039,N_7187);
xor U7398 (N_7398,N_7107,N_7062);
nor U7399 (N_7399,N_7188,N_7022);
nor U7400 (N_7400,N_7171,N_7082);
nand U7401 (N_7401,N_7218,N_7083);
xor U7402 (N_7402,N_7173,N_7226);
nor U7403 (N_7403,N_7122,N_7180);
nor U7404 (N_7404,N_7206,N_7032);
or U7405 (N_7405,N_7023,N_7249);
or U7406 (N_7406,N_7147,N_7180);
xnor U7407 (N_7407,N_7079,N_7107);
nor U7408 (N_7408,N_7064,N_7046);
nand U7409 (N_7409,N_7168,N_7033);
nor U7410 (N_7410,N_7167,N_7106);
xor U7411 (N_7411,N_7121,N_7243);
and U7412 (N_7412,N_7146,N_7050);
or U7413 (N_7413,N_7150,N_7024);
nor U7414 (N_7414,N_7011,N_7169);
nand U7415 (N_7415,N_7191,N_7205);
and U7416 (N_7416,N_7017,N_7022);
nand U7417 (N_7417,N_7102,N_7040);
or U7418 (N_7418,N_7176,N_7091);
or U7419 (N_7419,N_7144,N_7048);
xnor U7420 (N_7420,N_7078,N_7159);
xor U7421 (N_7421,N_7150,N_7217);
or U7422 (N_7422,N_7033,N_7055);
or U7423 (N_7423,N_7226,N_7162);
or U7424 (N_7424,N_7079,N_7093);
and U7425 (N_7425,N_7231,N_7056);
and U7426 (N_7426,N_7075,N_7201);
or U7427 (N_7427,N_7015,N_7114);
and U7428 (N_7428,N_7054,N_7224);
and U7429 (N_7429,N_7066,N_7214);
or U7430 (N_7430,N_7107,N_7049);
and U7431 (N_7431,N_7007,N_7173);
or U7432 (N_7432,N_7039,N_7161);
xnor U7433 (N_7433,N_7216,N_7171);
nor U7434 (N_7434,N_7048,N_7149);
xor U7435 (N_7435,N_7226,N_7047);
or U7436 (N_7436,N_7128,N_7220);
nor U7437 (N_7437,N_7199,N_7037);
nor U7438 (N_7438,N_7009,N_7065);
nor U7439 (N_7439,N_7208,N_7168);
nand U7440 (N_7440,N_7156,N_7060);
xor U7441 (N_7441,N_7050,N_7028);
xnor U7442 (N_7442,N_7061,N_7008);
nand U7443 (N_7443,N_7023,N_7118);
nand U7444 (N_7444,N_7114,N_7142);
xor U7445 (N_7445,N_7209,N_7031);
nand U7446 (N_7446,N_7079,N_7131);
nor U7447 (N_7447,N_7087,N_7075);
xor U7448 (N_7448,N_7002,N_7085);
xor U7449 (N_7449,N_7089,N_7227);
nor U7450 (N_7450,N_7158,N_7009);
nand U7451 (N_7451,N_7161,N_7241);
or U7452 (N_7452,N_7044,N_7015);
nor U7453 (N_7453,N_7192,N_7179);
and U7454 (N_7454,N_7171,N_7098);
or U7455 (N_7455,N_7247,N_7243);
xor U7456 (N_7456,N_7113,N_7131);
nor U7457 (N_7457,N_7074,N_7109);
and U7458 (N_7458,N_7215,N_7247);
xnor U7459 (N_7459,N_7230,N_7025);
xnor U7460 (N_7460,N_7186,N_7072);
or U7461 (N_7461,N_7124,N_7160);
xnor U7462 (N_7462,N_7114,N_7009);
and U7463 (N_7463,N_7202,N_7061);
or U7464 (N_7464,N_7216,N_7046);
nor U7465 (N_7465,N_7007,N_7246);
or U7466 (N_7466,N_7228,N_7222);
and U7467 (N_7467,N_7082,N_7048);
nor U7468 (N_7468,N_7189,N_7014);
or U7469 (N_7469,N_7216,N_7049);
or U7470 (N_7470,N_7108,N_7136);
or U7471 (N_7471,N_7016,N_7060);
and U7472 (N_7472,N_7208,N_7246);
nand U7473 (N_7473,N_7034,N_7089);
or U7474 (N_7474,N_7244,N_7205);
nor U7475 (N_7475,N_7062,N_7070);
xor U7476 (N_7476,N_7067,N_7148);
or U7477 (N_7477,N_7132,N_7213);
nand U7478 (N_7478,N_7080,N_7159);
and U7479 (N_7479,N_7236,N_7042);
and U7480 (N_7480,N_7170,N_7199);
or U7481 (N_7481,N_7209,N_7148);
xor U7482 (N_7482,N_7055,N_7164);
nand U7483 (N_7483,N_7193,N_7223);
nand U7484 (N_7484,N_7216,N_7151);
nor U7485 (N_7485,N_7035,N_7115);
xnor U7486 (N_7486,N_7000,N_7196);
nor U7487 (N_7487,N_7081,N_7105);
nor U7488 (N_7488,N_7047,N_7233);
and U7489 (N_7489,N_7233,N_7046);
nor U7490 (N_7490,N_7030,N_7163);
nand U7491 (N_7491,N_7163,N_7162);
nor U7492 (N_7492,N_7119,N_7166);
or U7493 (N_7493,N_7210,N_7224);
and U7494 (N_7494,N_7052,N_7047);
xor U7495 (N_7495,N_7022,N_7068);
nand U7496 (N_7496,N_7017,N_7200);
and U7497 (N_7497,N_7065,N_7115);
xor U7498 (N_7498,N_7036,N_7159);
nor U7499 (N_7499,N_7229,N_7136);
nand U7500 (N_7500,N_7354,N_7464);
or U7501 (N_7501,N_7287,N_7329);
xor U7502 (N_7502,N_7460,N_7258);
nand U7503 (N_7503,N_7421,N_7335);
nor U7504 (N_7504,N_7436,N_7259);
and U7505 (N_7505,N_7345,N_7267);
nor U7506 (N_7506,N_7364,N_7253);
xor U7507 (N_7507,N_7310,N_7461);
or U7508 (N_7508,N_7412,N_7428);
nand U7509 (N_7509,N_7397,N_7476);
xor U7510 (N_7510,N_7268,N_7434);
xnor U7511 (N_7511,N_7305,N_7328);
nor U7512 (N_7512,N_7493,N_7336);
nand U7513 (N_7513,N_7477,N_7290);
xor U7514 (N_7514,N_7313,N_7337);
xor U7515 (N_7515,N_7368,N_7250);
and U7516 (N_7516,N_7377,N_7358);
nand U7517 (N_7517,N_7447,N_7495);
nand U7518 (N_7518,N_7373,N_7296);
or U7519 (N_7519,N_7426,N_7485);
nand U7520 (N_7520,N_7449,N_7366);
xnor U7521 (N_7521,N_7362,N_7286);
and U7522 (N_7522,N_7439,N_7450);
nand U7523 (N_7523,N_7486,N_7312);
and U7524 (N_7524,N_7424,N_7378);
nor U7525 (N_7525,N_7279,N_7403);
xor U7526 (N_7526,N_7320,N_7443);
or U7527 (N_7527,N_7472,N_7479);
or U7528 (N_7528,N_7375,N_7456);
xor U7529 (N_7529,N_7445,N_7322);
and U7530 (N_7530,N_7490,N_7353);
nor U7531 (N_7531,N_7374,N_7355);
and U7532 (N_7532,N_7474,N_7384);
nor U7533 (N_7533,N_7441,N_7416);
nor U7534 (N_7534,N_7261,N_7380);
or U7535 (N_7535,N_7491,N_7357);
nand U7536 (N_7536,N_7467,N_7407);
and U7537 (N_7537,N_7420,N_7369);
nand U7538 (N_7538,N_7297,N_7352);
nor U7539 (N_7539,N_7282,N_7371);
nand U7540 (N_7540,N_7365,N_7321);
nor U7541 (N_7541,N_7307,N_7251);
and U7542 (N_7542,N_7478,N_7489);
nor U7543 (N_7543,N_7392,N_7315);
or U7544 (N_7544,N_7319,N_7399);
xor U7545 (N_7545,N_7482,N_7400);
or U7546 (N_7546,N_7265,N_7385);
nand U7547 (N_7547,N_7370,N_7414);
or U7548 (N_7548,N_7475,N_7404);
nand U7549 (N_7549,N_7338,N_7372);
nor U7550 (N_7550,N_7342,N_7376);
and U7551 (N_7551,N_7300,N_7281);
nand U7552 (N_7552,N_7360,N_7264);
xor U7553 (N_7553,N_7356,N_7272);
and U7554 (N_7554,N_7306,N_7276);
xor U7555 (N_7555,N_7344,N_7395);
and U7556 (N_7556,N_7388,N_7275);
or U7557 (N_7557,N_7273,N_7302);
nand U7558 (N_7558,N_7406,N_7325);
xnor U7559 (N_7559,N_7433,N_7346);
nand U7560 (N_7560,N_7418,N_7323);
nor U7561 (N_7561,N_7367,N_7348);
or U7562 (N_7562,N_7285,N_7314);
and U7563 (N_7563,N_7381,N_7289);
and U7564 (N_7564,N_7317,N_7410);
nand U7565 (N_7565,N_7484,N_7288);
or U7566 (N_7566,N_7442,N_7341);
nor U7567 (N_7567,N_7481,N_7311);
nand U7568 (N_7568,N_7382,N_7316);
nand U7569 (N_7569,N_7429,N_7334);
or U7570 (N_7570,N_7254,N_7387);
nor U7571 (N_7571,N_7270,N_7430);
and U7572 (N_7572,N_7396,N_7301);
or U7573 (N_7573,N_7263,N_7499);
nand U7574 (N_7574,N_7425,N_7440);
or U7575 (N_7575,N_7471,N_7409);
xor U7576 (N_7576,N_7350,N_7269);
xor U7577 (N_7577,N_7389,N_7298);
nor U7578 (N_7578,N_7332,N_7379);
xnor U7579 (N_7579,N_7359,N_7303);
nor U7580 (N_7580,N_7280,N_7257);
nor U7581 (N_7581,N_7393,N_7292);
xnor U7582 (N_7582,N_7262,N_7327);
nor U7583 (N_7583,N_7457,N_7427);
xor U7584 (N_7584,N_7483,N_7488);
nor U7585 (N_7585,N_7340,N_7274);
or U7586 (N_7586,N_7444,N_7331);
and U7587 (N_7587,N_7448,N_7452);
nand U7588 (N_7588,N_7487,N_7480);
xor U7589 (N_7589,N_7349,N_7413);
and U7590 (N_7590,N_7446,N_7496);
nor U7591 (N_7591,N_7309,N_7383);
xor U7592 (N_7592,N_7463,N_7438);
xor U7593 (N_7593,N_7347,N_7293);
nand U7594 (N_7594,N_7492,N_7437);
or U7595 (N_7595,N_7454,N_7401);
nor U7596 (N_7596,N_7498,N_7284);
nor U7597 (N_7597,N_7333,N_7419);
nor U7598 (N_7598,N_7455,N_7256);
nor U7599 (N_7599,N_7304,N_7283);
xnor U7600 (N_7600,N_7260,N_7473);
nand U7601 (N_7601,N_7398,N_7391);
xor U7602 (N_7602,N_7405,N_7266);
xor U7603 (N_7603,N_7255,N_7252);
xnor U7604 (N_7604,N_7423,N_7462);
xnor U7605 (N_7605,N_7469,N_7408);
or U7606 (N_7606,N_7390,N_7470);
and U7607 (N_7607,N_7324,N_7402);
or U7608 (N_7608,N_7326,N_7278);
or U7609 (N_7609,N_7432,N_7330);
and U7610 (N_7610,N_7343,N_7422);
or U7611 (N_7611,N_7466,N_7318);
nor U7612 (N_7612,N_7363,N_7435);
nor U7613 (N_7613,N_7291,N_7295);
nand U7614 (N_7614,N_7468,N_7394);
xor U7615 (N_7615,N_7411,N_7417);
xor U7616 (N_7616,N_7431,N_7277);
xor U7617 (N_7617,N_7415,N_7459);
or U7618 (N_7618,N_7453,N_7308);
and U7619 (N_7619,N_7339,N_7494);
or U7620 (N_7620,N_7458,N_7361);
nand U7621 (N_7621,N_7465,N_7497);
or U7622 (N_7622,N_7299,N_7451);
xor U7623 (N_7623,N_7386,N_7294);
and U7624 (N_7624,N_7351,N_7271);
and U7625 (N_7625,N_7428,N_7345);
nand U7626 (N_7626,N_7486,N_7259);
nor U7627 (N_7627,N_7397,N_7323);
nor U7628 (N_7628,N_7421,N_7466);
xor U7629 (N_7629,N_7272,N_7413);
or U7630 (N_7630,N_7271,N_7496);
nand U7631 (N_7631,N_7415,N_7406);
nor U7632 (N_7632,N_7461,N_7331);
and U7633 (N_7633,N_7474,N_7342);
and U7634 (N_7634,N_7371,N_7307);
or U7635 (N_7635,N_7322,N_7335);
or U7636 (N_7636,N_7285,N_7436);
nor U7637 (N_7637,N_7395,N_7282);
nand U7638 (N_7638,N_7400,N_7468);
and U7639 (N_7639,N_7473,N_7389);
or U7640 (N_7640,N_7418,N_7262);
xnor U7641 (N_7641,N_7307,N_7444);
and U7642 (N_7642,N_7462,N_7402);
xnor U7643 (N_7643,N_7474,N_7335);
xor U7644 (N_7644,N_7487,N_7349);
xor U7645 (N_7645,N_7274,N_7466);
nand U7646 (N_7646,N_7357,N_7309);
or U7647 (N_7647,N_7460,N_7413);
or U7648 (N_7648,N_7476,N_7405);
nand U7649 (N_7649,N_7453,N_7319);
nand U7650 (N_7650,N_7307,N_7431);
xnor U7651 (N_7651,N_7309,N_7294);
xor U7652 (N_7652,N_7283,N_7301);
xnor U7653 (N_7653,N_7346,N_7424);
nand U7654 (N_7654,N_7298,N_7378);
or U7655 (N_7655,N_7467,N_7309);
nor U7656 (N_7656,N_7273,N_7392);
nand U7657 (N_7657,N_7478,N_7281);
nand U7658 (N_7658,N_7346,N_7294);
and U7659 (N_7659,N_7436,N_7497);
xor U7660 (N_7660,N_7346,N_7262);
or U7661 (N_7661,N_7419,N_7261);
xor U7662 (N_7662,N_7472,N_7358);
nand U7663 (N_7663,N_7401,N_7386);
and U7664 (N_7664,N_7268,N_7256);
nor U7665 (N_7665,N_7256,N_7420);
and U7666 (N_7666,N_7469,N_7472);
nand U7667 (N_7667,N_7387,N_7260);
nor U7668 (N_7668,N_7456,N_7404);
and U7669 (N_7669,N_7345,N_7481);
or U7670 (N_7670,N_7330,N_7430);
nand U7671 (N_7671,N_7256,N_7495);
nor U7672 (N_7672,N_7322,N_7462);
or U7673 (N_7673,N_7385,N_7307);
xor U7674 (N_7674,N_7323,N_7419);
nor U7675 (N_7675,N_7402,N_7310);
nand U7676 (N_7676,N_7429,N_7487);
or U7677 (N_7677,N_7480,N_7272);
nor U7678 (N_7678,N_7331,N_7349);
nand U7679 (N_7679,N_7383,N_7482);
and U7680 (N_7680,N_7299,N_7287);
or U7681 (N_7681,N_7457,N_7484);
nand U7682 (N_7682,N_7380,N_7358);
and U7683 (N_7683,N_7419,N_7274);
xnor U7684 (N_7684,N_7448,N_7390);
and U7685 (N_7685,N_7345,N_7477);
xor U7686 (N_7686,N_7268,N_7390);
nor U7687 (N_7687,N_7477,N_7467);
or U7688 (N_7688,N_7378,N_7265);
nand U7689 (N_7689,N_7342,N_7324);
xnor U7690 (N_7690,N_7473,N_7326);
or U7691 (N_7691,N_7468,N_7449);
nand U7692 (N_7692,N_7347,N_7408);
nor U7693 (N_7693,N_7312,N_7365);
nor U7694 (N_7694,N_7342,N_7457);
nand U7695 (N_7695,N_7260,N_7440);
or U7696 (N_7696,N_7342,N_7423);
or U7697 (N_7697,N_7415,N_7326);
nor U7698 (N_7698,N_7270,N_7448);
and U7699 (N_7699,N_7445,N_7257);
and U7700 (N_7700,N_7361,N_7467);
nand U7701 (N_7701,N_7394,N_7494);
nand U7702 (N_7702,N_7345,N_7256);
nand U7703 (N_7703,N_7407,N_7329);
and U7704 (N_7704,N_7368,N_7479);
and U7705 (N_7705,N_7270,N_7352);
nor U7706 (N_7706,N_7447,N_7281);
xnor U7707 (N_7707,N_7451,N_7391);
xnor U7708 (N_7708,N_7474,N_7302);
and U7709 (N_7709,N_7333,N_7388);
or U7710 (N_7710,N_7407,N_7494);
or U7711 (N_7711,N_7405,N_7435);
nand U7712 (N_7712,N_7431,N_7317);
xnor U7713 (N_7713,N_7453,N_7491);
nor U7714 (N_7714,N_7439,N_7469);
and U7715 (N_7715,N_7398,N_7253);
and U7716 (N_7716,N_7334,N_7371);
or U7717 (N_7717,N_7469,N_7272);
or U7718 (N_7718,N_7405,N_7431);
xnor U7719 (N_7719,N_7440,N_7274);
nand U7720 (N_7720,N_7331,N_7441);
and U7721 (N_7721,N_7465,N_7297);
xor U7722 (N_7722,N_7389,N_7406);
or U7723 (N_7723,N_7313,N_7283);
or U7724 (N_7724,N_7316,N_7448);
nor U7725 (N_7725,N_7423,N_7345);
nand U7726 (N_7726,N_7499,N_7456);
or U7727 (N_7727,N_7267,N_7316);
or U7728 (N_7728,N_7305,N_7278);
nand U7729 (N_7729,N_7294,N_7265);
nor U7730 (N_7730,N_7489,N_7300);
and U7731 (N_7731,N_7440,N_7252);
or U7732 (N_7732,N_7325,N_7336);
nand U7733 (N_7733,N_7313,N_7445);
xor U7734 (N_7734,N_7433,N_7403);
nor U7735 (N_7735,N_7293,N_7372);
xnor U7736 (N_7736,N_7363,N_7472);
or U7737 (N_7737,N_7376,N_7418);
and U7738 (N_7738,N_7492,N_7458);
and U7739 (N_7739,N_7302,N_7352);
and U7740 (N_7740,N_7419,N_7301);
or U7741 (N_7741,N_7384,N_7265);
and U7742 (N_7742,N_7327,N_7359);
and U7743 (N_7743,N_7305,N_7452);
nand U7744 (N_7744,N_7358,N_7301);
or U7745 (N_7745,N_7337,N_7341);
nor U7746 (N_7746,N_7410,N_7368);
nand U7747 (N_7747,N_7485,N_7359);
xor U7748 (N_7748,N_7440,N_7262);
nand U7749 (N_7749,N_7406,N_7364);
nor U7750 (N_7750,N_7698,N_7510);
and U7751 (N_7751,N_7745,N_7593);
nor U7752 (N_7752,N_7734,N_7726);
xor U7753 (N_7753,N_7646,N_7507);
nand U7754 (N_7754,N_7628,N_7565);
or U7755 (N_7755,N_7689,N_7679);
xnor U7756 (N_7756,N_7638,N_7722);
or U7757 (N_7757,N_7647,N_7569);
or U7758 (N_7758,N_7559,N_7704);
xor U7759 (N_7759,N_7557,N_7516);
and U7760 (N_7760,N_7623,N_7571);
and U7761 (N_7761,N_7532,N_7552);
nor U7762 (N_7762,N_7687,N_7543);
and U7763 (N_7763,N_7680,N_7743);
and U7764 (N_7764,N_7564,N_7602);
nand U7765 (N_7765,N_7604,N_7728);
nand U7766 (N_7766,N_7735,N_7701);
or U7767 (N_7767,N_7749,N_7560);
nor U7768 (N_7768,N_7664,N_7581);
nand U7769 (N_7769,N_7671,N_7654);
nor U7770 (N_7770,N_7621,N_7586);
or U7771 (N_7771,N_7732,N_7556);
or U7772 (N_7772,N_7537,N_7637);
nand U7773 (N_7773,N_7530,N_7667);
or U7774 (N_7774,N_7607,N_7641);
xnor U7775 (N_7775,N_7632,N_7513);
nand U7776 (N_7776,N_7547,N_7694);
nand U7777 (N_7777,N_7619,N_7518);
or U7778 (N_7778,N_7582,N_7729);
and U7779 (N_7779,N_7611,N_7657);
and U7780 (N_7780,N_7691,N_7742);
xnor U7781 (N_7781,N_7551,N_7539);
xnor U7782 (N_7782,N_7662,N_7723);
nand U7783 (N_7783,N_7568,N_7653);
xor U7784 (N_7784,N_7739,N_7576);
xor U7785 (N_7785,N_7512,N_7548);
and U7786 (N_7786,N_7717,N_7716);
xor U7787 (N_7787,N_7522,N_7620);
xnor U7788 (N_7788,N_7606,N_7640);
nand U7789 (N_7789,N_7612,N_7738);
and U7790 (N_7790,N_7688,N_7655);
or U7791 (N_7791,N_7643,N_7613);
nor U7792 (N_7792,N_7578,N_7589);
nor U7793 (N_7793,N_7700,N_7709);
and U7794 (N_7794,N_7535,N_7703);
xor U7795 (N_7795,N_7696,N_7577);
and U7796 (N_7796,N_7675,N_7523);
nor U7797 (N_7797,N_7563,N_7708);
and U7798 (N_7798,N_7658,N_7651);
xor U7799 (N_7799,N_7545,N_7562);
xor U7800 (N_7800,N_7642,N_7546);
or U7801 (N_7801,N_7713,N_7501);
or U7802 (N_7802,N_7605,N_7618);
or U7803 (N_7803,N_7656,N_7674);
nand U7804 (N_7804,N_7681,N_7707);
or U7805 (N_7805,N_7528,N_7633);
or U7806 (N_7806,N_7711,N_7572);
and U7807 (N_7807,N_7744,N_7574);
or U7808 (N_7808,N_7629,N_7626);
xor U7809 (N_7809,N_7526,N_7685);
nor U7810 (N_7810,N_7660,N_7521);
or U7811 (N_7811,N_7673,N_7590);
and U7812 (N_7812,N_7599,N_7747);
xnor U7813 (N_7813,N_7666,N_7500);
nor U7814 (N_7814,N_7519,N_7668);
xor U7815 (N_7815,N_7587,N_7624);
nand U7816 (N_7816,N_7733,N_7692);
or U7817 (N_7817,N_7695,N_7533);
nand U7818 (N_7818,N_7731,N_7541);
and U7819 (N_7819,N_7514,N_7725);
nor U7820 (N_7820,N_7622,N_7614);
or U7821 (N_7821,N_7697,N_7580);
and U7822 (N_7822,N_7631,N_7588);
or U7823 (N_7823,N_7724,N_7506);
nor U7824 (N_7824,N_7555,N_7683);
and U7825 (N_7825,N_7720,N_7508);
and U7826 (N_7826,N_7567,N_7737);
nand U7827 (N_7827,N_7600,N_7625);
and U7828 (N_7828,N_7542,N_7594);
or U7829 (N_7829,N_7504,N_7736);
or U7830 (N_7830,N_7645,N_7693);
xnor U7831 (N_7831,N_7690,N_7598);
or U7832 (N_7832,N_7635,N_7648);
and U7833 (N_7833,N_7558,N_7509);
xor U7834 (N_7834,N_7634,N_7592);
nor U7835 (N_7835,N_7538,N_7601);
and U7836 (N_7836,N_7554,N_7505);
xor U7837 (N_7837,N_7584,N_7550);
and U7838 (N_7838,N_7677,N_7527);
and U7839 (N_7839,N_7603,N_7610);
or U7840 (N_7840,N_7615,N_7575);
nand U7841 (N_7841,N_7520,N_7570);
nand U7842 (N_7842,N_7748,N_7531);
and U7843 (N_7843,N_7650,N_7746);
nand U7844 (N_7844,N_7596,N_7740);
nor U7845 (N_7845,N_7682,N_7649);
and U7846 (N_7846,N_7665,N_7573);
and U7847 (N_7847,N_7718,N_7608);
xnor U7848 (N_7848,N_7699,N_7644);
and U7849 (N_7849,N_7659,N_7583);
and U7850 (N_7850,N_7670,N_7517);
nor U7851 (N_7851,N_7727,N_7515);
nor U7852 (N_7852,N_7715,N_7585);
xor U7853 (N_7853,N_7661,N_7524);
nand U7854 (N_7854,N_7676,N_7561);
nand U7855 (N_7855,N_7669,N_7553);
nand U7856 (N_7856,N_7705,N_7686);
or U7857 (N_7857,N_7549,N_7540);
and U7858 (N_7858,N_7597,N_7678);
nor U7859 (N_7859,N_7616,N_7702);
xor U7860 (N_7860,N_7714,N_7706);
nor U7861 (N_7861,N_7730,N_7721);
nand U7862 (N_7862,N_7636,N_7536);
and U7863 (N_7863,N_7595,N_7639);
xor U7864 (N_7864,N_7663,N_7503);
nor U7865 (N_7865,N_7511,N_7630);
and U7866 (N_7866,N_7529,N_7544);
xor U7867 (N_7867,N_7712,N_7609);
and U7868 (N_7868,N_7684,N_7525);
or U7869 (N_7869,N_7617,N_7672);
nor U7870 (N_7870,N_7627,N_7652);
and U7871 (N_7871,N_7719,N_7591);
xor U7872 (N_7872,N_7710,N_7741);
and U7873 (N_7873,N_7566,N_7502);
and U7874 (N_7874,N_7579,N_7534);
and U7875 (N_7875,N_7589,N_7696);
nand U7876 (N_7876,N_7613,N_7557);
nand U7877 (N_7877,N_7569,N_7719);
xor U7878 (N_7878,N_7592,N_7519);
nor U7879 (N_7879,N_7646,N_7738);
and U7880 (N_7880,N_7743,N_7639);
or U7881 (N_7881,N_7616,N_7638);
nor U7882 (N_7882,N_7560,N_7719);
nor U7883 (N_7883,N_7573,N_7529);
or U7884 (N_7884,N_7713,N_7603);
nor U7885 (N_7885,N_7519,N_7716);
nand U7886 (N_7886,N_7683,N_7689);
or U7887 (N_7887,N_7712,N_7735);
or U7888 (N_7888,N_7616,N_7601);
and U7889 (N_7889,N_7563,N_7588);
nor U7890 (N_7890,N_7524,N_7701);
nor U7891 (N_7891,N_7696,N_7618);
or U7892 (N_7892,N_7575,N_7709);
and U7893 (N_7893,N_7532,N_7643);
nand U7894 (N_7894,N_7615,N_7555);
xor U7895 (N_7895,N_7691,N_7733);
and U7896 (N_7896,N_7688,N_7701);
nor U7897 (N_7897,N_7642,N_7570);
and U7898 (N_7898,N_7651,N_7671);
or U7899 (N_7899,N_7744,N_7613);
xor U7900 (N_7900,N_7583,N_7697);
nand U7901 (N_7901,N_7506,N_7631);
and U7902 (N_7902,N_7603,N_7583);
xor U7903 (N_7903,N_7727,N_7550);
or U7904 (N_7904,N_7525,N_7683);
nor U7905 (N_7905,N_7520,N_7635);
nand U7906 (N_7906,N_7626,N_7727);
xnor U7907 (N_7907,N_7523,N_7594);
nor U7908 (N_7908,N_7567,N_7725);
nand U7909 (N_7909,N_7609,N_7599);
xor U7910 (N_7910,N_7657,N_7740);
nand U7911 (N_7911,N_7621,N_7682);
and U7912 (N_7912,N_7695,N_7570);
nor U7913 (N_7913,N_7526,N_7727);
nor U7914 (N_7914,N_7521,N_7687);
xnor U7915 (N_7915,N_7537,N_7710);
nand U7916 (N_7916,N_7687,N_7642);
xor U7917 (N_7917,N_7561,N_7565);
nor U7918 (N_7918,N_7623,N_7512);
xnor U7919 (N_7919,N_7621,N_7529);
and U7920 (N_7920,N_7559,N_7740);
or U7921 (N_7921,N_7726,N_7528);
nor U7922 (N_7922,N_7513,N_7623);
nand U7923 (N_7923,N_7724,N_7603);
or U7924 (N_7924,N_7740,N_7671);
xor U7925 (N_7925,N_7573,N_7506);
xnor U7926 (N_7926,N_7685,N_7687);
nand U7927 (N_7927,N_7733,N_7520);
nand U7928 (N_7928,N_7673,N_7565);
nand U7929 (N_7929,N_7688,N_7518);
or U7930 (N_7930,N_7716,N_7508);
and U7931 (N_7931,N_7672,N_7705);
nand U7932 (N_7932,N_7508,N_7741);
and U7933 (N_7933,N_7583,N_7658);
and U7934 (N_7934,N_7700,N_7603);
xor U7935 (N_7935,N_7541,N_7520);
nand U7936 (N_7936,N_7663,N_7647);
nor U7937 (N_7937,N_7540,N_7565);
nor U7938 (N_7938,N_7634,N_7713);
or U7939 (N_7939,N_7661,N_7634);
nand U7940 (N_7940,N_7691,N_7572);
xor U7941 (N_7941,N_7519,N_7685);
xnor U7942 (N_7942,N_7634,N_7696);
nor U7943 (N_7943,N_7527,N_7578);
or U7944 (N_7944,N_7642,N_7594);
nand U7945 (N_7945,N_7636,N_7730);
xor U7946 (N_7946,N_7550,N_7603);
nor U7947 (N_7947,N_7620,N_7653);
nor U7948 (N_7948,N_7648,N_7504);
and U7949 (N_7949,N_7550,N_7698);
nor U7950 (N_7950,N_7606,N_7734);
and U7951 (N_7951,N_7742,N_7549);
xor U7952 (N_7952,N_7742,N_7704);
xor U7953 (N_7953,N_7652,N_7522);
and U7954 (N_7954,N_7729,N_7682);
xor U7955 (N_7955,N_7628,N_7691);
xor U7956 (N_7956,N_7501,N_7621);
and U7957 (N_7957,N_7666,N_7571);
nor U7958 (N_7958,N_7653,N_7571);
nor U7959 (N_7959,N_7643,N_7574);
nor U7960 (N_7960,N_7576,N_7635);
xor U7961 (N_7961,N_7740,N_7695);
and U7962 (N_7962,N_7609,N_7522);
or U7963 (N_7963,N_7526,N_7536);
nor U7964 (N_7964,N_7571,N_7634);
or U7965 (N_7965,N_7705,N_7530);
and U7966 (N_7966,N_7726,N_7565);
and U7967 (N_7967,N_7513,N_7642);
nor U7968 (N_7968,N_7561,N_7741);
xor U7969 (N_7969,N_7602,N_7598);
xor U7970 (N_7970,N_7563,N_7707);
xnor U7971 (N_7971,N_7641,N_7522);
and U7972 (N_7972,N_7572,N_7727);
and U7973 (N_7973,N_7531,N_7532);
nand U7974 (N_7974,N_7590,N_7632);
xnor U7975 (N_7975,N_7561,N_7748);
nor U7976 (N_7976,N_7655,N_7747);
nand U7977 (N_7977,N_7617,N_7597);
nand U7978 (N_7978,N_7642,N_7653);
xor U7979 (N_7979,N_7621,N_7533);
nor U7980 (N_7980,N_7704,N_7548);
and U7981 (N_7981,N_7632,N_7666);
nand U7982 (N_7982,N_7631,N_7728);
nand U7983 (N_7983,N_7625,N_7599);
xor U7984 (N_7984,N_7583,N_7627);
nand U7985 (N_7985,N_7741,N_7676);
and U7986 (N_7986,N_7582,N_7608);
nor U7987 (N_7987,N_7680,N_7603);
nand U7988 (N_7988,N_7536,N_7653);
and U7989 (N_7989,N_7576,N_7688);
nor U7990 (N_7990,N_7599,N_7573);
nor U7991 (N_7991,N_7593,N_7717);
and U7992 (N_7992,N_7659,N_7627);
nor U7993 (N_7993,N_7714,N_7519);
nand U7994 (N_7994,N_7705,N_7736);
or U7995 (N_7995,N_7523,N_7738);
nor U7996 (N_7996,N_7579,N_7580);
xor U7997 (N_7997,N_7745,N_7619);
nand U7998 (N_7998,N_7641,N_7534);
xor U7999 (N_7999,N_7613,N_7528);
and U8000 (N_8000,N_7972,N_7874);
nand U8001 (N_8001,N_7992,N_7904);
nand U8002 (N_8002,N_7792,N_7888);
nand U8003 (N_8003,N_7833,N_7785);
xnor U8004 (N_8004,N_7879,N_7867);
and U8005 (N_8005,N_7980,N_7922);
nand U8006 (N_8006,N_7951,N_7887);
nor U8007 (N_8007,N_7801,N_7771);
and U8008 (N_8008,N_7805,N_7871);
nor U8009 (N_8009,N_7851,N_7819);
nor U8010 (N_8010,N_7962,N_7832);
nor U8011 (N_8011,N_7994,N_7956);
xor U8012 (N_8012,N_7966,N_7919);
nand U8013 (N_8013,N_7765,N_7979);
nor U8014 (N_8014,N_7913,N_7760);
xor U8015 (N_8015,N_7827,N_7866);
nor U8016 (N_8016,N_7897,N_7752);
or U8017 (N_8017,N_7820,N_7903);
or U8018 (N_8018,N_7842,N_7931);
or U8019 (N_8019,N_7935,N_7848);
and U8020 (N_8020,N_7877,N_7804);
or U8021 (N_8021,N_7818,N_7822);
xor U8022 (N_8022,N_7770,N_7876);
and U8023 (N_8023,N_7778,N_7774);
or U8024 (N_8024,N_7901,N_7787);
and U8025 (N_8025,N_7795,N_7756);
nor U8026 (N_8026,N_7939,N_7790);
nor U8027 (N_8027,N_7831,N_7784);
or U8028 (N_8028,N_7880,N_7912);
and U8029 (N_8029,N_7969,N_7996);
or U8030 (N_8030,N_7948,N_7862);
nand U8031 (N_8031,N_7967,N_7934);
xor U8032 (N_8032,N_7991,N_7970);
nand U8033 (N_8033,N_7961,N_7773);
nor U8034 (N_8034,N_7859,N_7834);
or U8035 (N_8035,N_7786,N_7872);
xnor U8036 (N_8036,N_7796,N_7989);
and U8037 (N_8037,N_7844,N_7830);
or U8038 (N_8038,N_7810,N_7797);
xnor U8039 (N_8039,N_7814,N_7767);
nor U8040 (N_8040,N_7769,N_7890);
xor U8041 (N_8041,N_7793,N_7998);
or U8042 (N_8042,N_7849,N_7963);
nand U8043 (N_8043,N_7825,N_7800);
xnor U8044 (N_8044,N_7855,N_7986);
and U8045 (N_8045,N_7853,N_7821);
xor U8046 (N_8046,N_7753,N_7858);
nand U8047 (N_8047,N_7780,N_7852);
or U8048 (N_8048,N_7828,N_7813);
and U8049 (N_8049,N_7794,N_7873);
and U8050 (N_8050,N_7987,N_7841);
and U8051 (N_8051,N_7905,N_7899);
nor U8052 (N_8052,N_7911,N_7781);
and U8053 (N_8053,N_7940,N_7918);
or U8054 (N_8054,N_7847,N_7840);
nor U8055 (N_8055,N_7789,N_7755);
nor U8056 (N_8056,N_7754,N_7910);
and U8057 (N_8057,N_7863,N_7788);
and U8058 (N_8058,N_7983,N_7772);
nor U8059 (N_8059,N_7898,N_7806);
nand U8060 (N_8060,N_7869,N_7809);
or U8061 (N_8061,N_7947,N_7791);
or U8062 (N_8062,N_7777,N_7955);
and U8063 (N_8063,N_7843,N_7977);
xor U8064 (N_8064,N_7757,N_7938);
and U8065 (N_8065,N_7836,N_7928);
xor U8066 (N_8066,N_7988,N_7953);
and U8067 (N_8067,N_7763,N_7895);
nand U8068 (N_8068,N_7826,N_7857);
or U8069 (N_8069,N_7875,N_7783);
nor U8070 (N_8070,N_7949,N_7817);
xnor U8071 (N_8071,N_7933,N_7926);
and U8072 (N_8072,N_7957,N_7802);
or U8073 (N_8073,N_7930,N_7960);
nor U8074 (N_8074,N_7835,N_7891);
or U8075 (N_8075,N_7838,N_7878);
or U8076 (N_8076,N_7982,N_7997);
and U8077 (N_8077,N_7837,N_7846);
xnor U8078 (N_8078,N_7968,N_7950);
and U8079 (N_8079,N_7975,N_7812);
or U8080 (N_8080,N_7807,N_7808);
nor U8081 (N_8081,N_7883,N_7750);
or U8082 (N_8082,N_7854,N_7782);
nor U8083 (N_8083,N_7965,N_7860);
nor U8084 (N_8084,N_7909,N_7892);
xnor U8085 (N_8085,N_7751,N_7758);
or U8086 (N_8086,N_7959,N_7929);
or U8087 (N_8087,N_7984,N_7954);
nor U8088 (N_8088,N_7824,N_7845);
and U8089 (N_8089,N_7973,N_7829);
nand U8090 (N_8090,N_7759,N_7946);
nand U8091 (N_8091,N_7945,N_7775);
or U8092 (N_8092,N_7896,N_7868);
or U8093 (N_8093,N_7850,N_7902);
xnor U8094 (N_8094,N_7811,N_7942);
and U8095 (N_8095,N_7976,N_7870);
and U8096 (N_8096,N_7971,N_7943);
xnor U8097 (N_8097,N_7861,N_7906);
or U8098 (N_8098,N_7764,N_7761);
nand U8099 (N_8099,N_7920,N_7974);
nor U8100 (N_8100,N_7856,N_7958);
nor U8101 (N_8101,N_7907,N_7839);
or U8102 (N_8102,N_7944,N_7889);
nand U8103 (N_8103,N_7978,N_7936);
and U8104 (N_8104,N_7925,N_7941);
nor U8105 (N_8105,N_7999,N_7816);
and U8106 (N_8106,N_7916,N_7884);
xor U8107 (N_8107,N_7865,N_7927);
nor U8108 (N_8108,N_7921,N_7981);
nor U8109 (N_8109,N_7937,N_7893);
nand U8110 (N_8110,N_7995,N_7815);
nor U8111 (N_8111,N_7924,N_7779);
nand U8112 (N_8112,N_7803,N_7894);
nand U8113 (N_8113,N_7799,N_7864);
nor U8114 (N_8114,N_7993,N_7990);
nor U8115 (N_8115,N_7882,N_7932);
nor U8116 (N_8116,N_7823,N_7923);
and U8117 (N_8117,N_7881,N_7798);
nor U8118 (N_8118,N_7886,N_7766);
nand U8119 (N_8119,N_7985,N_7762);
nand U8120 (N_8120,N_7917,N_7908);
or U8121 (N_8121,N_7915,N_7768);
nand U8122 (N_8122,N_7914,N_7900);
nor U8123 (N_8123,N_7952,N_7885);
or U8124 (N_8124,N_7776,N_7964);
and U8125 (N_8125,N_7772,N_7854);
or U8126 (N_8126,N_7937,N_7979);
xor U8127 (N_8127,N_7948,N_7915);
nand U8128 (N_8128,N_7774,N_7819);
or U8129 (N_8129,N_7945,N_7756);
nand U8130 (N_8130,N_7780,N_7813);
or U8131 (N_8131,N_7812,N_7984);
nand U8132 (N_8132,N_7777,N_7867);
and U8133 (N_8133,N_7777,N_7865);
nand U8134 (N_8134,N_7774,N_7809);
nor U8135 (N_8135,N_7988,N_7984);
nor U8136 (N_8136,N_7765,N_7835);
nor U8137 (N_8137,N_7819,N_7881);
nor U8138 (N_8138,N_7859,N_7819);
and U8139 (N_8139,N_7830,N_7789);
nand U8140 (N_8140,N_7774,N_7961);
nand U8141 (N_8141,N_7968,N_7767);
and U8142 (N_8142,N_7886,N_7991);
and U8143 (N_8143,N_7779,N_7993);
xor U8144 (N_8144,N_7997,N_7931);
and U8145 (N_8145,N_7875,N_7958);
nor U8146 (N_8146,N_7763,N_7972);
and U8147 (N_8147,N_7844,N_7851);
and U8148 (N_8148,N_7864,N_7938);
and U8149 (N_8149,N_7905,N_7893);
xnor U8150 (N_8150,N_7989,N_7985);
nor U8151 (N_8151,N_7787,N_7776);
xor U8152 (N_8152,N_7955,N_7755);
nand U8153 (N_8153,N_7847,N_7848);
xnor U8154 (N_8154,N_7987,N_7781);
nand U8155 (N_8155,N_7988,N_7811);
or U8156 (N_8156,N_7825,N_7824);
or U8157 (N_8157,N_7902,N_7913);
xnor U8158 (N_8158,N_7991,N_7864);
nand U8159 (N_8159,N_7766,N_7816);
or U8160 (N_8160,N_7945,N_7765);
xor U8161 (N_8161,N_7785,N_7953);
or U8162 (N_8162,N_7770,N_7899);
and U8163 (N_8163,N_7974,N_7859);
nand U8164 (N_8164,N_7841,N_7770);
xor U8165 (N_8165,N_7750,N_7955);
xor U8166 (N_8166,N_7826,N_7957);
and U8167 (N_8167,N_7985,N_7949);
nand U8168 (N_8168,N_7977,N_7996);
or U8169 (N_8169,N_7857,N_7909);
and U8170 (N_8170,N_7933,N_7844);
and U8171 (N_8171,N_7813,N_7966);
nand U8172 (N_8172,N_7915,N_7767);
nor U8173 (N_8173,N_7795,N_7990);
xnor U8174 (N_8174,N_7863,N_7943);
or U8175 (N_8175,N_7761,N_7936);
or U8176 (N_8176,N_7817,N_7833);
and U8177 (N_8177,N_7930,N_7890);
nand U8178 (N_8178,N_7932,N_7911);
nor U8179 (N_8179,N_7814,N_7967);
and U8180 (N_8180,N_7911,N_7931);
xor U8181 (N_8181,N_7810,N_7791);
xor U8182 (N_8182,N_7819,N_7997);
xnor U8183 (N_8183,N_7945,N_7813);
and U8184 (N_8184,N_7788,N_7848);
nand U8185 (N_8185,N_7900,N_7950);
nor U8186 (N_8186,N_7966,N_7994);
nand U8187 (N_8187,N_7926,N_7950);
and U8188 (N_8188,N_7821,N_7872);
nor U8189 (N_8189,N_7946,N_7855);
nor U8190 (N_8190,N_7786,N_7952);
or U8191 (N_8191,N_7830,N_7916);
or U8192 (N_8192,N_7795,N_7913);
nand U8193 (N_8193,N_7814,N_7824);
or U8194 (N_8194,N_7787,N_7965);
xor U8195 (N_8195,N_7765,N_7883);
and U8196 (N_8196,N_7798,N_7796);
xor U8197 (N_8197,N_7937,N_7847);
and U8198 (N_8198,N_7929,N_7835);
or U8199 (N_8199,N_7970,N_7773);
nor U8200 (N_8200,N_7783,N_7809);
and U8201 (N_8201,N_7828,N_7852);
or U8202 (N_8202,N_7997,N_7855);
or U8203 (N_8203,N_7788,N_7905);
nor U8204 (N_8204,N_7751,N_7841);
nand U8205 (N_8205,N_7764,N_7952);
and U8206 (N_8206,N_7814,N_7768);
xnor U8207 (N_8207,N_7831,N_7951);
or U8208 (N_8208,N_7939,N_7776);
and U8209 (N_8209,N_7892,N_7878);
xnor U8210 (N_8210,N_7873,N_7769);
xor U8211 (N_8211,N_7792,N_7910);
nor U8212 (N_8212,N_7860,N_7971);
and U8213 (N_8213,N_7932,N_7753);
nand U8214 (N_8214,N_7797,N_7849);
xnor U8215 (N_8215,N_7896,N_7780);
nor U8216 (N_8216,N_7798,N_7877);
nor U8217 (N_8217,N_7937,N_7878);
nor U8218 (N_8218,N_7780,N_7879);
nand U8219 (N_8219,N_7948,N_7870);
or U8220 (N_8220,N_7937,N_7904);
nand U8221 (N_8221,N_7947,N_7985);
nand U8222 (N_8222,N_7936,N_7777);
xnor U8223 (N_8223,N_7909,N_7862);
and U8224 (N_8224,N_7871,N_7894);
nor U8225 (N_8225,N_7928,N_7812);
xor U8226 (N_8226,N_7847,N_7793);
and U8227 (N_8227,N_7872,N_7820);
nor U8228 (N_8228,N_7790,N_7839);
and U8229 (N_8229,N_7768,N_7922);
xnor U8230 (N_8230,N_7764,N_7844);
nand U8231 (N_8231,N_7980,N_7770);
or U8232 (N_8232,N_7995,N_7884);
nand U8233 (N_8233,N_7974,N_7855);
or U8234 (N_8234,N_7816,N_7860);
nor U8235 (N_8235,N_7759,N_7878);
xor U8236 (N_8236,N_7783,N_7792);
and U8237 (N_8237,N_7804,N_7992);
and U8238 (N_8238,N_7959,N_7951);
xor U8239 (N_8239,N_7900,N_7815);
nor U8240 (N_8240,N_7924,N_7814);
and U8241 (N_8241,N_7891,N_7950);
and U8242 (N_8242,N_7817,N_7976);
xor U8243 (N_8243,N_7851,N_7839);
xnor U8244 (N_8244,N_7918,N_7983);
or U8245 (N_8245,N_7906,N_7899);
or U8246 (N_8246,N_7777,N_7946);
nand U8247 (N_8247,N_7983,N_7955);
nand U8248 (N_8248,N_7939,N_7817);
or U8249 (N_8249,N_7924,N_7939);
nand U8250 (N_8250,N_8106,N_8209);
or U8251 (N_8251,N_8164,N_8239);
xor U8252 (N_8252,N_8236,N_8098);
nor U8253 (N_8253,N_8223,N_8015);
or U8254 (N_8254,N_8060,N_8100);
and U8255 (N_8255,N_8027,N_8035);
nor U8256 (N_8256,N_8019,N_8123);
xnor U8257 (N_8257,N_8153,N_8119);
nand U8258 (N_8258,N_8232,N_8021);
nand U8259 (N_8259,N_8246,N_8029);
or U8260 (N_8260,N_8115,N_8125);
or U8261 (N_8261,N_8071,N_8079);
nand U8262 (N_8262,N_8216,N_8073);
or U8263 (N_8263,N_8101,N_8215);
and U8264 (N_8264,N_8137,N_8093);
or U8265 (N_8265,N_8247,N_8171);
and U8266 (N_8266,N_8003,N_8229);
nand U8267 (N_8267,N_8139,N_8046);
nor U8268 (N_8268,N_8032,N_8170);
and U8269 (N_8269,N_8110,N_8081);
and U8270 (N_8270,N_8054,N_8108);
or U8271 (N_8271,N_8152,N_8167);
nand U8272 (N_8272,N_8028,N_8002);
xor U8273 (N_8273,N_8127,N_8092);
xnor U8274 (N_8274,N_8086,N_8165);
or U8275 (N_8275,N_8234,N_8109);
nand U8276 (N_8276,N_8050,N_8243);
and U8277 (N_8277,N_8168,N_8180);
nor U8278 (N_8278,N_8175,N_8056);
nand U8279 (N_8279,N_8211,N_8131);
or U8280 (N_8280,N_8058,N_8169);
nor U8281 (N_8281,N_8087,N_8126);
xnor U8282 (N_8282,N_8096,N_8095);
nand U8283 (N_8283,N_8111,N_8117);
xor U8284 (N_8284,N_8065,N_8238);
and U8285 (N_8285,N_8121,N_8069);
nor U8286 (N_8286,N_8055,N_8136);
xnor U8287 (N_8287,N_8217,N_8141);
or U8288 (N_8288,N_8034,N_8160);
nor U8289 (N_8289,N_8059,N_8190);
nor U8290 (N_8290,N_8077,N_8072);
nor U8291 (N_8291,N_8147,N_8189);
xor U8292 (N_8292,N_8233,N_8205);
and U8293 (N_8293,N_8011,N_8207);
xnor U8294 (N_8294,N_8179,N_8241);
nor U8295 (N_8295,N_8157,N_8053);
and U8296 (N_8296,N_8161,N_8089);
or U8297 (N_8297,N_8154,N_8176);
and U8298 (N_8298,N_8016,N_8112);
and U8299 (N_8299,N_8074,N_8186);
nand U8300 (N_8300,N_8006,N_8178);
nor U8301 (N_8301,N_8138,N_8099);
nand U8302 (N_8302,N_8212,N_8222);
nand U8303 (N_8303,N_8064,N_8026);
and U8304 (N_8304,N_8018,N_8070);
or U8305 (N_8305,N_8103,N_8159);
xnor U8306 (N_8306,N_8200,N_8076);
xnor U8307 (N_8307,N_8094,N_8051);
or U8308 (N_8308,N_8067,N_8041);
xor U8309 (N_8309,N_8193,N_8184);
nand U8310 (N_8310,N_8085,N_8172);
and U8311 (N_8311,N_8210,N_8083);
or U8312 (N_8312,N_8090,N_8022);
and U8313 (N_8313,N_8155,N_8004);
nand U8314 (N_8314,N_8000,N_8057);
nand U8315 (N_8315,N_8088,N_8104);
nand U8316 (N_8316,N_8097,N_8230);
or U8317 (N_8317,N_8017,N_8005);
or U8318 (N_8318,N_8174,N_8078);
or U8319 (N_8319,N_8198,N_8197);
nor U8320 (N_8320,N_8033,N_8044);
and U8321 (N_8321,N_8196,N_8008);
nor U8322 (N_8322,N_8066,N_8105);
xnor U8323 (N_8323,N_8010,N_8128);
nand U8324 (N_8324,N_8062,N_8213);
nor U8325 (N_8325,N_8102,N_8208);
or U8326 (N_8326,N_8135,N_8226);
and U8327 (N_8327,N_8173,N_8091);
or U8328 (N_8328,N_8107,N_8195);
or U8329 (N_8329,N_8142,N_8231);
and U8330 (N_8330,N_8156,N_8237);
xnor U8331 (N_8331,N_8043,N_8151);
or U8332 (N_8332,N_8047,N_8012);
nor U8333 (N_8333,N_8129,N_8144);
and U8334 (N_8334,N_8235,N_8148);
nand U8335 (N_8335,N_8183,N_8052);
nand U8336 (N_8336,N_8218,N_8013);
nand U8337 (N_8337,N_8049,N_8202);
xor U8338 (N_8338,N_8166,N_8080);
nor U8339 (N_8339,N_8009,N_8162);
and U8340 (N_8340,N_8014,N_8206);
nand U8341 (N_8341,N_8158,N_8227);
nor U8342 (N_8342,N_8219,N_8201);
xnor U8343 (N_8343,N_8134,N_8038);
and U8344 (N_8344,N_8061,N_8225);
or U8345 (N_8345,N_8163,N_8140);
and U8346 (N_8346,N_8248,N_8113);
and U8347 (N_8347,N_8075,N_8084);
or U8348 (N_8348,N_8203,N_8036);
xor U8349 (N_8349,N_8191,N_8007);
nand U8350 (N_8350,N_8228,N_8181);
and U8351 (N_8351,N_8240,N_8045);
or U8352 (N_8352,N_8122,N_8187);
nor U8353 (N_8353,N_8177,N_8204);
and U8354 (N_8354,N_8224,N_8244);
xnor U8355 (N_8355,N_8040,N_8024);
and U8356 (N_8356,N_8242,N_8118);
nor U8357 (N_8357,N_8221,N_8023);
xnor U8358 (N_8358,N_8194,N_8120);
xnor U8359 (N_8359,N_8146,N_8132);
xor U8360 (N_8360,N_8249,N_8020);
nand U8361 (N_8361,N_8001,N_8082);
xor U8362 (N_8362,N_8245,N_8063);
nor U8363 (N_8363,N_8199,N_8116);
or U8364 (N_8364,N_8149,N_8042);
or U8365 (N_8365,N_8037,N_8182);
and U8366 (N_8366,N_8150,N_8220);
nor U8367 (N_8367,N_8192,N_8214);
and U8368 (N_8368,N_8030,N_8124);
or U8369 (N_8369,N_8031,N_8133);
and U8370 (N_8370,N_8185,N_8048);
nand U8371 (N_8371,N_8143,N_8145);
or U8372 (N_8372,N_8025,N_8039);
nand U8373 (N_8373,N_8188,N_8130);
or U8374 (N_8374,N_8068,N_8114);
and U8375 (N_8375,N_8015,N_8112);
xnor U8376 (N_8376,N_8047,N_8092);
and U8377 (N_8377,N_8157,N_8043);
or U8378 (N_8378,N_8060,N_8164);
xor U8379 (N_8379,N_8106,N_8208);
or U8380 (N_8380,N_8035,N_8111);
nor U8381 (N_8381,N_8018,N_8208);
or U8382 (N_8382,N_8006,N_8059);
nand U8383 (N_8383,N_8240,N_8042);
or U8384 (N_8384,N_8032,N_8204);
xnor U8385 (N_8385,N_8007,N_8071);
and U8386 (N_8386,N_8124,N_8074);
xnor U8387 (N_8387,N_8014,N_8039);
nand U8388 (N_8388,N_8160,N_8158);
or U8389 (N_8389,N_8117,N_8168);
and U8390 (N_8390,N_8226,N_8121);
and U8391 (N_8391,N_8117,N_8047);
or U8392 (N_8392,N_8113,N_8132);
xor U8393 (N_8393,N_8126,N_8013);
or U8394 (N_8394,N_8197,N_8217);
xnor U8395 (N_8395,N_8191,N_8128);
or U8396 (N_8396,N_8154,N_8190);
or U8397 (N_8397,N_8115,N_8199);
xor U8398 (N_8398,N_8226,N_8164);
xnor U8399 (N_8399,N_8020,N_8233);
and U8400 (N_8400,N_8075,N_8159);
nand U8401 (N_8401,N_8007,N_8009);
or U8402 (N_8402,N_8062,N_8001);
nand U8403 (N_8403,N_8016,N_8199);
nor U8404 (N_8404,N_8185,N_8197);
or U8405 (N_8405,N_8092,N_8099);
nand U8406 (N_8406,N_8008,N_8213);
and U8407 (N_8407,N_8137,N_8189);
xor U8408 (N_8408,N_8085,N_8123);
xnor U8409 (N_8409,N_8228,N_8217);
nor U8410 (N_8410,N_8230,N_8009);
nor U8411 (N_8411,N_8027,N_8119);
nor U8412 (N_8412,N_8079,N_8026);
or U8413 (N_8413,N_8026,N_8073);
and U8414 (N_8414,N_8249,N_8184);
xor U8415 (N_8415,N_8086,N_8208);
nand U8416 (N_8416,N_8066,N_8106);
nor U8417 (N_8417,N_8240,N_8010);
xor U8418 (N_8418,N_8105,N_8210);
xor U8419 (N_8419,N_8020,N_8075);
nand U8420 (N_8420,N_8018,N_8058);
or U8421 (N_8421,N_8246,N_8210);
nand U8422 (N_8422,N_8226,N_8036);
nand U8423 (N_8423,N_8167,N_8091);
xor U8424 (N_8424,N_8202,N_8230);
nor U8425 (N_8425,N_8185,N_8003);
and U8426 (N_8426,N_8002,N_8067);
xnor U8427 (N_8427,N_8080,N_8081);
xor U8428 (N_8428,N_8087,N_8010);
nor U8429 (N_8429,N_8230,N_8031);
nand U8430 (N_8430,N_8132,N_8061);
and U8431 (N_8431,N_8129,N_8164);
xnor U8432 (N_8432,N_8055,N_8188);
and U8433 (N_8433,N_8128,N_8177);
nand U8434 (N_8434,N_8068,N_8017);
or U8435 (N_8435,N_8078,N_8025);
nor U8436 (N_8436,N_8247,N_8137);
nand U8437 (N_8437,N_8064,N_8225);
nand U8438 (N_8438,N_8184,N_8130);
xnor U8439 (N_8439,N_8021,N_8208);
and U8440 (N_8440,N_8086,N_8068);
nand U8441 (N_8441,N_8034,N_8148);
xnor U8442 (N_8442,N_8186,N_8026);
xor U8443 (N_8443,N_8202,N_8062);
and U8444 (N_8444,N_8078,N_8171);
and U8445 (N_8445,N_8083,N_8188);
and U8446 (N_8446,N_8150,N_8021);
and U8447 (N_8447,N_8152,N_8019);
nor U8448 (N_8448,N_8009,N_8227);
or U8449 (N_8449,N_8177,N_8197);
xnor U8450 (N_8450,N_8084,N_8188);
nor U8451 (N_8451,N_8211,N_8185);
xor U8452 (N_8452,N_8005,N_8227);
or U8453 (N_8453,N_8237,N_8057);
nand U8454 (N_8454,N_8199,N_8210);
and U8455 (N_8455,N_8196,N_8220);
nand U8456 (N_8456,N_8058,N_8039);
xor U8457 (N_8457,N_8052,N_8149);
xnor U8458 (N_8458,N_8055,N_8035);
xnor U8459 (N_8459,N_8030,N_8192);
and U8460 (N_8460,N_8177,N_8117);
or U8461 (N_8461,N_8158,N_8052);
xor U8462 (N_8462,N_8028,N_8101);
nor U8463 (N_8463,N_8065,N_8086);
or U8464 (N_8464,N_8187,N_8084);
nand U8465 (N_8465,N_8132,N_8075);
nor U8466 (N_8466,N_8129,N_8085);
nand U8467 (N_8467,N_8022,N_8092);
and U8468 (N_8468,N_8016,N_8119);
nand U8469 (N_8469,N_8091,N_8121);
xnor U8470 (N_8470,N_8211,N_8115);
xor U8471 (N_8471,N_8010,N_8141);
nand U8472 (N_8472,N_8083,N_8052);
nand U8473 (N_8473,N_8113,N_8150);
or U8474 (N_8474,N_8098,N_8202);
nand U8475 (N_8475,N_8097,N_8246);
xnor U8476 (N_8476,N_8059,N_8228);
and U8477 (N_8477,N_8052,N_8147);
and U8478 (N_8478,N_8022,N_8193);
or U8479 (N_8479,N_8225,N_8184);
nor U8480 (N_8480,N_8019,N_8003);
or U8481 (N_8481,N_8122,N_8019);
xnor U8482 (N_8482,N_8175,N_8232);
xnor U8483 (N_8483,N_8219,N_8231);
nand U8484 (N_8484,N_8167,N_8121);
or U8485 (N_8485,N_8229,N_8220);
or U8486 (N_8486,N_8028,N_8033);
and U8487 (N_8487,N_8162,N_8121);
and U8488 (N_8488,N_8045,N_8086);
and U8489 (N_8489,N_8026,N_8232);
or U8490 (N_8490,N_8192,N_8110);
nand U8491 (N_8491,N_8206,N_8132);
or U8492 (N_8492,N_8160,N_8129);
nand U8493 (N_8493,N_8217,N_8231);
or U8494 (N_8494,N_8223,N_8048);
xnor U8495 (N_8495,N_8105,N_8152);
nor U8496 (N_8496,N_8001,N_8117);
or U8497 (N_8497,N_8065,N_8184);
xnor U8498 (N_8498,N_8010,N_8174);
xnor U8499 (N_8499,N_8205,N_8148);
nand U8500 (N_8500,N_8327,N_8433);
nand U8501 (N_8501,N_8300,N_8470);
or U8502 (N_8502,N_8342,N_8456);
or U8503 (N_8503,N_8460,N_8288);
xor U8504 (N_8504,N_8291,N_8398);
or U8505 (N_8505,N_8429,N_8446);
nand U8506 (N_8506,N_8266,N_8310);
or U8507 (N_8507,N_8413,N_8337);
or U8508 (N_8508,N_8445,N_8442);
nand U8509 (N_8509,N_8269,N_8478);
xnor U8510 (N_8510,N_8312,N_8280);
and U8511 (N_8511,N_8383,N_8307);
nand U8512 (N_8512,N_8338,N_8382);
nand U8513 (N_8513,N_8287,N_8279);
nand U8514 (N_8514,N_8302,N_8325);
nor U8515 (N_8515,N_8319,N_8360);
xor U8516 (N_8516,N_8362,N_8485);
and U8517 (N_8517,N_8309,N_8254);
or U8518 (N_8518,N_8306,N_8397);
nand U8519 (N_8519,N_8286,N_8355);
nor U8520 (N_8520,N_8381,N_8268);
or U8521 (N_8521,N_8444,N_8396);
xor U8522 (N_8522,N_8476,N_8466);
nand U8523 (N_8523,N_8469,N_8258);
xnor U8524 (N_8524,N_8465,N_8467);
nor U8525 (N_8525,N_8441,N_8384);
nand U8526 (N_8526,N_8411,N_8377);
or U8527 (N_8527,N_8452,N_8453);
nor U8528 (N_8528,N_8435,N_8353);
nor U8529 (N_8529,N_8499,N_8332);
nor U8530 (N_8530,N_8431,N_8263);
and U8531 (N_8531,N_8252,N_8428);
xor U8532 (N_8532,N_8359,N_8492);
xnor U8533 (N_8533,N_8474,N_8371);
or U8534 (N_8534,N_8289,N_8424);
nand U8535 (N_8535,N_8490,N_8494);
or U8536 (N_8536,N_8387,N_8255);
or U8537 (N_8537,N_8471,N_8451);
xor U8538 (N_8538,N_8294,N_8251);
nor U8539 (N_8539,N_8393,N_8409);
and U8540 (N_8540,N_8367,N_8295);
and U8541 (N_8541,N_8482,N_8361);
nand U8542 (N_8542,N_8285,N_8407);
and U8543 (N_8543,N_8496,N_8417);
or U8544 (N_8544,N_8329,N_8425);
nor U8545 (N_8545,N_8434,N_8366);
or U8546 (N_8546,N_8260,N_8489);
xor U8547 (N_8547,N_8497,N_8349);
xor U8548 (N_8548,N_8438,N_8498);
nor U8549 (N_8549,N_8418,N_8457);
or U8550 (N_8550,N_8394,N_8298);
or U8551 (N_8551,N_8278,N_8345);
or U8552 (N_8552,N_8473,N_8430);
or U8553 (N_8553,N_8399,N_8437);
nand U8554 (N_8554,N_8330,N_8380);
xnor U8555 (N_8555,N_8358,N_8282);
xor U8556 (N_8556,N_8369,N_8324);
nand U8557 (N_8557,N_8250,N_8270);
nor U8558 (N_8558,N_8322,N_8406);
xor U8559 (N_8559,N_8314,N_8326);
xnor U8560 (N_8560,N_8475,N_8386);
xnor U8561 (N_8561,N_8400,N_8283);
xnor U8562 (N_8562,N_8370,N_8459);
nor U8563 (N_8563,N_8480,N_8422);
nor U8564 (N_8564,N_8313,N_8363);
or U8565 (N_8565,N_8426,N_8305);
or U8566 (N_8566,N_8472,N_8373);
and U8567 (N_8567,N_8368,N_8292);
nor U8568 (N_8568,N_8331,N_8419);
xor U8569 (N_8569,N_8388,N_8341);
xnor U8570 (N_8570,N_8495,N_8253);
and U8571 (N_8571,N_8436,N_8454);
xor U8572 (N_8572,N_8448,N_8439);
nor U8573 (N_8573,N_8281,N_8262);
nor U8574 (N_8574,N_8346,N_8311);
nand U8575 (N_8575,N_8462,N_8317);
nand U8576 (N_8576,N_8450,N_8333);
nor U8577 (N_8577,N_8390,N_8423);
or U8578 (N_8578,N_8410,N_8443);
and U8579 (N_8579,N_8449,N_8491);
or U8580 (N_8580,N_8356,N_8412);
xnor U8581 (N_8581,N_8320,N_8316);
and U8582 (N_8582,N_8484,N_8343);
and U8583 (N_8583,N_8354,N_8339);
and U8584 (N_8584,N_8364,N_8464);
and U8585 (N_8585,N_8277,N_8376);
nand U8586 (N_8586,N_8372,N_8318);
nor U8587 (N_8587,N_8335,N_8273);
nor U8588 (N_8588,N_8308,N_8321);
nor U8589 (N_8589,N_8259,N_8458);
nand U8590 (N_8590,N_8481,N_8303);
xnor U8591 (N_8591,N_8290,N_8304);
and U8592 (N_8592,N_8389,N_8274);
or U8593 (N_8593,N_8477,N_8440);
nand U8594 (N_8594,N_8344,N_8402);
and U8595 (N_8595,N_8416,N_8348);
nand U8596 (N_8596,N_8301,N_8340);
xor U8597 (N_8597,N_8275,N_8403);
or U8598 (N_8598,N_8378,N_8493);
or U8599 (N_8599,N_8264,N_8427);
or U8600 (N_8600,N_8455,N_8271);
nand U8601 (N_8601,N_8486,N_8272);
and U8602 (N_8602,N_8432,N_8296);
and U8603 (N_8603,N_8463,N_8265);
nand U8604 (N_8604,N_8488,N_8276);
nor U8605 (N_8605,N_8487,N_8351);
or U8606 (N_8606,N_8415,N_8420);
nor U8607 (N_8607,N_8357,N_8352);
and U8608 (N_8608,N_8350,N_8297);
xnor U8609 (N_8609,N_8334,N_8483);
nor U8610 (N_8610,N_8421,N_8405);
xnor U8611 (N_8611,N_8256,N_8347);
and U8612 (N_8612,N_8392,N_8447);
xor U8613 (N_8613,N_8328,N_8375);
nand U8614 (N_8614,N_8336,N_8261);
nand U8615 (N_8615,N_8468,N_8374);
nor U8616 (N_8616,N_8293,N_8408);
and U8617 (N_8617,N_8315,N_8461);
and U8618 (N_8618,N_8299,N_8257);
nor U8619 (N_8619,N_8391,N_8379);
xor U8620 (N_8620,N_8479,N_8395);
nor U8621 (N_8621,N_8401,N_8404);
or U8622 (N_8622,N_8385,N_8365);
or U8623 (N_8623,N_8323,N_8284);
or U8624 (N_8624,N_8414,N_8267);
nor U8625 (N_8625,N_8407,N_8487);
xor U8626 (N_8626,N_8475,N_8497);
and U8627 (N_8627,N_8444,N_8355);
nand U8628 (N_8628,N_8364,N_8353);
xor U8629 (N_8629,N_8268,N_8380);
nor U8630 (N_8630,N_8368,N_8416);
xor U8631 (N_8631,N_8421,N_8298);
nor U8632 (N_8632,N_8455,N_8364);
or U8633 (N_8633,N_8365,N_8282);
and U8634 (N_8634,N_8263,N_8486);
nor U8635 (N_8635,N_8423,N_8496);
and U8636 (N_8636,N_8297,N_8420);
xor U8637 (N_8637,N_8460,N_8484);
nand U8638 (N_8638,N_8397,N_8448);
nor U8639 (N_8639,N_8449,N_8414);
xor U8640 (N_8640,N_8262,N_8474);
nor U8641 (N_8641,N_8262,N_8306);
or U8642 (N_8642,N_8368,N_8346);
nor U8643 (N_8643,N_8356,N_8376);
nor U8644 (N_8644,N_8296,N_8294);
nor U8645 (N_8645,N_8336,N_8415);
nand U8646 (N_8646,N_8424,N_8329);
or U8647 (N_8647,N_8400,N_8382);
nor U8648 (N_8648,N_8466,N_8434);
and U8649 (N_8649,N_8492,N_8481);
xnor U8650 (N_8650,N_8451,N_8379);
or U8651 (N_8651,N_8436,N_8255);
and U8652 (N_8652,N_8481,N_8261);
or U8653 (N_8653,N_8426,N_8462);
or U8654 (N_8654,N_8356,N_8484);
nand U8655 (N_8655,N_8427,N_8367);
xor U8656 (N_8656,N_8452,N_8439);
or U8657 (N_8657,N_8418,N_8490);
nand U8658 (N_8658,N_8323,N_8460);
xor U8659 (N_8659,N_8283,N_8406);
or U8660 (N_8660,N_8339,N_8315);
and U8661 (N_8661,N_8281,N_8434);
xnor U8662 (N_8662,N_8338,N_8453);
and U8663 (N_8663,N_8343,N_8262);
nor U8664 (N_8664,N_8399,N_8261);
or U8665 (N_8665,N_8261,N_8400);
nor U8666 (N_8666,N_8363,N_8268);
and U8667 (N_8667,N_8434,N_8365);
nand U8668 (N_8668,N_8460,N_8408);
nand U8669 (N_8669,N_8466,N_8481);
and U8670 (N_8670,N_8461,N_8375);
or U8671 (N_8671,N_8286,N_8493);
and U8672 (N_8672,N_8450,N_8296);
xnor U8673 (N_8673,N_8480,N_8383);
and U8674 (N_8674,N_8331,N_8362);
xor U8675 (N_8675,N_8418,N_8383);
xnor U8676 (N_8676,N_8498,N_8435);
and U8677 (N_8677,N_8294,N_8448);
xor U8678 (N_8678,N_8347,N_8436);
and U8679 (N_8679,N_8372,N_8347);
xor U8680 (N_8680,N_8291,N_8494);
nor U8681 (N_8681,N_8319,N_8351);
or U8682 (N_8682,N_8253,N_8379);
xor U8683 (N_8683,N_8447,N_8299);
xor U8684 (N_8684,N_8344,N_8473);
nand U8685 (N_8685,N_8429,N_8454);
nand U8686 (N_8686,N_8371,N_8448);
nand U8687 (N_8687,N_8284,N_8418);
or U8688 (N_8688,N_8301,N_8353);
nand U8689 (N_8689,N_8347,N_8434);
nor U8690 (N_8690,N_8368,N_8338);
nand U8691 (N_8691,N_8316,N_8255);
and U8692 (N_8692,N_8317,N_8398);
nand U8693 (N_8693,N_8299,N_8259);
xnor U8694 (N_8694,N_8252,N_8426);
xor U8695 (N_8695,N_8475,N_8385);
xnor U8696 (N_8696,N_8481,N_8468);
xor U8697 (N_8697,N_8395,N_8254);
or U8698 (N_8698,N_8360,N_8304);
nand U8699 (N_8699,N_8443,N_8302);
and U8700 (N_8700,N_8301,N_8300);
or U8701 (N_8701,N_8269,N_8304);
or U8702 (N_8702,N_8257,N_8315);
nor U8703 (N_8703,N_8408,N_8432);
xor U8704 (N_8704,N_8345,N_8437);
or U8705 (N_8705,N_8266,N_8302);
nor U8706 (N_8706,N_8352,N_8326);
nor U8707 (N_8707,N_8499,N_8402);
or U8708 (N_8708,N_8379,N_8400);
nor U8709 (N_8709,N_8289,N_8478);
or U8710 (N_8710,N_8276,N_8288);
xnor U8711 (N_8711,N_8459,N_8492);
and U8712 (N_8712,N_8497,N_8288);
or U8713 (N_8713,N_8250,N_8328);
or U8714 (N_8714,N_8285,N_8359);
nand U8715 (N_8715,N_8386,N_8499);
or U8716 (N_8716,N_8267,N_8478);
or U8717 (N_8717,N_8296,N_8379);
or U8718 (N_8718,N_8320,N_8420);
and U8719 (N_8719,N_8357,N_8324);
and U8720 (N_8720,N_8482,N_8481);
or U8721 (N_8721,N_8335,N_8498);
and U8722 (N_8722,N_8467,N_8459);
nand U8723 (N_8723,N_8327,N_8439);
xnor U8724 (N_8724,N_8433,N_8373);
nor U8725 (N_8725,N_8370,N_8385);
or U8726 (N_8726,N_8480,N_8262);
or U8727 (N_8727,N_8412,N_8458);
and U8728 (N_8728,N_8300,N_8314);
and U8729 (N_8729,N_8342,N_8499);
nor U8730 (N_8730,N_8411,N_8479);
nand U8731 (N_8731,N_8438,N_8333);
nor U8732 (N_8732,N_8339,N_8427);
xor U8733 (N_8733,N_8471,N_8290);
nor U8734 (N_8734,N_8310,N_8483);
nand U8735 (N_8735,N_8391,N_8359);
or U8736 (N_8736,N_8388,N_8278);
or U8737 (N_8737,N_8436,N_8419);
nand U8738 (N_8738,N_8278,N_8323);
nor U8739 (N_8739,N_8286,N_8351);
nand U8740 (N_8740,N_8378,N_8361);
nand U8741 (N_8741,N_8386,N_8322);
nand U8742 (N_8742,N_8266,N_8485);
and U8743 (N_8743,N_8475,N_8498);
xnor U8744 (N_8744,N_8340,N_8409);
nand U8745 (N_8745,N_8254,N_8345);
nor U8746 (N_8746,N_8379,N_8346);
nor U8747 (N_8747,N_8425,N_8334);
nand U8748 (N_8748,N_8353,N_8426);
nor U8749 (N_8749,N_8481,N_8279);
nor U8750 (N_8750,N_8531,N_8576);
or U8751 (N_8751,N_8674,N_8620);
nor U8752 (N_8752,N_8721,N_8544);
or U8753 (N_8753,N_8507,N_8600);
or U8754 (N_8754,N_8566,N_8680);
xnor U8755 (N_8755,N_8633,N_8505);
nor U8756 (N_8756,N_8520,N_8670);
nor U8757 (N_8757,N_8578,N_8725);
and U8758 (N_8758,N_8644,N_8693);
nand U8759 (N_8759,N_8603,N_8737);
nor U8760 (N_8760,N_8621,N_8573);
and U8761 (N_8761,N_8554,N_8589);
nand U8762 (N_8762,N_8515,N_8583);
nand U8763 (N_8763,N_8550,N_8524);
xnor U8764 (N_8764,N_8502,N_8614);
and U8765 (N_8765,N_8587,N_8658);
xor U8766 (N_8766,N_8581,N_8703);
nand U8767 (N_8767,N_8688,N_8555);
and U8768 (N_8768,N_8551,N_8729);
xor U8769 (N_8769,N_8570,N_8618);
nand U8770 (N_8770,N_8712,N_8749);
nor U8771 (N_8771,N_8637,N_8666);
or U8772 (N_8772,N_8536,N_8694);
and U8773 (N_8773,N_8707,N_8584);
and U8774 (N_8774,N_8696,N_8748);
or U8775 (N_8775,N_8636,N_8556);
nor U8776 (N_8776,N_8718,N_8728);
xnor U8777 (N_8777,N_8522,N_8529);
and U8778 (N_8778,N_8685,N_8663);
or U8779 (N_8779,N_8607,N_8501);
nand U8780 (N_8780,N_8526,N_8701);
nand U8781 (N_8781,N_8559,N_8738);
nand U8782 (N_8782,N_8653,N_8672);
or U8783 (N_8783,N_8604,N_8548);
nor U8784 (N_8784,N_8700,N_8683);
nand U8785 (N_8785,N_8572,N_8734);
or U8786 (N_8786,N_8588,N_8743);
or U8787 (N_8787,N_8617,N_8719);
and U8788 (N_8788,N_8552,N_8684);
xnor U8789 (N_8789,N_8528,N_8627);
and U8790 (N_8790,N_8730,N_8715);
nand U8791 (N_8791,N_8692,N_8597);
nor U8792 (N_8792,N_8652,N_8500);
and U8793 (N_8793,N_8648,N_8623);
nor U8794 (N_8794,N_8510,N_8537);
and U8795 (N_8795,N_8561,N_8586);
nor U8796 (N_8796,N_8558,N_8602);
nor U8797 (N_8797,N_8673,N_8532);
or U8798 (N_8798,N_8662,N_8521);
or U8799 (N_8799,N_8533,N_8651);
nor U8800 (N_8800,N_8699,N_8599);
or U8801 (N_8801,N_8682,N_8641);
nor U8802 (N_8802,N_8630,N_8654);
nor U8803 (N_8803,N_8562,N_8509);
and U8804 (N_8804,N_8628,N_8736);
nor U8805 (N_8805,N_8667,N_8690);
nand U8806 (N_8806,N_8545,N_8609);
nand U8807 (N_8807,N_8606,N_8676);
or U8808 (N_8808,N_8575,N_8540);
and U8809 (N_8809,N_8534,N_8669);
xnor U8810 (N_8810,N_8574,N_8514);
xor U8811 (N_8811,N_8677,N_8601);
or U8812 (N_8812,N_8634,N_8726);
or U8813 (N_8813,N_8649,N_8675);
or U8814 (N_8814,N_8741,N_8535);
nand U8815 (N_8815,N_8713,N_8733);
nor U8816 (N_8816,N_8625,N_8565);
and U8817 (N_8817,N_8527,N_8538);
nand U8818 (N_8818,N_8656,N_8513);
or U8819 (N_8819,N_8582,N_8643);
and U8820 (N_8820,N_8567,N_8580);
or U8821 (N_8821,N_8664,N_8632);
nor U8822 (N_8822,N_8516,N_8523);
or U8823 (N_8823,N_8506,N_8710);
or U8824 (N_8824,N_8747,N_8608);
nand U8825 (N_8825,N_8689,N_8503);
nand U8826 (N_8826,N_8731,N_8525);
nand U8827 (N_8827,N_8613,N_8705);
or U8828 (N_8828,N_8611,N_8563);
xnor U8829 (N_8829,N_8657,N_8504);
xor U8830 (N_8830,N_8708,N_8645);
and U8831 (N_8831,N_8619,N_8704);
nand U8832 (N_8832,N_8742,N_8724);
xnor U8833 (N_8833,N_8720,N_8592);
nand U8834 (N_8834,N_8711,N_8686);
or U8835 (N_8835,N_8542,N_8571);
nor U8836 (N_8836,N_8605,N_8569);
nand U8837 (N_8837,N_8629,N_8722);
or U8838 (N_8838,N_8596,N_8746);
nor U8839 (N_8839,N_8635,N_8547);
xor U8840 (N_8840,N_8650,N_8616);
nor U8841 (N_8841,N_8642,N_8671);
nand U8842 (N_8842,N_8665,N_8691);
and U8843 (N_8843,N_8744,N_8590);
nor U8844 (N_8844,N_8659,N_8511);
nor U8845 (N_8845,N_8622,N_8678);
nor U8846 (N_8846,N_8739,N_8647);
and U8847 (N_8847,N_8735,N_8557);
xnor U8848 (N_8848,N_8668,N_8591);
nand U8849 (N_8849,N_8518,N_8698);
nand U8850 (N_8850,N_8560,N_8661);
and U8851 (N_8851,N_8727,N_8530);
xnor U8852 (N_8852,N_8598,N_8626);
and U8853 (N_8853,N_8585,N_8695);
xnor U8854 (N_8854,N_8549,N_8702);
and U8855 (N_8855,N_8732,N_8508);
nor U8856 (N_8856,N_8517,N_8716);
or U8857 (N_8857,N_8723,N_8594);
and U8858 (N_8858,N_8745,N_8709);
xor U8859 (N_8859,N_8519,N_8660);
nor U8860 (N_8860,N_8595,N_8593);
or U8861 (N_8861,N_8541,N_8553);
nand U8862 (N_8862,N_8639,N_8697);
and U8863 (N_8863,N_8631,N_8546);
nor U8864 (N_8864,N_8714,N_8681);
nor U8865 (N_8865,N_8612,N_8577);
nand U8866 (N_8866,N_8706,N_8740);
or U8867 (N_8867,N_8512,N_8564);
xor U8868 (N_8868,N_8543,N_8679);
nand U8869 (N_8869,N_8640,N_8638);
nor U8870 (N_8870,N_8568,N_8655);
or U8871 (N_8871,N_8687,N_8615);
nand U8872 (N_8872,N_8610,N_8539);
nor U8873 (N_8873,N_8624,N_8579);
nand U8874 (N_8874,N_8646,N_8717);
nor U8875 (N_8875,N_8655,N_8703);
xnor U8876 (N_8876,N_8590,N_8710);
nor U8877 (N_8877,N_8589,N_8556);
nor U8878 (N_8878,N_8519,N_8524);
and U8879 (N_8879,N_8615,N_8633);
and U8880 (N_8880,N_8682,N_8729);
nand U8881 (N_8881,N_8527,N_8730);
nor U8882 (N_8882,N_8623,N_8586);
xnor U8883 (N_8883,N_8716,N_8738);
or U8884 (N_8884,N_8629,N_8679);
and U8885 (N_8885,N_8531,N_8509);
nor U8886 (N_8886,N_8695,N_8524);
or U8887 (N_8887,N_8670,N_8587);
or U8888 (N_8888,N_8539,N_8577);
nand U8889 (N_8889,N_8502,N_8720);
or U8890 (N_8890,N_8709,N_8500);
nor U8891 (N_8891,N_8551,N_8720);
nand U8892 (N_8892,N_8514,N_8579);
xor U8893 (N_8893,N_8578,N_8539);
and U8894 (N_8894,N_8633,N_8608);
nand U8895 (N_8895,N_8660,N_8702);
and U8896 (N_8896,N_8533,N_8652);
xnor U8897 (N_8897,N_8506,N_8623);
nor U8898 (N_8898,N_8735,N_8673);
xor U8899 (N_8899,N_8737,N_8649);
nand U8900 (N_8900,N_8620,N_8508);
or U8901 (N_8901,N_8639,N_8547);
nand U8902 (N_8902,N_8701,N_8515);
nand U8903 (N_8903,N_8693,N_8645);
and U8904 (N_8904,N_8628,N_8512);
nand U8905 (N_8905,N_8690,N_8747);
xor U8906 (N_8906,N_8614,N_8596);
xnor U8907 (N_8907,N_8714,N_8547);
xnor U8908 (N_8908,N_8648,N_8729);
nor U8909 (N_8909,N_8621,N_8607);
or U8910 (N_8910,N_8571,N_8506);
or U8911 (N_8911,N_8505,N_8613);
and U8912 (N_8912,N_8511,N_8678);
nand U8913 (N_8913,N_8691,N_8597);
nor U8914 (N_8914,N_8746,N_8502);
nor U8915 (N_8915,N_8702,N_8524);
xnor U8916 (N_8916,N_8502,N_8562);
nand U8917 (N_8917,N_8505,N_8641);
or U8918 (N_8918,N_8728,N_8694);
and U8919 (N_8919,N_8734,N_8511);
or U8920 (N_8920,N_8518,N_8531);
xnor U8921 (N_8921,N_8649,N_8524);
nor U8922 (N_8922,N_8543,N_8742);
xnor U8923 (N_8923,N_8526,N_8666);
or U8924 (N_8924,N_8670,N_8718);
nor U8925 (N_8925,N_8705,N_8738);
or U8926 (N_8926,N_8526,N_8565);
nor U8927 (N_8927,N_8652,N_8574);
or U8928 (N_8928,N_8529,N_8647);
xor U8929 (N_8929,N_8678,N_8713);
nand U8930 (N_8930,N_8719,N_8674);
nand U8931 (N_8931,N_8700,N_8550);
nor U8932 (N_8932,N_8657,N_8567);
nor U8933 (N_8933,N_8675,N_8744);
and U8934 (N_8934,N_8555,N_8696);
or U8935 (N_8935,N_8711,N_8712);
xor U8936 (N_8936,N_8663,N_8678);
nor U8937 (N_8937,N_8579,N_8591);
or U8938 (N_8938,N_8532,N_8559);
nand U8939 (N_8939,N_8561,N_8613);
or U8940 (N_8940,N_8718,N_8619);
nand U8941 (N_8941,N_8644,N_8536);
xnor U8942 (N_8942,N_8697,N_8663);
nor U8943 (N_8943,N_8579,N_8666);
or U8944 (N_8944,N_8712,N_8658);
and U8945 (N_8945,N_8524,N_8503);
nor U8946 (N_8946,N_8550,N_8749);
nand U8947 (N_8947,N_8552,N_8572);
nor U8948 (N_8948,N_8745,N_8551);
and U8949 (N_8949,N_8682,N_8701);
nor U8950 (N_8950,N_8659,N_8592);
or U8951 (N_8951,N_8592,N_8545);
and U8952 (N_8952,N_8507,N_8711);
nor U8953 (N_8953,N_8660,N_8614);
and U8954 (N_8954,N_8723,N_8504);
and U8955 (N_8955,N_8526,N_8616);
nor U8956 (N_8956,N_8577,N_8555);
xnor U8957 (N_8957,N_8573,N_8507);
nor U8958 (N_8958,N_8514,N_8682);
nand U8959 (N_8959,N_8500,N_8620);
nand U8960 (N_8960,N_8687,N_8660);
and U8961 (N_8961,N_8689,N_8550);
nor U8962 (N_8962,N_8639,N_8617);
xnor U8963 (N_8963,N_8534,N_8612);
nand U8964 (N_8964,N_8739,N_8533);
nor U8965 (N_8965,N_8645,N_8675);
nor U8966 (N_8966,N_8669,N_8729);
or U8967 (N_8967,N_8617,N_8559);
and U8968 (N_8968,N_8572,N_8627);
and U8969 (N_8969,N_8729,N_8511);
or U8970 (N_8970,N_8521,N_8538);
or U8971 (N_8971,N_8574,N_8616);
xnor U8972 (N_8972,N_8719,N_8668);
xnor U8973 (N_8973,N_8654,N_8675);
and U8974 (N_8974,N_8547,N_8669);
nand U8975 (N_8975,N_8598,N_8640);
nor U8976 (N_8976,N_8675,N_8552);
or U8977 (N_8977,N_8597,N_8670);
or U8978 (N_8978,N_8712,N_8740);
and U8979 (N_8979,N_8590,N_8746);
nor U8980 (N_8980,N_8730,N_8665);
and U8981 (N_8981,N_8531,N_8617);
and U8982 (N_8982,N_8522,N_8692);
and U8983 (N_8983,N_8704,N_8507);
xor U8984 (N_8984,N_8618,N_8532);
and U8985 (N_8985,N_8661,N_8584);
xor U8986 (N_8986,N_8537,N_8685);
xnor U8987 (N_8987,N_8648,N_8628);
nand U8988 (N_8988,N_8550,N_8703);
nand U8989 (N_8989,N_8519,N_8551);
xor U8990 (N_8990,N_8711,N_8715);
xor U8991 (N_8991,N_8664,N_8662);
or U8992 (N_8992,N_8521,N_8581);
nor U8993 (N_8993,N_8517,N_8623);
nor U8994 (N_8994,N_8558,N_8622);
and U8995 (N_8995,N_8681,N_8663);
xnor U8996 (N_8996,N_8534,N_8674);
nand U8997 (N_8997,N_8581,N_8540);
nand U8998 (N_8998,N_8525,N_8543);
nand U8999 (N_8999,N_8627,N_8664);
nor U9000 (N_9000,N_8983,N_8992);
and U9001 (N_9001,N_8990,N_8867);
nand U9002 (N_9002,N_8960,N_8920);
nor U9003 (N_9003,N_8945,N_8995);
nor U9004 (N_9004,N_8924,N_8833);
or U9005 (N_9005,N_8755,N_8810);
and U9006 (N_9006,N_8950,N_8851);
xnor U9007 (N_9007,N_8796,N_8793);
xnor U9008 (N_9008,N_8903,N_8963);
or U9009 (N_9009,N_8868,N_8962);
xor U9010 (N_9010,N_8877,N_8824);
nand U9011 (N_9011,N_8900,N_8958);
xor U9012 (N_9012,N_8979,N_8870);
xnor U9013 (N_9013,N_8993,N_8874);
nor U9014 (N_9014,N_8996,N_8754);
or U9015 (N_9015,N_8977,N_8803);
nor U9016 (N_9016,N_8927,N_8801);
or U9017 (N_9017,N_8842,N_8846);
nor U9018 (N_9018,N_8981,N_8914);
and U9019 (N_9019,N_8777,N_8951);
or U9020 (N_9020,N_8772,N_8885);
or U9021 (N_9021,N_8771,N_8837);
and U9022 (N_9022,N_8959,N_8802);
or U9023 (N_9023,N_8765,N_8858);
and U9024 (N_9024,N_8783,N_8843);
xnor U9025 (N_9025,N_8964,N_8999);
or U9026 (N_9026,N_8952,N_8826);
nand U9027 (N_9027,N_8781,N_8897);
xor U9028 (N_9028,N_8794,N_8967);
nand U9029 (N_9029,N_8855,N_8970);
xnor U9030 (N_9030,N_8789,N_8834);
or U9031 (N_9031,N_8982,N_8966);
xnor U9032 (N_9032,N_8938,N_8890);
nand U9033 (N_9033,N_8883,N_8998);
and U9034 (N_9034,N_8965,N_8812);
nand U9035 (N_9035,N_8814,N_8840);
xor U9036 (N_9036,N_8808,N_8784);
nand U9037 (N_9037,N_8969,N_8972);
nand U9038 (N_9038,N_8859,N_8813);
nand U9039 (N_9039,N_8854,N_8816);
nand U9040 (N_9040,N_8991,N_8929);
or U9041 (N_9041,N_8811,N_8778);
nor U9042 (N_9042,N_8844,N_8809);
or U9043 (N_9043,N_8880,N_8947);
nand U9044 (N_9044,N_8953,N_8864);
nand U9045 (N_9045,N_8861,N_8879);
and U9046 (N_9046,N_8909,N_8955);
or U9047 (N_9047,N_8762,N_8806);
xor U9048 (N_9048,N_8896,N_8946);
nor U9049 (N_9049,N_8761,N_8845);
xor U9050 (N_9050,N_8767,N_8876);
xnor U9051 (N_9051,N_8850,N_8984);
and U9052 (N_9052,N_8881,N_8912);
xor U9053 (N_9053,N_8830,N_8926);
xnor U9054 (N_9054,N_8799,N_8931);
and U9055 (N_9055,N_8974,N_8862);
and U9056 (N_9056,N_8863,N_8800);
xnor U9057 (N_9057,N_8935,N_8873);
nand U9058 (N_9058,N_8750,N_8886);
nand U9059 (N_9059,N_8857,N_8957);
nor U9060 (N_9060,N_8792,N_8988);
xor U9061 (N_9061,N_8758,N_8943);
nor U9062 (N_9062,N_8807,N_8928);
or U9063 (N_9063,N_8871,N_8847);
xor U9064 (N_9064,N_8889,N_8860);
or U9065 (N_9065,N_8875,N_8917);
and U9066 (N_9066,N_8786,N_8805);
nand U9067 (N_9067,N_8831,N_8911);
nand U9068 (N_9068,N_8753,N_8769);
or U9069 (N_9069,N_8756,N_8884);
and U9070 (N_9070,N_8825,N_8891);
and U9071 (N_9071,N_8828,N_8905);
nor U9072 (N_9072,N_8878,N_8848);
nor U9073 (N_9073,N_8785,N_8852);
nand U9074 (N_9074,N_8989,N_8898);
or U9075 (N_9075,N_8780,N_8866);
and U9076 (N_9076,N_8804,N_8934);
and U9077 (N_9077,N_8836,N_8894);
nor U9078 (N_9078,N_8788,N_8942);
and U9079 (N_9079,N_8978,N_8829);
nand U9080 (N_9080,N_8913,N_8770);
xor U9081 (N_9081,N_8779,N_8821);
xor U9082 (N_9082,N_8944,N_8930);
xor U9083 (N_9083,N_8768,N_8766);
or U9084 (N_9084,N_8752,N_8906);
nor U9085 (N_9085,N_8838,N_8902);
xor U9086 (N_9086,N_8976,N_8819);
nand U9087 (N_9087,N_8907,N_8910);
or U9088 (N_9088,N_8776,N_8835);
and U9089 (N_9089,N_8901,N_8787);
or U9090 (N_9090,N_8798,N_8791);
and U9091 (N_9091,N_8888,N_8773);
and U9092 (N_9092,N_8882,N_8908);
nor U9093 (N_9093,N_8940,N_8820);
nand U9094 (N_9094,N_8893,N_8763);
nor U9095 (N_9095,N_8887,N_8815);
nand U9096 (N_9096,N_8919,N_8975);
xor U9097 (N_9097,N_8818,N_8790);
or U9098 (N_9098,N_8980,N_8872);
and U9099 (N_9099,N_8823,N_8764);
nor U9100 (N_9100,N_8956,N_8941);
and U9101 (N_9101,N_8869,N_8922);
xnor U9102 (N_9102,N_8853,N_8892);
and U9103 (N_9103,N_8985,N_8915);
nor U9104 (N_9104,N_8827,N_8775);
nand U9105 (N_9105,N_8757,N_8817);
nand U9106 (N_9106,N_8895,N_8760);
xor U9107 (N_9107,N_8782,N_8971);
or U9108 (N_9108,N_8987,N_8936);
and U9109 (N_9109,N_8994,N_8797);
and U9110 (N_9110,N_8961,N_8923);
xnor U9111 (N_9111,N_8849,N_8997);
xnor U9112 (N_9112,N_8918,N_8973);
nor U9113 (N_9113,N_8759,N_8948);
or U9114 (N_9114,N_8856,N_8822);
or U9115 (N_9115,N_8774,N_8925);
and U9116 (N_9116,N_8841,N_8954);
nand U9117 (N_9117,N_8832,N_8921);
and U9118 (N_9118,N_8986,N_8939);
nand U9119 (N_9119,N_8932,N_8751);
or U9120 (N_9120,N_8933,N_8899);
or U9121 (N_9121,N_8968,N_8795);
or U9122 (N_9122,N_8916,N_8937);
xnor U9123 (N_9123,N_8865,N_8904);
xnor U9124 (N_9124,N_8949,N_8839);
and U9125 (N_9125,N_8944,N_8965);
or U9126 (N_9126,N_8789,N_8982);
nor U9127 (N_9127,N_8793,N_8862);
nand U9128 (N_9128,N_8865,N_8932);
xnor U9129 (N_9129,N_8879,N_8920);
nor U9130 (N_9130,N_8915,N_8758);
nor U9131 (N_9131,N_8871,N_8909);
nor U9132 (N_9132,N_8860,N_8847);
nor U9133 (N_9133,N_8851,N_8988);
nor U9134 (N_9134,N_8899,N_8800);
nand U9135 (N_9135,N_8938,N_8992);
xnor U9136 (N_9136,N_8966,N_8756);
and U9137 (N_9137,N_8786,N_8783);
and U9138 (N_9138,N_8783,N_8947);
xor U9139 (N_9139,N_8886,N_8910);
nor U9140 (N_9140,N_8834,N_8767);
or U9141 (N_9141,N_8904,N_8910);
or U9142 (N_9142,N_8943,N_8777);
or U9143 (N_9143,N_8758,N_8870);
or U9144 (N_9144,N_8789,N_8866);
nand U9145 (N_9145,N_8937,N_8763);
or U9146 (N_9146,N_8981,N_8940);
xnor U9147 (N_9147,N_8774,N_8988);
or U9148 (N_9148,N_8979,N_8763);
nand U9149 (N_9149,N_8915,N_8954);
xnor U9150 (N_9150,N_8812,N_8842);
xor U9151 (N_9151,N_8753,N_8877);
nor U9152 (N_9152,N_8879,N_8944);
or U9153 (N_9153,N_8876,N_8932);
or U9154 (N_9154,N_8842,N_8930);
nor U9155 (N_9155,N_8995,N_8946);
xor U9156 (N_9156,N_8870,N_8905);
nor U9157 (N_9157,N_8867,N_8971);
or U9158 (N_9158,N_8981,N_8876);
and U9159 (N_9159,N_8798,N_8829);
nand U9160 (N_9160,N_8869,N_8954);
or U9161 (N_9161,N_8868,N_8955);
or U9162 (N_9162,N_8918,N_8877);
or U9163 (N_9163,N_8833,N_8789);
nor U9164 (N_9164,N_8757,N_8953);
nor U9165 (N_9165,N_8925,N_8987);
nor U9166 (N_9166,N_8987,N_8826);
xnor U9167 (N_9167,N_8868,N_8844);
nor U9168 (N_9168,N_8761,N_8835);
and U9169 (N_9169,N_8838,N_8829);
xnor U9170 (N_9170,N_8759,N_8784);
nand U9171 (N_9171,N_8911,N_8984);
and U9172 (N_9172,N_8846,N_8790);
and U9173 (N_9173,N_8926,N_8958);
and U9174 (N_9174,N_8983,N_8906);
nand U9175 (N_9175,N_8958,N_8876);
nor U9176 (N_9176,N_8826,N_8834);
or U9177 (N_9177,N_8763,N_8790);
nand U9178 (N_9178,N_8960,N_8783);
nor U9179 (N_9179,N_8959,N_8985);
and U9180 (N_9180,N_8815,N_8762);
or U9181 (N_9181,N_8898,N_8964);
xnor U9182 (N_9182,N_8826,N_8785);
xnor U9183 (N_9183,N_8844,N_8848);
nand U9184 (N_9184,N_8841,N_8816);
or U9185 (N_9185,N_8751,N_8778);
nand U9186 (N_9186,N_8829,N_8750);
xnor U9187 (N_9187,N_8836,N_8819);
nor U9188 (N_9188,N_8844,N_8907);
nor U9189 (N_9189,N_8763,N_8809);
and U9190 (N_9190,N_8828,N_8795);
xnor U9191 (N_9191,N_8774,N_8969);
nor U9192 (N_9192,N_8853,N_8760);
nand U9193 (N_9193,N_8837,N_8805);
nand U9194 (N_9194,N_8764,N_8966);
and U9195 (N_9195,N_8787,N_8844);
and U9196 (N_9196,N_8826,N_8983);
and U9197 (N_9197,N_8913,N_8938);
nor U9198 (N_9198,N_8875,N_8784);
nor U9199 (N_9199,N_8905,N_8802);
nor U9200 (N_9200,N_8755,N_8986);
or U9201 (N_9201,N_8943,N_8754);
xnor U9202 (N_9202,N_8752,N_8807);
xnor U9203 (N_9203,N_8808,N_8934);
and U9204 (N_9204,N_8853,N_8756);
xor U9205 (N_9205,N_8853,N_8944);
nand U9206 (N_9206,N_8865,N_8908);
xor U9207 (N_9207,N_8983,N_8942);
xor U9208 (N_9208,N_8994,N_8990);
and U9209 (N_9209,N_8913,N_8999);
and U9210 (N_9210,N_8841,N_8753);
and U9211 (N_9211,N_8930,N_8991);
and U9212 (N_9212,N_8837,N_8758);
xor U9213 (N_9213,N_8849,N_8833);
or U9214 (N_9214,N_8958,N_8850);
xnor U9215 (N_9215,N_8866,N_8972);
xor U9216 (N_9216,N_8959,N_8813);
or U9217 (N_9217,N_8772,N_8974);
nand U9218 (N_9218,N_8888,N_8994);
and U9219 (N_9219,N_8822,N_8937);
or U9220 (N_9220,N_8909,N_8770);
nor U9221 (N_9221,N_8960,N_8814);
xnor U9222 (N_9222,N_8795,N_8831);
or U9223 (N_9223,N_8898,N_8965);
and U9224 (N_9224,N_8978,N_8876);
and U9225 (N_9225,N_8756,N_8796);
nand U9226 (N_9226,N_8957,N_8928);
and U9227 (N_9227,N_8824,N_8832);
nor U9228 (N_9228,N_8759,N_8952);
nand U9229 (N_9229,N_8833,N_8854);
nand U9230 (N_9230,N_8894,N_8912);
nand U9231 (N_9231,N_8956,N_8951);
nor U9232 (N_9232,N_8777,N_8938);
and U9233 (N_9233,N_8839,N_8752);
and U9234 (N_9234,N_8790,N_8816);
nand U9235 (N_9235,N_8862,N_8780);
nand U9236 (N_9236,N_8823,N_8803);
nand U9237 (N_9237,N_8906,N_8886);
and U9238 (N_9238,N_8904,N_8971);
or U9239 (N_9239,N_8763,N_8915);
or U9240 (N_9240,N_8793,N_8752);
nand U9241 (N_9241,N_8843,N_8908);
and U9242 (N_9242,N_8823,N_8872);
and U9243 (N_9243,N_8890,N_8919);
nor U9244 (N_9244,N_8795,N_8816);
nor U9245 (N_9245,N_8750,N_8802);
nor U9246 (N_9246,N_8872,N_8771);
nor U9247 (N_9247,N_8870,N_8819);
or U9248 (N_9248,N_8926,N_8891);
or U9249 (N_9249,N_8956,N_8937);
and U9250 (N_9250,N_9075,N_9135);
nor U9251 (N_9251,N_9206,N_9040);
or U9252 (N_9252,N_9172,N_9108);
xor U9253 (N_9253,N_9017,N_9195);
nor U9254 (N_9254,N_9177,N_9006);
xor U9255 (N_9255,N_9005,N_9096);
nor U9256 (N_9256,N_9104,N_9071);
or U9257 (N_9257,N_9154,N_9129);
xor U9258 (N_9258,N_9015,N_9150);
nor U9259 (N_9259,N_9182,N_9122);
or U9260 (N_9260,N_9180,N_9078);
and U9261 (N_9261,N_9019,N_9086);
nand U9262 (N_9262,N_9033,N_9021);
nand U9263 (N_9263,N_9160,N_9205);
nor U9264 (N_9264,N_9249,N_9197);
nor U9265 (N_9265,N_9179,N_9046);
xor U9266 (N_9266,N_9109,N_9052);
or U9267 (N_9267,N_9063,N_9087);
or U9268 (N_9268,N_9065,N_9169);
xor U9269 (N_9269,N_9213,N_9094);
or U9270 (N_9270,N_9217,N_9143);
nor U9271 (N_9271,N_9224,N_9051);
nand U9272 (N_9272,N_9147,N_9208);
nor U9273 (N_9273,N_9142,N_9126);
nand U9274 (N_9274,N_9089,N_9191);
or U9275 (N_9275,N_9153,N_9115);
xnor U9276 (N_9276,N_9136,N_9041);
nor U9277 (N_9277,N_9207,N_9002);
xnor U9278 (N_9278,N_9022,N_9238);
nand U9279 (N_9279,N_9060,N_9219);
nor U9280 (N_9280,N_9001,N_9134);
or U9281 (N_9281,N_9114,N_9008);
or U9282 (N_9282,N_9027,N_9178);
nor U9283 (N_9283,N_9010,N_9231);
and U9284 (N_9284,N_9175,N_9042);
nor U9285 (N_9285,N_9121,N_9050);
xor U9286 (N_9286,N_9196,N_9165);
xnor U9287 (N_9287,N_9088,N_9192);
and U9288 (N_9288,N_9045,N_9083);
nor U9289 (N_9289,N_9139,N_9116);
xor U9290 (N_9290,N_9221,N_9029);
and U9291 (N_9291,N_9112,N_9059);
or U9292 (N_9292,N_9119,N_9186);
and U9293 (N_9293,N_9157,N_9111);
or U9294 (N_9294,N_9009,N_9113);
or U9295 (N_9295,N_9039,N_9176);
nand U9296 (N_9296,N_9241,N_9077);
nand U9297 (N_9297,N_9144,N_9064);
xnor U9298 (N_9298,N_9235,N_9082);
xor U9299 (N_9299,N_9018,N_9090);
xnor U9300 (N_9300,N_9181,N_9067);
or U9301 (N_9301,N_9093,N_9124);
nor U9302 (N_9302,N_9034,N_9014);
nor U9303 (N_9303,N_9068,N_9201);
nand U9304 (N_9304,N_9155,N_9056);
nand U9305 (N_9305,N_9185,N_9161);
or U9306 (N_9306,N_9247,N_9248);
xor U9307 (N_9307,N_9228,N_9012);
or U9308 (N_9308,N_9100,N_9053);
nand U9309 (N_9309,N_9245,N_9101);
nor U9310 (N_9310,N_9007,N_9003);
or U9311 (N_9311,N_9133,N_9037);
and U9312 (N_9312,N_9092,N_9174);
or U9313 (N_9313,N_9229,N_9233);
or U9314 (N_9314,N_9216,N_9237);
nand U9315 (N_9315,N_9081,N_9117);
nand U9316 (N_9316,N_9159,N_9049);
xnor U9317 (N_9317,N_9244,N_9130);
nor U9318 (N_9318,N_9211,N_9242);
nand U9319 (N_9319,N_9025,N_9234);
xnor U9320 (N_9320,N_9200,N_9011);
and U9321 (N_9321,N_9079,N_9098);
and U9322 (N_9322,N_9204,N_9225);
xnor U9323 (N_9323,N_9183,N_9152);
nand U9324 (N_9324,N_9163,N_9214);
and U9325 (N_9325,N_9223,N_9031);
or U9326 (N_9326,N_9054,N_9120);
and U9327 (N_9327,N_9032,N_9230);
xnor U9328 (N_9328,N_9199,N_9057);
or U9329 (N_9329,N_9105,N_9131);
xor U9330 (N_9330,N_9220,N_9158);
and U9331 (N_9331,N_9103,N_9106);
or U9332 (N_9332,N_9194,N_9069);
and U9333 (N_9333,N_9023,N_9187);
nand U9334 (N_9334,N_9190,N_9074);
nand U9335 (N_9335,N_9102,N_9125);
nand U9336 (N_9336,N_9202,N_9149);
nor U9337 (N_9337,N_9128,N_9212);
or U9338 (N_9338,N_9210,N_9170);
nand U9339 (N_9339,N_9222,N_9076);
and U9340 (N_9340,N_9073,N_9091);
nor U9341 (N_9341,N_9061,N_9198);
xnor U9342 (N_9342,N_9004,N_9123);
or U9343 (N_9343,N_9099,N_9141);
nand U9344 (N_9344,N_9156,N_9028);
nor U9345 (N_9345,N_9189,N_9132);
nand U9346 (N_9346,N_9066,N_9193);
nor U9347 (N_9347,N_9227,N_9140);
nand U9348 (N_9348,N_9151,N_9110);
xnor U9349 (N_9349,N_9166,N_9055);
and U9350 (N_9350,N_9173,N_9226);
nand U9351 (N_9351,N_9072,N_9145);
nor U9352 (N_9352,N_9013,N_9026);
xor U9353 (N_9353,N_9162,N_9168);
xor U9354 (N_9354,N_9171,N_9240);
xor U9355 (N_9355,N_9215,N_9062);
nand U9356 (N_9356,N_9038,N_9164);
nor U9357 (N_9357,N_9030,N_9203);
and U9358 (N_9358,N_9035,N_9107);
or U9359 (N_9359,N_9044,N_9218);
nor U9360 (N_9360,N_9118,N_9232);
and U9361 (N_9361,N_9167,N_9048);
and U9362 (N_9362,N_9016,N_9239);
nor U9363 (N_9363,N_9127,N_9137);
nand U9364 (N_9364,N_9070,N_9184);
nor U9365 (N_9365,N_9243,N_9024);
nor U9366 (N_9366,N_9188,N_9036);
nand U9367 (N_9367,N_9043,N_9097);
xnor U9368 (N_9368,N_9080,N_9058);
xnor U9369 (N_9369,N_9209,N_9000);
nand U9370 (N_9370,N_9138,N_9047);
or U9371 (N_9371,N_9020,N_9095);
and U9372 (N_9372,N_9236,N_9084);
nor U9373 (N_9373,N_9148,N_9246);
nor U9374 (N_9374,N_9146,N_9085);
nand U9375 (N_9375,N_9046,N_9094);
xnor U9376 (N_9376,N_9231,N_9031);
xnor U9377 (N_9377,N_9035,N_9197);
and U9378 (N_9378,N_9133,N_9188);
and U9379 (N_9379,N_9140,N_9186);
nor U9380 (N_9380,N_9018,N_9216);
xor U9381 (N_9381,N_9096,N_9236);
nand U9382 (N_9382,N_9018,N_9244);
or U9383 (N_9383,N_9028,N_9138);
nor U9384 (N_9384,N_9209,N_9135);
nor U9385 (N_9385,N_9009,N_9172);
or U9386 (N_9386,N_9143,N_9141);
or U9387 (N_9387,N_9090,N_9188);
nand U9388 (N_9388,N_9055,N_9087);
nand U9389 (N_9389,N_9015,N_9012);
and U9390 (N_9390,N_9229,N_9161);
nor U9391 (N_9391,N_9202,N_9012);
xor U9392 (N_9392,N_9121,N_9033);
nor U9393 (N_9393,N_9100,N_9156);
and U9394 (N_9394,N_9125,N_9134);
and U9395 (N_9395,N_9017,N_9033);
xor U9396 (N_9396,N_9054,N_9147);
nor U9397 (N_9397,N_9190,N_9216);
or U9398 (N_9398,N_9123,N_9233);
xor U9399 (N_9399,N_9012,N_9077);
xnor U9400 (N_9400,N_9112,N_9142);
xnor U9401 (N_9401,N_9068,N_9049);
or U9402 (N_9402,N_9128,N_9073);
nor U9403 (N_9403,N_9044,N_9192);
xor U9404 (N_9404,N_9147,N_9101);
nand U9405 (N_9405,N_9055,N_9132);
nand U9406 (N_9406,N_9119,N_9192);
and U9407 (N_9407,N_9141,N_9144);
nor U9408 (N_9408,N_9210,N_9202);
nor U9409 (N_9409,N_9031,N_9083);
nor U9410 (N_9410,N_9113,N_9124);
or U9411 (N_9411,N_9103,N_9158);
nor U9412 (N_9412,N_9041,N_9240);
nand U9413 (N_9413,N_9144,N_9051);
nor U9414 (N_9414,N_9035,N_9154);
xor U9415 (N_9415,N_9041,N_9026);
nand U9416 (N_9416,N_9035,N_9215);
and U9417 (N_9417,N_9013,N_9229);
nand U9418 (N_9418,N_9179,N_9198);
nor U9419 (N_9419,N_9003,N_9061);
and U9420 (N_9420,N_9026,N_9174);
nand U9421 (N_9421,N_9026,N_9082);
nor U9422 (N_9422,N_9239,N_9172);
nand U9423 (N_9423,N_9198,N_9087);
xor U9424 (N_9424,N_9205,N_9210);
nor U9425 (N_9425,N_9180,N_9214);
and U9426 (N_9426,N_9004,N_9059);
nand U9427 (N_9427,N_9101,N_9081);
and U9428 (N_9428,N_9147,N_9034);
nor U9429 (N_9429,N_9239,N_9027);
or U9430 (N_9430,N_9095,N_9087);
nand U9431 (N_9431,N_9247,N_9098);
xnor U9432 (N_9432,N_9123,N_9141);
xor U9433 (N_9433,N_9089,N_9026);
or U9434 (N_9434,N_9238,N_9027);
or U9435 (N_9435,N_9145,N_9243);
xnor U9436 (N_9436,N_9206,N_9118);
nor U9437 (N_9437,N_9179,N_9139);
and U9438 (N_9438,N_9204,N_9205);
xnor U9439 (N_9439,N_9068,N_9142);
and U9440 (N_9440,N_9101,N_9076);
or U9441 (N_9441,N_9220,N_9029);
xnor U9442 (N_9442,N_9117,N_9126);
and U9443 (N_9443,N_9135,N_9098);
nand U9444 (N_9444,N_9196,N_9092);
xnor U9445 (N_9445,N_9088,N_9209);
and U9446 (N_9446,N_9179,N_9186);
xnor U9447 (N_9447,N_9210,N_9045);
xnor U9448 (N_9448,N_9112,N_9076);
nor U9449 (N_9449,N_9221,N_9036);
nor U9450 (N_9450,N_9037,N_9025);
nor U9451 (N_9451,N_9104,N_9208);
nand U9452 (N_9452,N_9013,N_9214);
nand U9453 (N_9453,N_9098,N_9000);
and U9454 (N_9454,N_9178,N_9028);
nor U9455 (N_9455,N_9160,N_9213);
nor U9456 (N_9456,N_9041,N_9161);
nor U9457 (N_9457,N_9223,N_9113);
nand U9458 (N_9458,N_9210,N_9133);
and U9459 (N_9459,N_9013,N_9003);
or U9460 (N_9460,N_9011,N_9091);
nand U9461 (N_9461,N_9230,N_9029);
and U9462 (N_9462,N_9196,N_9086);
nand U9463 (N_9463,N_9236,N_9247);
or U9464 (N_9464,N_9046,N_9089);
nand U9465 (N_9465,N_9030,N_9235);
nor U9466 (N_9466,N_9207,N_9087);
nand U9467 (N_9467,N_9147,N_9111);
and U9468 (N_9468,N_9172,N_9039);
xor U9469 (N_9469,N_9115,N_9139);
and U9470 (N_9470,N_9141,N_9238);
xnor U9471 (N_9471,N_9070,N_9195);
nand U9472 (N_9472,N_9120,N_9214);
nand U9473 (N_9473,N_9128,N_9090);
and U9474 (N_9474,N_9118,N_9237);
xor U9475 (N_9475,N_9054,N_9041);
xor U9476 (N_9476,N_9214,N_9109);
nand U9477 (N_9477,N_9241,N_9200);
nor U9478 (N_9478,N_9073,N_9044);
nand U9479 (N_9479,N_9047,N_9235);
xor U9480 (N_9480,N_9154,N_9234);
xnor U9481 (N_9481,N_9109,N_9105);
or U9482 (N_9482,N_9015,N_9116);
nor U9483 (N_9483,N_9197,N_9202);
xnor U9484 (N_9484,N_9089,N_9238);
xor U9485 (N_9485,N_9150,N_9215);
or U9486 (N_9486,N_9112,N_9099);
xnor U9487 (N_9487,N_9238,N_9234);
and U9488 (N_9488,N_9144,N_9242);
or U9489 (N_9489,N_9135,N_9114);
or U9490 (N_9490,N_9093,N_9164);
nor U9491 (N_9491,N_9105,N_9145);
and U9492 (N_9492,N_9208,N_9049);
xor U9493 (N_9493,N_9042,N_9047);
and U9494 (N_9494,N_9185,N_9123);
or U9495 (N_9495,N_9172,N_9138);
nand U9496 (N_9496,N_9199,N_9105);
nand U9497 (N_9497,N_9140,N_9081);
or U9498 (N_9498,N_9081,N_9130);
nor U9499 (N_9499,N_9237,N_9012);
xnor U9500 (N_9500,N_9427,N_9373);
and U9501 (N_9501,N_9393,N_9388);
or U9502 (N_9502,N_9443,N_9434);
nand U9503 (N_9503,N_9403,N_9347);
nor U9504 (N_9504,N_9317,N_9288);
and U9505 (N_9505,N_9266,N_9284);
or U9506 (N_9506,N_9265,N_9474);
nor U9507 (N_9507,N_9457,N_9310);
nor U9508 (N_9508,N_9428,N_9290);
nand U9509 (N_9509,N_9422,N_9256);
or U9510 (N_9510,N_9279,N_9329);
and U9511 (N_9511,N_9442,N_9400);
or U9512 (N_9512,N_9326,N_9351);
and U9513 (N_9513,N_9311,N_9405);
nor U9514 (N_9514,N_9287,N_9409);
xnor U9515 (N_9515,N_9435,N_9260);
or U9516 (N_9516,N_9466,N_9447);
nor U9517 (N_9517,N_9352,N_9426);
or U9518 (N_9518,N_9370,N_9316);
and U9519 (N_9519,N_9490,N_9470);
or U9520 (N_9520,N_9360,N_9268);
nand U9521 (N_9521,N_9449,N_9345);
nor U9522 (N_9522,N_9451,N_9424);
xor U9523 (N_9523,N_9332,N_9395);
nand U9524 (N_9524,N_9492,N_9301);
nand U9525 (N_9525,N_9253,N_9385);
nor U9526 (N_9526,N_9419,N_9402);
nor U9527 (N_9527,N_9357,N_9349);
xor U9528 (N_9528,N_9408,N_9483);
xor U9529 (N_9529,N_9366,N_9344);
or U9530 (N_9530,N_9448,N_9396);
nand U9531 (N_9531,N_9341,N_9337);
and U9532 (N_9532,N_9421,N_9312);
nor U9533 (N_9533,N_9465,N_9420);
or U9534 (N_9534,N_9440,N_9336);
nor U9535 (N_9535,N_9369,N_9304);
xor U9536 (N_9536,N_9278,N_9382);
xor U9537 (N_9537,N_9392,N_9418);
or U9538 (N_9538,N_9487,N_9273);
and U9539 (N_9539,N_9425,N_9378);
or U9540 (N_9540,N_9376,N_9295);
xnor U9541 (N_9541,N_9452,N_9323);
nor U9542 (N_9542,N_9251,N_9348);
or U9543 (N_9543,N_9404,N_9499);
nand U9544 (N_9544,N_9327,N_9430);
nor U9545 (N_9545,N_9309,N_9258);
nor U9546 (N_9546,N_9328,N_9495);
nand U9547 (N_9547,N_9263,N_9432);
nand U9548 (N_9548,N_9371,N_9441);
nor U9549 (N_9549,N_9285,N_9321);
or U9550 (N_9550,N_9383,N_9281);
or U9551 (N_9551,N_9485,N_9335);
and U9552 (N_9552,N_9294,N_9350);
nand U9553 (N_9553,N_9267,N_9363);
and U9554 (N_9554,N_9491,N_9429);
or U9555 (N_9555,N_9439,N_9386);
nand U9556 (N_9556,N_9473,N_9379);
xor U9557 (N_9557,N_9380,N_9413);
nor U9558 (N_9558,N_9291,N_9325);
and U9559 (N_9559,N_9320,N_9445);
nor U9560 (N_9560,N_9356,N_9459);
or U9561 (N_9561,N_9488,N_9282);
and U9562 (N_9562,N_9334,N_9368);
xnor U9563 (N_9563,N_9384,N_9272);
xnor U9564 (N_9564,N_9468,N_9481);
nor U9565 (N_9565,N_9477,N_9455);
and U9566 (N_9566,N_9478,N_9333);
or U9567 (N_9567,N_9330,N_9374);
nor U9568 (N_9568,N_9387,N_9472);
nand U9569 (N_9569,N_9493,N_9444);
or U9570 (N_9570,N_9375,N_9277);
nor U9571 (N_9571,N_9314,N_9324);
nand U9572 (N_9572,N_9359,N_9461);
nand U9573 (N_9573,N_9464,N_9437);
nand U9574 (N_9574,N_9283,N_9342);
xnor U9575 (N_9575,N_9399,N_9364);
or U9576 (N_9576,N_9254,N_9343);
nor U9577 (N_9577,N_9391,N_9454);
and U9578 (N_9578,N_9299,N_9257);
nand U9579 (N_9579,N_9262,N_9486);
and U9580 (N_9580,N_9471,N_9496);
xor U9581 (N_9581,N_9431,N_9479);
nand U9582 (N_9582,N_9264,N_9372);
nand U9583 (N_9583,N_9458,N_9280);
and U9584 (N_9584,N_9308,N_9469);
nand U9585 (N_9585,N_9367,N_9398);
nor U9586 (N_9586,N_9293,N_9340);
nand U9587 (N_9587,N_9410,N_9423);
nand U9588 (N_9588,N_9302,N_9298);
or U9589 (N_9589,N_9433,N_9275);
or U9590 (N_9590,N_9286,N_9497);
xor U9591 (N_9591,N_9353,N_9484);
and U9592 (N_9592,N_9255,N_9307);
nor U9593 (N_9593,N_9460,N_9259);
and U9594 (N_9594,N_9463,N_9494);
xor U9595 (N_9595,N_9456,N_9338);
and U9596 (N_9596,N_9475,N_9498);
nand U9597 (N_9597,N_9489,N_9306);
nor U9598 (N_9598,N_9361,N_9358);
and U9599 (N_9599,N_9397,N_9406);
or U9600 (N_9600,N_9271,N_9354);
and U9601 (N_9601,N_9365,N_9303);
and U9602 (N_9602,N_9453,N_9377);
xor U9603 (N_9603,N_9407,N_9482);
xor U9604 (N_9604,N_9417,N_9296);
or U9605 (N_9605,N_9252,N_9476);
nand U9606 (N_9606,N_9274,N_9346);
xor U9607 (N_9607,N_9480,N_9305);
or U9608 (N_9608,N_9355,N_9319);
or U9609 (N_9609,N_9446,N_9300);
nand U9610 (N_9610,N_9462,N_9438);
xnor U9611 (N_9611,N_9416,N_9401);
or U9612 (N_9612,N_9276,N_9269);
nand U9613 (N_9613,N_9331,N_9362);
nor U9614 (N_9614,N_9412,N_9389);
xor U9615 (N_9615,N_9322,N_9381);
nand U9616 (N_9616,N_9411,N_9339);
nor U9617 (N_9617,N_9318,N_9297);
xor U9618 (N_9618,N_9436,N_9270);
nor U9619 (N_9619,N_9467,N_9289);
nor U9620 (N_9620,N_9390,N_9292);
and U9621 (N_9621,N_9250,N_9414);
or U9622 (N_9622,N_9394,N_9261);
nand U9623 (N_9623,N_9313,N_9315);
nand U9624 (N_9624,N_9450,N_9415);
and U9625 (N_9625,N_9355,N_9371);
nand U9626 (N_9626,N_9364,N_9314);
or U9627 (N_9627,N_9448,N_9390);
nor U9628 (N_9628,N_9354,N_9322);
nand U9629 (N_9629,N_9381,N_9353);
xnor U9630 (N_9630,N_9495,N_9364);
nand U9631 (N_9631,N_9422,N_9349);
xnor U9632 (N_9632,N_9289,N_9293);
nand U9633 (N_9633,N_9444,N_9299);
nor U9634 (N_9634,N_9396,N_9466);
nor U9635 (N_9635,N_9499,N_9353);
nand U9636 (N_9636,N_9478,N_9309);
nor U9637 (N_9637,N_9480,N_9434);
or U9638 (N_9638,N_9350,N_9462);
nor U9639 (N_9639,N_9260,N_9371);
and U9640 (N_9640,N_9314,N_9290);
nor U9641 (N_9641,N_9384,N_9474);
or U9642 (N_9642,N_9433,N_9415);
nand U9643 (N_9643,N_9412,N_9479);
nor U9644 (N_9644,N_9258,N_9316);
and U9645 (N_9645,N_9433,N_9405);
and U9646 (N_9646,N_9251,N_9424);
and U9647 (N_9647,N_9283,N_9335);
or U9648 (N_9648,N_9384,N_9381);
nor U9649 (N_9649,N_9334,N_9296);
or U9650 (N_9650,N_9290,N_9355);
or U9651 (N_9651,N_9306,N_9380);
xor U9652 (N_9652,N_9370,N_9426);
nor U9653 (N_9653,N_9429,N_9350);
and U9654 (N_9654,N_9390,N_9356);
xnor U9655 (N_9655,N_9427,N_9483);
nor U9656 (N_9656,N_9279,N_9377);
or U9657 (N_9657,N_9421,N_9387);
xnor U9658 (N_9658,N_9438,N_9419);
nor U9659 (N_9659,N_9319,N_9264);
nor U9660 (N_9660,N_9321,N_9354);
nor U9661 (N_9661,N_9384,N_9411);
nand U9662 (N_9662,N_9368,N_9476);
or U9663 (N_9663,N_9464,N_9286);
or U9664 (N_9664,N_9420,N_9283);
xor U9665 (N_9665,N_9494,N_9323);
and U9666 (N_9666,N_9406,N_9474);
or U9667 (N_9667,N_9323,N_9356);
nand U9668 (N_9668,N_9434,N_9369);
nand U9669 (N_9669,N_9462,N_9277);
nor U9670 (N_9670,N_9381,N_9461);
xnor U9671 (N_9671,N_9415,N_9280);
and U9672 (N_9672,N_9416,N_9351);
and U9673 (N_9673,N_9397,N_9334);
xnor U9674 (N_9674,N_9258,N_9394);
nor U9675 (N_9675,N_9409,N_9474);
or U9676 (N_9676,N_9297,N_9345);
nand U9677 (N_9677,N_9375,N_9425);
xor U9678 (N_9678,N_9373,N_9417);
or U9679 (N_9679,N_9256,N_9303);
nand U9680 (N_9680,N_9362,N_9282);
and U9681 (N_9681,N_9419,N_9479);
nand U9682 (N_9682,N_9475,N_9458);
or U9683 (N_9683,N_9375,N_9272);
or U9684 (N_9684,N_9468,N_9463);
nand U9685 (N_9685,N_9289,N_9341);
and U9686 (N_9686,N_9413,N_9323);
or U9687 (N_9687,N_9262,N_9348);
nor U9688 (N_9688,N_9490,N_9419);
xnor U9689 (N_9689,N_9309,N_9405);
nor U9690 (N_9690,N_9463,N_9385);
and U9691 (N_9691,N_9250,N_9491);
nor U9692 (N_9692,N_9394,N_9458);
or U9693 (N_9693,N_9391,N_9422);
or U9694 (N_9694,N_9498,N_9389);
or U9695 (N_9695,N_9393,N_9497);
nor U9696 (N_9696,N_9259,N_9436);
nor U9697 (N_9697,N_9318,N_9361);
xnor U9698 (N_9698,N_9391,N_9337);
or U9699 (N_9699,N_9438,N_9333);
or U9700 (N_9700,N_9261,N_9389);
nand U9701 (N_9701,N_9260,N_9483);
and U9702 (N_9702,N_9414,N_9467);
or U9703 (N_9703,N_9489,N_9410);
or U9704 (N_9704,N_9334,N_9376);
and U9705 (N_9705,N_9465,N_9498);
nand U9706 (N_9706,N_9335,N_9339);
xor U9707 (N_9707,N_9305,N_9280);
nor U9708 (N_9708,N_9434,N_9292);
and U9709 (N_9709,N_9472,N_9473);
nand U9710 (N_9710,N_9304,N_9372);
nor U9711 (N_9711,N_9287,N_9403);
nand U9712 (N_9712,N_9414,N_9452);
and U9713 (N_9713,N_9493,N_9335);
or U9714 (N_9714,N_9425,N_9322);
xnor U9715 (N_9715,N_9334,N_9250);
nand U9716 (N_9716,N_9495,N_9482);
and U9717 (N_9717,N_9472,N_9363);
nand U9718 (N_9718,N_9409,N_9272);
or U9719 (N_9719,N_9353,N_9327);
xor U9720 (N_9720,N_9488,N_9375);
xor U9721 (N_9721,N_9261,N_9420);
nand U9722 (N_9722,N_9395,N_9380);
xor U9723 (N_9723,N_9363,N_9261);
nand U9724 (N_9724,N_9419,N_9272);
nand U9725 (N_9725,N_9282,N_9442);
xor U9726 (N_9726,N_9466,N_9287);
nor U9727 (N_9727,N_9316,N_9430);
nand U9728 (N_9728,N_9407,N_9295);
nand U9729 (N_9729,N_9271,N_9407);
and U9730 (N_9730,N_9313,N_9480);
and U9731 (N_9731,N_9422,N_9469);
nand U9732 (N_9732,N_9309,N_9414);
nor U9733 (N_9733,N_9357,N_9398);
and U9734 (N_9734,N_9314,N_9335);
xor U9735 (N_9735,N_9353,N_9431);
or U9736 (N_9736,N_9466,N_9329);
xnor U9737 (N_9737,N_9320,N_9489);
nor U9738 (N_9738,N_9305,N_9370);
nand U9739 (N_9739,N_9259,N_9320);
or U9740 (N_9740,N_9415,N_9328);
xnor U9741 (N_9741,N_9278,N_9338);
xnor U9742 (N_9742,N_9454,N_9430);
nand U9743 (N_9743,N_9282,N_9452);
and U9744 (N_9744,N_9425,N_9380);
or U9745 (N_9745,N_9423,N_9300);
nor U9746 (N_9746,N_9402,N_9413);
and U9747 (N_9747,N_9260,N_9294);
and U9748 (N_9748,N_9476,N_9393);
nand U9749 (N_9749,N_9432,N_9408);
nor U9750 (N_9750,N_9707,N_9574);
or U9751 (N_9751,N_9500,N_9665);
and U9752 (N_9752,N_9663,N_9542);
and U9753 (N_9753,N_9531,N_9738);
xnor U9754 (N_9754,N_9695,N_9546);
nor U9755 (N_9755,N_9632,N_9643);
xor U9756 (N_9756,N_9527,N_9514);
nand U9757 (N_9757,N_9691,N_9701);
xor U9758 (N_9758,N_9521,N_9660);
nand U9759 (N_9759,N_9645,N_9712);
nor U9760 (N_9760,N_9705,N_9621);
xor U9761 (N_9761,N_9749,N_9746);
or U9762 (N_9762,N_9614,N_9561);
nand U9763 (N_9763,N_9572,N_9680);
and U9764 (N_9764,N_9704,N_9578);
xor U9765 (N_9765,N_9615,N_9657);
xor U9766 (N_9766,N_9727,N_9523);
nor U9767 (N_9767,N_9510,N_9536);
and U9768 (N_9768,N_9553,N_9573);
nor U9769 (N_9769,N_9594,N_9736);
xor U9770 (N_9770,N_9700,N_9675);
nand U9771 (N_9771,N_9501,N_9575);
xnor U9772 (N_9772,N_9601,N_9733);
xor U9773 (N_9773,N_9607,N_9549);
or U9774 (N_9774,N_9728,N_9697);
nand U9775 (N_9775,N_9563,N_9658);
and U9776 (N_9776,N_9509,N_9581);
and U9777 (N_9777,N_9731,N_9659);
xnor U9778 (N_9778,N_9630,N_9584);
xnor U9779 (N_9779,N_9653,N_9708);
and U9780 (N_9780,N_9720,N_9623);
nor U9781 (N_9781,N_9566,N_9638);
and U9782 (N_9782,N_9714,N_9613);
xnor U9783 (N_9783,N_9689,N_9532);
and U9784 (N_9784,N_9508,N_9652);
or U9785 (N_9785,N_9577,N_9582);
nand U9786 (N_9786,N_9503,N_9661);
and U9787 (N_9787,N_9620,N_9543);
nor U9788 (N_9788,N_9526,N_9669);
xnor U9789 (N_9789,N_9539,N_9569);
nor U9790 (N_9790,N_9622,N_9648);
nand U9791 (N_9791,N_9512,N_9502);
nor U9792 (N_9792,N_9522,N_9627);
or U9793 (N_9793,N_9525,N_9618);
nor U9794 (N_9794,N_9692,N_9595);
or U9795 (N_9795,N_9541,N_9505);
nor U9796 (N_9796,N_9589,N_9585);
nor U9797 (N_9797,N_9676,N_9694);
nor U9798 (N_9798,N_9626,N_9698);
xnor U9799 (N_9799,N_9625,N_9646);
nand U9800 (N_9800,N_9565,N_9555);
nand U9801 (N_9801,N_9716,N_9504);
nor U9802 (N_9802,N_9709,N_9586);
and U9803 (N_9803,N_9723,N_9507);
nor U9804 (N_9804,N_9557,N_9511);
nand U9805 (N_9805,N_9516,N_9706);
nor U9806 (N_9806,N_9672,N_9591);
or U9807 (N_9807,N_9741,N_9673);
xor U9808 (N_9808,N_9711,N_9662);
or U9809 (N_9809,N_9664,N_9679);
nor U9810 (N_9810,N_9730,N_9671);
and U9811 (N_9811,N_9593,N_9550);
nor U9812 (N_9812,N_9740,N_9559);
nor U9813 (N_9813,N_9560,N_9538);
nor U9814 (N_9814,N_9629,N_9693);
nand U9815 (N_9815,N_9725,N_9631);
nand U9816 (N_9816,N_9639,N_9609);
nor U9817 (N_9817,N_9656,N_9592);
or U9818 (N_9818,N_9722,N_9544);
nor U9819 (N_9819,N_9612,N_9739);
nor U9820 (N_9820,N_9686,N_9713);
and U9821 (N_9821,N_9636,N_9644);
or U9822 (N_9822,N_9537,N_9718);
and U9823 (N_9823,N_9726,N_9696);
xor U9824 (N_9824,N_9576,N_9685);
nor U9825 (N_9825,N_9602,N_9558);
or U9826 (N_9826,N_9519,N_9535);
or U9827 (N_9827,N_9571,N_9617);
nand U9828 (N_9828,N_9640,N_9579);
xor U9829 (N_9829,N_9530,N_9628);
nor U9830 (N_9830,N_9674,N_9551);
or U9831 (N_9831,N_9688,N_9556);
or U9832 (N_9832,N_9655,N_9743);
nand U9833 (N_9833,N_9529,N_9647);
and U9834 (N_9834,N_9678,N_9506);
xor U9835 (N_9835,N_9682,N_9747);
xor U9836 (N_9836,N_9650,N_9524);
and U9837 (N_9837,N_9734,N_9515);
nor U9838 (N_9838,N_9732,N_9634);
nor U9839 (N_9839,N_9570,N_9635);
xnor U9840 (N_9840,N_9597,N_9721);
nand U9841 (N_9841,N_9681,N_9554);
or U9842 (N_9842,N_9668,N_9677);
or U9843 (N_9843,N_9654,N_9748);
xor U9844 (N_9844,N_9651,N_9580);
xor U9845 (N_9845,N_9642,N_9715);
nand U9846 (N_9846,N_9641,N_9603);
xor U9847 (N_9847,N_9667,N_9742);
xnor U9848 (N_9848,N_9710,N_9619);
or U9849 (N_9849,N_9552,N_9587);
or U9850 (N_9850,N_9590,N_9540);
and U9851 (N_9851,N_9568,N_9588);
and U9852 (N_9852,N_9610,N_9670);
nor U9853 (N_9853,N_9596,N_9548);
nor U9854 (N_9854,N_9611,N_9517);
nor U9855 (N_9855,N_9533,N_9518);
and U9856 (N_9856,N_9624,N_9744);
xnor U9857 (N_9857,N_9606,N_9684);
nand U9858 (N_9858,N_9717,N_9649);
or U9859 (N_9859,N_9724,N_9666);
nand U9860 (N_9860,N_9735,N_9513);
and U9861 (N_9861,N_9633,N_9547);
nor U9862 (N_9862,N_9745,N_9616);
nand U9863 (N_9863,N_9637,N_9583);
and U9864 (N_9864,N_9599,N_9545);
nand U9865 (N_9865,N_9608,N_9702);
xnor U9866 (N_9866,N_9699,N_9600);
nand U9867 (N_9867,N_9564,N_9562);
nor U9868 (N_9868,N_9683,N_9528);
or U9869 (N_9869,N_9719,N_9604);
xor U9870 (N_9870,N_9729,N_9520);
or U9871 (N_9871,N_9598,N_9703);
or U9872 (N_9872,N_9567,N_9737);
or U9873 (N_9873,N_9605,N_9690);
or U9874 (N_9874,N_9534,N_9687);
xor U9875 (N_9875,N_9514,N_9552);
and U9876 (N_9876,N_9605,N_9557);
nand U9877 (N_9877,N_9531,N_9733);
nand U9878 (N_9878,N_9507,N_9639);
and U9879 (N_9879,N_9674,N_9691);
nor U9880 (N_9880,N_9639,N_9739);
nand U9881 (N_9881,N_9684,N_9632);
and U9882 (N_9882,N_9506,N_9522);
nor U9883 (N_9883,N_9644,N_9589);
xor U9884 (N_9884,N_9506,N_9582);
xor U9885 (N_9885,N_9514,N_9546);
xnor U9886 (N_9886,N_9696,N_9669);
or U9887 (N_9887,N_9502,N_9679);
nor U9888 (N_9888,N_9634,N_9626);
xor U9889 (N_9889,N_9504,N_9591);
xor U9890 (N_9890,N_9657,N_9580);
and U9891 (N_9891,N_9662,N_9742);
xnor U9892 (N_9892,N_9519,N_9741);
and U9893 (N_9893,N_9655,N_9608);
and U9894 (N_9894,N_9658,N_9592);
or U9895 (N_9895,N_9607,N_9563);
or U9896 (N_9896,N_9623,N_9632);
nor U9897 (N_9897,N_9656,N_9709);
nor U9898 (N_9898,N_9564,N_9711);
and U9899 (N_9899,N_9721,N_9511);
and U9900 (N_9900,N_9719,N_9715);
nor U9901 (N_9901,N_9618,N_9503);
xnor U9902 (N_9902,N_9671,N_9624);
and U9903 (N_9903,N_9620,N_9647);
nand U9904 (N_9904,N_9713,N_9703);
or U9905 (N_9905,N_9709,N_9620);
xor U9906 (N_9906,N_9738,N_9608);
and U9907 (N_9907,N_9586,N_9502);
nand U9908 (N_9908,N_9698,N_9638);
nand U9909 (N_9909,N_9643,N_9501);
or U9910 (N_9910,N_9555,N_9708);
or U9911 (N_9911,N_9674,N_9519);
xor U9912 (N_9912,N_9501,N_9749);
nor U9913 (N_9913,N_9648,N_9615);
nand U9914 (N_9914,N_9652,N_9548);
and U9915 (N_9915,N_9536,N_9741);
and U9916 (N_9916,N_9685,N_9592);
or U9917 (N_9917,N_9644,N_9731);
or U9918 (N_9918,N_9585,N_9659);
nor U9919 (N_9919,N_9520,N_9568);
and U9920 (N_9920,N_9630,N_9705);
or U9921 (N_9921,N_9657,N_9586);
and U9922 (N_9922,N_9701,N_9635);
or U9923 (N_9923,N_9664,N_9501);
nor U9924 (N_9924,N_9727,N_9712);
nand U9925 (N_9925,N_9697,N_9705);
nand U9926 (N_9926,N_9524,N_9616);
or U9927 (N_9927,N_9551,N_9552);
or U9928 (N_9928,N_9536,N_9728);
or U9929 (N_9929,N_9716,N_9533);
nor U9930 (N_9930,N_9536,N_9500);
and U9931 (N_9931,N_9680,N_9681);
nor U9932 (N_9932,N_9602,N_9685);
and U9933 (N_9933,N_9523,N_9582);
xor U9934 (N_9934,N_9609,N_9544);
nor U9935 (N_9935,N_9729,N_9631);
or U9936 (N_9936,N_9718,N_9719);
and U9937 (N_9937,N_9691,N_9600);
nor U9938 (N_9938,N_9571,N_9526);
nand U9939 (N_9939,N_9674,N_9647);
nor U9940 (N_9940,N_9710,N_9712);
or U9941 (N_9941,N_9570,N_9660);
xor U9942 (N_9942,N_9545,N_9713);
nand U9943 (N_9943,N_9734,N_9536);
nor U9944 (N_9944,N_9629,N_9615);
xor U9945 (N_9945,N_9559,N_9749);
nand U9946 (N_9946,N_9705,N_9717);
nor U9947 (N_9947,N_9504,N_9569);
nand U9948 (N_9948,N_9748,N_9563);
nand U9949 (N_9949,N_9695,N_9739);
or U9950 (N_9950,N_9553,N_9696);
nor U9951 (N_9951,N_9615,N_9562);
xnor U9952 (N_9952,N_9621,N_9582);
nor U9953 (N_9953,N_9695,N_9534);
nand U9954 (N_9954,N_9589,N_9565);
or U9955 (N_9955,N_9574,N_9637);
nand U9956 (N_9956,N_9619,N_9517);
nor U9957 (N_9957,N_9693,N_9578);
or U9958 (N_9958,N_9620,N_9540);
xnor U9959 (N_9959,N_9576,N_9619);
or U9960 (N_9960,N_9641,N_9565);
nor U9961 (N_9961,N_9501,N_9592);
xor U9962 (N_9962,N_9702,N_9576);
xnor U9963 (N_9963,N_9704,N_9730);
or U9964 (N_9964,N_9675,N_9686);
nor U9965 (N_9965,N_9512,N_9727);
nand U9966 (N_9966,N_9709,N_9682);
and U9967 (N_9967,N_9605,N_9535);
and U9968 (N_9968,N_9720,N_9611);
xnor U9969 (N_9969,N_9734,N_9540);
xnor U9970 (N_9970,N_9722,N_9704);
nor U9971 (N_9971,N_9703,N_9534);
xor U9972 (N_9972,N_9509,N_9610);
xor U9973 (N_9973,N_9706,N_9544);
nand U9974 (N_9974,N_9743,N_9671);
xnor U9975 (N_9975,N_9545,N_9660);
or U9976 (N_9976,N_9594,N_9552);
nand U9977 (N_9977,N_9506,N_9586);
nor U9978 (N_9978,N_9585,N_9541);
nand U9979 (N_9979,N_9606,N_9729);
nand U9980 (N_9980,N_9678,N_9638);
nor U9981 (N_9981,N_9546,N_9540);
and U9982 (N_9982,N_9692,N_9579);
xor U9983 (N_9983,N_9651,N_9729);
nand U9984 (N_9984,N_9581,N_9729);
nor U9985 (N_9985,N_9517,N_9596);
nand U9986 (N_9986,N_9577,N_9640);
nand U9987 (N_9987,N_9624,N_9537);
xnor U9988 (N_9988,N_9699,N_9561);
xnor U9989 (N_9989,N_9645,N_9643);
nand U9990 (N_9990,N_9526,N_9749);
nand U9991 (N_9991,N_9638,N_9705);
xnor U9992 (N_9992,N_9575,N_9567);
and U9993 (N_9993,N_9686,N_9508);
or U9994 (N_9994,N_9735,N_9653);
or U9995 (N_9995,N_9670,N_9621);
nand U9996 (N_9996,N_9601,N_9712);
and U9997 (N_9997,N_9565,N_9642);
and U9998 (N_9998,N_9703,N_9731);
nand U9999 (N_9999,N_9645,N_9523);
or U10000 (N_10000,N_9821,N_9829);
nand U10001 (N_10001,N_9760,N_9846);
xnor U10002 (N_10002,N_9867,N_9816);
or U10003 (N_10003,N_9775,N_9853);
or U10004 (N_10004,N_9861,N_9927);
and U10005 (N_10005,N_9944,N_9822);
nand U10006 (N_10006,N_9759,N_9902);
nand U10007 (N_10007,N_9795,N_9848);
or U10008 (N_10008,N_9995,N_9788);
xor U10009 (N_10009,N_9807,N_9987);
xor U10010 (N_10010,N_9933,N_9928);
and U10011 (N_10011,N_9947,N_9826);
nand U10012 (N_10012,N_9994,N_9998);
nand U10013 (N_10013,N_9959,N_9828);
nand U10014 (N_10014,N_9809,N_9942);
xnor U10015 (N_10015,N_9852,N_9844);
nor U10016 (N_10016,N_9909,N_9907);
nor U10017 (N_10017,N_9893,N_9929);
and U10018 (N_10018,N_9873,N_9895);
or U10019 (N_10019,N_9990,N_9777);
nand U10020 (N_10020,N_9903,N_9818);
or U10021 (N_10021,N_9765,N_9940);
nand U10022 (N_10022,N_9803,N_9962);
and U10023 (N_10023,N_9989,N_9810);
nand U10024 (N_10024,N_9876,N_9796);
nand U10025 (N_10025,N_9780,N_9812);
or U10026 (N_10026,N_9868,N_9839);
xor U10027 (N_10027,N_9771,N_9783);
nand U10028 (N_10028,N_9865,N_9923);
or U10029 (N_10029,N_9988,N_9952);
and U10030 (N_10030,N_9789,N_9911);
xnor U10031 (N_10031,N_9896,N_9924);
nor U10032 (N_10032,N_9931,N_9756);
xor U10033 (N_10033,N_9958,N_9851);
xor U10034 (N_10034,N_9901,N_9761);
and U10035 (N_10035,N_9755,N_9953);
and U10036 (N_10036,N_9811,N_9872);
or U10037 (N_10037,N_9972,N_9824);
and U10038 (N_10038,N_9913,N_9831);
nor U10039 (N_10039,N_9770,N_9887);
xor U10040 (N_10040,N_9955,N_9763);
nand U10041 (N_10041,N_9830,N_9856);
xnor U10042 (N_10042,N_9773,N_9925);
xnor U10043 (N_10043,N_9941,N_9974);
nor U10044 (N_10044,N_9758,N_9936);
or U10045 (N_10045,N_9918,N_9782);
or U10046 (N_10046,N_9808,N_9769);
nor U10047 (N_10047,N_9900,N_9813);
nor U10048 (N_10048,N_9910,N_9875);
and U10049 (N_10049,N_9983,N_9916);
xnor U10050 (N_10050,N_9843,N_9915);
xor U10051 (N_10051,N_9835,N_9863);
xnor U10052 (N_10052,N_9871,N_9800);
xor U10053 (N_10053,N_9817,N_9975);
nand U10054 (N_10054,N_9791,N_9870);
nand U10055 (N_10055,N_9804,N_9914);
xnor U10056 (N_10056,N_9898,N_9966);
and U10057 (N_10057,N_9881,N_9957);
nor U10058 (N_10058,N_9982,N_9855);
and U10059 (N_10059,N_9781,N_9890);
nor U10060 (N_10060,N_9798,N_9930);
nor U10061 (N_10061,N_9885,N_9820);
and U10062 (N_10062,N_9778,N_9912);
nand U10063 (N_10063,N_9935,N_9869);
nand U10064 (N_10064,N_9946,N_9754);
or U10065 (N_10065,N_9978,N_9840);
xor U10066 (N_10066,N_9859,N_9794);
nor U10067 (N_10067,N_9834,N_9945);
xnor U10068 (N_10068,N_9787,N_9969);
nand U10069 (N_10069,N_9776,N_9973);
or U10070 (N_10070,N_9920,N_9797);
and U10071 (N_10071,N_9971,N_9779);
nand U10072 (N_10072,N_9979,N_9850);
xor U10073 (N_10073,N_9956,N_9841);
nor U10074 (N_10074,N_9950,N_9943);
nor U10075 (N_10075,N_9993,N_9792);
or U10076 (N_10076,N_9772,N_9805);
or U10077 (N_10077,N_9823,N_9836);
and U10078 (N_10078,N_9894,N_9751);
and U10079 (N_10079,N_9825,N_9784);
xnor U10080 (N_10080,N_9806,N_9926);
xor U10081 (N_10081,N_9768,N_9968);
or U10082 (N_10082,N_9985,N_9827);
nand U10083 (N_10083,N_9854,N_9984);
or U10084 (N_10084,N_9980,N_9981);
nand U10085 (N_10085,N_9889,N_9954);
nand U10086 (N_10086,N_9764,N_9802);
or U10087 (N_10087,N_9938,N_9961);
and U10088 (N_10088,N_9977,N_9858);
or U10089 (N_10089,N_9877,N_9874);
nand U10090 (N_10090,N_9767,N_9752);
xnor U10091 (N_10091,N_9837,N_9939);
and U10092 (N_10092,N_9908,N_9891);
or U10093 (N_10093,N_9880,N_9948);
xor U10094 (N_10094,N_9965,N_9857);
nand U10095 (N_10095,N_9904,N_9999);
and U10096 (N_10096,N_9847,N_9963);
nor U10097 (N_10097,N_9862,N_9917);
nor U10098 (N_10098,N_9919,N_9878);
nor U10099 (N_10099,N_9892,N_9864);
and U10100 (N_10100,N_9860,N_9976);
xnor U10101 (N_10101,N_9986,N_9785);
nor U10102 (N_10102,N_9786,N_9815);
xor U10103 (N_10103,N_9997,N_9879);
or U10104 (N_10104,N_9801,N_9814);
or U10105 (N_10105,N_9991,N_9883);
and U10106 (N_10106,N_9845,N_9757);
and U10107 (N_10107,N_9922,N_9932);
nor U10108 (N_10108,N_9967,N_9906);
nand U10109 (N_10109,N_9819,N_9934);
or U10110 (N_10110,N_9766,N_9970);
and U10111 (N_10111,N_9884,N_9937);
and U10112 (N_10112,N_9832,N_9949);
and U10113 (N_10113,N_9762,N_9951);
or U10114 (N_10114,N_9882,N_9921);
nor U10115 (N_10115,N_9964,N_9793);
or U10116 (N_10116,N_9753,N_9774);
nor U10117 (N_10117,N_9842,N_9849);
xor U10118 (N_10118,N_9899,N_9799);
nand U10119 (N_10119,N_9886,N_9866);
xor U10120 (N_10120,N_9888,N_9833);
or U10121 (N_10121,N_9790,N_9996);
nor U10122 (N_10122,N_9838,N_9992);
nand U10123 (N_10123,N_9750,N_9897);
nor U10124 (N_10124,N_9905,N_9960);
nor U10125 (N_10125,N_9821,N_9904);
nor U10126 (N_10126,N_9989,N_9915);
xor U10127 (N_10127,N_9878,N_9839);
nor U10128 (N_10128,N_9891,N_9881);
nand U10129 (N_10129,N_9969,N_9812);
and U10130 (N_10130,N_9869,N_9918);
nor U10131 (N_10131,N_9781,N_9823);
and U10132 (N_10132,N_9880,N_9828);
and U10133 (N_10133,N_9807,N_9804);
xor U10134 (N_10134,N_9942,N_9940);
and U10135 (N_10135,N_9878,N_9890);
nor U10136 (N_10136,N_9998,N_9927);
xor U10137 (N_10137,N_9857,N_9886);
xnor U10138 (N_10138,N_9769,N_9816);
nand U10139 (N_10139,N_9938,N_9779);
xnor U10140 (N_10140,N_9907,N_9929);
and U10141 (N_10141,N_9927,N_9951);
nor U10142 (N_10142,N_9756,N_9772);
nand U10143 (N_10143,N_9769,N_9869);
nor U10144 (N_10144,N_9859,N_9898);
and U10145 (N_10145,N_9759,N_9956);
and U10146 (N_10146,N_9766,N_9880);
or U10147 (N_10147,N_9804,N_9960);
or U10148 (N_10148,N_9913,N_9930);
nand U10149 (N_10149,N_9896,N_9823);
nor U10150 (N_10150,N_9764,N_9767);
nand U10151 (N_10151,N_9863,N_9852);
xnor U10152 (N_10152,N_9864,N_9773);
nand U10153 (N_10153,N_9987,N_9811);
nor U10154 (N_10154,N_9944,N_9785);
and U10155 (N_10155,N_9799,N_9833);
nor U10156 (N_10156,N_9956,N_9992);
xor U10157 (N_10157,N_9805,N_9972);
xnor U10158 (N_10158,N_9906,N_9805);
xnor U10159 (N_10159,N_9773,N_9900);
nor U10160 (N_10160,N_9902,N_9755);
and U10161 (N_10161,N_9790,N_9780);
or U10162 (N_10162,N_9986,N_9766);
nand U10163 (N_10163,N_9917,N_9764);
and U10164 (N_10164,N_9782,N_9800);
xor U10165 (N_10165,N_9821,N_9860);
nand U10166 (N_10166,N_9835,N_9928);
nor U10167 (N_10167,N_9760,N_9917);
nor U10168 (N_10168,N_9905,N_9766);
nand U10169 (N_10169,N_9919,N_9804);
nand U10170 (N_10170,N_9756,N_9911);
nor U10171 (N_10171,N_9932,N_9796);
or U10172 (N_10172,N_9810,N_9805);
or U10173 (N_10173,N_9976,N_9878);
nor U10174 (N_10174,N_9763,N_9793);
and U10175 (N_10175,N_9817,N_9781);
nor U10176 (N_10176,N_9886,N_9835);
xnor U10177 (N_10177,N_9991,N_9823);
nor U10178 (N_10178,N_9901,N_9990);
and U10179 (N_10179,N_9941,N_9831);
nand U10180 (N_10180,N_9827,N_9892);
and U10181 (N_10181,N_9814,N_9776);
or U10182 (N_10182,N_9897,N_9971);
or U10183 (N_10183,N_9909,N_9766);
xor U10184 (N_10184,N_9808,N_9854);
nand U10185 (N_10185,N_9777,N_9809);
and U10186 (N_10186,N_9923,N_9930);
nand U10187 (N_10187,N_9772,N_9939);
nor U10188 (N_10188,N_9790,N_9921);
or U10189 (N_10189,N_9886,N_9862);
or U10190 (N_10190,N_9832,N_9960);
or U10191 (N_10191,N_9963,N_9764);
and U10192 (N_10192,N_9982,N_9752);
xor U10193 (N_10193,N_9816,N_9797);
or U10194 (N_10194,N_9912,N_9751);
nor U10195 (N_10195,N_9791,N_9824);
xor U10196 (N_10196,N_9833,N_9807);
nor U10197 (N_10197,N_9869,N_9938);
nor U10198 (N_10198,N_9862,N_9911);
nand U10199 (N_10199,N_9768,N_9912);
nand U10200 (N_10200,N_9968,N_9875);
and U10201 (N_10201,N_9912,N_9763);
xor U10202 (N_10202,N_9850,N_9810);
nand U10203 (N_10203,N_9808,N_9929);
nor U10204 (N_10204,N_9990,N_9784);
nand U10205 (N_10205,N_9818,N_9879);
or U10206 (N_10206,N_9771,N_9881);
nand U10207 (N_10207,N_9868,N_9996);
nor U10208 (N_10208,N_9979,N_9891);
xnor U10209 (N_10209,N_9838,N_9880);
nand U10210 (N_10210,N_9797,N_9974);
xnor U10211 (N_10211,N_9945,N_9905);
nor U10212 (N_10212,N_9979,N_9937);
xnor U10213 (N_10213,N_9877,N_9777);
nand U10214 (N_10214,N_9971,N_9821);
and U10215 (N_10215,N_9899,N_9988);
xnor U10216 (N_10216,N_9875,N_9926);
nor U10217 (N_10217,N_9774,N_9987);
nor U10218 (N_10218,N_9987,N_9933);
or U10219 (N_10219,N_9937,N_9844);
nor U10220 (N_10220,N_9802,N_9820);
and U10221 (N_10221,N_9848,N_9957);
nor U10222 (N_10222,N_9927,N_9762);
xnor U10223 (N_10223,N_9891,N_9909);
nand U10224 (N_10224,N_9926,N_9776);
nand U10225 (N_10225,N_9980,N_9937);
or U10226 (N_10226,N_9973,N_9824);
and U10227 (N_10227,N_9958,N_9780);
and U10228 (N_10228,N_9854,N_9947);
or U10229 (N_10229,N_9960,N_9982);
nor U10230 (N_10230,N_9800,N_9836);
nor U10231 (N_10231,N_9920,N_9770);
nand U10232 (N_10232,N_9809,N_9988);
nand U10233 (N_10233,N_9949,N_9789);
or U10234 (N_10234,N_9895,N_9814);
nor U10235 (N_10235,N_9815,N_9856);
nor U10236 (N_10236,N_9877,N_9927);
nor U10237 (N_10237,N_9822,N_9934);
or U10238 (N_10238,N_9824,N_9847);
or U10239 (N_10239,N_9776,N_9767);
xnor U10240 (N_10240,N_9940,N_9901);
xnor U10241 (N_10241,N_9847,N_9892);
nand U10242 (N_10242,N_9775,N_9801);
nand U10243 (N_10243,N_9946,N_9832);
xor U10244 (N_10244,N_9772,N_9789);
nor U10245 (N_10245,N_9959,N_9933);
nand U10246 (N_10246,N_9793,N_9785);
nor U10247 (N_10247,N_9980,N_9935);
nand U10248 (N_10248,N_9987,N_9854);
nor U10249 (N_10249,N_9918,N_9877);
or U10250 (N_10250,N_10067,N_10124);
nor U10251 (N_10251,N_10145,N_10172);
or U10252 (N_10252,N_10135,N_10204);
xor U10253 (N_10253,N_10087,N_10000);
xor U10254 (N_10254,N_10032,N_10120);
xor U10255 (N_10255,N_10121,N_10035);
and U10256 (N_10256,N_10176,N_10239);
xnor U10257 (N_10257,N_10137,N_10225);
and U10258 (N_10258,N_10136,N_10112);
xor U10259 (N_10259,N_10233,N_10146);
and U10260 (N_10260,N_10127,N_10119);
or U10261 (N_10261,N_10184,N_10248);
nor U10262 (N_10262,N_10059,N_10048);
nand U10263 (N_10263,N_10181,N_10066);
xor U10264 (N_10264,N_10062,N_10235);
xor U10265 (N_10265,N_10208,N_10213);
nand U10266 (N_10266,N_10115,N_10011);
or U10267 (N_10267,N_10231,N_10168);
nand U10268 (N_10268,N_10132,N_10064);
xnor U10269 (N_10269,N_10243,N_10188);
xor U10270 (N_10270,N_10102,N_10244);
nor U10271 (N_10271,N_10015,N_10042);
and U10272 (N_10272,N_10221,N_10185);
or U10273 (N_10273,N_10074,N_10077);
and U10274 (N_10274,N_10163,N_10100);
nor U10275 (N_10275,N_10031,N_10018);
xnor U10276 (N_10276,N_10003,N_10187);
nor U10277 (N_10277,N_10060,N_10026);
or U10278 (N_10278,N_10073,N_10218);
xor U10279 (N_10279,N_10078,N_10023);
nor U10280 (N_10280,N_10098,N_10211);
xor U10281 (N_10281,N_10193,N_10104);
nand U10282 (N_10282,N_10099,N_10021);
nor U10283 (N_10283,N_10128,N_10084);
or U10284 (N_10284,N_10169,N_10151);
nor U10285 (N_10285,N_10045,N_10170);
nand U10286 (N_10286,N_10139,N_10116);
and U10287 (N_10287,N_10079,N_10105);
nand U10288 (N_10288,N_10182,N_10140);
and U10289 (N_10289,N_10072,N_10175);
and U10290 (N_10290,N_10006,N_10227);
xor U10291 (N_10291,N_10138,N_10070);
or U10292 (N_10292,N_10229,N_10126);
nor U10293 (N_10293,N_10008,N_10174);
and U10294 (N_10294,N_10232,N_10010);
nand U10295 (N_10295,N_10001,N_10061);
and U10296 (N_10296,N_10228,N_10052);
and U10297 (N_10297,N_10162,N_10224);
nand U10298 (N_10298,N_10220,N_10241);
or U10299 (N_10299,N_10009,N_10065);
nor U10300 (N_10300,N_10212,N_10028);
and U10301 (N_10301,N_10161,N_10216);
and U10302 (N_10302,N_10081,N_10201);
xnor U10303 (N_10303,N_10196,N_10198);
nor U10304 (N_10304,N_10049,N_10144);
and U10305 (N_10305,N_10171,N_10106);
or U10306 (N_10306,N_10056,N_10058);
or U10307 (N_10307,N_10155,N_10152);
nand U10308 (N_10308,N_10027,N_10095);
and U10309 (N_10309,N_10207,N_10071);
or U10310 (N_10310,N_10090,N_10205);
and U10311 (N_10311,N_10178,N_10055);
nor U10312 (N_10312,N_10157,N_10075);
or U10313 (N_10313,N_10160,N_10093);
nand U10314 (N_10314,N_10226,N_10051);
nand U10315 (N_10315,N_10223,N_10222);
or U10316 (N_10316,N_10020,N_10114);
nand U10317 (N_10317,N_10200,N_10177);
nor U10318 (N_10318,N_10167,N_10215);
or U10319 (N_10319,N_10016,N_10203);
xor U10320 (N_10320,N_10166,N_10123);
nor U10321 (N_10321,N_10063,N_10149);
nor U10322 (N_10322,N_10012,N_10110);
and U10323 (N_10323,N_10158,N_10113);
and U10324 (N_10324,N_10234,N_10085);
and U10325 (N_10325,N_10037,N_10014);
and U10326 (N_10326,N_10199,N_10034);
nand U10327 (N_10327,N_10044,N_10089);
and U10328 (N_10328,N_10013,N_10206);
nor U10329 (N_10329,N_10156,N_10019);
and U10330 (N_10330,N_10097,N_10080);
or U10331 (N_10331,N_10219,N_10125);
xor U10332 (N_10332,N_10133,N_10047);
or U10333 (N_10333,N_10165,N_10083);
or U10334 (N_10334,N_10154,N_10173);
nand U10335 (N_10335,N_10094,N_10148);
or U10336 (N_10336,N_10242,N_10164);
nor U10337 (N_10337,N_10039,N_10134);
nor U10338 (N_10338,N_10053,N_10030);
nand U10339 (N_10339,N_10109,N_10057);
nand U10340 (N_10340,N_10246,N_10101);
and U10341 (N_10341,N_10189,N_10025);
nand U10342 (N_10342,N_10118,N_10194);
and U10343 (N_10343,N_10091,N_10122);
or U10344 (N_10344,N_10143,N_10069);
nor U10345 (N_10345,N_10179,N_10017);
or U10346 (N_10346,N_10130,N_10108);
xnor U10347 (N_10347,N_10237,N_10197);
nand U10348 (N_10348,N_10022,N_10086);
or U10349 (N_10349,N_10142,N_10129);
nand U10350 (N_10350,N_10247,N_10043);
or U10351 (N_10351,N_10217,N_10159);
or U10352 (N_10352,N_10209,N_10041);
nand U10353 (N_10353,N_10190,N_10004);
or U10354 (N_10354,N_10050,N_10180);
and U10355 (N_10355,N_10238,N_10195);
xor U10356 (N_10356,N_10036,N_10040);
and U10357 (N_10357,N_10054,N_10214);
nor U10358 (N_10358,N_10153,N_10186);
nand U10359 (N_10359,N_10096,N_10007);
xnor U10360 (N_10360,N_10024,N_10103);
or U10361 (N_10361,N_10002,N_10150);
nor U10362 (N_10362,N_10107,N_10005);
and U10363 (N_10363,N_10236,N_10147);
or U10364 (N_10364,N_10183,N_10068);
nor U10365 (N_10365,N_10076,N_10029);
nor U10366 (N_10366,N_10240,N_10249);
or U10367 (N_10367,N_10088,N_10202);
and U10368 (N_10368,N_10210,N_10245);
and U10369 (N_10369,N_10111,N_10230);
nand U10370 (N_10370,N_10046,N_10033);
nor U10371 (N_10371,N_10082,N_10038);
xor U10372 (N_10372,N_10191,N_10192);
and U10373 (N_10373,N_10131,N_10117);
and U10374 (N_10374,N_10141,N_10092);
or U10375 (N_10375,N_10220,N_10016);
xor U10376 (N_10376,N_10133,N_10163);
and U10377 (N_10377,N_10088,N_10064);
or U10378 (N_10378,N_10052,N_10100);
or U10379 (N_10379,N_10092,N_10044);
or U10380 (N_10380,N_10187,N_10043);
xnor U10381 (N_10381,N_10180,N_10012);
or U10382 (N_10382,N_10031,N_10242);
nand U10383 (N_10383,N_10241,N_10105);
nand U10384 (N_10384,N_10070,N_10102);
and U10385 (N_10385,N_10186,N_10234);
xnor U10386 (N_10386,N_10131,N_10067);
nand U10387 (N_10387,N_10184,N_10075);
xor U10388 (N_10388,N_10173,N_10103);
xor U10389 (N_10389,N_10117,N_10027);
nor U10390 (N_10390,N_10100,N_10068);
and U10391 (N_10391,N_10188,N_10008);
nor U10392 (N_10392,N_10174,N_10029);
nor U10393 (N_10393,N_10091,N_10076);
or U10394 (N_10394,N_10097,N_10159);
nor U10395 (N_10395,N_10244,N_10008);
nand U10396 (N_10396,N_10244,N_10020);
or U10397 (N_10397,N_10240,N_10005);
nand U10398 (N_10398,N_10248,N_10110);
or U10399 (N_10399,N_10237,N_10049);
and U10400 (N_10400,N_10095,N_10050);
nor U10401 (N_10401,N_10210,N_10027);
or U10402 (N_10402,N_10080,N_10088);
and U10403 (N_10403,N_10019,N_10063);
nor U10404 (N_10404,N_10230,N_10075);
and U10405 (N_10405,N_10192,N_10149);
and U10406 (N_10406,N_10003,N_10135);
xnor U10407 (N_10407,N_10020,N_10130);
nand U10408 (N_10408,N_10020,N_10077);
nand U10409 (N_10409,N_10243,N_10080);
nand U10410 (N_10410,N_10230,N_10135);
and U10411 (N_10411,N_10111,N_10164);
or U10412 (N_10412,N_10217,N_10226);
or U10413 (N_10413,N_10064,N_10121);
xor U10414 (N_10414,N_10055,N_10219);
xnor U10415 (N_10415,N_10164,N_10002);
or U10416 (N_10416,N_10015,N_10241);
nand U10417 (N_10417,N_10178,N_10152);
or U10418 (N_10418,N_10030,N_10014);
or U10419 (N_10419,N_10148,N_10233);
nor U10420 (N_10420,N_10218,N_10232);
nand U10421 (N_10421,N_10096,N_10151);
nand U10422 (N_10422,N_10213,N_10103);
nand U10423 (N_10423,N_10226,N_10029);
or U10424 (N_10424,N_10166,N_10204);
nand U10425 (N_10425,N_10222,N_10163);
nor U10426 (N_10426,N_10019,N_10135);
xnor U10427 (N_10427,N_10143,N_10048);
xor U10428 (N_10428,N_10241,N_10185);
or U10429 (N_10429,N_10039,N_10179);
nand U10430 (N_10430,N_10074,N_10110);
nand U10431 (N_10431,N_10083,N_10204);
xnor U10432 (N_10432,N_10208,N_10156);
or U10433 (N_10433,N_10245,N_10211);
nand U10434 (N_10434,N_10187,N_10124);
xnor U10435 (N_10435,N_10091,N_10079);
xnor U10436 (N_10436,N_10151,N_10119);
or U10437 (N_10437,N_10186,N_10114);
and U10438 (N_10438,N_10225,N_10163);
xnor U10439 (N_10439,N_10016,N_10006);
nand U10440 (N_10440,N_10218,N_10032);
or U10441 (N_10441,N_10105,N_10184);
xnor U10442 (N_10442,N_10198,N_10093);
nand U10443 (N_10443,N_10198,N_10011);
nor U10444 (N_10444,N_10085,N_10162);
and U10445 (N_10445,N_10227,N_10109);
or U10446 (N_10446,N_10006,N_10106);
and U10447 (N_10447,N_10180,N_10084);
and U10448 (N_10448,N_10206,N_10203);
nand U10449 (N_10449,N_10157,N_10130);
nand U10450 (N_10450,N_10184,N_10084);
nand U10451 (N_10451,N_10060,N_10011);
nor U10452 (N_10452,N_10113,N_10166);
nand U10453 (N_10453,N_10216,N_10152);
xnor U10454 (N_10454,N_10177,N_10060);
or U10455 (N_10455,N_10037,N_10065);
and U10456 (N_10456,N_10201,N_10126);
nor U10457 (N_10457,N_10020,N_10242);
xor U10458 (N_10458,N_10211,N_10195);
or U10459 (N_10459,N_10179,N_10085);
xnor U10460 (N_10460,N_10157,N_10245);
and U10461 (N_10461,N_10124,N_10188);
nor U10462 (N_10462,N_10045,N_10114);
xnor U10463 (N_10463,N_10152,N_10031);
and U10464 (N_10464,N_10165,N_10201);
and U10465 (N_10465,N_10113,N_10104);
and U10466 (N_10466,N_10192,N_10116);
or U10467 (N_10467,N_10110,N_10222);
or U10468 (N_10468,N_10051,N_10152);
and U10469 (N_10469,N_10219,N_10052);
and U10470 (N_10470,N_10091,N_10248);
nor U10471 (N_10471,N_10056,N_10025);
xnor U10472 (N_10472,N_10221,N_10012);
xnor U10473 (N_10473,N_10003,N_10143);
xnor U10474 (N_10474,N_10095,N_10052);
xor U10475 (N_10475,N_10004,N_10067);
nor U10476 (N_10476,N_10130,N_10090);
xnor U10477 (N_10477,N_10113,N_10229);
nor U10478 (N_10478,N_10159,N_10215);
xnor U10479 (N_10479,N_10151,N_10078);
nor U10480 (N_10480,N_10095,N_10096);
and U10481 (N_10481,N_10006,N_10226);
nor U10482 (N_10482,N_10031,N_10029);
and U10483 (N_10483,N_10155,N_10178);
nor U10484 (N_10484,N_10095,N_10194);
nand U10485 (N_10485,N_10151,N_10192);
nor U10486 (N_10486,N_10169,N_10246);
xnor U10487 (N_10487,N_10109,N_10171);
xnor U10488 (N_10488,N_10222,N_10030);
nor U10489 (N_10489,N_10050,N_10037);
nor U10490 (N_10490,N_10086,N_10035);
nand U10491 (N_10491,N_10048,N_10116);
and U10492 (N_10492,N_10108,N_10134);
xor U10493 (N_10493,N_10163,N_10217);
nor U10494 (N_10494,N_10097,N_10186);
nor U10495 (N_10495,N_10090,N_10005);
xor U10496 (N_10496,N_10189,N_10091);
or U10497 (N_10497,N_10233,N_10107);
or U10498 (N_10498,N_10031,N_10060);
nand U10499 (N_10499,N_10151,N_10226);
xnor U10500 (N_10500,N_10317,N_10425);
nor U10501 (N_10501,N_10496,N_10490);
and U10502 (N_10502,N_10360,N_10277);
nor U10503 (N_10503,N_10497,N_10355);
nor U10504 (N_10504,N_10255,N_10303);
xnor U10505 (N_10505,N_10482,N_10256);
or U10506 (N_10506,N_10263,N_10295);
nor U10507 (N_10507,N_10310,N_10361);
and U10508 (N_10508,N_10286,N_10331);
xnor U10509 (N_10509,N_10393,N_10399);
nor U10510 (N_10510,N_10300,N_10294);
nand U10511 (N_10511,N_10391,N_10264);
and U10512 (N_10512,N_10440,N_10437);
nor U10513 (N_10513,N_10333,N_10441);
xor U10514 (N_10514,N_10311,N_10473);
xnor U10515 (N_10515,N_10357,N_10396);
xor U10516 (N_10516,N_10340,N_10252);
and U10517 (N_10517,N_10498,N_10327);
nor U10518 (N_10518,N_10292,N_10261);
nand U10519 (N_10519,N_10301,N_10459);
nor U10520 (N_10520,N_10332,N_10312);
xor U10521 (N_10521,N_10350,N_10345);
xor U10522 (N_10522,N_10417,N_10379);
nand U10523 (N_10523,N_10339,N_10401);
xnor U10524 (N_10524,N_10439,N_10318);
nand U10525 (N_10525,N_10398,N_10455);
and U10526 (N_10526,N_10383,N_10486);
or U10527 (N_10527,N_10328,N_10316);
and U10528 (N_10528,N_10403,N_10274);
xor U10529 (N_10529,N_10260,N_10374);
xor U10530 (N_10530,N_10409,N_10484);
nor U10531 (N_10531,N_10472,N_10422);
nand U10532 (N_10532,N_10481,N_10290);
and U10533 (N_10533,N_10358,N_10450);
or U10534 (N_10534,N_10352,N_10341);
or U10535 (N_10535,N_10412,N_10436);
xor U10536 (N_10536,N_10381,N_10414);
xor U10537 (N_10537,N_10298,N_10434);
nor U10538 (N_10538,N_10426,N_10429);
or U10539 (N_10539,N_10377,N_10489);
or U10540 (N_10540,N_10454,N_10424);
and U10541 (N_10541,N_10325,N_10467);
or U10542 (N_10542,N_10281,N_10308);
nor U10543 (N_10543,N_10433,N_10322);
and U10544 (N_10544,N_10423,N_10477);
xor U10545 (N_10545,N_10368,N_10289);
nand U10546 (N_10546,N_10428,N_10445);
and U10547 (N_10547,N_10373,N_10456);
nor U10548 (N_10548,N_10348,N_10468);
or U10549 (N_10549,N_10307,N_10461);
and U10550 (N_10550,N_10278,N_10478);
xor U10551 (N_10551,N_10287,N_10394);
or U10552 (N_10552,N_10465,N_10452);
xor U10553 (N_10553,N_10389,N_10280);
nand U10554 (N_10554,N_10458,N_10438);
xor U10555 (N_10555,N_10330,N_10251);
or U10556 (N_10556,N_10435,N_10375);
nor U10557 (N_10557,N_10343,N_10315);
or U10558 (N_10558,N_10250,N_10378);
or U10559 (N_10559,N_10356,N_10366);
or U10560 (N_10560,N_10432,N_10367);
or U10561 (N_10561,N_10272,N_10276);
nor U10562 (N_10562,N_10466,N_10408);
or U10563 (N_10563,N_10268,N_10476);
xor U10564 (N_10564,N_10411,N_10388);
or U10565 (N_10565,N_10314,N_10321);
xor U10566 (N_10566,N_10364,N_10320);
xor U10567 (N_10567,N_10338,N_10487);
xnor U10568 (N_10568,N_10460,N_10380);
xor U10569 (N_10569,N_10397,N_10479);
nand U10570 (N_10570,N_10386,N_10370);
nor U10571 (N_10571,N_10387,N_10362);
nand U10572 (N_10572,N_10447,N_10323);
xor U10573 (N_10573,N_10371,N_10329);
nand U10574 (N_10574,N_10336,N_10271);
nor U10575 (N_10575,N_10267,N_10449);
xnor U10576 (N_10576,N_10359,N_10363);
or U10577 (N_10577,N_10406,N_10353);
and U10578 (N_10578,N_10419,N_10495);
nand U10579 (N_10579,N_10384,N_10365);
or U10580 (N_10580,N_10291,N_10418);
nor U10581 (N_10581,N_10475,N_10376);
and U10582 (N_10582,N_10269,N_10257);
xor U10583 (N_10583,N_10313,N_10491);
nand U10584 (N_10584,N_10444,N_10347);
nand U10585 (N_10585,N_10342,N_10483);
nand U10586 (N_10586,N_10369,N_10453);
and U10587 (N_10587,N_10337,N_10283);
nor U10588 (N_10588,N_10488,N_10385);
or U10589 (N_10589,N_10259,N_10469);
nand U10590 (N_10590,N_10480,N_10265);
xnor U10591 (N_10591,N_10494,N_10297);
and U10592 (N_10592,N_10407,N_10354);
xor U10593 (N_10593,N_10326,N_10344);
nor U10594 (N_10594,N_10395,N_10442);
and U10595 (N_10595,N_10402,N_10416);
xor U10596 (N_10596,N_10253,N_10270);
nor U10597 (N_10597,N_10448,N_10427);
nand U10598 (N_10598,N_10346,N_10392);
nor U10599 (N_10599,N_10262,N_10420);
xor U10600 (N_10600,N_10485,N_10335);
and U10601 (N_10601,N_10443,N_10349);
nor U10602 (N_10602,N_10306,N_10254);
nand U10603 (N_10603,N_10470,N_10492);
and U10604 (N_10604,N_10299,N_10372);
nor U10605 (N_10605,N_10471,N_10351);
or U10606 (N_10606,N_10382,N_10304);
and U10607 (N_10607,N_10275,N_10457);
nand U10608 (N_10608,N_10309,N_10279);
or U10609 (N_10609,N_10463,N_10400);
nand U10610 (N_10610,N_10464,N_10390);
nor U10611 (N_10611,N_10334,N_10305);
xor U10612 (N_10612,N_10266,N_10430);
or U10613 (N_10613,N_10474,N_10451);
or U10614 (N_10614,N_10410,N_10405);
or U10615 (N_10615,N_10462,N_10293);
and U10616 (N_10616,N_10421,N_10493);
nor U10617 (N_10617,N_10413,N_10319);
nand U10618 (N_10618,N_10285,N_10302);
or U10619 (N_10619,N_10258,N_10282);
nand U10620 (N_10620,N_10324,N_10288);
xnor U10621 (N_10621,N_10431,N_10296);
or U10622 (N_10622,N_10273,N_10284);
or U10623 (N_10623,N_10446,N_10404);
and U10624 (N_10624,N_10415,N_10499);
xnor U10625 (N_10625,N_10254,N_10451);
and U10626 (N_10626,N_10311,N_10295);
and U10627 (N_10627,N_10256,N_10490);
nand U10628 (N_10628,N_10417,N_10304);
and U10629 (N_10629,N_10367,N_10343);
and U10630 (N_10630,N_10438,N_10258);
and U10631 (N_10631,N_10469,N_10290);
and U10632 (N_10632,N_10440,N_10326);
and U10633 (N_10633,N_10335,N_10496);
nor U10634 (N_10634,N_10390,N_10397);
or U10635 (N_10635,N_10416,N_10414);
or U10636 (N_10636,N_10333,N_10412);
and U10637 (N_10637,N_10362,N_10349);
nor U10638 (N_10638,N_10480,N_10447);
nor U10639 (N_10639,N_10384,N_10478);
nor U10640 (N_10640,N_10328,N_10266);
nand U10641 (N_10641,N_10419,N_10250);
nor U10642 (N_10642,N_10264,N_10404);
xor U10643 (N_10643,N_10325,N_10285);
nor U10644 (N_10644,N_10332,N_10409);
or U10645 (N_10645,N_10479,N_10407);
or U10646 (N_10646,N_10469,N_10358);
xnor U10647 (N_10647,N_10429,N_10277);
nor U10648 (N_10648,N_10319,N_10433);
or U10649 (N_10649,N_10487,N_10257);
nand U10650 (N_10650,N_10382,N_10451);
or U10651 (N_10651,N_10379,N_10479);
or U10652 (N_10652,N_10330,N_10264);
nand U10653 (N_10653,N_10312,N_10363);
nand U10654 (N_10654,N_10383,N_10391);
or U10655 (N_10655,N_10354,N_10250);
nand U10656 (N_10656,N_10417,N_10252);
or U10657 (N_10657,N_10262,N_10329);
xnor U10658 (N_10658,N_10280,N_10419);
nand U10659 (N_10659,N_10296,N_10338);
or U10660 (N_10660,N_10473,N_10370);
and U10661 (N_10661,N_10257,N_10366);
xor U10662 (N_10662,N_10353,N_10312);
or U10663 (N_10663,N_10284,N_10352);
nand U10664 (N_10664,N_10357,N_10466);
nand U10665 (N_10665,N_10332,N_10393);
or U10666 (N_10666,N_10371,N_10412);
nand U10667 (N_10667,N_10251,N_10364);
or U10668 (N_10668,N_10355,N_10420);
nand U10669 (N_10669,N_10374,N_10417);
nand U10670 (N_10670,N_10335,N_10363);
xnor U10671 (N_10671,N_10359,N_10267);
xnor U10672 (N_10672,N_10491,N_10259);
or U10673 (N_10673,N_10488,N_10474);
xnor U10674 (N_10674,N_10263,N_10464);
nor U10675 (N_10675,N_10286,N_10336);
nor U10676 (N_10676,N_10320,N_10275);
nand U10677 (N_10677,N_10266,N_10362);
nor U10678 (N_10678,N_10463,N_10473);
nor U10679 (N_10679,N_10400,N_10399);
and U10680 (N_10680,N_10298,N_10319);
nand U10681 (N_10681,N_10465,N_10263);
or U10682 (N_10682,N_10453,N_10435);
and U10683 (N_10683,N_10271,N_10353);
and U10684 (N_10684,N_10371,N_10283);
and U10685 (N_10685,N_10379,N_10378);
nand U10686 (N_10686,N_10251,N_10317);
nor U10687 (N_10687,N_10337,N_10279);
nand U10688 (N_10688,N_10484,N_10319);
and U10689 (N_10689,N_10384,N_10345);
or U10690 (N_10690,N_10463,N_10495);
xor U10691 (N_10691,N_10486,N_10467);
nand U10692 (N_10692,N_10363,N_10383);
xor U10693 (N_10693,N_10281,N_10362);
nor U10694 (N_10694,N_10373,N_10440);
xor U10695 (N_10695,N_10435,N_10306);
xnor U10696 (N_10696,N_10273,N_10323);
nand U10697 (N_10697,N_10281,N_10427);
nor U10698 (N_10698,N_10336,N_10466);
and U10699 (N_10699,N_10485,N_10316);
xor U10700 (N_10700,N_10465,N_10448);
and U10701 (N_10701,N_10398,N_10359);
nand U10702 (N_10702,N_10336,N_10403);
nand U10703 (N_10703,N_10429,N_10336);
and U10704 (N_10704,N_10489,N_10429);
xor U10705 (N_10705,N_10382,N_10317);
xor U10706 (N_10706,N_10415,N_10423);
or U10707 (N_10707,N_10485,N_10479);
nor U10708 (N_10708,N_10465,N_10493);
or U10709 (N_10709,N_10392,N_10489);
nand U10710 (N_10710,N_10368,N_10434);
nand U10711 (N_10711,N_10315,N_10464);
nand U10712 (N_10712,N_10355,N_10357);
and U10713 (N_10713,N_10395,N_10468);
xor U10714 (N_10714,N_10299,N_10308);
or U10715 (N_10715,N_10260,N_10377);
xnor U10716 (N_10716,N_10355,N_10414);
xor U10717 (N_10717,N_10342,N_10286);
xnor U10718 (N_10718,N_10380,N_10487);
nand U10719 (N_10719,N_10315,N_10395);
nand U10720 (N_10720,N_10337,N_10333);
or U10721 (N_10721,N_10264,N_10424);
nor U10722 (N_10722,N_10312,N_10418);
xnor U10723 (N_10723,N_10334,N_10363);
nand U10724 (N_10724,N_10316,N_10257);
nand U10725 (N_10725,N_10297,N_10313);
nand U10726 (N_10726,N_10499,N_10336);
nand U10727 (N_10727,N_10284,N_10260);
or U10728 (N_10728,N_10440,N_10391);
nor U10729 (N_10729,N_10354,N_10446);
xor U10730 (N_10730,N_10297,N_10497);
and U10731 (N_10731,N_10360,N_10351);
xor U10732 (N_10732,N_10440,N_10457);
or U10733 (N_10733,N_10317,N_10283);
and U10734 (N_10734,N_10399,N_10296);
nand U10735 (N_10735,N_10410,N_10442);
and U10736 (N_10736,N_10314,N_10387);
xnor U10737 (N_10737,N_10490,N_10319);
xor U10738 (N_10738,N_10253,N_10371);
xor U10739 (N_10739,N_10283,N_10355);
xor U10740 (N_10740,N_10455,N_10297);
xnor U10741 (N_10741,N_10394,N_10466);
nor U10742 (N_10742,N_10310,N_10265);
nor U10743 (N_10743,N_10428,N_10370);
and U10744 (N_10744,N_10482,N_10406);
xnor U10745 (N_10745,N_10321,N_10370);
or U10746 (N_10746,N_10432,N_10476);
nor U10747 (N_10747,N_10328,N_10273);
and U10748 (N_10748,N_10475,N_10450);
nor U10749 (N_10749,N_10453,N_10291);
or U10750 (N_10750,N_10598,N_10621);
nand U10751 (N_10751,N_10741,N_10556);
nand U10752 (N_10752,N_10716,N_10600);
and U10753 (N_10753,N_10531,N_10591);
or U10754 (N_10754,N_10667,N_10659);
and U10755 (N_10755,N_10589,N_10523);
and U10756 (N_10756,N_10625,N_10564);
or U10757 (N_10757,N_10525,N_10609);
xnor U10758 (N_10758,N_10677,N_10634);
nand U10759 (N_10759,N_10554,N_10595);
or U10760 (N_10760,N_10522,N_10666);
and U10761 (N_10761,N_10669,N_10579);
or U10762 (N_10762,N_10570,N_10652);
and U10763 (N_10763,N_10636,N_10664);
and U10764 (N_10764,N_10720,N_10562);
nor U10765 (N_10765,N_10673,N_10614);
or U10766 (N_10766,N_10628,N_10653);
and U10767 (N_10767,N_10566,N_10644);
nand U10768 (N_10768,N_10739,N_10622);
or U10769 (N_10769,N_10722,N_10578);
or U10770 (N_10770,N_10727,N_10708);
and U10771 (N_10771,N_10646,N_10545);
nand U10772 (N_10772,N_10701,N_10641);
and U10773 (N_10773,N_10707,N_10640);
or U10774 (N_10774,N_10599,N_10738);
and U10775 (N_10775,N_10699,N_10631);
and U10776 (N_10776,N_10513,N_10713);
nor U10777 (N_10777,N_10553,N_10530);
xor U10778 (N_10778,N_10617,N_10607);
and U10779 (N_10779,N_10558,N_10700);
and U10780 (N_10780,N_10696,N_10529);
nand U10781 (N_10781,N_10729,N_10674);
nand U10782 (N_10782,N_10593,N_10507);
or U10783 (N_10783,N_10612,N_10683);
or U10784 (N_10784,N_10662,N_10635);
or U10785 (N_10785,N_10538,N_10611);
and U10786 (N_10786,N_10670,N_10509);
or U10787 (N_10787,N_10528,N_10671);
or U10788 (N_10788,N_10505,N_10527);
nor U10789 (N_10789,N_10504,N_10552);
nand U10790 (N_10790,N_10569,N_10630);
and U10791 (N_10791,N_10603,N_10655);
or U10792 (N_10792,N_10637,N_10524);
and U10793 (N_10793,N_10592,N_10660);
and U10794 (N_10794,N_10686,N_10503);
nor U10795 (N_10795,N_10742,N_10672);
and U10796 (N_10796,N_10691,N_10502);
nand U10797 (N_10797,N_10689,N_10585);
or U10798 (N_10798,N_10731,N_10687);
nand U10799 (N_10799,N_10560,N_10732);
and U10800 (N_10800,N_10705,N_10661);
xnor U10801 (N_10801,N_10688,N_10548);
and U10802 (N_10802,N_10717,N_10718);
xnor U10803 (N_10803,N_10620,N_10702);
and U10804 (N_10804,N_10594,N_10535);
xnor U10805 (N_10805,N_10526,N_10656);
nor U10806 (N_10806,N_10645,N_10737);
or U10807 (N_10807,N_10643,N_10521);
xnor U10808 (N_10808,N_10561,N_10623);
and U10809 (N_10809,N_10719,N_10508);
and U10810 (N_10810,N_10710,N_10574);
or U10811 (N_10811,N_10632,N_10582);
and U10812 (N_10812,N_10565,N_10580);
or U10813 (N_10813,N_10743,N_10544);
or U10814 (N_10814,N_10735,N_10694);
and U10815 (N_10815,N_10546,N_10519);
xor U10816 (N_10816,N_10734,N_10557);
or U10817 (N_10817,N_10706,N_10629);
or U10818 (N_10818,N_10648,N_10744);
nor U10819 (N_10819,N_10668,N_10541);
xnor U10820 (N_10820,N_10539,N_10511);
nand U10821 (N_10821,N_10746,N_10606);
xor U10822 (N_10822,N_10638,N_10533);
nor U10823 (N_10823,N_10610,N_10559);
nand U10824 (N_10824,N_10692,N_10571);
nand U10825 (N_10825,N_10748,N_10682);
or U10826 (N_10826,N_10602,N_10517);
xnor U10827 (N_10827,N_10711,N_10730);
xnor U10828 (N_10828,N_10568,N_10726);
nand U10829 (N_10829,N_10615,N_10601);
and U10830 (N_10830,N_10654,N_10676);
and U10831 (N_10831,N_10551,N_10681);
nor U10832 (N_10832,N_10584,N_10572);
or U10833 (N_10833,N_10650,N_10693);
xor U10834 (N_10834,N_10613,N_10736);
nor U10835 (N_10835,N_10678,N_10555);
or U10836 (N_10836,N_10583,N_10532);
nor U10837 (N_10837,N_10596,N_10684);
and U10838 (N_10838,N_10604,N_10675);
and U10839 (N_10839,N_10709,N_10588);
nor U10840 (N_10840,N_10724,N_10616);
nor U10841 (N_10841,N_10590,N_10658);
nor U10842 (N_10842,N_10577,N_10714);
nor U10843 (N_10843,N_10639,N_10690);
and U10844 (N_10844,N_10704,N_10506);
nor U10845 (N_10845,N_10685,N_10633);
xnor U10846 (N_10846,N_10663,N_10665);
or U10847 (N_10847,N_10518,N_10728);
nand U10848 (N_10848,N_10597,N_10510);
nor U10849 (N_10849,N_10581,N_10725);
and U10850 (N_10850,N_10651,N_10550);
or U10851 (N_10851,N_10520,N_10624);
xor U10852 (N_10852,N_10586,N_10703);
and U10853 (N_10853,N_10647,N_10501);
nor U10854 (N_10854,N_10712,N_10549);
nand U10855 (N_10855,N_10642,N_10547);
nor U10856 (N_10856,N_10745,N_10567);
xor U10857 (N_10857,N_10747,N_10576);
and U10858 (N_10858,N_10680,N_10516);
xnor U10859 (N_10859,N_10512,N_10697);
nand U10860 (N_10860,N_10587,N_10515);
nor U10861 (N_10861,N_10540,N_10542);
or U10862 (N_10862,N_10698,N_10679);
nor U10863 (N_10863,N_10721,N_10605);
xor U10864 (N_10864,N_10537,N_10608);
nor U10865 (N_10865,N_10626,N_10627);
nand U10866 (N_10866,N_10575,N_10500);
xor U10867 (N_10867,N_10618,N_10563);
nor U10868 (N_10868,N_10657,N_10514);
nand U10869 (N_10869,N_10695,N_10536);
nor U10870 (N_10870,N_10715,N_10543);
or U10871 (N_10871,N_10619,N_10534);
xnor U10872 (N_10872,N_10573,N_10723);
xor U10873 (N_10873,N_10733,N_10649);
nand U10874 (N_10874,N_10749,N_10740);
xor U10875 (N_10875,N_10518,N_10703);
xnor U10876 (N_10876,N_10635,N_10656);
xor U10877 (N_10877,N_10536,N_10553);
nand U10878 (N_10878,N_10607,N_10736);
xnor U10879 (N_10879,N_10635,N_10652);
xnor U10880 (N_10880,N_10739,N_10666);
nor U10881 (N_10881,N_10646,N_10579);
nand U10882 (N_10882,N_10564,N_10728);
nor U10883 (N_10883,N_10562,N_10560);
nand U10884 (N_10884,N_10662,N_10596);
and U10885 (N_10885,N_10737,N_10599);
and U10886 (N_10886,N_10572,N_10588);
or U10887 (N_10887,N_10710,N_10582);
xor U10888 (N_10888,N_10604,N_10548);
and U10889 (N_10889,N_10695,N_10572);
and U10890 (N_10890,N_10584,N_10594);
or U10891 (N_10891,N_10689,N_10588);
or U10892 (N_10892,N_10598,N_10738);
nand U10893 (N_10893,N_10651,N_10542);
nand U10894 (N_10894,N_10700,N_10626);
and U10895 (N_10895,N_10638,N_10717);
xor U10896 (N_10896,N_10551,N_10675);
nor U10897 (N_10897,N_10560,N_10726);
nand U10898 (N_10898,N_10721,N_10636);
nor U10899 (N_10899,N_10573,N_10641);
xnor U10900 (N_10900,N_10514,N_10726);
nand U10901 (N_10901,N_10576,N_10671);
or U10902 (N_10902,N_10503,N_10707);
nand U10903 (N_10903,N_10577,N_10703);
xnor U10904 (N_10904,N_10555,N_10724);
xor U10905 (N_10905,N_10603,N_10563);
or U10906 (N_10906,N_10677,N_10663);
and U10907 (N_10907,N_10532,N_10626);
or U10908 (N_10908,N_10548,N_10590);
and U10909 (N_10909,N_10743,N_10538);
nor U10910 (N_10910,N_10574,N_10741);
nand U10911 (N_10911,N_10543,N_10545);
nor U10912 (N_10912,N_10582,N_10592);
xnor U10913 (N_10913,N_10513,N_10706);
nor U10914 (N_10914,N_10615,N_10729);
nor U10915 (N_10915,N_10541,N_10561);
or U10916 (N_10916,N_10545,N_10701);
and U10917 (N_10917,N_10656,N_10528);
xor U10918 (N_10918,N_10740,N_10636);
xor U10919 (N_10919,N_10739,N_10561);
or U10920 (N_10920,N_10631,N_10538);
and U10921 (N_10921,N_10706,N_10734);
nand U10922 (N_10922,N_10685,N_10728);
nor U10923 (N_10923,N_10535,N_10707);
and U10924 (N_10924,N_10500,N_10551);
and U10925 (N_10925,N_10621,N_10651);
or U10926 (N_10926,N_10598,N_10667);
nor U10927 (N_10927,N_10616,N_10505);
nand U10928 (N_10928,N_10716,N_10690);
and U10929 (N_10929,N_10554,N_10710);
xnor U10930 (N_10930,N_10690,N_10685);
and U10931 (N_10931,N_10595,N_10669);
and U10932 (N_10932,N_10574,N_10678);
nand U10933 (N_10933,N_10622,N_10534);
nor U10934 (N_10934,N_10560,N_10646);
and U10935 (N_10935,N_10589,N_10560);
xor U10936 (N_10936,N_10603,N_10626);
and U10937 (N_10937,N_10574,N_10521);
xnor U10938 (N_10938,N_10621,N_10724);
nor U10939 (N_10939,N_10687,N_10630);
or U10940 (N_10940,N_10601,N_10575);
or U10941 (N_10941,N_10709,N_10516);
or U10942 (N_10942,N_10529,N_10740);
xnor U10943 (N_10943,N_10520,N_10729);
nor U10944 (N_10944,N_10612,N_10730);
and U10945 (N_10945,N_10602,N_10553);
and U10946 (N_10946,N_10696,N_10646);
nor U10947 (N_10947,N_10634,N_10553);
or U10948 (N_10948,N_10558,N_10687);
nand U10949 (N_10949,N_10671,N_10511);
nor U10950 (N_10950,N_10524,N_10536);
xnor U10951 (N_10951,N_10638,N_10683);
or U10952 (N_10952,N_10741,N_10583);
nand U10953 (N_10953,N_10691,N_10504);
and U10954 (N_10954,N_10666,N_10672);
nand U10955 (N_10955,N_10543,N_10633);
or U10956 (N_10956,N_10668,N_10691);
or U10957 (N_10957,N_10733,N_10749);
nand U10958 (N_10958,N_10521,N_10640);
xnor U10959 (N_10959,N_10619,N_10593);
and U10960 (N_10960,N_10667,N_10619);
and U10961 (N_10961,N_10739,N_10742);
nor U10962 (N_10962,N_10718,N_10588);
xnor U10963 (N_10963,N_10524,N_10542);
nor U10964 (N_10964,N_10636,N_10676);
nand U10965 (N_10965,N_10695,N_10612);
xnor U10966 (N_10966,N_10609,N_10702);
xor U10967 (N_10967,N_10541,N_10577);
or U10968 (N_10968,N_10709,N_10511);
or U10969 (N_10969,N_10592,N_10713);
nand U10970 (N_10970,N_10727,N_10642);
xor U10971 (N_10971,N_10521,N_10675);
nor U10972 (N_10972,N_10587,N_10612);
xor U10973 (N_10973,N_10548,N_10684);
nand U10974 (N_10974,N_10543,N_10680);
or U10975 (N_10975,N_10631,N_10523);
nor U10976 (N_10976,N_10635,N_10692);
and U10977 (N_10977,N_10740,N_10589);
nand U10978 (N_10978,N_10572,N_10644);
and U10979 (N_10979,N_10686,N_10533);
xnor U10980 (N_10980,N_10548,N_10586);
xnor U10981 (N_10981,N_10516,N_10747);
xor U10982 (N_10982,N_10688,N_10545);
or U10983 (N_10983,N_10722,N_10559);
and U10984 (N_10984,N_10567,N_10748);
and U10985 (N_10985,N_10712,N_10507);
nand U10986 (N_10986,N_10501,N_10662);
nor U10987 (N_10987,N_10504,N_10683);
nand U10988 (N_10988,N_10593,N_10709);
or U10989 (N_10989,N_10672,N_10552);
nand U10990 (N_10990,N_10565,N_10619);
nor U10991 (N_10991,N_10642,N_10552);
or U10992 (N_10992,N_10518,N_10574);
nor U10993 (N_10993,N_10687,N_10662);
xnor U10994 (N_10994,N_10557,N_10632);
and U10995 (N_10995,N_10618,N_10580);
xor U10996 (N_10996,N_10622,N_10584);
and U10997 (N_10997,N_10519,N_10733);
or U10998 (N_10998,N_10625,N_10747);
and U10999 (N_10999,N_10621,N_10747);
xor U11000 (N_11000,N_10860,N_10903);
xnor U11001 (N_11001,N_10872,N_10871);
and U11002 (N_11002,N_10964,N_10882);
and U11003 (N_11003,N_10795,N_10974);
nand U11004 (N_11004,N_10932,N_10891);
or U11005 (N_11005,N_10951,N_10784);
and U11006 (N_11006,N_10815,N_10848);
nor U11007 (N_11007,N_10802,N_10855);
nand U11008 (N_11008,N_10813,N_10896);
nand U11009 (N_11009,N_10763,N_10806);
or U11010 (N_11010,N_10790,N_10949);
nor U11011 (N_11011,N_10805,N_10983);
nor U11012 (N_11012,N_10793,N_10809);
or U11013 (N_11013,N_10847,N_10846);
nor U11014 (N_11014,N_10935,N_10913);
nor U11015 (N_11015,N_10971,N_10826);
and U11016 (N_11016,N_10936,N_10839);
nand U11017 (N_11017,N_10859,N_10842);
nor U11018 (N_11018,N_10812,N_10844);
and U11019 (N_11019,N_10828,N_10798);
or U11020 (N_11020,N_10760,N_10782);
xor U11021 (N_11021,N_10781,N_10771);
or U11022 (N_11022,N_10814,N_10969);
xnor U11023 (N_11023,N_10884,N_10909);
or U11024 (N_11024,N_10888,N_10779);
xnor U11025 (N_11025,N_10856,N_10948);
nand U11026 (N_11026,N_10868,N_10989);
or U11027 (N_11027,N_10980,N_10845);
and U11028 (N_11028,N_10901,N_10907);
nand U11029 (N_11029,N_10934,N_10941);
or U11030 (N_11030,N_10968,N_10945);
nor U11031 (N_11031,N_10776,N_10836);
nand U11032 (N_11032,N_10834,N_10905);
xor U11033 (N_11033,N_10791,N_10774);
and U11034 (N_11034,N_10926,N_10900);
or U11035 (N_11035,N_10958,N_10800);
nand U11036 (N_11036,N_10962,N_10754);
nor U11037 (N_11037,N_10906,N_10981);
or U11038 (N_11038,N_10916,N_10887);
or U11039 (N_11039,N_10881,N_10994);
and U11040 (N_11040,N_10870,N_10915);
nor U11041 (N_11041,N_10973,N_10944);
nand U11042 (N_11042,N_10991,N_10825);
or U11043 (N_11043,N_10979,N_10765);
or U11044 (N_11044,N_10820,N_10853);
nor U11045 (N_11045,N_10922,N_10761);
nand U11046 (N_11046,N_10878,N_10823);
or U11047 (N_11047,N_10879,N_10863);
nand U11048 (N_11048,N_10854,N_10975);
xor U11049 (N_11049,N_10827,N_10972);
nor U11050 (N_11050,N_10775,N_10942);
nand U11051 (N_11051,N_10840,N_10889);
nand U11052 (N_11052,N_10957,N_10996);
or U11053 (N_11053,N_10822,N_10985);
nand U11054 (N_11054,N_10965,N_10769);
xor U11055 (N_11055,N_10787,N_10966);
nand U11056 (N_11056,N_10986,N_10877);
nor U11057 (N_11057,N_10780,N_10833);
and U11058 (N_11058,N_10954,N_10824);
nor U11059 (N_11059,N_10757,N_10858);
or U11060 (N_11060,N_10939,N_10883);
nand U11061 (N_11061,N_10838,N_10999);
nand U11062 (N_11062,N_10869,N_10947);
and U11063 (N_11063,N_10910,N_10931);
xor U11064 (N_11064,N_10912,N_10788);
nor U11065 (N_11065,N_10899,N_10865);
nand U11066 (N_11066,N_10946,N_10908);
nor U11067 (N_11067,N_10866,N_10914);
xor U11068 (N_11068,N_10956,N_10921);
or U11069 (N_11069,N_10799,N_10759);
nor U11070 (N_11070,N_10904,N_10995);
or U11071 (N_11071,N_10857,N_10753);
xnor U11072 (N_11072,N_10928,N_10778);
nand U11073 (N_11073,N_10864,N_10953);
nand U11074 (N_11074,N_10880,N_10886);
nand U11075 (N_11075,N_10758,N_10917);
nor U11076 (N_11076,N_10762,N_10938);
or U11077 (N_11077,N_10923,N_10821);
nand U11078 (N_11078,N_10930,N_10849);
or U11079 (N_11079,N_10893,N_10750);
nor U11080 (N_11080,N_10851,N_10919);
and U11081 (N_11081,N_10783,N_10818);
xor U11082 (N_11082,N_10770,N_10885);
and U11083 (N_11083,N_10876,N_10786);
nand U11084 (N_11084,N_10873,N_10852);
and U11085 (N_11085,N_10829,N_10803);
and U11086 (N_11086,N_10797,N_10807);
xnor U11087 (N_11087,N_10993,N_10929);
xor U11088 (N_11088,N_10832,N_10998);
xor U11089 (N_11089,N_10796,N_10772);
nor U11090 (N_11090,N_10943,N_10959);
nor U11091 (N_11091,N_10777,N_10940);
or U11092 (N_11092,N_10927,N_10835);
and U11093 (N_11093,N_10955,N_10816);
and U11094 (N_11094,N_10911,N_10830);
and U11095 (N_11095,N_10984,N_10850);
xor U11096 (N_11096,N_10920,N_10895);
xnor U11097 (N_11097,N_10841,N_10918);
nand U11098 (N_11098,N_10801,N_10867);
xnor U11099 (N_11099,N_10794,N_10768);
nand U11100 (N_11100,N_10766,N_10961);
nand U11101 (N_11101,N_10756,N_10764);
or U11102 (N_11102,N_10898,N_10752);
nor U11103 (N_11103,N_10890,N_10819);
and U11104 (N_11104,N_10804,N_10875);
and U11105 (N_11105,N_10789,N_10937);
or U11106 (N_11106,N_10963,N_10755);
nor U11107 (N_11107,N_10960,N_10987);
nand U11108 (N_11108,N_10976,N_10924);
nor U11109 (N_11109,N_10933,N_10952);
and U11110 (N_11110,N_10902,N_10831);
and U11111 (N_11111,N_10817,N_10892);
nor U11112 (N_11112,N_10767,N_10843);
xnor U11113 (N_11113,N_10977,N_10773);
xnor U11114 (N_11114,N_10950,N_10978);
and U11115 (N_11115,N_10874,N_10990);
nand U11116 (N_11116,N_10861,N_10967);
or U11117 (N_11117,N_10810,N_10811);
nand U11118 (N_11118,N_10862,N_10837);
or U11119 (N_11119,N_10970,N_10992);
xor U11120 (N_11120,N_10792,N_10897);
nand U11121 (N_11121,N_10785,N_10808);
or U11122 (N_11122,N_10925,N_10751);
xnor U11123 (N_11123,N_10982,N_10894);
and U11124 (N_11124,N_10997,N_10988);
nor U11125 (N_11125,N_10861,N_10791);
or U11126 (N_11126,N_10753,N_10835);
xnor U11127 (N_11127,N_10772,N_10962);
xor U11128 (N_11128,N_10762,N_10790);
nand U11129 (N_11129,N_10852,N_10999);
and U11130 (N_11130,N_10815,N_10864);
nor U11131 (N_11131,N_10946,N_10836);
xor U11132 (N_11132,N_10864,N_10965);
nor U11133 (N_11133,N_10804,N_10896);
xor U11134 (N_11134,N_10889,N_10763);
nand U11135 (N_11135,N_10885,N_10830);
or U11136 (N_11136,N_10808,N_10815);
nor U11137 (N_11137,N_10902,N_10852);
or U11138 (N_11138,N_10846,N_10886);
and U11139 (N_11139,N_10880,N_10798);
or U11140 (N_11140,N_10949,N_10978);
and U11141 (N_11141,N_10850,N_10794);
nor U11142 (N_11142,N_10965,N_10846);
nand U11143 (N_11143,N_10859,N_10941);
nand U11144 (N_11144,N_10849,N_10892);
and U11145 (N_11145,N_10756,N_10841);
and U11146 (N_11146,N_10779,N_10913);
or U11147 (N_11147,N_10928,N_10970);
nand U11148 (N_11148,N_10873,N_10921);
or U11149 (N_11149,N_10987,N_10884);
xor U11150 (N_11150,N_10880,N_10800);
or U11151 (N_11151,N_10761,N_10878);
or U11152 (N_11152,N_10873,N_10761);
or U11153 (N_11153,N_10954,N_10794);
nand U11154 (N_11154,N_10788,N_10950);
nor U11155 (N_11155,N_10764,N_10979);
and U11156 (N_11156,N_10998,N_10861);
xor U11157 (N_11157,N_10907,N_10828);
nand U11158 (N_11158,N_10764,N_10985);
and U11159 (N_11159,N_10846,N_10871);
nor U11160 (N_11160,N_10764,N_10837);
and U11161 (N_11161,N_10866,N_10861);
and U11162 (N_11162,N_10894,N_10834);
and U11163 (N_11163,N_10887,N_10918);
xor U11164 (N_11164,N_10963,N_10987);
or U11165 (N_11165,N_10853,N_10985);
xor U11166 (N_11166,N_10823,N_10821);
and U11167 (N_11167,N_10756,N_10900);
nor U11168 (N_11168,N_10907,N_10848);
and U11169 (N_11169,N_10919,N_10811);
nor U11170 (N_11170,N_10885,N_10971);
nand U11171 (N_11171,N_10761,N_10942);
nand U11172 (N_11172,N_10930,N_10785);
nand U11173 (N_11173,N_10808,N_10756);
nor U11174 (N_11174,N_10829,N_10995);
nor U11175 (N_11175,N_10913,N_10978);
and U11176 (N_11176,N_10759,N_10965);
or U11177 (N_11177,N_10952,N_10759);
xor U11178 (N_11178,N_10973,N_10774);
nor U11179 (N_11179,N_10784,N_10892);
nand U11180 (N_11180,N_10796,N_10923);
nand U11181 (N_11181,N_10888,N_10799);
nor U11182 (N_11182,N_10975,N_10762);
nor U11183 (N_11183,N_10929,N_10838);
or U11184 (N_11184,N_10795,N_10856);
and U11185 (N_11185,N_10777,N_10950);
nor U11186 (N_11186,N_10880,N_10839);
and U11187 (N_11187,N_10779,N_10865);
and U11188 (N_11188,N_10861,N_10812);
and U11189 (N_11189,N_10785,N_10873);
or U11190 (N_11190,N_10917,N_10776);
and U11191 (N_11191,N_10875,N_10985);
nand U11192 (N_11192,N_10850,N_10869);
or U11193 (N_11193,N_10906,N_10978);
and U11194 (N_11194,N_10944,N_10910);
or U11195 (N_11195,N_10754,N_10988);
nand U11196 (N_11196,N_10812,N_10881);
xor U11197 (N_11197,N_10756,N_10922);
xnor U11198 (N_11198,N_10771,N_10907);
and U11199 (N_11199,N_10894,N_10849);
or U11200 (N_11200,N_10759,N_10932);
and U11201 (N_11201,N_10819,N_10848);
and U11202 (N_11202,N_10842,N_10820);
and U11203 (N_11203,N_10781,N_10999);
nand U11204 (N_11204,N_10991,N_10890);
and U11205 (N_11205,N_10958,N_10872);
nand U11206 (N_11206,N_10814,N_10984);
xnor U11207 (N_11207,N_10825,N_10763);
and U11208 (N_11208,N_10886,N_10983);
and U11209 (N_11209,N_10870,N_10991);
nor U11210 (N_11210,N_10823,N_10974);
or U11211 (N_11211,N_10871,N_10960);
nor U11212 (N_11212,N_10819,N_10934);
and U11213 (N_11213,N_10897,N_10935);
xor U11214 (N_11214,N_10927,N_10762);
nand U11215 (N_11215,N_10934,N_10937);
nor U11216 (N_11216,N_10843,N_10846);
or U11217 (N_11217,N_10913,N_10771);
xnor U11218 (N_11218,N_10777,N_10837);
xnor U11219 (N_11219,N_10852,N_10764);
and U11220 (N_11220,N_10952,N_10816);
nand U11221 (N_11221,N_10804,N_10845);
or U11222 (N_11222,N_10765,N_10850);
xnor U11223 (N_11223,N_10949,N_10928);
xnor U11224 (N_11224,N_10882,N_10864);
nor U11225 (N_11225,N_10806,N_10981);
xnor U11226 (N_11226,N_10838,N_10757);
xnor U11227 (N_11227,N_10825,N_10847);
xor U11228 (N_11228,N_10955,N_10826);
or U11229 (N_11229,N_10806,N_10910);
xor U11230 (N_11230,N_10994,N_10977);
nand U11231 (N_11231,N_10925,N_10788);
and U11232 (N_11232,N_10813,N_10908);
xor U11233 (N_11233,N_10784,N_10880);
nand U11234 (N_11234,N_10822,N_10934);
xnor U11235 (N_11235,N_10825,N_10858);
or U11236 (N_11236,N_10887,N_10751);
xnor U11237 (N_11237,N_10923,N_10802);
xnor U11238 (N_11238,N_10976,N_10836);
and U11239 (N_11239,N_10884,N_10949);
xnor U11240 (N_11240,N_10919,N_10910);
or U11241 (N_11241,N_10766,N_10858);
and U11242 (N_11242,N_10873,N_10913);
and U11243 (N_11243,N_10796,N_10760);
or U11244 (N_11244,N_10806,N_10874);
nand U11245 (N_11245,N_10919,N_10953);
xnor U11246 (N_11246,N_10796,N_10914);
and U11247 (N_11247,N_10998,N_10888);
or U11248 (N_11248,N_10797,N_10949);
and U11249 (N_11249,N_10879,N_10900);
and U11250 (N_11250,N_11189,N_11070);
nand U11251 (N_11251,N_11209,N_11107);
nor U11252 (N_11252,N_11220,N_11001);
and U11253 (N_11253,N_11062,N_11112);
nor U11254 (N_11254,N_11221,N_11009);
nand U11255 (N_11255,N_11206,N_11030);
or U11256 (N_11256,N_11139,N_11008);
and U11257 (N_11257,N_11077,N_11205);
or U11258 (N_11258,N_11047,N_11126);
and U11259 (N_11259,N_11174,N_11129);
nor U11260 (N_11260,N_11188,N_11146);
xor U11261 (N_11261,N_11104,N_11054);
or U11262 (N_11262,N_11121,N_11072);
xnor U11263 (N_11263,N_11236,N_11076);
and U11264 (N_11264,N_11110,N_11242);
nor U11265 (N_11265,N_11195,N_11246);
nand U11266 (N_11266,N_11217,N_11010);
and U11267 (N_11267,N_11198,N_11184);
or U11268 (N_11268,N_11004,N_11153);
or U11269 (N_11269,N_11194,N_11210);
and U11270 (N_11270,N_11080,N_11244);
or U11271 (N_11271,N_11154,N_11237);
nor U11272 (N_11272,N_11056,N_11171);
xor U11273 (N_11273,N_11187,N_11045);
xor U11274 (N_11274,N_11101,N_11093);
or U11275 (N_11275,N_11224,N_11181);
or U11276 (N_11276,N_11197,N_11203);
and U11277 (N_11277,N_11175,N_11068);
nor U11278 (N_11278,N_11131,N_11167);
nor U11279 (N_11279,N_11243,N_11088);
or U11280 (N_11280,N_11018,N_11212);
or U11281 (N_11281,N_11202,N_11102);
nor U11282 (N_11282,N_11169,N_11066);
or U11283 (N_11283,N_11057,N_11151);
nand U11284 (N_11284,N_11035,N_11214);
nor U11285 (N_11285,N_11159,N_11114);
or U11286 (N_11286,N_11186,N_11204);
nand U11287 (N_11287,N_11097,N_11065);
and U11288 (N_11288,N_11201,N_11191);
and U11289 (N_11289,N_11133,N_11061);
or U11290 (N_11290,N_11003,N_11240);
xnor U11291 (N_11291,N_11041,N_11043);
xor U11292 (N_11292,N_11135,N_11157);
and U11293 (N_11293,N_11156,N_11039);
and U11294 (N_11294,N_11006,N_11090);
xnor U11295 (N_11295,N_11170,N_11031);
or U11296 (N_11296,N_11058,N_11111);
xor U11297 (N_11297,N_11032,N_11147);
nand U11298 (N_11298,N_11122,N_11150);
or U11299 (N_11299,N_11091,N_11231);
nand U11300 (N_11300,N_11086,N_11094);
xor U11301 (N_11301,N_11048,N_11109);
xnor U11302 (N_11302,N_11075,N_11046);
nand U11303 (N_11303,N_11179,N_11207);
and U11304 (N_11304,N_11143,N_11005);
nand U11305 (N_11305,N_11245,N_11084);
xor U11306 (N_11306,N_11222,N_11116);
nor U11307 (N_11307,N_11023,N_11185);
or U11308 (N_11308,N_11038,N_11160);
and U11309 (N_11309,N_11149,N_11055);
nand U11310 (N_11310,N_11002,N_11083);
or U11311 (N_11311,N_11248,N_11168);
or U11312 (N_11312,N_11063,N_11176);
or U11313 (N_11313,N_11108,N_11087);
or U11314 (N_11314,N_11162,N_11022);
and U11315 (N_11315,N_11105,N_11016);
nor U11316 (N_11316,N_11200,N_11144);
xnor U11317 (N_11317,N_11098,N_11042);
or U11318 (N_11318,N_11155,N_11029);
or U11319 (N_11319,N_11025,N_11044);
or U11320 (N_11320,N_11128,N_11113);
and U11321 (N_11321,N_11225,N_11082);
nand U11322 (N_11322,N_11040,N_11074);
nor U11323 (N_11323,N_11099,N_11213);
and U11324 (N_11324,N_11036,N_11199);
and U11325 (N_11325,N_11148,N_11052);
xor U11326 (N_11326,N_11081,N_11064);
nand U11327 (N_11327,N_11223,N_11019);
xnor U11328 (N_11328,N_11232,N_11172);
nor U11329 (N_11329,N_11049,N_11123);
xor U11330 (N_11330,N_11218,N_11132);
xor U11331 (N_11331,N_11024,N_11078);
nor U11332 (N_11332,N_11247,N_11051);
or U11333 (N_11333,N_11130,N_11161);
xor U11334 (N_11334,N_11060,N_11117);
xor U11335 (N_11335,N_11115,N_11000);
xor U11336 (N_11336,N_11228,N_11011);
or U11337 (N_11337,N_11014,N_11124);
nor U11338 (N_11338,N_11092,N_11141);
xor U11339 (N_11339,N_11026,N_11028);
and U11340 (N_11340,N_11208,N_11020);
or U11341 (N_11341,N_11069,N_11182);
and U11342 (N_11342,N_11089,N_11053);
xnor U11343 (N_11343,N_11071,N_11137);
or U11344 (N_11344,N_11178,N_11096);
nand U11345 (N_11345,N_11226,N_11079);
and U11346 (N_11346,N_11230,N_11012);
nor U11347 (N_11347,N_11067,N_11166);
nand U11348 (N_11348,N_11152,N_11190);
and U11349 (N_11349,N_11229,N_11100);
or U11350 (N_11350,N_11196,N_11033);
xnor U11351 (N_11351,N_11106,N_11120);
or U11352 (N_11352,N_11050,N_11164);
xor U11353 (N_11353,N_11118,N_11215);
and U11354 (N_11354,N_11173,N_11125);
and U11355 (N_11355,N_11017,N_11233);
xor U11356 (N_11356,N_11216,N_11145);
and U11357 (N_11357,N_11219,N_11021);
xnor U11358 (N_11358,N_11180,N_11027);
xor U11359 (N_11359,N_11193,N_11163);
and U11360 (N_11360,N_11158,N_11138);
or U11361 (N_11361,N_11095,N_11142);
and U11362 (N_11362,N_11059,N_11183);
xnor U11363 (N_11363,N_11238,N_11103);
nand U11364 (N_11364,N_11127,N_11136);
and U11365 (N_11365,N_11140,N_11073);
xor U11366 (N_11366,N_11015,N_11235);
or U11367 (N_11367,N_11134,N_11037);
nor U11368 (N_11368,N_11119,N_11034);
and U11369 (N_11369,N_11165,N_11013);
or U11370 (N_11370,N_11192,N_11239);
xor U11371 (N_11371,N_11211,N_11249);
nor U11372 (N_11372,N_11085,N_11241);
nand U11373 (N_11373,N_11227,N_11234);
xnor U11374 (N_11374,N_11007,N_11177);
nand U11375 (N_11375,N_11070,N_11058);
nor U11376 (N_11376,N_11114,N_11144);
or U11377 (N_11377,N_11158,N_11121);
xnor U11378 (N_11378,N_11151,N_11055);
nor U11379 (N_11379,N_11083,N_11041);
xnor U11380 (N_11380,N_11040,N_11042);
nand U11381 (N_11381,N_11173,N_11019);
xor U11382 (N_11382,N_11188,N_11160);
nor U11383 (N_11383,N_11077,N_11174);
or U11384 (N_11384,N_11007,N_11238);
nor U11385 (N_11385,N_11001,N_11014);
xor U11386 (N_11386,N_11151,N_11201);
xor U11387 (N_11387,N_11013,N_11105);
or U11388 (N_11388,N_11184,N_11196);
nor U11389 (N_11389,N_11054,N_11141);
or U11390 (N_11390,N_11000,N_11201);
nand U11391 (N_11391,N_11172,N_11248);
and U11392 (N_11392,N_11028,N_11141);
nor U11393 (N_11393,N_11162,N_11242);
xnor U11394 (N_11394,N_11001,N_11174);
xnor U11395 (N_11395,N_11104,N_11225);
and U11396 (N_11396,N_11130,N_11168);
nand U11397 (N_11397,N_11216,N_11210);
xnor U11398 (N_11398,N_11128,N_11015);
nand U11399 (N_11399,N_11205,N_11128);
and U11400 (N_11400,N_11076,N_11249);
and U11401 (N_11401,N_11178,N_11148);
and U11402 (N_11402,N_11194,N_11226);
and U11403 (N_11403,N_11203,N_11186);
nand U11404 (N_11404,N_11192,N_11119);
xnor U11405 (N_11405,N_11183,N_11111);
and U11406 (N_11406,N_11127,N_11050);
or U11407 (N_11407,N_11141,N_11175);
or U11408 (N_11408,N_11162,N_11083);
xnor U11409 (N_11409,N_11018,N_11050);
and U11410 (N_11410,N_11124,N_11119);
nand U11411 (N_11411,N_11110,N_11167);
and U11412 (N_11412,N_11169,N_11004);
xnor U11413 (N_11413,N_11231,N_11147);
nand U11414 (N_11414,N_11206,N_11221);
or U11415 (N_11415,N_11078,N_11101);
and U11416 (N_11416,N_11212,N_11143);
or U11417 (N_11417,N_11213,N_11013);
and U11418 (N_11418,N_11189,N_11073);
nor U11419 (N_11419,N_11039,N_11000);
xor U11420 (N_11420,N_11102,N_11160);
nor U11421 (N_11421,N_11107,N_11168);
and U11422 (N_11422,N_11034,N_11097);
nor U11423 (N_11423,N_11130,N_11025);
xnor U11424 (N_11424,N_11231,N_11144);
or U11425 (N_11425,N_11161,N_11096);
xor U11426 (N_11426,N_11043,N_11212);
nor U11427 (N_11427,N_11081,N_11206);
and U11428 (N_11428,N_11110,N_11108);
xnor U11429 (N_11429,N_11057,N_11165);
nor U11430 (N_11430,N_11207,N_11042);
nor U11431 (N_11431,N_11109,N_11063);
or U11432 (N_11432,N_11248,N_11074);
nor U11433 (N_11433,N_11145,N_11211);
xnor U11434 (N_11434,N_11245,N_11131);
nor U11435 (N_11435,N_11040,N_11078);
nor U11436 (N_11436,N_11134,N_11214);
and U11437 (N_11437,N_11127,N_11196);
or U11438 (N_11438,N_11089,N_11184);
and U11439 (N_11439,N_11237,N_11246);
and U11440 (N_11440,N_11128,N_11141);
nor U11441 (N_11441,N_11227,N_11003);
nor U11442 (N_11442,N_11075,N_11119);
nor U11443 (N_11443,N_11040,N_11036);
nand U11444 (N_11444,N_11002,N_11080);
nand U11445 (N_11445,N_11023,N_11167);
or U11446 (N_11446,N_11111,N_11210);
and U11447 (N_11447,N_11190,N_11145);
and U11448 (N_11448,N_11073,N_11063);
or U11449 (N_11449,N_11075,N_11030);
or U11450 (N_11450,N_11199,N_11198);
and U11451 (N_11451,N_11069,N_11044);
or U11452 (N_11452,N_11115,N_11076);
and U11453 (N_11453,N_11068,N_11050);
and U11454 (N_11454,N_11193,N_11112);
xnor U11455 (N_11455,N_11123,N_11041);
and U11456 (N_11456,N_11097,N_11108);
and U11457 (N_11457,N_11245,N_11114);
nor U11458 (N_11458,N_11068,N_11126);
xor U11459 (N_11459,N_11244,N_11177);
xnor U11460 (N_11460,N_11019,N_11035);
nor U11461 (N_11461,N_11230,N_11041);
and U11462 (N_11462,N_11130,N_11201);
nand U11463 (N_11463,N_11158,N_11029);
and U11464 (N_11464,N_11127,N_11091);
xor U11465 (N_11465,N_11053,N_11112);
and U11466 (N_11466,N_11182,N_11187);
nor U11467 (N_11467,N_11190,N_11054);
or U11468 (N_11468,N_11014,N_11240);
nand U11469 (N_11469,N_11217,N_11119);
nand U11470 (N_11470,N_11056,N_11210);
and U11471 (N_11471,N_11132,N_11027);
or U11472 (N_11472,N_11190,N_11014);
nand U11473 (N_11473,N_11204,N_11061);
xor U11474 (N_11474,N_11040,N_11213);
xor U11475 (N_11475,N_11204,N_11003);
nand U11476 (N_11476,N_11246,N_11098);
and U11477 (N_11477,N_11154,N_11184);
nand U11478 (N_11478,N_11061,N_11034);
nor U11479 (N_11479,N_11006,N_11237);
nor U11480 (N_11480,N_11149,N_11042);
and U11481 (N_11481,N_11078,N_11067);
and U11482 (N_11482,N_11088,N_11099);
nor U11483 (N_11483,N_11146,N_11239);
nand U11484 (N_11484,N_11061,N_11000);
nand U11485 (N_11485,N_11058,N_11035);
nor U11486 (N_11486,N_11222,N_11195);
and U11487 (N_11487,N_11196,N_11025);
or U11488 (N_11488,N_11219,N_11083);
nor U11489 (N_11489,N_11077,N_11133);
and U11490 (N_11490,N_11004,N_11046);
or U11491 (N_11491,N_11096,N_11233);
xor U11492 (N_11492,N_11005,N_11017);
xor U11493 (N_11493,N_11177,N_11212);
or U11494 (N_11494,N_11066,N_11125);
or U11495 (N_11495,N_11194,N_11109);
and U11496 (N_11496,N_11104,N_11043);
nor U11497 (N_11497,N_11032,N_11013);
nor U11498 (N_11498,N_11075,N_11160);
or U11499 (N_11499,N_11215,N_11229);
nor U11500 (N_11500,N_11359,N_11365);
nand U11501 (N_11501,N_11258,N_11494);
or U11502 (N_11502,N_11256,N_11456);
and U11503 (N_11503,N_11399,N_11452);
nor U11504 (N_11504,N_11489,N_11486);
and U11505 (N_11505,N_11336,N_11372);
nand U11506 (N_11506,N_11259,N_11270);
and U11507 (N_11507,N_11279,N_11318);
and U11508 (N_11508,N_11269,N_11324);
xnor U11509 (N_11509,N_11471,N_11499);
nand U11510 (N_11510,N_11402,N_11331);
nor U11511 (N_11511,N_11454,N_11284);
xor U11512 (N_11512,N_11420,N_11470);
or U11513 (N_11513,N_11304,N_11341);
nor U11514 (N_11514,N_11350,N_11337);
nand U11515 (N_11515,N_11493,N_11488);
or U11516 (N_11516,N_11396,N_11382);
or U11517 (N_11517,N_11432,N_11498);
nand U11518 (N_11518,N_11340,N_11475);
nor U11519 (N_11519,N_11381,N_11332);
xnor U11520 (N_11520,N_11405,N_11363);
and U11521 (N_11521,N_11491,N_11444);
and U11522 (N_11522,N_11398,N_11303);
xnor U11523 (N_11523,N_11266,N_11410);
nand U11524 (N_11524,N_11423,N_11315);
or U11525 (N_11525,N_11282,N_11403);
or U11526 (N_11526,N_11301,N_11251);
or U11527 (N_11527,N_11474,N_11371);
nand U11528 (N_11528,N_11278,N_11309);
xnor U11529 (N_11529,N_11465,N_11264);
nor U11530 (N_11530,N_11280,N_11422);
nand U11531 (N_11531,N_11453,N_11307);
or U11532 (N_11532,N_11473,N_11352);
nor U11533 (N_11533,N_11438,N_11286);
nand U11534 (N_11534,N_11276,N_11373);
or U11535 (N_11535,N_11448,N_11364);
and U11536 (N_11536,N_11391,N_11380);
nor U11537 (N_11537,N_11415,N_11294);
xnor U11538 (N_11538,N_11356,N_11466);
nor U11539 (N_11539,N_11333,N_11479);
or U11540 (N_11540,N_11327,N_11329);
nand U11541 (N_11541,N_11457,N_11497);
nand U11542 (N_11542,N_11417,N_11369);
nand U11543 (N_11543,N_11435,N_11370);
or U11544 (N_11544,N_11418,N_11482);
nand U11545 (N_11545,N_11468,N_11260);
nor U11546 (N_11546,N_11425,N_11358);
xor U11547 (N_11547,N_11447,N_11262);
nand U11548 (N_11548,N_11414,N_11459);
nor U11549 (N_11549,N_11461,N_11384);
or U11550 (N_11550,N_11427,N_11443);
and U11551 (N_11551,N_11411,N_11311);
or U11552 (N_11552,N_11317,N_11416);
xor U11553 (N_11553,N_11374,N_11393);
nand U11554 (N_11554,N_11330,N_11496);
nand U11555 (N_11555,N_11290,N_11334);
or U11556 (N_11556,N_11263,N_11426);
and U11557 (N_11557,N_11492,N_11409);
nand U11558 (N_11558,N_11392,N_11406);
xor U11559 (N_11559,N_11439,N_11419);
nand U11560 (N_11560,N_11275,N_11389);
or U11561 (N_11561,N_11395,N_11287);
nor U11562 (N_11562,N_11295,N_11344);
nor U11563 (N_11563,N_11285,N_11477);
nor U11564 (N_11564,N_11305,N_11430);
or U11565 (N_11565,N_11449,N_11351);
nor U11566 (N_11566,N_11267,N_11377);
and U11567 (N_11567,N_11292,N_11462);
nand U11568 (N_11568,N_11319,N_11478);
or U11569 (N_11569,N_11357,N_11273);
nand U11570 (N_11570,N_11272,N_11421);
xor U11571 (N_11571,N_11252,N_11431);
xor U11572 (N_11572,N_11366,N_11268);
or U11573 (N_11573,N_11480,N_11313);
and U11574 (N_11574,N_11451,N_11283);
xor U11575 (N_11575,N_11299,N_11361);
and U11576 (N_11576,N_11281,N_11433);
nand U11577 (N_11577,N_11345,N_11460);
and U11578 (N_11578,N_11441,N_11401);
xor U11579 (N_11579,N_11472,N_11436);
nand U11580 (N_11580,N_11490,N_11464);
and U11581 (N_11581,N_11469,N_11326);
xor U11582 (N_11582,N_11255,N_11310);
xor U11583 (N_11583,N_11434,N_11440);
xnor U11584 (N_11584,N_11306,N_11428);
xnor U11585 (N_11585,N_11288,N_11483);
nand U11586 (N_11586,N_11261,N_11348);
and U11587 (N_11587,N_11397,N_11376);
or U11588 (N_11588,N_11328,N_11323);
nor U11589 (N_11589,N_11298,N_11379);
or U11590 (N_11590,N_11322,N_11484);
or U11591 (N_11591,N_11346,N_11375);
xnor U11592 (N_11592,N_11387,N_11450);
xor U11593 (N_11593,N_11254,N_11293);
xnor U11594 (N_11594,N_11362,N_11343);
nand U11595 (N_11595,N_11400,N_11289);
xnor U11596 (N_11596,N_11442,N_11349);
or U11597 (N_11597,N_11386,N_11458);
nor U11598 (N_11598,N_11360,N_11388);
nand U11599 (N_11599,N_11412,N_11316);
or U11600 (N_11600,N_11320,N_11485);
nand U11601 (N_11601,N_11424,N_11445);
and U11602 (N_11602,N_11353,N_11312);
xnor U11603 (N_11603,N_11463,N_11495);
or U11604 (N_11604,N_11347,N_11277);
and U11605 (N_11605,N_11342,N_11476);
and U11606 (N_11606,N_11335,N_11429);
or U11607 (N_11607,N_11467,N_11297);
and U11608 (N_11608,N_11378,N_11437);
nor U11609 (N_11609,N_11339,N_11308);
nand U11610 (N_11610,N_11338,N_11354);
and U11611 (N_11611,N_11265,N_11253);
nor U11612 (N_11612,N_11408,N_11383);
nand U11613 (N_11613,N_11296,N_11257);
and U11614 (N_11614,N_11407,N_11274);
nor U11615 (N_11615,N_11271,N_11390);
xnor U11616 (N_11616,N_11446,N_11250);
nor U11617 (N_11617,N_11291,N_11487);
xnor U11618 (N_11618,N_11300,N_11321);
or U11619 (N_11619,N_11368,N_11455);
nand U11620 (N_11620,N_11325,N_11413);
and U11621 (N_11621,N_11355,N_11481);
or U11622 (N_11622,N_11394,N_11367);
or U11623 (N_11623,N_11314,N_11404);
and U11624 (N_11624,N_11302,N_11385);
and U11625 (N_11625,N_11274,N_11430);
and U11626 (N_11626,N_11413,N_11425);
xnor U11627 (N_11627,N_11423,N_11406);
nand U11628 (N_11628,N_11347,N_11457);
or U11629 (N_11629,N_11492,N_11283);
xor U11630 (N_11630,N_11470,N_11383);
or U11631 (N_11631,N_11432,N_11293);
nor U11632 (N_11632,N_11313,N_11419);
nor U11633 (N_11633,N_11299,N_11332);
xnor U11634 (N_11634,N_11254,N_11420);
and U11635 (N_11635,N_11309,N_11349);
nand U11636 (N_11636,N_11333,N_11252);
and U11637 (N_11637,N_11361,N_11452);
or U11638 (N_11638,N_11494,N_11296);
nor U11639 (N_11639,N_11376,N_11379);
and U11640 (N_11640,N_11460,N_11259);
nor U11641 (N_11641,N_11250,N_11372);
nor U11642 (N_11642,N_11374,N_11477);
nand U11643 (N_11643,N_11467,N_11489);
and U11644 (N_11644,N_11392,N_11496);
xnor U11645 (N_11645,N_11425,N_11312);
nand U11646 (N_11646,N_11499,N_11363);
or U11647 (N_11647,N_11419,N_11357);
xnor U11648 (N_11648,N_11285,N_11394);
and U11649 (N_11649,N_11355,N_11404);
nor U11650 (N_11650,N_11451,N_11475);
and U11651 (N_11651,N_11370,N_11362);
xnor U11652 (N_11652,N_11325,N_11415);
nor U11653 (N_11653,N_11332,N_11352);
xor U11654 (N_11654,N_11377,N_11324);
nor U11655 (N_11655,N_11485,N_11316);
and U11656 (N_11656,N_11444,N_11408);
nor U11657 (N_11657,N_11497,N_11326);
nand U11658 (N_11658,N_11368,N_11323);
xor U11659 (N_11659,N_11365,N_11333);
or U11660 (N_11660,N_11493,N_11402);
xnor U11661 (N_11661,N_11493,N_11293);
nand U11662 (N_11662,N_11395,N_11422);
nor U11663 (N_11663,N_11409,N_11282);
xor U11664 (N_11664,N_11342,N_11444);
xnor U11665 (N_11665,N_11268,N_11294);
and U11666 (N_11666,N_11380,N_11378);
or U11667 (N_11667,N_11278,N_11271);
nand U11668 (N_11668,N_11349,N_11409);
nand U11669 (N_11669,N_11358,N_11301);
nand U11670 (N_11670,N_11291,N_11419);
nand U11671 (N_11671,N_11399,N_11311);
or U11672 (N_11672,N_11477,N_11432);
nor U11673 (N_11673,N_11293,N_11424);
nand U11674 (N_11674,N_11288,N_11423);
xor U11675 (N_11675,N_11439,N_11413);
or U11676 (N_11676,N_11333,N_11317);
nor U11677 (N_11677,N_11354,N_11349);
nand U11678 (N_11678,N_11456,N_11414);
nor U11679 (N_11679,N_11374,N_11258);
and U11680 (N_11680,N_11389,N_11435);
nand U11681 (N_11681,N_11458,N_11486);
nor U11682 (N_11682,N_11260,N_11308);
and U11683 (N_11683,N_11404,N_11319);
nand U11684 (N_11684,N_11420,N_11297);
xnor U11685 (N_11685,N_11396,N_11309);
nand U11686 (N_11686,N_11331,N_11445);
and U11687 (N_11687,N_11367,N_11476);
and U11688 (N_11688,N_11492,N_11279);
nand U11689 (N_11689,N_11254,N_11328);
or U11690 (N_11690,N_11301,N_11342);
and U11691 (N_11691,N_11442,N_11481);
or U11692 (N_11692,N_11346,N_11378);
nand U11693 (N_11693,N_11254,N_11299);
xor U11694 (N_11694,N_11334,N_11415);
xnor U11695 (N_11695,N_11466,N_11451);
and U11696 (N_11696,N_11449,N_11267);
nor U11697 (N_11697,N_11396,N_11318);
and U11698 (N_11698,N_11281,N_11332);
or U11699 (N_11699,N_11428,N_11442);
nor U11700 (N_11700,N_11322,N_11462);
nor U11701 (N_11701,N_11488,N_11419);
nor U11702 (N_11702,N_11321,N_11394);
or U11703 (N_11703,N_11428,N_11342);
nand U11704 (N_11704,N_11351,N_11393);
or U11705 (N_11705,N_11343,N_11432);
and U11706 (N_11706,N_11308,N_11495);
nor U11707 (N_11707,N_11461,N_11368);
xor U11708 (N_11708,N_11401,N_11456);
nand U11709 (N_11709,N_11298,N_11467);
xnor U11710 (N_11710,N_11294,N_11326);
nand U11711 (N_11711,N_11385,N_11435);
xor U11712 (N_11712,N_11268,N_11482);
nor U11713 (N_11713,N_11332,N_11349);
nand U11714 (N_11714,N_11406,N_11282);
nor U11715 (N_11715,N_11391,N_11264);
nand U11716 (N_11716,N_11400,N_11320);
nand U11717 (N_11717,N_11401,N_11382);
nand U11718 (N_11718,N_11466,N_11291);
xnor U11719 (N_11719,N_11495,N_11335);
nor U11720 (N_11720,N_11341,N_11293);
xor U11721 (N_11721,N_11446,N_11378);
and U11722 (N_11722,N_11460,N_11367);
or U11723 (N_11723,N_11378,N_11425);
nor U11724 (N_11724,N_11469,N_11496);
or U11725 (N_11725,N_11447,N_11357);
or U11726 (N_11726,N_11355,N_11319);
and U11727 (N_11727,N_11427,N_11423);
xor U11728 (N_11728,N_11467,N_11441);
and U11729 (N_11729,N_11366,N_11397);
and U11730 (N_11730,N_11402,N_11371);
and U11731 (N_11731,N_11398,N_11331);
xor U11732 (N_11732,N_11466,N_11276);
nor U11733 (N_11733,N_11333,N_11463);
and U11734 (N_11734,N_11452,N_11321);
nor U11735 (N_11735,N_11475,N_11442);
or U11736 (N_11736,N_11284,N_11393);
or U11737 (N_11737,N_11285,N_11405);
or U11738 (N_11738,N_11400,N_11439);
xor U11739 (N_11739,N_11251,N_11471);
nand U11740 (N_11740,N_11390,N_11298);
and U11741 (N_11741,N_11298,N_11391);
xnor U11742 (N_11742,N_11382,N_11444);
or U11743 (N_11743,N_11325,N_11317);
nor U11744 (N_11744,N_11347,N_11452);
nand U11745 (N_11745,N_11481,N_11431);
nand U11746 (N_11746,N_11420,N_11328);
or U11747 (N_11747,N_11269,N_11274);
and U11748 (N_11748,N_11378,N_11394);
nand U11749 (N_11749,N_11354,N_11447);
nand U11750 (N_11750,N_11727,N_11520);
or U11751 (N_11751,N_11742,N_11525);
xor U11752 (N_11752,N_11553,N_11555);
or U11753 (N_11753,N_11711,N_11699);
nor U11754 (N_11754,N_11724,N_11579);
or U11755 (N_11755,N_11710,N_11708);
nand U11756 (N_11756,N_11530,N_11681);
nor U11757 (N_11757,N_11739,N_11734);
or U11758 (N_11758,N_11744,N_11573);
nand U11759 (N_11759,N_11630,N_11671);
nand U11760 (N_11760,N_11677,N_11745);
and U11761 (N_11761,N_11738,N_11693);
nand U11762 (N_11762,N_11552,N_11506);
or U11763 (N_11763,N_11574,N_11676);
xor U11764 (N_11764,N_11584,N_11690);
or U11765 (N_11765,N_11695,N_11501);
nand U11766 (N_11766,N_11649,N_11651);
xnor U11767 (N_11767,N_11604,N_11611);
xor U11768 (N_11768,N_11596,N_11568);
nand U11769 (N_11769,N_11578,N_11588);
xor U11770 (N_11770,N_11646,N_11500);
xnor U11771 (N_11771,N_11502,N_11533);
or U11772 (N_11772,N_11544,N_11624);
xor U11773 (N_11773,N_11562,N_11508);
xnor U11774 (N_11774,N_11600,N_11577);
xnor U11775 (N_11775,N_11661,N_11628);
nand U11776 (N_11776,N_11591,N_11593);
and U11777 (N_11777,N_11540,N_11507);
and U11778 (N_11778,N_11688,N_11747);
nand U11779 (N_11779,N_11720,N_11564);
and U11780 (N_11780,N_11670,N_11674);
nor U11781 (N_11781,N_11740,N_11602);
nand U11782 (N_11782,N_11598,N_11554);
nand U11783 (N_11783,N_11531,N_11510);
and U11784 (N_11784,N_11535,N_11513);
nand U11785 (N_11785,N_11615,N_11581);
xor U11786 (N_11786,N_11541,N_11650);
and U11787 (N_11787,N_11534,N_11580);
nor U11788 (N_11788,N_11639,N_11559);
and U11789 (N_11789,N_11539,N_11590);
nor U11790 (N_11790,N_11701,N_11567);
nor U11791 (N_11791,N_11503,N_11528);
nor U11792 (N_11792,N_11527,N_11666);
or U11793 (N_11793,N_11638,N_11730);
nand U11794 (N_11794,N_11705,N_11696);
xnor U11795 (N_11795,N_11697,N_11587);
nor U11796 (N_11796,N_11583,N_11620);
nor U11797 (N_11797,N_11655,N_11673);
or U11798 (N_11798,N_11709,N_11556);
xor U11799 (N_11799,N_11619,N_11537);
nor U11800 (N_11800,N_11504,N_11714);
and U11801 (N_11801,N_11576,N_11563);
nor U11802 (N_11802,N_11746,N_11692);
or U11803 (N_11803,N_11687,N_11737);
nand U11804 (N_11804,N_11678,N_11698);
and U11805 (N_11805,N_11606,N_11683);
nor U11806 (N_11806,N_11686,N_11728);
and U11807 (N_11807,N_11560,N_11523);
and U11808 (N_11808,N_11515,N_11684);
nand U11809 (N_11809,N_11643,N_11668);
xor U11810 (N_11810,N_11702,N_11667);
nor U11811 (N_11811,N_11631,N_11550);
and U11812 (N_11812,N_11542,N_11716);
and U11813 (N_11813,N_11521,N_11718);
nand U11814 (N_11814,N_11648,N_11543);
nand U11815 (N_11815,N_11538,N_11536);
or U11816 (N_11816,N_11572,N_11547);
xor U11817 (N_11817,N_11522,N_11597);
and U11818 (N_11818,N_11616,N_11675);
and U11819 (N_11819,N_11659,N_11548);
or U11820 (N_11820,N_11610,N_11685);
or U11821 (N_11821,N_11719,N_11715);
nand U11822 (N_11822,N_11735,N_11571);
and U11823 (N_11823,N_11617,N_11652);
nand U11824 (N_11824,N_11514,N_11749);
and U11825 (N_11825,N_11732,N_11601);
nand U11826 (N_11826,N_11656,N_11608);
xor U11827 (N_11827,N_11594,N_11725);
or U11828 (N_11828,N_11546,N_11558);
xor U11829 (N_11829,N_11634,N_11625);
or U11830 (N_11830,N_11703,N_11672);
and U11831 (N_11831,N_11733,N_11691);
xnor U11832 (N_11832,N_11633,N_11612);
and U11833 (N_11833,N_11595,N_11518);
nor U11834 (N_11834,N_11748,N_11641);
nor U11835 (N_11835,N_11529,N_11736);
nor U11836 (N_11836,N_11585,N_11603);
xor U11837 (N_11837,N_11645,N_11623);
and U11838 (N_11838,N_11614,N_11707);
nand U11839 (N_11839,N_11723,N_11582);
nand U11840 (N_11840,N_11660,N_11647);
nand U11841 (N_11841,N_11679,N_11729);
nor U11842 (N_11842,N_11519,N_11657);
or U11843 (N_11843,N_11524,N_11741);
or U11844 (N_11844,N_11629,N_11712);
nand U11845 (N_11845,N_11663,N_11653);
nor U11846 (N_11846,N_11517,N_11526);
xnor U11847 (N_11847,N_11613,N_11694);
nand U11848 (N_11848,N_11669,N_11644);
and U11849 (N_11849,N_11654,N_11516);
and U11850 (N_11850,N_11511,N_11607);
or U11851 (N_11851,N_11509,N_11658);
or U11852 (N_11852,N_11689,N_11704);
or U11853 (N_11853,N_11680,N_11575);
nor U11854 (N_11854,N_11599,N_11570);
nand U11855 (N_11855,N_11713,N_11549);
and U11856 (N_11856,N_11635,N_11665);
xor U11857 (N_11857,N_11589,N_11726);
xor U11858 (N_11858,N_11561,N_11565);
xnor U11859 (N_11859,N_11743,N_11700);
nor U11860 (N_11860,N_11731,N_11632);
or U11861 (N_11861,N_11627,N_11662);
and U11862 (N_11862,N_11586,N_11566);
or U11863 (N_11863,N_11717,N_11609);
and U11864 (N_11864,N_11706,N_11505);
and U11865 (N_11865,N_11569,N_11557);
xnor U11866 (N_11866,N_11722,N_11605);
and U11867 (N_11867,N_11636,N_11618);
and U11868 (N_11868,N_11664,N_11626);
nand U11869 (N_11869,N_11637,N_11512);
nand U11870 (N_11870,N_11721,N_11682);
nand U11871 (N_11871,N_11592,N_11532);
nand U11872 (N_11872,N_11621,N_11551);
and U11873 (N_11873,N_11642,N_11640);
nand U11874 (N_11874,N_11545,N_11622);
xor U11875 (N_11875,N_11583,N_11527);
nor U11876 (N_11876,N_11671,N_11694);
or U11877 (N_11877,N_11726,N_11524);
or U11878 (N_11878,N_11526,N_11660);
nand U11879 (N_11879,N_11609,N_11657);
and U11880 (N_11880,N_11541,N_11641);
nor U11881 (N_11881,N_11729,N_11736);
and U11882 (N_11882,N_11586,N_11558);
and U11883 (N_11883,N_11642,N_11689);
and U11884 (N_11884,N_11596,N_11514);
and U11885 (N_11885,N_11613,N_11544);
xor U11886 (N_11886,N_11526,N_11610);
xnor U11887 (N_11887,N_11676,N_11533);
xnor U11888 (N_11888,N_11739,N_11619);
nand U11889 (N_11889,N_11577,N_11650);
and U11890 (N_11890,N_11564,N_11567);
or U11891 (N_11891,N_11732,N_11597);
and U11892 (N_11892,N_11564,N_11504);
or U11893 (N_11893,N_11711,N_11740);
nor U11894 (N_11894,N_11680,N_11507);
and U11895 (N_11895,N_11572,N_11649);
or U11896 (N_11896,N_11542,N_11588);
nor U11897 (N_11897,N_11588,N_11689);
nor U11898 (N_11898,N_11685,N_11645);
nor U11899 (N_11899,N_11681,N_11649);
xnor U11900 (N_11900,N_11598,N_11548);
xor U11901 (N_11901,N_11508,N_11549);
nand U11902 (N_11902,N_11712,N_11709);
nand U11903 (N_11903,N_11657,N_11524);
nand U11904 (N_11904,N_11645,N_11692);
xnor U11905 (N_11905,N_11686,N_11552);
or U11906 (N_11906,N_11640,N_11600);
and U11907 (N_11907,N_11501,N_11538);
nor U11908 (N_11908,N_11593,N_11588);
xor U11909 (N_11909,N_11505,N_11509);
and U11910 (N_11910,N_11657,N_11625);
and U11911 (N_11911,N_11506,N_11530);
or U11912 (N_11912,N_11520,N_11583);
and U11913 (N_11913,N_11553,N_11576);
nor U11914 (N_11914,N_11593,N_11527);
nand U11915 (N_11915,N_11577,N_11642);
or U11916 (N_11916,N_11550,N_11515);
or U11917 (N_11917,N_11596,N_11658);
xnor U11918 (N_11918,N_11592,N_11606);
and U11919 (N_11919,N_11722,N_11661);
nor U11920 (N_11920,N_11691,N_11737);
or U11921 (N_11921,N_11733,N_11625);
and U11922 (N_11922,N_11667,N_11645);
nor U11923 (N_11923,N_11611,N_11630);
xor U11924 (N_11924,N_11514,N_11692);
and U11925 (N_11925,N_11555,N_11563);
nor U11926 (N_11926,N_11500,N_11644);
and U11927 (N_11927,N_11505,N_11563);
and U11928 (N_11928,N_11562,N_11517);
nand U11929 (N_11929,N_11584,N_11663);
xor U11930 (N_11930,N_11701,N_11606);
and U11931 (N_11931,N_11649,N_11538);
xnor U11932 (N_11932,N_11721,N_11528);
or U11933 (N_11933,N_11623,N_11552);
nand U11934 (N_11934,N_11685,N_11580);
xnor U11935 (N_11935,N_11572,N_11749);
nor U11936 (N_11936,N_11695,N_11500);
nand U11937 (N_11937,N_11526,N_11662);
nand U11938 (N_11938,N_11509,N_11689);
nor U11939 (N_11939,N_11673,N_11646);
nand U11940 (N_11940,N_11612,N_11680);
or U11941 (N_11941,N_11500,N_11582);
nand U11942 (N_11942,N_11539,N_11566);
or U11943 (N_11943,N_11637,N_11658);
and U11944 (N_11944,N_11575,N_11571);
nand U11945 (N_11945,N_11735,N_11620);
nor U11946 (N_11946,N_11502,N_11675);
and U11947 (N_11947,N_11555,N_11717);
xnor U11948 (N_11948,N_11661,N_11721);
nand U11949 (N_11949,N_11511,N_11519);
xnor U11950 (N_11950,N_11659,N_11628);
nor U11951 (N_11951,N_11681,N_11714);
and U11952 (N_11952,N_11732,N_11691);
xor U11953 (N_11953,N_11504,N_11557);
or U11954 (N_11954,N_11604,N_11592);
nand U11955 (N_11955,N_11697,N_11667);
and U11956 (N_11956,N_11570,N_11688);
xnor U11957 (N_11957,N_11717,N_11510);
nor U11958 (N_11958,N_11674,N_11600);
nand U11959 (N_11959,N_11504,N_11665);
or U11960 (N_11960,N_11546,N_11589);
xor U11961 (N_11961,N_11682,N_11555);
nor U11962 (N_11962,N_11637,N_11680);
nor U11963 (N_11963,N_11597,N_11669);
nand U11964 (N_11964,N_11523,N_11596);
and U11965 (N_11965,N_11549,N_11697);
or U11966 (N_11966,N_11634,N_11711);
or U11967 (N_11967,N_11715,N_11584);
nand U11968 (N_11968,N_11684,N_11577);
nor U11969 (N_11969,N_11661,N_11581);
nand U11970 (N_11970,N_11544,N_11524);
xor U11971 (N_11971,N_11594,N_11622);
nand U11972 (N_11972,N_11652,N_11534);
nor U11973 (N_11973,N_11617,N_11649);
xnor U11974 (N_11974,N_11515,N_11661);
xnor U11975 (N_11975,N_11671,N_11544);
and U11976 (N_11976,N_11726,N_11709);
or U11977 (N_11977,N_11669,N_11626);
xnor U11978 (N_11978,N_11738,N_11648);
nand U11979 (N_11979,N_11628,N_11684);
or U11980 (N_11980,N_11681,N_11601);
nor U11981 (N_11981,N_11593,N_11715);
and U11982 (N_11982,N_11648,N_11616);
nand U11983 (N_11983,N_11582,N_11586);
and U11984 (N_11984,N_11708,N_11734);
or U11985 (N_11985,N_11553,N_11606);
nor U11986 (N_11986,N_11622,N_11511);
or U11987 (N_11987,N_11545,N_11561);
and U11988 (N_11988,N_11693,N_11547);
nor U11989 (N_11989,N_11723,N_11702);
nor U11990 (N_11990,N_11731,N_11667);
or U11991 (N_11991,N_11692,N_11590);
or U11992 (N_11992,N_11686,N_11578);
xnor U11993 (N_11993,N_11532,N_11632);
and U11994 (N_11994,N_11532,N_11579);
and U11995 (N_11995,N_11520,N_11500);
xor U11996 (N_11996,N_11711,N_11679);
or U11997 (N_11997,N_11640,N_11533);
and U11998 (N_11998,N_11527,N_11704);
and U11999 (N_11999,N_11615,N_11616);
or U12000 (N_12000,N_11858,N_11876);
nand U12001 (N_12001,N_11822,N_11903);
nand U12002 (N_12002,N_11775,N_11849);
nor U12003 (N_12003,N_11875,N_11754);
nand U12004 (N_12004,N_11919,N_11826);
nor U12005 (N_12005,N_11940,N_11956);
or U12006 (N_12006,N_11998,N_11865);
nand U12007 (N_12007,N_11818,N_11761);
xor U12008 (N_12008,N_11817,N_11927);
or U12009 (N_12009,N_11837,N_11857);
or U12010 (N_12010,N_11778,N_11973);
and U12011 (N_12011,N_11871,N_11898);
nor U12012 (N_12012,N_11774,N_11877);
nand U12013 (N_12013,N_11772,N_11929);
nand U12014 (N_12014,N_11796,N_11989);
and U12015 (N_12015,N_11814,N_11937);
xor U12016 (N_12016,N_11983,N_11799);
and U12017 (N_12017,N_11951,N_11803);
nor U12018 (N_12018,N_11753,N_11808);
or U12019 (N_12019,N_11853,N_11889);
and U12020 (N_12020,N_11847,N_11873);
nand U12021 (N_12021,N_11966,N_11790);
xnor U12022 (N_12022,N_11985,N_11952);
xnor U12023 (N_12023,N_11982,N_11751);
xor U12024 (N_12024,N_11924,N_11773);
nand U12025 (N_12025,N_11820,N_11767);
xor U12026 (N_12026,N_11994,N_11816);
nand U12027 (N_12027,N_11827,N_11859);
and U12028 (N_12028,N_11913,N_11922);
nor U12029 (N_12029,N_11895,N_11801);
xor U12030 (N_12030,N_11992,N_11776);
and U12031 (N_12031,N_11917,N_11978);
nor U12032 (N_12032,N_11883,N_11750);
nor U12033 (N_12033,N_11806,N_11944);
nand U12034 (N_12034,N_11977,N_11974);
nor U12035 (N_12035,N_11906,N_11768);
nor U12036 (N_12036,N_11887,N_11984);
nand U12037 (N_12037,N_11804,N_11824);
or U12038 (N_12038,N_11894,N_11762);
and U12039 (N_12039,N_11935,N_11800);
or U12040 (N_12040,N_11884,N_11784);
or U12041 (N_12041,N_11972,N_11891);
and U12042 (N_12042,N_11901,N_11752);
and U12043 (N_12043,N_11797,N_11872);
nand U12044 (N_12044,N_11914,N_11925);
and U12045 (N_12045,N_11999,N_11771);
nand U12046 (N_12046,N_11829,N_11840);
nand U12047 (N_12047,N_11815,N_11830);
nand U12048 (N_12048,N_11967,N_11868);
nand U12049 (N_12049,N_11932,N_11856);
xnor U12050 (N_12050,N_11785,N_11809);
nand U12051 (N_12051,N_11961,N_11957);
nand U12052 (N_12052,N_11900,N_11834);
and U12053 (N_12053,N_11764,N_11802);
and U12054 (N_12054,N_11793,N_11791);
xor U12055 (N_12055,N_11947,N_11990);
and U12056 (N_12056,N_11941,N_11911);
and U12057 (N_12057,N_11788,N_11811);
xor U12058 (N_12058,N_11759,N_11787);
or U12059 (N_12059,N_11763,N_11867);
nand U12060 (N_12060,N_11958,N_11813);
xor U12061 (N_12061,N_11890,N_11869);
xor U12062 (N_12062,N_11833,N_11783);
xor U12063 (N_12063,N_11893,N_11907);
nor U12064 (N_12064,N_11879,N_11757);
nor U12065 (N_12065,N_11933,N_11888);
nor U12066 (N_12066,N_11968,N_11965);
nand U12067 (N_12067,N_11886,N_11920);
or U12068 (N_12068,N_11905,N_11786);
nand U12069 (N_12069,N_11792,N_11821);
or U12070 (N_12070,N_11777,N_11860);
xor U12071 (N_12071,N_11845,N_11831);
nand U12072 (N_12072,N_11874,N_11915);
nor U12073 (N_12073,N_11781,N_11904);
nor U12074 (N_12074,N_11918,N_11938);
nor U12075 (N_12075,N_11881,N_11844);
nand U12076 (N_12076,N_11769,N_11760);
nand U12077 (N_12077,N_11843,N_11916);
and U12078 (N_12078,N_11862,N_11842);
or U12079 (N_12079,N_11921,N_11943);
and U12080 (N_12080,N_11969,N_11758);
and U12081 (N_12081,N_11835,N_11836);
nand U12082 (N_12082,N_11839,N_11949);
and U12083 (N_12083,N_11948,N_11964);
or U12084 (N_12084,N_11995,N_11970);
nand U12085 (N_12085,N_11950,N_11945);
nor U12086 (N_12086,N_11988,N_11930);
or U12087 (N_12087,N_11812,N_11756);
xor U12088 (N_12088,N_11765,N_11980);
nand U12089 (N_12089,N_11854,N_11981);
or U12090 (N_12090,N_11880,N_11996);
and U12091 (N_12091,N_11882,N_11960);
xor U12092 (N_12092,N_11825,N_11838);
nand U12093 (N_12093,N_11782,N_11794);
xnor U12094 (N_12094,N_11976,N_11953);
and U12095 (N_12095,N_11975,N_11902);
nand U12096 (N_12096,N_11909,N_11766);
and U12097 (N_12097,N_11878,N_11851);
nand U12098 (N_12098,N_11850,N_11897);
nand U12099 (N_12099,N_11962,N_11912);
xnor U12100 (N_12100,N_11910,N_11848);
xor U12101 (N_12101,N_11819,N_11971);
nand U12102 (N_12102,N_11946,N_11846);
or U12103 (N_12103,N_11991,N_11789);
and U12104 (N_12104,N_11908,N_11928);
nand U12105 (N_12105,N_11855,N_11864);
nand U12106 (N_12106,N_11805,N_11863);
or U12107 (N_12107,N_11823,N_11993);
and U12108 (N_12108,N_11866,N_11899);
and U12109 (N_12109,N_11955,N_11828);
xor U12110 (N_12110,N_11896,N_11936);
xor U12111 (N_12111,N_11923,N_11987);
nor U12112 (N_12112,N_11795,N_11979);
nor U12113 (N_12113,N_11959,N_11939);
nor U12114 (N_12114,N_11832,N_11892);
or U12115 (N_12115,N_11755,N_11963);
nor U12116 (N_12116,N_11934,N_11841);
nand U12117 (N_12117,N_11807,N_11885);
nand U12118 (N_12118,N_11986,N_11779);
nor U12119 (N_12119,N_11954,N_11852);
nand U12120 (N_12120,N_11770,N_11780);
nand U12121 (N_12121,N_11870,N_11926);
or U12122 (N_12122,N_11861,N_11798);
xor U12123 (N_12123,N_11810,N_11997);
and U12124 (N_12124,N_11942,N_11931);
and U12125 (N_12125,N_11929,N_11796);
xnor U12126 (N_12126,N_11954,N_11992);
and U12127 (N_12127,N_11813,N_11837);
and U12128 (N_12128,N_11930,N_11882);
and U12129 (N_12129,N_11952,N_11939);
nor U12130 (N_12130,N_11944,N_11798);
nor U12131 (N_12131,N_11959,N_11771);
nor U12132 (N_12132,N_11895,N_11893);
and U12133 (N_12133,N_11847,N_11894);
xnor U12134 (N_12134,N_11833,N_11787);
nand U12135 (N_12135,N_11901,N_11821);
nand U12136 (N_12136,N_11840,N_11988);
nor U12137 (N_12137,N_11834,N_11928);
nor U12138 (N_12138,N_11771,N_11994);
and U12139 (N_12139,N_11958,N_11894);
or U12140 (N_12140,N_11800,N_11790);
nor U12141 (N_12141,N_11881,N_11750);
or U12142 (N_12142,N_11817,N_11798);
or U12143 (N_12143,N_11785,N_11988);
nand U12144 (N_12144,N_11933,N_11932);
or U12145 (N_12145,N_11930,N_11973);
and U12146 (N_12146,N_11827,N_11999);
and U12147 (N_12147,N_11850,N_11835);
nand U12148 (N_12148,N_11983,N_11961);
and U12149 (N_12149,N_11758,N_11781);
xor U12150 (N_12150,N_11853,N_11948);
and U12151 (N_12151,N_11820,N_11880);
or U12152 (N_12152,N_11946,N_11848);
xor U12153 (N_12153,N_11995,N_11910);
nand U12154 (N_12154,N_11831,N_11789);
nor U12155 (N_12155,N_11754,N_11847);
nor U12156 (N_12156,N_11878,N_11852);
nor U12157 (N_12157,N_11986,N_11871);
xnor U12158 (N_12158,N_11975,N_11861);
and U12159 (N_12159,N_11915,N_11943);
nand U12160 (N_12160,N_11883,N_11799);
nand U12161 (N_12161,N_11840,N_11899);
or U12162 (N_12162,N_11891,N_11859);
or U12163 (N_12163,N_11754,N_11781);
xnor U12164 (N_12164,N_11830,N_11939);
and U12165 (N_12165,N_11758,N_11914);
or U12166 (N_12166,N_11955,N_11997);
xnor U12167 (N_12167,N_11903,N_11791);
nand U12168 (N_12168,N_11934,N_11809);
xor U12169 (N_12169,N_11944,N_11787);
and U12170 (N_12170,N_11823,N_11917);
and U12171 (N_12171,N_11769,N_11905);
or U12172 (N_12172,N_11863,N_11919);
nand U12173 (N_12173,N_11768,N_11814);
nand U12174 (N_12174,N_11909,N_11835);
nand U12175 (N_12175,N_11877,N_11865);
nand U12176 (N_12176,N_11962,N_11887);
nor U12177 (N_12177,N_11827,N_11969);
nand U12178 (N_12178,N_11851,N_11809);
nand U12179 (N_12179,N_11754,N_11955);
and U12180 (N_12180,N_11773,N_11987);
or U12181 (N_12181,N_11979,N_11997);
or U12182 (N_12182,N_11808,N_11758);
xnor U12183 (N_12183,N_11906,N_11840);
or U12184 (N_12184,N_11767,N_11913);
nor U12185 (N_12185,N_11787,N_11753);
nor U12186 (N_12186,N_11946,N_11853);
or U12187 (N_12187,N_11863,N_11813);
nor U12188 (N_12188,N_11929,N_11945);
nand U12189 (N_12189,N_11923,N_11953);
nand U12190 (N_12190,N_11762,N_11998);
nor U12191 (N_12191,N_11852,N_11771);
and U12192 (N_12192,N_11859,N_11912);
nand U12193 (N_12193,N_11952,N_11963);
nor U12194 (N_12194,N_11951,N_11777);
nand U12195 (N_12195,N_11775,N_11787);
or U12196 (N_12196,N_11975,N_11862);
nor U12197 (N_12197,N_11880,N_11867);
xor U12198 (N_12198,N_11919,N_11801);
or U12199 (N_12199,N_11943,N_11820);
or U12200 (N_12200,N_11770,N_11927);
nand U12201 (N_12201,N_11810,N_11845);
nor U12202 (N_12202,N_11766,N_11895);
and U12203 (N_12203,N_11930,N_11790);
xor U12204 (N_12204,N_11900,N_11868);
nor U12205 (N_12205,N_11964,N_11812);
xor U12206 (N_12206,N_11901,N_11956);
and U12207 (N_12207,N_11911,N_11763);
xnor U12208 (N_12208,N_11874,N_11969);
and U12209 (N_12209,N_11929,N_11854);
nor U12210 (N_12210,N_11829,N_11806);
or U12211 (N_12211,N_11987,N_11977);
xnor U12212 (N_12212,N_11904,N_11811);
nand U12213 (N_12213,N_11883,N_11843);
or U12214 (N_12214,N_11874,N_11862);
xnor U12215 (N_12215,N_11976,N_11810);
xor U12216 (N_12216,N_11891,N_11801);
xor U12217 (N_12217,N_11753,N_11866);
nor U12218 (N_12218,N_11959,N_11999);
or U12219 (N_12219,N_11993,N_11845);
nand U12220 (N_12220,N_11978,N_11889);
or U12221 (N_12221,N_11777,N_11764);
or U12222 (N_12222,N_11832,N_11932);
nand U12223 (N_12223,N_11882,N_11908);
and U12224 (N_12224,N_11984,N_11752);
and U12225 (N_12225,N_11851,N_11988);
nand U12226 (N_12226,N_11818,N_11927);
xor U12227 (N_12227,N_11984,N_11941);
and U12228 (N_12228,N_11873,N_11792);
nor U12229 (N_12229,N_11901,N_11822);
xor U12230 (N_12230,N_11854,N_11802);
nor U12231 (N_12231,N_11966,N_11843);
nand U12232 (N_12232,N_11900,N_11931);
or U12233 (N_12233,N_11889,N_11914);
xor U12234 (N_12234,N_11853,N_11868);
xnor U12235 (N_12235,N_11978,N_11810);
and U12236 (N_12236,N_11812,N_11981);
xnor U12237 (N_12237,N_11940,N_11907);
and U12238 (N_12238,N_11847,N_11959);
and U12239 (N_12239,N_11823,N_11774);
nand U12240 (N_12240,N_11758,N_11807);
nor U12241 (N_12241,N_11841,N_11973);
xor U12242 (N_12242,N_11896,N_11962);
or U12243 (N_12243,N_11887,N_11843);
nor U12244 (N_12244,N_11752,N_11809);
or U12245 (N_12245,N_11758,N_11901);
and U12246 (N_12246,N_11987,N_11798);
or U12247 (N_12247,N_11774,N_11829);
or U12248 (N_12248,N_11951,N_11769);
nand U12249 (N_12249,N_11840,N_11946);
xnor U12250 (N_12250,N_12136,N_12060);
or U12251 (N_12251,N_12134,N_12096);
nand U12252 (N_12252,N_12037,N_12123);
or U12253 (N_12253,N_12210,N_12156);
or U12254 (N_12254,N_12099,N_12174);
nand U12255 (N_12255,N_12049,N_12157);
nor U12256 (N_12256,N_12073,N_12158);
and U12257 (N_12257,N_12044,N_12125);
or U12258 (N_12258,N_12149,N_12105);
xnor U12259 (N_12259,N_12195,N_12238);
nand U12260 (N_12260,N_12208,N_12040);
nor U12261 (N_12261,N_12102,N_12169);
nor U12262 (N_12262,N_12237,N_12046);
and U12263 (N_12263,N_12217,N_12212);
nor U12264 (N_12264,N_12047,N_12178);
and U12265 (N_12265,N_12038,N_12150);
xor U12266 (N_12266,N_12233,N_12110);
xor U12267 (N_12267,N_12072,N_12222);
nor U12268 (N_12268,N_12041,N_12152);
or U12269 (N_12269,N_12207,N_12243);
xnor U12270 (N_12270,N_12194,N_12161);
nor U12271 (N_12271,N_12114,N_12120);
and U12272 (N_12272,N_12187,N_12234);
or U12273 (N_12273,N_12124,N_12209);
xor U12274 (N_12274,N_12227,N_12028);
and U12275 (N_12275,N_12067,N_12220);
nor U12276 (N_12276,N_12200,N_12019);
or U12277 (N_12277,N_12062,N_12221);
nor U12278 (N_12278,N_12192,N_12190);
nor U12279 (N_12279,N_12085,N_12117);
or U12280 (N_12280,N_12081,N_12104);
xor U12281 (N_12281,N_12170,N_12188);
and U12282 (N_12282,N_12057,N_12100);
and U12283 (N_12283,N_12131,N_12162);
xnor U12284 (N_12284,N_12132,N_12051);
nor U12285 (N_12285,N_12166,N_12130);
nand U12286 (N_12286,N_12016,N_12020);
or U12287 (N_12287,N_12053,N_12108);
and U12288 (N_12288,N_12246,N_12167);
nand U12289 (N_12289,N_12086,N_12168);
or U12290 (N_12290,N_12155,N_12230);
nand U12291 (N_12291,N_12186,N_12177);
nand U12292 (N_12292,N_12055,N_12010);
and U12293 (N_12293,N_12247,N_12014);
nor U12294 (N_12294,N_12148,N_12127);
or U12295 (N_12295,N_12244,N_12018);
or U12296 (N_12296,N_12185,N_12201);
xnor U12297 (N_12297,N_12023,N_12043);
and U12298 (N_12298,N_12141,N_12024);
nor U12299 (N_12299,N_12008,N_12199);
or U12300 (N_12300,N_12021,N_12203);
nand U12301 (N_12301,N_12068,N_12214);
nand U12302 (N_12302,N_12173,N_12142);
or U12303 (N_12303,N_12121,N_12082);
or U12304 (N_12304,N_12113,N_12112);
nor U12305 (N_12305,N_12075,N_12074);
nor U12306 (N_12306,N_12025,N_12163);
and U12307 (N_12307,N_12058,N_12129);
and U12308 (N_12308,N_12229,N_12126);
or U12309 (N_12309,N_12071,N_12064);
xor U12310 (N_12310,N_12029,N_12245);
nand U12311 (N_12311,N_12140,N_12191);
nor U12312 (N_12312,N_12183,N_12223);
xor U12313 (N_12313,N_12009,N_12181);
nand U12314 (N_12314,N_12045,N_12239);
and U12315 (N_12315,N_12034,N_12248);
or U12316 (N_12316,N_12035,N_12015);
nor U12317 (N_12317,N_12002,N_12103);
or U12318 (N_12318,N_12241,N_12143);
xor U12319 (N_12319,N_12116,N_12080);
xor U12320 (N_12320,N_12118,N_12011);
nor U12321 (N_12321,N_12059,N_12013);
xnor U12322 (N_12322,N_12228,N_12176);
nand U12323 (N_12323,N_12033,N_12189);
xnor U12324 (N_12324,N_12109,N_12030);
nand U12325 (N_12325,N_12079,N_12159);
nand U12326 (N_12326,N_12165,N_12111);
nor U12327 (N_12327,N_12083,N_12098);
and U12328 (N_12328,N_12061,N_12171);
or U12329 (N_12329,N_12135,N_12095);
nor U12330 (N_12330,N_12048,N_12240);
xnor U12331 (N_12331,N_12145,N_12092);
xnor U12332 (N_12332,N_12146,N_12231);
xnor U12333 (N_12333,N_12115,N_12225);
and U12334 (N_12334,N_12242,N_12069);
nand U12335 (N_12335,N_12000,N_12179);
or U12336 (N_12336,N_12003,N_12001);
xor U12337 (N_12337,N_12006,N_12084);
and U12338 (N_12338,N_12097,N_12215);
and U12339 (N_12339,N_12042,N_12147);
nor U12340 (N_12340,N_12172,N_12107);
nor U12341 (N_12341,N_12219,N_12218);
nand U12342 (N_12342,N_12235,N_12022);
xor U12343 (N_12343,N_12036,N_12206);
nor U12344 (N_12344,N_12232,N_12122);
and U12345 (N_12345,N_12106,N_12224);
and U12346 (N_12346,N_12026,N_12182);
nor U12347 (N_12347,N_12128,N_12091);
xnor U12348 (N_12348,N_12004,N_12198);
and U12349 (N_12349,N_12090,N_12196);
xor U12350 (N_12350,N_12052,N_12101);
xnor U12351 (N_12351,N_12088,N_12050);
and U12352 (N_12352,N_12216,N_12063);
and U12353 (N_12353,N_12249,N_12087);
nor U12354 (N_12354,N_12031,N_12093);
or U12355 (N_12355,N_12054,N_12184);
nand U12356 (N_12356,N_12236,N_12077);
xor U12357 (N_12357,N_12160,N_12007);
or U12358 (N_12358,N_12211,N_12180);
nor U12359 (N_12359,N_12151,N_12164);
and U12360 (N_12360,N_12154,N_12193);
nand U12361 (N_12361,N_12137,N_12226);
or U12362 (N_12362,N_12138,N_12133);
or U12363 (N_12363,N_12204,N_12078);
nand U12364 (N_12364,N_12144,N_12027);
and U12365 (N_12365,N_12012,N_12032);
or U12366 (N_12366,N_12175,N_12153);
nand U12367 (N_12367,N_12094,N_12205);
nor U12368 (N_12368,N_12070,N_12213);
and U12369 (N_12369,N_12065,N_12089);
nor U12370 (N_12370,N_12056,N_12119);
xnor U12371 (N_12371,N_12202,N_12017);
nand U12372 (N_12372,N_12039,N_12005);
nor U12373 (N_12373,N_12197,N_12139);
nor U12374 (N_12374,N_12076,N_12066);
or U12375 (N_12375,N_12133,N_12033);
and U12376 (N_12376,N_12193,N_12139);
xnor U12377 (N_12377,N_12186,N_12150);
nor U12378 (N_12378,N_12027,N_12132);
nand U12379 (N_12379,N_12221,N_12068);
xor U12380 (N_12380,N_12195,N_12067);
nand U12381 (N_12381,N_12074,N_12022);
nor U12382 (N_12382,N_12035,N_12089);
nand U12383 (N_12383,N_12050,N_12179);
xor U12384 (N_12384,N_12238,N_12016);
or U12385 (N_12385,N_12050,N_12121);
nand U12386 (N_12386,N_12034,N_12055);
and U12387 (N_12387,N_12027,N_12169);
or U12388 (N_12388,N_12033,N_12240);
nor U12389 (N_12389,N_12075,N_12209);
nand U12390 (N_12390,N_12139,N_12182);
nor U12391 (N_12391,N_12057,N_12238);
xnor U12392 (N_12392,N_12010,N_12167);
and U12393 (N_12393,N_12111,N_12146);
nand U12394 (N_12394,N_12144,N_12003);
nand U12395 (N_12395,N_12089,N_12245);
nor U12396 (N_12396,N_12114,N_12028);
or U12397 (N_12397,N_12241,N_12149);
or U12398 (N_12398,N_12168,N_12110);
nor U12399 (N_12399,N_12082,N_12013);
nand U12400 (N_12400,N_12247,N_12244);
or U12401 (N_12401,N_12171,N_12120);
nor U12402 (N_12402,N_12028,N_12113);
nand U12403 (N_12403,N_12055,N_12174);
or U12404 (N_12404,N_12081,N_12135);
xnor U12405 (N_12405,N_12179,N_12184);
nor U12406 (N_12406,N_12195,N_12006);
or U12407 (N_12407,N_12098,N_12202);
xor U12408 (N_12408,N_12065,N_12187);
xnor U12409 (N_12409,N_12236,N_12075);
nand U12410 (N_12410,N_12218,N_12245);
nor U12411 (N_12411,N_12214,N_12212);
and U12412 (N_12412,N_12194,N_12153);
and U12413 (N_12413,N_12145,N_12034);
nor U12414 (N_12414,N_12057,N_12017);
or U12415 (N_12415,N_12224,N_12125);
nor U12416 (N_12416,N_12137,N_12062);
and U12417 (N_12417,N_12079,N_12121);
nand U12418 (N_12418,N_12230,N_12164);
nand U12419 (N_12419,N_12109,N_12174);
and U12420 (N_12420,N_12225,N_12085);
nand U12421 (N_12421,N_12063,N_12120);
or U12422 (N_12422,N_12131,N_12170);
or U12423 (N_12423,N_12094,N_12082);
or U12424 (N_12424,N_12007,N_12015);
nor U12425 (N_12425,N_12164,N_12041);
xor U12426 (N_12426,N_12085,N_12007);
or U12427 (N_12427,N_12211,N_12170);
or U12428 (N_12428,N_12249,N_12050);
and U12429 (N_12429,N_12238,N_12113);
nand U12430 (N_12430,N_12091,N_12216);
and U12431 (N_12431,N_12047,N_12061);
xor U12432 (N_12432,N_12236,N_12073);
nand U12433 (N_12433,N_12159,N_12104);
xnor U12434 (N_12434,N_12097,N_12143);
and U12435 (N_12435,N_12075,N_12168);
nand U12436 (N_12436,N_12028,N_12176);
nor U12437 (N_12437,N_12041,N_12091);
nand U12438 (N_12438,N_12084,N_12113);
nand U12439 (N_12439,N_12108,N_12119);
nand U12440 (N_12440,N_12002,N_12041);
xnor U12441 (N_12441,N_12035,N_12066);
or U12442 (N_12442,N_12103,N_12120);
nand U12443 (N_12443,N_12072,N_12186);
and U12444 (N_12444,N_12090,N_12103);
and U12445 (N_12445,N_12215,N_12020);
xor U12446 (N_12446,N_12228,N_12081);
or U12447 (N_12447,N_12080,N_12161);
and U12448 (N_12448,N_12120,N_12002);
nand U12449 (N_12449,N_12146,N_12216);
nor U12450 (N_12450,N_12107,N_12202);
nand U12451 (N_12451,N_12101,N_12117);
nor U12452 (N_12452,N_12226,N_12100);
nand U12453 (N_12453,N_12092,N_12201);
xor U12454 (N_12454,N_12064,N_12202);
nand U12455 (N_12455,N_12010,N_12066);
and U12456 (N_12456,N_12121,N_12160);
xnor U12457 (N_12457,N_12189,N_12178);
and U12458 (N_12458,N_12024,N_12105);
and U12459 (N_12459,N_12207,N_12038);
and U12460 (N_12460,N_12198,N_12249);
and U12461 (N_12461,N_12035,N_12131);
and U12462 (N_12462,N_12181,N_12133);
nor U12463 (N_12463,N_12025,N_12203);
xor U12464 (N_12464,N_12122,N_12171);
xor U12465 (N_12465,N_12031,N_12073);
xnor U12466 (N_12466,N_12059,N_12206);
xor U12467 (N_12467,N_12144,N_12132);
or U12468 (N_12468,N_12110,N_12225);
or U12469 (N_12469,N_12167,N_12099);
or U12470 (N_12470,N_12082,N_12127);
and U12471 (N_12471,N_12040,N_12046);
and U12472 (N_12472,N_12243,N_12116);
nand U12473 (N_12473,N_12174,N_12197);
nor U12474 (N_12474,N_12016,N_12215);
and U12475 (N_12475,N_12092,N_12041);
and U12476 (N_12476,N_12126,N_12239);
nand U12477 (N_12477,N_12117,N_12205);
or U12478 (N_12478,N_12230,N_12029);
nand U12479 (N_12479,N_12114,N_12156);
nand U12480 (N_12480,N_12243,N_12087);
or U12481 (N_12481,N_12085,N_12241);
nand U12482 (N_12482,N_12058,N_12092);
xnor U12483 (N_12483,N_12147,N_12115);
xnor U12484 (N_12484,N_12162,N_12177);
xor U12485 (N_12485,N_12092,N_12103);
xnor U12486 (N_12486,N_12121,N_12074);
or U12487 (N_12487,N_12007,N_12062);
xnor U12488 (N_12488,N_12110,N_12191);
and U12489 (N_12489,N_12203,N_12076);
nor U12490 (N_12490,N_12118,N_12108);
or U12491 (N_12491,N_12013,N_12026);
and U12492 (N_12492,N_12193,N_12179);
nor U12493 (N_12493,N_12213,N_12084);
or U12494 (N_12494,N_12098,N_12128);
xnor U12495 (N_12495,N_12204,N_12248);
xor U12496 (N_12496,N_12107,N_12103);
xor U12497 (N_12497,N_12172,N_12065);
xor U12498 (N_12498,N_12110,N_12045);
and U12499 (N_12499,N_12199,N_12226);
xor U12500 (N_12500,N_12416,N_12349);
xnor U12501 (N_12501,N_12442,N_12341);
and U12502 (N_12502,N_12309,N_12461);
and U12503 (N_12503,N_12449,N_12375);
xor U12504 (N_12504,N_12268,N_12258);
nand U12505 (N_12505,N_12293,N_12318);
nand U12506 (N_12506,N_12418,N_12270);
nand U12507 (N_12507,N_12274,N_12321);
nand U12508 (N_12508,N_12443,N_12494);
and U12509 (N_12509,N_12451,N_12407);
xnor U12510 (N_12510,N_12422,N_12426);
and U12511 (N_12511,N_12291,N_12356);
or U12512 (N_12512,N_12402,N_12350);
and U12513 (N_12513,N_12339,N_12295);
nand U12514 (N_12514,N_12464,N_12421);
or U12515 (N_12515,N_12287,N_12381);
or U12516 (N_12516,N_12317,N_12450);
nand U12517 (N_12517,N_12272,N_12476);
or U12518 (N_12518,N_12305,N_12300);
and U12519 (N_12519,N_12338,N_12495);
xor U12520 (N_12520,N_12403,N_12331);
nand U12521 (N_12521,N_12286,N_12490);
or U12522 (N_12522,N_12297,N_12279);
and U12523 (N_12523,N_12444,N_12362);
xor U12524 (N_12524,N_12492,N_12352);
or U12525 (N_12525,N_12313,N_12322);
nand U12526 (N_12526,N_12281,N_12430);
and U12527 (N_12527,N_12376,N_12377);
or U12528 (N_12528,N_12342,N_12265);
or U12529 (N_12529,N_12334,N_12499);
or U12530 (N_12530,N_12327,N_12435);
xor U12531 (N_12531,N_12343,N_12471);
nor U12532 (N_12532,N_12311,N_12480);
or U12533 (N_12533,N_12353,N_12389);
nand U12534 (N_12534,N_12283,N_12367);
and U12535 (N_12535,N_12436,N_12459);
and U12536 (N_12536,N_12384,N_12371);
and U12537 (N_12537,N_12429,N_12257);
nor U12538 (N_12538,N_12346,N_12386);
xnor U12539 (N_12539,N_12397,N_12278);
xor U12540 (N_12540,N_12340,N_12292);
and U12541 (N_12541,N_12487,N_12423);
or U12542 (N_12542,N_12332,N_12348);
or U12543 (N_12543,N_12280,N_12361);
and U12544 (N_12544,N_12351,N_12453);
or U12545 (N_12545,N_12387,N_12411);
and U12546 (N_12546,N_12428,N_12304);
xor U12547 (N_12547,N_12329,N_12456);
and U12548 (N_12548,N_12432,N_12269);
or U12549 (N_12549,N_12315,N_12282);
nor U12550 (N_12550,N_12468,N_12474);
nor U12551 (N_12551,N_12485,N_12398);
xor U12552 (N_12552,N_12488,N_12379);
and U12553 (N_12553,N_12445,N_12424);
nand U12554 (N_12554,N_12333,N_12306);
or U12555 (N_12555,N_12308,N_12363);
and U12556 (N_12556,N_12395,N_12344);
nand U12557 (N_12557,N_12314,N_12307);
nand U12558 (N_12558,N_12335,N_12462);
and U12559 (N_12559,N_12498,N_12441);
and U12560 (N_12560,N_12369,N_12417);
nand U12561 (N_12561,N_12290,N_12326);
and U12562 (N_12562,N_12271,N_12275);
and U12563 (N_12563,N_12368,N_12483);
nor U12564 (N_12564,N_12415,N_12382);
xor U12565 (N_12565,N_12408,N_12277);
and U12566 (N_12566,N_12320,N_12405);
and U12567 (N_12567,N_12469,N_12460);
and U12568 (N_12568,N_12285,N_12372);
xnor U12569 (N_12569,N_12253,N_12373);
and U12570 (N_12570,N_12284,N_12431);
xnor U12571 (N_12571,N_12425,N_12433);
or U12572 (N_12572,N_12336,N_12319);
nor U12573 (N_12573,N_12414,N_12404);
nand U12574 (N_12574,N_12380,N_12259);
or U12575 (N_12575,N_12496,N_12472);
or U12576 (N_12576,N_12448,N_12458);
xor U12577 (N_12577,N_12486,N_12410);
nand U12578 (N_12578,N_12470,N_12301);
and U12579 (N_12579,N_12374,N_12267);
and U12580 (N_12580,N_12359,N_12427);
nor U12581 (N_12581,N_12330,N_12446);
and U12582 (N_12582,N_12289,N_12252);
nand U12583 (N_12583,N_12262,N_12264);
or U12584 (N_12584,N_12288,N_12481);
and U12585 (N_12585,N_12260,N_12325);
and U12586 (N_12586,N_12463,N_12254);
or U12587 (N_12587,N_12392,N_12294);
or U12588 (N_12588,N_12316,N_12452);
xnor U12589 (N_12589,N_12312,N_12357);
or U12590 (N_12590,N_12365,N_12337);
nand U12591 (N_12591,N_12296,N_12457);
nor U12592 (N_12592,N_12302,N_12491);
nand U12593 (N_12593,N_12303,N_12482);
or U12594 (N_12594,N_12256,N_12420);
and U12595 (N_12595,N_12385,N_12355);
nor U12596 (N_12596,N_12255,N_12412);
nor U12597 (N_12597,N_12455,N_12378);
xnor U12598 (N_12598,N_12401,N_12383);
or U12599 (N_12599,N_12419,N_12347);
nor U12600 (N_12600,N_12261,N_12406);
nor U12601 (N_12601,N_12388,N_12489);
nand U12602 (N_12602,N_12447,N_12366);
xor U12603 (N_12603,N_12394,N_12413);
xor U12604 (N_12604,N_12323,N_12479);
or U12605 (N_12605,N_12467,N_12263);
and U12606 (N_12606,N_12299,N_12493);
and U12607 (N_12607,N_12251,N_12391);
and U12608 (N_12608,N_12437,N_12250);
xnor U12609 (N_12609,N_12298,N_12400);
xor U12610 (N_12610,N_12328,N_12310);
nand U12611 (N_12611,N_12390,N_12454);
nand U12612 (N_12612,N_12364,N_12473);
nand U12613 (N_12613,N_12358,N_12399);
nand U12614 (N_12614,N_12409,N_12438);
nand U12615 (N_12615,N_12477,N_12345);
nor U12616 (N_12616,N_12484,N_12440);
and U12617 (N_12617,N_12466,N_12273);
nor U12618 (N_12618,N_12370,N_12393);
nand U12619 (N_12619,N_12465,N_12276);
nor U12620 (N_12620,N_12475,N_12396);
nand U12621 (N_12621,N_12497,N_12360);
xor U12622 (N_12622,N_12324,N_12266);
or U12623 (N_12623,N_12434,N_12478);
xor U12624 (N_12624,N_12354,N_12439);
nor U12625 (N_12625,N_12422,N_12413);
and U12626 (N_12626,N_12434,N_12369);
or U12627 (N_12627,N_12278,N_12318);
xor U12628 (N_12628,N_12488,N_12311);
or U12629 (N_12629,N_12483,N_12497);
nand U12630 (N_12630,N_12373,N_12488);
nand U12631 (N_12631,N_12419,N_12294);
and U12632 (N_12632,N_12343,N_12399);
xor U12633 (N_12633,N_12352,N_12411);
and U12634 (N_12634,N_12429,N_12392);
nand U12635 (N_12635,N_12470,N_12345);
xnor U12636 (N_12636,N_12396,N_12263);
nor U12637 (N_12637,N_12379,N_12388);
nand U12638 (N_12638,N_12402,N_12265);
xor U12639 (N_12639,N_12435,N_12276);
nor U12640 (N_12640,N_12409,N_12348);
xor U12641 (N_12641,N_12262,N_12352);
and U12642 (N_12642,N_12487,N_12349);
nor U12643 (N_12643,N_12403,N_12328);
and U12644 (N_12644,N_12445,N_12281);
nor U12645 (N_12645,N_12456,N_12264);
or U12646 (N_12646,N_12285,N_12344);
and U12647 (N_12647,N_12377,N_12413);
nor U12648 (N_12648,N_12314,N_12353);
nand U12649 (N_12649,N_12311,N_12309);
nor U12650 (N_12650,N_12476,N_12329);
xor U12651 (N_12651,N_12419,N_12297);
nand U12652 (N_12652,N_12464,N_12285);
nand U12653 (N_12653,N_12411,N_12255);
nand U12654 (N_12654,N_12444,N_12286);
and U12655 (N_12655,N_12251,N_12430);
nand U12656 (N_12656,N_12336,N_12266);
nor U12657 (N_12657,N_12281,N_12493);
nand U12658 (N_12658,N_12420,N_12332);
nand U12659 (N_12659,N_12305,N_12326);
or U12660 (N_12660,N_12332,N_12303);
xnor U12661 (N_12661,N_12371,N_12463);
and U12662 (N_12662,N_12414,N_12460);
and U12663 (N_12663,N_12440,N_12446);
or U12664 (N_12664,N_12415,N_12253);
or U12665 (N_12665,N_12467,N_12397);
xor U12666 (N_12666,N_12322,N_12397);
xor U12667 (N_12667,N_12461,N_12437);
and U12668 (N_12668,N_12250,N_12472);
xor U12669 (N_12669,N_12291,N_12396);
nor U12670 (N_12670,N_12491,N_12328);
nand U12671 (N_12671,N_12473,N_12256);
xnor U12672 (N_12672,N_12356,N_12270);
and U12673 (N_12673,N_12446,N_12275);
nor U12674 (N_12674,N_12491,N_12416);
and U12675 (N_12675,N_12383,N_12444);
xnor U12676 (N_12676,N_12434,N_12424);
nor U12677 (N_12677,N_12276,N_12437);
or U12678 (N_12678,N_12358,N_12396);
or U12679 (N_12679,N_12412,N_12267);
and U12680 (N_12680,N_12480,N_12482);
xnor U12681 (N_12681,N_12273,N_12252);
or U12682 (N_12682,N_12362,N_12471);
or U12683 (N_12683,N_12386,N_12331);
and U12684 (N_12684,N_12493,N_12380);
nand U12685 (N_12685,N_12362,N_12306);
or U12686 (N_12686,N_12364,N_12279);
xnor U12687 (N_12687,N_12286,N_12393);
or U12688 (N_12688,N_12346,N_12456);
nand U12689 (N_12689,N_12354,N_12447);
and U12690 (N_12690,N_12376,N_12328);
and U12691 (N_12691,N_12482,N_12443);
nand U12692 (N_12692,N_12316,N_12414);
nor U12693 (N_12693,N_12290,N_12271);
or U12694 (N_12694,N_12286,N_12470);
xnor U12695 (N_12695,N_12428,N_12457);
nor U12696 (N_12696,N_12425,N_12298);
or U12697 (N_12697,N_12436,N_12272);
nor U12698 (N_12698,N_12488,N_12362);
or U12699 (N_12699,N_12346,N_12487);
and U12700 (N_12700,N_12493,N_12295);
and U12701 (N_12701,N_12443,N_12428);
and U12702 (N_12702,N_12390,N_12359);
nand U12703 (N_12703,N_12334,N_12421);
or U12704 (N_12704,N_12275,N_12278);
or U12705 (N_12705,N_12422,N_12459);
xnor U12706 (N_12706,N_12411,N_12473);
nor U12707 (N_12707,N_12337,N_12321);
nor U12708 (N_12708,N_12345,N_12316);
nor U12709 (N_12709,N_12468,N_12443);
or U12710 (N_12710,N_12450,N_12436);
xnor U12711 (N_12711,N_12452,N_12338);
xnor U12712 (N_12712,N_12421,N_12263);
or U12713 (N_12713,N_12260,N_12402);
nand U12714 (N_12714,N_12434,N_12493);
and U12715 (N_12715,N_12341,N_12397);
and U12716 (N_12716,N_12383,N_12375);
nand U12717 (N_12717,N_12455,N_12477);
or U12718 (N_12718,N_12356,N_12460);
nor U12719 (N_12719,N_12348,N_12279);
xnor U12720 (N_12720,N_12414,N_12478);
nor U12721 (N_12721,N_12366,N_12378);
or U12722 (N_12722,N_12380,N_12262);
xnor U12723 (N_12723,N_12307,N_12285);
xnor U12724 (N_12724,N_12480,N_12454);
nor U12725 (N_12725,N_12395,N_12495);
nor U12726 (N_12726,N_12443,N_12419);
nand U12727 (N_12727,N_12346,N_12337);
xor U12728 (N_12728,N_12418,N_12491);
and U12729 (N_12729,N_12273,N_12394);
or U12730 (N_12730,N_12250,N_12276);
nand U12731 (N_12731,N_12319,N_12425);
or U12732 (N_12732,N_12471,N_12429);
or U12733 (N_12733,N_12251,N_12444);
or U12734 (N_12734,N_12454,N_12364);
or U12735 (N_12735,N_12487,N_12439);
nand U12736 (N_12736,N_12320,N_12269);
and U12737 (N_12737,N_12456,N_12284);
nand U12738 (N_12738,N_12452,N_12270);
xnor U12739 (N_12739,N_12411,N_12256);
nand U12740 (N_12740,N_12369,N_12288);
nand U12741 (N_12741,N_12431,N_12342);
nand U12742 (N_12742,N_12268,N_12315);
nand U12743 (N_12743,N_12290,N_12474);
xnor U12744 (N_12744,N_12281,N_12434);
nand U12745 (N_12745,N_12280,N_12336);
nand U12746 (N_12746,N_12355,N_12319);
nor U12747 (N_12747,N_12371,N_12453);
nor U12748 (N_12748,N_12364,N_12375);
xnor U12749 (N_12749,N_12423,N_12333);
nor U12750 (N_12750,N_12717,N_12610);
nor U12751 (N_12751,N_12510,N_12558);
xor U12752 (N_12752,N_12687,N_12611);
and U12753 (N_12753,N_12516,N_12708);
or U12754 (N_12754,N_12730,N_12654);
and U12755 (N_12755,N_12570,N_12580);
or U12756 (N_12756,N_12672,N_12636);
or U12757 (N_12757,N_12598,N_12551);
nor U12758 (N_12758,N_12603,N_12606);
nor U12759 (N_12759,N_12573,N_12615);
or U12760 (N_12760,N_12557,N_12582);
nand U12761 (N_12761,N_12550,N_12502);
and U12762 (N_12762,N_12547,N_12536);
xnor U12763 (N_12763,N_12662,N_12583);
xnor U12764 (N_12764,N_12545,N_12569);
xnor U12765 (N_12765,N_12650,N_12509);
and U12766 (N_12766,N_12725,N_12519);
nand U12767 (N_12767,N_12713,N_12741);
or U12768 (N_12768,N_12588,N_12686);
and U12769 (N_12769,N_12571,N_12566);
nand U12770 (N_12770,N_12620,N_12609);
and U12771 (N_12771,N_12556,N_12714);
and U12772 (N_12772,N_12638,N_12653);
nor U12773 (N_12773,N_12539,N_12549);
or U12774 (N_12774,N_12711,N_12702);
or U12775 (N_12775,N_12601,N_12734);
nor U12776 (N_12776,N_12621,N_12712);
xnor U12777 (N_12777,N_12561,N_12529);
or U12778 (N_12778,N_12572,N_12612);
and U12779 (N_12779,N_12727,N_12581);
nand U12780 (N_12780,N_12693,N_12590);
nand U12781 (N_12781,N_12507,N_12733);
nand U12782 (N_12782,N_12591,N_12523);
xnor U12783 (N_12783,N_12701,N_12640);
or U12784 (N_12784,N_12520,N_12522);
or U12785 (N_12785,N_12739,N_12697);
and U12786 (N_12786,N_12512,N_12500);
or U12787 (N_12787,N_12565,N_12614);
nor U12788 (N_12788,N_12674,N_12746);
or U12789 (N_12789,N_12553,N_12552);
xor U12790 (N_12790,N_12651,N_12732);
and U12791 (N_12791,N_12532,N_12664);
or U12792 (N_12792,N_12544,N_12625);
or U12793 (N_12793,N_12682,N_12709);
nand U12794 (N_12794,N_12635,N_12528);
and U12795 (N_12795,N_12575,N_12542);
and U12796 (N_12796,N_12629,N_12681);
or U12797 (N_12797,N_12623,N_12698);
or U12798 (N_12798,N_12579,N_12728);
or U12799 (N_12799,N_12587,N_12619);
xor U12800 (N_12800,N_12645,N_12658);
nand U12801 (N_12801,N_12597,N_12505);
nand U12802 (N_12802,N_12576,N_12726);
nor U12803 (N_12803,N_12548,N_12652);
nor U12804 (N_12804,N_12639,N_12604);
nor U12805 (N_12805,N_12517,N_12724);
nor U12806 (N_12806,N_12666,N_12624);
nand U12807 (N_12807,N_12524,N_12718);
xor U12808 (N_12808,N_12628,N_12663);
or U12809 (N_12809,N_12596,N_12670);
xnor U12810 (N_12810,N_12568,N_12616);
nand U12811 (N_12811,N_12655,N_12715);
xnor U12812 (N_12812,N_12634,N_12649);
or U12813 (N_12813,N_12703,N_12515);
xnor U12814 (N_12814,N_12690,N_12630);
xor U12815 (N_12815,N_12659,N_12667);
nand U12816 (N_12816,N_12538,N_12656);
nor U12817 (N_12817,N_12541,N_12593);
xor U12818 (N_12818,N_12647,N_12503);
or U12819 (N_12819,N_12744,N_12683);
or U12820 (N_12820,N_12720,N_12748);
nor U12821 (N_12821,N_12560,N_12595);
nor U12822 (N_12822,N_12736,N_12525);
nor U12823 (N_12823,N_12501,N_12511);
nor U12824 (N_12824,N_12513,N_12742);
and U12825 (N_12825,N_12680,N_12564);
and U12826 (N_12826,N_12694,N_12584);
nor U12827 (N_12827,N_12695,N_12745);
nand U12828 (N_12828,N_12688,N_12673);
and U12829 (N_12829,N_12578,N_12618);
or U12830 (N_12830,N_12735,N_12675);
nor U12831 (N_12831,N_12531,N_12710);
nor U12832 (N_12832,N_12617,N_12622);
nand U12833 (N_12833,N_12506,N_12643);
nor U12834 (N_12834,N_12665,N_12669);
and U12835 (N_12835,N_12692,N_12671);
nand U12836 (N_12836,N_12535,N_12716);
or U12837 (N_12837,N_12696,N_12642);
or U12838 (N_12838,N_12546,N_12705);
nand U12839 (N_12839,N_12626,N_12534);
or U12840 (N_12840,N_12648,N_12677);
nor U12841 (N_12841,N_12592,N_12719);
or U12842 (N_12842,N_12721,N_12599);
xor U12843 (N_12843,N_12685,N_12530);
nand U12844 (N_12844,N_12608,N_12737);
or U12845 (N_12845,N_12700,N_12585);
nor U12846 (N_12846,N_12504,N_12577);
nor U12847 (N_12847,N_12526,N_12521);
and U12848 (N_12848,N_12644,N_12699);
xor U12849 (N_12849,N_12633,N_12738);
xnor U12850 (N_12850,N_12707,N_12678);
or U12851 (N_12851,N_12613,N_12518);
or U12852 (N_12852,N_12508,N_12605);
or U12853 (N_12853,N_12627,N_12676);
or U12854 (N_12854,N_12563,N_12722);
xnor U12855 (N_12855,N_12740,N_12706);
nor U12856 (N_12856,N_12631,N_12729);
and U12857 (N_12857,N_12747,N_12749);
or U12858 (N_12858,N_12555,N_12657);
and U12859 (N_12859,N_12562,N_12586);
nor U12860 (N_12860,N_12723,N_12533);
xor U12861 (N_12861,N_12684,N_12567);
or U12862 (N_12862,N_12646,N_12607);
or U12863 (N_12863,N_12641,N_12527);
xnor U12864 (N_12864,N_12731,N_12514);
and U12865 (N_12865,N_12540,N_12559);
nand U12866 (N_12866,N_12660,N_12632);
nand U12867 (N_12867,N_12600,N_12589);
nor U12868 (N_12868,N_12594,N_12689);
or U12869 (N_12869,N_12554,N_12661);
xor U12870 (N_12870,N_12602,N_12704);
xnor U12871 (N_12871,N_12668,N_12543);
and U12872 (N_12872,N_12537,N_12743);
or U12873 (N_12873,N_12691,N_12574);
nor U12874 (N_12874,N_12637,N_12679);
and U12875 (N_12875,N_12562,N_12728);
xnor U12876 (N_12876,N_12703,N_12502);
xor U12877 (N_12877,N_12616,N_12703);
or U12878 (N_12878,N_12685,N_12553);
and U12879 (N_12879,N_12717,N_12615);
xnor U12880 (N_12880,N_12647,N_12600);
and U12881 (N_12881,N_12723,N_12566);
nand U12882 (N_12882,N_12530,N_12533);
xor U12883 (N_12883,N_12547,N_12637);
xor U12884 (N_12884,N_12659,N_12672);
or U12885 (N_12885,N_12550,N_12600);
nor U12886 (N_12886,N_12514,N_12526);
nor U12887 (N_12887,N_12677,N_12681);
xor U12888 (N_12888,N_12502,N_12715);
nor U12889 (N_12889,N_12727,N_12630);
or U12890 (N_12890,N_12639,N_12694);
xnor U12891 (N_12891,N_12552,N_12538);
or U12892 (N_12892,N_12691,N_12724);
xor U12893 (N_12893,N_12679,N_12623);
nand U12894 (N_12894,N_12719,N_12529);
and U12895 (N_12895,N_12698,N_12576);
nand U12896 (N_12896,N_12710,N_12530);
nor U12897 (N_12897,N_12713,N_12654);
nor U12898 (N_12898,N_12685,N_12593);
nor U12899 (N_12899,N_12516,N_12701);
or U12900 (N_12900,N_12668,N_12640);
and U12901 (N_12901,N_12530,N_12612);
xnor U12902 (N_12902,N_12614,N_12670);
or U12903 (N_12903,N_12741,N_12653);
xor U12904 (N_12904,N_12547,N_12511);
xnor U12905 (N_12905,N_12574,N_12628);
or U12906 (N_12906,N_12698,N_12537);
and U12907 (N_12907,N_12628,N_12664);
nand U12908 (N_12908,N_12521,N_12540);
nor U12909 (N_12909,N_12535,N_12686);
nand U12910 (N_12910,N_12654,N_12532);
or U12911 (N_12911,N_12612,N_12714);
and U12912 (N_12912,N_12633,N_12547);
nand U12913 (N_12913,N_12716,N_12654);
or U12914 (N_12914,N_12742,N_12605);
nor U12915 (N_12915,N_12723,N_12526);
or U12916 (N_12916,N_12599,N_12594);
and U12917 (N_12917,N_12692,N_12613);
and U12918 (N_12918,N_12700,N_12645);
or U12919 (N_12919,N_12581,N_12571);
and U12920 (N_12920,N_12589,N_12585);
nor U12921 (N_12921,N_12552,N_12716);
nand U12922 (N_12922,N_12601,N_12508);
and U12923 (N_12923,N_12608,N_12686);
xnor U12924 (N_12924,N_12576,N_12521);
nand U12925 (N_12925,N_12629,N_12633);
nand U12926 (N_12926,N_12576,N_12711);
or U12927 (N_12927,N_12726,N_12743);
or U12928 (N_12928,N_12659,N_12504);
and U12929 (N_12929,N_12746,N_12547);
xnor U12930 (N_12930,N_12575,N_12506);
nor U12931 (N_12931,N_12550,N_12526);
nor U12932 (N_12932,N_12687,N_12696);
nand U12933 (N_12933,N_12724,N_12580);
and U12934 (N_12934,N_12690,N_12721);
nor U12935 (N_12935,N_12697,N_12656);
nand U12936 (N_12936,N_12541,N_12685);
xnor U12937 (N_12937,N_12741,N_12674);
or U12938 (N_12938,N_12706,N_12748);
xnor U12939 (N_12939,N_12732,N_12713);
xnor U12940 (N_12940,N_12502,N_12714);
or U12941 (N_12941,N_12580,N_12643);
nor U12942 (N_12942,N_12723,N_12628);
and U12943 (N_12943,N_12519,N_12631);
and U12944 (N_12944,N_12722,N_12664);
nor U12945 (N_12945,N_12523,N_12562);
or U12946 (N_12946,N_12677,N_12539);
nand U12947 (N_12947,N_12746,N_12506);
nor U12948 (N_12948,N_12566,N_12506);
nor U12949 (N_12949,N_12567,N_12738);
or U12950 (N_12950,N_12531,N_12628);
and U12951 (N_12951,N_12602,N_12630);
or U12952 (N_12952,N_12533,N_12684);
and U12953 (N_12953,N_12665,N_12581);
nand U12954 (N_12954,N_12711,N_12526);
or U12955 (N_12955,N_12567,N_12579);
nor U12956 (N_12956,N_12605,N_12529);
or U12957 (N_12957,N_12748,N_12687);
and U12958 (N_12958,N_12740,N_12651);
and U12959 (N_12959,N_12740,N_12519);
nor U12960 (N_12960,N_12517,N_12646);
or U12961 (N_12961,N_12564,N_12678);
nand U12962 (N_12962,N_12631,N_12656);
and U12963 (N_12963,N_12518,N_12729);
and U12964 (N_12964,N_12553,N_12647);
and U12965 (N_12965,N_12742,N_12686);
nor U12966 (N_12966,N_12739,N_12606);
nand U12967 (N_12967,N_12503,N_12556);
nand U12968 (N_12968,N_12731,N_12726);
or U12969 (N_12969,N_12621,N_12726);
or U12970 (N_12970,N_12743,N_12720);
xor U12971 (N_12971,N_12527,N_12543);
xnor U12972 (N_12972,N_12529,N_12665);
and U12973 (N_12973,N_12688,N_12566);
nor U12974 (N_12974,N_12608,N_12747);
xnor U12975 (N_12975,N_12739,N_12524);
xnor U12976 (N_12976,N_12504,N_12501);
or U12977 (N_12977,N_12638,N_12522);
xor U12978 (N_12978,N_12629,N_12648);
nor U12979 (N_12979,N_12656,N_12514);
nand U12980 (N_12980,N_12644,N_12596);
nand U12981 (N_12981,N_12648,N_12532);
or U12982 (N_12982,N_12588,N_12551);
and U12983 (N_12983,N_12744,N_12589);
xnor U12984 (N_12984,N_12502,N_12729);
nand U12985 (N_12985,N_12579,N_12505);
xor U12986 (N_12986,N_12523,N_12712);
nor U12987 (N_12987,N_12580,N_12717);
nand U12988 (N_12988,N_12507,N_12655);
nor U12989 (N_12989,N_12707,N_12658);
or U12990 (N_12990,N_12501,N_12500);
nand U12991 (N_12991,N_12652,N_12522);
nand U12992 (N_12992,N_12507,N_12644);
nor U12993 (N_12993,N_12705,N_12732);
nand U12994 (N_12994,N_12536,N_12684);
xor U12995 (N_12995,N_12721,N_12614);
xor U12996 (N_12996,N_12556,N_12532);
and U12997 (N_12997,N_12594,N_12669);
xnor U12998 (N_12998,N_12643,N_12523);
nand U12999 (N_12999,N_12573,N_12639);
and U13000 (N_13000,N_12913,N_12846);
or U13001 (N_13001,N_12863,N_12988);
nand U13002 (N_13002,N_12902,N_12932);
nor U13003 (N_13003,N_12948,N_12969);
and U13004 (N_13004,N_12965,N_12938);
xnor U13005 (N_13005,N_12839,N_12873);
and U13006 (N_13006,N_12981,N_12882);
nand U13007 (N_13007,N_12867,N_12996);
and U13008 (N_13008,N_12957,N_12876);
nand U13009 (N_13009,N_12827,N_12764);
or U13010 (N_13010,N_12844,N_12755);
and U13011 (N_13011,N_12833,N_12875);
or U13012 (N_13012,N_12900,N_12884);
xor U13013 (N_13013,N_12872,N_12776);
and U13014 (N_13014,N_12992,N_12923);
nor U13015 (N_13015,N_12877,N_12917);
or U13016 (N_13016,N_12958,N_12936);
and U13017 (N_13017,N_12920,N_12836);
or U13018 (N_13018,N_12995,N_12999);
nand U13019 (N_13019,N_12780,N_12823);
nor U13020 (N_13020,N_12950,N_12960);
xor U13021 (N_13021,N_12757,N_12997);
and U13022 (N_13022,N_12942,N_12753);
or U13023 (N_13023,N_12750,N_12811);
xor U13024 (N_13024,N_12962,N_12946);
and U13025 (N_13025,N_12794,N_12987);
or U13026 (N_13026,N_12984,N_12982);
and U13027 (N_13027,N_12929,N_12849);
and U13028 (N_13028,N_12881,N_12928);
xor U13029 (N_13029,N_12765,N_12752);
or U13030 (N_13030,N_12887,N_12908);
nor U13031 (N_13031,N_12799,N_12885);
nand U13032 (N_13032,N_12842,N_12864);
nand U13033 (N_13033,N_12904,N_12991);
nor U13034 (N_13034,N_12985,N_12859);
xor U13035 (N_13035,N_12855,N_12933);
nand U13036 (N_13036,N_12898,N_12800);
or U13037 (N_13037,N_12886,N_12801);
and U13038 (N_13038,N_12993,N_12935);
or U13039 (N_13039,N_12767,N_12769);
and U13040 (N_13040,N_12869,N_12955);
and U13041 (N_13041,N_12857,N_12921);
or U13042 (N_13042,N_12834,N_12854);
xor U13043 (N_13043,N_12952,N_12943);
or U13044 (N_13044,N_12968,N_12813);
nor U13045 (N_13045,N_12840,N_12761);
nor U13046 (N_13046,N_12797,N_12848);
xor U13047 (N_13047,N_12889,N_12994);
or U13048 (N_13048,N_12934,N_12922);
or U13049 (N_13049,N_12914,N_12961);
and U13050 (N_13050,N_12810,N_12916);
and U13051 (N_13051,N_12878,N_12816);
nor U13052 (N_13052,N_12819,N_12828);
nor U13053 (N_13053,N_12911,N_12861);
nor U13054 (N_13054,N_12959,N_12870);
or U13055 (N_13055,N_12924,N_12835);
nor U13056 (N_13056,N_12807,N_12894);
xnor U13057 (N_13057,N_12975,N_12758);
or U13058 (N_13058,N_12785,N_12815);
nand U13059 (N_13059,N_12927,N_12754);
nor U13060 (N_13060,N_12830,N_12788);
nor U13061 (N_13061,N_12970,N_12897);
nor U13062 (N_13062,N_12890,N_12817);
nand U13063 (N_13063,N_12760,N_12778);
xor U13064 (N_13064,N_12947,N_12820);
nand U13065 (N_13065,N_12998,N_12803);
xor U13066 (N_13066,N_12806,N_12845);
nand U13067 (N_13067,N_12901,N_12847);
or U13068 (N_13068,N_12805,N_12774);
nand U13069 (N_13069,N_12903,N_12974);
nor U13070 (N_13070,N_12852,N_12972);
nor U13071 (N_13071,N_12796,N_12931);
nor U13072 (N_13072,N_12787,N_12909);
nand U13073 (N_13073,N_12910,N_12953);
nor U13074 (N_13074,N_12763,N_12808);
and U13075 (N_13075,N_12895,N_12971);
and U13076 (N_13076,N_12851,N_12779);
or U13077 (N_13077,N_12980,N_12989);
xnor U13078 (N_13078,N_12777,N_12949);
nor U13079 (N_13079,N_12966,N_12918);
xor U13080 (N_13080,N_12751,N_12814);
nor U13081 (N_13081,N_12809,N_12892);
and U13082 (N_13082,N_12944,N_12945);
or U13083 (N_13083,N_12896,N_12979);
nor U13084 (N_13084,N_12899,N_12940);
nor U13085 (N_13085,N_12825,N_12926);
and U13086 (N_13086,N_12919,N_12838);
nand U13087 (N_13087,N_12858,N_12866);
or U13088 (N_13088,N_12783,N_12762);
and U13089 (N_13089,N_12853,N_12860);
xor U13090 (N_13090,N_12791,N_12963);
and U13091 (N_13091,N_12812,N_12951);
xnor U13092 (N_13092,N_12781,N_12880);
or U13093 (N_13093,N_12990,N_12804);
nor U13094 (N_13094,N_12891,N_12802);
nand U13095 (N_13095,N_12826,N_12879);
and U13096 (N_13096,N_12850,N_12862);
and U13097 (N_13097,N_12865,N_12956);
nand U13098 (N_13098,N_12930,N_12954);
nor U13099 (N_13099,N_12907,N_12789);
nor U13100 (N_13100,N_12888,N_12795);
nor U13101 (N_13101,N_12977,N_12983);
xor U13102 (N_13102,N_12906,N_12868);
and U13103 (N_13103,N_12768,N_12772);
and U13104 (N_13104,N_12883,N_12837);
nor U13105 (N_13105,N_12784,N_12832);
xor U13106 (N_13106,N_12905,N_12871);
or U13107 (N_13107,N_12798,N_12831);
nand U13108 (N_13108,N_12782,N_12937);
and U13109 (N_13109,N_12915,N_12964);
xnor U13110 (N_13110,N_12976,N_12756);
nand U13111 (N_13111,N_12821,N_12978);
xor U13112 (N_13112,N_12967,N_12792);
nor U13113 (N_13113,N_12824,N_12759);
and U13114 (N_13114,N_12766,N_12843);
nand U13115 (N_13115,N_12770,N_12939);
nand U13116 (N_13116,N_12874,N_12912);
and U13117 (N_13117,N_12941,N_12925);
and U13118 (N_13118,N_12818,N_12856);
or U13119 (N_13119,N_12773,N_12775);
nor U13120 (N_13120,N_12771,N_12790);
and U13121 (N_13121,N_12786,N_12822);
or U13122 (N_13122,N_12793,N_12973);
xnor U13123 (N_13123,N_12829,N_12986);
and U13124 (N_13124,N_12841,N_12893);
and U13125 (N_13125,N_12891,N_12985);
and U13126 (N_13126,N_12962,N_12765);
xnor U13127 (N_13127,N_12935,N_12985);
and U13128 (N_13128,N_12894,N_12757);
or U13129 (N_13129,N_12989,N_12982);
xor U13130 (N_13130,N_12940,N_12987);
nor U13131 (N_13131,N_12889,N_12881);
or U13132 (N_13132,N_12836,N_12793);
xnor U13133 (N_13133,N_12783,N_12811);
nand U13134 (N_13134,N_12973,N_12937);
and U13135 (N_13135,N_12833,N_12845);
nand U13136 (N_13136,N_12952,N_12926);
and U13137 (N_13137,N_12824,N_12815);
and U13138 (N_13138,N_12959,N_12830);
or U13139 (N_13139,N_12929,N_12754);
xnor U13140 (N_13140,N_12833,N_12998);
xnor U13141 (N_13141,N_12877,N_12787);
and U13142 (N_13142,N_12818,N_12858);
or U13143 (N_13143,N_12824,N_12849);
and U13144 (N_13144,N_12884,N_12894);
or U13145 (N_13145,N_12953,N_12784);
nand U13146 (N_13146,N_12826,N_12918);
or U13147 (N_13147,N_12821,N_12858);
or U13148 (N_13148,N_12882,N_12993);
or U13149 (N_13149,N_12768,N_12998);
nand U13150 (N_13150,N_12893,N_12997);
xnor U13151 (N_13151,N_12798,N_12936);
or U13152 (N_13152,N_12930,N_12780);
or U13153 (N_13153,N_12957,N_12754);
or U13154 (N_13154,N_12826,N_12921);
xor U13155 (N_13155,N_12989,N_12993);
nand U13156 (N_13156,N_12928,N_12829);
and U13157 (N_13157,N_12953,N_12825);
or U13158 (N_13158,N_12879,N_12965);
nor U13159 (N_13159,N_12753,N_12926);
nand U13160 (N_13160,N_12999,N_12936);
nor U13161 (N_13161,N_12904,N_12788);
and U13162 (N_13162,N_12792,N_12966);
and U13163 (N_13163,N_12823,N_12953);
nand U13164 (N_13164,N_12781,N_12969);
or U13165 (N_13165,N_12985,N_12816);
or U13166 (N_13166,N_12887,N_12834);
xor U13167 (N_13167,N_12945,N_12876);
nor U13168 (N_13168,N_12789,N_12970);
and U13169 (N_13169,N_12965,N_12815);
nor U13170 (N_13170,N_12947,N_12809);
and U13171 (N_13171,N_12819,N_12786);
or U13172 (N_13172,N_12827,N_12919);
nand U13173 (N_13173,N_12834,N_12838);
nor U13174 (N_13174,N_12890,N_12946);
and U13175 (N_13175,N_12890,N_12990);
and U13176 (N_13176,N_12889,N_12885);
nor U13177 (N_13177,N_12794,N_12955);
nor U13178 (N_13178,N_12872,N_12939);
and U13179 (N_13179,N_12977,N_12789);
and U13180 (N_13180,N_12840,N_12898);
nor U13181 (N_13181,N_12855,N_12931);
nand U13182 (N_13182,N_12939,N_12844);
nor U13183 (N_13183,N_12915,N_12780);
or U13184 (N_13184,N_12874,N_12989);
nor U13185 (N_13185,N_12811,N_12764);
or U13186 (N_13186,N_12990,N_12869);
or U13187 (N_13187,N_12922,N_12897);
nand U13188 (N_13188,N_12923,N_12826);
xnor U13189 (N_13189,N_12828,N_12922);
xnor U13190 (N_13190,N_12770,N_12840);
nor U13191 (N_13191,N_12986,N_12921);
xor U13192 (N_13192,N_12816,N_12798);
nand U13193 (N_13193,N_12854,N_12944);
or U13194 (N_13194,N_12793,N_12878);
xnor U13195 (N_13195,N_12898,N_12875);
or U13196 (N_13196,N_12953,N_12796);
xor U13197 (N_13197,N_12899,N_12852);
xnor U13198 (N_13198,N_12791,N_12850);
nand U13199 (N_13199,N_12899,N_12818);
and U13200 (N_13200,N_12965,N_12801);
or U13201 (N_13201,N_12785,N_12819);
or U13202 (N_13202,N_12834,N_12859);
xnor U13203 (N_13203,N_12966,N_12973);
xor U13204 (N_13204,N_12901,N_12751);
or U13205 (N_13205,N_12891,N_12852);
nor U13206 (N_13206,N_12784,N_12910);
or U13207 (N_13207,N_12872,N_12818);
or U13208 (N_13208,N_12905,N_12967);
xor U13209 (N_13209,N_12932,N_12892);
nor U13210 (N_13210,N_12829,N_12931);
nand U13211 (N_13211,N_12931,N_12819);
nand U13212 (N_13212,N_12909,N_12833);
and U13213 (N_13213,N_12815,N_12996);
or U13214 (N_13214,N_12752,N_12901);
and U13215 (N_13215,N_12782,N_12961);
xor U13216 (N_13216,N_12780,N_12893);
and U13217 (N_13217,N_12878,N_12982);
and U13218 (N_13218,N_12855,N_12980);
and U13219 (N_13219,N_12985,N_12817);
or U13220 (N_13220,N_12763,N_12812);
nand U13221 (N_13221,N_12995,N_12868);
nand U13222 (N_13222,N_12975,N_12790);
or U13223 (N_13223,N_12871,N_12790);
and U13224 (N_13224,N_12796,N_12867);
or U13225 (N_13225,N_12884,N_12759);
nand U13226 (N_13226,N_12799,N_12761);
xor U13227 (N_13227,N_12820,N_12924);
nor U13228 (N_13228,N_12912,N_12915);
nand U13229 (N_13229,N_12857,N_12996);
nor U13230 (N_13230,N_12998,N_12951);
and U13231 (N_13231,N_12870,N_12957);
xor U13232 (N_13232,N_12857,N_12830);
or U13233 (N_13233,N_12792,N_12870);
xnor U13234 (N_13234,N_12965,N_12884);
xor U13235 (N_13235,N_12855,N_12959);
nand U13236 (N_13236,N_12797,N_12920);
or U13237 (N_13237,N_12910,N_12886);
nor U13238 (N_13238,N_12965,N_12845);
nor U13239 (N_13239,N_12788,N_12902);
and U13240 (N_13240,N_12852,N_12927);
or U13241 (N_13241,N_12770,N_12769);
and U13242 (N_13242,N_12927,N_12946);
and U13243 (N_13243,N_12835,N_12964);
nor U13244 (N_13244,N_12872,N_12843);
or U13245 (N_13245,N_12803,N_12929);
xnor U13246 (N_13246,N_12788,N_12996);
xor U13247 (N_13247,N_12933,N_12987);
and U13248 (N_13248,N_12904,N_12856);
nor U13249 (N_13249,N_12990,N_12904);
or U13250 (N_13250,N_13170,N_13152);
nand U13251 (N_13251,N_13133,N_13234);
or U13252 (N_13252,N_13168,N_13218);
nand U13253 (N_13253,N_13182,N_13031);
and U13254 (N_13254,N_13085,N_13070);
nor U13255 (N_13255,N_13221,N_13057);
nor U13256 (N_13256,N_13173,N_13093);
and U13257 (N_13257,N_13224,N_13248);
or U13258 (N_13258,N_13108,N_13016);
and U13259 (N_13259,N_13112,N_13180);
nor U13260 (N_13260,N_13008,N_13179);
nand U13261 (N_13261,N_13190,N_13134);
nor U13262 (N_13262,N_13153,N_13096);
and U13263 (N_13263,N_13088,N_13158);
xnor U13264 (N_13264,N_13147,N_13155);
nand U13265 (N_13265,N_13172,N_13222);
and U13266 (N_13266,N_13240,N_13056);
nor U13267 (N_13267,N_13192,N_13074);
xnor U13268 (N_13268,N_13103,N_13200);
nor U13269 (N_13269,N_13142,N_13051);
xor U13270 (N_13270,N_13012,N_13003);
nand U13271 (N_13271,N_13052,N_13166);
or U13272 (N_13272,N_13117,N_13061);
xor U13273 (N_13273,N_13092,N_13191);
or U13274 (N_13274,N_13111,N_13073);
nor U13275 (N_13275,N_13014,N_13068);
nor U13276 (N_13276,N_13027,N_13163);
nor U13277 (N_13277,N_13030,N_13019);
nor U13278 (N_13278,N_13042,N_13135);
xor U13279 (N_13279,N_13232,N_13069);
nand U13280 (N_13280,N_13000,N_13001);
or U13281 (N_13281,N_13032,N_13138);
nor U13282 (N_13282,N_13087,N_13165);
or U13283 (N_13283,N_13102,N_13143);
nor U13284 (N_13284,N_13037,N_13215);
or U13285 (N_13285,N_13109,N_13053);
nand U13286 (N_13286,N_13207,N_13214);
or U13287 (N_13287,N_13004,N_13178);
nand U13288 (N_13288,N_13022,N_13098);
and U13289 (N_13289,N_13212,N_13033);
nand U13290 (N_13290,N_13047,N_13148);
nand U13291 (N_13291,N_13038,N_13078);
and U13292 (N_13292,N_13020,N_13169);
and U13293 (N_13293,N_13045,N_13136);
nand U13294 (N_13294,N_13041,N_13246);
nor U13295 (N_13295,N_13089,N_13036);
or U13296 (N_13296,N_13116,N_13189);
and U13297 (N_13297,N_13177,N_13125);
nor U13298 (N_13298,N_13137,N_13225);
and U13299 (N_13299,N_13006,N_13100);
and U13300 (N_13300,N_13118,N_13231);
and U13301 (N_13301,N_13219,N_13079);
or U13302 (N_13302,N_13119,N_13216);
xor U13303 (N_13303,N_13198,N_13241);
nor U13304 (N_13304,N_13059,N_13181);
nor U13305 (N_13305,N_13186,N_13115);
nand U13306 (N_13306,N_13199,N_13164);
nor U13307 (N_13307,N_13120,N_13196);
nand U13308 (N_13308,N_13054,N_13249);
nor U13309 (N_13309,N_13245,N_13151);
and U13310 (N_13310,N_13082,N_13028);
xor U13311 (N_13311,N_13201,N_13140);
or U13312 (N_13312,N_13127,N_13065);
nor U13313 (N_13313,N_13139,N_13183);
nand U13314 (N_13314,N_13145,N_13185);
nand U13315 (N_13315,N_13066,N_13113);
and U13316 (N_13316,N_13007,N_13050);
and U13317 (N_13317,N_13205,N_13097);
and U13318 (N_13318,N_13157,N_13105);
xnor U13319 (N_13319,N_13141,N_13247);
nand U13320 (N_13320,N_13058,N_13086);
nand U13321 (N_13321,N_13084,N_13174);
nor U13322 (N_13322,N_13130,N_13203);
xor U13323 (N_13323,N_13154,N_13067);
xor U13324 (N_13324,N_13126,N_13043);
nor U13325 (N_13325,N_13076,N_13062);
xnor U13326 (N_13326,N_13211,N_13023);
or U13327 (N_13327,N_13159,N_13220);
xor U13328 (N_13328,N_13226,N_13077);
xor U13329 (N_13329,N_13167,N_13040);
or U13330 (N_13330,N_13081,N_13204);
nor U13331 (N_13331,N_13160,N_13121);
xnor U13332 (N_13332,N_13099,N_13029);
nand U13333 (N_13333,N_13094,N_13015);
or U13334 (N_13334,N_13090,N_13146);
or U13335 (N_13335,N_13026,N_13188);
or U13336 (N_13336,N_13128,N_13018);
nor U13337 (N_13337,N_13110,N_13083);
and U13338 (N_13338,N_13044,N_13104);
and U13339 (N_13339,N_13176,N_13239);
nand U13340 (N_13340,N_13197,N_13024);
and U13341 (N_13341,N_13123,N_13237);
and U13342 (N_13342,N_13209,N_13161);
nor U13343 (N_13343,N_13049,N_13064);
nand U13344 (N_13344,N_13171,N_13242);
nor U13345 (N_13345,N_13005,N_13213);
xnor U13346 (N_13346,N_13010,N_13114);
and U13347 (N_13347,N_13101,N_13144);
nand U13348 (N_13348,N_13075,N_13236);
nand U13349 (N_13349,N_13039,N_13095);
nor U13350 (N_13350,N_13063,N_13129);
xor U13351 (N_13351,N_13150,N_13208);
xor U13352 (N_13352,N_13046,N_13187);
nor U13353 (N_13353,N_13048,N_13210);
and U13354 (N_13354,N_13235,N_13217);
xor U13355 (N_13355,N_13233,N_13080);
and U13356 (N_13356,N_13107,N_13021);
or U13357 (N_13357,N_13230,N_13122);
xnor U13358 (N_13358,N_13002,N_13206);
xnor U13359 (N_13359,N_13244,N_13132);
nand U13360 (N_13360,N_13195,N_13156);
nor U13361 (N_13361,N_13091,N_13223);
nand U13362 (N_13362,N_13071,N_13193);
and U13363 (N_13363,N_13013,N_13227);
and U13364 (N_13364,N_13162,N_13106);
nor U13365 (N_13365,N_13072,N_13149);
nand U13366 (N_13366,N_13243,N_13238);
nor U13367 (N_13367,N_13034,N_13194);
and U13368 (N_13368,N_13175,N_13202);
nor U13369 (N_13369,N_13011,N_13131);
and U13370 (N_13370,N_13184,N_13228);
or U13371 (N_13371,N_13124,N_13060);
nand U13372 (N_13372,N_13009,N_13035);
nand U13373 (N_13373,N_13017,N_13229);
xor U13374 (N_13374,N_13055,N_13025);
nand U13375 (N_13375,N_13155,N_13237);
and U13376 (N_13376,N_13228,N_13066);
xnor U13377 (N_13377,N_13205,N_13086);
nand U13378 (N_13378,N_13076,N_13053);
nor U13379 (N_13379,N_13029,N_13157);
or U13380 (N_13380,N_13088,N_13134);
nand U13381 (N_13381,N_13089,N_13000);
nand U13382 (N_13382,N_13042,N_13027);
nor U13383 (N_13383,N_13015,N_13231);
xnor U13384 (N_13384,N_13177,N_13140);
or U13385 (N_13385,N_13226,N_13021);
nor U13386 (N_13386,N_13028,N_13229);
nor U13387 (N_13387,N_13191,N_13233);
or U13388 (N_13388,N_13127,N_13134);
or U13389 (N_13389,N_13125,N_13007);
nor U13390 (N_13390,N_13144,N_13206);
nor U13391 (N_13391,N_13035,N_13022);
xor U13392 (N_13392,N_13071,N_13014);
nand U13393 (N_13393,N_13248,N_13110);
or U13394 (N_13394,N_13075,N_13093);
xnor U13395 (N_13395,N_13065,N_13169);
or U13396 (N_13396,N_13109,N_13082);
nand U13397 (N_13397,N_13132,N_13140);
nor U13398 (N_13398,N_13143,N_13139);
nand U13399 (N_13399,N_13132,N_13137);
or U13400 (N_13400,N_13049,N_13067);
nor U13401 (N_13401,N_13218,N_13050);
nand U13402 (N_13402,N_13207,N_13155);
xor U13403 (N_13403,N_13022,N_13070);
and U13404 (N_13404,N_13032,N_13196);
xnor U13405 (N_13405,N_13053,N_13239);
nand U13406 (N_13406,N_13139,N_13165);
nand U13407 (N_13407,N_13039,N_13019);
or U13408 (N_13408,N_13025,N_13053);
nor U13409 (N_13409,N_13070,N_13182);
nor U13410 (N_13410,N_13198,N_13224);
nand U13411 (N_13411,N_13047,N_13103);
or U13412 (N_13412,N_13140,N_13049);
or U13413 (N_13413,N_13038,N_13054);
or U13414 (N_13414,N_13110,N_13004);
nor U13415 (N_13415,N_13218,N_13148);
nand U13416 (N_13416,N_13231,N_13053);
or U13417 (N_13417,N_13140,N_13191);
or U13418 (N_13418,N_13241,N_13179);
and U13419 (N_13419,N_13095,N_13099);
xnor U13420 (N_13420,N_13154,N_13229);
xnor U13421 (N_13421,N_13152,N_13017);
nand U13422 (N_13422,N_13020,N_13077);
xnor U13423 (N_13423,N_13199,N_13030);
or U13424 (N_13424,N_13104,N_13056);
and U13425 (N_13425,N_13064,N_13176);
nand U13426 (N_13426,N_13235,N_13030);
and U13427 (N_13427,N_13059,N_13214);
xor U13428 (N_13428,N_13151,N_13230);
nand U13429 (N_13429,N_13001,N_13016);
or U13430 (N_13430,N_13235,N_13089);
nand U13431 (N_13431,N_13199,N_13144);
and U13432 (N_13432,N_13033,N_13221);
nand U13433 (N_13433,N_13124,N_13171);
or U13434 (N_13434,N_13062,N_13128);
nand U13435 (N_13435,N_13172,N_13125);
and U13436 (N_13436,N_13135,N_13248);
and U13437 (N_13437,N_13213,N_13030);
nor U13438 (N_13438,N_13172,N_13003);
nand U13439 (N_13439,N_13109,N_13013);
nand U13440 (N_13440,N_13160,N_13143);
and U13441 (N_13441,N_13137,N_13243);
or U13442 (N_13442,N_13058,N_13129);
and U13443 (N_13443,N_13124,N_13011);
nand U13444 (N_13444,N_13171,N_13075);
xnor U13445 (N_13445,N_13032,N_13021);
xnor U13446 (N_13446,N_13109,N_13112);
xor U13447 (N_13447,N_13128,N_13086);
nor U13448 (N_13448,N_13223,N_13143);
or U13449 (N_13449,N_13090,N_13156);
nor U13450 (N_13450,N_13019,N_13137);
nor U13451 (N_13451,N_13090,N_13064);
nand U13452 (N_13452,N_13074,N_13213);
or U13453 (N_13453,N_13041,N_13156);
xnor U13454 (N_13454,N_13156,N_13089);
xnor U13455 (N_13455,N_13222,N_13199);
xor U13456 (N_13456,N_13165,N_13146);
nand U13457 (N_13457,N_13095,N_13156);
nor U13458 (N_13458,N_13192,N_13190);
xnor U13459 (N_13459,N_13176,N_13164);
xnor U13460 (N_13460,N_13009,N_13224);
or U13461 (N_13461,N_13101,N_13098);
nand U13462 (N_13462,N_13224,N_13139);
and U13463 (N_13463,N_13169,N_13090);
or U13464 (N_13464,N_13225,N_13105);
or U13465 (N_13465,N_13111,N_13115);
nand U13466 (N_13466,N_13190,N_13011);
and U13467 (N_13467,N_13128,N_13031);
and U13468 (N_13468,N_13209,N_13114);
or U13469 (N_13469,N_13064,N_13127);
or U13470 (N_13470,N_13015,N_13173);
nand U13471 (N_13471,N_13127,N_13221);
xnor U13472 (N_13472,N_13210,N_13239);
and U13473 (N_13473,N_13190,N_13010);
and U13474 (N_13474,N_13104,N_13030);
nand U13475 (N_13475,N_13224,N_13023);
nand U13476 (N_13476,N_13083,N_13018);
nor U13477 (N_13477,N_13094,N_13061);
nor U13478 (N_13478,N_13181,N_13209);
xor U13479 (N_13479,N_13121,N_13147);
and U13480 (N_13480,N_13026,N_13152);
xnor U13481 (N_13481,N_13225,N_13136);
xnor U13482 (N_13482,N_13000,N_13145);
nand U13483 (N_13483,N_13156,N_13010);
xnor U13484 (N_13484,N_13114,N_13146);
nor U13485 (N_13485,N_13043,N_13211);
nor U13486 (N_13486,N_13011,N_13132);
nor U13487 (N_13487,N_13113,N_13076);
nand U13488 (N_13488,N_13193,N_13033);
nand U13489 (N_13489,N_13082,N_13024);
nand U13490 (N_13490,N_13008,N_13174);
and U13491 (N_13491,N_13166,N_13164);
nand U13492 (N_13492,N_13231,N_13011);
or U13493 (N_13493,N_13029,N_13073);
nor U13494 (N_13494,N_13081,N_13083);
and U13495 (N_13495,N_13221,N_13234);
nand U13496 (N_13496,N_13053,N_13064);
and U13497 (N_13497,N_13129,N_13197);
nand U13498 (N_13498,N_13218,N_13000);
and U13499 (N_13499,N_13179,N_13234);
or U13500 (N_13500,N_13397,N_13290);
and U13501 (N_13501,N_13264,N_13497);
nor U13502 (N_13502,N_13322,N_13467);
or U13503 (N_13503,N_13328,N_13426);
xnor U13504 (N_13504,N_13259,N_13289);
xnor U13505 (N_13505,N_13427,N_13317);
and U13506 (N_13506,N_13443,N_13472);
nor U13507 (N_13507,N_13311,N_13492);
nand U13508 (N_13508,N_13498,N_13447);
nor U13509 (N_13509,N_13457,N_13367);
and U13510 (N_13510,N_13361,N_13280);
or U13511 (N_13511,N_13465,N_13488);
and U13512 (N_13512,N_13484,N_13310);
and U13513 (N_13513,N_13454,N_13373);
and U13514 (N_13514,N_13262,N_13325);
or U13515 (N_13515,N_13345,N_13282);
nor U13516 (N_13516,N_13384,N_13480);
and U13517 (N_13517,N_13323,N_13257);
and U13518 (N_13518,N_13283,N_13483);
or U13519 (N_13519,N_13318,N_13471);
nand U13520 (N_13520,N_13390,N_13366);
or U13521 (N_13521,N_13255,N_13309);
nand U13522 (N_13522,N_13250,N_13331);
xnor U13523 (N_13523,N_13334,N_13370);
or U13524 (N_13524,N_13391,N_13319);
or U13525 (N_13525,N_13461,N_13332);
nor U13526 (N_13526,N_13269,N_13336);
and U13527 (N_13527,N_13495,N_13327);
and U13528 (N_13528,N_13413,N_13288);
nor U13529 (N_13529,N_13307,N_13409);
nand U13530 (N_13530,N_13416,N_13481);
nand U13531 (N_13531,N_13450,N_13470);
xor U13532 (N_13532,N_13347,N_13275);
xnor U13533 (N_13533,N_13440,N_13439);
nand U13534 (N_13534,N_13417,N_13482);
and U13535 (N_13535,N_13385,N_13441);
or U13536 (N_13536,N_13435,N_13422);
or U13537 (N_13537,N_13379,N_13365);
and U13538 (N_13538,N_13496,N_13256);
and U13539 (N_13539,N_13281,N_13329);
xnor U13540 (N_13540,N_13460,N_13359);
nor U13541 (N_13541,N_13434,N_13350);
and U13542 (N_13542,N_13466,N_13306);
or U13543 (N_13543,N_13272,N_13414);
xor U13544 (N_13544,N_13375,N_13316);
nor U13545 (N_13545,N_13287,N_13491);
nand U13546 (N_13546,N_13418,N_13456);
and U13547 (N_13547,N_13448,N_13320);
xor U13548 (N_13548,N_13267,N_13485);
and U13549 (N_13549,N_13442,N_13438);
or U13550 (N_13550,N_13342,N_13295);
nand U13551 (N_13551,N_13458,N_13389);
nand U13552 (N_13552,N_13446,N_13380);
and U13553 (N_13553,N_13343,N_13278);
or U13554 (N_13554,N_13252,N_13392);
nand U13555 (N_13555,N_13285,N_13261);
xnor U13556 (N_13556,N_13321,N_13398);
or U13557 (N_13557,N_13253,N_13411);
nand U13558 (N_13558,N_13301,N_13377);
nand U13559 (N_13559,N_13308,N_13358);
nor U13560 (N_13560,N_13400,N_13314);
or U13561 (N_13561,N_13304,N_13363);
and U13562 (N_13562,N_13421,N_13284);
nand U13563 (N_13563,N_13432,N_13337);
nand U13564 (N_13564,N_13431,N_13452);
or U13565 (N_13565,N_13300,N_13338);
or U13566 (N_13566,N_13277,N_13473);
nor U13567 (N_13567,N_13401,N_13464);
and U13568 (N_13568,N_13490,N_13424);
nand U13569 (N_13569,N_13399,N_13364);
xor U13570 (N_13570,N_13462,N_13403);
or U13571 (N_13571,N_13425,N_13368);
xor U13572 (N_13572,N_13305,N_13296);
xnor U13573 (N_13573,N_13386,N_13410);
nor U13574 (N_13574,N_13339,N_13265);
and U13575 (N_13575,N_13333,N_13459);
xor U13576 (N_13576,N_13362,N_13293);
nor U13577 (N_13577,N_13335,N_13451);
xnor U13578 (N_13578,N_13372,N_13455);
nor U13579 (N_13579,N_13344,N_13312);
or U13580 (N_13580,N_13346,N_13486);
xnor U13581 (N_13581,N_13388,N_13408);
nand U13582 (N_13582,N_13376,N_13374);
and U13583 (N_13583,N_13349,N_13326);
or U13584 (N_13584,N_13393,N_13378);
nand U13585 (N_13585,N_13297,N_13294);
nor U13586 (N_13586,N_13268,N_13348);
nand U13587 (N_13587,N_13251,N_13475);
xnor U13588 (N_13588,N_13354,N_13499);
and U13589 (N_13589,N_13436,N_13313);
nand U13590 (N_13590,N_13254,N_13406);
xnor U13591 (N_13591,N_13260,N_13355);
xor U13592 (N_13592,N_13276,N_13286);
or U13593 (N_13593,N_13382,N_13415);
and U13594 (N_13594,N_13453,N_13352);
and U13595 (N_13595,N_13468,N_13412);
or U13596 (N_13596,N_13353,N_13477);
nor U13597 (N_13597,N_13429,N_13394);
xnor U13598 (N_13598,N_13351,N_13299);
and U13599 (N_13599,N_13356,N_13387);
xnor U13600 (N_13600,N_13493,N_13273);
nand U13601 (N_13601,N_13271,N_13487);
nor U13602 (N_13602,N_13430,N_13423);
or U13603 (N_13603,N_13478,N_13371);
or U13604 (N_13604,N_13266,N_13469);
nand U13605 (N_13605,N_13476,N_13395);
nor U13606 (N_13606,N_13405,N_13489);
or U13607 (N_13607,N_13463,N_13433);
and U13608 (N_13608,N_13291,N_13292);
nor U13609 (N_13609,N_13428,N_13396);
xnor U13610 (N_13610,N_13258,N_13340);
xor U13611 (N_13611,N_13279,N_13445);
and U13612 (N_13612,N_13324,N_13444);
nand U13613 (N_13613,N_13302,N_13369);
nand U13614 (N_13614,N_13420,N_13270);
nand U13615 (N_13615,N_13404,N_13298);
xor U13616 (N_13616,N_13315,N_13330);
nor U13617 (N_13617,N_13494,N_13479);
xnor U13618 (N_13618,N_13341,N_13419);
nor U13619 (N_13619,N_13383,N_13274);
xnor U13620 (N_13620,N_13360,N_13449);
and U13621 (N_13621,N_13407,N_13263);
xor U13622 (N_13622,N_13402,N_13381);
xnor U13623 (N_13623,N_13437,N_13357);
nand U13624 (N_13624,N_13474,N_13303);
and U13625 (N_13625,N_13253,N_13388);
and U13626 (N_13626,N_13496,N_13345);
nand U13627 (N_13627,N_13274,N_13356);
xor U13628 (N_13628,N_13383,N_13345);
and U13629 (N_13629,N_13412,N_13254);
nand U13630 (N_13630,N_13417,N_13308);
and U13631 (N_13631,N_13439,N_13484);
nand U13632 (N_13632,N_13291,N_13410);
nor U13633 (N_13633,N_13471,N_13365);
xnor U13634 (N_13634,N_13352,N_13327);
or U13635 (N_13635,N_13340,N_13352);
xnor U13636 (N_13636,N_13286,N_13466);
nand U13637 (N_13637,N_13467,N_13319);
nor U13638 (N_13638,N_13452,N_13370);
or U13639 (N_13639,N_13343,N_13308);
nor U13640 (N_13640,N_13490,N_13277);
and U13641 (N_13641,N_13298,N_13309);
nand U13642 (N_13642,N_13303,N_13351);
xnor U13643 (N_13643,N_13330,N_13404);
nand U13644 (N_13644,N_13455,N_13267);
nor U13645 (N_13645,N_13275,N_13446);
nor U13646 (N_13646,N_13436,N_13379);
nand U13647 (N_13647,N_13296,N_13307);
nand U13648 (N_13648,N_13368,N_13415);
nand U13649 (N_13649,N_13404,N_13289);
nand U13650 (N_13650,N_13491,N_13387);
xor U13651 (N_13651,N_13327,N_13464);
nor U13652 (N_13652,N_13289,N_13333);
xor U13653 (N_13653,N_13349,N_13396);
and U13654 (N_13654,N_13377,N_13417);
xnor U13655 (N_13655,N_13479,N_13256);
xnor U13656 (N_13656,N_13262,N_13419);
nor U13657 (N_13657,N_13280,N_13370);
nor U13658 (N_13658,N_13343,N_13459);
and U13659 (N_13659,N_13367,N_13313);
xor U13660 (N_13660,N_13270,N_13396);
or U13661 (N_13661,N_13368,N_13359);
and U13662 (N_13662,N_13459,N_13370);
nand U13663 (N_13663,N_13401,N_13318);
and U13664 (N_13664,N_13322,N_13336);
and U13665 (N_13665,N_13310,N_13457);
nor U13666 (N_13666,N_13438,N_13382);
and U13667 (N_13667,N_13336,N_13335);
and U13668 (N_13668,N_13319,N_13396);
and U13669 (N_13669,N_13423,N_13458);
and U13670 (N_13670,N_13499,N_13430);
nand U13671 (N_13671,N_13325,N_13334);
nor U13672 (N_13672,N_13445,N_13365);
or U13673 (N_13673,N_13283,N_13346);
xor U13674 (N_13674,N_13441,N_13380);
nand U13675 (N_13675,N_13366,N_13276);
nor U13676 (N_13676,N_13494,N_13302);
nand U13677 (N_13677,N_13362,N_13320);
and U13678 (N_13678,N_13388,N_13437);
nor U13679 (N_13679,N_13454,N_13387);
nand U13680 (N_13680,N_13434,N_13295);
and U13681 (N_13681,N_13443,N_13331);
or U13682 (N_13682,N_13460,N_13382);
nor U13683 (N_13683,N_13257,N_13393);
and U13684 (N_13684,N_13314,N_13405);
and U13685 (N_13685,N_13466,N_13427);
or U13686 (N_13686,N_13379,N_13396);
or U13687 (N_13687,N_13499,N_13331);
and U13688 (N_13688,N_13418,N_13353);
xnor U13689 (N_13689,N_13375,N_13360);
nor U13690 (N_13690,N_13400,N_13455);
and U13691 (N_13691,N_13388,N_13382);
or U13692 (N_13692,N_13498,N_13372);
nor U13693 (N_13693,N_13295,N_13343);
xnor U13694 (N_13694,N_13468,N_13328);
and U13695 (N_13695,N_13390,N_13270);
or U13696 (N_13696,N_13412,N_13341);
or U13697 (N_13697,N_13335,N_13482);
nor U13698 (N_13698,N_13291,N_13386);
nor U13699 (N_13699,N_13420,N_13259);
or U13700 (N_13700,N_13484,N_13377);
xnor U13701 (N_13701,N_13318,N_13388);
nand U13702 (N_13702,N_13343,N_13495);
xnor U13703 (N_13703,N_13448,N_13309);
and U13704 (N_13704,N_13291,N_13354);
or U13705 (N_13705,N_13449,N_13250);
nor U13706 (N_13706,N_13451,N_13433);
nand U13707 (N_13707,N_13340,N_13480);
nor U13708 (N_13708,N_13329,N_13423);
xor U13709 (N_13709,N_13358,N_13419);
nand U13710 (N_13710,N_13354,N_13426);
or U13711 (N_13711,N_13302,N_13487);
nor U13712 (N_13712,N_13370,N_13400);
or U13713 (N_13713,N_13251,N_13443);
nor U13714 (N_13714,N_13374,N_13290);
and U13715 (N_13715,N_13272,N_13327);
nor U13716 (N_13716,N_13486,N_13255);
or U13717 (N_13717,N_13423,N_13366);
nor U13718 (N_13718,N_13342,N_13290);
or U13719 (N_13719,N_13291,N_13435);
nor U13720 (N_13720,N_13265,N_13419);
and U13721 (N_13721,N_13397,N_13473);
nor U13722 (N_13722,N_13422,N_13418);
and U13723 (N_13723,N_13265,N_13253);
nand U13724 (N_13724,N_13448,N_13357);
nor U13725 (N_13725,N_13277,N_13442);
or U13726 (N_13726,N_13344,N_13369);
or U13727 (N_13727,N_13329,N_13417);
nand U13728 (N_13728,N_13327,N_13433);
nor U13729 (N_13729,N_13388,N_13480);
and U13730 (N_13730,N_13429,N_13493);
nand U13731 (N_13731,N_13499,N_13439);
and U13732 (N_13732,N_13347,N_13354);
nand U13733 (N_13733,N_13479,N_13410);
nand U13734 (N_13734,N_13385,N_13293);
xor U13735 (N_13735,N_13464,N_13324);
nand U13736 (N_13736,N_13323,N_13288);
nor U13737 (N_13737,N_13262,N_13335);
nor U13738 (N_13738,N_13487,N_13353);
nand U13739 (N_13739,N_13459,N_13253);
nor U13740 (N_13740,N_13339,N_13463);
and U13741 (N_13741,N_13418,N_13457);
and U13742 (N_13742,N_13283,N_13417);
xnor U13743 (N_13743,N_13276,N_13359);
or U13744 (N_13744,N_13253,N_13311);
and U13745 (N_13745,N_13290,N_13438);
nor U13746 (N_13746,N_13432,N_13382);
nor U13747 (N_13747,N_13384,N_13294);
and U13748 (N_13748,N_13336,N_13384);
or U13749 (N_13749,N_13414,N_13321);
nand U13750 (N_13750,N_13699,N_13500);
nor U13751 (N_13751,N_13705,N_13569);
xor U13752 (N_13752,N_13546,N_13619);
or U13753 (N_13753,N_13670,N_13642);
nor U13754 (N_13754,N_13706,N_13543);
nand U13755 (N_13755,N_13680,N_13544);
and U13756 (N_13756,N_13721,N_13559);
and U13757 (N_13757,N_13741,N_13735);
or U13758 (N_13758,N_13577,N_13505);
nand U13759 (N_13759,N_13593,N_13573);
and U13760 (N_13760,N_13687,N_13726);
and U13761 (N_13761,N_13531,N_13635);
nand U13762 (N_13762,N_13677,N_13638);
nand U13763 (N_13763,N_13691,N_13737);
or U13764 (N_13764,N_13742,N_13600);
nand U13765 (N_13765,N_13719,N_13659);
nand U13766 (N_13766,N_13740,N_13612);
nor U13767 (N_13767,N_13566,N_13506);
xor U13768 (N_13768,N_13567,N_13665);
and U13769 (N_13769,N_13633,N_13604);
nand U13770 (N_13770,N_13613,N_13651);
nand U13771 (N_13771,N_13652,N_13524);
nand U13772 (N_13772,N_13607,N_13729);
or U13773 (N_13773,N_13647,N_13654);
or U13774 (N_13774,N_13663,N_13707);
nand U13775 (N_13775,N_13636,N_13644);
nor U13776 (N_13776,N_13526,N_13556);
nor U13777 (N_13777,N_13689,N_13530);
or U13778 (N_13778,N_13621,N_13716);
or U13779 (N_13779,N_13669,N_13591);
nand U13780 (N_13780,N_13645,N_13601);
nor U13781 (N_13781,N_13535,N_13534);
nand U13782 (N_13782,N_13503,N_13587);
nand U13783 (N_13783,N_13743,N_13712);
nand U13784 (N_13784,N_13568,N_13734);
nand U13785 (N_13785,N_13649,N_13510);
and U13786 (N_13786,N_13722,N_13529);
nand U13787 (N_13787,N_13521,N_13615);
nand U13788 (N_13788,N_13558,N_13702);
nor U13789 (N_13789,N_13727,N_13516);
or U13790 (N_13790,N_13545,N_13572);
and U13791 (N_13791,N_13552,N_13576);
nor U13792 (N_13792,N_13748,N_13578);
nor U13793 (N_13793,N_13720,N_13536);
nor U13794 (N_13794,N_13730,N_13731);
nand U13795 (N_13795,N_13682,N_13562);
nand U13796 (N_13796,N_13634,N_13527);
nor U13797 (N_13797,N_13513,N_13581);
nand U13798 (N_13798,N_13664,N_13629);
or U13799 (N_13799,N_13584,N_13708);
nor U13800 (N_13800,N_13704,N_13686);
xor U13801 (N_13801,N_13523,N_13632);
xor U13802 (N_13802,N_13700,N_13668);
and U13803 (N_13803,N_13690,N_13598);
or U13804 (N_13804,N_13745,N_13518);
nand U13805 (N_13805,N_13501,N_13672);
nor U13806 (N_13806,N_13724,N_13557);
or U13807 (N_13807,N_13564,N_13693);
nand U13808 (N_13808,N_13588,N_13627);
nor U13809 (N_13809,N_13599,N_13650);
nand U13810 (N_13810,N_13733,N_13504);
xor U13811 (N_13811,N_13739,N_13596);
nor U13812 (N_13812,N_13695,N_13628);
xnor U13813 (N_13813,N_13514,N_13565);
nand U13814 (N_13814,N_13641,N_13608);
xor U13815 (N_13815,N_13508,N_13595);
and U13816 (N_13816,N_13614,N_13698);
nor U13817 (N_13817,N_13571,N_13616);
nor U13818 (N_13818,N_13512,N_13656);
nand U13819 (N_13819,N_13648,N_13592);
xor U13820 (N_13820,N_13609,N_13711);
nor U13821 (N_13821,N_13519,N_13671);
nor U13822 (N_13822,N_13550,N_13703);
nor U13823 (N_13823,N_13646,N_13688);
and U13824 (N_13824,N_13582,N_13723);
nor U13825 (N_13825,N_13639,N_13709);
and U13826 (N_13826,N_13620,N_13554);
or U13827 (N_13827,N_13553,N_13736);
xnor U13828 (N_13828,N_13549,N_13579);
xnor U13829 (N_13829,N_13622,N_13625);
or U13830 (N_13830,N_13580,N_13610);
and U13831 (N_13831,N_13681,N_13533);
nor U13832 (N_13832,N_13570,N_13710);
nor U13833 (N_13833,N_13657,N_13575);
and U13834 (N_13834,N_13714,N_13747);
nand U13835 (N_13835,N_13744,N_13597);
or U13836 (N_13836,N_13548,N_13630);
nand U13837 (N_13837,N_13653,N_13713);
nor U13838 (N_13838,N_13583,N_13603);
xnor U13839 (N_13839,N_13611,N_13738);
xnor U13840 (N_13840,N_13509,N_13697);
or U13841 (N_13841,N_13602,N_13667);
xnor U13842 (N_13842,N_13502,N_13666);
or U13843 (N_13843,N_13637,N_13574);
or U13844 (N_13844,N_13585,N_13746);
or U13845 (N_13845,N_13675,N_13547);
nor U13846 (N_13846,N_13684,N_13617);
xnor U13847 (N_13847,N_13662,N_13749);
nand U13848 (N_13848,N_13658,N_13643);
xor U13849 (N_13849,N_13555,N_13624);
nor U13850 (N_13850,N_13542,N_13674);
xnor U13851 (N_13851,N_13605,N_13732);
nand U13852 (N_13852,N_13586,N_13678);
and U13853 (N_13853,N_13685,N_13589);
or U13854 (N_13854,N_13520,N_13660);
xor U13855 (N_13855,N_13692,N_13717);
xnor U13856 (N_13856,N_13528,N_13551);
and U13857 (N_13857,N_13694,N_13718);
nor U13858 (N_13858,N_13661,N_13563);
xnor U13859 (N_13859,N_13525,N_13631);
nor U13860 (N_13860,N_13541,N_13515);
nor U13861 (N_13861,N_13701,N_13623);
xor U13862 (N_13862,N_13560,N_13626);
nand U13863 (N_13863,N_13673,N_13683);
nor U13864 (N_13864,N_13511,N_13696);
nor U13865 (N_13865,N_13561,N_13594);
nor U13866 (N_13866,N_13640,N_13676);
xor U13867 (N_13867,N_13715,N_13618);
or U13868 (N_13868,N_13538,N_13522);
nand U13869 (N_13869,N_13539,N_13540);
nand U13870 (N_13870,N_13537,N_13606);
or U13871 (N_13871,N_13517,N_13679);
nand U13872 (N_13872,N_13590,N_13728);
or U13873 (N_13873,N_13532,N_13725);
nand U13874 (N_13874,N_13655,N_13507);
nor U13875 (N_13875,N_13725,N_13740);
xor U13876 (N_13876,N_13603,N_13501);
or U13877 (N_13877,N_13659,N_13575);
nor U13878 (N_13878,N_13645,N_13581);
nand U13879 (N_13879,N_13581,N_13598);
xnor U13880 (N_13880,N_13681,N_13593);
xor U13881 (N_13881,N_13614,N_13635);
or U13882 (N_13882,N_13707,N_13690);
and U13883 (N_13883,N_13746,N_13620);
or U13884 (N_13884,N_13721,N_13556);
nand U13885 (N_13885,N_13672,N_13697);
or U13886 (N_13886,N_13587,N_13601);
xor U13887 (N_13887,N_13680,N_13535);
xor U13888 (N_13888,N_13599,N_13601);
nand U13889 (N_13889,N_13581,N_13728);
nor U13890 (N_13890,N_13701,N_13539);
xor U13891 (N_13891,N_13621,N_13508);
nand U13892 (N_13892,N_13681,N_13547);
or U13893 (N_13893,N_13631,N_13725);
nand U13894 (N_13894,N_13625,N_13662);
xnor U13895 (N_13895,N_13587,N_13708);
nand U13896 (N_13896,N_13683,N_13573);
xnor U13897 (N_13897,N_13736,N_13665);
xor U13898 (N_13898,N_13746,N_13697);
xor U13899 (N_13899,N_13630,N_13578);
xor U13900 (N_13900,N_13511,N_13714);
xor U13901 (N_13901,N_13554,N_13577);
nor U13902 (N_13902,N_13646,N_13587);
or U13903 (N_13903,N_13719,N_13589);
and U13904 (N_13904,N_13550,N_13628);
nor U13905 (N_13905,N_13647,N_13512);
or U13906 (N_13906,N_13607,N_13546);
nor U13907 (N_13907,N_13527,N_13617);
xnor U13908 (N_13908,N_13632,N_13587);
and U13909 (N_13909,N_13625,N_13583);
or U13910 (N_13910,N_13529,N_13651);
nand U13911 (N_13911,N_13715,N_13673);
and U13912 (N_13912,N_13525,N_13732);
xor U13913 (N_13913,N_13622,N_13623);
and U13914 (N_13914,N_13553,N_13674);
or U13915 (N_13915,N_13605,N_13621);
and U13916 (N_13916,N_13511,N_13629);
nor U13917 (N_13917,N_13647,N_13673);
xor U13918 (N_13918,N_13745,N_13692);
or U13919 (N_13919,N_13634,N_13680);
nand U13920 (N_13920,N_13617,N_13669);
or U13921 (N_13921,N_13586,N_13563);
or U13922 (N_13922,N_13744,N_13506);
nor U13923 (N_13923,N_13629,N_13678);
nand U13924 (N_13924,N_13503,N_13606);
or U13925 (N_13925,N_13709,N_13601);
or U13926 (N_13926,N_13664,N_13730);
nor U13927 (N_13927,N_13572,N_13634);
nand U13928 (N_13928,N_13735,N_13737);
or U13929 (N_13929,N_13620,N_13640);
xnor U13930 (N_13930,N_13681,N_13662);
xor U13931 (N_13931,N_13662,N_13676);
and U13932 (N_13932,N_13575,N_13623);
or U13933 (N_13933,N_13643,N_13606);
nand U13934 (N_13934,N_13729,N_13651);
and U13935 (N_13935,N_13661,N_13577);
or U13936 (N_13936,N_13507,N_13549);
or U13937 (N_13937,N_13530,N_13625);
and U13938 (N_13938,N_13609,N_13611);
nor U13939 (N_13939,N_13605,N_13692);
or U13940 (N_13940,N_13583,N_13637);
or U13941 (N_13941,N_13583,N_13719);
or U13942 (N_13942,N_13648,N_13657);
xor U13943 (N_13943,N_13726,N_13667);
nor U13944 (N_13944,N_13676,N_13547);
nor U13945 (N_13945,N_13686,N_13579);
xnor U13946 (N_13946,N_13682,N_13586);
or U13947 (N_13947,N_13663,N_13717);
and U13948 (N_13948,N_13531,N_13615);
and U13949 (N_13949,N_13573,N_13608);
nand U13950 (N_13950,N_13543,N_13682);
nor U13951 (N_13951,N_13662,N_13666);
and U13952 (N_13952,N_13565,N_13748);
and U13953 (N_13953,N_13635,N_13507);
nand U13954 (N_13954,N_13600,N_13521);
and U13955 (N_13955,N_13672,N_13650);
and U13956 (N_13956,N_13500,N_13737);
nand U13957 (N_13957,N_13606,N_13745);
and U13958 (N_13958,N_13707,N_13601);
and U13959 (N_13959,N_13658,N_13654);
or U13960 (N_13960,N_13562,N_13538);
nand U13961 (N_13961,N_13677,N_13718);
nor U13962 (N_13962,N_13560,N_13741);
nor U13963 (N_13963,N_13672,N_13647);
xor U13964 (N_13964,N_13700,N_13636);
or U13965 (N_13965,N_13664,N_13718);
and U13966 (N_13966,N_13517,N_13704);
xnor U13967 (N_13967,N_13510,N_13677);
or U13968 (N_13968,N_13687,N_13597);
nor U13969 (N_13969,N_13513,N_13575);
nor U13970 (N_13970,N_13518,N_13746);
nand U13971 (N_13971,N_13542,N_13594);
nor U13972 (N_13972,N_13728,N_13645);
nor U13973 (N_13973,N_13654,N_13638);
nand U13974 (N_13974,N_13648,N_13582);
nor U13975 (N_13975,N_13725,N_13666);
xnor U13976 (N_13976,N_13722,N_13603);
or U13977 (N_13977,N_13610,N_13631);
and U13978 (N_13978,N_13541,N_13545);
and U13979 (N_13979,N_13566,N_13624);
nor U13980 (N_13980,N_13719,N_13715);
and U13981 (N_13981,N_13633,N_13623);
nand U13982 (N_13982,N_13632,N_13571);
or U13983 (N_13983,N_13550,N_13720);
nor U13984 (N_13984,N_13736,N_13526);
and U13985 (N_13985,N_13649,N_13739);
nand U13986 (N_13986,N_13570,N_13729);
nor U13987 (N_13987,N_13627,N_13655);
or U13988 (N_13988,N_13681,N_13609);
xor U13989 (N_13989,N_13527,N_13623);
and U13990 (N_13990,N_13517,N_13701);
or U13991 (N_13991,N_13603,N_13518);
or U13992 (N_13992,N_13682,N_13733);
nor U13993 (N_13993,N_13706,N_13712);
and U13994 (N_13994,N_13507,N_13739);
nand U13995 (N_13995,N_13539,N_13542);
and U13996 (N_13996,N_13642,N_13722);
nor U13997 (N_13997,N_13746,N_13735);
and U13998 (N_13998,N_13516,N_13613);
or U13999 (N_13999,N_13711,N_13589);
and U14000 (N_14000,N_13969,N_13881);
or U14001 (N_14001,N_13766,N_13992);
and U14002 (N_14002,N_13800,N_13948);
or U14003 (N_14003,N_13941,N_13939);
nor U14004 (N_14004,N_13798,N_13998);
or U14005 (N_14005,N_13809,N_13901);
nor U14006 (N_14006,N_13808,N_13756);
and U14007 (N_14007,N_13973,N_13949);
xnor U14008 (N_14008,N_13841,N_13818);
nand U14009 (N_14009,N_13765,N_13916);
nand U14010 (N_14010,N_13976,N_13794);
nand U14011 (N_14011,N_13986,N_13855);
nor U14012 (N_14012,N_13968,N_13950);
nor U14013 (N_14013,N_13990,N_13930);
nor U14014 (N_14014,N_13918,N_13959);
nor U14015 (N_14015,N_13757,N_13753);
or U14016 (N_14016,N_13825,N_13868);
xnor U14017 (N_14017,N_13829,N_13801);
nor U14018 (N_14018,N_13910,N_13854);
xnor U14019 (N_14019,N_13819,N_13997);
or U14020 (N_14020,N_13919,N_13859);
nand U14021 (N_14021,N_13844,N_13759);
xor U14022 (N_14022,N_13848,N_13871);
nand U14023 (N_14023,N_13850,N_13775);
xnor U14024 (N_14024,N_13758,N_13987);
and U14025 (N_14025,N_13983,N_13900);
and U14026 (N_14026,N_13928,N_13851);
or U14027 (N_14027,N_13909,N_13863);
nor U14028 (N_14028,N_13838,N_13956);
nand U14029 (N_14029,N_13932,N_13920);
and U14030 (N_14030,N_13776,N_13913);
and U14031 (N_14031,N_13926,N_13942);
nor U14032 (N_14032,N_13872,N_13862);
and U14033 (N_14033,N_13857,N_13887);
xor U14034 (N_14034,N_13787,N_13791);
xor U14035 (N_14035,N_13889,N_13937);
nand U14036 (N_14036,N_13828,N_13830);
nand U14037 (N_14037,N_13917,N_13891);
or U14038 (N_14038,N_13799,N_13897);
or U14039 (N_14039,N_13784,N_13898);
or U14040 (N_14040,N_13955,N_13849);
nand U14041 (N_14041,N_13905,N_13778);
nor U14042 (N_14042,N_13780,N_13944);
xor U14043 (N_14043,N_13996,N_13972);
nand U14044 (N_14044,N_13852,N_13988);
nand U14045 (N_14045,N_13879,N_13790);
and U14046 (N_14046,N_13878,N_13893);
xnor U14047 (N_14047,N_13755,N_13962);
or U14048 (N_14048,N_13783,N_13824);
or U14049 (N_14049,N_13903,N_13772);
or U14050 (N_14050,N_13875,N_13888);
and U14051 (N_14051,N_13974,N_13895);
xnor U14052 (N_14052,N_13779,N_13938);
nor U14053 (N_14053,N_13923,N_13985);
xor U14054 (N_14054,N_13995,N_13979);
and U14055 (N_14055,N_13813,N_13989);
nand U14056 (N_14056,N_13795,N_13853);
xor U14057 (N_14057,N_13977,N_13951);
or U14058 (N_14058,N_13991,N_13876);
xnor U14059 (N_14059,N_13936,N_13880);
xnor U14060 (N_14060,N_13820,N_13822);
or U14061 (N_14061,N_13884,N_13954);
or U14062 (N_14062,N_13856,N_13922);
xnor U14063 (N_14063,N_13833,N_13858);
xnor U14064 (N_14064,N_13817,N_13894);
and U14065 (N_14065,N_13981,N_13821);
or U14066 (N_14066,N_13842,N_13786);
nand U14067 (N_14067,N_13877,N_13964);
nor U14068 (N_14068,N_13843,N_13940);
nand U14069 (N_14069,N_13911,N_13797);
nand U14070 (N_14070,N_13957,N_13999);
and U14071 (N_14071,N_13835,N_13978);
nand U14072 (N_14072,N_13761,N_13965);
nand U14073 (N_14073,N_13945,N_13793);
or U14074 (N_14074,N_13792,N_13924);
xor U14075 (N_14075,N_13807,N_13946);
nor U14076 (N_14076,N_13796,N_13806);
or U14077 (N_14077,N_13914,N_13760);
nand U14078 (N_14078,N_13904,N_13993);
nor U14079 (N_14079,N_13768,N_13823);
or U14080 (N_14080,N_13840,N_13802);
and U14081 (N_14081,N_13931,N_13812);
nor U14082 (N_14082,N_13788,N_13831);
xnor U14083 (N_14083,N_13980,N_13912);
nor U14084 (N_14084,N_13927,N_13921);
xor U14085 (N_14085,N_13885,N_13805);
nand U14086 (N_14086,N_13754,N_13929);
nor U14087 (N_14087,N_13750,N_13867);
xor U14088 (N_14088,N_13899,N_13984);
nor U14089 (N_14089,N_13845,N_13751);
or U14090 (N_14090,N_13896,N_13781);
xnor U14091 (N_14091,N_13767,N_13803);
xnor U14092 (N_14092,N_13902,N_13870);
xnor U14093 (N_14093,N_13960,N_13907);
or U14094 (N_14094,N_13816,N_13811);
or U14095 (N_14095,N_13763,N_13752);
nor U14096 (N_14096,N_13883,N_13782);
and U14097 (N_14097,N_13873,N_13785);
nand U14098 (N_14098,N_13769,N_13860);
xor U14099 (N_14099,N_13771,N_13804);
nor U14100 (N_14100,N_13963,N_13961);
nor U14101 (N_14101,N_13815,N_13846);
and U14102 (N_14102,N_13847,N_13839);
xnor U14103 (N_14103,N_13886,N_13975);
or U14104 (N_14104,N_13827,N_13836);
or U14105 (N_14105,N_13762,N_13934);
and U14106 (N_14106,N_13952,N_13777);
nor U14107 (N_14107,N_13869,N_13943);
and U14108 (N_14108,N_13864,N_13933);
nand U14109 (N_14109,N_13810,N_13789);
or U14110 (N_14110,N_13832,N_13826);
or U14111 (N_14111,N_13770,N_13892);
nand U14112 (N_14112,N_13890,N_13970);
and U14113 (N_14113,N_13774,N_13882);
and U14114 (N_14114,N_13967,N_13865);
nand U14115 (N_14115,N_13994,N_13925);
nand U14116 (N_14116,N_13837,N_13915);
nand U14117 (N_14117,N_13971,N_13908);
and U14118 (N_14118,N_13874,N_13814);
nor U14119 (N_14119,N_13866,N_13982);
xor U14120 (N_14120,N_13773,N_13764);
nand U14121 (N_14121,N_13834,N_13906);
and U14122 (N_14122,N_13935,N_13861);
and U14123 (N_14123,N_13947,N_13958);
or U14124 (N_14124,N_13966,N_13953);
nand U14125 (N_14125,N_13896,N_13834);
and U14126 (N_14126,N_13899,N_13782);
or U14127 (N_14127,N_13763,N_13871);
nor U14128 (N_14128,N_13907,N_13890);
xnor U14129 (N_14129,N_13968,N_13876);
or U14130 (N_14130,N_13791,N_13918);
xor U14131 (N_14131,N_13824,N_13890);
nand U14132 (N_14132,N_13812,N_13851);
and U14133 (N_14133,N_13788,N_13913);
or U14134 (N_14134,N_13755,N_13816);
or U14135 (N_14135,N_13846,N_13847);
or U14136 (N_14136,N_13984,N_13869);
xnor U14137 (N_14137,N_13781,N_13892);
nor U14138 (N_14138,N_13887,N_13828);
and U14139 (N_14139,N_13793,N_13818);
nor U14140 (N_14140,N_13977,N_13982);
or U14141 (N_14141,N_13999,N_13852);
xnor U14142 (N_14142,N_13817,N_13879);
nor U14143 (N_14143,N_13817,N_13764);
xor U14144 (N_14144,N_13968,N_13787);
nor U14145 (N_14145,N_13964,N_13832);
and U14146 (N_14146,N_13865,N_13966);
nor U14147 (N_14147,N_13876,N_13937);
or U14148 (N_14148,N_13864,N_13898);
and U14149 (N_14149,N_13943,N_13989);
and U14150 (N_14150,N_13838,N_13848);
or U14151 (N_14151,N_13792,N_13833);
and U14152 (N_14152,N_13980,N_13924);
and U14153 (N_14153,N_13879,N_13815);
or U14154 (N_14154,N_13997,N_13798);
or U14155 (N_14155,N_13873,N_13797);
and U14156 (N_14156,N_13862,N_13965);
nand U14157 (N_14157,N_13924,N_13838);
and U14158 (N_14158,N_13906,N_13913);
nor U14159 (N_14159,N_13906,N_13895);
and U14160 (N_14160,N_13830,N_13936);
and U14161 (N_14161,N_13832,N_13887);
nor U14162 (N_14162,N_13860,N_13938);
nor U14163 (N_14163,N_13877,N_13896);
nand U14164 (N_14164,N_13784,N_13932);
xor U14165 (N_14165,N_13791,N_13806);
nor U14166 (N_14166,N_13867,N_13980);
xor U14167 (N_14167,N_13926,N_13923);
or U14168 (N_14168,N_13834,N_13868);
and U14169 (N_14169,N_13954,N_13910);
nor U14170 (N_14170,N_13770,N_13912);
or U14171 (N_14171,N_13837,N_13880);
nor U14172 (N_14172,N_13914,N_13902);
nand U14173 (N_14173,N_13776,N_13910);
or U14174 (N_14174,N_13918,N_13939);
xor U14175 (N_14175,N_13970,N_13987);
nand U14176 (N_14176,N_13833,N_13905);
xnor U14177 (N_14177,N_13778,N_13946);
nand U14178 (N_14178,N_13987,N_13866);
xnor U14179 (N_14179,N_13768,N_13977);
or U14180 (N_14180,N_13753,N_13934);
or U14181 (N_14181,N_13996,N_13753);
xor U14182 (N_14182,N_13937,N_13946);
nor U14183 (N_14183,N_13820,N_13864);
nand U14184 (N_14184,N_13943,N_13919);
nor U14185 (N_14185,N_13885,N_13763);
xor U14186 (N_14186,N_13854,N_13889);
nand U14187 (N_14187,N_13837,N_13779);
or U14188 (N_14188,N_13819,N_13767);
xnor U14189 (N_14189,N_13832,N_13820);
nor U14190 (N_14190,N_13963,N_13834);
nor U14191 (N_14191,N_13828,N_13794);
and U14192 (N_14192,N_13971,N_13973);
nor U14193 (N_14193,N_13752,N_13987);
or U14194 (N_14194,N_13966,N_13786);
nand U14195 (N_14195,N_13934,N_13861);
nor U14196 (N_14196,N_13983,N_13891);
and U14197 (N_14197,N_13941,N_13897);
or U14198 (N_14198,N_13872,N_13819);
and U14199 (N_14199,N_13933,N_13904);
nand U14200 (N_14200,N_13896,N_13978);
or U14201 (N_14201,N_13977,N_13928);
or U14202 (N_14202,N_13985,N_13951);
nor U14203 (N_14203,N_13808,N_13919);
xnor U14204 (N_14204,N_13828,N_13799);
or U14205 (N_14205,N_13940,N_13917);
xnor U14206 (N_14206,N_13998,N_13752);
or U14207 (N_14207,N_13984,N_13986);
xor U14208 (N_14208,N_13832,N_13778);
nor U14209 (N_14209,N_13915,N_13808);
xor U14210 (N_14210,N_13848,N_13962);
and U14211 (N_14211,N_13769,N_13838);
nor U14212 (N_14212,N_13827,N_13808);
xor U14213 (N_14213,N_13812,N_13950);
nand U14214 (N_14214,N_13775,N_13836);
nand U14215 (N_14215,N_13807,N_13941);
nor U14216 (N_14216,N_13920,N_13813);
nor U14217 (N_14217,N_13793,N_13890);
nand U14218 (N_14218,N_13759,N_13791);
xor U14219 (N_14219,N_13793,N_13905);
or U14220 (N_14220,N_13984,N_13828);
nand U14221 (N_14221,N_13906,N_13833);
nand U14222 (N_14222,N_13938,N_13880);
or U14223 (N_14223,N_13826,N_13970);
nand U14224 (N_14224,N_13970,N_13966);
nor U14225 (N_14225,N_13807,N_13873);
or U14226 (N_14226,N_13980,N_13892);
nand U14227 (N_14227,N_13887,N_13896);
or U14228 (N_14228,N_13808,N_13971);
and U14229 (N_14229,N_13984,N_13942);
and U14230 (N_14230,N_13855,N_13762);
xnor U14231 (N_14231,N_13970,N_13955);
nor U14232 (N_14232,N_13876,N_13816);
nor U14233 (N_14233,N_13783,N_13776);
xnor U14234 (N_14234,N_13843,N_13897);
and U14235 (N_14235,N_13931,N_13797);
nor U14236 (N_14236,N_13894,N_13840);
nor U14237 (N_14237,N_13869,N_13876);
or U14238 (N_14238,N_13866,N_13952);
nand U14239 (N_14239,N_13935,N_13936);
nor U14240 (N_14240,N_13810,N_13801);
and U14241 (N_14241,N_13894,N_13775);
or U14242 (N_14242,N_13933,N_13994);
and U14243 (N_14243,N_13926,N_13964);
and U14244 (N_14244,N_13862,N_13970);
or U14245 (N_14245,N_13796,N_13988);
or U14246 (N_14246,N_13788,N_13845);
nand U14247 (N_14247,N_13793,N_13995);
and U14248 (N_14248,N_13932,N_13830);
nor U14249 (N_14249,N_13808,N_13806);
and U14250 (N_14250,N_14051,N_14122);
nor U14251 (N_14251,N_14174,N_14195);
and U14252 (N_14252,N_14097,N_14237);
nand U14253 (N_14253,N_14190,N_14091);
or U14254 (N_14254,N_14032,N_14184);
nand U14255 (N_14255,N_14008,N_14206);
nor U14256 (N_14256,N_14223,N_14131);
nor U14257 (N_14257,N_14039,N_14110);
nor U14258 (N_14258,N_14069,N_14128);
or U14259 (N_14259,N_14020,N_14001);
nand U14260 (N_14260,N_14210,N_14155);
nand U14261 (N_14261,N_14086,N_14046);
nand U14262 (N_14262,N_14041,N_14166);
nand U14263 (N_14263,N_14243,N_14026);
xor U14264 (N_14264,N_14140,N_14170);
or U14265 (N_14265,N_14227,N_14240);
nor U14266 (N_14266,N_14102,N_14221);
xnor U14267 (N_14267,N_14191,N_14149);
xor U14268 (N_14268,N_14065,N_14027);
xnor U14269 (N_14269,N_14212,N_14014);
and U14270 (N_14270,N_14104,N_14031);
nor U14271 (N_14271,N_14093,N_14241);
xnor U14272 (N_14272,N_14007,N_14134);
and U14273 (N_14273,N_14179,N_14211);
nor U14274 (N_14274,N_14066,N_14245);
or U14275 (N_14275,N_14204,N_14129);
or U14276 (N_14276,N_14124,N_14025);
xor U14277 (N_14277,N_14100,N_14151);
xnor U14278 (N_14278,N_14022,N_14111);
and U14279 (N_14279,N_14006,N_14207);
and U14280 (N_14280,N_14139,N_14067);
nand U14281 (N_14281,N_14000,N_14150);
nor U14282 (N_14282,N_14197,N_14157);
and U14283 (N_14283,N_14083,N_14017);
or U14284 (N_14284,N_14165,N_14021);
xor U14285 (N_14285,N_14082,N_14012);
or U14286 (N_14286,N_14004,N_14037);
nor U14287 (N_14287,N_14118,N_14231);
and U14288 (N_14288,N_14219,N_14103);
and U14289 (N_14289,N_14060,N_14003);
nor U14290 (N_14290,N_14099,N_14224);
nor U14291 (N_14291,N_14028,N_14144);
or U14292 (N_14292,N_14145,N_14002);
nor U14293 (N_14293,N_14222,N_14096);
and U14294 (N_14294,N_14249,N_14218);
or U14295 (N_14295,N_14143,N_14246);
xnor U14296 (N_14296,N_14036,N_14234);
and U14297 (N_14297,N_14239,N_14013);
xor U14298 (N_14298,N_14119,N_14076);
or U14299 (N_14299,N_14203,N_14087);
xor U14300 (N_14300,N_14117,N_14085);
nor U14301 (N_14301,N_14167,N_14229);
nor U14302 (N_14302,N_14054,N_14044);
xnor U14303 (N_14303,N_14029,N_14169);
nor U14304 (N_14304,N_14200,N_14090);
nor U14305 (N_14305,N_14189,N_14214);
xnor U14306 (N_14306,N_14205,N_14141);
or U14307 (N_14307,N_14146,N_14057);
xnor U14308 (N_14308,N_14137,N_14005);
xnor U14309 (N_14309,N_14194,N_14136);
xor U14310 (N_14310,N_14156,N_14130);
or U14311 (N_14311,N_14064,N_14063);
or U14312 (N_14312,N_14115,N_14228);
nor U14313 (N_14313,N_14043,N_14225);
nor U14314 (N_14314,N_14162,N_14132);
or U14315 (N_14315,N_14192,N_14233);
xnor U14316 (N_14316,N_14138,N_14154);
xnor U14317 (N_14317,N_14078,N_14107);
or U14318 (N_14318,N_14176,N_14024);
or U14319 (N_14319,N_14161,N_14055);
or U14320 (N_14320,N_14070,N_14216);
or U14321 (N_14321,N_14153,N_14010);
xnor U14322 (N_14322,N_14125,N_14120);
nor U14323 (N_14323,N_14053,N_14018);
xor U14324 (N_14324,N_14244,N_14186);
nand U14325 (N_14325,N_14198,N_14177);
and U14326 (N_14326,N_14185,N_14199);
and U14327 (N_14327,N_14202,N_14073);
xor U14328 (N_14328,N_14109,N_14236);
nor U14329 (N_14329,N_14158,N_14220);
nor U14330 (N_14330,N_14188,N_14175);
and U14331 (N_14331,N_14193,N_14180);
xnor U14332 (N_14332,N_14232,N_14114);
nor U14333 (N_14333,N_14123,N_14133);
nor U14334 (N_14334,N_14088,N_14048);
nand U14335 (N_14335,N_14112,N_14226);
or U14336 (N_14336,N_14173,N_14011);
nor U14337 (N_14337,N_14023,N_14038);
and U14338 (N_14338,N_14019,N_14235);
nand U14339 (N_14339,N_14079,N_14035);
or U14340 (N_14340,N_14159,N_14095);
nand U14341 (N_14341,N_14181,N_14047);
and U14342 (N_14342,N_14075,N_14142);
nor U14343 (N_14343,N_14101,N_14217);
nand U14344 (N_14344,N_14016,N_14113);
nand U14345 (N_14345,N_14121,N_14196);
nor U14346 (N_14346,N_14030,N_14147);
and U14347 (N_14347,N_14209,N_14248);
xnor U14348 (N_14348,N_14061,N_14126);
or U14349 (N_14349,N_14108,N_14247);
nor U14350 (N_14350,N_14106,N_14152);
or U14351 (N_14351,N_14171,N_14084);
nand U14352 (N_14352,N_14094,N_14071);
xor U14353 (N_14353,N_14077,N_14116);
xnor U14354 (N_14354,N_14148,N_14033);
nand U14355 (N_14355,N_14050,N_14074);
and U14356 (N_14356,N_14052,N_14230);
xor U14357 (N_14357,N_14182,N_14049);
xor U14358 (N_14358,N_14009,N_14163);
nand U14359 (N_14359,N_14105,N_14034);
xnor U14360 (N_14360,N_14058,N_14164);
and U14361 (N_14361,N_14056,N_14135);
nor U14362 (N_14362,N_14238,N_14068);
or U14363 (N_14363,N_14187,N_14089);
xnor U14364 (N_14364,N_14183,N_14072);
nor U14365 (N_14365,N_14042,N_14201);
xor U14366 (N_14366,N_14098,N_14092);
or U14367 (N_14367,N_14040,N_14242);
nor U14368 (N_14368,N_14215,N_14172);
nand U14369 (N_14369,N_14081,N_14080);
nand U14370 (N_14370,N_14168,N_14045);
xor U14371 (N_14371,N_14178,N_14213);
nor U14372 (N_14372,N_14062,N_14208);
nand U14373 (N_14373,N_14015,N_14059);
or U14374 (N_14374,N_14160,N_14127);
nand U14375 (N_14375,N_14123,N_14037);
nor U14376 (N_14376,N_14171,N_14118);
xnor U14377 (N_14377,N_14125,N_14172);
nor U14378 (N_14378,N_14223,N_14127);
or U14379 (N_14379,N_14071,N_14230);
or U14380 (N_14380,N_14165,N_14036);
nor U14381 (N_14381,N_14124,N_14062);
or U14382 (N_14382,N_14215,N_14236);
and U14383 (N_14383,N_14072,N_14201);
nand U14384 (N_14384,N_14024,N_14156);
and U14385 (N_14385,N_14011,N_14086);
and U14386 (N_14386,N_14194,N_14247);
or U14387 (N_14387,N_14195,N_14179);
nand U14388 (N_14388,N_14059,N_14105);
and U14389 (N_14389,N_14146,N_14142);
nand U14390 (N_14390,N_14071,N_14127);
nor U14391 (N_14391,N_14243,N_14113);
xor U14392 (N_14392,N_14047,N_14225);
xor U14393 (N_14393,N_14182,N_14057);
or U14394 (N_14394,N_14080,N_14056);
xnor U14395 (N_14395,N_14221,N_14184);
or U14396 (N_14396,N_14218,N_14245);
and U14397 (N_14397,N_14084,N_14188);
xor U14398 (N_14398,N_14197,N_14122);
and U14399 (N_14399,N_14185,N_14203);
and U14400 (N_14400,N_14026,N_14212);
nor U14401 (N_14401,N_14031,N_14137);
or U14402 (N_14402,N_14199,N_14143);
xor U14403 (N_14403,N_14005,N_14033);
nand U14404 (N_14404,N_14009,N_14102);
xnor U14405 (N_14405,N_14204,N_14016);
nand U14406 (N_14406,N_14004,N_14021);
nand U14407 (N_14407,N_14026,N_14103);
nor U14408 (N_14408,N_14117,N_14069);
or U14409 (N_14409,N_14025,N_14131);
and U14410 (N_14410,N_14222,N_14145);
xor U14411 (N_14411,N_14126,N_14181);
nor U14412 (N_14412,N_14149,N_14010);
and U14413 (N_14413,N_14242,N_14090);
xnor U14414 (N_14414,N_14073,N_14124);
nor U14415 (N_14415,N_14239,N_14057);
or U14416 (N_14416,N_14084,N_14172);
and U14417 (N_14417,N_14035,N_14099);
xnor U14418 (N_14418,N_14174,N_14138);
and U14419 (N_14419,N_14032,N_14017);
or U14420 (N_14420,N_14216,N_14009);
xnor U14421 (N_14421,N_14152,N_14195);
or U14422 (N_14422,N_14133,N_14058);
nor U14423 (N_14423,N_14049,N_14181);
and U14424 (N_14424,N_14129,N_14053);
and U14425 (N_14425,N_14183,N_14134);
and U14426 (N_14426,N_14219,N_14032);
or U14427 (N_14427,N_14141,N_14077);
or U14428 (N_14428,N_14147,N_14063);
nor U14429 (N_14429,N_14145,N_14213);
and U14430 (N_14430,N_14180,N_14222);
xor U14431 (N_14431,N_14235,N_14142);
nand U14432 (N_14432,N_14243,N_14046);
or U14433 (N_14433,N_14113,N_14186);
xnor U14434 (N_14434,N_14030,N_14003);
nor U14435 (N_14435,N_14088,N_14047);
nor U14436 (N_14436,N_14158,N_14205);
nand U14437 (N_14437,N_14247,N_14229);
xnor U14438 (N_14438,N_14063,N_14107);
nor U14439 (N_14439,N_14047,N_14086);
nor U14440 (N_14440,N_14029,N_14231);
nand U14441 (N_14441,N_14146,N_14085);
or U14442 (N_14442,N_14216,N_14235);
or U14443 (N_14443,N_14143,N_14105);
nor U14444 (N_14444,N_14227,N_14178);
xor U14445 (N_14445,N_14119,N_14147);
and U14446 (N_14446,N_14164,N_14037);
xor U14447 (N_14447,N_14220,N_14238);
or U14448 (N_14448,N_14247,N_14053);
and U14449 (N_14449,N_14069,N_14011);
and U14450 (N_14450,N_14067,N_14151);
nor U14451 (N_14451,N_14207,N_14219);
xor U14452 (N_14452,N_14237,N_14057);
xor U14453 (N_14453,N_14061,N_14018);
nand U14454 (N_14454,N_14003,N_14193);
xnor U14455 (N_14455,N_14005,N_14017);
nor U14456 (N_14456,N_14046,N_14248);
xnor U14457 (N_14457,N_14244,N_14157);
xor U14458 (N_14458,N_14193,N_14229);
or U14459 (N_14459,N_14111,N_14094);
nand U14460 (N_14460,N_14100,N_14185);
or U14461 (N_14461,N_14142,N_14052);
xor U14462 (N_14462,N_14168,N_14093);
nor U14463 (N_14463,N_14079,N_14004);
xor U14464 (N_14464,N_14140,N_14107);
nand U14465 (N_14465,N_14142,N_14152);
nand U14466 (N_14466,N_14144,N_14186);
nor U14467 (N_14467,N_14063,N_14144);
nand U14468 (N_14468,N_14033,N_14132);
xnor U14469 (N_14469,N_14135,N_14218);
or U14470 (N_14470,N_14060,N_14224);
nor U14471 (N_14471,N_14150,N_14169);
or U14472 (N_14472,N_14029,N_14217);
xor U14473 (N_14473,N_14166,N_14210);
and U14474 (N_14474,N_14029,N_14171);
or U14475 (N_14475,N_14188,N_14128);
and U14476 (N_14476,N_14134,N_14217);
or U14477 (N_14477,N_14104,N_14175);
or U14478 (N_14478,N_14167,N_14224);
xor U14479 (N_14479,N_14074,N_14035);
and U14480 (N_14480,N_14154,N_14176);
and U14481 (N_14481,N_14180,N_14183);
xnor U14482 (N_14482,N_14051,N_14196);
or U14483 (N_14483,N_14155,N_14054);
nor U14484 (N_14484,N_14048,N_14138);
nor U14485 (N_14485,N_14243,N_14144);
or U14486 (N_14486,N_14072,N_14015);
and U14487 (N_14487,N_14073,N_14011);
nor U14488 (N_14488,N_14128,N_14168);
nor U14489 (N_14489,N_14065,N_14082);
and U14490 (N_14490,N_14062,N_14166);
xnor U14491 (N_14491,N_14239,N_14064);
or U14492 (N_14492,N_14054,N_14062);
and U14493 (N_14493,N_14113,N_14131);
or U14494 (N_14494,N_14110,N_14243);
nand U14495 (N_14495,N_14202,N_14064);
nand U14496 (N_14496,N_14011,N_14128);
nand U14497 (N_14497,N_14120,N_14212);
xor U14498 (N_14498,N_14180,N_14192);
xnor U14499 (N_14499,N_14100,N_14136);
and U14500 (N_14500,N_14405,N_14308);
or U14501 (N_14501,N_14366,N_14499);
or U14502 (N_14502,N_14256,N_14387);
xnor U14503 (N_14503,N_14435,N_14395);
nor U14504 (N_14504,N_14461,N_14365);
or U14505 (N_14505,N_14425,N_14282);
nor U14506 (N_14506,N_14351,N_14289);
nor U14507 (N_14507,N_14454,N_14414);
or U14508 (N_14508,N_14310,N_14474);
xor U14509 (N_14509,N_14274,N_14498);
nand U14510 (N_14510,N_14327,N_14406);
and U14511 (N_14511,N_14350,N_14369);
or U14512 (N_14512,N_14300,N_14312);
xor U14513 (N_14513,N_14400,N_14285);
nand U14514 (N_14514,N_14403,N_14401);
and U14515 (N_14515,N_14311,N_14367);
nand U14516 (N_14516,N_14415,N_14298);
nand U14517 (N_14517,N_14456,N_14421);
xor U14518 (N_14518,N_14412,N_14373);
nor U14519 (N_14519,N_14441,N_14331);
or U14520 (N_14520,N_14437,N_14330);
and U14521 (N_14521,N_14294,N_14480);
xor U14522 (N_14522,N_14303,N_14397);
or U14523 (N_14523,N_14463,N_14320);
and U14524 (N_14524,N_14464,N_14445);
nor U14525 (N_14525,N_14388,N_14278);
and U14526 (N_14526,N_14460,N_14264);
and U14527 (N_14527,N_14283,N_14384);
and U14528 (N_14528,N_14432,N_14270);
xor U14529 (N_14529,N_14391,N_14426);
nor U14530 (N_14530,N_14375,N_14396);
xnor U14531 (N_14531,N_14496,N_14255);
xor U14532 (N_14532,N_14494,N_14433);
nand U14533 (N_14533,N_14321,N_14313);
nor U14534 (N_14534,N_14402,N_14329);
and U14535 (N_14535,N_14355,N_14328);
nand U14536 (N_14536,N_14483,N_14385);
nand U14537 (N_14537,N_14322,N_14446);
and U14538 (N_14538,N_14469,N_14343);
nand U14539 (N_14539,N_14348,N_14389);
xnor U14540 (N_14540,N_14491,N_14339);
nor U14541 (N_14541,N_14409,N_14394);
or U14542 (N_14542,N_14299,N_14301);
xnor U14543 (N_14543,N_14453,N_14497);
xor U14544 (N_14544,N_14377,N_14353);
nand U14545 (N_14545,N_14413,N_14368);
xnor U14546 (N_14546,N_14309,N_14419);
nor U14547 (N_14547,N_14281,N_14346);
nand U14548 (N_14548,N_14380,N_14418);
and U14549 (N_14549,N_14318,N_14315);
nor U14550 (N_14550,N_14493,N_14363);
and U14551 (N_14551,N_14332,N_14408);
nor U14552 (N_14552,N_14489,N_14471);
or U14553 (N_14553,N_14467,N_14374);
or U14554 (N_14554,N_14317,N_14361);
nand U14555 (N_14555,N_14338,N_14345);
or U14556 (N_14556,N_14268,N_14470);
or U14557 (N_14557,N_14280,N_14444);
nor U14558 (N_14558,N_14428,N_14344);
nor U14559 (N_14559,N_14487,N_14319);
or U14560 (N_14560,N_14360,N_14307);
or U14561 (N_14561,N_14447,N_14475);
and U14562 (N_14562,N_14459,N_14443);
or U14563 (N_14563,N_14481,N_14424);
xor U14564 (N_14564,N_14265,N_14258);
and U14565 (N_14565,N_14286,N_14257);
nor U14566 (N_14566,N_14485,N_14482);
xnor U14567 (N_14567,N_14290,N_14416);
nand U14568 (N_14568,N_14357,N_14293);
nor U14569 (N_14569,N_14383,N_14334);
nor U14570 (N_14570,N_14466,N_14295);
nor U14571 (N_14571,N_14336,N_14254);
and U14572 (N_14572,N_14381,N_14275);
and U14573 (N_14573,N_14362,N_14347);
xnor U14574 (N_14574,N_14392,N_14448);
and U14575 (N_14575,N_14455,N_14349);
nor U14576 (N_14576,N_14382,N_14273);
or U14577 (N_14577,N_14468,N_14324);
nor U14578 (N_14578,N_14335,N_14305);
nand U14579 (N_14579,N_14422,N_14266);
or U14580 (N_14580,N_14476,N_14279);
nand U14581 (N_14581,N_14252,N_14284);
xnor U14582 (N_14582,N_14378,N_14276);
or U14583 (N_14583,N_14462,N_14407);
xnor U14584 (N_14584,N_14423,N_14302);
xor U14585 (N_14585,N_14261,N_14304);
nand U14586 (N_14586,N_14393,N_14404);
and U14587 (N_14587,N_14417,N_14452);
and U14588 (N_14588,N_14398,N_14288);
nor U14589 (N_14589,N_14271,N_14352);
xnor U14590 (N_14590,N_14314,N_14478);
and U14591 (N_14591,N_14364,N_14267);
and U14592 (N_14592,N_14386,N_14439);
nor U14593 (N_14593,N_14420,N_14442);
nand U14594 (N_14594,N_14372,N_14259);
and U14595 (N_14595,N_14465,N_14296);
nand U14596 (N_14596,N_14434,N_14370);
and U14597 (N_14597,N_14292,N_14488);
and U14598 (N_14598,N_14251,N_14262);
nor U14599 (N_14599,N_14495,N_14333);
and U14600 (N_14600,N_14371,N_14427);
or U14601 (N_14601,N_14340,N_14399);
and U14602 (N_14602,N_14341,N_14287);
nor U14603 (N_14603,N_14376,N_14451);
xnor U14604 (N_14604,N_14306,N_14325);
nand U14605 (N_14605,N_14316,N_14356);
xor U14606 (N_14606,N_14450,N_14337);
xor U14607 (N_14607,N_14253,N_14297);
or U14608 (N_14608,N_14429,N_14477);
nand U14609 (N_14609,N_14277,N_14354);
nor U14610 (N_14610,N_14479,N_14438);
or U14611 (N_14611,N_14492,N_14359);
nor U14612 (N_14612,N_14291,N_14323);
or U14613 (N_14613,N_14457,N_14342);
nor U14614 (N_14614,N_14473,N_14326);
or U14615 (N_14615,N_14436,N_14484);
xnor U14616 (N_14616,N_14379,N_14449);
nor U14617 (N_14617,N_14458,N_14430);
nand U14618 (N_14618,N_14410,N_14260);
xnor U14619 (N_14619,N_14486,N_14358);
nor U14620 (N_14620,N_14272,N_14411);
or U14621 (N_14621,N_14250,N_14431);
xnor U14622 (N_14622,N_14390,N_14269);
or U14623 (N_14623,N_14490,N_14263);
and U14624 (N_14624,N_14440,N_14472);
nor U14625 (N_14625,N_14299,N_14451);
nand U14626 (N_14626,N_14415,N_14499);
and U14627 (N_14627,N_14323,N_14497);
nand U14628 (N_14628,N_14470,N_14389);
nor U14629 (N_14629,N_14470,N_14289);
xnor U14630 (N_14630,N_14330,N_14441);
nand U14631 (N_14631,N_14425,N_14445);
or U14632 (N_14632,N_14452,N_14460);
and U14633 (N_14633,N_14491,N_14349);
nor U14634 (N_14634,N_14407,N_14260);
xnor U14635 (N_14635,N_14477,N_14271);
and U14636 (N_14636,N_14346,N_14479);
xor U14637 (N_14637,N_14261,N_14323);
xnor U14638 (N_14638,N_14449,N_14392);
nand U14639 (N_14639,N_14347,N_14292);
nand U14640 (N_14640,N_14477,N_14321);
and U14641 (N_14641,N_14407,N_14469);
or U14642 (N_14642,N_14300,N_14357);
and U14643 (N_14643,N_14437,N_14268);
and U14644 (N_14644,N_14386,N_14322);
and U14645 (N_14645,N_14471,N_14469);
or U14646 (N_14646,N_14422,N_14411);
nand U14647 (N_14647,N_14427,N_14296);
and U14648 (N_14648,N_14292,N_14301);
and U14649 (N_14649,N_14266,N_14346);
or U14650 (N_14650,N_14373,N_14294);
xnor U14651 (N_14651,N_14262,N_14268);
nand U14652 (N_14652,N_14307,N_14293);
and U14653 (N_14653,N_14396,N_14414);
nand U14654 (N_14654,N_14262,N_14458);
nand U14655 (N_14655,N_14365,N_14436);
nor U14656 (N_14656,N_14397,N_14451);
xnor U14657 (N_14657,N_14298,N_14386);
xnor U14658 (N_14658,N_14292,N_14378);
nand U14659 (N_14659,N_14477,N_14373);
xor U14660 (N_14660,N_14465,N_14439);
xor U14661 (N_14661,N_14304,N_14442);
nor U14662 (N_14662,N_14276,N_14268);
xnor U14663 (N_14663,N_14399,N_14266);
nand U14664 (N_14664,N_14473,N_14300);
xnor U14665 (N_14665,N_14456,N_14345);
xnor U14666 (N_14666,N_14409,N_14370);
and U14667 (N_14667,N_14295,N_14306);
and U14668 (N_14668,N_14379,N_14292);
nor U14669 (N_14669,N_14344,N_14425);
and U14670 (N_14670,N_14317,N_14406);
xnor U14671 (N_14671,N_14447,N_14251);
and U14672 (N_14672,N_14272,N_14391);
xor U14673 (N_14673,N_14465,N_14484);
nor U14674 (N_14674,N_14385,N_14499);
nand U14675 (N_14675,N_14260,N_14325);
or U14676 (N_14676,N_14417,N_14455);
or U14677 (N_14677,N_14343,N_14405);
or U14678 (N_14678,N_14361,N_14432);
nor U14679 (N_14679,N_14389,N_14495);
xor U14680 (N_14680,N_14447,N_14252);
nor U14681 (N_14681,N_14368,N_14260);
nand U14682 (N_14682,N_14391,N_14261);
nor U14683 (N_14683,N_14482,N_14314);
nor U14684 (N_14684,N_14305,N_14475);
nand U14685 (N_14685,N_14486,N_14467);
xor U14686 (N_14686,N_14415,N_14259);
or U14687 (N_14687,N_14333,N_14254);
or U14688 (N_14688,N_14325,N_14356);
nand U14689 (N_14689,N_14393,N_14419);
nand U14690 (N_14690,N_14338,N_14356);
xor U14691 (N_14691,N_14264,N_14477);
or U14692 (N_14692,N_14403,N_14297);
nand U14693 (N_14693,N_14387,N_14424);
nor U14694 (N_14694,N_14335,N_14407);
xor U14695 (N_14695,N_14456,N_14461);
or U14696 (N_14696,N_14348,N_14357);
xor U14697 (N_14697,N_14476,N_14250);
nand U14698 (N_14698,N_14346,N_14381);
and U14699 (N_14699,N_14490,N_14359);
xnor U14700 (N_14700,N_14415,N_14426);
nand U14701 (N_14701,N_14493,N_14343);
nor U14702 (N_14702,N_14377,N_14410);
xor U14703 (N_14703,N_14403,N_14267);
or U14704 (N_14704,N_14416,N_14357);
nor U14705 (N_14705,N_14296,N_14277);
and U14706 (N_14706,N_14338,N_14405);
and U14707 (N_14707,N_14260,N_14371);
and U14708 (N_14708,N_14491,N_14309);
nand U14709 (N_14709,N_14447,N_14302);
xnor U14710 (N_14710,N_14307,N_14446);
nor U14711 (N_14711,N_14298,N_14286);
nand U14712 (N_14712,N_14317,N_14430);
nor U14713 (N_14713,N_14250,N_14399);
or U14714 (N_14714,N_14256,N_14352);
nor U14715 (N_14715,N_14283,N_14267);
nor U14716 (N_14716,N_14371,N_14309);
xor U14717 (N_14717,N_14417,N_14384);
nand U14718 (N_14718,N_14431,N_14427);
and U14719 (N_14719,N_14461,N_14442);
xnor U14720 (N_14720,N_14266,N_14429);
nand U14721 (N_14721,N_14477,N_14478);
and U14722 (N_14722,N_14329,N_14478);
or U14723 (N_14723,N_14276,N_14388);
xnor U14724 (N_14724,N_14391,N_14439);
and U14725 (N_14725,N_14447,N_14474);
xnor U14726 (N_14726,N_14370,N_14351);
xnor U14727 (N_14727,N_14340,N_14490);
nand U14728 (N_14728,N_14414,N_14451);
nor U14729 (N_14729,N_14495,N_14418);
nor U14730 (N_14730,N_14321,N_14467);
or U14731 (N_14731,N_14449,N_14270);
and U14732 (N_14732,N_14452,N_14441);
xor U14733 (N_14733,N_14465,N_14453);
nor U14734 (N_14734,N_14440,N_14280);
nand U14735 (N_14735,N_14330,N_14335);
or U14736 (N_14736,N_14471,N_14451);
xnor U14737 (N_14737,N_14450,N_14331);
xnor U14738 (N_14738,N_14420,N_14287);
or U14739 (N_14739,N_14432,N_14321);
or U14740 (N_14740,N_14250,N_14324);
nand U14741 (N_14741,N_14250,N_14284);
nor U14742 (N_14742,N_14264,N_14368);
and U14743 (N_14743,N_14310,N_14271);
and U14744 (N_14744,N_14432,N_14376);
and U14745 (N_14745,N_14347,N_14413);
xor U14746 (N_14746,N_14468,N_14415);
or U14747 (N_14747,N_14271,N_14331);
xor U14748 (N_14748,N_14262,N_14371);
or U14749 (N_14749,N_14370,N_14397);
nor U14750 (N_14750,N_14602,N_14661);
nor U14751 (N_14751,N_14622,N_14545);
xnor U14752 (N_14752,N_14615,N_14650);
or U14753 (N_14753,N_14646,N_14575);
nand U14754 (N_14754,N_14662,N_14532);
and U14755 (N_14755,N_14742,N_14673);
nor U14756 (N_14756,N_14749,N_14630);
xnor U14757 (N_14757,N_14583,N_14693);
nor U14758 (N_14758,N_14632,N_14550);
xnor U14759 (N_14759,N_14507,N_14525);
nor U14760 (N_14760,N_14704,N_14599);
or U14761 (N_14761,N_14741,N_14644);
xnor U14762 (N_14762,N_14537,N_14614);
nand U14763 (N_14763,N_14597,N_14730);
xnor U14764 (N_14764,N_14648,N_14732);
xor U14765 (N_14765,N_14544,N_14581);
or U14766 (N_14766,N_14682,N_14692);
and U14767 (N_14767,N_14721,N_14551);
and U14768 (N_14768,N_14707,N_14524);
or U14769 (N_14769,N_14720,N_14715);
or U14770 (N_14770,N_14556,N_14509);
nor U14771 (N_14771,N_14670,N_14685);
and U14772 (N_14772,N_14530,N_14526);
nor U14773 (N_14773,N_14563,N_14511);
or U14774 (N_14774,N_14686,N_14580);
and U14775 (N_14775,N_14728,N_14631);
or U14776 (N_14776,N_14633,N_14691);
xor U14777 (N_14777,N_14688,N_14744);
or U14778 (N_14778,N_14561,N_14642);
nor U14779 (N_14779,N_14578,N_14586);
and U14780 (N_14780,N_14598,N_14706);
xor U14781 (N_14781,N_14645,N_14664);
or U14782 (N_14782,N_14547,N_14536);
and U14783 (N_14783,N_14501,N_14699);
and U14784 (N_14784,N_14566,N_14625);
or U14785 (N_14785,N_14500,N_14723);
xnor U14786 (N_14786,N_14619,N_14674);
or U14787 (N_14787,N_14624,N_14710);
xnor U14788 (N_14788,N_14565,N_14639);
or U14789 (N_14789,N_14683,N_14609);
or U14790 (N_14790,N_14542,N_14521);
xor U14791 (N_14791,N_14520,N_14652);
nand U14792 (N_14792,N_14716,N_14560);
xor U14793 (N_14793,N_14747,N_14726);
or U14794 (N_14794,N_14522,N_14513);
nand U14795 (N_14795,N_14591,N_14668);
nor U14796 (N_14796,N_14745,N_14568);
xnor U14797 (N_14797,N_14594,N_14606);
nor U14798 (N_14798,N_14651,N_14623);
nor U14799 (N_14799,N_14512,N_14535);
or U14800 (N_14800,N_14722,N_14736);
xnor U14801 (N_14801,N_14548,N_14667);
nor U14802 (N_14802,N_14640,N_14653);
xor U14803 (N_14803,N_14641,N_14666);
nand U14804 (N_14804,N_14539,N_14684);
nor U14805 (N_14805,N_14689,N_14637);
or U14806 (N_14806,N_14617,N_14610);
and U14807 (N_14807,N_14600,N_14677);
or U14808 (N_14808,N_14712,N_14601);
nand U14809 (N_14809,N_14713,N_14654);
nor U14810 (N_14810,N_14517,N_14636);
xnor U14811 (N_14811,N_14621,N_14574);
nor U14812 (N_14812,N_14678,N_14502);
or U14813 (N_14813,N_14717,N_14572);
nor U14814 (N_14814,N_14629,N_14739);
nor U14815 (N_14815,N_14703,N_14660);
nand U14816 (N_14816,N_14675,N_14529);
nand U14817 (N_14817,N_14705,N_14604);
and U14818 (N_14818,N_14527,N_14523);
or U14819 (N_14819,N_14719,N_14571);
nor U14820 (N_14820,N_14725,N_14557);
or U14821 (N_14821,N_14538,N_14634);
nand U14822 (N_14822,N_14595,N_14649);
or U14823 (N_14823,N_14679,N_14553);
nand U14824 (N_14824,N_14737,N_14743);
xor U14825 (N_14825,N_14733,N_14540);
xnor U14826 (N_14826,N_14588,N_14697);
and U14827 (N_14827,N_14570,N_14573);
nand U14828 (N_14828,N_14549,N_14596);
and U14829 (N_14829,N_14554,N_14626);
xor U14830 (N_14830,N_14638,N_14504);
or U14831 (N_14831,N_14543,N_14603);
or U14832 (N_14832,N_14687,N_14593);
xnor U14833 (N_14833,N_14738,N_14711);
and U14834 (N_14834,N_14665,N_14718);
and U14835 (N_14835,N_14607,N_14559);
and U14836 (N_14836,N_14647,N_14681);
and U14837 (N_14837,N_14671,N_14735);
and U14838 (N_14838,N_14531,N_14505);
nor U14839 (N_14839,N_14616,N_14659);
nor U14840 (N_14840,N_14635,N_14672);
nand U14841 (N_14841,N_14727,N_14676);
nand U14842 (N_14842,N_14655,N_14714);
nor U14843 (N_14843,N_14669,N_14579);
and U14844 (N_14844,N_14695,N_14734);
or U14845 (N_14845,N_14533,N_14567);
and U14846 (N_14846,N_14541,N_14518);
or U14847 (N_14847,N_14577,N_14709);
and U14848 (N_14848,N_14611,N_14748);
or U14849 (N_14849,N_14508,N_14643);
and U14850 (N_14850,N_14576,N_14680);
xnor U14851 (N_14851,N_14503,N_14585);
nand U14852 (N_14852,N_14590,N_14569);
and U14853 (N_14853,N_14528,N_14584);
nor U14854 (N_14854,N_14562,N_14708);
xor U14855 (N_14855,N_14627,N_14582);
nand U14856 (N_14856,N_14663,N_14519);
nor U14857 (N_14857,N_14620,N_14564);
and U14858 (N_14858,N_14514,N_14558);
nand U14859 (N_14859,N_14534,N_14605);
or U14860 (N_14860,N_14516,N_14612);
and U14861 (N_14861,N_14618,N_14656);
or U14862 (N_14862,N_14552,N_14592);
and U14863 (N_14863,N_14658,N_14613);
and U14864 (N_14864,N_14724,N_14701);
or U14865 (N_14865,N_14628,N_14587);
xnor U14866 (N_14866,N_14698,N_14555);
or U14867 (N_14867,N_14506,N_14694);
nand U14868 (N_14868,N_14731,N_14700);
nand U14869 (N_14869,N_14589,N_14657);
nor U14870 (N_14870,N_14729,N_14546);
xnor U14871 (N_14871,N_14746,N_14510);
or U14872 (N_14872,N_14740,N_14702);
xnor U14873 (N_14873,N_14608,N_14690);
xnor U14874 (N_14874,N_14696,N_14515);
and U14875 (N_14875,N_14590,N_14527);
xnor U14876 (N_14876,N_14729,N_14628);
and U14877 (N_14877,N_14740,N_14534);
nor U14878 (N_14878,N_14501,N_14697);
nand U14879 (N_14879,N_14550,N_14596);
and U14880 (N_14880,N_14568,N_14715);
or U14881 (N_14881,N_14733,N_14675);
or U14882 (N_14882,N_14635,N_14708);
and U14883 (N_14883,N_14720,N_14697);
and U14884 (N_14884,N_14523,N_14692);
nand U14885 (N_14885,N_14655,N_14575);
and U14886 (N_14886,N_14748,N_14656);
nand U14887 (N_14887,N_14511,N_14679);
or U14888 (N_14888,N_14673,N_14656);
and U14889 (N_14889,N_14594,N_14655);
or U14890 (N_14890,N_14541,N_14622);
nor U14891 (N_14891,N_14736,N_14527);
nor U14892 (N_14892,N_14541,N_14587);
nand U14893 (N_14893,N_14747,N_14715);
nor U14894 (N_14894,N_14728,N_14724);
nor U14895 (N_14895,N_14573,N_14548);
and U14896 (N_14896,N_14518,N_14516);
or U14897 (N_14897,N_14669,N_14638);
or U14898 (N_14898,N_14599,N_14505);
nor U14899 (N_14899,N_14736,N_14580);
nand U14900 (N_14900,N_14606,N_14514);
nor U14901 (N_14901,N_14508,N_14628);
or U14902 (N_14902,N_14643,N_14578);
nor U14903 (N_14903,N_14594,N_14532);
and U14904 (N_14904,N_14626,N_14525);
and U14905 (N_14905,N_14683,N_14537);
or U14906 (N_14906,N_14660,N_14520);
xnor U14907 (N_14907,N_14697,N_14614);
and U14908 (N_14908,N_14705,N_14622);
and U14909 (N_14909,N_14528,N_14643);
nand U14910 (N_14910,N_14629,N_14636);
and U14911 (N_14911,N_14716,N_14722);
and U14912 (N_14912,N_14503,N_14727);
and U14913 (N_14913,N_14645,N_14572);
or U14914 (N_14914,N_14672,N_14578);
or U14915 (N_14915,N_14632,N_14647);
and U14916 (N_14916,N_14729,N_14595);
or U14917 (N_14917,N_14514,N_14632);
xnor U14918 (N_14918,N_14657,N_14678);
xor U14919 (N_14919,N_14608,N_14703);
nor U14920 (N_14920,N_14701,N_14720);
xor U14921 (N_14921,N_14700,N_14681);
or U14922 (N_14922,N_14604,N_14684);
nand U14923 (N_14923,N_14541,N_14630);
nand U14924 (N_14924,N_14539,N_14705);
nor U14925 (N_14925,N_14735,N_14626);
nand U14926 (N_14926,N_14650,N_14577);
nand U14927 (N_14927,N_14737,N_14722);
nor U14928 (N_14928,N_14738,N_14701);
xor U14929 (N_14929,N_14642,N_14749);
nand U14930 (N_14930,N_14654,N_14511);
or U14931 (N_14931,N_14526,N_14664);
nand U14932 (N_14932,N_14569,N_14700);
nor U14933 (N_14933,N_14680,N_14684);
nor U14934 (N_14934,N_14601,N_14733);
nand U14935 (N_14935,N_14630,N_14570);
xor U14936 (N_14936,N_14563,N_14659);
and U14937 (N_14937,N_14596,N_14580);
nand U14938 (N_14938,N_14576,N_14706);
nand U14939 (N_14939,N_14715,N_14604);
nor U14940 (N_14940,N_14721,N_14662);
or U14941 (N_14941,N_14731,N_14604);
nor U14942 (N_14942,N_14532,N_14629);
nor U14943 (N_14943,N_14726,N_14713);
and U14944 (N_14944,N_14527,N_14516);
xor U14945 (N_14945,N_14748,N_14630);
nand U14946 (N_14946,N_14718,N_14659);
xor U14947 (N_14947,N_14581,N_14687);
nor U14948 (N_14948,N_14555,N_14582);
xnor U14949 (N_14949,N_14504,N_14583);
nor U14950 (N_14950,N_14711,N_14532);
nand U14951 (N_14951,N_14589,N_14663);
nand U14952 (N_14952,N_14673,N_14581);
or U14953 (N_14953,N_14725,N_14540);
nor U14954 (N_14954,N_14707,N_14596);
and U14955 (N_14955,N_14624,N_14679);
nor U14956 (N_14956,N_14519,N_14616);
and U14957 (N_14957,N_14675,N_14512);
and U14958 (N_14958,N_14544,N_14600);
nand U14959 (N_14959,N_14653,N_14525);
nand U14960 (N_14960,N_14608,N_14738);
nand U14961 (N_14961,N_14509,N_14506);
and U14962 (N_14962,N_14569,N_14589);
nor U14963 (N_14963,N_14606,N_14571);
and U14964 (N_14964,N_14665,N_14609);
xnor U14965 (N_14965,N_14651,N_14711);
nand U14966 (N_14966,N_14611,N_14731);
or U14967 (N_14967,N_14641,N_14693);
and U14968 (N_14968,N_14607,N_14522);
or U14969 (N_14969,N_14503,N_14673);
nand U14970 (N_14970,N_14672,N_14687);
nand U14971 (N_14971,N_14627,N_14688);
nor U14972 (N_14972,N_14628,N_14724);
xor U14973 (N_14973,N_14681,N_14654);
and U14974 (N_14974,N_14600,N_14518);
xnor U14975 (N_14975,N_14739,N_14674);
nand U14976 (N_14976,N_14661,N_14702);
and U14977 (N_14977,N_14642,N_14604);
xnor U14978 (N_14978,N_14550,N_14690);
and U14979 (N_14979,N_14674,N_14575);
nor U14980 (N_14980,N_14560,N_14681);
or U14981 (N_14981,N_14640,N_14630);
xor U14982 (N_14982,N_14565,N_14573);
and U14983 (N_14983,N_14649,N_14668);
or U14984 (N_14984,N_14638,N_14629);
nand U14985 (N_14985,N_14730,N_14678);
and U14986 (N_14986,N_14689,N_14569);
or U14987 (N_14987,N_14516,N_14708);
xnor U14988 (N_14988,N_14513,N_14597);
nand U14989 (N_14989,N_14538,N_14697);
and U14990 (N_14990,N_14574,N_14578);
or U14991 (N_14991,N_14683,N_14569);
and U14992 (N_14992,N_14692,N_14561);
xor U14993 (N_14993,N_14731,N_14584);
and U14994 (N_14994,N_14591,N_14584);
and U14995 (N_14995,N_14587,N_14663);
or U14996 (N_14996,N_14594,N_14745);
nor U14997 (N_14997,N_14530,N_14604);
nor U14998 (N_14998,N_14699,N_14537);
nor U14999 (N_14999,N_14739,N_14712);
and UO_0 (O_0,N_14992,N_14905);
or UO_1 (O_1,N_14769,N_14934);
nor UO_2 (O_2,N_14790,N_14820);
or UO_3 (O_3,N_14877,N_14796);
xor UO_4 (O_4,N_14948,N_14809);
and UO_5 (O_5,N_14823,N_14837);
or UO_6 (O_6,N_14861,N_14800);
nand UO_7 (O_7,N_14920,N_14806);
or UO_8 (O_8,N_14856,N_14901);
xor UO_9 (O_9,N_14828,N_14761);
or UO_10 (O_10,N_14960,N_14838);
xnor UO_11 (O_11,N_14989,N_14768);
and UO_12 (O_12,N_14902,N_14950);
nand UO_13 (O_13,N_14914,N_14762);
and UO_14 (O_14,N_14954,N_14967);
and UO_15 (O_15,N_14883,N_14864);
nor UO_16 (O_16,N_14813,N_14835);
nor UO_17 (O_17,N_14816,N_14787);
nor UO_18 (O_18,N_14918,N_14965);
or UO_19 (O_19,N_14781,N_14840);
or UO_20 (O_20,N_14939,N_14943);
or UO_21 (O_21,N_14855,N_14925);
or UO_22 (O_22,N_14897,N_14824);
nand UO_23 (O_23,N_14789,N_14894);
or UO_24 (O_24,N_14770,N_14872);
nor UO_25 (O_25,N_14750,N_14944);
nand UO_26 (O_26,N_14827,N_14871);
nand UO_27 (O_27,N_14926,N_14974);
xor UO_28 (O_28,N_14988,N_14869);
or UO_29 (O_29,N_14910,N_14912);
xnor UO_30 (O_30,N_14915,N_14839);
xor UO_31 (O_31,N_14756,N_14945);
or UO_32 (O_32,N_14962,N_14969);
or UO_33 (O_33,N_14999,N_14981);
or UO_34 (O_34,N_14830,N_14868);
or UO_35 (O_35,N_14972,N_14807);
xor UO_36 (O_36,N_14975,N_14968);
and UO_37 (O_37,N_14986,N_14777);
nand UO_38 (O_38,N_14997,N_14983);
xnor UO_39 (O_39,N_14977,N_14998);
or UO_40 (O_40,N_14832,N_14793);
nand UO_41 (O_41,N_14956,N_14859);
nor UO_42 (O_42,N_14775,N_14848);
xnor UO_43 (O_43,N_14985,N_14963);
xor UO_44 (O_44,N_14792,N_14845);
nand UO_45 (O_45,N_14879,N_14980);
nand UO_46 (O_46,N_14996,N_14755);
xnor UO_47 (O_47,N_14825,N_14888);
or UO_48 (O_48,N_14971,N_14922);
and UO_49 (O_49,N_14862,N_14782);
nand UO_50 (O_50,N_14976,N_14913);
or UO_51 (O_51,N_14812,N_14929);
xor UO_52 (O_52,N_14849,N_14919);
or UO_53 (O_53,N_14936,N_14810);
or UO_54 (O_54,N_14779,N_14909);
nand UO_55 (O_55,N_14904,N_14784);
and UO_56 (O_56,N_14785,N_14966);
and UO_57 (O_57,N_14842,N_14884);
nor UO_58 (O_58,N_14937,N_14941);
or UO_59 (O_59,N_14771,N_14766);
nand UO_60 (O_60,N_14819,N_14763);
or UO_61 (O_61,N_14895,N_14942);
xor UO_62 (O_62,N_14927,N_14878);
xnor UO_63 (O_63,N_14978,N_14911);
or UO_64 (O_64,N_14958,N_14955);
or UO_65 (O_65,N_14858,N_14931);
nor UO_66 (O_66,N_14778,N_14951);
nand UO_67 (O_67,N_14882,N_14860);
nand UO_68 (O_68,N_14984,N_14814);
or UO_69 (O_69,N_14818,N_14938);
nor UO_70 (O_70,N_14794,N_14921);
nand UO_71 (O_71,N_14853,N_14788);
or UO_72 (O_72,N_14887,N_14893);
nor UO_73 (O_73,N_14906,N_14822);
nand UO_74 (O_74,N_14854,N_14767);
or UO_75 (O_75,N_14876,N_14908);
nand UO_76 (O_76,N_14940,N_14765);
nor UO_77 (O_77,N_14896,N_14973);
and UO_78 (O_78,N_14804,N_14817);
nand UO_79 (O_79,N_14844,N_14892);
nor UO_80 (O_80,N_14783,N_14791);
xnor UO_81 (O_81,N_14760,N_14851);
nor UO_82 (O_82,N_14841,N_14776);
xnor UO_83 (O_83,N_14970,N_14885);
and UO_84 (O_84,N_14875,N_14917);
and UO_85 (O_85,N_14863,N_14933);
and UO_86 (O_86,N_14852,N_14786);
xor UO_87 (O_87,N_14898,N_14886);
xnor UO_88 (O_88,N_14991,N_14773);
nand UO_89 (O_89,N_14964,N_14959);
nand UO_90 (O_90,N_14881,N_14952);
xor UO_91 (O_91,N_14774,N_14752);
nand UO_92 (O_92,N_14847,N_14801);
nand UO_93 (O_93,N_14759,N_14754);
nor UO_94 (O_94,N_14994,N_14753);
nor UO_95 (O_95,N_14826,N_14873);
or UO_96 (O_96,N_14982,N_14949);
xor UO_97 (O_97,N_14799,N_14757);
xnor UO_98 (O_98,N_14870,N_14993);
or UO_99 (O_99,N_14798,N_14836);
nand UO_100 (O_100,N_14990,N_14815);
and UO_101 (O_101,N_14808,N_14903);
xor UO_102 (O_102,N_14865,N_14821);
or UO_103 (O_103,N_14907,N_14946);
nor UO_104 (O_104,N_14843,N_14803);
xnor UO_105 (O_105,N_14850,N_14772);
or UO_106 (O_106,N_14758,N_14957);
nor UO_107 (O_107,N_14995,N_14834);
xnor UO_108 (O_108,N_14890,N_14795);
and UO_109 (O_109,N_14866,N_14916);
or UO_110 (O_110,N_14924,N_14805);
or UO_111 (O_111,N_14857,N_14928);
or UO_112 (O_112,N_14979,N_14899);
nor UO_113 (O_113,N_14797,N_14867);
and UO_114 (O_114,N_14953,N_14935);
xnor UO_115 (O_115,N_14880,N_14930);
nor UO_116 (O_116,N_14829,N_14846);
and UO_117 (O_117,N_14947,N_14802);
or UO_118 (O_118,N_14831,N_14889);
and UO_119 (O_119,N_14811,N_14780);
nor UO_120 (O_120,N_14923,N_14874);
or UO_121 (O_121,N_14932,N_14751);
or UO_122 (O_122,N_14891,N_14900);
xor UO_123 (O_123,N_14833,N_14987);
xnor UO_124 (O_124,N_14764,N_14961);
or UO_125 (O_125,N_14764,N_14814);
or UO_126 (O_126,N_14894,N_14857);
xnor UO_127 (O_127,N_14872,N_14889);
xor UO_128 (O_128,N_14887,N_14879);
and UO_129 (O_129,N_14982,N_14940);
or UO_130 (O_130,N_14875,N_14833);
xnor UO_131 (O_131,N_14838,N_14890);
nor UO_132 (O_132,N_14887,N_14884);
nor UO_133 (O_133,N_14976,N_14838);
nor UO_134 (O_134,N_14924,N_14823);
or UO_135 (O_135,N_14961,N_14936);
or UO_136 (O_136,N_14776,N_14942);
xor UO_137 (O_137,N_14854,N_14775);
or UO_138 (O_138,N_14750,N_14909);
or UO_139 (O_139,N_14905,N_14954);
or UO_140 (O_140,N_14780,N_14917);
or UO_141 (O_141,N_14988,N_14945);
xnor UO_142 (O_142,N_14841,N_14949);
and UO_143 (O_143,N_14812,N_14825);
and UO_144 (O_144,N_14820,N_14988);
and UO_145 (O_145,N_14972,N_14825);
nand UO_146 (O_146,N_14863,N_14751);
and UO_147 (O_147,N_14864,N_14903);
xnor UO_148 (O_148,N_14905,N_14847);
nor UO_149 (O_149,N_14910,N_14882);
nor UO_150 (O_150,N_14850,N_14833);
nand UO_151 (O_151,N_14774,N_14909);
and UO_152 (O_152,N_14892,N_14951);
nand UO_153 (O_153,N_14807,N_14961);
nor UO_154 (O_154,N_14816,N_14756);
xnor UO_155 (O_155,N_14816,N_14826);
and UO_156 (O_156,N_14900,N_14754);
and UO_157 (O_157,N_14829,N_14912);
nand UO_158 (O_158,N_14940,N_14846);
and UO_159 (O_159,N_14923,N_14776);
nand UO_160 (O_160,N_14964,N_14819);
or UO_161 (O_161,N_14795,N_14809);
and UO_162 (O_162,N_14876,N_14930);
or UO_163 (O_163,N_14783,N_14775);
xor UO_164 (O_164,N_14822,N_14902);
or UO_165 (O_165,N_14857,N_14977);
nand UO_166 (O_166,N_14755,N_14808);
and UO_167 (O_167,N_14835,N_14969);
nand UO_168 (O_168,N_14828,N_14783);
or UO_169 (O_169,N_14828,N_14774);
and UO_170 (O_170,N_14869,N_14909);
nand UO_171 (O_171,N_14986,N_14823);
nand UO_172 (O_172,N_14903,N_14752);
nor UO_173 (O_173,N_14933,N_14907);
nand UO_174 (O_174,N_14897,N_14757);
nor UO_175 (O_175,N_14884,N_14931);
or UO_176 (O_176,N_14750,N_14843);
nor UO_177 (O_177,N_14926,N_14855);
nor UO_178 (O_178,N_14848,N_14880);
and UO_179 (O_179,N_14893,N_14894);
xor UO_180 (O_180,N_14797,N_14980);
nand UO_181 (O_181,N_14959,N_14797);
xnor UO_182 (O_182,N_14983,N_14825);
and UO_183 (O_183,N_14789,N_14885);
nand UO_184 (O_184,N_14757,N_14768);
and UO_185 (O_185,N_14956,N_14851);
nand UO_186 (O_186,N_14864,N_14782);
or UO_187 (O_187,N_14988,N_14895);
xnor UO_188 (O_188,N_14917,N_14968);
and UO_189 (O_189,N_14817,N_14972);
or UO_190 (O_190,N_14793,N_14831);
or UO_191 (O_191,N_14910,N_14903);
and UO_192 (O_192,N_14949,N_14976);
and UO_193 (O_193,N_14831,N_14821);
or UO_194 (O_194,N_14809,N_14787);
and UO_195 (O_195,N_14763,N_14751);
nand UO_196 (O_196,N_14825,N_14950);
nand UO_197 (O_197,N_14763,N_14958);
nor UO_198 (O_198,N_14986,N_14806);
or UO_199 (O_199,N_14930,N_14891);
xor UO_200 (O_200,N_14970,N_14987);
or UO_201 (O_201,N_14926,N_14901);
nand UO_202 (O_202,N_14847,N_14840);
or UO_203 (O_203,N_14974,N_14982);
nand UO_204 (O_204,N_14864,N_14763);
or UO_205 (O_205,N_14949,N_14765);
and UO_206 (O_206,N_14791,N_14961);
or UO_207 (O_207,N_14780,N_14962);
and UO_208 (O_208,N_14785,N_14999);
nor UO_209 (O_209,N_14912,N_14985);
xnor UO_210 (O_210,N_14939,N_14820);
xnor UO_211 (O_211,N_14891,N_14967);
xnor UO_212 (O_212,N_14964,N_14838);
xnor UO_213 (O_213,N_14904,N_14862);
and UO_214 (O_214,N_14864,N_14771);
nor UO_215 (O_215,N_14990,N_14890);
nor UO_216 (O_216,N_14951,N_14986);
and UO_217 (O_217,N_14951,N_14960);
xor UO_218 (O_218,N_14978,N_14957);
nor UO_219 (O_219,N_14981,N_14775);
or UO_220 (O_220,N_14966,N_14866);
and UO_221 (O_221,N_14877,N_14803);
nor UO_222 (O_222,N_14930,N_14826);
xor UO_223 (O_223,N_14846,N_14826);
nand UO_224 (O_224,N_14798,N_14925);
and UO_225 (O_225,N_14833,N_14827);
or UO_226 (O_226,N_14966,N_14910);
xor UO_227 (O_227,N_14764,N_14903);
nor UO_228 (O_228,N_14950,N_14845);
or UO_229 (O_229,N_14993,N_14780);
and UO_230 (O_230,N_14861,N_14867);
nor UO_231 (O_231,N_14979,N_14862);
xnor UO_232 (O_232,N_14857,N_14953);
nand UO_233 (O_233,N_14800,N_14893);
and UO_234 (O_234,N_14971,N_14833);
nand UO_235 (O_235,N_14805,N_14954);
or UO_236 (O_236,N_14916,N_14803);
or UO_237 (O_237,N_14946,N_14861);
or UO_238 (O_238,N_14784,N_14926);
and UO_239 (O_239,N_14800,N_14810);
and UO_240 (O_240,N_14784,N_14999);
xnor UO_241 (O_241,N_14781,N_14834);
and UO_242 (O_242,N_14951,N_14842);
xnor UO_243 (O_243,N_14868,N_14997);
and UO_244 (O_244,N_14926,N_14873);
nor UO_245 (O_245,N_14926,N_14990);
nor UO_246 (O_246,N_14971,N_14811);
and UO_247 (O_247,N_14980,N_14818);
nand UO_248 (O_248,N_14906,N_14762);
xor UO_249 (O_249,N_14861,N_14875);
xor UO_250 (O_250,N_14987,N_14930);
xnor UO_251 (O_251,N_14976,N_14841);
or UO_252 (O_252,N_14792,N_14920);
and UO_253 (O_253,N_14874,N_14888);
or UO_254 (O_254,N_14766,N_14763);
nand UO_255 (O_255,N_14755,N_14824);
or UO_256 (O_256,N_14773,N_14969);
nor UO_257 (O_257,N_14894,N_14768);
or UO_258 (O_258,N_14877,N_14829);
and UO_259 (O_259,N_14814,N_14979);
nand UO_260 (O_260,N_14906,N_14871);
or UO_261 (O_261,N_14909,N_14829);
and UO_262 (O_262,N_14761,N_14926);
or UO_263 (O_263,N_14988,N_14807);
nand UO_264 (O_264,N_14975,N_14947);
or UO_265 (O_265,N_14918,N_14896);
xnor UO_266 (O_266,N_14963,N_14824);
nand UO_267 (O_267,N_14754,N_14875);
xor UO_268 (O_268,N_14822,N_14859);
or UO_269 (O_269,N_14987,N_14975);
xnor UO_270 (O_270,N_14815,N_14874);
or UO_271 (O_271,N_14991,N_14783);
nand UO_272 (O_272,N_14918,N_14949);
xnor UO_273 (O_273,N_14847,N_14879);
nand UO_274 (O_274,N_14991,N_14875);
and UO_275 (O_275,N_14885,N_14754);
nand UO_276 (O_276,N_14847,N_14877);
and UO_277 (O_277,N_14968,N_14775);
and UO_278 (O_278,N_14834,N_14922);
or UO_279 (O_279,N_14941,N_14812);
xnor UO_280 (O_280,N_14811,N_14912);
and UO_281 (O_281,N_14884,N_14882);
nand UO_282 (O_282,N_14802,N_14841);
xor UO_283 (O_283,N_14961,N_14783);
nor UO_284 (O_284,N_14771,N_14880);
and UO_285 (O_285,N_14775,N_14928);
or UO_286 (O_286,N_14945,N_14882);
nand UO_287 (O_287,N_14907,N_14792);
nor UO_288 (O_288,N_14917,N_14845);
nand UO_289 (O_289,N_14786,N_14870);
nor UO_290 (O_290,N_14939,N_14803);
xor UO_291 (O_291,N_14797,N_14759);
or UO_292 (O_292,N_14757,N_14921);
xor UO_293 (O_293,N_14852,N_14916);
or UO_294 (O_294,N_14940,N_14752);
nor UO_295 (O_295,N_14754,N_14837);
and UO_296 (O_296,N_14988,N_14792);
nor UO_297 (O_297,N_14977,N_14940);
nand UO_298 (O_298,N_14944,N_14802);
or UO_299 (O_299,N_14918,N_14968);
nand UO_300 (O_300,N_14898,N_14973);
and UO_301 (O_301,N_14994,N_14907);
nor UO_302 (O_302,N_14894,N_14972);
and UO_303 (O_303,N_14889,N_14882);
nor UO_304 (O_304,N_14905,N_14766);
nand UO_305 (O_305,N_14965,N_14846);
and UO_306 (O_306,N_14916,N_14874);
xor UO_307 (O_307,N_14972,N_14782);
and UO_308 (O_308,N_14813,N_14850);
or UO_309 (O_309,N_14905,N_14999);
or UO_310 (O_310,N_14925,N_14837);
and UO_311 (O_311,N_14926,N_14911);
and UO_312 (O_312,N_14826,N_14986);
or UO_313 (O_313,N_14851,N_14878);
or UO_314 (O_314,N_14954,N_14775);
or UO_315 (O_315,N_14929,N_14761);
nand UO_316 (O_316,N_14926,N_14892);
and UO_317 (O_317,N_14833,N_14959);
nand UO_318 (O_318,N_14866,N_14962);
or UO_319 (O_319,N_14872,N_14794);
or UO_320 (O_320,N_14820,N_14892);
nor UO_321 (O_321,N_14778,N_14841);
nand UO_322 (O_322,N_14931,N_14829);
or UO_323 (O_323,N_14879,N_14763);
or UO_324 (O_324,N_14871,N_14847);
and UO_325 (O_325,N_14892,N_14827);
nor UO_326 (O_326,N_14818,N_14766);
and UO_327 (O_327,N_14781,N_14779);
nor UO_328 (O_328,N_14782,N_14905);
or UO_329 (O_329,N_14949,N_14810);
xor UO_330 (O_330,N_14788,N_14782);
xnor UO_331 (O_331,N_14860,N_14822);
nand UO_332 (O_332,N_14992,N_14955);
nand UO_333 (O_333,N_14942,N_14900);
or UO_334 (O_334,N_14873,N_14793);
xor UO_335 (O_335,N_14891,N_14882);
xor UO_336 (O_336,N_14801,N_14961);
xor UO_337 (O_337,N_14957,N_14759);
and UO_338 (O_338,N_14797,N_14838);
and UO_339 (O_339,N_14976,N_14921);
nand UO_340 (O_340,N_14813,N_14918);
and UO_341 (O_341,N_14816,N_14913);
xnor UO_342 (O_342,N_14851,N_14960);
nor UO_343 (O_343,N_14984,N_14874);
nand UO_344 (O_344,N_14831,N_14988);
or UO_345 (O_345,N_14849,N_14978);
xnor UO_346 (O_346,N_14826,N_14791);
xor UO_347 (O_347,N_14882,N_14879);
or UO_348 (O_348,N_14959,N_14993);
nor UO_349 (O_349,N_14778,N_14862);
or UO_350 (O_350,N_14752,N_14904);
xor UO_351 (O_351,N_14760,N_14962);
xor UO_352 (O_352,N_14753,N_14918);
xnor UO_353 (O_353,N_14954,N_14940);
nor UO_354 (O_354,N_14913,N_14897);
or UO_355 (O_355,N_14846,N_14866);
xnor UO_356 (O_356,N_14757,N_14874);
nand UO_357 (O_357,N_14868,N_14989);
nand UO_358 (O_358,N_14839,N_14809);
and UO_359 (O_359,N_14889,N_14858);
xor UO_360 (O_360,N_14812,N_14756);
nor UO_361 (O_361,N_14941,N_14790);
and UO_362 (O_362,N_14862,N_14843);
and UO_363 (O_363,N_14847,N_14962);
xnor UO_364 (O_364,N_14989,N_14908);
nand UO_365 (O_365,N_14829,N_14989);
xnor UO_366 (O_366,N_14853,N_14887);
xnor UO_367 (O_367,N_14805,N_14766);
nand UO_368 (O_368,N_14843,N_14857);
or UO_369 (O_369,N_14840,N_14887);
xor UO_370 (O_370,N_14844,N_14888);
nor UO_371 (O_371,N_14837,N_14994);
and UO_372 (O_372,N_14862,N_14968);
nand UO_373 (O_373,N_14797,N_14978);
or UO_374 (O_374,N_14930,N_14997);
and UO_375 (O_375,N_14843,N_14994);
nor UO_376 (O_376,N_14915,N_14976);
xor UO_377 (O_377,N_14982,N_14892);
nand UO_378 (O_378,N_14926,N_14824);
or UO_379 (O_379,N_14841,N_14796);
xnor UO_380 (O_380,N_14902,N_14827);
nor UO_381 (O_381,N_14964,N_14968);
and UO_382 (O_382,N_14782,N_14764);
and UO_383 (O_383,N_14832,N_14955);
and UO_384 (O_384,N_14956,N_14818);
or UO_385 (O_385,N_14969,N_14857);
xor UO_386 (O_386,N_14848,N_14750);
nor UO_387 (O_387,N_14903,N_14918);
nand UO_388 (O_388,N_14971,N_14929);
nand UO_389 (O_389,N_14990,N_14857);
nand UO_390 (O_390,N_14750,N_14966);
nor UO_391 (O_391,N_14779,N_14959);
nor UO_392 (O_392,N_14932,N_14970);
and UO_393 (O_393,N_14999,N_14982);
and UO_394 (O_394,N_14902,N_14759);
xor UO_395 (O_395,N_14914,N_14871);
nand UO_396 (O_396,N_14759,N_14900);
nor UO_397 (O_397,N_14876,N_14879);
xnor UO_398 (O_398,N_14809,N_14894);
or UO_399 (O_399,N_14947,N_14974);
xnor UO_400 (O_400,N_14927,N_14793);
xor UO_401 (O_401,N_14921,N_14866);
or UO_402 (O_402,N_14969,N_14958);
nor UO_403 (O_403,N_14815,N_14797);
xnor UO_404 (O_404,N_14864,N_14766);
nand UO_405 (O_405,N_14871,N_14919);
or UO_406 (O_406,N_14756,N_14778);
xor UO_407 (O_407,N_14967,N_14884);
nand UO_408 (O_408,N_14766,N_14944);
xor UO_409 (O_409,N_14766,N_14758);
or UO_410 (O_410,N_14781,N_14849);
nand UO_411 (O_411,N_14902,N_14771);
nand UO_412 (O_412,N_14780,N_14788);
or UO_413 (O_413,N_14976,N_14985);
xor UO_414 (O_414,N_14871,N_14928);
nand UO_415 (O_415,N_14767,N_14948);
nor UO_416 (O_416,N_14953,N_14961);
nand UO_417 (O_417,N_14975,N_14903);
nor UO_418 (O_418,N_14871,N_14789);
and UO_419 (O_419,N_14755,N_14826);
xor UO_420 (O_420,N_14898,N_14787);
nor UO_421 (O_421,N_14902,N_14762);
or UO_422 (O_422,N_14934,N_14920);
xnor UO_423 (O_423,N_14785,N_14857);
and UO_424 (O_424,N_14899,N_14938);
and UO_425 (O_425,N_14789,N_14754);
nand UO_426 (O_426,N_14762,N_14870);
xor UO_427 (O_427,N_14942,N_14981);
nor UO_428 (O_428,N_14782,N_14952);
nor UO_429 (O_429,N_14789,N_14874);
and UO_430 (O_430,N_14854,N_14962);
or UO_431 (O_431,N_14825,N_14842);
and UO_432 (O_432,N_14830,N_14976);
or UO_433 (O_433,N_14847,N_14949);
xnor UO_434 (O_434,N_14825,N_14829);
and UO_435 (O_435,N_14826,N_14931);
xor UO_436 (O_436,N_14910,N_14997);
or UO_437 (O_437,N_14928,N_14826);
and UO_438 (O_438,N_14995,N_14790);
nand UO_439 (O_439,N_14845,N_14760);
or UO_440 (O_440,N_14939,N_14897);
xnor UO_441 (O_441,N_14948,N_14887);
and UO_442 (O_442,N_14849,N_14958);
and UO_443 (O_443,N_14964,N_14989);
xnor UO_444 (O_444,N_14838,N_14977);
nand UO_445 (O_445,N_14901,N_14888);
nor UO_446 (O_446,N_14998,N_14982);
xnor UO_447 (O_447,N_14933,N_14948);
nand UO_448 (O_448,N_14822,N_14833);
xnor UO_449 (O_449,N_14865,N_14911);
nand UO_450 (O_450,N_14911,N_14854);
xnor UO_451 (O_451,N_14914,N_14975);
and UO_452 (O_452,N_14917,N_14771);
xor UO_453 (O_453,N_14783,N_14811);
nand UO_454 (O_454,N_14960,N_14996);
nor UO_455 (O_455,N_14798,N_14921);
nor UO_456 (O_456,N_14751,N_14954);
nand UO_457 (O_457,N_14991,N_14835);
or UO_458 (O_458,N_14799,N_14761);
nand UO_459 (O_459,N_14818,N_14848);
nor UO_460 (O_460,N_14919,N_14806);
xnor UO_461 (O_461,N_14808,N_14818);
or UO_462 (O_462,N_14955,N_14947);
xor UO_463 (O_463,N_14959,N_14950);
and UO_464 (O_464,N_14845,N_14894);
nor UO_465 (O_465,N_14954,N_14956);
and UO_466 (O_466,N_14898,N_14968);
and UO_467 (O_467,N_14891,N_14777);
nor UO_468 (O_468,N_14867,N_14964);
nand UO_469 (O_469,N_14900,N_14863);
xor UO_470 (O_470,N_14960,N_14822);
or UO_471 (O_471,N_14923,N_14796);
nor UO_472 (O_472,N_14862,N_14881);
nand UO_473 (O_473,N_14760,N_14954);
nand UO_474 (O_474,N_14900,N_14791);
and UO_475 (O_475,N_14807,N_14936);
nand UO_476 (O_476,N_14756,N_14860);
and UO_477 (O_477,N_14882,N_14940);
xor UO_478 (O_478,N_14920,N_14826);
nand UO_479 (O_479,N_14893,N_14750);
or UO_480 (O_480,N_14782,N_14790);
nor UO_481 (O_481,N_14828,N_14859);
or UO_482 (O_482,N_14803,N_14874);
nor UO_483 (O_483,N_14878,N_14947);
nor UO_484 (O_484,N_14850,N_14920);
or UO_485 (O_485,N_14876,N_14922);
and UO_486 (O_486,N_14935,N_14974);
xnor UO_487 (O_487,N_14899,N_14820);
and UO_488 (O_488,N_14976,N_14845);
and UO_489 (O_489,N_14802,N_14826);
nand UO_490 (O_490,N_14925,N_14861);
nand UO_491 (O_491,N_14970,N_14867);
and UO_492 (O_492,N_14777,N_14801);
xnor UO_493 (O_493,N_14832,N_14855);
and UO_494 (O_494,N_14888,N_14913);
and UO_495 (O_495,N_14860,N_14787);
nand UO_496 (O_496,N_14885,N_14913);
xnor UO_497 (O_497,N_14919,N_14788);
xor UO_498 (O_498,N_14875,N_14817);
nor UO_499 (O_499,N_14770,N_14867);
and UO_500 (O_500,N_14871,N_14840);
nand UO_501 (O_501,N_14995,N_14785);
and UO_502 (O_502,N_14832,N_14815);
nor UO_503 (O_503,N_14768,N_14818);
and UO_504 (O_504,N_14766,N_14867);
nor UO_505 (O_505,N_14784,N_14817);
xnor UO_506 (O_506,N_14896,N_14924);
and UO_507 (O_507,N_14822,N_14965);
or UO_508 (O_508,N_14761,N_14790);
xnor UO_509 (O_509,N_14836,N_14918);
nand UO_510 (O_510,N_14829,N_14995);
nand UO_511 (O_511,N_14827,N_14935);
and UO_512 (O_512,N_14861,N_14945);
nor UO_513 (O_513,N_14834,N_14847);
or UO_514 (O_514,N_14771,N_14894);
nor UO_515 (O_515,N_14884,N_14927);
xor UO_516 (O_516,N_14972,N_14987);
or UO_517 (O_517,N_14894,N_14777);
nand UO_518 (O_518,N_14797,N_14839);
nor UO_519 (O_519,N_14847,N_14812);
or UO_520 (O_520,N_14866,N_14838);
nor UO_521 (O_521,N_14883,N_14986);
and UO_522 (O_522,N_14864,N_14777);
and UO_523 (O_523,N_14901,N_14920);
nor UO_524 (O_524,N_14919,N_14845);
and UO_525 (O_525,N_14922,N_14868);
or UO_526 (O_526,N_14927,N_14798);
or UO_527 (O_527,N_14932,N_14819);
xnor UO_528 (O_528,N_14893,N_14755);
nor UO_529 (O_529,N_14805,N_14932);
or UO_530 (O_530,N_14786,N_14825);
xor UO_531 (O_531,N_14757,N_14761);
xor UO_532 (O_532,N_14912,N_14922);
and UO_533 (O_533,N_14910,N_14878);
nand UO_534 (O_534,N_14855,N_14789);
nand UO_535 (O_535,N_14941,N_14772);
nor UO_536 (O_536,N_14893,N_14824);
or UO_537 (O_537,N_14998,N_14989);
nand UO_538 (O_538,N_14945,N_14754);
xor UO_539 (O_539,N_14751,N_14817);
and UO_540 (O_540,N_14822,N_14924);
or UO_541 (O_541,N_14897,N_14978);
and UO_542 (O_542,N_14791,N_14976);
or UO_543 (O_543,N_14819,N_14807);
or UO_544 (O_544,N_14989,N_14909);
nand UO_545 (O_545,N_14797,N_14998);
nand UO_546 (O_546,N_14807,N_14928);
or UO_547 (O_547,N_14804,N_14986);
nand UO_548 (O_548,N_14973,N_14826);
nor UO_549 (O_549,N_14955,N_14840);
xnor UO_550 (O_550,N_14867,N_14788);
or UO_551 (O_551,N_14952,N_14808);
and UO_552 (O_552,N_14949,N_14937);
or UO_553 (O_553,N_14834,N_14952);
nor UO_554 (O_554,N_14856,N_14889);
nor UO_555 (O_555,N_14937,N_14818);
nor UO_556 (O_556,N_14760,N_14792);
or UO_557 (O_557,N_14966,N_14791);
and UO_558 (O_558,N_14807,N_14895);
and UO_559 (O_559,N_14783,N_14952);
nor UO_560 (O_560,N_14782,N_14923);
or UO_561 (O_561,N_14953,N_14919);
or UO_562 (O_562,N_14813,N_14899);
xnor UO_563 (O_563,N_14793,N_14789);
xor UO_564 (O_564,N_14929,N_14979);
xnor UO_565 (O_565,N_14880,N_14844);
nor UO_566 (O_566,N_14941,N_14890);
xnor UO_567 (O_567,N_14842,N_14801);
xor UO_568 (O_568,N_14821,N_14764);
and UO_569 (O_569,N_14892,N_14877);
and UO_570 (O_570,N_14943,N_14956);
or UO_571 (O_571,N_14868,N_14773);
or UO_572 (O_572,N_14922,N_14993);
nand UO_573 (O_573,N_14862,N_14888);
xor UO_574 (O_574,N_14802,N_14775);
and UO_575 (O_575,N_14964,N_14909);
and UO_576 (O_576,N_14818,N_14862);
or UO_577 (O_577,N_14761,N_14944);
and UO_578 (O_578,N_14962,N_14945);
xor UO_579 (O_579,N_14829,N_14925);
nand UO_580 (O_580,N_14912,N_14871);
nor UO_581 (O_581,N_14968,N_14895);
and UO_582 (O_582,N_14955,N_14975);
and UO_583 (O_583,N_14785,N_14771);
and UO_584 (O_584,N_14889,N_14811);
nor UO_585 (O_585,N_14798,N_14946);
and UO_586 (O_586,N_14787,N_14942);
nor UO_587 (O_587,N_14848,N_14955);
nand UO_588 (O_588,N_14888,N_14795);
xor UO_589 (O_589,N_14812,N_14947);
nor UO_590 (O_590,N_14929,N_14796);
xor UO_591 (O_591,N_14816,N_14818);
and UO_592 (O_592,N_14846,N_14772);
nor UO_593 (O_593,N_14772,N_14842);
xor UO_594 (O_594,N_14868,N_14751);
nor UO_595 (O_595,N_14839,N_14793);
nor UO_596 (O_596,N_14994,N_14847);
xor UO_597 (O_597,N_14856,N_14861);
nand UO_598 (O_598,N_14882,N_14876);
xnor UO_599 (O_599,N_14845,N_14821);
xnor UO_600 (O_600,N_14769,N_14809);
xnor UO_601 (O_601,N_14971,N_14830);
nor UO_602 (O_602,N_14956,N_14774);
nor UO_603 (O_603,N_14866,N_14857);
nor UO_604 (O_604,N_14789,N_14853);
nand UO_605 (O_605,N_14842,N_14936);
or UO_606 (O_606,N_14819,N_14867);
or UO_607 (O_607,N_14938,N_14963);
nor UO_608 (O_608,N_14999,N_14753);
nand UO_609 (O_609,N_14839,N_14922);
and UO_610 (O_610,N_14775,N_14914);
nand UO_611 (O_611,N_14877,N_14789);
nand UO_612 (O_612,N_14834,N_14757);
and UO_613 (O_613,N_14890,N_14823);
nor UO_614 (O_614,N_14941,N_14853);
and UO_615 (O_615,N_14987,N_14850);
nand UO_616 (O_616,N_14991,N_14809);
nand UO_617 (O_617,N_14959,N_14931);
nor UO_618 (O_618,N_14924,N_14934);
nor UO_619 (O_619,N_14971,N_14787);
xnor UO_620 (O_620,N_14858,N_14828);
or UO_621 (O_621,N_14883,N_14882);
nor UO_622 (O_622,N_14894,N_14950);
nor UO_623 (O_623,N_14874,N_14946);
nand UO_624 (O_624,N_14856,N_14975);
nor UO_625 (O_625,N_14861,N_14838);
or UO_626 (O_626,N_14752,N_14786);
nor UO_627 (O_627,N_14893,N_14891);
nand UO_628 (O_628,N_14974,N_14894);
or UO_629 (O_629,N_14752,N_14753);
nor UO_630 (O_630,N_14808,N_14913);
or UO_631 (O_631,N_14777,N_14878);
or UO_632 (O_632,N_14945,N_14759);
nand UO_633 (O_633,N_14856,N_14785);
nor UO_634 (O_634,N_14949,N_14792);
nor UO_635 (O_635,N_14756,N_14894);
and UO_636 (O_636,N_14923,N_14913);
xor UO_637 (O_637,N_14943,N_14804);
nand UO_638 (O_638,N_14779,N_14960);
nand UO_639 (O_639,N_14937,N_14791);
nor UO_640 (O_640,N_14896,N_14945);
xor UO_641 (O_641,N_14945,N_14825);
xor UO_642 (O_642,N_14971,N_14968);
nand UO_643 (O_643,N_14950,N_14849);
xor UO_644 (O_644,N_14952,N_14809);
and UO_645 (O_645,N_14972,N_14841);
nor UO_646 (O_646,N_14970,N_14774);
nor UO_647 (O_647,N_14978,N_14872);
nand UO_648 (O_648,N_14877,N_14922);
nor UO_649 (O_649,N_14947,N_14969);
xnor UO_650 (O_650,N_14966,N_14904);
nand UO_651 (O_651,N_14778,N_14908);
or UO_652 (O_652,N_14784,N_14916);
nor UO_653 (O_653,N_14773,N_14886);
and UO_654 (O_654,N_14757,N_14993);
nor UO_655 (O_655,N_14777,N_14903);
nand UO_656 (O_656,N_14930,N_14879);
nor UO_657 (O_657,N_14842,N_14913);
xnor UO_658 (O_658,N_14868,N_14939);
or UO_659 (O_659,N_14870,N_14869);
or UO_660 (O_660,N_14938,N_14826);
and UO_661 (O_661,N_14949,N_14957);
nor UO_662 (O_662,N_14793,N_14997);
or UO_663 (O_663,N_14794,N_14803);
nand UO_664 (O_664,N_14758,N_14796);
nor UO_665 (O_665,N_14786,N_14773);
nor UO_666 (O_666,N_14912,N_14776);
nor UO_667 (O_667,N_14859,N_14837);
or UO_668 (O_668,N_14963,N_14781);
xor UO_669 (O_669,N_14864,N_14811);
xnor UO_670 (O_670,N_14909,N_14948);
nor UO_671 (O_671,N_14895,N_14824);
nor UO_672 (O_672,N_14854,N_14836);
nand UO_673 (O_673,N_14861,N_14827);
nor UO_674 (O_674,N_14948,N_14992);
or UO_675 (O_675,N_14823,N_14964);
or UO_676 (O_676,N_14918,N_14859);
or UO_677 (O_677,N_14866,N_14961);
or UO_678 (O_678,N_14926,N_14816);
and UO_679 (O_679,N_14923,N_14891);
nand UO_680 (O_680,N_14788,N_14894);
nor UO_681 (O_681,N_14850,N_14873);
nand UO_682 (O_682,N_14965,N_14815);
xor UO_683 (O_683,N_14763,N_14895);
nand UO_684 (O_684,N_14880,N_14917);
nand UO_685 (O_685,N_14810,N_14791);
nand UO_686 (O_686,N_14979,N_14799);
nand UO_687 (O_687,N_14984,N_14987);
xnor UO_688 (O_688,N_14823,N_14884);
nor UO_689 (O_689,N_14934,N_14806);
and UO_690 (O_690,N_14821,N_14788);
and UO_691 (O_691,N_14990,N_14953);
and UO_692 (O_692,N_14845,N_14902);
xor UO_693 (O_693,N_14814,N_14793);
nor UO_694 (O_694,N_14966,N_14967);
nor UO_695 (O_695,N_14895,N_14970);
nor UO_696 (O_696,N_14811,N_14983);
and UO_697 (O_697,N_14794,N_14785);
and UO_698 (O_698,N_14916,N_14793);
nor UO_699 (O_699,N_14772,N_14847);
nor UO_700 (O_700,N_14971,N_14997);
and UO_701 (O_701,N_14843,N_14755);
or UO_702 (O_702,N_14809,N_14812);
nor UO_703 (O_703,N_14804,N_14872);
xor UO_704 (O_704,N_14995,N_14963);
nand UO_705 (O_705,N_14979,N_14839);
and UO_706 (O_706,N_14803,N_14986);
and UO_707 (O_707,N_14827,N_14777);
xnor UO_708 (O_708,N_14811,N_14816);
nand UO_709 (O_709,N_14818,N_14750);
xnor UO_710 (O_710,N_14952,N_14939);
xnor UO_711 (O_711,N_14992,N_14835);
and UO_712 (O_712,N_14942,N_14939);
xor UO_713 (O_713,N_14958,N_14852);
xnor UO_714 (O_714,N_14966,N_14809);
and UO_715 (O_715,N_14823,N_14832);
xor UO_716 (O_716,N_14875,N_14855);
or UO_717 (O_717,N_14946,N_14901);
and UO_718 (O_718,N_14912,N_14939);
or UO_719 (O_719,N_14905,N_14818);
or UO_720 (O_720,N_14795,N_14937);
nor UO_721 (O_721,N_14796,N_14948);
nor UO_722 (O_722,N_14896,N_14776);
and UO_723 (O_723,N_14862,N_14855);
nor UO_724 (O_724,N_14764,N_14801);
or UO_725 (O_725,N_14859,N_14818);
xor UO_726 (O_726,N_14898,N_14937);
xnor UO_727 (O_727,N_14913,N_14938);
xnor UO_728 (O_728,N_14779,N_14753);
nand UO_729 (O_729,N_14862,N_14998);
nor UO_730 (O_730,N_14766,N_14980);
nor UO_731 (O_731,N_14767,N_14768);
or UO_732 (O_732,N_14852,N_14859);
nor UO_733 (O_733,N_14872,N_14893);
nor UO_734 (O_734,N_14957,N_14817);
nor UO_735 (O_735,N_14974,N_14816);
nor UO_736 (O_736,N_14779,N_14924);
or UO_737 (O_737,N_14940,N_14845);
xor UO_738 (O_738,N_14799,N_14918);
and UO_739 (O_739,N_14847,N_14904);
nor UO_740 (O_740,N_14997,N_14940);
nor UO_741 (O_741,N_14893,N_14866);
and UO_742 (O_742,N_14900,N_14837);
xor UO_743 (O_743,N_14805,N_14861);
xnor UO_744 (O_744,N_14880,N_14960);
and UO_745 (O_745,N_14976,N_14818);
or UO_746 (O_746,N_14827,N_14880);
nor UO_747 (O_747,N_14809,N_14763);
or UO_748 (O_748,N_14907,N_14924);
and UO_749 (O_749,N_14800,N_14801);
nand UO_750 (O_750,N_14764,N_14959);
xor UO_751 (O_751,N_14850,N_14874);
xor UO_752 (O_752,N_14889,N_14762);
nor UO_753 (O_753,N_14964,N_14984);
xor UO_754 (O_754,N_14806,N_14834);
and UO_755 (O_755,N_14970,N_14791);
nand UO_756 (O_756,N_14920,N_14973);
and UO_757 (O_757,N_14850,N_14957);
xnor UO_758 (O_758,N_14801,N_14992);
xnor UO_759 (O_759,N_14961,N_14805);
nor UO_760 (O_760,N_14854,N_14966);
and UO_761 (O_761,N_14877,N_14761);
nand UO_762 (O_762,N_14862,N_14988);
or UO_763 (O_763,N_14985,N_14787);
and UO_764 (O_764,N_14758,N_14779);
or UO_765 (O_765,N_14826,N_14810);
nand UO_766 (O_766,N_14786,N_14763);
xnor UO_767 (O_767,N_14949,N_14972);
or UO_768 (O_768,N_14795,N_14964);
or UO_769 (O_769,N_14785,N_14950);
nand UO_770 (O_770,N_14956,N_14868);
nor UO_771 (O_771,N_14758,N_14847);
nand UO_772 (O_772,N_14821,N_14908);
xor UO_773 (O_773,N_14774,N_14898);
or UO_774 (O_774,N_14926,N_14835);
and UO_775 (O_775,N_14986,N_14750);
xor UO_776 (O_776,N_14884,N_14981);
or UO_777 (O_777,N_14937,N_14800);
and UO_778 (O_778,N_14980,N_14765);
xnor UO_779 (O_779,N_14760,N_14859);
or UO_780 (O_780,N_14810,N_14918);
and UO_781 (O_781,N_14865,N_14951);
or UO_782 (O_782,N_14893,N_14832);
nand UO_783 (O_783,N_14843,N_14953);
xnor UO_784 (O_784,N_14928,N_14787);
xor UO_785 (O_785,N_14804,N_14933);
nand UO_786 (O_786,N_14906,N_14986);
nand UO_787 (O_787,N_14810,N_14992);
and UO_788 (O_788,N_14862,N_14820);
xnor UO_789 (O_789,N_14981,N_14991);
nor UO_790 (O_790,N_14923,N_14800);
xor UO_791 (O_791,N_14876,N_14987);
and UO_792 (O_792,N_14852,N_14850);
nand UO_793 (O_793,N_14899,N_14961);
nand UO_794 (O_794,N_14795,N_14801);
nand UO_795 (O_795,N_14807,N_14863);
xnor UO_796 (O_796,N_14968,N_14904);
and UO_797 (O_797,N_14770,N_14781);
xnor UO_798 (O_798,N_14774,N_14837);
or UO_799 (O_799,N_14790,N_14976);
xor UO_800 (O_800,N_14770,N_14883);
and UO_801 (O_801,N_14969,N_14751);
nand UO_802 (O_802,N_14781,N_14848);
nor UO_803 (O_803,N_14767,N_14887);
nor UO_804 (O_804,N_14819,N_14750);
and UO_805 (O_805,N_14950,N_14806);
and UO_806 (O_806,N_14874,N_14832);
and UO_807 (O_807,N_14925,N_14845);
and UO_808 (O_808,N_14813,N_14796);
xnor UO_809 (O_809,N_14806,N_14771);
or UO_810 (O_810,N_14807,N_14838);
nor UO_811 (O_811,N_14800,N_14764);
nand UO_812 (O_812,N_14956,N_14897);
nor UO_813 (O_813,N_14846,N_14921);
xor UO_814 (O_814,N_14953,N_14966);
nand UO_815 (O_815,N_14826,N_14862);
or UO_816 (O_816,N_14815,N_14757);
nand UO_817 (O_817,N_14968,N_14825);
xor UO_818 (O_818,N_14790,N_14989);
nor UO_819 (O_819,N_14922,N_14924);
nor UO_820 (O_820,N_14935,N_14945);
and UO_821 (O_821,N_14810,N_14875);
xor UO_822 (O_822,N_14980,N_14834);
xnor UO_823 (O_823,N_14751,N_14885);
or UO_824 (O_824,N_14981,N_14919);
nor UO_825 (O_825,N_14937,N_14985);
nand UO_826 (O_826,N_14797,N_14802);
nand UO_827 (O_827,N_14867,N_14975);
xor UO_828 (O_828,N_14890,N_14779);
nor UO_829 (O_829,N_14886,N_14881);
or UO_830 (O_830,N_14785,N_14911);
xnor UO_831 (O_831,N_14991,N_14976);
and UO_832 (O_832,N_14945,N_14845);
xor UO_833 (O_833,N_14934,N_14961);
nor UO_834 (O_834,N_14933,N_14999);
xor UO_835 (O_835,N_14773,N_14881);
or UO_836 (O_836,N_14888,N_14918);
or UO_837 (O_837,N_14883,N_14756);
and UO_838 (O_838,N_14840,N_14976);
xnor UO_839 (O_839,N_14991,N_14822);
xnor UO_840 (O_840,N_14965,N_14790);
nor UO_841 (O_841,N_14920,N_14897);
and UO_842 (O_842,N_14762,N_14883);
xor UO_843 (O_843,N_14767,N_14972);
xor UO_844 (O_844,N_14964,N_14818);
or UO_845 (O_845,N_14866,N_14799);
nor UO_846 (O_846,N_14988,N_14864);
nor UO_847 (O_847,N_14853,N_14912);
nand UO_848 (O_848,N_14918,N_14982);
xnor UO_849 (O_849,N_14904,N_14812);
xor UO_850 (O_850,N_14807,N_14926);
xnor UO_851 (O_851,N_14921,N_14937);
and UO_852 (O_852,N_14941,N_14858);
nor UO_853 (O_853,N_14906,N_14957);
xnor UO_854 (O_854,N_14826,N_14889);
nand UO_855 (O_855,N_14846,N_14926);
nand UO_856 (O_856,N_14933,N_14868);
nand UO_857 (O_857,N_14850,N_14979);
and UO_858 (O_858,N_14824,N_14977);
nand UO_859 (O_859,N_14865,N_14979);
nor UO_860 (O_860,N_14788,N_14808);
and UO_861 (O_861,N_14926,N_14934);
or UO_862 (O_862,N_14846,N_14901);
nand UO_863 (O_863,N_14997,N_14803);
and UO_864 (O_864,N_14828,N_14807);
nand UO_865 (O_865,N_14987,N_14881);
and UO_866 (O_866,N_14849,N_14927);
nand UO_867 (O_867,N_14819,N_14846);
xor UO_868 (O_868,N_14777,N_14797);
and UO_869 (O_869,N_14832,N_14784);
or UO_870 (O_870,N_14874,N_14961);
nor UO_871 (O_871,N_14990,N_14956);
nand UO_872 (O_872,N_14914,N_14938);
xor UO_873 (O_873,N_14885,N_14791);
and UO_874 (O_874,N_14983,N_14928);
nor UO_875 (O_875,N_14870,N_14998);
or UO_876 (O_876,N_14940,N_14794);
xor UO_877 (O_877,N_14996,N_14949);
or UO_878 (O_878,N_14790,N_14847);
or UO_879 (O_879,N_14868,N_14898);
and UO_880 (O_880,N_14898,N_14880);
and UO_881 (O_881,N_14902,N_14758);
and UO_882 (O_882,N_14902,N_14911);
nor UO_883 (O_883,N_14932,N_14788);
nand UO_884 (O_884,N_14772,N_14965);
nand UO_885 (O_885,N_14923,N_14952);
nor UO_886 (O_886,N_14770,N_14868);
xnor UO_887 (O_887,N_14980,N_14895);
and UO_888 (O_888,N_14992,N_14858);
or UO_889 (O_889,N_14936,N_14958);
nand UO_890 (O_890,N_14763,N_14868);
or UO_891 (O_891,N_14991,N_14982);
xnor UO_892 (O_892,N_14918,N_14923);
nand UO_893 (O_893,N_14870,N_14834);
xnor UO_894 (O_894,N_14883,N_14889);
and UO_895 (O_895,N_14983,N_14927);
and UO_896 (O_896,N_14977,N_14969);
nand UO_897 (O_897,N_14812,N_14907);
or UO_898 (O_898,N_14760,N_14944);
and UO_899 (O_899,N_14855,N_14929);
nand UO_900 (O_900,N_14807,N_14767);
nor UO_901 (O_901,N_14830,N_14791);
xnor UO_902 (O_902,N_14859,N_14782);
nand UO_903 (O_903,N_14851,N_14957);
xor UO_904 (O_904,N_14768,N_14754);
xnor UO_905 (O_905,N_14801,N_14948);
nor UO_906 (O_906,N_14756,N_14807);
and UO_907 (O_907,N_14855,N_14842);
nand UO_908 (O_908,N_14788,N_14985);
nand UO_909 (O_909,N_14781,N_14951);
xor UO_910 (O_910,N_14945,N_14897);
nor UO_911 (O_911,N_14921,N_14872);
nand UO_912 (O_912,N_14754,N_14827);
xor UO_913 (O_913,N_14795,N_14950);
xnor UO_914 (O_914,N_14965,N_14829);
nor UO_915 (O_915,N_14753,N_14896);
xnor UO_916 (O_916,N_14908,N_14837);
or UO_917 (O_917,N_14768,N_14996);
xnor UO_918 (O_918,N_14953,N_14997);
or UO_919 (O_919,N_14956,N_14891);
nand UO_920 (O_920,N_14786,N_14751);
or UO_921 (O_921,N_14940,N_14860);
nor UO_922 (O_922,N_14857,N_14954);
xor UO_923 (O_923,N_14929,N_14962);
nor UO_924 (O_924,N_14945,N_14956);
nor UO_925 (O_925,N_14858,N_14891);
and UO_926 (O_926,N_14788,N_14895);
and UO_927 (O_927,N_14756,N_14925);
xnor UO_928 (O_928,N_14843,N_14938);
or UO_929 (O_929,N_14754,N_14819);
nor UO_930 (O_930,N_14956,N_14819);
nand UO_931 (O_931,N_14870,N_14945);
nor UO_932 (O_932,N_14973,N_14854);
or UO_933 (O_933,N_14901,N_14949);
and UO_934 (O_934,N_14804,N_14906);
and UO_935 (O_935,N_14972,N_14988);
and UO_936 (O_936,N_14828,N_14837);
and UO_937 (O_937,N_14754,N_14866);
or UO_938 (O_938,N_14809,N_14887);
nor UO_939 (O_939,N_14936,N_14959);
nand UO_940 (O_940,N_14950,N_14909);
nand UO_941 (O_941,N_14908,N_14854);
nand UO_942 (O_942,N_14947,N_14786);
nand UO_943 (O_943,N_14769,N_14944);
xnor UO_944 (O_944,N_14813,N_14854);
nor UO_945 (O_945,N_14871,N_14941);
and UO_946 (O_946,N_14782,N_14964);
xor UO_947 (O_947,N_14785,N_14763);
or UO_948 (O_948,N_14935,N_14984);
nor UO_949 (O_949,N_14947,N_14847);
xnor UO_950 (O_950,N_14795,N_14840);
nand UO_951 (O_951,N_14914,N_14892);
nand UO_952 (O_952,N_14973,N_14874);
xnor UO_953 (O_953,N_14787,N_14818);
nand UO_954 (O_954,N_14951,N_14760);
and UO_955 (O_955,N_14980,N_14947);
or UO_956 (O_956,N_14844,N_14860);
nand UO_957 (O_957,N_14843,N_14870);
xnor UO_958 (O_958,N_14844,N_14900);
and UO_959 (O_959,N_14900,N_14815);
nand UO_960 (O_960,N_14828,N_14993);
nor UO_961 (O_961,N_14821,N_14989);
nand UO_962 (O_962,N_14817,N_14823);
or UO_963 (O_963,N_14897,N_14976);
or UO_964 (O_964,N_14921,N_14969);
and UO_965 (O_965,N_14949,N_14846);
or UO_966 (O_966,N_14870,N_14879);
or UO_967 (O_967,N_14889,N_14950);
nor UO_968 (O_968,N_14892,N_14756);
xnor UO_969 (O_969,N_14984,N_14751);
or UO_970 (O_970,N_14839,N_14765);
nor UO_971 (O_971,N_14892,N_14988);
xor UO_972 (O_972,N_14952,N_14760);
xnor UO_973 (O_973,N_14805,N_14951);
nand UO_974 (O_974,N_14835,N_14890);
nor UO_975 (O_975,N_14933,N_14959);
xor UO_976 (O_976,N_14873,N_14809);
xnor UO_977 (O_977,N_14995,N_14850);
or UO_978 (O_978,N_14874,N_14921);
and UO_979 (O_979,N_14863,N_14767);
and UO_980 (O_980,N_14765,N_14800);
or UO_981 (O_981,N_14786,N_14836);
nor UO_982 (O_982,N_14862,N_14986);
nor UO_983 (O_983,N_14875,N_14907);
and UO_984 (O_984,N_14938,N_14893);
and UO_985 (O_985,N_14811,N_14965);
and UO_986 (O_986,N_14944,N_14956);
nand UO_987 (O_987,N_14965,N_14776);
and UO_988 (O_988,N_14963,N_14998);
nand UO_989 (O_989,N_14786,N_14817);
nor UO_990 (O_990,N_14753,N_14929);
nor UO_991 (O_991,N_14835,N_14757);
xnor UO_992 (O_992,N_14906,N_14868);
or UO_993 (O_993,N_14915,N_14859);
or UO_994 (O_994,N_14899,N_14781);
nand UO_995 (O_995,N_14877,N_14819);
or UO_996 (O_996,N_14985,N_14983);
nor UO_997 (O_997,N_14882,N_14806);
and UO_998 (O_998,N_14817,N_14881);
nand UO_999 (O_999,N_14862,N_14926);
nand UO_1000 (O_1000,N_14920,N_14959);
nand UO_1001 (O_1001,N_14918,N_14864);
or UO_1002 (O_1002,N_14808,N_14950);
xnor UO_1003 (O_1003,N_14940,N_14920);
nor UO_1004 (O_1004,N_14759,N_14809);
nand UO_1005 (O_1005,N_14988,N_14986);
xnor UO_1006 (O_1006,N_14958,N_14832);
nand UO_1007 (O_1007,N_14790,N_14792);
xnor UO_1008 (O_1008,N_14935,N_14936);
nand UO_1009 (O_1009,N_14938,N_14960);
and UO_1010 (O_1010,N_14783,N_14998);
xor UO_1011 (O_1011,N_14894,N_14848);
and UO_1012 (O_1012,N_14872,N_14865);
or UO_1013 (O_1013,N_14751,N_14929);
and UO_1014 (O_1014,N_14917,N_14923);
xor UO_1015 (O_1015,N_14992,N_14791);
or UO_1016 (O_1016,N_14948,N_14775);
nand UO_1017 (O_1017,N_14757,N_14776);
and UO_1018 (O_1018,N_14786,N_14809);
nor UO_1019 (O_1019,N_14752,N_14815);
nand UO_1020 (O_1020,N_14964,N_14751);
xor UO_1021 (O_1021,N_14814,N_14973);
nand UO_1022 (O_1022,N_14882,N_14815);
and UO_1023 (O_1023,N_14862,N_14751);
nand UO_1024 (O_1024,N_14966,N_14994);
nor UO_1025 (O_1025,N_14911,N_14887);
nor UO_1026 (O_1026,N_14870,N_14898);
and UO_1027 (O_1027,N_14870,N_14829);
nor UO_1028 (O_1028,N_14822,N_14890);
xnor UO_1029 (O_1029,N_14783,N_14766);
nor UO_1030 (O_1030,N_14751,N_14914);
nand UO_1031 (O_1031,N_14825,N_14758);
nand UO_1032 (O_1032,N_14789,N_14895);
nand UO_1033 (O_1033,N_14849,N_14907);
nand UO_1034 (O_1034,N_14866,N_14906);
nor UO_1035 (O_1035,N_14892,N_14848);
or UO_1036 (O_1036,N_14959,N_14877);
nor UO_1037 (O_1037,N_14893,N_14954);
and UO_1038 (O_1038,N_14832,N_14957);
and UO_1039 (O_1039,N_14915,N_14808);
nand UO_1040 (O_1040,N_14963,N_14888);
xor UO_1041 (O_1041,N_14769,N_14880);
or UO_1042 (O_1042,N_14949,N_14856);
nand UO_1043 (O_1043,N_14840,N_14915);
and UO_1044 (O_1044,N_14799,N_14947);
nand UO_1045 (O_1045,N_14830,N_14913);
xnor UO_1046 (O_1046,N_14977,N_14938);
nand UO_1047 (O_1047,N_14972,N_14845);
nand UO_1048 (O_1048,N_14799,N_14949);
and UO_1049 (O_1049,N_14885,N_14801);
nand UO_1050 (O_1050,N_14893,N_14909);
nor UO_1051 (O_1051,N_14951,N_14798);
nor UO_1052 (O_1052,N_14758,N_14976);
or UO_1053 (O_1053,N_14982,N_14768);
or UO_1054 (O_1054,N_14946,N_14801);
nor UO_1055 (O_1055,N_14974,N_14830);
nor UO_1056 (O_1056,N_14845,N_14962);
nor UO_1057 (O_1057,N_14892,N_14787);
xor UO_1058 (O_1058,N_14783,N_14850);
xor UO_1059 (O_1059,N_14765,N_14903);
nor UO_1060 (O_1060,N_14912,N_14891);
or UO_1061 (O_1061,N_14797,N_14808);
xor UO_1062 (O_1062,N_14909,N_14769);
or UO_1063 (O_1063,N_14985,N_14757);
and UO_1064 (O_1064,N_14777,N_14887);
nor UO_1065 (O_1065,N_14830,N_14847);
nand UO_1066 (O_1066,N_14827,N_14993);
xnor UO_1067 (O_1067,N_14926,N_14868);
and UO_1068 (O_1068,N_14820,N_14755);
nor UO_1069 (O_1069,N_14840,N_14891);
or UO_1070 (O_1070,N_14884,N_14828);
nor UO_1071 (O_1071,N_14901,N_14821);
or UO_1072 (O_1072,N_14989,N_14996);
or UO_1073 (O_1073,N_14818,N_14996);
or UO_1074 (O_1074,N_14807,N_14897);
or UO_1075 (O_1075,N_14853,N_14820);
xnor UO_1076 (O_1076,N_14802,N_14960);
or UO_1077 (O_1077,N_14929,N_14799);
nand UO_1078 (O_1078,N_14956,N_14871);
or UO_1079 (O_1079,N_14884,N_14767);
and UO_1080 (O_1080,N_14947,N_14928);
nand UO_1081 (O_1081,N_14924,N_14935);
and UO_1082 (O_1082,N_14970,N_14824);
xor UO_1083 (O_1083,N_14986,N_14867);
xnor UO_1084 (O_1084,N_14913,N_14960);
or UO_1085 (O_1085,N_14872,N_14806);
xnor UO_1086 (O_1086,N_14867,N_14996);
nand UO_1087 (O_1087,N_14925,N_14792);
nand UO_1088 (O_1088,N_14995,N_14836);
or UO_1089 (O_1089,N_14958,N_14880);
nor UO_1090 (O_1090,N_14824,N_14901);
or UO_1091 (O_1091,N_14858,N_14818);
or UO_1092 (O_1092,N_14973,N_14879);
xor UO_1093 (O_1093,N_14891,N_14821);
nand UO_1094 (O_1094,N_14959,N_14888);
and UO_1095 (O_1095,N_14874,N_14872);
and UO_1096 (O_1096,N_14864,N_14928);
or UO_1097 (O_1097,N_14767,N_14835);
nor UO_1098 (O_1098,N_14948,N_14777);
xnor UO_1099 (O_1099,N_14995,N_14936);
and UO_1100 (O_1100,N_14790,N_14910);
xnor UO_1101 (O_1101,N_14944,N_14757);
and UO_1102 (O_1102,N_14862,N_14842);
and UO_1103 (O_1103,N_14906,N_14886);
nor UO_1104 (O_1104,N_14887,N_14758);
xor UO_1105 (O_1105,N_14988,N_14989);
and UO_1106 (O_1106,N_14828,N_14812);
nor UO_1107 (O_1107,N_14769,N_14851);
and UO_1108 (O_1108,N_14919,N_14757);
or UO_1109 (O_1109,N_14841,N_14835);
nor UO_1110 (O_1110,N_14971,N_14770);
or UO_1111 (O_1111,N_14797,N_14966);
xnor UO_1112 (O_1112,N_14959,N_14751);
or UO_1113 (O_1113,N_14943,N_14903);
nand UO_1114 (O_1114,N_14893,N_14850);
or UO_1115 (O_1115,N_14785,N_14769);
nor UO_1116 (O_1116,N_14854,N_14855);
xnor UO_1117 (O_1117,N_14885,N_14876);
nor UO_1118 (O_1118,N_14962,N_14767);
nand UO_1119 (O_1119,N_14834,N_14949);
and UO_1120 (O_1120,N_14924,N_14949);
nor UO_1121 (O_1121,N_14998,N_14910);
and UO_1122 (O_1122,N_14993,N_14950);
nor UO_1123 (O_1123,N_14978,N_14891);
nor UO_1124 (O_1124,N_14954,N_14968);
xnor UO_1125 (O_1125,N_14821,N_14954);
and UO_1126 (O_1126,N_14771,N_14861);
nor UO_1127 (O_1127,N_14759,N_14785);
nand UO_1128 (O_1128,N_14919,N_14963);
nand UO_1129 (O_1129,N_14867,N_14869);
nand UO_1130 (O_1130,N_14894,N_14943);
and UO_1131 (O_1131,N_14993,N_14851);
nand UO_1132 (O_1132,N_14771,N_14815);
nor UO_1133 (O_1133,N_14920,N_14835);
and UO_1134 (O_1134,N_14828,N_14770);
or UO_1135 (O_1135,N_14895,N_14989);
or UO_1136 (O_1136,N_14982,N_14778);
nor UO_1137 (O_1137,N_14943,N_14986);
nand UO_1138 (O_1138,N_14820,N_14855);
nor UO_1139 (O_1139,N_14896,N_14856);
xnor UO_1140 (O_1140,N_14852,N_14883);
or UO_1141 (O_1141,N_14836,N_14787);
xor UO_1142 (O_1142,N_14967,N_14866);
or UO_1143 (O_1143,N_14934,N_14857);
nand UO_1144 (O_1144,N_14847,N_14894);
or UO_1145 (O_1145,N_14936,N_14960);
xnor UO_1146 (O_1146,N_14871,N_14990);
and UO_1147 (O_1147,N_14984,N_14846);
xor UO_1148 (O_1148,N_14809,N_14843);
nand UO_1149 (O_1149,N_14982,N_14837);
nor UO_1150 (O_1150,N_14846,N_14963);
or UO_1151 (O_1151,N_14959,N_14958);
or UO_1152 (O_1152,N_14857,N_14853);
nor UO_1153 (O_1153,N_14947,N_14826);
or UO_1154 (O_1154,N_14958,N_14761);
xor UO_1155 (O_1155,N_14882,N_14753);
nor UO_1156 (O_1156,N_14999,N_14959);
nand UO_1157 (O_1157,N_14876,N_14871);
or UO_1158 (O_1158,N_14872,N_14816);
and UO_1159 (O_1159,N_14949,N_14951);
nand UO_1160 (O_1160,N_14779,N_14852);
or UO_1161 (O_1161,N_14811,N_14961);
and UO_1162 (O_1162,N_14823,N_14998);
nor UO_1163 (O_1163,N_14942,N_14817);
or UO_1164 (O_1164,N_14944,N_14860);
and UO_1165 (O_1165,N_14813,N_14911);
nor UO_1166 (O_1166,N_14775,N_14852);
nand UO_1167 (O_1167,N_14993,N_14829);
nand UO_1168 (O_1168,N_14802,N_14894);
or UO_1169 (O_1169,N_14879,N_14822);
nor UO_1170 (O_1170,N_14875,N_14902);
and UO_1171 (O_1171,N_14845,N_14973);
and UO_1172 (O_1172,N_14911,N_14760);
or UO_1173 (O_1173,N_14967,N_14889);
nand UO_1174 (O_1174,N_14857,N_14821);
or UO_1175 (O_1175,N_14858,N_14946);
and UO_1176 (O_1176,N_14794,N_14994);
xnor UO_1177 (O_1177,N_14992,N_14808);
nand UO_1178 (O_1178,N_14861,N_14831);
nor UO_1179 (O_1179,N_14899,N_14883);
or UO_1180 (O_1180,N_14916,N_14992);
or UO_1181 (O_1181,N_14752,N_14846);
nor UO_1182 (O_1182,N_14880,N_14804);
nor UO_1183 (O_1183,N_14811,N_14926);
nand UO_1184 (O_1184,N_14875,N_14893);
and UO_1185 (O_1185,N_14799,N_14768);
or UO_1186 (O_1186,N_14914,N_14999);
xnor UO_1187 (O_1187,N_14814,N_14834);
and UO_1188 (O_1188,N_14922,N_14812);
and UO_1189 (O_1189,N_14978,N_14830);
nor UO_1190 (O_1190,N_14927,N_14823);
and UO_1191 (O_1191,N_14871,N_14867);
or UO_1192 (O_1192,N_14801,N_14772);
nand UO_1193 (O_1193,N_14958,N_14991);
and UO_1194 (O_1194,N_14814,N_14931);
xnor UO_1195 (O_1195,N_14886,N_14888);
xnor UO_1196 (O_1196,N_14769,N_14750);
or UO_1197 (O_1197,N_14776,N_14754);
nand UO_1198 (O_1198,N_14941,N_14919);
xor UO_1199 (O_1199,N_14752,N_14760);
nand UO_1200 (O_1200,N_14780,N_14938);
xnor UO_1201 (O_1201,N_14956,N_14896);
nor UO_1202 (O_1202,N_14794,N_14810);
xor UO_1203 (O_1203,N_14794,N_14829);
nand UO_1204 (O_1204,N_14956,N_14762);
nor UO_1205 (O_1205,N_14891,N_14761);
xor UO_1206 (O_1206,N_14766,N_14886);
and UO_1207 (O_1207,N_14900,N_14950);
and UO_1208 (O_1208,N_14811,N_14968);
xor UO_1209 (O_1209,N_14760,N_14896);
xnor UO_1210 (O_1210,N_14828,N_14835);
or UO_1211 (O_1211,N_14941,N_14900);
nand UO_1212 (O_1212,N_14949,N_14818);
xnor UO_1213 (O_1213,N_14975,N_14845);
nand UO_1214 (O_1214,N_14970,N_14929);
or UO_1215 (O_1215,N_14946,N_14753);
nand UO_1216 (O_1216,N_14960,N_14959);
nand UO_1217 (O_1217,N_14927,N_14940);
nand UO_1218 (O_1218,N_14912,N_14810);
xor UO_1219 (O_1219,N_14771,N_14976);
or UO_1220 (O_1220,N_14896,N_14928);
and UO_1221 (O_1221,N_14848,N_14780);
and UO_1222 (O_1222,N_14877,N_14795);
xor UO_1223 (O_1223,N_14903,N_14970);
or UO_1224 (O_1224,N_14954,N_14988);
xnor UO_1225 (O_1225,N_14808,N_14949);
nand UO_1226 (O_1226,N_14900,N_14886);
or UO_1227 (O_1227,N_14993,N_14875);
nand UO_1228 (O_1228,N_14752,N_14799);
nand UO_1229 (O_1229,N_14900,N_14882);
nand UO_1230 (O_1230,N_14781,N_14846);
or UO_1231 (O_1231,N_14995,N_14861);
nand UO_1232 (O_1232,N_14997,N_14851);
xnor UO_1233 (O_1233,N_14942,N_14759);
nand UO_1234 (O_1234,N_14821,N_14920);
or UO_1235 (O_1235,N_14762,N_14831);
xnor UO_1236 (O_1236,N_14960,N_14917);
and UO_1237 (O_1237,N_14876,N_14757);
xnor UO_1238 (O_1238,N_14861,N_14978);
and UO_1239 (O_1239,N_14869,N_14830);
nand UO_1240 (O_1240,N_14871,N_14907);
nand UO_1241 (O_1241,N_14873,N_14758);
nor UO_1242 (O_1242,N_14929,N_14770);
or UO_1243 (O_1243,N_14829,N_14798);
and UO_1244 (O_1244,N_14943,N_14785);
or UO_1245 (O_1245,N_14851,N_14902);
nand UO_1246 (O_1246,N_14979,N_14926);
xnor UO_1247 (O_1247,N_14988,N_14920);
nor UO_1248 (O_1248,N_14878,N_14847);
nand UO_1249 (O_1249,N_14759,N_14911);
nand UO_1250 (O_1250,N_14899,N_14913);
or UO_1251 (O_1251,N_14940,N_14888);
nand UO_1252 (O_1252,N_14959,N_14883);
xnor UO_1253 (O_1253,N_14922,N_14964);
nor UO_1254 (O_1254,N_14948,N_14958);
xor UO_1255 (O_1255,N_14851,N_14778);
xor UO_1256 (O_1256,N_14941,N_14993);
or UO_1257 (O_1257,N_14948,N_14919);
and UO_1258 (O_1258,N_14961,N_14877);
nand UO_1259 (O_1259,N_14957,N_14890);
and UO_1260 (O_1260,N_14872,N_14923);
or UO_1261 (O_1261,N_14785,N_14833);
or UO_1262 (O_1262,N_14905,N_14885);
or UO_1263 (O_1263,N_14859,N_14884);
and UO_1264 (O_1264,N_14822,N_14985);
nor UO_1265 (O_1265,N_14962,N_14830);
nand UO_1266 (O_1266,N_14889,N_14873);
nand UO_1267 (O_1267,N_14969,N_14926);
nand UO_1268 (O_1268,N_14815,N_14778);
nand UO_1269 (O_1269,N_14853,N_14880);
and UO_1270 (O_1270,N_14931,N_14915);
or UO_1271 (O_1271,N_14891,N_14759);
or UO_1272 (O_1272,N_14799,N_14986);
nor UO_1273 (O_1273,N_14877,N_14758);
or UO_1274 (O_1274,N_14977,N_14933);
and UO_1275 (O_1275,N_14890,N_14864);
and UO_1276 (O_1276,N_14845,N_14808);
and UO_1277 (O_1277,N_14795,N_14943);
xor UO_1278 (O_1278,N_14895,N_14828);
nand UO_1279 (O_1279,N_14888,N_14951);
or UO_1280 (O_1280,N_14992,N_14794);
nor UO_1281 (O_1281,N_14756,N_14870);
nand UO_1282 (O_1282,N_14812,N_14781);
nor UO_1283 (O_1283,N_14816,N_14878);
nor UO_1284 (O_1284,N_14762,N_14898);
nand UO_1285 (O_1285,N_14784,N_14991);
and UO_1286 (O_1286,N_14941,N_14792);
and UO_1287 (O_1287,N_14774,N_14768);
nor UO_1288 (O_1288,N_14896,N_14884);
nor UO_1289 (O_1289,N_14921,N_14947);
nand UO_1290 (O_1290,N_14888,N_14919);
and UO_1291 (O_1291,N_14884,N_14955);
or UO_1292 (O_1292,N_14847,N_14935);
and UO_1293 (O_1293,N_14884,N_14814);
nand UO_1294 (O_1294,N_14902,N_14835);
nor UO_1295 (O_1295,N_14920,N_14896);
and UO_1296 (O_1296,N_14833,N_14813);
nand UO_1297 (O_1297,N_14984,N_14992);
or UO_1298 (O_1298,N_14850,N_14808);
and UO_1299 (O_1299,N_14985,N_14902);
xor UO_1300 (O_1300,N_14887,N_14964);
and UO_1301 (O_1301,N_14970,N_14757);
nand UO_1302 (O_1302,N_14916,N_14812);
xor UO_1303 (O_1303,N_14765,N_14823);
nor UO_1304 (O_1304,N_14997,N_14861);
or UO_1305 (O_1305,N_14934,N_14849);
xnor UO_1306 (O_1306,N_14816,N_14765);
nor UO_1307 (O_1307,N_14837,N_14978);
nor UO_1308 (O_1308,N_14887,N_14914);
or UO_1309 (O_1309,N_14753,N_14847);
nand UO_1310 (O_1310,N_14896,N_14796);
and UO_1311 (O_1311,N_14838,N_14830);
nand UO_1312 (O_1312,N_14773,N_14996);
nor UO_1313 (O_1313,N_14807,N_14766);
xor UO_1314 (O_1314,N_14753,N_14892);
nor UO_1315 (O_1315,N_14845,N_14999);
or UO_1316 (O_1316,N_14962,N_14839);
xnor UO_1317 (O_1317,N_14871,N_14891);
or UO_1318 (O_1318,N_14894,N_14805);
nor UO_1319 (O_1319,N_14955,N_14925);
or UO_1320 (O_1320,N_14783,N_14982);
nand UO_1321 (O_1321,N_14790,N_14920);
and UO_1322 (O_1322,N_14902,N_14888);
or UO_1323 (O_1323,N_14889,N_14868);
or UO_1324 (O_1324,N_14994,N_14856);
nand UO_1325 (O_1325,N_14769,N_14888);
and UO_1326 (O_1326,N_14791,N_14860);
and UO_1327 (O_1327,N_14752,N_14811);
nand UO_1328 (O_1328,N_14771,N_14777);
nand UO_1329 (O_1329,N_14861,N_14873);
or UO_1330 (O_1330,N_14813,N_14996);
xnor UO_1331 (O_1331,N_14818,N_14753);
xor UO_1332 (O_1332,N_14796,N_14898);
or UO_1333 (O_1333,N_14869,N_14770);
nor UO_1334 (O_1334,N_14787,N_14820);
nor UO_1335 (O_1335,N_14754,N_14947);
or UO_1336 (O_1336,N_14810,N_14770);
nand UO_1337 (O_1337,N_14881,N_14972);
nor UO_1338 (O_1338,N_14877,N_14817);
nand UO_1339 (O_1339,N_14762,N_14903);
xnor UO_1340 (O_1340,N_14985,N_14794);
or UO_1341 (O_1341,N_14965,N_14867);
nand UO_1342 (O_1342,N_14934,N_14775);
and UO_1343 (O_1343,N_14937,N_14963);
nand UO_1344 (O_1344,N_14850,N_14895);
xnor UO_1345 (O_1345,N_14859,N_14927);
xnor UO_1346 (O_1346,N_14786,N_14933);
nor UO_1347 (O_1347,N_14892,N_14987);
and UO_1348 (O_1348,N_14813,N_14818);
or UO_1349 (O_1349,N_14970,N_14799);
and UO_1350 (O_1350,N_14967,N_14990);
nor UO_1351 (O_1351,N_14844,N_14842);
nand UO_1352 (O_1352,N_14883,N_14873);
nand UO_1353 (O_1353,N_14880,N_14786);
nand UO_1354 (O_1354,N_14801,N_14786);
xnor UO_1355 (O_1355,N_14883,N_14755);
nor UO_1356 (O_1356,N_14932,N_14923);
or UO_1357 (O_1357,N_14799,N_14988);
nor UO_1358 (O_1358,N_14934,N_14753);
xnor UO_1359 (O_1359,N_14857,N_14768);
and UO_1360 (O_1360,N_14869,N_14766);
xor UO_1361 (O_1361,N_14850,N_14993);
nor UO_1362 (O_1362,N_14867,N_14758);
and UO_1363 (O_1363,N_14974,N_14985);
nand UO_1364 (O_1364,N_14820,N_14893);
or UO_1365 (O_1365,N_14874,N_14963);
or UO_1366 (O_1366,N_14874,N_14812);
nand UO_1367 (O_1367,N_14935,N_14980);
nor UO_1368 (O_1368,N_14870,N_14985);
xor UO_1369 (O_1369,N_14854,N_14986);
or UO_1370 (O_1370,N_14853,N_14868);
xor UO_1371 (O_1371,N_14861,N_14803);
nor UO_1372 (O_1372,N_14842,N_14932);
nor UO_1373 (O_1373,N_14958,N_14899);
or UO_1374 (O_1374,N_14908,N_14795);
xor UO_1375 (O_1375,N_14769,N_14939);
nand UO_1376 (O_1376,N_14906,N_14832);
or UO_1377 (O_1377,N_14806,N_14791);
nor UO_1378 (O_1378,N_14906,N_14827);
nor UO_1379 (O_1379,N_14814,N_14933);
or UO_1380 (O_1380,N_14936,N_14898);
or UO_1381 (O_1381,N_14804,N_14952);
nor UO_1382 (O_1382,N_14852,N_14758);
and UO_1383 (O_1383,N_14996,N_14952);
nor UO_1384 (O_1384,N_14928,N_14754);
xor UO_1385 (O_1385,N_14939,N_14919);
and UO_1386 (O_1386,N_14767,N_14900);
and UO_1387 (O_1387,N_14919,N_14805);
nor UO_1388 (O_1388,N_14840,N_14773);
xor UO_1389 (O_1389,N_14844,N_14810);
nand UO_1390 (O_1390,N_14922,N_14885);
nand UO_1391 (O_1391,N_14853,N_14778);
and UO_1392 (O_1392,N_14895,N_14961);
xnor UO_1393 (O_1393,N_14982,N_14752);
and UO_1394 (O_1394,N_14806,N_14859);
nand UO_1395 (O_1395,N_14951,N_14788);
or UO_1396 (O_1396,N_14757,N_14794);
xor UO_1397 (O_1397,N_14996,N_14966);
or UO_1398 (O_1398,N_14865,N_14980);
nor UO_1399 (O_1399,N_14784,N_14792);
nor UO_1400 (O_1400,N_14920,N_14950);
or UO_1401 (O_1401,N_14799,N_14916);
xnor UO_1402 (O_1402,N_14800,N_14856);
and UO_1403 (O_1403,N_14932,N_14988);
or UO_1404 (O_1404,N_14768,N_14971);
xnor UO_1405 (O_1405,N_14825,N_14803);
nor UO_1406 (O_1406,N_14841,N_14753);
xnor UO_1407 (O_1407,N_14823,N_14766);
xor UO_1408 (O_1408,N_14943,N_14851);
and UO_1409 (O_1409,N_14989,N_14955);
nor UO_1410 (O_1410,N_14958,N_14881);
nand UO_1411 (O_1411,N_14930,N_14910);
nor UO_1412 (O_1412,N_14814,N_14996);
nor UO_1413 (O_1413,N_14914,N_14761);
xor UO_1414 (O_1414,N_14757,N_14925);
xnor UO_1415 (O_1415,N_14940,N_14906);
nor UO_1416 (O_1416,N_14848,N_14836);
xnor UO_1417 (O_1417,N_14861,N_14950);
xnor UO_1418 (O_1418,N_14878,N_14802);
and UO_1419 (O_1419,N_14902,N_14928);
and UO_1420 (O_1420,N_14948,N_14853);
xor UO_1421 (O_1421,N_14819,N_14761);
and UO_1422 (O_1422,N_14981,N_14911);
xor UO_1423 (O_1423,N_14855,N_14813);
nand UO_1424 (O_1424,N_14917,N_14848);
or UO_1425 (O_1425,N_14922,N_14921);
or UO_1426 (O_1426,N_14785,N_14912);
or UO_1427 (O_1427,N_14846,N_14934);
and UO_1428 (O_1428,N_14919,N_14859);
nand UO_1429 (O_1429,N_14804,N_14977);
or UO_1430 (O_1430,N_14901,N_14862);
nor UO_1431 (O_1431,N_14912,N_14837);
nor UO_1432 (O_1432,N_14869,N_14791);
xor UO_1433 (O_1433,N_14887,N_14918);
and UO_1434 (O_1434,N_14814,N_14981);
or UO_1435 (O_1435,N_14988,N_14868);
and UO_1436 (O_1436,N_14988,N_14832);
nand UO_1437 (O_1437,N_14948,N_14912);
nor UO_1438 (O_1438,N_14889,N_14792);
and UO_1439 (O_1439,N_14798,N_14986);
xnor UO_1440 (O_1440,N_14813,N_14937);
or UO_1441 (O_1441,N_14878,N_14954);
nand UO_1442 (O_1442,N_14963,N_14806);
or UO_1443 (O_1443,N_14780,N_14910);
xnor UO_1444 (O_1444,N_14765,N_14803);
nand UO_1445 (O_1445,N_14927,N_14963);
nor UO_1446 (O_1446,N_14964,N_14969);
and UO_1447 (O_1447,N_14905,N_14926);
nand UO_1448 (O_1448,N_14786,N_14871);
xnor UO_1449 (O_1449,N_14764,N_14806);
xor UO_1450 (O_1450,N_14900,N_14940);
nor UO_1451 (O_1451,N_14979,N_14869);
or UO_1452 (O_1452,N_14971,N_14781);
xnor UO_1453 (O_1453,N_14886,N_14774);
xor UO_1454 (O_1454,N_14979,N_14998);
or UO_1455 (O_1455,N_14928,N_14817);
xor UO_1456 (O_1456,N_14869,N_14896);
nand UO_1457 (O_1457,N_14998,N_14757);
xnor UO_1458 (O_1458,N_14838,N_14791);
nor UO_1459 (O_1459,N_14930,N_14995);
and UO_1460 (O_1460,N_14886,N_14943);
nor UO_1461 (O_1461,N_14767,N_14766);
nor UO_1462 (O_1462,N_14820,N_14872);
and UO_1463 (O_1463,N_14944,N_14845);
xnor UO_1464 (O_1464,N_14974,N_14869);
or UO_1465 (O_1465,N_14849,N_14890);
nor UO_1466 (O_1466,N_14844,N_14867);
nor UO_1467 (O_1467,N_14833,N_14806);
xor UO_1468 (O_1468,N_14827,N_14877);
nor UO_1469 (O_1469,N_14854,N_14827);
nand UO_1470 (O_1470,N_14766,N_14828);
xnor UO_1471 (O_1471,N_14759,N_14875);
xnor UO_1472 (O_1472,N_14850,N_14914);
xnor UO_1473 (O_1473,N_14841,N_14799);
xnor UO_1474 (O_1474,N_14961,N_14876);
or UO_1475 (O_1475,N_14954,N_14813);
nor UO_1476 (O_1476,N_14973,N_14818);
xor UO_1477 (O_1477,N_14952,N_14941);
xor UO_1478 (O_1478,N_14772,N_14834);
xor UO_1479 (O_1479,N_14809,N_14885);
nand UO_1480 (O_1480,N_14922,N_14983);
or UO_1481 (O_1481,N_14921,N_14756);
nand UO_1482 (O_1482,N_14780,N_14961);
nor UO_1483 (O_1483,N_14892,N_14836);
nor UO_1484 (O_1484,N_14813,N_14753);
and UO_1485 (O_1485,N_14751,N_14999);
or UO_1486 (O_1486,N_14970,N_14893);
nand UO_1487 (O_1487,N_14829,N_14755);
xor UO_1488 (O_1488,N_14872,N_14787);
or UO_1489 (O_1489,N_14753,N_14846);
xor UO_1490 (O_1490,N_14759,N_14803);
or UO_1491 (O_1491,N_14928,N_14829);
and UO_1492 (O_1492,N_14908,N_14845);
and UO_1493 (O_1493,N_14974,N_14978);
xor UO_1494 (O_1494,N_14790,N_14812);
and UO_1495 (O_1495,N_14933,N_14929);
and UO_1496 (O_1496,N_14979,N_14972);
nand UO_1497 (O_1497,N_14884,N_14865);
or UO_1498 (O_1498,N_14892,N_14772);
xor UO_1499 (O_1499,N_14982,N_14782);
xnor UO_1500 (O_1500,N_14823,N_14997);
nand UO_1501 (O_1501,N_14952,N_14937);
nand UO_1502 (O_1502,N_14828,N_14755);
nand UO_1503 (O_1503,N_14908,N_14877);
xnor UO_1504 (O_1504,N_14962,N_14859);
nand UO_1505 (O_1505,N_14941,N_14827);
or UO_1506 (O_1506,N_14838,N_14965);
nor UO_1507 (O_1507,N_14977,N_14828);
and UO_1508 (O_1508,N_14766,N_14778);
and UO_1509 (O_1509,N_14912,N_14929);
or UO_1510 (O_1510,N_14934,N_14975);
xor UO_1511 (O_1511,N_14912,N_14806);
xnor UO_1512 (O_1512,N_14897,N_14943);
nor UO_1513 (O_1513,N_14907,N_14947);
nand UO_1514 (O_1514,N_14781,N_14998);
and UO_1515 (O_1515,N_14799,N_14856);
and UO_1516 (O_1516,N_14951,N_14944);
xor UO_1517 (O_1517,N_14811,N_14928);
and UO_1518 (O_1518,N_14979,N_14906);
and UO_1519 (O_1519,N_14838,N_14783);
and UO_1520 (O_1520,N_14809,N_14923);
or UO_1521 (O_1521,N_14946,N_14938);
nor UO_1522 (O_1522,N_14914,N_14863);
nand UO_1523 (O_1523,N_14797,N_14817);
or UO_1524 (O_1524,N_14964,N_14754);
xor UO_1525 (O_1525,N_14983,N_14837);
and UO_1526 (O_1526,N_14909,N_14986);
and UO_1527 (O_1527,N_14861,N_14809);
xnor UO_1528 (O_1528,N_14809,N_14791);
nor UO_1529 (O_1529,N_14940,N_14879);
and UO_1530 (O_1530,N_14843,N_14872);
nand UO_1531 (O_1531,N_14835,N_14914);
and UO_1532 (O_1532,N_14965,N_14950);
nor UO_1533 (O_1533,N_14770,N_14816);
nor UO_1534 (O_1534,N_14752,N_14750);
nand UO_1535 (O_1535,N_14881,N_14966);
or UO_1536 (O_1536,N_14821,N_14964);
nor UO_1537 (O_1537,N_14897,N_14942);
and UO_1538 (O_1538,N_14771,N_14833);
nand UO_1539 (O_1539,N_14990,N_14783);
and UO_1540 (O_1540,N_14811,N_14890);
xnor UO_1541 (O_1541,N_14896,N_14925);
xnor UO_1542 (O_1542,N_14896,N_14894);
nand UO_1543 (O_1543,N_14963,N_14801);
and UO_1544 (O_1544,N_14908,N_14919);
and UO_1545 (O_1545,N_14767,N_14868);
xnor UO_1546 (O_1546,N_14763,N_14811);
xor UO_1547 (O_1547,N_14980,N_14903);
nand UO_1548 (O_1548,N_14990,N_14812);
nand UO_1549 (O_1549,N_14967,N_14807);
and UO_1550 (O_1550,N_14772,N_14787);
or UO_1551 (O_1551,N_14857,N_14960);
xor UO_1552 (O_1552,N_14762,N_14918);
nand UO_1553 (O_1553,N_14990,N_14823);
nand UO_1554 (O_1554,N_14771,N_14936);
nand UO_1555 (O_1555,N_14858,N_14765);
or UO_1556 (O_1556,N_14866,N_14970);
and UO_1557 (O_1557,N_14837,N_14914);
xnor UO_1558 (O_1558,N_14752,N_14958);
nand UO_1559 (O_1559,N_14785,N_14916);
nand UO_1560 (O_1560,N_14834,N_14864);
or UO_1561 (O_1561,N_14856,N_14955);
and UO_1562 (O_1562,N_14989,N_14901);
and UO_1563 (O_1563,N_14914,N_14753);
xnor UO_1564 (O_1564,N_14996,N_14918);
or UO_1565 (O_1565,N_14838,N_14788);
or UO_1566 (O_1566,N_14953,N_14806);
xnor UO_1567 (O_1567,N_14829,N_14864);
and UO_1568 (O_1568,N_14945,N_14891);
xnor UO_1569 (O_1569,N_14963,N_14913);
or UO_1570 (O_1570,N_14840,N_14759);
nand UO_1571 (O_1571,N_14923,N_14865);
and UO_1572 (O_1572,N_14781,N_14830);
nand UO_1573 (O_1573,N_14946,N_14829);
nand UO_1574 (O_1574,N_14791,N_14864);
xor UO_1575 (O_1575,N_14773,N_14860);
xor UO_1576 (O_1576,N_14942,N_14797);
xor UO_1577 (O_1577,N_14871,N_14765);
nand UO_1578 (O_1578,N_14970,N_14918);
xor UO_1579 (O_1579,N_14758,N_14813);
and UO_1580 (O_1580,N_14822,N_14754);
xor UO_1581 (O_1581,N_14945,N_14998);
nor UO_1582 (O_1582,N_14958,N_14796);
xor UO_1583 (O_1583,N_14812,N_14953);
or UO_1584 (O_1584,N_14885,N_14931);
xor UO_1585 (O_1585,N_14954,N_14950);
xor UO_1586 (O_1586,N_14848,N_14956);
nand UO_1587 (O_1587,N_14842,N_14870);
or UO_1588 (O_1588,N_14820,N_14941);
nor UO_1589 (O_1589,N_14892,N_14922);
nand UO_1590 (O_1590,N_14902,N_14943);
nand UO_1591 (O_1591,N_14991,N_14986);
nand UO_1592 (O_1592,N_14909,N_14943);
or UO_1593 (O_1593,N_14881,N_14954);
and UO_1594 (O_1594,N_14989,N_14850);
and UO_1595 (O_1595,N_14760,N_14934);
or UO_1596 (O_1596,N_14897,N_14765);
xnor UO_1597 (O_1597,N_14847,N_14766);
or UO_1598 (O_1598,N_14832,N_14915);
and UO_1599 (O_1599,N_14770,N_14765);
or UO_1600 (O_1600,N_14797,N_14963);
and UO_1601 (O_1601,N_14898,N_14835);
and UO_1602 (O_1602,N_14932,N_14960);
or UO_1603 (O_1603,N_14867,N_14985);
nor UO_1604 (O_1604,N_14982,N_14753);
xor UO_1605 (O_1605,N_14958,N_14910);
nand UO_1606 (O_1606,N_14912,N_14795);
nor UO_1607 (O_1607,N_14858,N_14999);
and UO_1608 (O_1608,N_14919,N_14774);
and UO_1609 (O_1609,N_14996,N_14963);
xnor UO_1610 (O_1610,N_14832,N_14962);
or UO_1611 (O_1611,N_14756,N_14955);
or UO_1612 (O_1612,N_14791,N_14769);
or UO_1613 (O_1613,N_14945,N_14964);
nand UO_1614 (O_1614,N_14839,N_14767);
or UO_1615 (O_1615,N_14765,N_14978);
xnor UO_1616 (O_1616,N_14782,N_14999);
and UO_1617 (O_1617,N_14823,N_14865);
or UO_1618 (O_1618,N_14922,N_14856);
nor UO_1619 (O_1619,N_14844,N_14881);
and UO_1620 (O_1620,N_14814,N_14927);
nor UO_1621 (O_1621,N_14996,N_14805);
nor UO_1622 (O_1622,N_14948,N_14868);
or UO_1623 (O_1623,N_14926,N_14830);
xor UO_1624 (O_1624,N_14819,N_14966);
nand UO_1625 (O_1625,N_14932,N_14955);
xor UO_1626 (O_1626,N_14968,N_14899);
nand UO_1627 (O_1627,N_14823,N_14770);
and UO_1628 (O_1628,N_14836,N_14951);
nor UO_1629 (O_1629,N_14772,N_14844);
nand UO_1630 (O_1630,N_14766,N_14953);
or UO_1631 (O_1631,N_14991,N_14946);
xor UO_1632 (O_1632,N_14840,N_14934);
and UO_1633 (O_1633,N_14953,N_14774);
xnor UO_1634 (O_1634,N_14928,N_14901);
or UO_1635 (O_1635,N_14847,N_14755);
xor UO_1636 (O_1636,N_14863,N_14838);
nand UO_1637 (O_1637,N_14930,N_14917);
nor UO_1638 (O_1638,N_14930,N_14941);
nand UO_1639 (O_1639,N_14857,N_14856);
nand UO_1640 (O_1640,N_14904,N_14870);
xor UO_1641 (O_1641,N_14846,N_14894);
nor UO_1642 (O_1642,N_14839,N_14782);
nand UO_1643 (O_1643,N_14806,N_14889);
xor UO_1644 (O_1644,N_14889,N_14776);
nand UO_1645 (O_1645,N_14912,N_14901);
nor UO_1646 (O_1646,N_14943,N_14970);
and UO_1647 (O_1647,N_14819,N_14924);
nor UO_1648 (O_1648,N_14770,N_14924);
and UO_1649 (O_1649,N_14926,N_14963);
nand UO_1650 (O_1650,N_14798,N_14766);
xor UO_1651 (O_1651,N_14826,N_14871);
or UO_1652 (O_1652,N_14753,N_14883);
nand UO_1653 (O_1653,N_14787,N_14891);
nor UO_1654 (O_1654,N_14753,N_14796);
nand UO_1655 (O_1655,N_14946,N_14847);
and UO_1656 (O_1656,N_14974,N_14871);
nand UO_1657 (O_1657,N_14764,N_14992);
or UO_1658 (O_1658,N_14881,N_14832);
nand UO_1659 (O_1659,N_14822,N_14794);
or UO_1660 (O_1660,N_14988,N_14891);
and UO_1661 (O_1661,N_14923,N_14797);
nand UO_1662 (O_1662,N_14751,N_14891);
xnor UO_1663 (O_1663,N_14878,N_14757);
xnor UO_1664 (O_1664,N_14805,N_14819);
and UO_1665 (O_1665,N_14867,N_14948);
xnor UO_1666 (O_1666,N_14855,N_14943);
and UO_1667 (O_1667,N_14804,N_14923);
nor UO_1668 (O_1668,N_14767,N_14880);
nor UO_1669 (O_1669,N_14797,N_14889);
nor UO_1670 (O_1670,N_14769,N_14925);
and UO_1671 (O_1671,N_14929,N_14890);
and UO_1672 (O_1672,N_14919,N_14860);
or UO_1673 (O_1673,N_14795,N_14757);
or UO_1674 (O_1674,N_14962,N_14939);
nor UO_1675 (O_1675,N_14853,N_14937);
xnor UO_1676 (O_1676,N_14832,N_14789);
or UO_1677 (O_1677,N_14980,N_14855);
or UO_1678 (O_1678,N_14845,N_14752);
xor UO_1679 (O_1679,N_14840,N_14752);
and UO_1680 (O_1680,N_14826,N_14842);
xor UO_1681 (O_1681,N_14792,N_14812);
nor UO_1682 (O_1682,N_14952,N_14800);
xnor UO_1683 (O_1683,N_14950,N_14769);
nand UO_1684 (O_1684,N_14931,N_14821);
nor UO_1685 (O_1685,N_14944,N_14875);
nor UO_1686 (O_1686,N_14971,N_14901);
and UO_1687 (O_1687,N_14877,N_14986);
nand UO_1688 (O_1688,N_14965,N_14985);
xnor UO_1689 (O_1689,N_14888,N_14757);
and UO_1690 (O_1690,N_14771,N_14918);
or UO_1691 (O_1691,N_14953,N_14968);
nor UO_1692 (O_1692,N_14879,N_14818);
xnor UO_1693 (O_1693,N_14777,N_14953);
nor UO_1694 (O_1694,N_14988,N_14928);
nor UO_1695 (O_1695,N_14772,N_14888);
nor UO_1696 (O_1696,N_14937,N_14847);
and UO_1697 (O_1697,N_14949,N_14875);
nor UO_1698 (O_1698,N_14955,N_14966);
and UO_1699 (O_1699,N_14991,N_14854);
or UO_1700 (O_1700,N_14991,N_14762);
or UO_1701 (O_1701,N_14872,N_14989);
and UO_1702 (O_1702,N_14931,N_14773);
xor UO_1703 (O_1703,N_14800,N_14849);
nand UO_1704 (O_1704,N_14872,N_14932);
or UO_1705 (O_1705,N_14920,N_14908);
nand UO_1706 (O_1706,N_14868,N_14905);
nor UO_1707 (O_1707,N_14773,N_14807);
nand UO_1708 (O_1708,N_14934,N_14892);
xnor UO_1709 (O_1709,N_14822,N_14946);
nand UO_1710 (O_1710,N_14941,N_14762);
and UO_1711 (O_1711,N_14914,N_14981);
xor UO_1712 (O_1712,N_14805,N_14875);
or UO_1713 (O_1713,N_14795,N_14874);
and UO_1714 (O_1714,N_14989,N_14776);
nand UO_1715 (O_1715,N_14939,N_14886);
or UO_1716 (O_1716,N_14965,N_14762);
and UO_1717 (O_1717,N_14903,N_14955);
and UO_1718 (O_1718,N_14810,N_14972);
or UO_1719 (O_1719,N_14779,N_14759);
or UO_1720 (O_1720,N_14777,N_14789);
or UO_1721 (O_1721,N_14993,N_14848);
and UO_1722 (O_1722,N_14843,N_14846);
and UO_1723 (O_1723,N_14751,N_14852);
and UO_1724 (O_1724,N_14762,N_14968);
xor UO_1725 (O_1725,N_14787,N_14841);
nand UO_1726 (O_1726,N_14998,N_14777);
nand UO_1727 (O_1727,N_14854,N_14814);
nand UO_1728 (O_1728,N_14906,N_14820);
and UO_1729 (O_1729,N_14846,N_14757);
xnor UO_1730 (O_1730,N_14941,N_14798);
nor UO_1731 (O_1731,N_14876,N_14770);
nand UO_1732 (O_1732,N_14799,N_14967);
or UO_1733 (O_1733,N_14816,N_14903);
and UO_1734 (O_1734,N_14863,N_14912);
and UO_1735 (O_1735,N_14775,N_14864);
and UO_1736 (O_1736,N_14868,N_14953);
nand UO_1737 (O_1737,N_14917,N_14763);
xor UO_1738 (O_1738,N_14920,N_14779);
nor UO_1739 (O_1739,N_14958,N_14916);
nand UO_1740 (O_1740,N_14876,N_14874);
or UO_1741 (O_1741,N_14818,N_14798);
or UO_1742 (O_1742,N_14814,N_14867);
nor UO_1743 (O_1743,N_14912,N_14990);
nor UO_1744 (O_1744,N_14912,N_14945);
and UO_1745 (O_1745,N_14952,N_14947);
and UO_1746 (O_1746,N_14979,N_14798);
nor UO_1747 (O_1747,N_14991,N_14900);
nand UO_1748 (O_1748,N_14959,N_14823);
or UO_1749 (O_1749,N_14898,N_14942);
nor UO_1750 (O_1750,N_14803,N_14752);
nand UO_1751 (O_1751,N_14855,N_14885);
nor UO_1752 (O_1752,N_14765,N_14896);
xor UO_1753 (O_1753,N_14772,N_14881);
and UO_1754 (O_1754,N_14830,N_14756);
xnor UO_1755 (O_1755,N_14808,N_14769);
and UO_1756 (O_1756,N_14786,N_14755);
and UO_1757 (O_1757,N_14936,N_14844);
nand UO_1758 (O_1758,N_14753,N_14754);
or UO_1759 (O_1759,N_14752,N_14916);
xor UO_1760 (O_1760,N_14940,N_14933);
nand UO_1761 (O_1761,N_14807,N_14971);
nor UO_1762 (O_1762,N_14791,N_14910);
and UO_1763 (O_1763,N_14860,N_14843);
nand UO_1764 (O_1764,N_14949,N_14993);
nand UO_1765 (O_1765,N_14900,N_14814);
nand UO_1766 (O_1766,N_14783,N_14860);
nand UO_1767 (O_1767,N_14886,N_14755);
and UO_1768 (O_1768,N_14873,N_14958);
nor UO_1769 (O_1769,N_14834,N_14792);
or UO_1770 (O_1770,N_14827,N_14952);
or UO_1771 (O_1771,N_14860,N_14885);
nand UO_1772 (O_1772,N_14862,N_14879);
nor UO_1773 (O_1773,N_14917,N_14815);
nor UO_1774 (O_1774,N_14756,N_14879);
xor UO_1775 (O_1775,N_14944,N_14853);
or UO_1776 (O_1776,N_14939,N_14910);
and UO_1777 (O_1777,N_14935,N_14763);
nor UO_1778 (O_1778,N_14955,N_14753);
xor UO_1779 (O_1779,N_14895,N_14981);
or UO_1780 (O_1780,N_14917,N_14835);
nand UO_1781 (O_1781,N_14973,N_14856);
or UO_1782 (O_1782,N_14878,N_14933);
nor UO_1783 (O_1783,N_14795,N_14984);
and UO_1784 (O_1784,N_14957,N_14968);
nand UO_1785 (O_1785,N_14799,N_14924);
nor UO_1786 (O_1786,N_14840,N_14897);
or UO_1787 (O_1787,N_14964,N_14794);
and UO_1788 (O_1788,N_14880,N_14763);
nand UO_1789 (O_1789,N_14828,N_14925);
and UO_1790 (O_1790,N_14843,N_14868);
or UO_1791 (O_1791,N_14860,N_14839);
nand UO_1792 (O_1792,N_14909,N_14903);
and UO_1793 (O_1793,N_14918,N_14932);
or UO_1794 (O_1794,N_14854,N_14857);
xor UO_1795 (O_1795,N_14926,N_14866);
or UO_1796 (O_1796,N_14844,N_14944);
xnor UO_1797 (O_1797,N_14972,N_14899);
nand UO_1798 (O_1798,N_14922,N_14779);
nor UO_1799 (O_1799,N_14778,N_14939);
nor UO_1800 (O_1800,N_14936,N_14879);
nor UO_1801 (O_1801,N_14888,N_14796);
nor UO_1802 (O_1802,N_14997,N_14838);
nor UO_1803 (O_1803,N_14846,N_14913);
xor UO_1804 (O_1804,N_14943,N_14961);
nor UO_1805 (O_1805,N_14911,N_14792);
nand UO_1806 (O_1806,N_14847,N_14873);
nand UO_1807 (O_1807,N_14936,N_14804);
nand UO_1808 (O_1808,N_14925,N_14796);
or UO_1809 (O_1809,N_14842,N_14974);
nor UO_1810 (O_1810,N_14880,N_14876);
nor UO_1811 (O_1811,N_14911,N_14974);
xnor UO_1812 (O_1812,N_14944,N_14839);
or UO_1813 (O_1813,N_14955,N_14950);
and UO_1814 (O_1814,N_14758,N_14967);
or UO_1815 (O_1815,N_14851,N_14832);
or UO_1816 (O_1816,N_14953,N_14907);
and UO_1817 (O_1817,N_14936,N_14820);
and UO_1818 (O_1818,N_14874,N_14802);
or UO_1819 (O_1819,N_14998,N_14857);
nand UO_1820 (O_1820,N_14912,N_14783);
xor UO_1821 (O_1821,N_14988,N_14752);
or UO_1822 (O_1822,N_14769,N_14968);
or UO_1823 (O_1823,N_14998,N_14773);
or UO_1824 (O_1824,N_14940,N_14949);
or UO_1825 (O_1825,N_14992,N_14772);
and UO_1826 (O_1826,N_14921,N_14810);
and UO_1827 (O_1827,N_14968,N_14980);
xor UO_1828 (O_1828,N_14899,N_14840);
xor UO_1829 (O_1829,N_14874,N_14792);
xor UO_1830 (O_1830,N_14769,N_14949);
or UO_1831 (O_1831,N_14941,N_14894);
and UO_1832 (O_1832,N_14752,N_14972);
or UO_1833 (O_1833,N_14905,N_14792);
xor UO_1834 (O_1834,N_14767,N_14933);
or UO_1835 (O_1835,N_14807,N_14935);
or UO_1836 (O_1836,N_14858,N_14780);
and UO_1837 (O_1837,N_14765,N_14881);
nor UO_1838 (O_1838,N_14844,N_14986);
nor UO_1839 (O_1839,N_14840,N_14911);
or UO_1840 (O_1840,N_14921,N_14981);
nor UO_1841 (O_1841,N_14862,N_14997);
nand UO_1842 (O_1842,N_14906,N_14761);
or UO_1843 (O_1843,N_14815,N_14945);
and UO_1844 (O_1844,N_14862,N_14908);
or UO_1845 (O_1845,N_14984,N_14762);
or UO_1846 (O_1846,N_14826,N_14803);
and UO_1847 (O_1847,N_14902,N_14780);
nor UO_1848 (O_1848,N_14924,N_14872);
nor UO_1849 (O_1849,N_14803,N_14754);
nand UO_1850 (O_1850,N_14912,N_14764);
nor UO_1851 (O_1851,N_14805,N_14971);
nand UO_1852 (O_1852,N_14931,N_14909);
xnor UO_1853 (O_1853,N_14807,N_14835);
nor UO_1854 (O_1854,N_14851,N_14812);
nand UO_1855 (O_1855,N_14906,N_14776);
nor UO_1856 (O_1856,N_14953,N_14934);
xnor UO_1857 (O_1857,N_14778,N_14962);
xnor UO_1858 (O_1858,N_14874,N_14875);
or UO_1859 (O_1859,N_14962,N_14927);
or UO_1860 (O_1860,N_14915,N_14800);
xor UO_1861 (O_1861,N_14984,N_14921);
nand UO_1862 (O_1862,N_14870,N_14908);
and UO_1863 (O_1863,N_14931,N_14788);
nor UO_1864 (O_1864,N_14909,N_14858);
or UO_1865 (O_1865,N_14837,N_14888);
or UO_1866 (O_1866,N_14835,N_14925);
xnor UO_1867 (O_1867,N_14784,N_14853);
or UO_1868 (O_1868,N_14769,N_14907);
nor UO_1869 (O_1869,N_14821,N_14773);
xnor UO_1870 (O_1870,N_14778,N_14953);
and UO_1871 (O_1871,N_14759,N_14952);
or UO_1872 (O_1872,N_14987,N_14770);
xor UO_1873 (O_1873,N_14805,N_14901);
nand UO_1874 (O_1874,N_14785,N_14874);
and UO_1875 (O_1875,N_14929,N_14804);
and UO_1876 (O_1876,N_14908,N_14952);
nor UO_1877 (O_1877,N_14779,N_14837);
xor UO_1878 (O_1878,N_14938,N_14754);
or UO_1879 (O_1879,N_14942,N_14982);
and UO_1880 (O_1880,N_14752,N_14860);
and UO_1881 (O_1881,N_14756,N_14918);
or UO_1882 (O_1882,N_14774,N_14967);
and UO_1883 (O_1883,N_14910,N_14795);
nor UO_1884 (O_1884,N_14908,N_14886);
nand UO_1885 (O_1885,N_14760,N_14968);
and UO_1886 (O_1886,N_14973,N_14998);
nand UO_1887 (O_1887,N_14795,N_14829);
nor UO_1888 (O_1888,N_14968,N_14869);
nor UO_1889 (O_1889,N_14882,N_14817);
or UO_1890 (O_1890,N_14892,N_14858);
xnor UO_1891 (O_1891,N_14803,N_14888);
xnor UO_1892 (O_1892,N_14891,N_14892);
xor UO_1893 (O_1893,N_14895,N_14893);
nand UO_1894 (O_1894,N_14815,N_14820);
nor UO_1895 (O_1895,N_14952,N_14794);
xor UO_1896 (O_1896,N_14812,N_14843);
or UO_1897 (O_1897,N_14903,N_14872);
and UO_1898 (O_1898,N_14816,N_14901);
nor UO_1899 (O_1899,N_14898,N_14938);
nor UO_1900 (O_1900,N_14948,N_14800);
or UO_1901 (O_1901,N_14966,N_14927);
nor UO_1902 (O_1902,N_14928,N_14884);
and UO_1903 (O_1903,N_14972,N_14908);
and UO_1904 (O_1904,N_14940,N_14867);
nor UO_1905 (O_1905,N_14859,N_14846);
xor UO_1906 (O_1906,N_14941,N_14832);
nor UO_1907 (O_1907,N_14851,N_14876);
xor UO_1908 (O_1908,N_14848,N_14762);
or UO_1909 (O_1909,N_14792,N_14751);
nor UO_1910 (O_1910,N_14996,N_14776);
xnor UO_1911 (O_1911,N_14980,N_14969);
nor UO_1912 (O_1912,N_14796,N_14818);
nand UO_1913 (O_1913,N_14985,N_14866);
nand UO_1914 (O_1914,N_14950,N_14791);
and UO_1915 (O_1915,N_14851,N_14967);
nor UO_1916 (O_1916,N_14869,N_14865);
nor UO_1917 (O_1917,N_14953,N_14841);
nor UO_1918 (O_1918,N_14934,N_14754);
nor UO_1919 (O_1919,N_14881,N_14828);
or UO_1920 (O_1920,N_14885,N_14901);
or UO_1921 (O_1921,N_14932,N_14852);
nor UO_1922 (O_1922,N_14830,N_14903);
and UO_1923 (O_1923,N_14839,N_14941);
or UO_1924 (O_1924,N_14938,N_14903);
or UO_1925 (O_1925,N_14791,N_14929);
nor UO_1926 (O_1926,N_14881,N_14810);
and UO_1927 (O_1927,N_14995,N_14760);
or UO_1928 (O_1928,N_14845,N_14949);
or UO_1929 (O_1929,N_14981,N_14778);
nand UO_1930 (O_1930,N_14908,N_14969);
xnor UO_1931 (O_1931,N_14913,N_14833);
and UO_1932 (O_1932,N_14979,N_14921);
xor UO_1933 (O_1933,N_14962,N_14914);
or UO_1934 (O_1934,N_14947,N_14810);
nor UO_1935 (O_1935,N_14940,N_14881);
nand UO_1936 (O_1936,N_14862,N_14860);
nand UO_1937 (O_1937,N_14972,N_14812);
nand UO_1938 (O_1938,N_14864,N_14951);
or UO_1939 (O_1939,N_14775,N_14771);
nor UO_1940 (O_1940,N_14771,N_14938);
xor UO_1941 (O_1941,N_14754,N_14933);
and UO_1942 (O_1942,N_14807,N_14946);
or UO_1943 (O_1943,N_14943,N_14862);
nand UO_1944 (O_1944,N_14974,N_14888);
or UO_1945 (O_1945,N_14994,N_14821);
nor UO_1946 (O_1946,N_14992,N_14783);
or UO_1947 (O_1947,N_14846,N_14831);
nor UO_1948 (O_1948,N_14817,N_14998);
nor UO_1949 (O_1949,N_14995,N_14860);
and UO_1950 (O_1950,N_14916,N_14946);
or UO_1951 (O_1951,N_14857,N_14898);
nor UO_1952 (O_1952,N_14817,N_14927);
xor UO_1953 (O_1953,N_14863,N_14761);
nor UO_1954 (O_1954,N_14920,N_14840);
nand UO_1955 (O_1955,N_14774,N_14957);
or UO_1956 (O_1956,N_14961,N_14886);
or UO_1957 (O_1957,N_14942,N_14988);
or UO_1958 (O_1958,N_14826,N_14892);
xor UO_1959 (O_1959,N_14852,N_14986);
or UO_1960 (O_1960,N_14754,N_14988);
or UO_1961 (O_1961,N_14897,N_14758);
and UO_1962 (O_1962,N_14977,N_14862);
nand UO_1963 (O_1963,N_14961,N_14995);
and UO_1964 (O_1964,N_14841,N_14792);
or UO_1965 (O_1965,N_14983,N_14955);
xnor UO_1966 (O_1966,N_14907,N_14887);
nand UO_1967 (O_1967,N_14761,N_14949);
nand UO_1968 (O_1968,N_14901,N_14997);
or UO_1969 (O_1969,N_14941,N_14947);
and UO_1970 (O_1970,N_14929,N_14943);
xor UO_1971 (O_1971,N_14905,N_14933);
xor UO_1972 (O_1972,N_14970,N_14850);
nand UO_1973 (O_1973,N_14896,N_14901);
or UO_1974 (O_1974,N_14765,N_14953);
and UO_1975 (O_1975,N_14751,N_14814);
nor UO_1976 (O_1976,N_14825,N_14761);
nand UO_1977 (O_1977,N_14866,N_14804);
nand UO_1978 (O_1978,N_14882,N_14828);
or UO_1979 (O_1979,N_14842,N_14796);
nor UO_1980 (O_1980,N_14860,N_14881);
and UO_1981 (O_1981,N_14824,N_14921);
xnor UO_1982 (O_1982,N_14796,N_14996);
nand UO_1983 (O_1983,N_14866,N_14796);
and UO_1984 (O_1984,N_14780,N_14817);
and UO_1985 (O_1985,N_14961,N_14852);
and UO_1986 (O_1986,N_14927,N_14758);
xnor UO_1987 (O_1987,N_14922,N_14972);
and UO_1988 (O_1988,N_14831,N_14856);
nor UO_1989 (O_1989,N_14760,N_14836);
xnor UO_1990 (O_1990,N_14944,N_14807);
xnor UO_1991 (O_1991,N_14985,N_14959);
and UO_1992 (O_1992,N_14802,N_14778);
and UO_1993 (O_1993,N_14815,N_14753);
or UO_1994 (O_1994,N_14881,N_14911);
or UO_1995 (O_1995,N_14784,N_14781);
nand UO_1996 (O_1996,N_14802,N_14861);
nor UO_1997 (O_1997,N_14750,N_14844);
nand UO_1998 (O_1998,N_14879,N_14898);
and UO_1999 (O_1999,N_14794,N_14978);
endmodule