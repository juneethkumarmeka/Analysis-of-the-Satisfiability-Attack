module basic_500_3000_500_50_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_123,In_52);
and U1 (N_1,In_18,In_165);
nor U2 (N_2,In_88,In_480);
nand U3 (N_3,In_285,In_348);
or U4 (N_4,In_99,In_58);
and U5 (N_5,In_73,In_316);
or U6 (N_6,In_335,In_320);
or U7 (N_7,In_353,In_27);
and U8 (N_8,In_309,In_15);
and U9 (N_9,In_93,In_278);
nand U10 (N_10,In_262,In_171);
and U11 (N_11,In_45,In_478);
and U12 (N_12,In_307,In_382);
nor U13 (N_13,In_232,In_421);
nor U14 (N_14,In_223,In_358);
xor U15 (N_15,In_184,In_94);
nor U16 (N_16,In_4,In_314);
or U17 (N_17,In_56,In_35);
nand U18 (N_18,In_22,In_218);
nor U19 (N_19,In_60,In_362);
or U20 (N_20,In_124,In_202);
nand U21 (N_21,In_279,In_192);
nor U22 (N_22,In_283,In_393);
and U23 (N_23,In_406,In_433);
or U24 (N_24,In_152,In_38);
nor U25 (N_25,In_288,In_33);
nor U26 (N_26,In_310,In_442);
and U27 (N_27,In_221,In_380);
nor U28 (N_28,In_264,In_384);
and U29 (N_29,In_44,In_343);
nor U30 (N_30,In_456,In_313);
xor U31 (N_31,In_117,In_249);
nand U32 (N_32,In_397,In_14);
or U33 (N_33,In_426,In_95);
nand U34 (N_34,In_304,In_120);
and U35 (N_35,In_39,In_328);
or U36 (N_36,In_332,In_427);
or U37 (N_37,In_55,In_143);
nor U38 (N_38,In_220,In_338);
xnor U39 (N_39,In_319,In_377);
nand U40 (N_40,In_325,In_114);
nor U41 (N_41,In_365,In_371);
or U42 (N_42,In_403,In_386);
nand U43 (N_43,In_451,In_102);
xnor U44 (N_44,In_241,In_373);
nor U45 (N_45,In_396,In_20);
nand U46 (N_46,In_398,In_460);
nor U47 (N_47,In_179,In_199);
xor U48 (N_48,In_477,In_248);
or U49 (N_49,In_11,In_441);
nand U50 (N_50,In_231,In_315);
and U51 (N_51,In_96,In_49);
xor U52 (N_52,In_312,In_268);
xor U53 (N_53,In_208,In_467);
nor U54 (N_54,In_475,In_493);
nor U55 (N_55,In_369,In_90);
nand U56 (N_56,In_274,In_244);
nor U57 (N_57,In_470,In_383);
and U58 (N_58,In_200,In_79);
or U59 (N_59,In_280,In_352);
nor U60 (N_60,In_207,In_8);
nand U61 (N_61,In_404,In_156);
nand U62 (N_62,In_381,In_211);
and U63 (N_63,In_78,In_306);
and U64 (N_64,In_144,N_57);
and U65 (N_65,In_28,In_337);
nor U66 (N_66,In_121,In_9);
and U67 (N_67,In_215,In_254);
nand U68 (N_68,In_158,In_154);
and U69 (N_69,In_497,In_284);
nor U70 (N_70,In_75,In_111);
nand U71 (N_71,In_351,In_130);
and U72 (N_72,In_445,In_340);
nand U73 (N_73,In_226,In_370);
or U74 (N_74,In_360,In_455);
nand U75 (N_75,In_435,N_35);
nor U76 (N_76,In_177,N_25);
nor U77 (N_77,In_203,In_62);
and U78 (N_78,In_481,In_63);
or U79 (N_79,In_206,In_449);
xnor U80 (N_80,N_38,In_260);
nor U81 (N_81,N_10,In_84);
and U82 (N_82,In_374,In_141);
or U83 (N_83,N_7,In_212);
nand U84 (N_84,In_23,N_4);
nor U85 (N_85,In_105,In_482);
nand U86 (N_86,In_0,In_263);
or U87 (N_87,In_305,In_350);
nand U88 (N_88,In_333,In_188);
nand U89 (N_89,In_321,N_14);
or U90 (N_90,In_401,In_399);
xnor U91 (N_91,In_331,In_48);
or U92 (N_92,In_185,N_51);
xnor U93 (N_93,In_378,In_245);
xnor U94 (N_94,N_36,In_483);
nor U95 (N_95,In_425,In_363);
or U96 (N_96,In_295,In_109);
xnor U97 (N_97,In_388,In_339);
nor U98 (N_98,In_224,In_228);
or U99 (N_99,In_34,In_159);
or U100 (N_100,In_489,In_443);
nand U101 (N_101,In_222,In_466);
nor U102 (N_102,In_308,In_303);
and U103 (N_103,In_178,In_347);
nor U104 (N_104,In_133,In_327);
or U105 (N_105,In_457,In_420);
nand U106 (N_106,N_9,In_468);
and U107 (N_107,In_19,In_160);
nand U108 (N_108,In_6,In_10);
nand U109 (N_109,In_1,In_108);
and U110 (N_110,In_82,N_52);
or U111 (N_111,In_235,In_80);
nand U112 (N_112,In_463,In_415);
nor U113 (N_113,In_499,In_118);
nand U114 (N_114,In_453,N_30);
nor U115 (N_115,In_436,In_31);
and U116 (N_116,In_336,In_70);
nor U117 (N_117,In_67,N_26);
nand U118 (N_118,In_287,In_491);
nand U119 (N_119,In_193,In_42);
or U120 (N_120,N_19,In_155);
or U121 (N_121,N_62,In_204);
and U122 (N_122,In_92,In_417);
or U123 (N_123,In_418,N_1);
and U124 (N_124,In_100,In_276);
nor U125 (N_125,In_391,In_153);
and U126 (N_126,N_42,In_345);
nand U127 (N_127,In_234,In_251);
nor U128 (N_128,N_15,In_85);
nand U129 (N_129,In_140,N_17);
nand U130 (N_130,N_61,In_301);
nand U131 (N_131,In_135,In_157);
or U132 (N_132,In_190,In_71);
nand U133 (N_133,In_492,In_7);
or U134 (N_134,In_488,In_172);
nand U135 (N_135,N_72,In_299);
and U136 (N_136,In_17,In_410);
nand U137 (N_137,In_269,N_83);
and U138 (N_138,In_237,In_324);
nand U139 (N_139,N_99,In_405);
nor U140 (N_140,In_407,N_5);
xnor U141 (N_141,In_447,In_173);
or U142 (N_142,In_496,In_372);
nor U143 (N_143,In_261,N_49);
nand U144 (N_144,In_122,In_484);
nand U145 (N_145,In_246,In_69);
and U146 (N_146,N_81,In_13);
and U147 (N_147,In_424,In_334);
nor U148 (N_148,In_103,In_472);
xor U149 (N_149,In_30,N_106);
and U150 (N_150,N_27,N_48);
nand U151 (N_151,In_209,In_474);
or U152 (N_152,In_476,In_469);
nor U153 (N_153,N_8,N_117);
nor U154 (N_154,In_87,In_494);
nor U155 (N_155,N_103,N_43);
and U156 (N_156,In_430,N_89);
or U157 (N_157,In_116,In_342);
nor U158 (N_158,In_180,In_253);
nand U159 (N_159,In_162,In_230);
nor U160 (N_160,In_290,In_250);
and U161 (N_161,In_164,In_240);
or U162 (N_162,N_70,In_317);
nor U163 (N_163,N_53,N_114);
and U164 (N_164,N_37,N_46);
and U165 (N_165,In_458,In_289);
or U166 (N_166,In_361,In_329);
or U167 (N_167,In_68,In_486);
or U168 (N_168,In_349,N_31);
nor U169 (N_169,In_225,In_359);
nand U170 (N_170,N_88,N_3);
and U171 (N_171,N_108,N_40);
or U172 (N_172,N_24,In_213);
and U173 (N_173,In_46,In_473);
nor U174 (N_174,In_217,N_13);
and U175 (N_175,N_23,In_367);
and U176 (N_176,In_129,In_36);
xor U177 (N_177,In_138,N_22);
nor U178 (N_178,In_330,In_166);
and U179 (N_179,In_110,In_270);
nor U180 (N_180,In_267,N_126);
or U181 (N_181,N_163,In_292);
and U182 (N_182,In_125,N_148);
nor U183 (N_183,In_148,N_110);
and U184 (N_184,N_142,N_116);
or U185 (N_185,N_125,In_196);
xor U186 (N_186,N_16,N_120);
and U187 (N_187,In_265,N_45);
nor U188 (N_188,In_65,N_135);
nand U189 (N_189,In_302,N_162);
nor U190 (N_190,N_98,N_59);
or U191 (N_191,In_216,N_85);
nand U192 (N_192,In_252,In_387);
xnor U193 (N_193,N_155,In_64);
nand U194 (N_194,In_400,In_437);
or U195 (N_195,In_411,In_408);
nor U196 (N_196,In_356,N_111);
nor U197 (N_197,In_89,In_236);
nor U198 (N_198,In_149,N_122);
nand U199 (N_199,N_56,In_368);
nand U200 (N_200,In_448,In_139);
nor U201 (N_201,N_96,In_97);
and U202 (N_202,In_182,In_136);
nand U203 (N_203,In_275,N_86);
and U204 (N_204,In_194,In_311);
and U205 (N_205,N_164,In_454);
nor U206 (N_206,N_33,N_146);
or U207 (N_207,N_28,N_178);
and U208 (N_208,N_118,In_459);
xnor U209 (N_209,N_84,In_197);
nor U210 (N_210,N_136,N_158);
nand U211 (N_211,N_71,In_465);
and U212 (N_212,In_169,In_72);
xor U213 (N_213,In_247,N_140);
nor U214 (N_214,In_440,In_47);
and U215 (N_215,In_32,In_357);
and U216 (N_216,In_341,In_239);
xnor U217 (N_217,N_138,In_490);
and U218 (N_218,In_323,N_141);
or U219 (N_219,N_93,N_100);
or U220 (N_220,In_344,In_375);
and U221 (N_221,In_40,In_385);
xor U222 (N_222,In_438,In_366);
xnor U223 (N_223,N_60,In_498);
nand U224 (N_224,N_119,In_189);
and U225 (N_225,In_66,N_18);
and U226 (N_226,N_161,In_205);
and U227 (N_227,N_172,In_434);
or U228 (N_228,N_133,N_2);
nor U229 (N_229,N_54,N_115);
nand U230 (N_230,N_174,In_322);
and U231 (N_231,In_146,In_346);
or U232 (N_232,N_166,In_495);
or U233 (N_233,In_266,In_214);
nand U234 (N_234,N_68,N_145);
xnor U235 (N_235,N_41,In_57);
nor U236 (N_236,In_175,In_429);
xor U237 (N_237,N_109,In_198);
nor U238 (N_238,In_127,In_227);
and U239 (N_239,In_462,In_53);
nand U240 (N_240,N_234,N_179);
nand U241 (N_241,In_113,N_6);
nor U242 (N_242,In_422,In_29);
nor U243 (N_243,In_170,In_163);
nor U244 (N_244,In_176,N_206);
or U245 (N_245,N_193,In_439);
nor U246 (N_246,N_80,In_150);
nor U247 (N_247,N_123,In_412);
and U248 (N_248,N_149,In_416);
and U249 (N_249,In_271,N_101);
and U250 (N_250,In_392,N_184);
nand U251 (N_251,In_296,In_168);
xor U252 (N_252,N_227,N_104);
and U253 (N_253,N_213,In_101);
nand U254 (N_254,In_233,N_230);
nor U255 (N_255,In_258,In_147);
and U256 (N_256,In_259,N_233);
nor U257 (N_257,In_376,N_130);
or U258 (N_258,In_77,In_293);
nor U259 (N_259,N_90,In_137);
nand U260 (N_260,N_121,In_119);
and U261 (N_261,In_485,In_54);
nor U262 (N_262,N_127,N_55);
or U263 (N_263,N_165,In_255);
or U264 (N_264,In_43,N_79);
nor U265 (N_265,In_419,N_204);
and U266 (N_266,N_207,N_34);
nor U267 (N_267,In_59,N_92);
and U268 (N_268,In_151,N_195);
nor U269 (N_269,N_105,In_61);
nand U270 (N_270,In_402,N_223);
nand U271 (N_271,In_195,N_44);
nand U272 (N_272,N_194,N_0);
nor U273 (N_273,N_63,N_58);
or U274 (N_274,In_106,N_94);
nor U275 (N_275,N_168,In_16);
or U276 (N_276,In_187,N_232);
and U277 (N_277,N_107,In_76);
nor U278 (N_278,In_98,In_142);
xnor U279 (N_279,N_78,N_159);
or U280 (N_280,In_134,N_160);
nand U281 (N_281,N_185,N_50);
and U282 (N_282,In_115,N_186);
or U283 (N_283,N_102,N_228);
xnor U284 (N_284,N_189,In_326);
and U285 (N_285,N_73,N_69);
nand U286 (N_286,In_395,N_231);
or U287 (N_287,In_256,In_25);
or U288 (N_288,In_242,N_180);
or U289 (N_289,N_113,In_291);
nor U290 (N_290,N_144,In_2);
or U291 (N_291,N_167,In_452);
nand U292 (N_292,N_217,N_188);
nor U293 (N_293,N_29,N_202);
nand U294 (N_294,N_154,N_239);
and U295 (N_295,N_238,In_300);
nand U296 (N_296,N_150,In_431);
or U297 (N_297,N_182,N_124);
nand U298 (N_298,In_277,N_47);
xor U299 (N_299,In_297,In_229);
or U300 (N_300,N_97,N_219);
nor U301 (N_301,N_128,N_151);
nand U302 (N_302,N_240,N_143);
xor U303 (N_303,In_354,N_245);
nand U304 (N_304,In_281,N_74);
or U305 (N_305,In_379,N_290);
nor U306 (N_306,N_281,In_446);
nand U307 (N_307,N_226,N_269);
or U308 (N_308,In_74,N_267);
nand U309 (N_309,N_205,N_147);
and U310 (N_310,N_152,In_364);
and U311 (N_311,In_191,In_479);
and U312 (N_312,In_37,In_12);
or U313 (N_313,N_279,In_128);
nor U314 (N_314,In_243,In_81);
nor U315 (N_315,N_255,N_77);
and U316 (N_316,In_26,N_285);
nand U317 (N_317,In_273,N_224);
or U318 (N_318,N_278,N_236);
or U319 (N_319,In_414,N_289);
and U320 (N_320,In_272,N_218);
or U321 (N_321,In_201,N_212);
or U322 (N_322,N_32,In_461);
nor U323 (N_323,In_83,N_192);
nand U324 (N_324,N_216,N_173);
nand U325 (N_325,In_51,In_219);
nand U326 (N_326,N_265,N_262);
nand U327 (N_327,N_258,N_20);
and U328 (N_328,In_282,In_257);
or U329 (N_329,N_131,In_450);
or U330 (N_330,N_237,N_264);
xor U331 (N_331,N_266,In_181);
and U332 (N_332,N_137,N_273);
or U333 (N_333,N_67,In_428);
or U334 (N_334,In_107,N_291);
and U335 (N_335,N_246,N_211);
or U336 (N_336,N_251,N_39);
or U337 (N_337,In_210,N_76);
nor U338 (N_338,N_12,In_174);
nand U339 (N_339,N_87,N_260);
and U340 (N_340,N_177,N_210);
and U341 (N_341,In_471,In_390);
nor U342 (N_342,N_214,N_156);
nand U343 (N_343,In_3,N_271);
xnor U344 (N_344,N_277,N_229);
xor U345 (N_345,N_298,N_201);
nor U346 (N_346,N_181,In_487);
xor U347 (N_347,N_175,In_444);
nor U348 (N_348,N_241,In_41);
or U349 (N_349,N_209,N_295);
and U350 (N_350,N_75,N_199);
nor U351 (N_351,In_423,N_243);
or U352 (N_352,N_242,In_238);
or U353 (N_353,In_413,In_298);
nand U354 (N_354,N_197,N_221);
and U355 (N_355,In_186,N_191);
xor U356 (N_356,N_247,N_257);
or U357 (N_357,N_284,N_275);
nand U358 (N_358,N_190,In_389);
and U359 (N_359,In_132,N_268);
or U360 (N_360,N_139,N_337);
nor U361 (N_361,N_319,N_296);
nand U362 (N_362,N_95,N_318);
xor U363 (N_363,N_333,N_235);
and U364 (N_364,N_312,N_309);
and U365 (N_365,In_91,N_344);
and U366 (N_366,In_112,N_331);
xnor U367 (N_367,N_305,N_326);
and U368 (N_368,In_294,N_263);
nand U369 (N_369,N_346,N_329);
nand U370 (N_370,N_261,N_338);
xor U371 (N_371,N_339,In_104);
xor U372 (N_372,N_297,N_350);
and U373 (N_373,N_65,N_82);
nor U374 (N_374,N_208,In_432);
or U375 (N_375,N_313,N_287);
or U376 (N_376,N_358,N_248);
xor U377 (N_377,N_276,N_153);
and U378 (N_378,N_335,N_336);
and U379 (N_379,N_293,N_215);
nor U380 (N_380,In_318,N_355);
and U381 (N_381,In_50,N_129);
nor U382 (N_382,N_256,In_286);
nand U383 (N_383,N_316,N_307);
and U384 (N_384,N_198,N_314);
nand U385 (N_385,N_203,N_171);
xnor U386 (N_386,N_308,N_222);
nor U387 (N_387,N_270,N_157);
nand U388 (N_388,In_86,N_310);
and U389 (N_389,N_340,N_170);
nand U390 (N_390,N_286,N_252);
or U391 (N_391,N_21,N_323);
nand U392 (N_392,N_304,N_283);
nor U393 (N_393,In_24,N_183);
or U394 (N_394,In_355,N_306);
and U395 (N_395,N_64,In_126);
nand U396 (N_396,N_352,N_169);
or U397 (N_397,In_409,N_225);
and U398 (N_398,N_348,N_317);
and U399 (N_399,N_176,N_280);
nor U400 (N_400,N_332,N_343);
nor U401 (N_401,N_300,N_341);
or U402 (N_402,N_66,N_349);
nand U403 (N_403,N_347,N_134);
and U404 (N_404,N_299,In_394);
and U405 (N_405,N_249,N_334);
nand U406 (N_406,N_354,N_325);
and U407 (N_407,N_357,N_345);
or U408 (N_408,N_259,In_5);
nand U409 (N_409,N_328,N_327);
or U410 (N_410,In_183,N_294);
and U411 (N_411,N_272,N_91);
nor U412 (N_412,N_311,N_244);
xnor U413 (N_413,In_161,N_112);
nand U414 (N_414,N_359,N_200);
nor U415 (N_415,In_145,N_288);
or U416 (N_416,In_131,N_301);
nand U417 (N_417,N_196,N_220);
nor U418 (N_418,In_21,N_356);
or U419 (N_419,N_321,N_330);
xnor U420 (N_420,N_187,N_370);
nand U421 (N_421,N_389,N_418);
and U422 (N_422,N_374,N_397);
nand U423 (N_423,N_368,N_417);
nor U424 (N_424,N_383,N_363);
or U425 (N_425,N_360,N_342);
and U426 (N_426,N_403,N_353);
nor U427 (N_427,N_379,N_386);
or U428 (N_428,N_398,N_292);
nor U429 (N_429,N_315,N_324);
nor U430 (N_430,N_351,N_419);
nor U431 (N_431,N_378,N_392);
nor U432 (N_432,N_410,N_384);
or U433 (N_433,N_380,N_416);
or U434 (N_434,N_399,N_302);
and U435 (N_435,N_409,N_250);
and U436 (N_436,N_412,N_254);
xor U437 (N_437,N_253,N_362);
or U438 (N_438,N_393,N_365);
and U439 (N_439,N_413,N_396);
or U440 (N_440,N_303,N_372);
or U441 (N_441,N_11,N_369);
nand U442 (N_442,N_376,N_401);
or U443 (N_443,N_364,N_400);
xnor U444 (N_444,N_361,N_394);
and U445 (N_445,N_274,N_391);
xor U446 (N_446,N_406,N_373);
nand U447 (N_447,In_167,N_387);
and U448 (N_448,N_382,N_377);
or U449 (N_449,N_385,N_402);
nand U450 (N_450,N_415,N_371);
nor U451 (N_451,N_411,N_367);
nor U452 (N_452,N_407,N_320);
and U453 (N_453,N_388,N_390);
or U454 (N_454,N_408,N_322);
nor U455 (N_455,N_405,N_381);
nand U456 (N_456,N_414,N_132);
nand U457 (N_457,N_375,In_464);
nor U458 (N_458,N_395,N_404);
and U459 (N_459,N_366,N_282);
nor U460 (N_460,N_391,N_390);
nor U461 (N_461,N_408,N_342);
or U462 (N_462,N_410,N_351);
and U463 (N_463,N_418,N_412);
nand U464 (N_464,N_415,N_351);
or U465 (N_465,N_403,N_372);
or U466 (N_466,N_388,N_342);
xnor U467 (N_467,N_368,N_132);
xnor U468 (N_468,N_254,N_386);
nor U469 (N_469,N_390,N_396);
or U470 (N_470,N_415,N_401);
nand U471 (N_471,N_410,N_414);
and U472 (N_472,N_390,N_250);
or U473 (N_473,N_418,N_373);
nand U474 (N_474,N_342,N_393);
and U475 (N_475,N_363,N_391);
and U476 (N_476,N_11,N_401);
nor U477 (N_477,N_395,N_282);
nand U478 (N_478,N_416,N_417);
nor U479 (N_479,N_324,N_396);
nand U480 (N_480,N_473,N_463);
and U481 (N_481,N_429,N_448);
and U482 (N_482,N_425,N_476);
and U483 (N_483,N_433,N_468);
nor U484 (N_484,N_437,N_443);
or U485 (N_485,N_455,N_469);
xor U486 (N_486,N_461,N_444);
or U487 (N_487,N_428,N_420);
xnor U488 (N_488,N_458,N_467);
nor U489 (N_489,N_472,N_452);
and U490 (N_490,N_440,N_427);
or U491 (N_491,N_453,N_445);
and U492 (N_492,N_441,N_471);
nor U493 (N_493,N_451,N_462);
nand U494 (N_494,N_439,N_466);
and U495 (N_495,N_465,N_454);
or U496 (N_496,N_479,N_475);
xor U497 (N_497,N_421,N_474);
xor U498 (N_498,N_449,N_460);
xor U499 (N_499,N_477,N_432);
nand U500 (N_500,N_435,N_434);
nor U501 (N_501,N_446,N_447);
or U502 (N_502,N_422,N_423);
or U503 (N_503,N_431,N_438);
nor U504 (N_504,N_457,N_426);
and U505 (N_505,N_478,N_470);
or U506 (N_506,N_424,N_456);
or U507 (N_507,N_464,N_430);
and U508 (N_508,N_450,N_459);
nand U509 (N_509,N_442,N_436);
and U510 (N_510,N_420,N_447);
nor U511 (N_511,N_465,N_467);
or U512 (N_512,N_425,N_462);
nand U513 (N_513,N_444,N_455);
and U514 (N_514,N_466,N_453);
nor U515 (N_515,N_476,N_469);
and U516 (N_516,N_459,N_427);
and U517 (N_517,N_450,N_435);
xnor U518 (N_518,N_433,N_444);
nand U519 (N_519,N_458,N_436);
nor U520 (N_520,N_435,N_433);
nand U521 (N_521,N_463,N_431);
nor U522 (N_522,N_468,N_436);
nor U523 (N_523,N_458,N_434);
and U524 (N_524,N_465,N_479);
or U525 (N_525,N_442,N_474);
or U526 (N_526,N_432,N_424);
and U527 (N_527,N_437,N_477);
or U528 (N_528,N_429,N_453);
nor U529 (N_529,N_429,N_464);
nor U530 (N_530,N_477,N_466);
nand U531 (N_531,N_438,N_424);
and U532 (N_532,N_471,N_432);
and U533 (N_533,N_455,N_468);
or U534 (N_534,N_439,N_451);
or U535 (N_535,N_449,N_442);
nor U536 (N_536,N_442,N_447);
xnor U537 (N_537,N_440,N_445);
nand U538 (N_538,N_474,N_434);
nand U539 (N_539,N_453,N_477);
nor U540 (N_540,N_497,N_535);
nor U541 (N_541,N_499,N_500);
and U542 (N_542,N_522,N_526);
and U543 (N_543,N_487,N_510);
or U544 (N_544,N_521,N_502);
xor U545 (N_545,N_491,N_516);
or U546 (N_546,N_525,N_486);
nand U547 (N_547,N_504,N_488);
nand U548 (N_548,N_483,N_481);
nor U549 (N_549,N_538,N_520);
nor U550 (N_550,N_505,N_519);
and U551 (N_551,N_529,N_537);
nor U552 (N_552,N_515,N_524);
nor U553 (N_553,N_539,N_518);
nand U554 (N_554,N_528,N_501);
or U555 (N_555,N_512,N_508);
nand U556 (N_556,N_531,N_523);
or U557 (N_557,N_533,N_480);
or U558 (N_558,N_489,N_485);
nor U559 (N_559,N_509,N_534);
nor U560 (N_560,N_530,N_513);
nor U561 (N_561,N_498,N_495);
nor U562 (N_562,N_517,N_511);
and U563 (N_563,N_507,N_527);
or U564 (N_564,N_503,N_532);
nand U565 (N_565,N_494,N_482);
and U566 (N_566,N_493,N_490);
nor U567 (N_567,N_492,N_484);
nor U568 (N_568,N_496,N_514);
or U569 (N_569,N_536,N_506);
nand U570 (N_570,N_536,N_523);
or U571 (N_571,N_508,N_496);
nor U572 (N_572,N_514,N_512);
nor U573 (N_573,N_499,N_526);
or U574 (N_574,N_539,N_527);
and U575 (N_575,N_529,N_538);
and U576 (N_576,N_490,N_517);
or U577 (N_577,N_510,N_497);
nand U578 (N_578,N_528,N_529);
nand U579 (N_579,N_505,N_485);
and U580 (N_580,N_493,N_520);
nand U581 (N_581,N_498,N_519);
nor U582 (N_582,N_538,N_482);
nand U583 (N_583,N_520,N_528);
nor U584 (N_584,N_481,N_503);
nor U585 (N_585,N_486,N_527);
and U586 (N_586,N_527,N_493);
xor U587 (N_587,N_511,N_514);
nor U588 (N_588,N_493,N_517);
xnor U589 (N_589,N_480,N_506);
or U590 (N_590,N_518,N_482);
nor U591 (N_591,N_496,N_513);
and U592 (N_592,N_511,N_534);
nor U593 (N_593,N_517,N_484);
nand U594 (N_594,N_504,N_517);
or U595 (N_595,N_515,N_495);
xnor U596 (N_596,N_503,N_499);
and U597 (N_597,N_520,N_517);
nor U598 (N_598,N_525,N_488);
nor U599 (N_599,N_490,N_489);
and U600 (N_600,N_582,N_552);
and U601 (N_601,N_586,N_564);
nor U602 (N_602,N_592,N_547);
or U603 (N_603,N_585,N_550);
nor U604 (N_604,N_540,N_598);
xnor U605 (N_605,N_583,N_590);
nand U606 (N_606,N_553,N_577);
and U607 (N_607,N_578,N_554);
and U608 (N_608,N_572,N_571);
nand U609 (N_609,N_595,N_570);
and U610 (N_610,N_549,N_597);
nor U611 (N_611,N_545,N_568);
and U612 (N_612,N_575,N_593);
nand U613 (N_613,N_561,N_567);
nand U614 (N_614,N_569,N_556);
and U615 (N_615,N_557,N_591);
nor U616 (N_616,N_596,N_543);
and U617 (N_617,N_551,N_555);
xor U618 (N_618,N_589,N_541);
and U619 (N_619,N_548,N_544);
nor U620 (N_620,N_559,N_581);
or U621 (N_621,N_560,N_563);
nor U622 (N_622,N_573,N_584);
or U623 (N_623,N_580,N_587);
nand U624 (N_624,N_562,N_588);
and U625 (N_625,N_566,N_542);
or U626 (N_626,N_576,N_565);
nand U627 (N_627,N_579,N_558);
or U628 (N_628,N_599,N_594);
xnor U629 (N_629,N_574,N_546);
xor U630 (N_630,N_598,N_548);
xor U631 (N_631,N_587,N_545);
xor U632 (N_632,N_568,N_571);
or U633 (N_633,N_556,N_562);
or U634 (N_634,N_574,N_594);
nand U635 (N_635,N_576,N_548);
nor U636 (N_636,N_552,N_546);
xor U637 (N_637,N_548,N_547);
nand U638 (N_638,N_563,N_586);
and U639 (N_639,N_546,N_550);
and U640 (N_640,N_587,N_548);
nand U641 (N_641,N_556,N_586);
nand U642 (N_642,N_596,N_588);
nor U643 (N_643,N_566,N_587);
and U644 (N_644,N_581,N_585);
nor U645 (N_645,N_552,N_598);
nor U646 (N_646,N_583,N_549);
xnor U647 (N_647,N_569,N_557);
nor U648 (N_648,N_573,N_554);
xnor U649 (N_649,N_571,N_570);
and U650 (N_650,N_563,N_593);
nand U651 (N_651,N_578,N_589);
nor U652 (N_652,N_564,N_544);
nand U653 (N_653,N_553,N_554);
nor U654 (N_654,N_581,N_553);
and U655 (N_655,N_591,N_558);
xnor U656 (N_656,N_560,N_549);
nor U657 (N_657,N_550,N_575);
or U658 (N_658,N_586,N_570);
or U659 (N_659,N_570,N_547);
nor U660 (N_660,N_649,N_656);
nand U661 (N_661,N_613,N_631);
nand U662 (N_662,N_608,N_648);
or U663 (N_663,N_607,N_645);
nand U664 (N_664,N_619,N_647);
nand U665 (N_665,N_616,N_654);
nand U666 (N_666,N_623,N_622);
nand U667 (N_667,N_626,N_615);
nand U668 (N_668,N_641,N_617);
nor U669 (N_669,N_625,N_612);
and U670 (N_670,N_633,N_610);
and U671 (N_671,N_637,N_602);
nand U672 (N_672,N_639,N_636);
or U673 (N_673,N_600,N_652);
and U674 (N_674,N_643,N_644);
and U675 (N_675,N_621,N_638);
or U676 (N_676,N_618,N_629);
xnor U677 (N_677,N_635,N_651);
xor U678 (N_678,N_601,N_653);
nor U679 (N_679,N_614,N_620);
nand U680 (N_680,N_658,N_657);
and U681 (N_681,N_604,N_605);
or U682 (N_682,N_630,N_609);
xnor U683 (N_683,N_627,N_603);
xor U684 (N_684,N_624,N_659);
nor U685 (N_685,N_642,N_632);
xnor U686 (N_686,N_628,N_606);
nor U687 (N_687,N_650,N_646);
nand U688 (N_688,N_640,N_634);
and U689 (N_689,N_655,N_611);
nand U690 (N_690,N_641,N_623);
or U691 (N_691,N_631,N_617);
nor U692 (N_692,N_645,N_642);
nor U693 (N_693,N_616,N_601);
nor U694 (N_694,N_610,N_650);
nand U695 (N_695,N_645,N_600);
nor U696 (N_696,N_655,N_601);
or U697 (N_697,N_656,N_647);
nor U698 (N_698,N_615,N_659);
nor U699 (N_699,N_628,N_643);
and U700 (N_700,N_609,N_632);
or U701 (N_701,N_619,N_608);
nor U702 (N_702,N_603,N_649);
nand U703 (N_703,N_611,N_651);
nand U704 (N_704,N_658,N_615);
nand U705 (N_705,N_608,N_629);
xor U706 (N_706,N_624,N_632);
or U707 (N_707,N_607,N_633);
or U708 (N_708,N_640,N_610);
and U709 (N_709,N_639,N_656);
or U710 (N_710,N_628,N_636);
nand U711 (N_711,N_639,N_625);
xnor U712 (N_712,N_606,N_651);
and U713 (N_713,N_600,N_628);
nand U714 (N_714,N_655,N_603);
or U715 (N_715,N_645,N_625);
or U716 (N_716,N_614,N_629);
nand U717 (N_717,N_638,N_612);
nand U718 (N_718,N_640,N_608);
and U719 (N_719,N_635,N_648);
nor U720 (N_720,N_702,N_685);
or U721 (N_721,N_682,N_708);
and U722 (N_722,N_660,N_710);
nand U723 (N_723,N_677,N_679);
nor U724 (N_724,N_706,N_699);
nor U725 (N_725,N_680,N_698);
nand U726 (N_726,N_671,N_666);
nand U727 (N_727,N_670,N_715);
nor U728 (N_728,N_673,N_686);
and U729 (N_729,N_668,N_712);
nor U730 (N_730,N_663,N_696);
nand U731 (N_731,N_678,N_694);
nand U732 (N_732,N_716,N_705);
nand U733 (N_733,N_697,N_695);
and U734 (N_734,N_711,N_681);
nor U735 (N_735,N_701,N_717);
nand U736 (N_736,N_661,N_719);
or U737 (N_737,N_669,N_667);
nor U738 (N_738,N_700,N_688);
nand U739 (N_739,N_704,N_674);
and U740 (N_740,N_687,N_692);
nor U741 (N_741,N_664,N_713);
or U742 (N_742,N_714,N_707);
xnor U743 (N_743,N_718,N_689);
nand U744 (N_744,N_693,N_675);
nand U745 (N_745,N_665,N_690);
and U746 (N_746,N_676,N_684);
and U747 (N_747,N_709,N_683);
and U748 (N_748,N_672,N_662);
or U749 (N_749,N_703,N_691);
nor U750 (N_750,N_663,N_707);
or U751 (N_751,N_711,N_709);
nand U752 (N_752,N_698,N_708);
and U753 (N_753,N_677,N_715);
nand U754 (N_754,N_700,N_712);
or U755 (N_755,N_688,N_680);
nand U756 (N_756,N_699,N_669);
or U757 (N_757,N_715,N_709);
or U758 (N_758,N_664,N_710);
nand U759 (N_759,N_668,N_682);
nor U760 (N_760,N_687,N_695);
or U761 (N_761,N_702,N_714);
or U762 (N_762,N_690,N_674);
nor U763 (N_763,N_661,N_678);
and U764 (N_764,N_714,N_674);
nand U765 (N_765,N_660,N_696);
and U766 (N_766,N_701,N_714);
nor U767 (N_767,N_717,N_666);
and U768 (N_768,N_714,N_664);
xor U769 (N_769,N_673,N_705);
and U770 (N_770,N_706,N_712);
and U771 (N_771,N_701,N_679);
nand U772 (N_772,N_661,N_703);
nand U773 (N_773,N_696,N_662);
nor U774 (N_774,N_702,N_679);
nor U775 (N_775,N_663,N_714);
and U776 (N_776,N_714,N_719);
nor U777 (N_777,N_706,N_663);
nor U778 (N_778,N_714,N_665);
nor U779 (N_779,N_695,N_696);
and U780 (N_780,N_721,N_735);
and U781 (N_781,N_755,N_767);
nor U782 (N_782,N_756,N_764);
nand U783 (N_783,N_733,N_777);
and U784 (N_784,N_732,N_724);
and U785 (N_785,N_760,N_737);
and U786 (N_786,N_725,N_741);
nand U787 (N_787,N_745,N_779);
nor U788 (N_788,N_722,N_772);
nand U789 (N_789,N_751,N_774);
or U790 (N_790,N_765,N_738);
nand U791 (N_791,N_734,N_743);
xor U792 (N_792,N_740,N_730);
xnor U793 (N_793,N_778,N_752);
and U794 (N_794,N_747,N_746);
nand U795 (N_795,N_723,N_769);
and U796 (N_796,N_757,N_775);
nor U797 (N_797,N_748,N_736);
xor U798 (N_798,N_728,N_771);
or U799 (N_799,N_768,N_773);
and U800 (N_800,N_739,N_770);
or U801 (N_801,N_750,N_731);
xor U802 (N_802,N_744,N_729);
and U803 (N_803,N_761,N_727);
and U804 (N_804,N_776,N_753);
nand U805 (N_805,N_766,N_763);
and U806 (N_806,N_754,N_758);
nand U807 (N_807,N_742,N_749);
and U808 (N_808,N_726,N_720);
or U809 (N_809,N_762,N_759);
nor U810 (N_810,N_743,N_776);
or U811 (N_811,N_741,N_745);
nand U812 (N_812,N_735,N_766);
or U813 (N_813,N_770,N_726);
or U814 (N_814,N_735,N_779);
nand U815 (N_815,N_763,N_753);
nand U816 (N_816,N_759,N_763);
nor U817 (N_817,N_748,N_738);
nand U818 (N_818,N_726,N_761);
nand U819 (N_819,N_735,N_761);
nand U820 (N_820,N_732,N_751);
or U821 (N_821,N_763,N_758);
or U822 (N_822,N_752,N_734);
xor U823 (N_823,N_740,N_779);
nor U824 (N_824,N_775,N_727);
nand U825 (N_825,N_766,N_742);
nor U826 (N_826,N_767,N_777);
nand U827 (N_827,N_761,N_731);
nand U828 (N_828,N_765,N_724);
and U829 (N_829,N_752,N_735);
nor U830 (N_830,N_747,N_757);
and U831 (N_831,N_720,N_770);
nand U832 (N_832,N_773,N_759);
nand U833 (N_833,N_773,N_766);
or U834 (N_834,N_723,N_755);
xor U835 (N_835,N_764,N_732);
nand U836 (N_836,N_727,N_725);
nor U837 (N_837,N_767,N_731);
or U838 (N_838,N_772,N_741);
or U839 (N_839,N_725,N_734);
and U840 (N_840,N_806,N_829);
and U841 (N_841,N_828,N_798);
or U842 (N_842,N_804,N_822);
and U843 (N_843,N_830,N_796);
and U844 (N_844,N_808,N_831);
xor U845 (N_845,N_816,N_817);
nor U846 (N_846,N_780,N_791);
nor U847 (N_847,N_781,N_792);
nand U848 (N_848,N_787,N_805);
and U849 (N_849,N_832,N_834);
and U850 (N_850,N_826,N_790);
nand U851 (N_851,N_800,N_799);
or U852 (N_852,N_838,N_794);
or U853 (N_853,N_784,N_810);
and U854 (N_854,N_818,N_807);
nand U855 (N_855,N_809,N_786);
and U856 (N_856,N_839,N_835);
and U857 (N_857,N_783,N_823);
and U858 (N_858,N_793,N_827);
or U859 (N_859,N_812,N_801);
nand U860 (N_860,N_820,N_814);
xnor U861 (N_861,N_819,N_785);
nand U862 (N_862,N_824,N_797);
and U863 (N_863,N_837,N_821);
nor U864 (N_864,N_836,N_815);
and U865 (N_865,N_833,N_813);
and U866 (N_866,N_825,N_803);
nand U867 (N_867,N_788,N_789);
nor U868 (N_868,N_811,N_782);
nand U869 (N_869,N_795,N_802);
nor U870 (N_870,N_792,N_804);
or U871 (N_871,N_783,N_815);
or U872 (N_872,N_798,N_811);
or U873 (N_873,N_834,N_816);
nor U874 (N_874,N_824,N_785);
or U875 (N_875,N_809,N_816);
xor U876 (N_876,N_827,N_816);
nand U877 (N_877,N_785,N_789);
xor U878 (N_878,N_785,N_809);
nor U879 (N_879,N_799,N_823);
and U880 (N_880,N_829,N_811);
nand U881 (N_881,N_825,N_823);
nor U882 (N_882,N_793,N_820);
or U883 (N_883,N_798,N_795);
or U884 (N_884,N_783,N_832);
and U885 (N_885,N_836,N_817);
or U886 (N_886,N_822,N_823);
nor U887 (N_887,N_791,N_827);
nor U888 (N_888,N_815,N_809);
nand U889 (N_889,N_826,N_813);
and U890 (N_890,N_826,N_834);
nor U891 (N_891,N_788,N_798);
and U892 (N_892,N_798,N_839);
and U893 (N_893,N_815,N_808);
xnor U894 (N_894,N_802,N_792);
nand U895 (N_895,N_803,N_830);
or U896 (N_896,N_819,N_838);
nor U897 (N_897,N_792,N_797);
or U898 (N_898,N_822,N_795);
or U899 (N_899,N_784,N_828);
nand U900 (N_900,N_878,N_852);
and U901 (N_901,N_886,N_848);
or U902 (N_902,N_872,N_888);
nor U903 (N_903,N_856,N_877);
nand U904 (N_904,N_873,N_858);
nand U905 (N_905,N_862,N_857);
nand U906 (N_906,N_844,N_899);
or U907 (N_907,N_882,N_849);
nor U908 (N_908,N_885,N_896);
nand U909 (N_909,N_850,N_842);
nand U910 (N_910,N_861,N_840);
nand U911 (N_911,N_887,N_865);
and U912 (N_912,N_889,N_853);
or U913 (N_913,N_894,N_890);
xnor U914 (N_914,N_866,N_895);
or U915 (N_915,N_854,N_879);
nor U916 (N_916,N_841,N_892);
nand U917 (N_917,N_898,N_864);
xor U918 (N_918,N_867,N_880);
and U919 (N_919,N_869,N_843);
nor U920 (N_920,N_846,N_847);
nand U921 (N_921,N_863,N_860);
and U922 (N_922,N_881,N_870);
nor U923 (N_923,N_875,N_891);
and U924 (N_924,N_876,N_883);
nor U925 (N_925,N_874,N_871);
or U926 (N_926,N_893,N_851);
nor U927 (N_927,N_859,N_884);
nor U928 (N_928,N_897,N_845);
nor U929 (N_929,N_868,N_855);
and U930 (N_930,N_858,N_849);
or U931 (N_931,N_865,N_848);
and U932 (N_932,N_864,N_888);
and U933 (N_933,N_851,N_858);
nor U934 (N_934,N_849,N_896);
nor U935 (N_935,N_849,N_873);
nor U936 (N_936,N_892,N_845);
and U937 (N_937,N_893,N_858);
or U938 (N_938,N_896,N_844);
and U939 (N_939,N_858,N_840);
xnor U940 (N_940,N_890,N_854);
and U941 (N_941,N_841,N_891);
and U942 (N_942,N_871,N_844);
xnor U943 (N_943,N_851,N_880);
and U944 (N_944,N_889,N_857);
and U945 (N_945,N_891,N_861);
or U946 (N_946,N_863,N_895);
or U947 (N_947,N_853,N_883);
nor U948 (N_948,N_869,N_881);
nand U949 (N_949,N_880,N_841);
nor U950 (N_950,N_854,N_842);
and U951 (N_951,N_873,N_860);
and U952 (N_952,N_881,N_847);
nor U953 (N_953,N_887,N_864);
or U954 (N_954,N_896,N_898);
or U955 (N_955,N_879,N_877);
and U956 (N_956,N_889,N_852);
or U957 (N_957,N_892,N_848);
or U958 (N_958,N_861,N_875);
and U959 (N_959,N_869,N_848);
or U960 (N_960,N_954,N_946);
nand U961 (N_961,N_903,N_909);
nand U962 (N_962,N_902,N_952);
or U963 (N_963,N_908,N_901);
or U964 (N_964,N_937,N_951);
or U965 (N_965,N_912,N_923);
or U966 (N_966,N_905,N_943);
xor U967 (N_967,N_915,N_956);
or U968 (N_968,N_957,N_935);
or U969 (N_969,N_945,N_925);
or U970 (N_970,N_959,N_928);
and U971 (N_971,N_911,N_918);
nand U972 (N_972,N_947,N_944);
nor U973 (N_973,N_920,N_906);
or U974 (N_974,N_917,N_900);
nor U975 (N_975,N_924,N_936);
and U976 (N_976,N_929,N_916);
and U977 (N_977,N_949,N_919);
nor U978 (N_978,N_933,N_931);
nand U979 (N_979,N_926,N_907);
nor U980 (N_980,N_922,N_941);
nor U981 (N_981,N_948,N_913);
or U982 (N_982,N_955,N_938);
nand U983 (N_983,N_921,N_904);
or U984 (N_984,N_910,N_932);
nor U985 (N_985,N_958,N_939);
and U986 (N_986,N_940,N_927);
or U987 (N_987,N_953,N_914);
xnor U988 (N_988,N_942,N_930);
and U989 (N_989,N_950,N_934);
and U990 (N_990,N_937,N_956);
xnor U991 (N_991,N_926,N_912);
xor U992 (N_992,N_918,N_917);
xor U993 (N_993,N_949,N_907);
xor U994 (N_994,N_902,N_910);
and U995 (N_995,N_939,N_957);
xor U996 (N_996,N_929,N_949);
xnor U997 (N_997,N_937,N_923);
nand U998 (N_998,N_902,N_936);
xnor U999 (N_999,N_953,N_952);
nor U1000 (N_1000,N_925,N_922);
or U1001 (N_1001,N_905,N_912);
nand U1002 (N_1002,N_942,N_917);
nand U1003 (N_1003,N_953,N_903);
nand U1004 (N_1004,N_954,N_950);
and U1005 (N_1005,N_912,N_945);
nand U1006 (N_1006,N_912,N_930);
nand U1007 (N_1007,N_941,N_926);
and U1008 (N_1008,N_946,N_934);
and U1009 (N_1009,N_956,N_911);
or U1010 (N_1010,N_921,N_928);
and U1011 (N_1011,N_955,N_905);
nand U1012 (N_1012,N_938,N_912);
xor U1013 (N_1013,N_943,N_944);
nand U1014 (N_1014,N_905,N_907);
xnor U1015 (N_1015,N_916,N_910);
xnor U1016 (N_1016,N_940,N_923);
nor U1017 (N_1017,N_944,N_918);
and U1018 (N_1018,N_930,N_908);
nor U1019 (N_1019,N_930,N_915);
nor U1020 (N_1020,N_975,N_1012);
and U1021 (N_1021,N_995,N_985);
and U1022 (N_1022,N_987,N_961);
or U1023 (N_1023,N_1008,N_999);
xor U1024 (N_1024,N_1018,N_969);
nand U1025 (N_1025,N_1001,N_972);
nor U1026 (N_1026,N_965,N_996);
or U1027 (N_1027,N_986,N_962);
nor U1028 (N_1028,N_973,N_1003);
xnor U1029 (N_1029,N_978,N_982);
nor U1030 (N_1030,N_1005,N_991);
and U1031 (N_1031,N_979,N_1002);
and U1032 (N_1032,N_1019,N_997);
and U1033 (N_1033,N_989,N_968);
nor U1034 (N_1034,N_976,N_1014);
or U1035 (N_1035,N_971,N_1013);
nor U1036 (N_1036,N_983,N_1011);
nand U1037 (N_1037,N_990,N_966);
and U1038 (N_1038,N_993,N_980);
xnor U1039 (N_1039,N_977,N_1017);
nand U1040 (N_1040,N_984,N_1006);
and U1041 (N_1041,N_1016,N_1004);
or U1042 (N_1042,N_967,N_1007);
nor U1043 (N_1043,N_988,N_963);
nor U1044 (N_1044,N_1015,N_998);
nor U1045 (N_1045,N_960,N_1009);
or U1046 (N_1046,N_1000,N_974);
xor U1047 (N_1047,N_992,N_981);
nand U1048 (N_1048,N_970,N_964);
nor U1049 (N_1049,N_1010,N_994);
and U1050 (N_1050,N_999,N_1004);
nand U1051 (N_1051,N_973,N_1011);
or U1052 (N_1052,N_979,N_992);
and U1053 (N_1053,N_1009,N_1018);
nand U1054 (N_1054,N_995,N_1016);
and U1055 (N_1055,N_1007,N_983);
and U1056 (N_1056,N_997,N_994);
or U1057 (N_1057,N_1017,N_976);
nor U1058 (N_1058,N_1005,N_1015);
nor U1059 (N_1059,N_967,N_970);
nand U1060 (N_1060,N_1019,N_1012);
or U1061 (N_1061,N_999,N_981);
nand U1062 (N_1062,N_968,N_1005);
and U1063 (N_1063,N_976,N_1016);
nand U1064 (N_1064,N_1013,N_967);
or U1065 (N_1065,N_1019,N_1011);
and U1066 (N_1066,N_987,N_992);
and U1067 (N_1067,N_974,N_962);
and U1068 (N_1068,N_970,N_983);
nor U1069 (N_1069,N_977,N_968);
nand U1070 (N_1070,N_976,N_988);
nand U1071 (N_1071,N_969,N_1011);
and U1072 (N_1072,N_1003,N_960);
nand U1073 (N_1073,N_985,N_983);
nand U1074 (N_1074,N_969,N_1007);
nor U1075 (N_1075,N_964,N_1011);
xnor U1076 (N_1076,N_1017,N_974);
or U1077 (N_1077,N_970,N_1005);
or U1078 (N_1078,N_1018,N_992);
and U1079 (N_1079,N_1013,N_1019);
nor U1080 (N_1080,N_1025,N_1056);
xor U1081 (N_1081,N_1052,N_1028);
nor U1082 (N_1082,N_1069,N_1040);
nor U1083 (N_1083,N_1043,N_1039);
nor U1084 (N_1084,N_1021,N_1051);
nand U1085 (N_1085,N_1060,N_1027);
xnor U1086 (N_1086,N_1048,N_1068);
and U1087 (N_1087,N_1065,N_1020);
nand U1088 (N_1088,N_1041,N_1058);
or U1089 (N_1089,N_1061,N_1042);
nand U1090 (N_1090,N_1054,N_1071);
or U1091 (N_1091,N_1049,N_1075);
or U1092 (N_1092,N_1055,N_1029);
nor U1093 (N_1093,N_1074,N_1036);
or U1094 (N_1094,N_1022,N_1079);
or U1095 (N_1095,N_1078,N_1050);
and U1096 (N_1096,N_1077,N_1034);
nor U1097 (N_1097,N_1046,N_1031);
nand U1098 (N_1098,N_1035,N_1024);
xnor U1099 (N_1099,N_1063,N_1072);
or U1100 (N_1100,N_1064,N_1044);
or U1101 (N_1101,N_1059,N_1076);
and U1102 (N_1102,N_1033,N_1066);
and U1103 (N_1103,N_1053,N_1057);
nor U1104 (N_1104,N_1032,N_1038);
or U1105 (N_1105,N_1067,N_1030);
or U1106 (N_1106,N_1045,N_1037);
nand U1107 (N_1107,N_1047,N_1023);
nand U1108 (N_1108,N_1062,N_1070);
nor U1109 (N_1109,N_1073,N_1026);
nand U1110 (N_1110,N_1034,N_1038);
xor U1111 (N_1111,N_1077,N_1057);
and U1112 (N_1112,N_1074,N_1044);
or U1113 (N_1113,N_1078,N_1029);
nor U1114 (N_1114,N_1067,N_1073);
or U1115 (N_1115,N_1043,N_1079);
nor U1116 (N_1116,N_1079,N_1028);
xor U1117 (N_1117,N_1079,N_1057);
and U1118 (N_1118,N_1046,N_1030);
xnor U1119 (N_1119,N_1049,N_1079);
nand U1120 (N_1120,N_1029,N_1056);
or U1121 (N_1121,N_1041,N_1028);
nand U1122 (N_1122,N_1023,N_1026);
nor U1123 (N_1123,N_1040,N_1070);
nor U1124 (N_1124,N_1026,N_1047);
or U1125 (N_1125,N_1046,N_1077);
nor U1126 (N_1126,N_1028,N_1022);
and U1127 (N_1127,N_1074,N_1078);
or U1128 (N_1128,N_1072,N_1061);
nor U1129 (N_1129,N_1075,N_1046);
or U1130 (N_1130,N_1035,N_1030);
nor U1131 (N_1131,N_1031,N_1067);
nand U1132 (N_1132,N_1045,N_1044);
or U1133 (N_1133,N_1064,N_1063);
nor U1134 (N_1134,N_1044,N_1030);
or U1135 (N_1135,N_1054,N_1036);
nand U1136 (N_1136,N_1023,N_1050);
nor U1137 (N_1137,N_1031,N_1059);
nand U1138 (N_1138,N_1062,N_1037);
nand U1139 (N_1139,N_1061,N_1048);
nor U1140 (N_1140,N_1132,N_1127);
nor U1141 (N_1141,N_1093,N_1124);
nor U1142 (N_1142,N_1099,N_1082);
nand U1143 (N_1143,N_1104,N_1131);
nand U1144 (N_1144,N_1121,N_1136);
or U1145 (N_1145,N_1128,N_1120);
nor U1146 (N_1146,N_1080,N_1118);
or U1147 (N_1147,N_1097,N_1137);
nand U1148 (N_1148,N_1085,N_1102);
nor U1149 (N_1149,N_1101,N_1092);
and U1150 (N_1150,N_1084,N_1123);
xnor U1151 (N_1151,N_1139,N_1109);
nor U1152 (N_1152,N_1115,N_1114);
or U1153 (N_1153,N_1107,N_1083);
nor U1154 (N_1154,N_1090,N_1126);
nor U1155 (N_1155,N_1089,N_1086);
nand U1156 (N_1156,N_1125,N_1112);
xor U1157 (N_1157,N_1095,N_1103);
or U1158 (N_1158,N_1098,N_1135);
and U1159 (N_1159,N_1100,N_1122);
nor U1160 (N_1160,N_1088,N_1096);
or U1161 (N_1161,N_1129,N_1110);
or U1162 (N_1162,N_1133,N_1081);
nor U1163 (N_1163,N_1106,N_1091);
or U1164 (N_1164,N_1094,N_1130);
and U1165 (N_1165,N_1138,N_1134);
and U1166 (N_1166,N_1108,N_1105);
nor U1167 (N_1167,N_1113,N_1119);
and U1168 (N_1168,N_1116,N_1117);
or U1169 (N_1169,N_1111,N_1087);
nor U1170 (N_1170,N_1094,N_1095);
nand U1171 (N_1171,N_1125,N_1137);
nor U1172 (N_1172,N_1132,N_1094);
nor U1173 (N_1173,N_1111,N_1138);
and U1174 (N_1174,N_1125,N_1129);
or U1175 (N_1175,N_1082,N_1124);
or U1176 (N_1176,N_1133,N_1110);
or U1177 (N_1177,N_1116,N_1104);
nor U1178 (N_1178,N_1091,N_1138);
nand U1179 (N_1179,N_1117,N_1129);
nor U1180 (N_1180,N_1125,N_1093);
nor U1181 (N_1181,N_1138,N_1133);
nor U1182 (N_1182,N_1101,N_1119);
nand U1183 (N_1183,N_1139,N_1099);
and U1184 (N_1184,N_1084,N_1080);
xnor U1185 (N_1185,N_1083,N_1128);
and U1186 (N_1186,N_1107,N_1129);
and U1187 (N_1187,N_1087,N_1130);
nand U1188 (N_1188,N_1125,N_1130);
and U1189 (N_1189,N_1110,N_1123);
nor U1190 (N_1190,N_1106,N_1098);
or U1191 (N_1191,N_1116,N_1101);
nand U1192 (N_1192,N_1115,N_1096);
and U1193 (N_1193,N_1087,N_1139);
nand U1194 (N_1194,N_1115,N_1111);
nand U1195 (N_1195,N_1092,N_1099);
nand U1196 (N_1196,N_1112,N_1084);
xnor U1197 (N_1197,N_1136,N_1113);
and U1198 (N_1198,N_1115,N_1113);
nand U1199 (N_1199,N_1084,N_1108);
nor U1200 (N_1200,N_1199,N_1143);
nor U1201 (N_1201,N_1142,N_1192);
nand U1202 (N_1202,N_1168,N_1178);
nor U1203 (N_1203,N_1162,N_1172);
nand U1204 (N_1204,N_1183,N_1197);
nand U1205 (N_1205,N_1169,N_1165);
nor U1206 (N_1206,N_1179,N_1188);
nand U1207 (N_1207,N_1186,N_1195);
xor U1208 (N_1208,N_1190,N_1166);
nor U1209 (N_1209,N_1157,N_1176);
nor U1210 (N_1210,N_1163,N_1155);
nor U1211 (N_1211,N_1150,N_1144);
or U1212 (N_1212,N_1196,N_1177);
or U1213 (N_1213,N_1175,N_1174);
or U1214 (N_1214,N_1140,N_1173);
and U1215 (N_1215,N_1147,N_1160);
nor U1216 (N_1216,N_1158,N_1151);
nand U1217 (N_1217,N_1156,N_1181);
nand U1218 (N_1218,N_1149,N_1152);
nand U1219 (N_1219,N_1182,N_1161);
and U1220 (N_1220,N_1191,N_1187);
or U1221 (N_1221,N_1154,N_1146);
and U1222 (N_1222,N_1193,N_1153);
nand U1223 (N_1223,N_1198,N_1185);
nand U1224 (N_1224,N_1145,N_1171);
nor U1225 (N_1225,N_1189,N_1141);
and U1226 (N_1226,N_1180,N_1164);
nand U1227 (N_1227,N_1148,N_1184);
or U1228 (N_1228,N_1167,N_1159);
or U1229 (N_1229,N_1194,N_1170);
nand U1230 (N_1230,N_1142,N_1199);
or U1231 (N_1231,N_1174,N_1160);
nor U1232 (N_1232,N_1194,N_1162);
or U1233 (N_1233,N_1180,N_1143);
or U1234 (N_1234,N_1191,N_1183);
nor U1235 (N_1235,N_1172,N_1198);
nor U1236 (N_1236,N_1144,N_1193);
and U1237 (N_1237,N_1151,N_1152);
nor U1238 (N_1238,N_1144,N_1178);
nor U1239 (N_1239,N_1177,N_1180);
or U1240 (N_1240,N_1158,N_1170);
or U1241 (N_1241,N_1184,N_1150);
nand U1242 (N_1242,N_1148,N_1182);
and U1243 (N_1243,N_1140,N_1145);
and U1244 (N_1244,N_1176,N_1186);
and U1245 (N_1245,N_1176,N_1191);
or U1246 (N_1246,N_1148,N_1156);
or U1247 (N_1247,N_1141,N_1150);
nand U1248 (N_1248,N_1181,N_1192);
nand U1249 (N_1249,N_1148,N_1172);
nand U1250 (N_1250,N_1186,N_1178);
nor U1251 (N_1251,N_1179,N_1146);
or U1252 (N_1252,N_1191,N_1188);
nand U1253 (N_1253,N_1187,N_1169);
and U1254 (N_1254,N_1185,N_1188);
nor U1255 (N_1255,N_1158,N_1198);
xnor U1256 (N_1256,N_1197,N_1172);
xor U1257 (N_1257,N_1176,N_1163);
nor U1258 (N_1258,N_1173,N_1187);
and U1259 (N_1259,N_1182,N_1185);
nor U1260 (N_1260,N_1220,N_1231);
nand U1261 (N_1261,N_1201,N_1204);
and U1262 (N_1262,N_1250,N_1209);
nor U1263 (N_1263,N_1208,N_1207);
or U1264 (N_1264,N_1249,N_1243);
and U1265 (N_1265,N_1232,N_1256);
or U1266 (N_1266,N_1234,N_1241);
xnor U1267 (N_1267,N_1237,N_1235);
nand U1268 (N_1268,N_1206,N_1225);
or U1269 (N_1269,N_1222,N_1212);
and U1270 (N_1270,N_1257,N_1244);
and U1271 (N_1271,N_1217,N_1200);
xor U1272 (N_1272,N_1229,N_1223);
and U1273 (N_1273,N_1245,N_1238);
nor U1274 (N_1274,N_1205,N_1242);
and U1275 (N_1275,N_1254,N_1213);
and U1276 (N_1276,N_1202,N_1210);
nor U1277 (N_1277,N_1259,N_1233);
or U1278 (N_1278,N_1216,N_1224);
or U1279 (N_1279,N_1214,N_1219);
nor U1280 (N_1280,N_1226,N_1227);
or U1281 (N_1281,N_1253,N_1240);
nor U1282 (N_1282,N_1246,N_1215);
and U1283 (N_1283,N_1258,N_1255);
and U1284 (N_1284,N_1230,N_1228);
or U1285 (N_1285,N_1236,N_1218);
and U1286 (N_1286,N_1211,N_1252);
nand U1287 (N_1287,N_1203,N_1251);
or U1288 (N_1288,N_1239,N_1221);
nor U1289 (N_1289,N_1248,N_1247);
or U1290 (N_1290,N_1242,N_1248);
or U1291 (N_1291,N_1224,N_1244);
nor U1292 (N_1292,N_1212,N_1251);
nor U1293 (N_1293,N_1245,N_1216);
nand U1294 (N_1294,N_1209,N_1227);
nand U1295 (N_1295,N_1259,N_1237);
nor U1296 (N_1296,N_1253,N_1230);
nor U1297 (N_1297,N_1218,N_1233);
or U1298 (N_1298,N_1252,N_1253);
nor U1299 (N_1299,N_1238,N_1257);
nand U1300 (N_1300,N_1229,N_1226);
or U1301 (N_1301,N_1253,N_1228);
nand U1302 (N_1302,N_1235,N_1244);
nand U1303 (N_1303,N_1232,N_1247);
or U1304 (N_1304,N_1235,N_1255);
xnor U1305 (N_1305,N_1211,N_1259);
nand U1306 (N_1306,N_1254,N_1200);
xor U1307 (N_1307,N_1237,N_1231);
or U1308 (N_1308,N_1236,N_1213);
xor U1309 (N_1309,N_1253,N_1238);
or U1310 (N_1310,N_1221,N_1203);
or U1311 (N_1311,N_1230,N_1251);
nand U1312 (N_1312,N_1213,N_1256);
and U1313 (N_1313,N_1233,N_1244);
or U1314 (N_1314,N_1252,N_1258);
or U1315 (N_1315,N_1256,N_1204);
or U1316 (N_1316,N_1247,N_1206);
and U1317 (N_1317,N_1219,N_1229);
xor U1318 (N_1318,N_1245,N_1215);
nor U1319 (N_1319,N_1209,N_1215);
nand U1320 (N_1320,N_1260,N_1317);
or U1321 (N_1321,N_1303,N_1271);
nor U1322 (N_1322,N_1273,N_1265);
and U1323 (N_1323,N_1272,N_1307);
and U1324 (N_1324,N_1295,N_1270);
or U1325 (N_1325,N_1289,N_1269);
or U1326 (N_1326,N_1306,N_1262);
nand U1327 (N_1327,N_1286,N_1267);
nor U1328 (N_1328,N_1281,N_1283);
and U1329 (N_1329,N_1288,N_1309);
and U1330 (N_1330,N_1284,N_1266);
nor U1331 (N_1331,N_1314,N_1274);
or U1332 (N_1332,N_1312,N_1296);
or U1333 (N_1333,N_1292,N_1300);
nor U1334 (N_1334,N_1311,N_1308);
nor U1335 (N_1335,N_1294,N_1299);
nor U1336 (N_1336,N_1297,N_1298);
nand U1337 (N_1337,N_1310,N_1263);
or U1338 (N_1338,N_1261,N_1291);
and U1339 (N_1339,N_1276,N_1313);
xnor U1340 (N_1340,N_1315,N_1277);
or U1341 (N_1341,N_1282,N_1318);
and U1342 (N_1342,N_1285,N_1319);
or U1343 (N_1343,N_1304,N_1290);
or U1344 (N_1344,N_1275,N_1316);
nand U1345 (N_1345,N_1268,N_1278);
nand U1346 (N_1346,N_1301,N_1305);
nand U1347 (N_1347,N_1302,N_1280);
nor U1348 (N_1348,N_1287,N_1293);
nand U1349 (N_1349,N_1264,N_1279);
nand U1350 (N_1350,N_1266,N_1272);
and U1351 (N_1351,N_1292,N_1319);
nand U1352 (N_1352,N_1317,N_1319);
or U1353 (N_1353,N_1286,N_1315);
and U1354 (N_1354,N_1318,N_1260);
xnor U1355 (N_1355,N_1274,N_1270);
or U1356 (N_1356,N_1288,N_1305);
or U1357 (N_1357,N_1301,N_1272);
nor U1358 (N_1358,N_1293,N_1291);
or U1359 (N_1359,N_1266,N_1296);
or U1360 (N_1360,N_1304,N_1319);
nor U1361 (N_1361,N_1269,N_1272);
or U1362 (N_1362,N_1284,N_1278);
and U1363 (N_1363,N_1295,N_1280);
or U1364 (N_1364,N_1299,N_1264);
nand U1365 (N_1365,N_1304,N_1299);
or U1366 (N_1366,N_1260,N_1292);
and U1367 (N_1367,N_1291,N_1310);
or U1368 (N_1368,N_1317,N_1294);
nand U1369 (N_1369,N_1308,N_1297);
xnor U1370 (N_1370,N_1308,N_1277);
or U1371 (N_1371,N_1308,N_1313);
and U1372 (N_1372,N_1298,N_1282);
or U1373 (N_1373,N_1272,N_1264);
and U1374 (N_1374,N_1312,N_1268);
nor U1375 (N_1375,N_1291,N_1284);
or U1376 (N_1376,N_1290,N_1316);
nand U1377 (N_1377,N_1268,N_1303);
xor U1378 (N_1378,N_1318,N_1276);
or U1379 (N_1379,N_1313,N_1303);
nand U1380 (N_1380,N_1323,N_1347);
and U1381 (N_1381,N_1364,N_1352);
and U1382 (N_1382,N_1362,N_1360);
and U1383 (N_1383,N_1349,N_1325);
nor U1384 (N_1384,N_1375,N_1324);
nand U1385 (N_1385,N_1377,N_1378);
and U1386 (N_1386,N_1340,N_1331);
and U1387 (N_1387,N_1350,N_1334);
or U1388 (N_1388,N_1327,N_1365);
or U1389 (N_1389,N_1348,N_1345);
or U1390 (N_1390,N_1354,N_1330);
nor U1391 (N_1391,N_1370,N_1335);
and U1392 (N_1392,N_1367,N_1333);
and U1393 (N_1393,N_1379,N_1359);
or U1394 (N_1394,N_1329,N_1357);
nor U1395 (N_1395,N_1374,N_1342);
or U1396 (N_1396,N_1353,N_1376);
nor U1397 (N_1397,N_1363,N_1356);
nor U1398 (N_1398,N_1344,N_1343);
nor U1399 (N_1399,N_1368,N_1358);
nor U1400 (N_1400,N_1328,N_1369);
nor U1401 (N_1401,N_1336,N_1339);
xor U1402 (N_1402,N_1321,N_1373);
or U1403 (N_1403,N_1338,N_1322);
or U1404 (N_1404,N_1320,N_1332);
nor U1405 (N_1405,N_1346,N_1326);
nand U1406 (N_1406,N_1366,N_1372);
or U1407 (N_1407,N_1351,N_1341);
nand U1408 (N_1408,N_1355,N_1371);
nand U1409 (N_1409,N_1361,N_1337);
nand U1410 (N_1410,N_1323,N_1358);
nand U1411 (N_1411,N_1353,N_1368);
and U1412 (N_1412,N_1351,N_1379);
and U1413 (N_1413,N_1329,N_1323);
xnor U1414 (N_1414,N_1327,N_1328);
nor U1415 (N_1415,N_1368,N_1346);
and U1416 (N_1416,N_1373,N_1365);
nor U1417 (N_1417,N_1329,N_1358);
or U1418 (N_1418,N_1353,N_1329);
and U1419 (N_1419,N_1340,N_1325);
nand U1420 (N_1420,N_1322,N_1328);
or U1421 (N_1421,N_1340,N_1339);
and U1422 (N_1422,N_1338,N_1368);
and U1423 (N_1423,N_1350,N_1328);
nor U1424 (N_1424,N_1338,N_1331);
nand U1425 (N_1425,N_1371,N_1357);
xor U1426 (N_1426,N_1378,N_1333);
nor U1427 (N_1427,N_1325,N_1357);
nor U1428 (N_1428,N_1328,N_1336);
or U1429 (N_1429,N_1344,N_1372);
or U1430 (N_1430,N_1325,N_1337);
or U1431 (N_1431,N_1361,N_1322);
and U1432 (N_1432,N_1374,N_1341);
nor U1433 (N_1433,N_1330,N_1339);
nand U1434 (N_1434,N_1337,N_1321);
or U1435 (N_1435,N_1365,N_1364);
or U1436 (N_1436,N_1372,N_1331);
nor U1437 (N_1437,N_1344,N_1377);
or U1438 (N_1438,N_1335,N_1332);
or U1439 (N_1439,N_1362,N_1350);
nor U1440 (N_1440,N_1412,N_1424);
nand U1441 (N_1441,N_1393,N_1413);
nand U1442 (N_1442,N_1434,N_1385);
nand U1443 (N_1443,N_1405,N_1388);
nor U1444 (N_1444,N_1425,N_1384);
or U1445 (N_1445,N_1398,N_1382);
nor U1446 (N_1446,N_1406,N_1404);
and U1447 (N_1447,N_1414,N_1430);
xor U1448 (N_1448,N_1399,N_1436);
nor U1449 (N_1449,N_1416,N_1418);
or U1450 (N_1450,N_1387,N_1420);
and U1451 (N_1451,N_1391,N_1429);
xor U1452 (N_1452,N_1433,N_1421);
and U1453 (N_1453,N_1415,N_1396);
xor U1454 (N_1454,N_1435,N_1397);
nand U1455 (N_1455,N_1380,N_1417);
or U1456 (N_1456,N_1426,N_1400);
nand U1457 (N_1457,N_1427,N_1423);
nor U1458 (N_1458,N_1437,N_1390);
nor U1459 (N_1459,N_1386,N_1383);
nor U1460 (N_1460,N_1438,N_1408);
and U1461 (N_1461,N_1403,N_1381);
or U1462 (N_1462,N_1395,N_1439);
or U1463 (N_1463,N_1409,N_1410);
or U1464 (N_1464,N_1432,N_1392);
or U1465 (N_1465,N_1419,N_1402);
nand U1466 (N_1466,N_1407,N_1431);
nor U1467 (N_1467,N_1411,N_1422);
and U1468 (N_1468,N_1389,N_1428);
nand U1469 (N_1469,N_1401,N_1394);
nor U1470 (N_1470,N_1420,N_1430);
or U1471 (N_1471,N_1389,N_1409);
and U1472 (N_1472,N_1399,N_1435);
xnor U1473 (N_1473,N_1395,N_1387);
nor U1474 (N_1474,N_1389,N_1397);
xnor U1475 (N_1475,N_1381,N_1399);
nand U1476 (N_1476,N_1426,N_1425);
nand U1477 (N_1477,N_1393,N_1424);
nor U1478 (N_1478,N_1439,N_1408);
nor U1479 (N_1479,N_1380,N_1438);
and U1480 (N_1480,N_1394,N_1432);
and U1481 (N_1481,N_1386,N_1437);
xnor U1482 (N_1482,N_1403,N_1398);
or U1483 (N_1483,N_1381,N_1433);
or U1484 (N_1484,N_1398,N_1409);
and U1485 (N_1485,N_1388,N_1398);
nand U1486 (N_1486,N_1401,N_1381);
nand U1487 (N_1487,N_1381,N_1429);
nand U1488 (N_1488,N_1429,N_1405);
and U1489 (N_1489,N_1389,N_1419);
and U1490 (N_1490,N_1418,N_1385);
nor U1491 (N_1491,N_1401,N_1438);
nand U1492 (N_1492,N_1411,N_1437);
and U1493 (N_1493,N_1433,N_1397);
and U1494 (N_1494,N_1381,N_1392);
or U1495 (N_1495,N_1389,N_1423);
nand U1496 (N_1496,N_1422,N_1407);
and U1497 (N_1497,N_1418,N_1432);
and U1498 (N_1498,N_1401,N_1390);
or U1499 (N_1499,N_1419,N_1421);
xnor U1500 (N_1500,N_1467,N_1485);
nand U1501 (N_1501,N_1457,N_1488);
and U1502 (N_1502,N_1481,N_1451);
nand U1503 (N_1503,N_1497,N_1492);
and U1504 (N_1504,N_1480,N_1447);
nor U1505 (N_1505,N_1445,N_1450);
xor U1506 (N_1506,N_1499,N_1459);
xor U1507 (N_1507,N_1476,N_1477);
or U1508 (N_1508,N_1474,N_1441);
or U1509 (N_1509,N_1482,N_1469);
or U1510 (N_1510,N_1468,N_1493);
xnor U1511 (N_1511,N_1495,N_1498);
or U1512 (N_1512,N_1454,N_1463);
xnor U1513 (N_1513,N_1462,N_1496);
nor U1514 (N_1514,N_1452,N_1456);
nand U1515 (N_1515,N_1461,N_1478);
and U1516 (N_1516,N_1483,N_1464);
nand U1517 (N_1517,N_1470,N_1448);
or U1518 (N_1518,N_1443,N_1465);
nor U1519 (N_1519,N_1442,N_1440);
or U1520 (N_1520,N_1487,N_1490);
nor U1521 (N_1521,N_1460,N_1453);
or U1522 (N_1522,N_1484,N_1491);
nor U1523 (N_1523,N_1446,N_1494);
nor U1524 (N_1524,N_1444,N_1475);
and U1525 (N_1525,N_1455,N_1473);
nand U1526 (N_1526,N_1479,N_1458);
and U1527 (N_1527,N_1472,N_1486);
and U1528 (N_1528,N_1466,N_1471);
nand U1529 (N_1529,N_1489,N_1449);
or U1530 (N_1530,N_1483,N_1490);
nor U1531 (N_1531,N_1488,N_1478);
or U1532 (N_1532,N_1489,N_1469);
nor U1533 (N_1533,N_1457,N_1452);
nand U1534 (N_1534,N_1498,N_1455);
or U1535 (N_1535,N_1454,N_1480);
nand U1536 (N_1536,N_1482,N_1458);
and U1537 (N_1537,N_1494,N_1466);
nor U1538 (N_1538,N_1478,N_1484);
or U1539 (N_1539,N_1468,N_1447);
or U1540 (N_1540,N_1442,N_1473);
xor U1541 (N_1541,N_1484,N_1440);
nor U1542 (N_1542,N_1449,N_1460);
and U1543 (N_1543,N_1482,N_1488);
nand U1544 (N_1544,N_1476,N_1453);
nor U1545 (N_1545,N_1469,N_1456);
nor U1546 (N_1546,N_1447,N_1472);
xor U1547 (N_1547,N_1489,N_1446);
or U1548 (N_1548,N_1455,N_1499);
nand U1549 (N_1549,N_1470,N_1476);
or U1550 (N_1550,N_1461,N_1447);
nand U1551 (N_1551,N_1454,N_1445);
and U1552 (N_1552,N_1448,N_1494);
nand U1553 (N_1553,N_1448,N_1496);
nand U1554 (N_1554,N_1494,N_1468);
nor U1555 (N_1555,N_1483,N_1461);
and U1556 (N_1556,N_1440,N_1499);
or U1557 (N_1557,N_1440,N_1469);
xor U1558 (N_1558,N_1451,N_1463);
nand U1559 (N_1559,N_1461,N_1494);
or U1560 (N_1560,N_1535,N_1548);
nor U1561 (N_1561,N_1540,N_1533);
nor U1562 (N_1562,N_1549,N_1507);
nand U1563 (N_1563,N_1521,N_1534);
or U1564 (N_1564,N_1553,N_1552);
or U1565 (N_1565,N_1513,N_1539);
nand U1566 (N_1566,N_1547,N_1514);
and U1567 (N_1567,N_1541,N_1504);
nand U1568 (N_1568,N_1538,N_1502);
nor U1569 (N_1569,N_1511,N_1527);
nor U1570 (N_1570,N_1520,N_1529);
and U1571 (N_1571,N_1515,N_1530);
nand U1572 (N_1572,N_1528,N_1557);
nand U1573 (N_1573,N_1555,N_1523);
and U1574 (N_1574,N_1531,N_1512);
or U1575 (N_1575,N_1532,N_1554);
nor U1576 (N_1576,N_1546,N_1526);
or U1577 (N_1577,N_1542,N_1551);
nand U1578 (N_1578,N_1508,N_1518);
and U1579 (N_1579,N_1500,N_1556);
nand U1580 (N_1580,N_1543,N_1503);
xor U1581 (N_1581,N_1537,N_1501);
and U1582 (N_1582,N_1522,N_1506);
nand U1583 (N_1583,N_1524,N_1525);
nand U1584 (N_1584,N_1544,N_1516);
nor U1585 (N_1585,N_1559,N_1545);
or U1586 (N_1586,N_1505,N_1519);
and U1587 (N_1587,N_1558,N_1536);
and U1588 (N_1588,N_1509,N_1517);
nand U1589 (N_1589,N_1510,N_1550);
xnor U1590 (N_1590,N_1554,N_1559);
nand U1591 (N_1591,N_1510,N_1534);
and U1592 (N_1592,N_1534,N_1544);
nor U1593 (N_1593,N_1548,N_1551);
or U1594 (N_1594,N_1534,N_1555);
nand U1595 (N_1595,N_1518,N_1514);
nor U1596 (N_1596,N_1550,N_1518);
nand U1597 (N_1597,N_1559,N_1546);
or U1598 (N_1598,N_1545,N_1553);
xor U1599 (N_1599,N_1502,N_1537);
or U1600 (N_1600,N_1523,N_1546);
nor U1601 (N_1601,N_1514,N_1519);
nor U1602 (N_1602,N_1527,N_1540);
nand U1603 (N_1603,N_1526,N_1508);
and U1604 (N_1604,N_1543,N_1528);
and U1605 (N_1605,N_1549,N_1556);
xnor U1606 (N_1606,N_1534,N_1527);
or U1607 (N_1607,N_1533,N_1534);
nand U1608 (N_1608,N_1539,N_1526);
and U1609 (N_1609,N_1522,N_1512);
or U1610 (N_1610,N_1500,N_1559);
or U1611 (N_1611,N_1557,N_1544);
nand U1612 (N_1612,N_1504,N_1512);
or U1613 (N_1613,N_1544,N_1545);
or U1614 (N_1614,N_1536,N_1502);
or U1615 (N_1615,N_1516,N_1533);
nor U1616 (N_1616,N_1528,N_1550);
xnor U1617 (N_1617,N_1506,N_1517);
nor U1618 (N_1618,N_1506,N_1512);
and U1619 (N_1619,N_1555,N_1532);
and U1620 (N_1620,N_1586,N_1588);
and U1621 (N_1621,N_1580,N_1611);
or U1622 (N_1622,N_1608,N_1592);
nand U1623 (N_1623,N_1615,N_1603);
nor U1624 (N_1624,N_1571,N_1597);
nand U1625 (N_1625,N_1564,N_1619);
nor U1626 (N_1626,N_1617,N_1563);
or U1627 (N_1627,N_1593,N_1589);
and U1628 (N_1628,N_1587,N_1567);
xor U1629 (N_1629,N_1604,N_1577);
nor U1630 (N_1630,N_1596,N_1618);
nor U1631 (N_1631,N_1606,N_1560);
or U1632 (N_1632,N_1612,N_1610);
nor U1633 (N_1633,N_1585,N_1590);
nand U1634 (N_1634,N_1566,N_1572);
or U1635 (N_1635,N_1583,N_1562);
nor U1636 (N_1636,N_1574,N_1599);
nor U1637 (N_1637,N_1600,N_1576);
and U1638 (N_1638,N_1565,N_1578);
nand U1639 (N_1639,N_1605,N_1601);
and U1640 (N_1640,N_1602,N_1609);
xor U1641 (N_1641,N_1568,N_1614);
and U1642 (N_1642,N_1613,N_1616);
and U1643 (N_1643,N_1573,N_1584);
xnor U1644 (N_1644,N_1579,N_1570);
or U1645 (N_1645,N_1598,N_1581);
nand U1646 (N_1646,N_1607,N_1594);
and U1647 (N_1647,N_1575,N_1591);
or U1648 (N_1648,N_1561,N_1569);
nor U1649 (N_1649,N_1595,N_1582);
nand U1650 (N_1650,N_1618,N_1567);
nand U1651 (N_1651,N_1574,N_1565);
nand U1652 (N_1652,N_1588,N_1594);
nand U1653 (N_1653,N_1583,N_1590);
nand U1654 (N_1654,N_1569,N_1578);
or U1655 (N_1655,N_1605,N_1616);
or U1656 (N_1656,N_1604,N_1568);
nand U1657 (N_1657,N_1561,N_1606);
and U1658 (N_1658,N_1571,N_1567);
nand U1659 (N_1659,N_1570,N_1617);
and U1660 (N_1660,N_1607,N_1578);
nor U1661 (N_1661,N_1561,N_1605);
nand U1662 (N_1662,N_1566,N_1583);
nand U1663 (N_1663,N_1611,N_1585);
nor U1664 (N_1664,N_1587,N_1581);
nand U1665 (N_1665,N_1608,N_1614);
and U1666 (N_1666,N_1576,N_1569);
nor U1667 (N_1667,N_1586,N_1591);
nand U1668 (N_1668,N_1564,N_1585);
or U1669 (N_1669,N_1615,N_1613);
nand U1670 (N_1670,N_1565,N_1571);
nand U1671 (N_1671,N_1580,N_1612);
xnor U1672 (N_1672,N_1581,N_1616);
nand U1673 (N_1673,N_1582,N_1579);
nand U1674 (N_1674,N_1565,N_1585);
or U1675 (N_1675,N_1582,N_1616);
nor U1676 (N_1676,N_1560,N_1590);
nor U1677 (N_1677,N_1593,N_1561);
nand U1678 (N_1678,N_1617,N_1593);
xor U1679 (N_1679,N_1598,N_1611);
and U1680 (N_1680,N_1675,N_1659);
or U1681 (N_1681,N_1629,N_1674);
and U1682 (N_1682,N_1624,N_1648);
or U1683 (N_1683,N_1670,N_1637);
nand U1684 (N_1684,N_1655,N_1651);
nand U1685 (N_1685,N_1625,N_1667);
and U1686 (N_1686,N_1638,N_1644);
or U1687 (N_1687,N_1633,N_1669);
nor U1688 (N_1688,N_1631,N_1650);
and U1689 (N_1689,N_1623,N_1656);
and U1690 (N_1690,N_1635,N_1672);
and U1691 (N_1691,N_1643,N_1661);
xor U1692 (N_1692,N_1627,N_1630);
nor U1693 (N_1693,N_1658,N_1634);
or U1694 (N_1694,N_1636,N_1646);
xnor U1695 (N_1695,N_1673,N_1632);
and U1696 (N_1696,N_1671,N_1641);
and U1697 (N_1697,N_1626,N_1657);
xor U1698 (N_1698,N_1677,N_1663);
and U1699 (N_1699,N_1679,N_1642);
nor U1700 (N_1700,N_1647,N_1628);
nand U1701 (N_1701,N_1640,N_1662);
nand U1702 (N_1702,N_1654,N_1653);
and U1703 (N_1703,N_1666,N_1660);
xnor U1704 (N_1704,N_1621,N_1620);
or U1705 (N_1705,N_1678,N_1649);
and U1706 (N_1706,N_1668,N_1639);
and U1707 (N_1707,N_1665,N_1664);
nand U1708 (N_1708,N_1652,N_1622);
nand U1709 (N_1709,N_1645,N_1676);
or U1710 (N_1710,N_1668,N_1620);
nand U1711 (N_1711,N_1637,N_1663);
nor U1712 (N_1712,N_1629,N_1662);
nor U1713 (N_1713,N_1635,N_1649);
xnor U1714 (N_1714,N_1679,N_1636);
nand U1715 (N_1715,N_1654,N_1656);
nor U1716 (N_1716,N_1678,N_1651);
nand U1717 (N_1717,N_1648,N_1655);
and U1718 (N_1718,N_1645,N_1667);
nand U1719 (N_1719,N_1631,N_1638);
or U1720 (N_1720,N_1673,N_1650);
nor U1721 (N_1721,N_1644,N_1673);
nor U1722 (N_1722,N_1631,N_1633);
and U1723 (N_1723,N_1674,N_1640);
and U1724 (N_1724,N_1671,N_1656);
or U1725 (N_1725,N_1655,N_1644);
nor U1726 (N_1726,N_1668,N_1657);
and U1727 (N_1727,N_1679,N_1634);
and U1728 (N_1728,N_1655,N_1662);
nand U1729 (N_1729,N_1626,N_1676);
or U1730 (N_1730,N_1635,N_1640);
nand U1731 (N_1731,N_1624,N_1646);
nand U1732 (N_1732,N_1636,N_1641);
xnor U1733 (N_1733,N_1667,N_1649);
nand U1734 (N_1734,N_1669,N_1674);
nand U1735 (N_1735,N_1632,N_1645);
nor U1736 (N_1736,N_1621,N_1624);
nand U1737 (N_1737,N_1639,N_1674);
or U1738 (N_1738,N_1627,N_1640);
nand U1739 (N_1739,N_1670,N_1641);
nand U1740 (N_1740,N_1701,N_1733);
or U1741 (N_1741,N_1727,N_1687);
or U1742 (N_1742,N_1717,N_1681);
or U1743 (N_1743,N_1730,N_1715);
and U1744 (N_1744,N_1697,N_1724);
xor U1745 (N_1745,N_1707,N_1692);
or U1746 (N_1746,N_1722,N_1738);
nand U1747 (N_1747,N_1709,N_1739);
or U1748 (N_1748,N_1699,N_1682);
and U1749 (N_1749,N_1736,N_1685);
and U1750 (N_1750,N_1686,N_1710);
nand U1751 (N_1751,N_1696,N_1728);
or U1752 (N_1752,N_1691,N_1693);
xor U1753 (N_1753,N_1731,N_1725);
and U1754 (N_1754,N_1689,N_1700);
nand U1755 (N_1755,N_1737,N_1713);
xnor U1756 (N_1756,N_1698,N_1723);
nor U1757 (N_1757,N_1694,N_1708);
or U1758 (N_1758,N_1719,N_1680);
nor U1759 (N_1759,N_1688,N_1712);
and U1760 (N_1760,N_1732,N_1703);
nor U1761 (N_1761,N_1705,N_1695);
xor U1762 (N_1762,N_1711,N_1706);
nor U1763 (N_1763,N_1716,N_1683);
or U1764 (N_1764,N_1714,N_1735);
xor U1765 (N_1765,N_1718,N_1690);
nor U1766 (N_1766,N_1704,N_1729);
and U1767 (N_1767,N_1720,N_1734);
and U1768 (N_1768,N_1721,N_1702);
and U1769 (N_1769,N_1726,N_1684);
or U1770 (N_1770,N_1685,N_1727);
xnor U1771 (N_1771,N_1732,N_1724);
nand U1772 (N_1772,N_1692,N_1721);
xor U1773 (N_1773,N_1680,N_1732);
nor U1774 (N_1774,N_1697,N_1716);
or U1775 (N_1775,N_1697,N_1738);
nand U1776 (N_1776,N_1736,N_1712);
nor U1777 (N_1777,N_1730,N_1729);
nand U1778 (N_1778,N_1703,N_1721);
and U1779 (N_1779,N_1697,N_1704);
nand U1780 (N_1780,N_1736,N_1739);
nand U1781 (N_1781,N_1717,N_1707);
nor U1782 (N_1782,N_1708,N_1722);
xor U1783 (N_1783,N_1717,N_1718);
and U1784 (N_1784,N_1705,N_1734);
and U1785 (N_1785,N_1730,N_1698);
or U1786 (N_1786,N_1735,N_1712);
nor U1787 (N_1787,N_1701,N_1692);
nand U1788 (N_1788,N_1718,N_1713);
nand U1789 (N_1789,N_1700,N_1709);
nor U1790 (N_1790,N_1722,N_1731);
nor U1791 (N_1791,N_1695,N_1716);
xor U1792 (N_1792,N_1718,N_1730);
and U1793 (N_1793,N_1702,N_1685);
nand U1794 (N_1794,N_1739,N_1735);
and U1795 (N_1795,N_1738,N_1708);
or U1796 (N_1796,N_1714,N_1736);
and U1797 (N_1797,N_1684,N_1728);
and U1798 (N_1798,N_1693,N_1736);
nor U1799 (N_1799,N_1698,N_1734);
or U1800 (N_1800,N_1779,N_1752);
nor U1801 (N_1801,N_1792,N_1780);
and U1802 (N_1802,N_1748,N_1795);
or U1803 (N_1803,N_1789,N_1761);
and U1804 (N_1804,N_1778,N_1767);
xnor U1805 (N_1805,N_1753,N_1770);
nand U1806 (N_1806,N_1783,N_1786);
nand U1807 (N_1807,N_1790,N_1762);
nor U1808 (N_1808,N_1776,N_1746);
nor U1809 (N_1809,N_1798,N_1757);
nand U1810 (N_1810,N_1774,N_1797);
xor U1811 (N_1811,N_1799,N_1787);
nand U1812 (N_1812,N_1766,N_1754);
xor U1813 (N_1813,N_1743,N_1744);
and U1814 (N_1814,N_1788,N_1759);
nor U1815 (N_1815,N_1760,N_1771);
nor U1816 (N_1816,N_1769,N_1796);
or U1817 (N_1817,N_1747,N_1742);
and U1818 (N_1818,N_1750,N_1765);
nand U1819 (N_1819,N_1741,N_1749);
and U1820 (N_1820,N_1758,N_1785);
nor U1821 (N_1821,N_1756,N_1781);
and U1822 (N_1822,N_1782,N_1793);
and U1823 (N_1823,N_1740,N_1794);
nand U1824 (N_1824,N_1775,N_1745);
or U1825 (N_1825,N_1755,N_1773);
nand U1826 (N_1826,N_1777,N_1751);
xnor U1827 (N_1827,N_1784,N_1763);
or U1828 (N_1828,N_1772,N_1791);
and U1829 (N_1829,N_1768,N_1764);
nor U1830 (N_1830,N_1773,N_1792);
nor U1831 (N_1831,N_1788,N_1799);
nor U1832 (N_1832,N_1776,N_1741);
and U1833 (N_1833,N_1778,N_1744);
and U1834 (N_1834,N_1789,N_1771);
and U1835 (N_1835,N_1756,N_1772);
xnor U1836 (N_1836,N_1757,N_1773);
and U1837 (N_1837,N_1750,N_1773);
xnor U1838 (N_1838,N_1766,N_1789);
or U1839 (N_1839,N_1750,N_1777);
and U1840 (N_1840,N_1765,N_1793);
xor U1841 (N_1841,N_1756,N_1755);
xor U1842 (N_1842,N_1794,N_1752);
xor U1843 (N_1843,N_1766,N_1740);
and U1844 (N_1844,N_1744,N_1768);
nor U1845 (N_1845,N_1773,N_1780);
and U1846 (N_1846,N_1749,N_1799);
nor U1847 (N_1847,N_1760,N_1791);
nor U1848 (N_1848,N_1779,N_1791);
or U1849 (N_1849,N_1780,N_1759);
nand U1850 (N_1850,N_1778,N_1795);
or U1851 (N_1851,N_1779,N_1756);
nor U1852 (N_1852,N_1770,N_1747);
or U1853 (N_1853,N_1782,N_1742);
and U1854 (N_1854,N_1758,N_1781);
nor U1855 (N_1855,N_1774,N_1795);
nor U1856 (N_1856,N_1773,N_1782);
nand U1857 (N_1857,N_1751,N_1744);
and U1858 (N_1858,N_1744,N_1790);
and U1859 (N_1859,N_1770,N_1743);
or U1860 (N_1860,N_1808,N_1835);
xor U1861 (N_1861,N_1816,N_1833);
and U1862 (N_1862,N_1836,N_1850);
nand U1863 (N_1863,N_1831,N_1814);
xor U1864 (N_1864,N_1834,N_1807);
nor U1865 (N_1865,N_1825,N_1855);
and U1866 (N_1866,N_1819,N_1846);
nor U1867 (N_1867,N_1815,N_1854);
nand U1868 (N_1868,N_1820,N_1811);
or U1869 (N_1869,N_1847,N_1822);
nand U1870 (N_1870,N_1824,N_1841);
nand U1871 (N_1871,N_1828,N_1826);
or U1872 (N_1872,N_1842,N_1801);
nor U1873 (N_1873,N_1856,N_1803);
and U1874 (N_1874,N_1817,N_1821);
and U1875 (N_1875,N_1818,N_1857);
nand U1876 (N_1876,N_1838,N_1853);
or U1877 (N_1877,N_1851,N_1802);
nor U1878 (N_1878,N_1813,N_1810);
or U1879 (N_1879,N_1804,N_1830);
or U1880 (N_1880,N_1840,N_1845);
nor U1881 (N_1881,N_1843,N_1844);
xor U1882 (N_1882,N_1827,N_1806);
nand U1883 (N_1883,N_1812,N_1837);
or U1884 (N_1884,N_1829,N_1805);
xnor U1885 (N_1885,N_1848,N_1832);
nand U1886 (N_1886,N_1823,N_1800);
nand U1887 (N_1887,N_1809,N_1839);
and U1888 (N_1888,N_1852,N_1859);
nand U1889 (N_1889,N_1849,N_1858);
nor U1890 (N_1890,N_1832,N_1843);
or U1891 (N_1891,N_1845,N_1819);
xnor U1892 (N_1892,N_1826,N_1804);
or U1893 (N_1893,N_1851,N_1855);
or U1894 (N_1894,N_1841,N_1817);
nand U1895 (N_1895,N_1811,N_1816);
nand U1896 (N_1896,N_1816,N_1857);
nand U1897 (N_1897,N_1834,N_1857);
or U1898 (N_1898,N_1818,N_1842);
or U1899 (N_1899,N_1833,N_1830);
nand U1900 (N_1900,N_1821,N_1825);
and U1901 (N_1901,N_1837,N_1830);
nor U1902 (N_1902,N_1832,N_1807);
or U1903 (N_1903,N_1832,N_1823);
nor U1904 (N_1904,N_1858,N_1852);
nand U1905 (N_1905,N_1807,N_1804);
nor U1906 (N_1906,N_1809,N_1859);
nand U1907 (N_1907,N_1802,N_1808);
nor U1908 (N_1908,N_1829,N_1801);
xor U1909 (N_1909,N_1857,N_1819);
nand U1910 (N_1910,N_1848,N_1807);
xor U1911 (N_1911,N_1839,N_1820);
nand U1912 (N_1912,N_1814,N_1823);
nor U1913 (N_1913,N_1845,N_1830);
nand U1914 (N_1914,N_1848,N_1839);
and U1915 (N_1915,N_1802,N_1813);
nor U1916 (N_1916,N_1803,N_1817);
nor U1917 (N_1917,N_1851,N_1858);
and U1918 (N_1918,N_1820,N_1854);
nor U1919 (N_1919,N_1846,N_1839);
xor U1920 (N_1920,N_1910,N_1873);
and U1921 (N_1921,N_1862,N_1880);
or U1922 (N_1922,N_1885,N_1915);
nor U1923 (N_1923,N_1906,N_1893);
nor U1924 (N_1924,N_1913,N_1874);
nand U1925 (N_1925,N_1869,N_1914);
or U1926 (N_1926,N_1909,N_1875);
and U1927 (N_1927,N_1877,N_1898);
nor U1928 (N_1928,N_1878,N_1908);
nor U1929 (N_1929,N_1882,N_1871);
nor U1930 (N_1930,N_1891,N_1865);
and U1931 (N_1931,N_1870,N_1881);
and U1932 (N_1932,N_1905,N_1884);
and U1933 (N_1933,N_1868,N_1867);
and U1934 (N_1934,N_1864,N_1911);
and U1935 (N_1935,N_1916,N_1907);
xnor U1936 (N_1936,N_1903,N_1894);
nor U1937 (N_1937,N_1902,N_1861);
nor U1938 (N_1938,N_1899,N_1888);
and U1939 (N_1939,N_1887,N_1912);
nand U1940 (N_1940,N_1901,N_1863);
xor U1941 (N_1941,N_1918,N_1879);
nor U1942 (N_1942,N_1897,N_1904);
xnor U1943 (N_1943,N_1866,N_1900);
nor U1944 (N_1944,N_1889,N_1895);
nand U1945 (N_1945,N_1883,N_1860);
nand U1946 (N_1946,N_1919,N_1886);
or U1947 (N_1947,N_1890,N_1917);
nand U1948 (N_1948,N_1876,N_1872);
nand U1949 (N_1949,N_1896,N_1892);
nor U1950 (N_1950,N_1876,N_1869);
nand U1951 (N_1951,N_1900,N_1895);
and U1952 (N_1952,N_1868,N_1917);
or U1953 (N_1953,N_1914,N_1874);
and U1954 (N_1954,N_1891,N_1880);
and U1955 (N_1955,N_1908,N_1865);
nor U1956 (N_1956,N_1903,N_1871);
nand U1957 (N_1957,N_1884,N_1890);
nand U1958 (N_1958,N_1897,N_1878);
nor U1959 (N_1959,N_1874,N_1907);
and U1960 (N_1960,N_1901,N_1878);
nor U1961 (N_1961,N_1893,N_1888);
nor U1962 (N_1962,N_1910,N_1913);
and U1963 (N_1963,N_1894,N_1868);
and U1964 (N_1964,N_1919,N_1870);
and U1965 (N_1965,N_1908,N_1899);
nand U1966 (N_1966,N_1880,N_1904);
nand U1967 (N_1967,N_1883,N_1892);
or U1968 (N_1968,N_1876,N_1902);
xor U1969 (N_1969,N_1913,N_1903);
and U1970 (N_1970,N_1899,N_1868);
and U1971 (N_1971,N_1900,N_1884);
xnor U1972 (N_1972,N_1917,N_1881);
and U1973 (N_1973,N_1860,N_1889);
nand U1974 (N_1974,N_1916,N_1908);
and U1975 (N_1975,N_1874,N_1911);
and U1976 (N_1976,N_1881,N_1905);
and U1977 (N_1977,N_1887,N_1916);
nand U1978 (N_1978,N_1872,N_1881);
and U1979 (N_1979,N_1905,N_1894);
nor U1980 (N_1980,N_1971,N_1963);
xnor U1981 (N_1981,N_1952,N_1935);
or U1982 (N_1982,N_1979,N_1967);
nand U1983 (N_1983,N_1946,N_1932);
nand U1984 (N_1984,N_1944,N_1973);
nand U1985 (N_1985,N_1947,N_1942);
and U1986 (N_1986,N_1941,N_1931);
nor U1987 (N_1987,N_1970,N_1927);
or U1988 (N_1988,N_1958,N_1969);
or U1989 (N_1989,N_1933,N_1928);
or U1990 (N_1990,N_1976,N_1930);
nand U1991 (N_1991,N_1925,N_1968);
nor U1992 (N_1992,N_1950,N_1951);
nor U1993 (N_1993,N_1953,N_1923);
or U1994 (N_1994,N_1964,N_1978);
and U1995 (N_1995,N_1977,N_1948);
nor U1996 (N_1996,N_1962,N_1939);
and U1997 (N_1997,N_1960,N_1966);
and U1998 (N_1998,N_1921,N_1972);
nand U1999 (N_1999,N_1922,N_1924);
or U2000 (N_2000,N_1920,N_1926);
nand U2001 (N_2001,N_1965,N_1957);
nor U2002 (N_2002,N_1934,N_1940);
or U2003 (N_2003,N_1945,N_1961);
nand U2004 (N_2004,N_1943,N_1936);
or U2005 (N_2005,N_1949,N_1959);
nand U2006 (N_2006,N_1929,N_1937);
or U2007 (N_2007,N_1938,N_1956);
or U2008 (N_2008,N_1954,N_1955);
and U2009 (N_2009,N_1974,N_1975);
nand U2010 (N_2010,N_1923,N_1926);
nand U2011 (N_2011,N_1951,N_1942);
nor U2012 (N_2012,N_1946,N_1929);
and U2013 (N_2013,N_1943,N_1975);
xnor U2014 (N_2014,N_1936,N_1945);
or U2015 (N_2015,N_1926,N_1953);
nand U2016 (N_2016,N_1970,N_1954);
nor U2017 (N_2017,N_1936,N_1976);
nor U2018 (N_2018,N_1942,N_1979);
and U2019 (N_2019,N_1924,N_1965);
nor U2020 (N_2020,N_1926,N_1934);
xnor U2021 (N_2021,N_1950,N_1923);
and U2022 (N_2022,N_1943,N_1965);
nor U2023 (N_2023,N_1962,N_1977);
or U2024 (N_2024,N_1967,N_1945);
nor U2025 (N_2025,N_1948,N_1961);
and U2026 (N_2026,N_1958,N_1932);
xnor U2027 (N_2027,N_1928,N_1955);
and U2028 (N_2028,N_1942,N_1949);
nand U2029 (N_2029,N_1925,N_1951);
nor U2030 (N_2030,N_1959,N_1950);
nor U2031 (N_2031,N_1943,N_1962);
and U2032 (N_2032,N_1967,N_1949);
nor U2033 (N_2033,N_1972,N_1957);
nand U2034 (N_2034,N_1956,N_1947);
nand U2035 (N_2035,N_1922,N_1943);
nand U2036 (N_2036,N_1935,N_1940);
or U2037 (N_2037,N_1957,N_1945);
and U2038 (N_2038,N_1951,N_1939);
nand U2039 (N_2039,N_1950,N_1967);
xnor U2040 (N_2040,N_2029,N_1981);
or U2041 (N_2041,N_2017,N_2007);
nor U2042 (N_2042,N_1998,N_2003);
nor U2043 (N_2043,N_2005,N_2015);
nand U2044 (N_2044,N_2018,N_2036);
and U2045 (N_2045,N_2027,N_2034);
or U2046 (N_2046,N_2013,N_2024);
nand U2047 (N_2047,N_2016,N_2025);
nor U2048 (N_2048,N_2012,N_1980);
or U2049 (N_2049,N_1996,N_2008);
nand U2050 (N_2050,N_2023,N_2019);
xor U2051 (N_2051,N_2037,N_2028);
and U2052 (N_2052,N_1999,N_2010);
nor U2053 (N_2053,N_2038,N_2004);
and U2054 (N_2054,N_1989,N_1983);
nand U2055 (N_2055,N_2009,N_2035);
and U2056 (N_2056,N_1990,N_2021);
or U2057 (N_2057,N_1984,N_2006);
nand U2058 (N_2058,N_2033,N_2011);
or U2059 (N_2059,N_2002,N_2020);
or U2060 (N_2060,N_1997,N_2000);
or U2061 (N_2061,N_1986,N_1995);
or U2062 (N_2062,N_1987,N_1994);
nand U2063 (N_2063,N_2031,N_1991);
nor U2064 (N_2064,N_1993,N_1988);
nand U2065 (N_2065,N_2026,N_2014);
or U2066 (N_2066,N_2022,N_2030);
nand U2067 (N_2067,N_2001,N_2032);
or U2068 (N_2068,N_2039,N_1985);
and U2069 (N_2069,N_1982,N_1992);
or U2070 (N_2070,N_1986,N_2034);
nor U2071 (N_2071,N_2033,N_1999);
nor U2072 (N_2072,N_1992,N_2012);
or U2073 (N_2073,N_2016,N_2024);
or U2074 (N_2074,N_2037,N_2023);
and U2075 (N_2075,N_1988,N_2029);
nand U2076 (N_2076,N_2009,N_2024);
or U2077 (N_2077,N_1980,N_1984);
and U2078 (N_2078,N_2011,N_2034);
nor U2079 (N_2079,N_1990,N_1995);
and U2080 (N_2080,N_2025,N_2003);
nand U2081 (N_2081,N_2025,N_2039);
nand U2082 (N_2082,N_2014,N_2032);
and U2083 (N_2083,N_2006,N_2027);
and U2084 (N_2084,N_1983,N_2025);
xnor U2085 (N_2085,N_1997,N_2019);
and U2086 (N_2086,N_2024,N_2021);
xor U2087 (N_2087,N_2024,N_1982);
nand U2088 (N_2088,N_2034,N_1998);
or U2089 (N_2089,N_2003,N_1985);
xor U2090 (N_2090,N_2002,N_2026);
nor U2091 (N_2091,N_1986,N_2015);
nor U2092 (N_2092,N_2038,N_1994);
xor U2093 (N_2093,N_2025,N_1980);
nor U2094 (N_2094,N_1983,N_2011);
nor U2095 (N_2095,N_2000,N_2006);
or U2096 (N_2096,N_2003,N_2019);
or U2097 (N_2097,N_2012,N_2032);
nor U2098 (N_2098,N_1993,N_2001);
nand U2099 (N_2099,N_2035,N_2034);
nand U2100 (N_2100,N_2040,N_2043);
xor U2101 (N_2101,N_2070,N_2076);
nand U2102 (N_2102,N_2056,N_2051);
nor U2103 (N_2103,N_2057,N_2074);
or U2104 (N_2104,N_2071,N_2068);
or U2105 (N_2105,N_2058,N_2088);
and U2106 (N_2106,N_2097,N_2045);
and U2107 (N_2107,N_2087,N_2080);
or U2108 (N_2108,N_2072,N_2093);
nand U2109 (N_2109,N_2098,N_2089);
or U2110 (N_2110,N_2084,N_2044);
and U2111 (N_2111,N_2047,N_2082);
nand U2112 (N_2112,N_2063,N_2050);
xor U2113 (N_2113,N_2095,N_2086);
nor U2114 (N_2114,N_2055,N_2090);
or U2115 (N_2115,N_2061,N_2099);
nor U2116 (N_2116,N_2060,N_2062);
nand U2117 (N_2117,N_2052,N_2064);
nand U2118 (N_2118,N_2077,N_2065);
or U2119 (N_2119,N_2083,N_2079);
or U2120 (N_2120,N_2066,N_2073);
xor U2121 (N_2121,N_2094,N_2096);
nor U2122 (N_2122,N_2053,N_2092);
xnor U2123 (N_2123,N_2048,N_2041);
nand U2124 (N_2124,N_2042,N_2067);
and U2125 (N_2125,N_2091,N_2046);
or U2126 (N_2126,N_2075,N_2054);
nand U2127 (N_2127,N_2078,N_2081);
nor U2128 (N_2128,N_2069,N_2049);
or U2129 (N_2129,N_2059,N_2085);
nor U2130 (N_2130,N_2067,N_2089);
xnor U2131 (N_2131,N_2051,N_2049);
and U2132 (N_2132,N_2081,N_2066);
nor U2133 (N_2133,N_2080,N_2055);
nor U2134 (N_2134,N_2087,N_2047);
or U2135 (N_2135,N_2085,N_2078);
and U2136 (N_2136,N_2046,N_2075);
nor U2137 (N_2137,N_2086,N_2077);
nand U2138 (N_2138,N_2086,N_2070);
nand U2139 (N_2139,N_2085,N_2080);
and U2140 (N_2140,N_2072,N_2092);
and U2141 (N_2141,N_2053,N_2099);
and U2142 (N_2142,N_2052,N_2042);
or U2143 (N_2143,N_2083,N_2075);
xnor U2144 (N_2144,N_2065,N_2055);
and U2145 (N_2145,N_2090,N_2094);
and U2146 (N_2146,N_2042,N_2073);
nand U2147 (N_2147,N_2061,N_2052);
nor U2148 (N_2148,N_2095,N_2053);
or U2149 (N_2149,N_2068,N_2091);
and U2150 (N_2150,N_2094,N_2085);
and U2151 (N_2151,N_2042,N_2098);
or U2152 (N_2152,N_2050,N_2067);
and U2153 (N_2153,N_2057,N_2045);
nor U2154 (N_2154,N_2076,N_2079);
nand U2155 (N_2155,N_2051,N_2087);
and U2156 (N_2156,N_2072,N_2067);
nor U2157 (N_2157,N_2094,N_2044);
and U2158 (N_2158,N_2063,N_2047);
and U2159 (N_2159,N_2066,N_2068);
or U2160 (N_2160,N_2105,N_2100);
nand U2161 (N_2161,N_2140,N_2159);
and U2162 (N_2162,N_2109,N_2108);
and U2163 (N_2163,N_2154,N_2143);
or U2164 (N_2164,N_2133,N_2128);
nand U2165 (N_2165,N_2148,N_2146);
nand U2166 (N_2166,N_2135,N_2149);
or U2167 (N_2167,N_2104,N_2145);
and U2168 (N_2168,N_2119,N_2147);
nand U2169 (N_2169,N_2117,N_2125);
or U2170 (N_2170,N_2120,N_2102);
or U2171 (N_2171,N_2153,N_2121);
and U2172 (N_2172,N_2113,N_2107);
nand U2173 (N_2173,N_2126,N_2112);
and U2174 (N_2174,N_2101,N_2142);
nand U2175 (N_2175,N_2118,N_2139);
nor U2176 (N_2176,N_2103,N_2131);
nand U2177 (N_2177,N_2137,N_2132);
nand U2178 (N_2178,N_2130,N_2134);
or U2179 (N_2179,N_2136,N_2138);
nand U2180 (N_2180,N_2157,N_2150);
nor U2181 (N_2181,N_2155,N_2144);
nand U2182 (N_2182,N_2110,N_2111);
xor U2183 (N_2183,N_2124,N_2127);
or U2184 (N_2184,N_2116,N_2151);
or U2185 (N_2185,N_2106,N_2152);
and U2186 (N_2186,N_2115,N_2123);
nor U2187 (N_2187,N_2158,N_2141);
nor U2188 (N_2188,N_2129,N_2122);
and U2189 (N_2189,N_2156,N_2114);
xor U2190 (N_2190,N_2103,N_2141);
and U2191 (N_2191,N_2148,N_2149);
or U2192 (N_2192,N_2144,N_2124);
nor U2193 (N_2193,N_2102,N_2129);
and U2194 (N_2194,N_2145,N_2158);
nand U2195 (N_2195,N_2115,N_2134);
nor U2196 (N_2196,N_2131,N_2141);
xor U2197 (N_2197,N_2141,N_2101);
or U2198 (N_2198,N_2112,N_2139);
nand U2199 (N_2199,N_2128,N_2114);
xnor U2200 (N_2200,N_2159,N_2152);
and U2201 (N_2201,N_2105,N_2137);
nor U2202 (N_2202,N_2107,N_2106);
nand U2203 (N_2203,N_2123,N_2127);
or U2204 (N_2204,N_2108,N_2122);
xnor U2205 (N_2205,N_2140,N_2116);
nand U2206 (N_2206,N_2126,N_2159);
nor U2207 (N_2207,N_2102,N_2147);
nand U2208 (N_2208,N_2121,N_2124);
nor U2209 (N_2209,N_2145,N_2125);
and U2210 (N_2210,N_2159,N_2119);
nand U2211 (N_2211,N_2133,N_2132);
xnor U2212 (N_2212,N_2122,N_2132);
nor U2213 (N_2213,N_2122,N_2110);
nor U2214 (N_2214,N_2109,N_2113);
nor U2215 (N_2215,N_2158,N_2146);
or U2216 (N_2216,N_2149,N_2145);
and U2217 (N_2217,N_2147,N_2127);
nand U2218 (N_2218,N_2127,N_2139);
nand U2219 (N_2219,N_2154,N_2102);
or U2220 (N_2220,N_2205,N_2176);
nand U2221 (N_2221,N_2165,N_2187);
and U2222 (N_2222,N_2173,N_2164);
nand U2223 (N_2223,N_2195,N_2166);
or U2224 (N_2224,N_2183,N_2168);
nor U2225 (N_2225,N_2215,N_2177);
or U2226 (N_2226,N_2161,N_2206);
and U2227 (N_2227,N_2210,N_2180);
or U2228 (N_2228,N_2171,N_2217);
nand U2229 (N_2229,N_2208,N_2169);
nand U2230 (N_2230,N_2209,N_2197);
xnor U2231 (N_2231,N_2181,N_2213);
and U2232 (N_2232,N_2179,N_2200);
nand U2233 (N_2233,N_2216,N_2184);
and U2234 (N_2234,N_2174,N_2193);
nand U2235 (N_2235,N_2212,N_2198);
and U2236 (N_2236,N_2218,N_2194);
nor U2237 (N_2237,N_2182,N_2178);
or U2238 (N_2238,N_2162,N_2167);
nand U2239 (N_2239,N_2219,N_2202);
nor U2240 (N_2240,N_2190,N_2191);
or U2241 (N_2241,N_2186,N_2211);
and U2242 (N_2242,N_2207,N_2204);
and U2243 (N_2243,N_2196,N_2203);
nand U2244 (N_2244,N_2214,N_2163);
nor U2245 (N_2245,N_2189,N_2199);
or U2246 (N_2246,N_2172,N_2192);
nand U2247 (N_2247,N_2201,N_2188);
xor U2248 (N_2248,N_2175,N_2185);
and U2249 (N_2249,N_2160,N_2170);
nor U2250 (N_2250,N_2204,N_2182);
nand U2251 (N_2251,N_2209,N_2167);
and U2252 (N_2252,N_2190,N_2162);
and U2253 (N_2253,N_2175,N_2164);
and U2254 (N_2254,N_2215,N_2167);
or U2255 (N_2255,N_2199,N_2194);
or U2256 (N_2256,N_2181,N_2170);
xor U2257 (N_2257,N_2160,N_2184);
or U2258 (N_2258,N_2202,N_2217);
and U2259 (N_2259,N_2169,N_2191);
or U2260 (N_2260,N_2163,N_2160);
or U2261 (N_2261,N_2206,N_2179);
or U2262 (N_2262,N_2206,N_2164);
xor U2263 (N_2263,N_2174,N_2204);
or U2264 (N_2264,N_2193,N_2216);
and U2265 (N_2265,N_2186,N_2191);
xnor U2266 (N_2266,N_2181,N_2194);
nand U2267 (N_2267,N_2195,N_2176);
or U2268 (N_2268,N_2162,N_2188);
nand U2269 (N_2269,N_2202,N_2188);
nand U2270 (N_2270,N_2174,N_2207);
and U2271 (N_2271,N_2168,N_2182);
nor U2272 (N_2272,N_2180,N_2172);
nor U2273 (N_2273,N_2200,N_2161);
nand U2274 (N_2274,N_2201,N_2166);
nand U2275 (N_2275,N_2181,N_2203);
nor U2276 (N_2276,N_2198,N_2209);
and U2277 (N_2277,N_2211,N_2198);
nand U2278 (N_2278,N_2175,N_2176);
or U2279 (N_2279,N_2174,N_2164);
or U2280 (N_2280,N_2264,N_2234);
xor U2281 (N_2281,N_2222,N_2246);
nor U2282 (N_2282,N_2278,N_2261);
nand U2283 (N_2283,N_2263,N_2237);
or U2284 (N_2284,N_2274,N_2276);
and U2285 (N_2285,N_2271,N_2268);
and U2286 (N_2286,N_2241,N_2252);
and U2287 (N_2287,N_2227,N_2254);
nor U2288 (N_2288,N_2226,N_2250);
or U2289 (N_2289,N_2243,N_2231);
and U2290 (N_2290,N_2236,N_2251);
nor U2291 (N_2291,N_2228,N_2260);
nor U2292 (N_2292,N_2238,N_2223);
nand U2293 (N_2293,N_2258,N_2259);
nand U2294 (N_2294,N_2262,N_2242);
xnor U2295 (N_2295,N_2244,N_2267);
nand U2296 (N_2296,N_2249,N_2256);
nor U2297 (N_2297,N_2233,N_2277);
or U2298 (N_2298,N_2224,N_2229);
nand U2299 (N_2299,N_2240,N_2253);
nand U2300 (N_2300,N_2279,N_2272);
nand U2301 (N_2301,N_2273,N_2270);
nor U2302 (N_2302,N_2220,N_2269);
and U2303 (N_2303,N_2230,N_2232);
nand U2304 (N_2304,N_2255,N_2247);
nor U2305 (N_2305,N_2275,N_2221);
nor U2306 (N_2306,N_2257,N_2225);
and U2307 (N_2307,N_2266,N_2239);
nand U2308 (N_2308,N_2265,N_2248);
nor U2309 (N_2309,N_2245,N_2235);
nand U2310 (N_2310,N_2250,N_2235);
xnor U2311 (N_2311,N_2240,N_2252);
or U2312 (N_2312,N_2224,N_2258);
xor U2313 (N_2313,N_2257,N_2226);
and U2314 (N_2314,N_2269,N_2234);
nor U2315 (N_2315,N_2243,N_2220);
nand U2316 (N_2316,N_2235,N_2221);
and U2317 (N_2317,N_2225,N_2272);
or U2318 (N_2318,N_2247,N_2273);
and U2319 (N_2319,N_2273,N_2241);
and U2320 (N_2320,N_2242,N_2221);
nand U2321 (N_2321,N_2254,N_2251);
or U2322 (N_2322,N_2246,N_2250);
nand U2323 (N_2323,N_2237,N_2225);
or U2324 (N_2324,N_2246,N_2273);
or U2325 (N_2325,N_2240,N_2226);
and U2326 (N_2326,N_2270,N_2260);
nand U2327 (N_2327,N_2248,N_2225);
nor U2328 (N_2328,N_2228,N_2253);
nor U2329 (N_2329,N_2261,N_2245);
nor U2330 (N_2330,N_2270,N_2239);
and U2331 (N_2331,N_2237,N_2266);
and U2332 (N_2332,N_2243,N_2230);
and U2333 (N_2333,N_2250,N_2237);
and U2334 (N_2334,N_2226,N_2234);
nor U2335 (N_2335,N_2252,N_2265);
nor U2336 (N_2336,N_2259,N_2252);
and U2337 (N_2337,N_2264,N_2262);
xnor U2338 (N_2338,N_2260,N_2241);
nor U2339 (N_2339,N_2274,N_2267);
nand U2340 (N_2340,N_2329,N_2288);
and U2341 (N_2341,N_2318,N_2292);
or U2342 (N_2342,N_2337,N_2305);
or U2343 (N_2343,N_2334,N_2313);
nand U2344 (N_2344,N_2324,N_2332);
nand U2345 (N_2345,N_2336,N_2289);
and U2346 (N_2346,N_2287,N_2303);
nand U2347 (N_2347,N_2290,N_2322);
nor U2348 (N_2348,N_2309,N_2319);
nand U2349 (N_2349,N_2298,N_2302);
nand U2350 (N_2350,N_2304,N_2339);
nor U2351 (N_2351,N_2280,N_2284);
or U2352 (N_2352,N_2297,N_2328);
and U2353 (N_2353,N_2335,N_2312);
nand U2354 (N_2354,N_2301,N_2311);
nor U2355 (N_2355,N_2294,N_2295);
nor U2356 (N_2356,N_2300,N_2306);
and U2357 (N_2357,N_2281,N_2314);
nor U2358 (N_2358,N_2283,N_2327);
xnor U2359 (N_2359,N_2338,N_2296);
and U2360 (N_2360,N_2325,N_2323);
nand U2361 (N_2361,N_2321,N_2285);
and U2362 (N_2362,N_2315,N_2310);
nand U2363 (N_2363,N_2320,N_2316);
and U2364 (N_2364,N_2286,N_2317);
nor U2365 (N_2365,N_2333,N_2293);
nor U2366 (N_2366,N_2291,N_2299);
xnor U2367 (N_2367,N_2330,N_2331);
nand U2368 (N_2368,N_2308,N_2326);
and U2369 (N_2369,N_2307,N_2282);
nand U2370 (N_2370,N_2306,N_2325);
and U2371 (N_2371,N_2327,N_2321);
nand U2372 (N_2372,N_2289,N_2333);
nor U2373 (N_2373,N_2337,N_2333);
nor U2374 (N_2374,N_2290,N_2324);
nand U2375 (N_2375,N_2287,N_2331);
and U2376 (N_2376,N_2323,N_2294);
nor U2377 (N_2377,N_2316,N_2294);
and U2378 (N_2378,N_2313,N_2306);
nor U2379 (N_2379,N_2315,N_2316);
nor U2380 (N_2380,N_2299,N_2312);
nor U2381 (N_2381,N_2323,N_2330);
nand U2382 (N_2382,N_2329,N_2317);
and U2383 (N_2383,N_2302,N_2292);
nand U2384 (N_2384,N_2306,N_2290);
or U2385 (N_2385,N_2316,N_2285);
nand U2386 (N_2386,N_2319,N_2329);
and U2387 (N_2387,N_2308,N_2333);
and U2388 (N_2388,N_2337,N_2339);
or U2389 (N_2389,N_2285,N_2309);
or U2390 (N_2390,N_2300,N_2291);
nor U2391 (N_2391,N_2311,N_2334);
nor U2392 (N_2392,N_2299,N_2331);
and U2393 (N_2393,N_2325,N_2300);
nand U2394 (N_2394,N_2307,N_2333);
xnor U2395 (N_2395,N_2319,N_2289);
nor U2396 (N_2396,N_2289,N_2331);
nor U2397 (N_2397,N_2316,N_2292);
and U2398 (N_2398,N_2311,N_2338);
or U2399 (N_2399,N_2316,N_2322);
nor U2400 (N_2400,N_2379,N_2367);
xor U2401 (N_2401,N_2381,N_2393);
nand U2402 (N_2402,N_2360,N_2399);
nand U2403 (N_2403,N_2385,N_2342);
nand U2404 (N_2404,N_2387,N_2346);
or U2405 (N_2405,N_2372,N_2364);
or U2406 (N_2406,N_2340,N_2396);
and U2407 (N_2407,N_2370,N_2391);
nand U2408 (N_2408,N_2394,N_2350);
nor U2409 (N_2409,N_2369,N_2377);
xor U2410 (N_2410,N_2366,N_2352);
xor U2411 (N_2411,N_2395,N_2362);
or U2412 (N_2412,N_2398,N_2382);
nor U2413 (N_2413,N_2373,N_2392);
nand U2414 (N_2414,N_2371,N_2374);
and U2415 (N_2415,N_2365,N_2353);
nor U2416 (N_2416,N_2349,N_2368);
or U2417 (N_2417,N_2361,N_2344);
or U2418 (N_2418,N_2376,N_2348);
or U2419 (N_2419,N_2386,N_2390);
and U2420 (N_2420,N_2383,N_2389);
xnor U2421 (N_2421,N_2375,N_2341);
or U2422 (N_2422,N_2355,N_2351);
or U2423 (N_2423,N_2397,N_2358);
xnor U2424 (N_2424,N_2363,N_2357);
nand U2425 (N_2425,N_2378,N_2345);
nor U2426 (N_2426,N_2380,N_2384);
or U2427 (N_2427,N_2354,N_2347);
and U2428 (N_2428,N_2356,N_2388);
nand U2429 (N_2429,N_2343,N_2359);
nand U2430 (N_2430,N_2394,N_2360);
and U2431 (N_2431,N_2396,N_2398);
and U2432 (N_2432,N_2372,N_2388);
and U2433 (N_2433,N_2349,N_2378);
or U2434 (N_2434,N_2382,N_2385);
nor U2435 (N_2435,N_2348,N_2344);
and U2436 (N_2436,N_2347,N_2355);
nand U2437 (N_2437,N_2388,N_2381);
and U2438 (N_2438,N_2372,N_2379);
nand U2439 (N_2439,N_2384,N_2390);
and U2440 (N_2440,N_2379,N_2376);
and U2441 (N_2441,N_2389,N_2385);
nand U2442 (N_2442,N_2394,N_2382);
xnor U2443 (N_2443,N_2362,N_2342);
xor U2444 (N_2444,N_2367,N_2391);
nor U2445 (N_2445,N_2345,N_2362);
or U2446 (N_2446,N_2358,N_2344);
nor U2447 (N_2447,N_2352,N_2375);
and U2448 (N_2448,N_2371,N_2378);
nor U2449 (N_2449,N_2387,N_2383);
or U2450 (N_2450,N_2385,N_2391);
xor U2451 (N_2451,N_2363,N_2344);
nand U2452 (N_2452,N_2354,N_2369);
nor U2453 (N_2453,N_2389,N_2342);
nand U2454 (N_2454,N_2345,N_2387);
xor U2455 (N_2455,N_2386,N_2360);
xnor U2456 (N_2456,N_2349,N_2377);
nor U2457 (N_2457,N_2362,N_2393);
nor U2458 (N_2458,N_2384,N_2388);
nand U2459 (N_2459,N_2343,N_2355);
nor U2460 (N_2460,N_2449,N_2430);
nand U2461 (N_2461,N_2401,N_2408);
nand U2462 (N_2462,N_2419,N_2421);
nand U2463 (N_2463,N_2434,N_2433);
xor U2464 (N_2464,N_2446,N_2445);
and U2465 (N_2465,N_2428,N_2400);
xor U2466 (N_2466,N_2439,N_2432);
xor U2467 (N_2467,N_2431,N_2423);
or U2468 (N_2468,N_2457,N_2443);
and U2469 (N_2469,N_2453,N_2442);
nor U2470 (N_2470,N_2426,N_2436);
or U2471 (N_2471,N_2456,N_2410);
nor U2472 (N_2472,N_2407,N_2422);
and U2473 (N_2473,N_2403,N_2452);
nand U2474 (N_2474,N_2440,N_2404);
nand U2475 (N_2475,N_2458,N_2412);
xnor U2476 (N_2476,N_2437,N_2406);
or U2477 (N_2477,N_2450,N_2416);
and U2478 (N_2478,N_2402,N_2455);
nand U2479 (N_2479,N_2447,N_2427);
nor U2480 (N_2480,N_2454,N_2425);
or U2481 (N_2481,N_2459,N_2418);
nor U2482 (N_2482,N_2405,N_2413);
and U2483 (N_2483,N_2417,N_2444);
nor U2484 (N_2484,N_2438,N_2441);
or U2485 (N_2485,N_2448,N_2429);
and U2486 (N_2486,N_2415,N_2451);
nor U2487 (N_2487,N_2420,N_2414);
and U2488 (N_2488,N_2424,N_2411);
and U2489 (N_2489,N_2435,N_2409);
or U2490 (N_2490,N_2408,N_2431);
and U2491 (N_2491,N_2403,N_2418);
nand U2492 (N_2492,N_2424,N_2417);
and U2493 (N_2493,N_2438,N_2402);
nor U2494 (N_2494,N_2443,N_2416);
xor U2495 (N_2495,N_2454,N_2445);
nor U2496 (N_2496,N_2428,N_2443);
nor U2497 (N_2497,N_2454,N_2442);
and U2498 (N_2498,N_2411,N_2410);
nor U2499 (N_2499,N_2421,N_2414);
and U2500 (N_2500,N_2439,N_2452);
or U2501 (N_2501,N_2455,N_2452);
nor U2502 (N_2502,N_2412,N_2426);
or U2503 (N_2503,N_2448,N_2403);
nor U2504 (N_2504,N_2459,N_2442);
and U2505 (N_2505,N_2427,N_2426);
nor U2506 (N_2506,N_2415,N_2417);
xor U2507 (N_2507,N_2438,N_2430);
xnor U2508 (N_2508,N_2400,N_2450);
and U2509 (N_2509,N_2425,N_2408);
nand U2510 (N_2510,N_2417,N_2401);
nor U2511 (N_2511,N_2403,N_2429);
nor U2512 (N_2512,N_2401,N_2440);
nor U2513 (N_2513,N_2435,N_2428);
or U2514 (N_2514,N_2459,N_2438);
and U2515 (N_2515,N_2450,N_2455);
nor U2516 (N_2516,N_2419,N_2456);
or U2517 (N_2517,N_2440,N_2455);
nand U2518 (N_2518,N_2435,N_2434);
nor U2519 (N_2519,N_2414,N_2403);
and U2520 (N_2520,N_2465,N_2475);
xor U2521 (N_2521,N_2485,N_2461);
and U2522 (N_2522,N_2469,N_2463);
or U2523 (N_2523,N_2496,N_2491);
nand U2524 (N_2524,N_2498,N_2509);
nor U2525 (N_2525,N_2482,N_2500);
and U2526 (N_2526,N_2510,N_2488);
nor U2527 (N_2527,N_2478,N_2468);
and U2528 (N_2528,N_2519,N_2503);
or U2529 (N_2529,N_2472,N_2466);
and U2530 (N_2530,N_2517,N_2513);
or U2531 (N_2531,N_2518,N_2473);
and U2532 (N_2532,N_2487,N_2484);
or U2533 (N_2533,N_2481,N_2508);
and U2534 (N_2534,N_2486,N_2501);
or U2535 (N_2535,N_2477,N_2511);
nand U2536 (N_2536,N_2506,N_2515);
or U2537 (N_2537,N_2507,N_2476);
nand U2538 (N_2538,N_2505,N_2467);
or U2539 (N_2539,N_2460,N_2493);
nand U2540 (N_2540,N_2497,N_2495);
nand U2541 (N_2541,N_2499,N_2502);
and U2542 (N_2542,N_2516,N_2489);
and U2543 (N_2543,N_2492,N_2480);
or U2544 (N_2544,N_2471,N_2483);
and U2545 (N_2545,N_2490,N_2512);
and U2546 (N_2546,N_2464,N_2462);
and U2547 (N_2547,N_2504,N_2474);
and U2548 (N_2548,N_2494,N_2514);
and U2549 (N_2549,N_2470,N_2479);
nor U2550 (N_2550,N_2495,N_2488);
xnor U2551 (N_2551,N_2481,N_2461);
nor U2552 (N_2552,N_2488,N_2502);
xnor U2553 (N_2553,N_2474,N_2471);
xnor U2554 (N_2554,N_2485,N_2513);
nand U2555 (N_2555,N_2478,N_2508);
and U2556 (N_2556,N_2508,N_2491);
nand U2557 (N_2557,N_2482,N_2464);
or U2558 (N_2558,N_2506,N_2466);
and U2559 (N_2559,N_2463,N_2506);
nor U2560 (N_2560,N_2516,N_2517);
or U2561 (N_2561,N_2471,N_2460);
and U2562 (N_2562,N_2508,N_2471);
xnor U2563 (N_2563,N_2516,N_2461);
and U2564 (N_2564,N_2497,N_2468);
and U2565 (N_2565,N_2507,N_2498);
and U2566 (N_2566,N_2477,N_2479);
or U2567 (N_2567,N_2515,N_2484);
nor U2568 (N_2568,N_2493,N_2509);
nand U2569 (N_2569,N_2468,N_2466);
nor U2570 (N_2570,N_2461,N_2463);
nor U2571 (N_2571,N_2461,N_2466);
nor U2572 (N_2572,N_2509,N_2475);
nand U2573 (N_2573,N_2470,N_2501);
or U2574 (N_2574,N_2470,N_2504);
nor U2575 (N_2575,N_2517,N_2471);
nand U2576 (N_2576,N_2517,N_2476);
nor U2577 (N_2577,N_2477,N_2507);
xor U2578 (N_2578,N_2465,N_2505);
nand U2579 (N_2579,N_2468,N_2519);
nor U2580 (N_2580,N_2545,N_2522);
nand U2581 (N_2581,N_2556,N_2523);
or U2582 (N_2582,N_2546,N_2532);
or U2583 (N_2583,N_2552,N_2550);
and U2584 (N_2584,N_2539,N_2564);
nand U2585 (N_2585,N_2529,N_2566);
and U2586 (N_2586,N_2538,N_2561);
nand U2587 (N_2587,N_2531,N_2535);
and U2588 (N_2588,N_2577,N_2568);
or U2589 (N_2589,N_2534,N_2527);
nor U2590 (N_2590,N_2526,N_2524);
nand U2591 (N_2591,N_2576,N_2528);
nand U2592 (N_2592,N_2547,N_2548);
nand U2593 (N_2593,N_2559,N_2553);
nand U2594 (N_2594,N_2536,N_2544);
and U2595 (N_2595,N_2572,N_2562);
or U2596 (N_2596,N_2543,N_2571);
and U2597 (N_2597,N_2551,N_2530);
nand U2598 (N_2598,N_2541,N_2549);
nand U2599 (N_2599,N_2525,N_2560);
nor U2600 (N_2600,N_2542,N_2563);
and U2601 (N_2601,N_2555,N_2537);
nand U2602 (N_2602,N_2558,N_2521);
xor U2603 (N_2603,N_2554,N_2570);
or U2604 (N_2604,N_2569,N_2520);
and U2605 (N_2605,N_2579,N_2565);
or U2606 (N_2606,N_2574,N_2540);
nor U2607 (N_2607,N_2578,N_2575);
nand U2608 (N_2608,N_2573,N_2533);
and U2609 (N_2609,N_2567,N_2557);
nand U2610 (N_2610,N_2557,N_2563);
or U2611 (N_2611,N_2559,N_2530);
or U2612 (N_2612,N_2554,N_2540);
nor U2613 (N_2613,N_2541,N_2552);
or U2614 (N_2614,N_2533,N_2537);
and U2615 (N_2615,N_2542,N_2535);
and U2616 (N_2616,N_2540,N_2542);
nor U2617 (N_2617,N_2539,N_2561);
nand U2618 (N_2618,N_2542,N_2574);
nand U2619 (N_2619,N_2520,N_2561);
or U2620 (N_2620,N_2562,N_2529);
or U2621 (N_2621,N_2521,N_2535);
or U2622 (N_2622,N_2569,N_2527);
nand U2623 (N_2623,N_2550,N_2529);
or U2624 (N_2624,N_2561,N_2537);
or U2625 (N_2625,N_2538,N_2552);
nor U2626 (N_2626,N_2531,N_2562);
nand U2627 (N_2627,N_2576,N_2530);
or U2628 (N_2628,N_2533,N_2534);
or U2629 (N_2629,N_2526,N_2578);
nand U2630 (N_2630,N_2520,N_2574);
and U2631 (N_2631,N_2548,N_2536);
xor U2632 (N_2632,N_2533,N_2566);
or U2633 (N_2633,N_2520,N_2545);
and U2634 (N_2634,N_2555,N_2525);
or U2635 (N_2635,N_2572,N_2530);
or U2636 (N_2636,N_2540,N_2520);
and U2637 (N_2637,N_2540,N_2558);
and U2638 (N_2638,N_2531,N_2573);
xor U2639 (N_2639,N_2537,N_2557);
nand U2640 (N_2640,N_2639,N_2582);
xnor U2641 (N_2641,N_2617,N_2596);
nand U2642 (N_2642,N_2590,N_2602);
and U2643 (N_2643,N_2634,N_2625);
and U2644 (N_2644,N_2583,N_2588);
nor U2645 (N_2645,N_2587,N_2629);
and U2646 (N_2646,N_2624,N_2609);
xnor U2647 (N_2647,N_2599,N_2593);
or U2648 (N_2648,N_2605,N_2585);
xor U2649 (N_2649,N_2616,N_2586);
nand U2650 (N_2650,N_2628,N_2633);
nand U2651 (N_2651,N_2595,N_2613);
nand U2652 (N_2652,N_2607,N_2621);
nor U2653 (N_2653,N_2614,N_2615);
xnor U2654 (N_2654,N_2603,N_2580);
or U2655 (N_2655,N_2635,N_2598);
and U2656 (N_2656,N_2626,N_2611);
or U2657 (N_2657,N_2589,N_2592);
xnor U2658 (N_2658,N_2594,N_2601);
nor U2659 (N_2659,N_2630,N_2622);
nor U2660 (N_2660,N_2600,N_2591);
and U2661 (N_2661,N_2608,N_2636);
or U2662 (N_2662,N_2581,N_2627);
nor U2663 (N_2663,N_2637,N_2604);
nor U2664 (N_2664,N_2638,N_2631);
xnor U2665 (N_2665,N_2618,N_2619);
or U2666 (N_2666,N_2606,N_2612);
xnor U2667 (N_2667,N_2597,N_2623);
nor U2668 (N_2668,N_2584,N_2610);
or U2669 (N_2669,N_2620,N_2632);
nand U2670 (N_2670,N_2604,N_2598);
and U2671 (N_2671,N_2629,N_2596);
nand U2672 (N_2672,N_2592,N_2603);
nand U2673 (N_2673,N_2585,N_2595);
nor U2674 (N_2674,N_2619,N_2625);
xnor U2675 (N_2675,N_2616,N_2608);
or U2676 (N_2676,N_2580,N_2621);
xnor U2677 (N_2677,N_2604,N_2587);
nand U2678 (N_2678,N_2627,N_2621);
and U2679 (N_2679,N_2612,N_2629);
nor U2680 (N_2680,N_2596,N_2580);
and U2681 (N_2681,N_2595,N_2614);
nand U2682 (N_2682,N_2582,N_2618);
and U2683 (N_2683,N_2601,N_2631);
nand U2684 (N_2684,N_2638,N_2582);
nor U2685 (N_2685,N_2639,N_2600);
or U2686 (N_2686,N_2620,N_2596);
and U2687 (N_2687,N_2609,N_2581);
and U2688 (N_2688,N_2589,N_2582);
nor U2689 (N_2689,N_2613,N_2614);
nor U2690 (N_2690,N_2632,N_2602);
or U2691 (N_2691,N_2586,N_2625);
nand U2692 (N_2692,N_2638,N_2601);
nand U2693 (N_2693,N_2638,N_2610);
and U2694 (N_2694,N_2598,N_2586);
nor U2695 (N_2695,N_2622,N_2620);
nand U2696 (N_2696,N_2615,N_2639);
or U2697 (N_2697,N_2609,N_2636);
xor U2698 (N_2698,N_2629,N_2613);
nand U2699 (N_2699,N_2632,N_2583);
nand U2700 (N_2700,N_2654,N_2656);
nand U2701 (N_2701,N_2665,N_2667);
nand U2702 (N_2702,N_2686,N_2640);
and U2703 (N_2703,N_2683,N_2663);
or U2704 (N_2704,N_2669,N_2681);
and U2705 (N_2705,N_2648,N_2678);
and U2706 (N_2706,N_2680,N_2668);
nor U2707 (N_2707,N_2679,N_2658);
nand U2708 (N_2708,N_2650,N_2647);
and U2709 (N_2709,N_2660,N_2674);
xor U2710 (N_2710,N_2670,N_2699);
or U2711 (N_2711,N_2645,N_2689);
and U2712 (N_2712,N_2690,N_2661);
nor U2713 (N_2713,N_2646,N_2673);
or U2714 (N_2714,N_2653,N_2694);
or U2715 (N_2715,N_2693,N_2642);
and U2716 (N_2716,N_2698,N_2697);
nand U2717 (N_2717,N_2687,N_2685);
nand U2718 (N_2718,N_2664,N_2643);
or U2719 (N_2719,N_2696,N_2677);
nand U2720 (N_2720,N_2641,N_2666);
and U2721 (N_2721,N_2662,N_2695);
and U2722 (N_2722,N_2682,N_2688);
xnor U2723 (N_2723,N_2675,N_2644);
nand U2724 (N_2724,N_2655,N_2671);
and U2725 (N_2725,N_2652,N_2676);
xnor U2726 (N_2726,N_2649,N_2692);
xnor U2727 (N_2727,N_2659,N_2684);
nand U2728 (N_2728,N_2657,N_2691);
and U2729 (N_2729,N_2651,N_2672);
nor U2730 (N_2730,N_2669,N_2691);
and U2731 (N_2731,N_2699,N_2684);
and U2732 (N_2732,N_2654,N_2685);
nand U2733 (N_2733,N_2681,N_2691);
nor U2734 (N_2734,N_2663,N_2677);
nor U2735 (N_2735,N_2684,N_2648);
xnor U2736 (N_2736,N_2647,N_2665);
or U2737 (N_2737,N_2647,N_2684);
xor U2738 (N_2738,N_2674,N_2689);
nand U2739 (N_2739,N_2675,N_2660);
nor U2740 (N_2740,N_2683,N_2699);
or U2741 (N_2741,N_2653,N_2677);
and U2742 (N_2742,N_2642,N_2671);
nand U2743 (N_2743,N_2685,N_2681);
nor U2744 (N_2744,N_2690,N_2691);
nand U2745 (N_2745,N_2695,N_2670);
and U2746 (N_2746,N_2684,N_2642);
and U2747 (N_2747,N_2690,N_2672);
or U2748 (N_2748,N_2679,N_2652);
and U2749 (N_2749,N_2666,N_2691);
and U2750 (N_2750,N_2678,N_2680);
nand U2751 (N_2751,N_2659,N_2651);
or U2752 (N_2752,N_2661,N_2691);
xnor U2753 (N_2753,N_2685,N_2652);
nand U2754 (N_2754,N_2678,N_2646);
or U2755 (N_2755,N_2673,N_2692);
and U2756 (N_2756,N_2650,N_2679);
nor U2757 (N_2757,N_2680,N_2687);
nand U2758 (N_2758,N_2687,N_2672);
or U2759 (N_2759,N_2669,N_2673);
and U2760 (N_2760,N_2751,N_2745);
nor U2761 (N_2761,N_2707,N_2728);
and U2762 (N_2762,N_2755,N_2754);
and U2763 (N_2763,N_2739,N_2723);
and U2764 (N_2764,N_2703,N_2731);
or U2765 (N_2765,N_2725,N_2717);
and U2766 (N_2766,N_2756,N_2716);
and U2767 (N_2767,N_2737,N_2714);
nand U2768 (N_2768,N_2726,N_2722);
or U2769 (N_2769,N_2721,N_2710);
nand U2770 (N_2770,N_2711,N_2747);
or U2771 (N_2771,N_2704,N_2740);
nand U2772 (N_2772,N_2724,N_2733);
and U2773 (N_2773,N_2750,N_2759);
or U2774 (N_2774,N_2749,N_2757);
nand U2775 (N_2775,N_2753,N_2752);
nor U2776 (N_2776,N_2727,N_2709);
and U2777 (N_2777,N_2732,N_2743);
nand U2778 (N_2778,N_2734,N_2748);
or U2779 (N_2779,N_2713,N_2746);
and U2780 (N_2780,N_2708,N_2736);
or U2781 (N_2781,N_2742,N_2701);
nor U2782 (N_2782,N_2705,N_2735);
nand U2783 (N_2783,N_2702,N_2700);
nor U2784 (N_2784,N_2720,N_2741);
xnor U2785 (N_2785,N_2758,N_2744);
nor U2786 (N_2786,N_2738,N_2706);
nor U2787 (N_2787,N_2719,N_2712);
and U2788 (N_2788,N_2729,N_2730);
nand U2789 (N_2789,N_2718,N_2715);
nand U2790 (N_2790,N_2755,N_2721);
xnor U2791 (N_2791,N_2715,N_2702);
or U2792 (N_2792,N_2740,N_2715);
nand U2793 (N_2793,N_2716,N_2730);
nand U2794 (N_2794,N_2728,N_2716);
and U2795 (N_2795,N_2718,N_2735);
and U2796 (N_2796,N_2720,N_2753);
nand U2797 (N_2797,N_2741,N_2716);
xnor U2798 (N_2798,N_2719,N_2708);
nand U2799 (N_2799,N_2754,N_2748);
nor U2800 (N_2800,N_2713,N_2706);
xnor U2801 (N_2801,N_2710,N_2744);
nor U2802 (N_2802,N_2705,N_2750);
and U2803 (N_2803,N_2748,N_2731);
nand U2804 (N_2804,N_2716,N_2715);
or U2805 (N_2805,N_2734,N_2726);
xnor U2806 (N_2806,N_2700,N_2753);
nor U2807 (N_2807,N_2740,N_2712);
nand U2808 (N_2808,N_2742,N_2739);
nor U2809 (N_2809,N_2741,N_2723);
xnor U2810 (N_2810,N_2731,N_2744);
xor U2811 (N_2811,N_2755,N_2725);
or U2812 (N_2812,N_2746,N_2735);
nor U2813 (N_2813,N_2721,N_2716);
or U2814 (N_2814,N_2747,N_2735);
and U2815 (N_2815,N_2700,N_2732);
nand U2816 (N_2816,N_2702,N_2714);
nor U2817 (N_2817,N_2755,N_2746);
nand U2818 (N_2818,N_2757,N_2703);
nand U2819 (N_2819,N_2706,N_2730);
and U2820 (N_2820,N_2781,N_2809);
and U2821 (N_2821,N_2796,N_2798);
and U2822 (N_2822,N_2789,N_2801);
and U2823 (N_2823,N_2764,N_2816);
and U2824 (N_2824,N_2800,N_2776);
nor U2825 (N_2825,N_2779,N_2786);
xor U2826 (N_2826,N_2784,N_2807);
xor U2827 (N_2827,N_2788,N_2768);
nor U2828 (N_2828,N_2780,N_2783);
nor U2829 (N_2829,N_2775,N_2782);
and U2830 (N_2830,N_2762,N_2805);
and U2831 (N_2831,N_2760,N_2813);
xor U2832 (N_2832,N_2777,N_2791);
nor U2833 (N_2833,N_2804,N_2792);
nor U2834 (N_2834,N_2812,N_2770);
nor U2835 (N_2835,N_2810,N_2811);
and U2836 (N_2836,N_2772,N_2802);
xnor U2837 (N_2837,N_2771,N_2799);
and U2838 (N_2838,N_2818,N_2819);
and U2839 (N_2839,N_2774,N_2790);
or U2840 (N_2840,N_2778,N_2803);
and U2841 (N_2841,N_2806,N_2769);
nor U2842 (N_2842,N_2773,N_2766);
nor U2843 (N_2843,N_2795,N_2785);
xor U2844 (N_2844,N_2767,N_2765);
nor U2845 (N_2845,N_2793,N_2763);
nor U2846 (N_2846,N_2794,N_2817);
nor U2847 (N_2847,N_2787,N_2761);
nand U2848 (N_2848,N_2815,N_2814);
or U2849 (N_2849,N_2808,N_2797);
nand U2850 (N_2850,N_2807,N_2768);
nor U2851 (N_2851,N_2807,N_2808);
nor U2852 (N_2852,N_2760,N_2768);
and U2853 (N_2853,N_2786,N_2808);
and U2854 (N_2854,N_2772,N_2797);
or U2855 (N_2855,N_2808,N_2778);
nand U2856 (N_2856,N_2810,N_2765);
nand U2857 (N_2857,N_2764,N_2774);
nor U2858 (N_2858,N_2765,N_2775);
nor U2859 (N_2859,N_2783,N_2811);
or U2860 (N_2860,N_2807,N_2797);
xor U2861 (N_2861,N_2809,N_2819);
nor U2862 (N_2862,N_2762,N_2804);
and U2863 (N_2863,N_2817,N_2762);
xnor U2864 (N_2864,N_2800,N_2761);
nand U2865 (N_2865,N_2803,N_2776);
nor U2866 (N_2866,N_2792,N_2775);
xnor U2867 (N_2867,N_2817,N_2768);
nor U2868 (N_2868,N_2785,N_2810);
or U2869 (N_2869,N_2806,N_2780);
or U2870 (N_2870,N_2798,N_2799);
and U2871 (N_2871,N_2774,N_2761);
nor U2872 (N_2872,N_2776,N_2811);
nand U2873 (N_2873,N_2798,N_2810);
nor U2874 (N_2874,N_2804,N_2810);
xnor U2875 (N_2875,N_2777,N_2815);
or U2876 (N_2876,N_2790,N_2798);
xnor U2877 (N_2877,N_2815,N_2772);
xnor U2878 (N_2878,N_2818,N_2784);
nand U2879 (N_2879,N_2765,N_2816);
or U2880 (N_2880,N_2879,N_2822);
or U2881 (N_2881,N_2863,N_2851);
and U2882 (N_2882,N_2837,N_2856);
nor U2883 (N_2883,N_2875,N_2830);
nand U2884 (N_2884,N_2878,N_2840);
nand U2885 (N_2885,N_2829,N_2864);
and U2886 (N_2886,N_2834,N_2877);
xnor U2887 (N_2887,N_2841,N_2876);
nor U2888 (N_2888,N_2839,N_2849);
or U2889 (N_2889,N_2855,N_2860);
and U2890 (N_2890,N_2871,N_2873);
or U2891 (N_2891,N_2842,N_2825);
and U2892 (N_2892,N_2854,N_2831);
or U2893 (N_2893,N_2852,N_2838);
or U2894 (N_2894,N_2858,N_2823);
or U2895 (N_2895,N_2828,N_2862);
nor U2896 (N_2896,N_2850,N_2869);
or U2897 (N_2897,N_2843,N_2827);
nor U2898 (N_2898,N_2824,N_2874);
xor U2899 (N_2899,N_2859,N_2833);
and U2900 (N_2900,N_2821,N_2835);
nor U2901 (N_2901,N_2857,N_2865);
and U2902 (N_2902,N_2853,N_2847);
and U2903 (N_2903,N_2845,N_2846);
nand U2904 (N_2904,N_2848,N_2844);
or U2905 (N_2905,N_2820,N_2867);
nor U2906 (N_2906,N_2836,N_2832);
nor U2907 (N_2907,N_2868,N_2861);
nor U2908 (N_2908,N_2872,N_2866);
and U2909 (N_2909,N_2826,N_2870);
nand U2910 (N_2910,N_2833,N_2851);
nand U2911 (N_2911,N_2825,N_2820);
xor U2912 (N_2912,N_2868,N_2826);
nor U2913 (N_2913,N_2826,N_2871);
nand U2914 (N_2914,N_2829,N_2840);
nor U2915 (N_2915,N_2873,N_2872);
or U2916 (N_2916,N_2877,N_2858);
nand U2917 (N_2917,N_2848,N_2875);
nand U2918 (N_2918,N_2870,N_2835);
and U2919 (N_2919,N_2855,N_2868);
or U2920 (N_2920,N_2872,N_2827);
nor U2921 (N_2921,N_2866,N_2852);
nand U2922 (N_2922,N_2873,N_2827);
nor U2923 (N_2923,N_2863,N_2836);
nor U2924 (N_2924,N_2870,N_2850);
or U2925 (N_2925,N_2858,N_2847);
nor U2926 (N_2926,N_2826,N_2851);
nor U2927 (N_2927,N_2831,N_2836);
nor U2928 (N_2928,N_2867,N_2838);
and U2929 (N_2929,N_2839,N_2858);
nor U2930 (N_2930,N_2842,N_2848);
and U2931 (N_2931,N_2868,N_2866);
and U2932 (N_2932,N_2871,N_2840);
nor U2933 (N_2933,N_2821,N_2865);
or U2934 (N_2934,N_2869,N_2835);
nand U2935 (N_2935,N_2838,N_2874);
and U2936 (N_2936,N_2867,N_2841);
or U2937 (N_2937,N_2859,N_2860);
nand U2938 (N_2938,N_2870,N_2827);
xor U2939 (N_2939,N_2835,N_2860);
nand U2940 (N_2940,N_2895,N_2900);
and U2941 (N_2941,N_2938,N_2914);
or U2942 (N_2942,N_2885,N_2925);
nand U2943 (N_2943,N_2933,N_2929);
nand U2944 (N_2944,N_2928,N_2897);
or U2945 (N_2945,N_2922,N_2891);
and U2946 (N_2946,N_2884,N_2883);
and U2947 (N_2947,N_2912,N_2936);
nor U2948 (N_2948,N_2917,N_2909);
nand U2949 (N_2949,N_2923,N_2939);
xor U2950 (N_2950,N_2899,N_2898);
xnor U2951 (N_2951,N_2913,N_2888);
or U2952 (N_2952,N_2918,N_2927);
or U2953 (N_2953,N_2880,N_2881);
and U2954 (N_2954,N_2889,N_2905);
nand U2955 (N_2955,N_2937,N_2934);
nand U2956 (N_2956,N_2903,N_2894);
or U2957 (N_2957,N_2908,N_2910);
nand U2958 (N_2958,N_2907,N_2882);
nor U2959 (N_2959,N_2911,N_2930);
nor U2960 (N_2960,N_2887,N_2919);
nor U2961 (N_2961,N_2906,N_2901);
or U2962 (N_2962,N_2931,N_2916);
and U2963 (N_2963,N_2924,N_2890);
or U2964 (N_2964,N_2902,N_2904);
nand U2965 (N_2965,N_2921,N_2892);
xor U2966 (N_2966,N_2896,N_2893);
nor U2967 (N_2967,N_2915,N_2932);
and U2968 (N_2968,N_2926,N_2920);
xnor U2969 (N_2969,N_2935,N_2886);
nand U2970 (N_2970,N_2905,N_2914);
nor U2971 (N_2971,N_2890,N_2892);
or U2972 (N_2972,N_2910,N_2926);
nor U2973 (N_2973,N_2890,N_2901);
or U2974 (N_2974,N_2924,N_2897);
nor U2975 (N_2975,N_2899,N_2886);
and U2976 (N_2976,N_2899,N_2934);
or U2977 (N_2977,N_2900,N_2904);
and U2978 (N_2978,N_2889,N_2907);
nand U2979 (N_2979,N_2906,N_2909);
or U2980 (N_2980,N_2934,N_2885);
nor U2981 (N_2981,N_2910,N_2920);
nor U2982 (N_2982,N_2887,N_2915);
nor U2983 (N_2983,N_2892,N_2919);
xnor U2984 (N_2984,N_2880,N_2899);
and U2985 (N_2985,N_2900,N_2880);
nor U2986 (N_2986,N_2933,N_2907);
nand U2987 (N_2987,N_2908,N_2893);
or U2988 (N_2988,N_2919,N_2912);
xnor U2989 (N_2989,N_2931,N_2935);
nand U2990 (N_2990,N_2885,N_2910);
and U2991 (N_2991,N_2928,N_2938);
and U2992 (N_2992,N_2920,N_2922);
xnor U2993 (N_2993,N_2922,N_2897);
nor U2994 (N_2994,N_2910,N_2891);
nand U2995 (N_2995,N_2890,N_2894);
or U2996 (N_2996,N_2918,N_2935);
nand U2997 (N_2997,N_2880,N_2896);
xnor U2998 (N_2998,N_2933,N_2888);
or U2999 (N_2999,N_2900,N_2886);
or UO_0 (O_0,N_2999,N_2977);
or UO_1 (O_1,N_2996,N_2949);
or UO_2 (O_2,N_2964,N_2974);
nand UO_3 (O_3,N_2969,N_2976);
xor UO_4 (O_4,N_2962,N_2954);
nor UO_5 (O_5,N_2981,N_2988);
xnor UO_6 (O_6,N_2987,N_2968);
xnor UO_7 (O_7,N_2941,N_2948);
or UO_8 (O_8,N_2958,N_2944);
nor UO_9 (O_9,N_2963,N_2955);
xor UO_10 (O_10,N_2943,N_2959);
and UO_11 (O_11,N_2947,N_2985);
and UO_12 (O_12,N_2952,N_2993);
xor UO_13 (O_13,N_2978,N_2990);
or UO_14 (O_14,N_2995,N_2965);
and UO_15 (O_15,N_2980,N_2992);
and UO_16 (O_16,N_2982,N_2950);
nand UO_17 (O_17,N_2970,N_2942);
nand UO_18 (O_18,N_2972,N_2975);
nand UO_19 (O_19,N_2971,N_2953);
or UO_20 (O_20,N_2967,N_2994);
nor UO_21 (O_21,N_2957,N_2984);
nor UO_22 (O_22,N_2979,N_2966);
nor UO_23 (O_23,N_2983,N_2960);
xnor UO_24 (O_24,N_2998,N_2951);
nand UO_25 (O_25,N_2940,N_2946);
or UO_26 (O_26,N_2986,N_2961);
xor UO_27 (O_27,N_2997,N_2973);
nor UO_28 (O_28,N_2956,N_2989);
nor UO_29 (O_29,N_2991,N_2945);
nand UO_30 (O_30,N_2945,N_2962);
and UO_31 (O_31,N_2947,N_2961);
nand UO_32 (O_32,N_2947,N_2963);
and UO_33 (O_33,N_2988,N_2973);
nand UO_34 (O_34,N_2970,N_2948);
nor UO_35 (O_35,N_2998,N_2972);
nand UO_36 (O_36,N_2948,N_2960);
nand UO_37 (O_37,N_2950,N_2981);
nor UO_38 (O_38,N_2943,N_2948);
xnor UO_39 (O_39,N_2951,N_2944);
and UO_40 (O_40,N_2986,N_2996);
or UO_41 (O_41,N_2961,N_2960);
or UO_42 (O_42,N_2949,N_2963);
and UO_43 (O_43,N_2962,N_2964);
nand UO_44 (O_44,N_2941,N_2964);
or UO_45 (O_45,N_2999,N_2979);
nand UO_46 (O_46,N_2998,N_2975);
and UO_47 (O_47,N_2941,N_2940);
xnor UO_48 (O_48,N_2945,N_2967);
and UO_49 (O_49,N_2981,N_2962);
xor UO_50 (O_50,N_2975,N_2947);
and UO_51 (O_51,N_2949,N_2965);
or UO_52 (O_52,N_2965,N_2976);
nor UO_53 (O_53,N_2980,N_2950);
nor UO_54 (O_54,N_2955,N_2999);
and UO_55 (O_55,N_2949,N_2966);
nand UO_56 (O_56,N_2993,N_2996);
nor UO_57 (O_57,N_2948,N_2952);
xor UO_58 (O_58,N_2958,N_2965);
and UO_59 (O_59,N_2958,N_2961);
or UO_60 (O_60,N_2966,N_2984);
xor UO_61 (O_61,N_2960,N_2975);
nor UO_62 (O_62,N_2940,N_2955);
nor UO_63 (O_63,N_2972,N_2961);
or UO_64 (O_64,N_2976,N_2986);
or UO_65 (O_65,N_2942,N_2972);
nand UO_66 (O_66,N_2963,N_2975);
nor UO_67 (O_67,N_2970,N_2958);
and UO_68 (O_68,N_2977,N_2978);
nor UO_69 (O_69,N_2952,N_2979);
or UO_70 (O_70,N_2986,N_2967);
nand UO_71 (O_71,N_2988,N_2979);
nor UO_72 (O_72,N_2945,N_2958);
nand UO_73 (O_73,N_2971,N_2988);
nor UO_74 (O_74,N_2991,N_2972);
or UO_75 (O_75,N_2959,N_2985);
and UO_76 (O_76,N_2982,N_2972);
nand UO_77 (O_77,N_2989,N_2966);
nor UO_78 (O_78,N_2974,N_2971);
nor UO_79 (O_79,N_2951,N_2943);
or UO_80 (O_80,N_2996,N_2984);
or UO_81 (O_81,N_2969,N_2981);
or UO_82 (O_82,N_2995,N_2968);
or UO_83 (O_83,N_2954,N_2992);
nand UO_84 (O_84,N_2973,N_2941);
and UO_85 (O_85,N_2946,N_2973);
or UO_86 (O_86,N_2955,N_2969);
and UO_87 (O_87,N_2958,N_2991);
nor UO_88 (O_88,N_2981,N_2967);
nand UO_89 (O_89,N_2960,N_2969);
nor UO_90 (O_90,N_2951,N_2997);
nor UO_91 (O_91,N_2947,N_2993);
or UO_92 (O_92,N_2958,N_2986);
or UO_93 (O_93,N_2972,N_2979);
and UO_94 (O_94,N_2998,N_2964);
nor UO_95 (O_95,N_2998,N_2982);
nand UO_96 (O_96,N_2948,N_2995);
nand UO_97 (O_97,N_2967,N_2983);
and UO_98 (O_98,N_2985,N_2975);
nor UO_99 (O_99,N_2942,N_2989);
xor UO_100 (O_100,N_2945,N_2957);
nand UO_101 (O_101,N_2948,N_2958);
nand UO_102 (O_102,N_2966,N_2955);
or UO_103 (O_103,N_2979,N_2965);
nor UO_104 (O_104,N_2984,N_2946);
or UO_105 (O_105,N_2967,N_2950);
or UO_106 (O_106,N_2951,N_2973);
nor UO_107 (O_107,N_2954,N_2942);
and UO_108 (O_108,N_2948,N_2981);
nor UO_109 (O_109,N_2945,N_2966);
or UO_110 (O_110,N_2966,N_2983);
xor UO_111 (O_111,N_2993,N_2960);
and UO_112 (O_112,N_2950,N_2962);
nand UO_113 (O_113,N_2974,N_2988);
and UO_114 (O_114,N_2956,N_2983);
and UO_115 (O_115,N_2951,N_2969);
nor UO_116 (O_116,N_2981,N_2971);
nor UO_117 (O_117,N_2951,N_2948);
and UO_118 (O_118,N_2974,N_2956);
or UO_119 (O_119,N_2969,N_2945);
nor UO_120 (O_120,N_2978,N_2984);
nor UO_121 (O_121,N_2988,N_2951);
and UO_122 (O_122,N_2959,N_2995);
nand UO_123 (O_123,N_2982,N_2999);
nand UO_124 (O_124,N_2989,N_2951);
or UO_125 (O_125,N_2966,N_2998);
xnor UO_126 (O_126,N_2972,N_2999);
and UO_127 (O_127,N_2992,N_2997);
nand UO_128 (O_128,N_2981,N_2947);
or UO_129 (O_129,N_2968,N_2969);
nand UO_130 (O_130,N_2967,N_2989);
and UO_131 (O_131,N_2990,N_2971);
nand UO_132 (O_132,N_2984,N_2991);
or UO_133 (O_133,N_2974,N_2976);
and UO_134 (O_134,N_2968,N_2945);
nand UO_135 (O_135,N_2976,N_2970);
and UO_136 (O_136,N_2994,N_2991);
and UO_137 (O_137,N_2967,N_2955);
or UO_138 (O_138,N_2942,N_2955);
nor UO_139 (O_139,N_2977,N_2998);
nor UO_140 (O_140,N_2948,N_2963);
or UO_141 (O_141,N_2976,N_2943);
nor UO_142 (O_142,N_2967,N_2966);
nor UO_143 (O_143,N_2961,N_2978);
nor UO_144 (O_144,N_2942,N_2968);
nor UO_145 (O_145,N_2945,N_2979);
and UO_146 (O_146,N_2977,N_2958);
nand UO_147 (O_147,N_2941,N_2974);
or UO_148 (O_148,N_2987,N_2941);
and UO_149 (O_149,N_2956,N_2944);
nand UO_150 (O_150,N_2964,N_2983);
and UO_151 (O_151,N_2973,N_2987);
and UO_152 (O_152,N_2999,N_2987);
nand UO_153 (O_153,N_2973,N_2948);
nand UO_154 (O_154,N_2946,N_2983);
and UO_155 (O_155,N_2982,N_2976);
or UO_156 (O_156,N_2988,N_2945);
nand UO_157 (O_157,N_2979,N_2956);
nand UO_158 (O_158,N_2982,N_2995);
or UO_159 (O_159,N_2960,N_2994);
nand UO_160 (O_160,N_2964,N_2992);
and UO_161 (O_161,N_2959,N_2979);
or UO_162 (O_162,N_2999,N_2953);
or UO_163 (O_163,N_2956,N_2993);
or UO_164 (O_164,N_2979,N_2967);
or UO_165 (O_165,N_2953,N_2984);
nand UO_166 (O_166,N_2963,N_2952);
and UO_167 (O_167,N_2965,N_2989);
or UO_168 (O_168,N_2944,N_2969);
xor UO_169 (O_169,N_2940,N_2995);
nor UO_170 (O_170,N_2954,N_2981);
nand UO_171 (O_171,N_2962,N_2963);
and UO_172 (O_172,N_2942,N_2978);
nand UO_173 (O_173,N_2989,N_2997);
nor UO_174 (O_174,N_2988,N_2996);
and UO_175 (O_175,N_2994,N_2993);
and UO_176 (O_176,N_2998,N_2990);
nand UO_177 (O_177,N_2988,N_2963);
and UO_178 (O_178,N_2948,N_2992);
and UO_179 (O_179,N_2979,N_2983);
nor UO_180 (O_180,N_2949,N_2988);
nor UO_181 (O_181,N_2962,N_2944);
or UO_182 (O_182,N_2996,N_2969);
nand UO_183 (O_183,N_2982,N_2986);
nor UO_184 (O_184,N_2995,N_2997);
or UO_185 (O_185,N_2997,N_2950);
or UO_186 (O_186,N_2956,N_2973);
nor UO_187 (O_187,N_2941,N_2945);
nand UO_188 (O_188,N_2941,N_2969);
nand UO_189 (O_189,N_2994,N_2986);
nor UO_190 (O_190,N_2983,N_2952);
nor UO_191 (O_191,N_2944,N_2961);
nor UO_192 (O_192,N_2959,N_2994);
nand UO_193 (O_193,N_2982,N_2961);
nand UO_194 (O_194,N_2956,N_2999);
or UO_195 (O_195,N_2941,N_2947);
nor UO_196 (O_196,N_2966,N_2977);
or UO_197 (O_197,N_2940,N_2952);
nor UO_198 (O_198,N_2973,N_2957);
nand UO_199 (O_199,N_2993,N_2971);
and UO_200 (O_200,N_2999,N_2992);
xnor UO_201 (O_201,N_2978,N_2991);
nand UO_202 (O_202,N_2970,N_2998);
xor UO_203 (O_203,N_2979,N_2953);
or UO_204 (O_204,N_2994,N_2961);
or UO_205 (O_205,N_2944,N_2943);
nand UO_206 (O_206,N_2966,N_2954);
nand UO_207 (O_207,N_2952,N_2988);
and UO_208 (O_208,N_2957,N_2996);
xor UO_209 (O_209,N_2958,N_2995);
nor UO_210 (O_210,N_2956,N_2970);
or UO_211 (O_211,N_2965,N_2961);
or UO_212 (O_212,N_2999,N_2998);
and UO_213 (O_213,N_2956,N_2955);
nor UO_214 (O_214,N_2964,N_2996);
and UO_215 (O_215,N_2968,N_2979);
nand UO_216 (O_216,N_2964,N_2955);
nor UO_217 (O_217,N_2973,N_2953);
or UO_218 (O_218,N_2975,N_2999);
xor UO_219 (O_219,N_2976,N_2989);
or UO_220 (O_220,N_2947,N_2979);
and UO_221 (O_221,N_2954,N_2952);
nand UO_222 (O_222,N_2995,N_2950);
nor UO_223 (O_223,N_2978,N_2995);
or UO_224 (O_224,N_2961,N_2955);
xnor UO_225 (O_225,N_2964,N_2987);
nand UO_226 (O_226,N_2985,N_2961);
xor UO_227 (O_227,N_2968,N_2996);
and UO_228 (O_228,N_2969,N_2943);
and UO_229 (O_229,N_2952,N_2995);
and UO_230 (O_230,N_2983,N_2969);
nor UO_231 (O_231,N_2996,N_2995);
nor UO_232 (O_232,N_2953,N_2957);
and UO_233 (O_233,N_2980,N_2976);
and UO_234 (O_234,N_2992,N_2968);
and UO_235 (O_235,N_2987,N_2986);
nand UO_236 (O_236,N_2961,N_2989);
nor UO_237 (O_237,N_2948,N_2987);
or UO_238 (O_238,N_2964,N_2954);
nor UO_239 (O_239,N_2957,N_2961);
and UO_240 (O_240,N_2944,N_2949);
or UO_241 (O_241,N_2956,N_2957);
nor UO_242 (O_242,N_2946,N_2965);
and UO_243 (O_243,N_2940,N_2961);
and UO_244 (O_244,N_2950,N_2949);
nor UO_245 (O_245,N_2990,N_2959);
and UO_246 (O_246,N_2950,N_2969);
or UO_247 (O_247,N_2963,N_2957);
nand UO_248 (O_248,N_2942,N_2986);
nor UO_249 (O_249,N_2990,N_2957);
xnor UO_250 (O_250,N_2970,N_2992);
nand UO_251 (O_251,N_2952,N_2996);
or UO_252 (O_252,N_2993,N_2943);
xor UO_253 (O_253,N_2987,N_2985);
xor UO_254 (O_254,N_2970,N_2964);
or UO_255 (O_255,N_2980,N_2952);
xor UO_256 (O_256,N_2948,N_2945);
nor UO_257 (O_257,N_2959,N_2946);
nor UO_258 (O_258,N_2944,N_2994);
nor UO_259 (O_259,N_2947,N_2946);
or UO_260 (O_260,N_2974,N_2945);
nand UO_261 (O_261,N_2970,N_2949);
nand UO_262 (O_262,N_2946,N_2970);
xor UO_263 (O_263,N_2954,N_2957);
and UO_264 (O_264,N_2992,N_2991);
or UO_265 (O_265,N_2995,N_2990);
or UO_266 (O_266,N_2970,N_2960);
and UO_267 (O_267,N_2952,N_2971);
or UO_268 (O_268,N_2973,N_2947);
nand UO_269 (O_269,N_2957,N_2980);
nand UO_270 (O_270,N_2945,N_2980);
and UO_271 (O_271,N_2974,N_2961);
nor UO_272 (O_272,N_2980,N_2965);
xor UO_273 (O_273,N_2982,N_2947);
or UO_274 (O_274,N_2972,N_2994);
and UO_275 (O_275,N_2947,N_2984);
nor UO_276 (O_276,N_2942,N_2960);
or UO_277 (O_277,N_2957,N_2950);
nor UO_278 (O_278,N_2981,N_2940);
xnor UO_279 (O_279,N_2960,N_2999);
and UO_280 (O_280,N_2940,N_2950);
and UO_281 (O_281,N_2955,N_2985);
xor UO_282 (O_282,N_2962,N_2956);
nor UO_283 (O_283,N_2978,N_2950);
and UO_284 (O_284,N_2940,N_2963);
nor UO_285 (O_285,N_2958,N_2989);
nor UO_286 (O_286,N_2980,N_2973);
and UO_287 (O_287,N_2993,N_2951);
nor UO_288 (O_288,N_2941,N_2965);
or UO_289 (O_289,N_2949,N_2997);
nor UO_290 (O_290,N_2991,N_2960);
nor UO_291 (O_291,N_2968,N_2997);
or UO_292 (O_292,N_2960,N_2955);
nor UO_293 (O_293,N_2985,N_2965);
or UO_294 (O_294,N_2942,N_2993);
or UO_295 (O_295,N_2999,N_2986);
xnor UO_296 (O_296,N_2986,N_2977);
nand UO_297 (O_297,N_2982,N_2996);
nor UO_298 (O_298,N_2944,N_2966);
xnor UO_299 (O_299,N_2948,N_2997);
nor UO_300 (O_300,N_2984,N_2948);
and UO_301 (O_301,N_2977,N_2971);
or UO_302 (O_302,N_2996,N_2948);
and UO_303 (O_303,N_2965,N_2970);
nand UO_304 (O_304,N_2980,N_2947);
nor UO_305 (O_305,N_2972,N_2997);
nand UO_306 (O_306,N_2954,N_2982);
nand UO_307 (O_307,N_2967,N_2944);
and UO_308 (O_308,N_2995,N_2943);
or UO_309 (O_309,N_2960,N_2982);
and UO_310 (O_310,N_2953,N_2960);
or UO_311 (O_311,N_2985,N_2973);
xor UO_312 (O_312,N_2954,N_2995);
nand UO_313 (O_313,N_2945,N_2982);
nand UO_314 (O_314,N_2991,N_2999);
or UO_315 (O_315,N_2947,N_2952);
or UO_316 (O_316,N_2987,N_2975);
nand UO_317 (O_317,N_2985,N_2997);
nand UO_318 (O_318,N_2978,N_2952);
nand UO_319 (O_319,N_2990,N_2963);
nand UO_320 (O_320,N_2968,N_2986);
or UO_321 (O_321,N_2955,N_2972);
and UO_322 (O_322,N_2992,N_2971);
nand UO_323 (O_323,N_2984,N_2987);
or UO_324 (O_324,N_2992,N_2972);
or UO_325 (O_325,N_2966,N_2995);
nand UO_326 (O_326,N_2954,N_2984);
nand UO_327 (O_327,N_2999,N_2988);
or UO_328 (O_328,N_2990,N_2980);
or UO_329 (O_329,N_2957,N_2997);
xnor UO_330 (O_330,N_2964,N_2978);
nand UO_331 (O_331,N_2945,N_2949);
nand UO_332 (O_332,N_2998,N_2994);
nor UO_333 (O_333,N_2951,N_2952);
or UO_334 (O_334,N_2950,N_2999);
nor UO_335 (O_335,N_2941,N_2992);
nand UO_336 (O_336,N_2945,N_2990);
or UO_337 (O_337,N_2946,N_2997);
xor UO_338 (O_338,N_2994,N_2943);
or UO_339 (O_339,N_2976,N_2997);
and UO_340 (O_340,N_2989,N_2996);
nand UO_341 (O_341,N_2941,N_2953);
and UO_342 (O_342,N_2953,N_2980);
and UO_343 (O_343,N_2967,N_2982);
nor UO_344 (O_344,N_2966,N_2965);
nand UO_345 (O_345,N_2991,N_2993);
nor UO_346 (O_346,N_2966,N_2974);
nor UO_347 (O_347,N_2940,N_2988);
nand UO_348 (O_348,N_2957,N_2959);
or UO_349 (O_349,N_2993,N_2966);
or UO_350 (O_350,N_2970,N_2972);
nor UO_351 (O_351,N_2976,N_2945);
and UO_352 (O_352,N_2965,N_2957);
nor UO_353 (O_353,N_2968,N_2963);
or UO_354 (O_354,N_2970,N_2993);
nor UO_355 (O_355,N_2945,N_2999);
and UO_356 (O_356,N_2971,N_2957);
xnor UO_357 (O_357,N_2998,N_2983);
nand UO_358 (O_358,N_2941,N_2967);
or UO_359 (O_359,N_2960,N_2977);
nand UO_360 (O_360,N_2971,N_2950);
or UO_361 (O_361,N_2993,N_2940);
or UO_362 (O_362,N_2945,N_2997);
and UO_363 (O_363,N_2968,N_2966);
xor UO_364 (O_364,N_2995,N_2991);
or UO_365 (O_365,N_2955,N_2949);
and UO_366 (O_366,N_2958,N_2984);
and UO_367 (O_367,N_2963,N_2976);
nand UO_368 (O_368,N_2965,N_2996);
or UO_369 (O_369,N_2969,N_2973);
and UO_370 (O_370,N_2941,N_2960);
nand UO_371 (O_371,N_2961,N_2951);
or UO_372 (O_372,N_2950,N_2996);
nand UO_373 (O_373,N_2996,N_2980);
nor UO_374 (O_374,N_2974,N_2963);
nand UO_375 (O_375,N_2958,N_2952);
nand UO_376 (O_376,N_2950,N_2989);
or UO_377 (O_377,N_2973,N_2994);
or UO_378 (O_378,N_2950,N_2952);
nor UO_379 (O_379,N_2960,N_2966);
xnor UO_380 (O_380,N_2990,N_2940);
nand UO_381 (O_381,N_2986,N_2971);
xor UO_382 (O_382,N_2985,N_2988);
and UO_383 (O_383,N_2947,N_2953);
and UO_384 (O_384,N_2977,N_2982);
and UO_385 (O_385,N_2950,N_2951);
and UO_386 (O_386,N_2985,N_2949);
or UO_387 (O_387,N_2985,N_2982);
nor UO_388 (O_388,N_2971,N_2994);
nor UO_389 (O_389,N_2973,N_2996);
nor UO_390 (O_390,N_2953,N_2978);
nor UO_391 (O_391,N_2967,N_2959);
xnor UO_392 (O_392,N_2961,N_2993);
nand UO_393 (O_393,N_2973,N_2978);
nand UO_394 (O_394,N_2977,N_2946);
or UO_395 (O_395,N_2995,N_2980);
nor UO_396 (O_396,N_2946,N_2954);
xor UO_397 (O_397,N_2988,N_2965);
or UO_398 (O_398,N_2940,N_2965);
nand UO_399 (O_399,N_2999,N_2993);
xnor UO_400 (O_400,N_2980,N_2998);
nor UO_401 (O_401,N_2974,N_2959);
and UO_402 (O_402,N_2994,N_2963);
and UO_403 (O_403,N_2950,N_2988);
nor UO_404 (O_404,N_2983,N_2972);
nor UO_405 (O_405,N_2979,N_2986);
nor UO_406 (O_406,N_2961,N_2996);
xor UO_407 (O_407,N_2944,N_2971);
xnor UO_408 (O_408,N_2945,N_2952);
and UO_409 (O_409,N_2966,N_2943);
nand UO_410 (O_410,N_2987,N_2979);
and UO_411 (O_411,N_2949,N_2973);
nor UO_412 (O_412,N_2973,N_2989);
nor UO_413 (O_413,N_2997,N_2943);
and UO_414 (O_414,N_2991,N_2961);
xnor UO_415 (O_415,N_2949,N_2983);
or UO_416 (O_416,N_2953,N_2988);
nand UO_417 (O_417,N_2999,N_2946);
and UO_418 (O_418,N_2981,N_2977);
and UO_419 (O_419,N_2961,N_2963);
or UO_420 (O_420,N_2999,N_2980);
and UO_421 (O_421,N_2983,N_2945);
nor UO_422 (O_422,N_2998,N_2956);
and UO_423 (O_423,N_2985,N_2993);
or UO_424 (O_424,N_2952,N_2977);
nand UO_425 (O_425,N_2962,N_2977);
and UO_426 (O_426,N_2997,N_2967);
or UO_427 (O_427,N_2947,N_2995);
nor UO_428 (O_428,N_2961,N_2976);
xnor UO_429 (O_429,N_2944,N_2947);
nor UO_430 (O_430,N_2985,N_2954);
xnor UO_431 (O_431,N_2944,N_2960);
nand UO_432 (O_432,N_2996,N_2940);
nor UO_433 (O_433,N_2980,N_2956);
and UO_434 (O_434,N_2984,N_2974);
nand UO_435 (O_435,N_2958,N_2993);
nor UO_436 (O_436,N_2983,N_2963);
or UO_437 (O_437,N_2987,N_2949);
and UO_438 (O_438,N_2948,N_2957);
nand UO_439 (O_439,N_2960,N_2986);
nor UO_440 (O_440,N_2984,N_2972);
nand UO_441 (O_441,N_2990,N_2982);
nand UO_442 (O_442,N_2961,N_2998);
and UO_443 (O_443,N_2996,N_2963);
or UO_444 (O_444,N_2970,N_2984);
xor UO_445 (O_445,N_2955,N_2975);
xnor UO_446 (O_446,N_2983,N_2947);
or UO_447 (O_447,N_2958,N_2971);
or UO_448 (O_448,N_2956,N_2988);
and UO_449 (O_449,N_2955,N_2944);
and UO_450 (O_450,N_2971,N_2983);
and UO_451 (O_451,N_2995,N_2949);
nor UO_452 (O_452,N_2984,N_2965);
nor UO_453 (O_453,N_2984,N_2993);
nand UO_454 (O_454,N_2952,N_2994);
nand UO_455 (O_455,N_2962,N_2996);
nor UO_456 (O_456,N_2948,N_2968);
nand UO_457 (O_457,N_2957,N_2993);
or UO_458 (O_458,N_2973,N_2958);
nor UO_459 (O_459,N_2996,N_2966);
xor UO_460 (O_460,N_2999,N_2962);
nand UO_461 (O_461,N_2973,N_2976);
nand UO_462 (O_462,N_2984,N_2997);
xor UO_463 (O_463,N_2988,N_2992);
or UO_464 (O_464,N_2940,N_2956);
nand UO_465 (O_465,N_2949,N_2971);
nor UO_466 (O_466,N_2974,N_2986);
nand UO_467 (O_467,N_2970,N_2995);
xnor UO_468 (O_468,N_2963,N_2985);
or UO_469 (O_469,N_2943,N_2974);
xor UO_470 (O_470,N_2946,N_2972);
nor UO_471 (O_471,N_2969,N_2966);
and UO_472 (O_472,N_2972,N_2965);
nand UO_473 (O_473,N_2974,N_2954);
and UO_474 (O_474,N_2971,N_2959);
nor UO_475 (O_475,N_2993,N_2955);
nor UO_476 (O_476,N_2949,N_2946);
nor UO_477 (O_477,N_2965,N_2969);
nand UO_478 (O_478,N_2981,N_2986);
or UO_479 (O_479,N_2998,N_2985);
nor UO_480 (O_480,N_2983,N_2973);
and UO_481 (O_481,N_2977,N_2993);
nor UO_482 (O_482,N_2962,N_2973);
or UO_483 (O_483,N_2970,N_2990);
and UO_484 (O_484,N_2948,N_2982);
nand UO_485 (O_485,N_2987,N_2989);
nand UO_486 (O_486,N_2946,N_2981);
nor UO_487 (O_487,N_2943,N_2991);
and UO_488 (O_488,N_2945,N_2963);
nor UO_489 (O_489,N_2983,N_2984);
and UO_490 (O_490,N_2961,N_2952);
nand UO_491 (O_491,N_2978,N_2996);
or UO_492 (O_492,N_2976,N_2996);
nand UO_493 (O_493,N_2942,N_2999);
nor UO_494 (O_494,N_2989,N_2998);
nand UO_495 (O_495,N_2975,N_2995);
and UO_496 (O_496,N_2958,N_2972);
or UO_497 (O_497,N_2942,N_2990);
nand UO_498 (O_498,N_2976,N_2962);
xor UO_499 (O_499,N_2964,N_2977);
endmodule