module basic_1500_15000_2000_5_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_655,In_535);
nand U1 (N_1,In_552,In_281);
or U2 (N_2,In_784,In_1017);
nand U3 (N_3,In_1426,In_258);
or U4 (N_4,In_1182,In_116);
and U5 (N_5,In_764,In_686);
or U6 (N_6,In_894,In_423);
and U7 (N_7,In_297,In_488);
or U8 (N_8,In_805,In_1271);
or U9 (N_9,In_804,In_324);
or U10 (N_10,In_1206,In_1181);
nor U11 (N_11,In_68,In_528);
nor U12 (N_12,In_348,In_1115);
nor U13 (N_13,In_1278,In_895);
nor U14 (N_14,In_1214,In_953);
nand U15 (N_15,In_869,In_219);
or U16 (N_16,In_151,In_77);
nor U17 (N_17,In_1338,In_407);
or U18 (N_18,In_1368,In_582);
nand U19 (N_19,In_502,In_768);
nor U20 (N_20,In_1228,In_347);
nand U21 (N_21,In_404,In_1216);
and U22 (N_22,In_903,In_1085);
nor U23 (N_23,In_825,In_388);
xor U24 (N_24,In_451,In_538);
and U25 (N_25,In_1498,In_820);
nand U26 (N_26,In_1298,In_976);
nor U27 (N_27,In_911,In_834);
or U28 (N_28,In_932,In_1264);
nor U29 (N_29,In_1275,In_1412);
or U30 (N_30,In_1185,In_442);
nand U31 (N_31,In_449,In_386);
nor U32 (N_32,In_402,In_844);
or U33 (N_33,In_997,In_1053);
nand U34 (N_34,In_42,In_1337);
or U35 (N_35,In_1048,In_833);
nor U36 (N_36,In_1287,In_958);
nand U37 (N_37,In_26,In_456);
nand U38 (N_38,In_1025,In_1388);
nand U39 (N_39,In_53,In_1478);
or U40 (N_40,In_909,In_1403);
or U41 (N_41,In_419,In_1477);
nand U42 (N_42,In_536,In_479);
or U43 (N_43,In_1193,In_1101);
nand U44 (N_44,In_921,In_1232);
or U45 (N_45,In_271,In_1109);
and U46 (N_46,In_622,In_573);
and U47 (N_47,In_584,In_509);
or U48 (N_48,In_852,In_1459);
nand U49 (N_49,In_1179,In_1496);
or U50 (N_50,In_802,In_485);
nand U51 (N_51,In_1312,In_890);
or U52 (N_52,In_1333,In_865);
nor U53 (N_53,In_856,In_530);
or U54 (N_54,In_1261,In_154);
nor U55 (N_55,In_177,In_689);
nand U56 (N_56,In_999,In_1421);
or U57 (N_57,In_195,In_1133);
xor U58 (N_58,In_356,In_62);
and U59 (N_59,In_170,In_306);
and U60 (N_60,In_902,In_1094);
nor U61 (N_61,In_1032,In_13);
nand U62 (N_62,In_525,In_1370);
and U63 (N_63,In_631,In_832);
or U64 (N_64,In_1313,In_827);
nor U65 (N_65,In_105,In_357);
nor U66 (N_66,In_632,In_648);
and U67 (N_67,In_10,In_685);
xnor U68 (N_68,In_720,In_1082);
nor U69 (N_69,In_1122,In_1146);
nand U70 (N_70,In_123,In_916);
and U71 (N_71,In_938,In_524);
and U72 (N_72,In_1078,In_668);
and U73 (N_73,In_490,In_1325);
nand U74 (N_74,In_973,In_311);
or U75 (N_75,In_100,In_396);
nand U76 (N_76,In_421,In_948);
nor U77 (N_77,In_907,In_1425);
nor U78 (N_78,In_1492,In_194);
nand U79 (N_79,In_30,In_1162);
or U80 (N_80,In_355,In_1174);
and U81 (N_81,In_82,In_1359);
nand U82 (N_82,In_1307,In_83);
nor U83 (N_83,In_893,In_694);
or U84 (N_84,In_98,In_1234);
nand U85 (N_85,In_307,In_558);
nor U86 (N_86,In_724,In_63);
nor U87 (N_87,In_46,In_149);
xnor U88 (N_88,In_1279,In_1166);
nand U89 (N_89,In_366,In_203);
nor U90 (N_90,In_1090,In_130);
and U91 (N_91,In_540,In_70);
xnor U92 (N_92,In_732,In_708);
nand U93 (N_93,In_1251,In_1341);
and U94 (N_94,In_1246,In_437);
or U95 (N_95,In_1176,In_1314);
or U96 (N_96,In_1355,In_1168);
nor U97 (N_97,In_596,In_1343);
or U98 (N_98,In_1473,In_1250);
and U99 (N_99,In_36,In_494);
and U100 (N_100,In_572,In_1136);
and U101 (N_101,In_405,In_1449);
nand U102 (N_102,In_433,In_860);
and U103 (N_103,In_137,In_445);
nor U104 (N_104,In_164,In_1083);
and U105 (N_105,In_216,In_108);
nand U106 (N_106,In_1366,In_1469);
xnor U107 (N_107,In_246,In_415);
nor U108 (N_108,In_308,In_735);
nand U109 (N_109,In_291,In_606);
and U110 (N_110,In_889,In_369);
or U111 (N_111,In_150,In_1494);
and U112 (N_112,In_168,In_393);
and U113 (N_113,In_1191,In_787);
nor U114 (N_114,In_892,In_910);
or U115 (N_115,In_942,In_153);
and U116 (N_116,In_770,In_736);
nand U117 (N_117,In_416,In_1143);
or U118 (N_118,In_1467,In_862);
and U119 (N_119,In_132,In_1295);
nor U120 (N_120,In_1060,In_237);
nand U121 (N_121,In_481,In_1223);
xnor U122 (N_122,In_568,In_672);
nand U123 (N_123,In_794,In_1153);
nor U124 (N_124,In_1108,In_522);
and U125 (N_125,In_1335,In_1192);
nand U126 (N_126,In_33,In_217);
and U127 (N_127,In_891,In_1224);
nor U128 (N_128,In_319,In_830);
or U129 (N_129,In_813,In_377);
nor U130 (N_130,In_1465,In_1126);
and U131 (N_131,In_586,In_915);
nor U132 (N_132,In_1009,In_197);
or U133 (N_133,In_460,In_330);
nor U134 (N_134,In_495,In_811);
and U135 (N_135,In_1006,In_1015);
nand U136 (N_136,In_293,In_1242);
nand U137 (N_137,In_854,In_1407);
and U138 (N_138,In_1187,In_1356);
nand U139 (N_139,In_145,In_139);
nand U140 (N_140,In_1054,In_702);
or U141 (N_141,In_290,In_1297);
or U142 (N_142,In_66,In_1437);
nor U143 (N_143,In_1117,In_1020);
and U144 (N_144,In_1257,In_96);
or U145 (N_145,In_409,In_230);
nor U146 (N_146,In_1064,In_1172);
xnor U147 (N_147,In_635,In_607);
nor U148 (N_148,In_256,In_111);
and U149 (N_149,In_165,In_1120);
nor U150 (N_150,In_774,In_1189);
or U151 (N_151,In_1266,In_273);
nand U152 (N_152,In_269,In_174);
and U153 (N_153,In_619,In_43);
nand U154 (N_154,In_1180,In_876);
xor U155 (N_155,In_615,In_1353);
nand U156 (N_156,In_993,In_904);
nor U157 (N_157,In_384,In_268);
and U158 (N_158,In_920,In_969);
nor U159 (N_159,In_341,In_1365);
and U160 (N_160,In_86,In_581);
nor U161 (N_161,In_812,In_294);
or U162 (N_162,In_80,In_714);
or U163 (N_163,In_1023,In_692);
or U164 (N_164,In_842,In_730);
xor U165 (N_165,In_381,In_867);
nand U166 (N_166,In_1345,In_400);
and U167 (N_167,In_641,In_674);
nand U168 (N_168,In_143,In_122);
and U169 (N_169,In_1373,In_767);
or U170 (N_170,In_1489,In_576);
and U171 (N_171,In_444,In_262);
nor U172 (N_172,In_1210,In_778);
and U173 (N_173,In_761,In_241);
and U174 (N_174,In_851,In_799);
nor U175 (N_175,In_472,In_1288);
nand U176 (N_176,In_1034,In_288);
xnor U177 (N_177,In_1079,In_140);
nor U178 (N_178,In_979,In_747);
and U179 (N_179,In_253,In_1317);
and U180 (N_180,In_1376,In_331);
xnor U181 (N_181,In_1367,In_984);
nor U182 (N_182,In_777,In_380);
and U183 (N_183,In_1169,In_275);
xnor U184 (N_184,In_1039,In_191);
nor U185 (N_185,In_299,In_908);
nand U186 (N_186,In_226,In_376);
or U187 (N_187,In_1374,In_335);
or U188 (N_188,In_157,In_1051);
nand U189 (N_189,In_874,In_977);
nor U190 (N_190,In_700,In_541);
and U191 (N_191,In_960,In_1480);
nand U192 (N_192,In_49,In_387);
nor U193 (N_193,In_1419,In_1091);
and U194 (N_194,In_755,In_1123);
nand U195 (N_195,In_414,In_1424);
nor U196 (N_196,In_283,In_469);
or U197 (N_197,In_1453,In_882);
nand U198 (N_198,In_225,In_1217);
and U199 (N_199,In_295,In_1003);
and U200 (N_200,In_662,In_629);
and U201 (N_201,In_1385,In_658);
and U202 (N_202,In_1022,In_37);
nand U203 (N_203,In_630,In_688);
or U204 (N_204,In_232,In_775);
or U205 (N_205,In_1225,In_944);
xnor U206 (N_206,In_1429,In_1215);
xnor U207 (N_207,In_1147,In_1229);
nand U208 (N_208,In_782,In_554);
or U209 (N_209,In_507,In_744);
and U210 (N_210,In_261,In_990);
nor U211 (N_211,In_408,In_871);
xor U212 (N_212,In_801,In_360);
nor U213 (N_213,In_1283,In_721);
and U214 (N_214,In_881,In_1445);
nor U215 (N_215,In_248,In_1381);
and U216 (N_216,In_1163,In_521);
or U217 (N_217,In_265,In_468);
nand U218 (N_218,In_41,In_925);
nand U219 (N_219,In_710,In_1004);
nand U220 (N_220,In_503,In_1451);
or U221 (N_221,In_1326,In_266);
nand U222 (N_222,In_553,In_762);
and U223 (N_223,In_1139,In_455);
or U224 (N_224,In_337,In_305);
nor U225 (N_225,In_873,In_1141);
or U226 (N_226,In_900,In_315);
nand U227 (N_227,In_1131,In_185);
nand U228 (N_228,In_382,In_1482);
and U229 (N_229,In_1301,In_814);
or U230 (N_230,In_38,In_1292);
and U231 (N_231,In_189,In_1463);
nor U232 (N_232,In_85,In_564);
or U233 (N_233,In_646,In_7);
and U234 (N_234,In_642,In_363);
and U235 (N_235,In_975,In_312);
nor U236 (N_236,In_872,In_1285);
and U237 (N_237,In_1235,In_625);
and U238 (N_238,In_660,In_1401);
nand U239 (N_239,In_1427,In_698);
nand U240 (N_240,In_1018,In_310);
or U241 (N_241,In_1436,In_1156);
and U242 (N_242,In_1331,In_1164);
nand U243 (N_243,In_547,In_901);
and U244 (N_244,In_87,In_284);
or U245 (N_245,In_1442,In_201);
or U246 (N_246,In_1397,In_850);
nand U247 (N_247,In_543,In_167);
or U248 (N_248,In_1487,In_1342);
or U249 (N_249,In_722,In_716);
or U250 (N_250,In_1222,In_613);
nand U251 (N_251,In_78,In_438);
and U252 (N_252,In_304,In_1323);
or U253 (N_253,In_459,In_1396);
or U254 (N_254,In_1076,In_487);
nand U255 (N_255,In_1457,In_542);
nand U256 (N_256,In_886,In_647);
nor U257 (N_257,In_1204,In_705);
nand U258 (N_258,In_1456,In_649);
xnor U259 (N_259,In_179,In_440);
and U260 (N_260,In_412,In_1072);
and U261 (N_261,In_486,In_796);
xnor U262 (N_262,In_371,In_788);
and U263 (N_263,In_1304,In_952);
or U264 (N_264,In_1227,In_922);
xnor U265 (N_265,In_967,In_828);
nand U266 (N_266,In_97,In_501);
or U267 (N_267,In_950,In_354);
or U268 (N_268,In_336,In_417);
nor U269 (N_269,In_652,In_756);
and U270 (N_270,In_1272,In_1140);
and U271 (N_271,In_220,In_1357);
or U272 (N_272,In_1371,In_949);
and U273 (N_273,In_1208,In_994);
and U274 (N_274,In_25,In_598);
nand U275 (N_275,In_144,In_379);
or U276 (N_276,In_1086,In_1254);
nor U277 (N_277,In_592,In_588);
nand U278 (N_278,In_1431,In_1132);
xor U279 (N_279,In_966,In_654);
nand U280 (N_280,In_1050,In_1065);
or U281 (N_281,In_1081,In_1479);
or U282 (N_282,In_657,In_726);
nand U283 (N_283,In_771,In_3);
nor U284 (N_284,In_1256,In_1125);
or U285 (N_285,In_936,In_845);
or U286 (N_286,In_389,In_21);
nand U287 (N_287,In_537,In_439);
and U288 (N_288,In_411,In_699);
nor U289 (N_289,In_656,In_651);
xor U290 (N_290,In_1190,In_1061);
or U291 (N_291,In_1361,In_741);
nor U292 (N_292,In_680,In_260);
and U293 (N_293,In_1226,In_1387);
or U294 (N_294,In_687,In_1339);
or U295 (N_295,In_1096,In_90);
and U296 (N_296,In_1280,In_595);
and U297 (N_297,In_992,In_339);
xnor U298 (N_298,In_465,In_309);
or U299 (N_299,In_1201,In_684);
and U300 (N_300,In_1129,In_988);
and U301 (N_301,In_110,In_579);
or U302 (N_302,In_323,In_514);
nand U303 (N_303,In_640,In_670);
nand U304 (N_304,In_769,In_1438);
and U305 (N_305,In_798,In_561);
xnor U306 (N_306,In_559,In_218);
nand U307 (N_307,In_1055,In_1399);
nand U308 (N_308,In_156,In_757);
or U309 (N_309,In_1276,In_54);
or U310 (N_310,In_1230,In_1466);
or U311 (N_311,In_51,In_557);
nand U312 (N_312,In_1268,In_9);
nor U313 (N_313,In_1071,In_1319);
and U314 (N_314,In_1499,In_951);
and U315 (N_315,In_1238,In_192);
nor U316 (N_316,In_1041,In_1493);
and U317 (N_317,In_1178,In_1443);
and U318 (N_318,In_752,In_180);
xor U319 (N_319,In_1395,In_1416);
nand U320 (N_320,In_1218,In_986);
and U321 (N_321,In_600,In_527);
or U322 (N_322,In_780,In_1252);
nand U323 (N_323,In_677,In_864);
and U324 (N_324,In_974,In_1379);
or U325 (N_325,In_120,In_106);
nor U326 (N_326,In_597,In_663);
nand U327 (N_327,In_962,In_879);
and U328 (N_328,In_758,In_1000);
nor U329 (N_329,In_718,In_1130);
xor U330 (N_330,In_797,In_1236);
or U331 (N_331,In_1111,In_1336);
or U332 (N_332,In_94,In_238);
nand U333 (N_333,In_512,In_1121);
xor U334 (N_334,In_280,In_493);
and U335 (N_335,In_1349,In_1057);
and U336 (N_336,In_534,In_1420);
nor U337 (N_337,In_1102,In_34);
nor U338 (N_338,In_1274,In_76);
nand U339 (N_339,In_1321,In_461);
nor U340 (N_340,In_127,In_239);
or U341 (N_341,In_743,In_1157);
nor U342 (N_342,In_1046,In_661);
nand U343 (N_343,In_1290,In_603);
and U344 (N_344,In_751,In_996);
nor U345 (N_345,In_803,In_448);
nor U346 (N_346,In_1471,In_591);
nor U347 (N_347,In_399,In_102);
and U348 (N_348,In_861,In_420);
nand U349 (N_349,In_945,In_723);
nand U350 (N_350,In_413,In_1422);
nor U351 (N_351,In_1155,In_1033);
nor U352 (N_352,In_1294,In_637);
nor U353 (N_353,In_683,In_759);
nand U354 (N_354,In_1188,In_822);
nor U355 (N_355,In_52,In_1028);
or U356 (N_356,In_274,In_224);
or U357 (N_357,In_1398,In_1144);
nor U358 (N_358,In_1291,In_859);
or U359 (N_359,In_624,In_1194);
nor U360 (N_360,In_1418,In_1151);
nand U361 (N_361,In_551,In_482);
nor U362 (N_362,In_1198,In_1106);
nor U363 (N_363,In_807,In_362);
nor U364 (N_364,In_887,In_772);
nand U365 (N_365,In_749,In_590);
nor U366 (N_366,In_313,In_334);
nor U367 (N_367,In_1148,In_678);
or U368 (N_368,In_1383,In_270);
nand U369 (N_369,In_1423,In_121);
or U370 (N_370,In_286,In_4);
xnor U371 (N_371,In_231,In_571);
or U372 (N_372,In_1249,In_1152);
nand U373 (N_373,In_429,In_817);
nor U374 (N_374,In_212,In_1415);
or U375 (N_375,In_1002,In_113);
nor U376 (N_376,In_888,In_1363);
or U377 (N_377,In_245,In_555);
and U378 (N_378,In_843,In_653);
xor U379 (N_379,In_40,In_352);
or U380 (N_380,In_228,In_1461);
nand U381 (N_381,In_816,In_991);
or U382 (N_382,In_240,In_322);
and U383 (N_383,In_620,In_972);
nor U384 (N_384,In_866,In_1042);
and U385 (N_385,In_931,In_957);
or U386 (N_386,In_1329,In_1052);
or U387 (N_387,In_81,In_981);
or U388 (N_388,In_1328,In_1432);
xnor U389 (N_389,In_329,In_659);
or U390 (N_390,In_466,In_518);
or U391 (N_391,In_1289,In_679);
nor U392 (N_392,In_1233,In_675);
or U393 (N_393,In_1118,In_346);
or U394 (N_394,In_727,In_1137);
or U395 (N_395,In_1265,In_1351);
xor U396 (N_396,In_691,In_385);
xnor U397 (N_397,In_1012,In_390);
nor U398 (N_398,In_1458,In_178);
nand U399 (N_399,In_665,In_1213);
nand U400 (N_400,In_282,In_594);
and U401 (N_401,In_940,In_1391);
nor U402 (N_402,In_474,In_1262);
xnor U403 (N_403,In_673,In_1200);
nand U404 (N_404,In_546,In_878);
and U405 (N_405,In_202,In_325);
or U406 (N_406,In_1142,In_792);
or U407 (N_407,In_358,In_126);
nor U408 (N_408,In_955,In_1497);
nand U409 (N_409,In_27,In_1134);
nor U410 (N_410,In_574,In_134);
and U411 (N_411,In_112,In_221);
nand U412 (N_412,In_61,In_549);
xor U413 (N_413,In_585,In_835);
nor U414 (N_414,In_1293,In_1400);
and U415 (N_415,In_162,In_877);
nand U416 (N_416,In_896,In_913);
xor U417 (N_417,In_14,In_707);
nor U418 (N_418,In_1177,In_1145);
xnor U419 (N_419,In_1173,In_72);
and U420 (N_420,In_434,In_58);
or U421 (N_421,In_454,In_841);
or U422 (N_422,In_158,In_183);
and U423 (N_423,In_808,In_351);
nand U424 (N_424,In_457,In_750);
nand U425 (N_425,In_1447,In_129);
nor U426 (N_426,In_578,In_905);
and U427 (N_427,In_939,In_2);
and U428 (N_428,In_1462,In_1452);
nand U429 (N_429,In_1460,In_884);
nand U430 (N_430,In_252,In_166);
or U431 (N_431,In_148,In_298);
nor U432 (N_432,In_0,In_15);
and U433 (N_433,In_234,In_1043);
nor U434 (N_434,In_318,In_941);
nor U435 (N_435,In_1026,In_463);
nor U436 (N_436,In_1414,In_1116);
nor U437 (N_437,In_1024,In_1001);
xor U438 (N_438,In_519,In_1089);
nor U439 (N_439,In_806,In_181);
nand U440 (N_440,In_1183,In_1488);
nand U441 (N_441,In_163,In_147);
or U442 (N_442,In_853,In_1303);
or U443 (N_443,In_608,In_1175);
nand U444 (N_444,In_633,In_1170);
nor U445 (N_445,In_8,In_489);
and U446 (N_446,In_483,In_359);
or U447 (N_447,In_99,In_1029);
or U448 (N_448,In_1197,In_760);
or U449 (N_449,In_75,In_497);
and U450 (N_450,In_1092,In_365);
or U451 (N_451,In_16,In_863);
nor U452 (N_452,In_985,In_1481);
nor U453 (N_453,In_1350,In_636);
nand U454 (N_454,In_1240,In_1375);
or U455 (N_455,In_471,In_1160);
and U456 (N_456,In_715,In_31);
nand U457 (N_457,In_1430,In_847);
xnor U458 (N_458,In_676,In_343);
xnor U459 (N_459,In_243,In_161);
nor U460 (N_460,In_1411,In_826);
nor U461 (N_461,In_701,In_1327);
nand U462 (N_462,In_169,In_198);
nand U463 (N_463,In_1062,In_1404);
xor U464 (N_464,In_621,In_184);
nand U465 (N_465,In_119,In_109);
nand U466 (N_466,In_289,In_589);
and U467 (N_467,In_1409,In_114);
xor U468 (N_468,In_943,In_435);
and U469 (N_469,In_84,In_961);
nand U470 (N_470,In_79,In_55);
and U471 (N_471,In_783,In_1073);
nor U472 (N_472,In_781,In_666);
nand U473 (N_473,In_1058,In_510);
and U474 (N_474,In_1069,In_508);
nand U475 (N_475,In_171,In_1195);
and U476 (N_476,In_1455,In_645);
xor U477 (N_477,In_569,In_11);
or U478 (N_478,In_1007,In_906);
nand U479 (N_479,In_1241,In_210);
nand U480 (N_480,In_831,In_550);
nor U481 (N_481,In_855,In_1159);
xor U482 (N_482,In_1282,In_1446);
nor U483 (N_483,In_946,In_930);
nand U484 (N_484,In_1267,In_556);
or U485 (N_485,In_1444,In_1358);
nor U486 (N_486,In_763,In_447);
nor U487 (N_487,In_155,In_1439);
or U488 (N_488,In_1258,In_1309);
nor U489 (N_489,In_965,In_18);
and U490 (N_490,In_350,In_917);
or U491 (N_491,In_731,In_247);
nand U492 (N_492,In_1410,In_1346);
or U493 (N_493,In_1302,In_1348);
nor U494 (N_494,In_136,In_565);
or U495 (N_495,In_506,In_1119);
xor U496 (N_496,In_733,In_172);
or U497 (N_497,In_104,In_35);
and U498 (N_498,In_1382,In_623);
nand U499 (N_499,In_1105,In_250);
nor U500 (N_500,In_1296,In_563);
nor U501 (N_501,In_1113,In_74);
or U502 (N_502,In_5,In_1202);
and U503 (N_503,In_924,In_837);
nor U504 (N_504,In_1372,In_1435);
or U505 (N_505,In_1299,In_264);
nand U506 (N_506,In_1027,In_492);
and U507 (N_507,In_819,In_712);
or U508 (N_508,In_278,In_316);
nor U509 (N_509,In_345,In_968);
or U510 (N_510,In_1286,In_103);
or U511 (N_511,In_1114,In_317);
or U512 (N_512,In_1138,In_374);
or U513 (N_513,In_251,In_327);
or U514 (N_514,In_1205,In_182);
and U515 (N_515,In_840,In_328);
or U516 (N_516,In_1088,In_314);
xor U517 (N_517,In_1011,In_395);
nor U518 (N_518,In_124,In_361);
or U519 (N_519,In_511,In_899);
nor U520 (N_520,In_664,In_1248);
nor U521 (N_521,In_593,In_1247);
and U522 (N_522,In_987,In_272);
nand U523 (N_523,In_539,In_818);
nand U524 (N_524,In_186,In_809);
nand U525 (N_525,In_681,In_1450);
and U526 (N_526,In_477,In_406);
or U527 (N_527,In_1104,In_418);
or U528 (N_528,In_276,In_1402);
nand U529 (N_529,In_995,In_233);
nand U530 (N_530,In_709,In_279);
nor U531 (N_531,In_779,In_650);
or U532 (N_532,In_1386,In_566);
xnor U533 (N_533,In_200,In_410);
nor U534 (N_534,In_333,In_1310);
nand U535 (N_535,In_734,In_1334);
xor U536 (N_536,In_1253,In_443);
xor U537 (N_537,In_934,In_1209);
nand U538 (N_538,In_173,In_1047);
nor U539 (N_539,In_602,In_1199);
xnor U540 (N_540,In_1038,In_1378);
or U541 (N_541,In_146,In_1220);
nand U542 (N_542,In_669,In_1080);
and U543 (N_543,In_285,In_1084);
and U544 (N_544,In_473,In_32);
nor U545 (N_545,In_858,In_1270);
or U546 (N_546,In_65,In_131);
nor U547 (N_547,In_257,In_1219);
and U548 (N_548,In_926,In_728);
nor U549 (N_549,In_207,In_342);
nor U550 (N_550,In_898,In_821);
or U551 (N_551,In_1394,In_22);
nor U552 (N_552,In_242,In_1077);
or U553 (N_553,In_1428,In_128);
xnor U554 (N_554,In_23,In_857);
nor U555 (N_555,In_452,In_790);
nand U556 (N_556,In_627,In_1390);
nand U557 (N_557,In_56,In_703);
and U558 (N_558,In_773,In_1040);
nor U559 (N_559,In_222,In_1324);
nand U560 (N_560,In_745,In_970);
or U561 (N_561,In_462,In_1221);
xnor U562 (N_562,In_725,In_159);
nor U563 (N_563,In_254,In_1016);
nand U564 (N_564,In_338,In_259);
nand U565 (N_565,In_1049,In_671);
nand U566 (N_566,In_368,In_1008);
nor U567 (N_567,In_1269,In_875);
xnor U568 (N_568,In_19,In_800);
and U569 (N_569,In_1149,In_667);
nor U570 (N_570,In_432,In_142);
and U571 (N_571,In_1408,In_523);
or U572 (N_572,In_634,In_378);
or U573 (N_573,In_836,In_918);
xnor U574 (N_574,In_526,In_24);
nor U575 (N_575,In_1005,In_1360);
and U576 (N_576,In_1044,In_1259);
nor U577 (N_577,In_209,In_141);
xor U578 (N_578,In_1380,In_639);
and U579 (N_579,In_383,In_1161);
nand U580 (N_580,In_1237,In_1485);
nor U581 (N_581,In_1330,In_1263);
nor U582 (N_582,In_971,In_1068);
nor U583 (N_583,In_560,In_880);
xnor U584 (N_584,In_1306,In_1318);
nor U585 (N_585,In_344,In_1203);
nand U586 (N_586,In_544,In_989);
nand U587 (N_587,In_101,In_1167);
nor U588 (N_588,In_504,In_321);
or U589 (N_589,In_978,In_364);
and U590 (N_590,In_1475,In_263);
or U591 (N_591,In_176,In_815);
xnor U592 (N_592,In_738,In_998);
xor U593 (N_593,In_403,In_643);
or U594 (N_594,In_1135,In_1243);
or U595 (N_595,In_1124,In_824);
or U596 (N_596,In_199,In_59);
xor U597 (N_597,In_1244,In_1472);
or U598 (N_598,In_187,In_107);
nand U599 (N_599,In_287,In_255);
nand U600 (N_600,In_391,In_1483);
nor U601 (N_601,In_964,In_1103);
or U602 (N_602,In_1030,In_422);
and U603 (N_603,In_1308,In_1434);
nor U604 (N_604,In_614,In_425);
xor U605 (N_605,In_12,In_1448);
or U606 (N_606,In_138,In_1171);
and U607 (N_607,In_60,In_244);
and U608 (N_608,In_50,In_789);
or U609 (N_609,In_742,In_1031);
or U610 (N_610,In_303,In_436);
nand U611 (N_611,In_1316,In_870);
nand U612 (N_612,In_1255,In_1186);
nand U613 (N_613,In_980,In_118);
or U614 (N_614,In_426,In_513);
and U615 (N_615,In_545,In_92);
and U616 (N_616,In_93,In_706);
or U617 (N_617,In_1245,In_476);
and U618 (N_618,In_480,In_1491);
xnor U619 (N_619,In_64,In_580);
or U620 (N_620,In_496,In_17);
or U621 (N_621,In_223,In_193);
or U622 (N_622,In_737,In_117);
or U623 (N_623,In_296,In_39);
or U624 (N_624,In_1484,In_301);
nor U625 (N_625,In_1154,In_793);
and U626 (N_626,In_1100,In_1212);
nand U627 (N_627,In_713,In_1045);
or U628 (N_628,In_601,In_227);
and U629 (N_629,In_532,In_1417);
xnor U630 (N_630,In_57,In_1184);
or U631 (N_631,In_441,In_1464);
nand U632 (N_632,In_1150,In_498);
and U633 (N_633,In_605,In_729);
nor U634 (N_634,In_928,In_1158);
or U635 (N_635,In_1098,In_611);
and U636 (N_636,In_567,In_1433);
nand U637 (N_637,In_67,In_1281);
xnor U638 (N_638,In_954,In_267);
and U639 (N_639,In_91,In_125);
or U640 (N_640,In_933,In_823);
nand U641 (N_641,In_475,In_353);
or U642 (N_642,In_982,In_927);
and U643 (N_643,In_1354,In_458);
nand U644 (N_644,In_89,In_587);
nand U645 (N_645,In_849,In_533);
or U646 (N_646,In_214,In_947);
and U647 (N_647,In_912,In_20);
and U648 (N_648,In_776,In_1300);
or U649 (N_649,In_484,In_95);
or U650 (N_650,In_1273,In_326);
nor U651 (N_651,In_88,In_1490);
or U652 (N_652,In_548,In_609);
xor U653 (N_653,In_848,In_711);
nand U654 (N_654,In_914,In_215);
or U655 (N_655,In_919,In_1093);
nand U656 (N_656,In_48,In_372);
and U657 (N_657,In_1389,In_1441);
nand U658 (N_658,In_1392,In_1128);
nand U659 (N_659,In_1036,In_229);
nand U660 (N_660,In_446,In_401);
and U661 (N_661,In_204,In_746);
nor U662 (N_662,In_577,In_517);
or U663 (N_663,In_1231,In_1066);
and U664 (N_664,In_152,In_29);
and U665 (N_665,In_1284,In_320);
nand U666 (N_666,In_765,In_616);
or U667 (N_667,In_1305,In_375);
xnor U668 (N_668,In_428,In_367);
nand U669 (N_669,In_575,In_935);
or U670 (N_670,In_520,In_1311);
xor U671 (N_671,In_188,In_1239);
and U672 (N_672,In_397,In_846);
nand U673 (N_673,In_300,In_1107);
or U674 (N_674,In_531,In_697);
nor U675 (N_675,In_69,In_349);
or U676 (N_676,In_740,In_1352);
nand U677 (N_677,In_205,In_160);
nor U678 (N_678,In_1468,In_838);
xnor U679 (N_679,In_505,In_638);
xor U680 (N_680,In_500,In_236);
nand U681 (N_681,In_467,In_529);
or U682 (N_682,In_1405,In_424);
and U683 (N_683,In_1440,In_1087);
and U684 (N_684,In_719,In_431);
xnor U685 (N_685,In_430,In_753);
and U686 (N_686,In_478,In_1364);
or U687 (N_687,In_516,In_44);
nor U688 (N_688,In_373,In_612);
and U689 (N_689,In_427,In_135);
nand U690 (N_690,In_1495,In_1);
nand U691 (N_691,In_766,In_1377);
or U692 (N_692,In_73,In_213);
nor U693 (N_693,In_617,In_883);
and U694 (N_694,In_983,In_292);
or U695 (N_695,In_1059,In_1362);
nor U696 (N_696,In_1019,In_717);
nor U697 (N_697,In_1260,In_1035);
nor U698 (N_698,In_453,In_1406);
nand U699 (N_699,In_133,In_332);
and U700 (N_700,In_175,In_610);
and U701 (N_701,In_1369,In_470);
nand U702 (N_702,In_206,In_1277);
and U703 (N_703,In_1127,In_515);
nand U704 (N_704,In_929,In_1021);
xnor U705 (N_705,In_583,In_1332);
xor U706 (N_706,In_839,In_618);
and U707 (N_707,In_696,In_211);
nand U708 (N_708,In_1454,In_695);
or U709 (N_709,In_1322,In_1070);
or U710 (N_710,In_464,In_1112);
or U711 (N_711,In_47,In_249);
and U712 (N_712,In_1099,In_1010);
nor U713 (N_713,In_690,In_1095);
nand U714 (N_714,In_795,In_786);
and U715 (N_715,In_277,In_1110);
or U716 (N_716,In_739,In_754);
nand U717 (N_717,In_392,In_302);
nor U718 (N_718,In_1486,In_1207);
and U719 (N_719,In_6,In_959);
or U720 (N_720,In_810,In_1211);
and U721 (N_721,In_1470,In_748);
xnor U722 (N_722,In_1075,In_604);
nand U723 (N_723,In_704,In_1344);
nor U724 (N_724,In_1347,In_394);
nand U725 (N_725,In_1097,In_682);
or U726 (N_726,In_963,In_937);
nand U727 (N_727,In_693,In_450);
and U728 (N_728,In_562,In_923);
and U729 (N_729,In_791,In_115);
nor U730 (N_730,In_1196,In_897);
or U731 (N_731,In_499,In_370);
or U732 (N_732,In_1013,In_1067);
or U733 (N_733,In_340,In_644);
xnor U734 (N_734,In_190,In_235);
nand U735 (N_735,In_1037,In_1315);
or U736 (N_736,In_1476,In_1474);
nand U737 (N_737,In_1340,In_1320);
nor U738 (N_738,In_956,In_1014);
nand U739 (N_739,In_71,In_868);
xnor U740 (N_740,In_1384,In_599);
or U741 (N_741,In_1393,In_1063);
or U742 (N_742,In_196,In_1413);
nand U743 (N_743,In_45,In_785);
nand U744 (N_744,In_1056,In_885);
and U745 (N_745,In_628,In_1074);
nor U746 (N_746,In_1165,In_491);
and U747 (N_747,In_829,In_626);
or U748 (N_748,In_570,In_398);
nor U749 (N_749,In_28,In_208);
and U750 (N_750,In_776,In_340);
nor U751 (N_751,In_1052,In_1108);
nor U752 (N_752,In_250,In_387);
and U753 (N_753,In_265,In_1407);
nand U754 (N_754,In_806,In_141);
and U755 (N_755,In_1337,In_1064);
and U756 (N_756,In_808,In_384);
or U757 (N_757,In_608,In_1463);
or U758 (N_758,In_203,In_18);
nand U759 (N_759,In_1245,In_603);
xor U760 (N_760,In_740,In_1466);
nor U761 (N_761,In_813,In_18);
and U762 (N_762,In_264,In_1478);
xor U763 (N_763,In_149,In_1069);
nor U764 (N_764,In_1296,In_402);
and U765 (N_765,In_655,In_237);
and U766 (N_766,In_1012,In_177);
xor U767 (N_767,In_1326,In_643);
nor U768 (N_768,In_1132,In_509);
and U769 (N_769,In_1320,In_748);
and U770 (N_770,In_744,In_1160);
nor U771 (N_771,In_694,In_1405);
or U772 (N_772,In_630,In_253);
nand U773 (N_773,In_1146,In_1428);
or U774 (N_774,In_414,In_1102);
xor U775 (N_775,In_1149,In_1237);
nand U776 (N_776,In_1034,In_1124);
xor U777 (N_777,In_795,In_538);
nand U778 (N_778,In_1352,In_465);
nor U779 (N_779,In_668,In_463);
nand U780 (N_780,In_544,In_880);
or U781 (N_781,In_511,In_709);
and U782 (N_782,In_98,In_650);
nand U783 (N_783,In_319,In_282);
xor U784 (N_784,In_1298,In_11);
xnor U785 (N_785,In_904,In_999);
nand U786 (N_786,In_1160,In_1477);
or U787 (N_787,In_235,In_852);
or U788 (N_788,In_1110,In_1458);
xnor U789 (N_789,In_168,In_1237);
and U790 (N_790,In_1134,In_1108);
nand U791 (N_791,In_77,In_82);
and U792 (N_792,In_623,In_686);
or U793 (N_793,In_105,In_579);
xnor U794 (N_794,In_396,In_628);
and U795 (N_795,In_474,In_668);
and U796 (N_796,In_481,In_309);
nand U797 (N_797,In_534,In_728);
or U798 (N_798,In_203,In_1277);
or U799 (N_799,In_298,In_156);
and U800 (N_800,In_1102,In_948);
nor U801 (N_801,In_759,In_974);
and U802 (N_802,In_778,In_1196);
nand U803 (N_803,In_1364,In_301);
nor U804 (N_804,In_913,In_304);
or U805 (N_805,In_1288,In_1048);
and U806 (N_806,In_205,In_783);
nor U807 (N_807,In_944,In_829);
or U808 (N_808,In_940,In_1494);
or U809 (N_809,In_67,In_806);
xor U810 (N_810,In_242,In_55);
or U811 (N_811,In_1073,In_708);
nand U812 (N_812,In_61,In_1034);
xor U813 (N_813,In_25,In_10);
and U814 (N_814,In_18,In_541);
and U815 (N_815,In_319,In_1322);
nor U816 (N_816,In_868,In_1223);
nand U817 (N_817,In_759,In_1349);
and U818 (N_818,In_1156,In_981);
nor U819 (N_819,In_1068,In_25);
or U820 (N_820,In_1482,In_553);
or U821 (N_821,In_455,In_627);
and U822 (N_822,In_1191,In_614);
and U823 (N_823,In_1432,In_793);
and U824 (N_824,In_1246,In_111);
nand U825 (N_825,In_1225,In_1330);
nor U826 (N_826,In_691,In_406);
nand U827 (N_827,In_747,In_1233);
or U828 (N_828,In_216,In_219);
and U829 (N_829,In_1221,In_841);
or U830 (N_830,In_288,In_216);
and U831 (N_831,In_563,In_1026);
or U832 (N_832,In_1031,In_1474);
nor U833 (N_833,In_1204,In_358);
or U834 (N_834,In_572,In_926);
and U835 (N_835,In_362,In_626);
or U836 (N_836,In_127,In_275);
xor U837 (N_837,In_759,In_1033);
xnor U838 (N_838,In_227,In_548);
and U839 (N_839,In_868,In_968);
and U840 (N_840,In_921,In_648);
or U841 (N_841,In_319,In_1346);
or U842 (N_842,In_193,In_1193);
or U843 (N_843,In_1070,In_52);
or U844 (N_844,In_1444,In_821);
nand U845 (N_845,In_1239,In_427);
nor U846 (N_846,In_57,In_978);
nand U847 (N_847,In_1110,In_624);
nand U848 (N_848,In_708,In_198);
nand U849 (N_849,In_1005,In_1001);
or U850 (N_850,In_935,In_1455);
xor U851 (N_851,In_292,In_319);
nor U852 (N_852,In_414,In_934);
xnor U853 (N_853,In_1364,In_1106);
nor U854 (N_854,In_1376,In_515);
nor U855 (N_855,In_390,In_619);
nor U856 (N_856,In_657,In_899);
nor U857 (N_857,In_1261,In_1230);
nand U858 (N_858,In_1453,In_266);
or U859 (N_859,In_1044,In_979);
nor U860 (N_860,In_1473,In_41);
and U861 (N_861,In_539,In_1228);
or U862 (N_862,In_172,In_720);
nand U863 (N_863,In_321,In_978);
xor U864 (N_864,In_1062,In_1286);
nand U865 (N_865,In_1490,In_348);
nand U866 (N_866,In_937,In_385);
nand U867 (N_867,In_958,In_1407);
or U868 (N_868,In_328,In_1100);
or U869 (N_869,In_318,In_160);
nor U870 (N_870,In_1440,In_126);
or U871 (N_871,In_1447,In_1403);
xor U872 (N_872,In_1203,In_1163);
or U873 (N_873,In_1438,In_872);
or U874 (N_874,In_1043,In_970);
nor U875 (N_875,In_1056,In_144);
and U876 (N_876,In_937,In_442);
xnor U877 (N_877,In_1129,In_1132);
xor U878 (N_878,In_256,In_576);
nand U879 (N_879,In_719,In_393);
and U880 (N_880,In_808,In_1364);
nor U881 (N_881,In_312,In_807);
nor U882 (N_882,In_808,In_1235);
xor U883 (N_883,In_403,In_123);
and U884 (N_884,In_1158,In_1030);
and U885 (N_885,In_1073,In_1276);
or U886 (N_886,In_559,In_1184);
and U887 (N_887,In_263,In_1350);
nand U888 (N_888,In_542,In_1086);
nor U889 (N_889,In_1281,In_937);
nor U890 (N_890,In_374,In_283);
nand U891 (N_891,In_1053,In_301);
and U892 (N_892,In_928,In_1083);
nand U893 (N_893,In_112,In_1146);
or U894 (N_894,In_1471,In_1167);
nand U895 (N_895,In_1076,In_516);
nand U896 (N_896,In_799,In_138);
or U897 (N_897,In_1287,In_260);
or U898 (N_898,In_421,In_448);
and U899 (N_899,In_817,In_209);
nand U900 (N_900,In_779,In_8);
and U901 (N_901,In_1317,In_407);
nor U902 (N_902,In_69,In_1242);
and U903 (N_903,In_1242,In_1196);
nand U904 (N_904,In_678,In_133);
xor U905 (N_905,In_1213,In_257);
xnor U906 (N_906,In_1353,In_767);
and U907 (N_907,In_241,In_801);
and U908 (N_908,In_1171,In_1000);
xnor U909 (N_909,In_887,In_1421);
or U910 (N_910,In_541,In_272);
nand U911 (N_911,In_925,In_631);
nor U912 (N_912,In_1267,In_39);
or U913 (N_913,In_524,In_1488);
and U914 (N_914,In_1363,In_942);
nand U915 (N_915,In_17,In_1332);
nand U916 (N_916,In_316,In_960);
nand U917 (N_917,In_164,In_659);
nand U918 (N_918,In_101,In_1297);
nor U919 (N_919,In_1268,In_1467);
or U920 (N_920,In_1379,In_1024);
or U921 (N_921,In_926,In_390);
or U922 (N_922,In_990,In_311);
or U923 (N_923,In_55,In_272);
nand U924 (N_924,In_884,In_877);
nand U925 (N_925,In_1100,In_1087);
or U926 (N_926,In_1326,In_906);
or U927 (N_927,In_52,In_98);
nor U928 (N_928,In_1049,In_1064);
nand U929 (N_929,In_727,In_350);
nor U930 (N_930,In_995,In_351);
or U931 (N_931,In_746,In_1087);
nand U932 (N_932,In_214,In_1315);
and U933 (N_933,In_630,In_430);
nor U934 (N_934,In_370,In_301);
or U935 (N_935,In_686,In_453);
nand U936 (N_936,In_946,In_466);
or U937 (N_937,In_28,In_1045);
or U938 (N_938,In_874,In_212);
nor U939 (N_939,In_87,In_198);
nand U940 (N_940,In_2,In_367);
nor U941 (N_941,In_949,In_618);
or U942 (N_942,In_1474,In_1078);
nand U943 (N_943,In_1261,In_797);
nor U944 (N_944,In_796,In_863);
or U945 (N_945,In_1412,In_779);
nor U946 (N_946,In_756,In_930);
and U947 (N_947,In_137,In_430);
and U948 (N_948,In_1224,In_239);
or U949 (N_949,In_1491,In_1113);
nor U950 (N_950,In_936,In_1471);
nand U951 (N_951,In_232,In_7);
or U952 (N_952,In_166,In_658);
xnor U953 (N_953,In_1344,In_1230);
or U954 (N_954,In_472,In_605);
and U955 (N_955,In_47,In_456);
and U956 (N_956,In_1408,In_399);
nor U957 (N_957,In_970,In_1254);
or U958 (N_958,In_833,In_911);
nor U959 (N_959,In_1348,In_922);
nand U960 (N_960,In_98,In_1300);
and U961 (N_961,In_1037,In_893);
or U962 (N_962,In_829,In_280);
or U963 (N_963,In_179,In_65);
xnor U964 (N_964,In_1263,In_1051);
xnor U965 (N_965,In_233,In_256);
nor U966 (N_966,In_565,In_661);
nor U967 (N_967,In_1223,In_79);
xnor U968 (N_968,In_1184,In_783);
nor U969 (N_969,In_601,In_440);
and U970 (N_970,In_228,In_750);
or U971 (N_971,In_482,In_904);
xnor U972 (N_972,In_1205,In_796);
nor U973 (N_973,In_1435,In_130);
nand U974 (N_974,In_358,In_956);
or U975 (N_975,In_100,In_1440);
xnor U976 (N_976,In_244,In_293);
nor U977 (N_977,In_831,In_824);
nor U978 (N_978,In_1159,In_1441);
xnor U979 (N_979,In_586,In_1127);
nor U980 (N_980,In_1072,In_1182);
and U981 (N_981,In_1496,In_808);
nand U982 (N_982,In_694,In_1120);
and U983 (N_983,In_1431,In_490);
or U984 (N_984,In_58,In_1269);
xnor U985 (N_985,In_517,In_101);
nand U986 (N_986,In_1332,In_1104);
xnor U987 (N_987,In_1187,In_1202);
or U988 (N_988,In_382,In_816);
and U989 (N_989,In_1404,In_679);
or U990 (N_990,In_882,In_969);
xor U991 (N_991,In_143,In_1312);
and U992 (N_992,In_506,In_933);
and U993 (N_993,In_83,In_752);
nor U994 (N_994,In_1400,In_653);
nand U995 (N_995,In_1265,In_1458);
xnor U996 (N_996,In_1223,In_1434);
and U997 (N_997,In_1267,In_1413);
and U998 (N_998,In_503,In_1134);
nor U999 (N_999,In_1134,In_960);
nor U1000 (N_1000,In_1308,In_442);
nor U1001 (N_1001,In_1337,In_151);
and U1002 (N_1002,In_1354,In_167);
or U1003 (N_1003,In_17,In_1471);
nand U1004 (N_1004,In_1358,In_900);
and U1005 (N_1005,In_1344,In_1335);
nor U1006 (N_1006,In_825,In_845);
nor U1007 (N_1007,In_1489,In_41);
or U1008 (N_1008,In_1354,In_1157);
xnor U1009 (N_1009,In_902,In_932);
xnor U1010 (N_1010,In_698,In_486);
nand U1011 (N_1011,In_346,In_1200);
nand U1012 (N_1012,In_142,In_486);
and U1013 (N_1013,In_236,In_1325);
and U1014 (N_1014,In_20,In_169);
nand U1015 (N_1015,In_165,In_927);
nand U1016 (N_1016,In_253,In_49);
nand U1017 (N_1017,In_719,In_554);
and U1018 (N_1018,In_166,In_997);
nand U1019 (N_1019,In_345,In_1382);
and U1020 (N_1020,In_1308,In_17);
and U1021 (N_1021,In_763,In_5);
or U1022 (N_1022,In_530,In_1210);
nand U1023 (N_1023,In_889,In_501);
and U1024 (N_1024,In_155,In_1235);
and U1025 (N_1025,In_129,In_175);
nand U1026 (N_1026,In_981,In_628);
nand U1027 (N_1027,In_642,In_130);
and U1028 (N_1028,In_1130,In_899);
nand U1029 (N_1029,In_760,In_654);
nor U1030 (N_1030,In_758,In_611);
nor U1031 (N_1031,In_232,In_842);
or U1032 (N_1032,In_1106,In_240);
nor U1033 (N_1033,In_1490,In_263);
or U1034 (N_1034,In_1460,In_61);
nor U1035 (N_1035,In_812,In_1232);
and U1036 (N_1036,In_186,In_1133);
and U1037 (N_1037,In_1457,In_1084);
nand U1038 (N_1038,In_635,In_1081);
xnor U1039 (N_1039,In_1301,In_706);
xnor U1040 (N_1040,In_1276,In_1339);
nand U1041 (N_1041,In_591,In_1151);
or U1042 (N_1042,In_901,In_776);
nor U1043 (N_1043,In_1442,In_804);
and U1044 (N_1044,In_1182,In_309);
or U1045 (N_1045,In_1440,In_426);
nand U1046 (N_1046,In_616,In_768);
nor U1047 (N_1047,In_113,In_1424);
or U1048 (N_1048,In_393,In_445);
or U1049 (N_1049,In_1053,In_853);
or U1050 (N_1050,In_1270,In_1195);
and U1051 (N_1051,In_869,In_382);
and U1052 (N_1052,In_508,In_372);
and U1053 (N_1053,In_1492,In_100);
or U1054 (N_1054,In_84,In_404);
or U1055 (N_1055,In_174,In_40);
or U1056 (N_1056,In_1426,In_790);
nor U1057 (N_1057,In_229,In_1129);
nand U1058 (N_1058,In_191,In_633);
or U1059 (N_1059,In_923,In_947);
or U1060 (N_1060,In_964,In_1175);
nor U1061 (N_1061,In_242,In_819);
and U1062 (N_1062,In_174,In_1357);
xnor U1063 (N_1063,In_808,In_184);
or U1064 (N_1064,In_710,In_1349);
xor U1065 (N_1065,In_79,In_883);
xnor U1066 (N_1066,In_1013,In_558);
nand U1067 (N_1067,In_1072,In_48);
nand U1068 (N_1068,In_398,In_1384);
and U1069 (N_1069,In_509,In_686);
and U1070 (N_1070,In_274,In_1133);
xnor U1071 (N_1071,In_0,In_210);
nand U1072 (N_1072,In_1106,In_784);
nand U1073 (N_1073,In_1213,In_878);
and U1074 (N_1074,In_582,In_1160);
or U1075 (N_1075,In_778,In_730);
nor U1076 (N_1076,In_884,In_419);
or U1077 (N_1077,In_742,In_397);
or U1078 (N_1078,In_521,In_100);
or U1079 (N_1079,In_768,In_20);
and U1080 (N_1080,In_1326,In_532);
nand U1081 (N_1081,In_48,In_830);
nor U1082 (N_1082,In_239,In_1406);
xnor U1083 (N_1083,In_659,In_1115);
xor U1084 (N_1084,In_606,In_1266);
nor U1085 (N_1085,In_142,In_156);
nand U1086 (N_1086,In_156,In_556);
nand U1087 (N_1087,In_337,In_264);
nor U1088 (N_1088,In_554,In_873);
or U1089 (N_1089,In_471,In_594);
and U1090 (N_1090,In_1400,In_1004);
or U1091 (N_1091,In_967,In_1082);
or U1092 (N_1092,In_574,In_1444);
xor U1093 (N_1093,In_1432,In_424);
nor U1094 (N_1094,In_251,In_1028);
nand U1095 (N_1095,In_533,In_1343);
or U1096 (N_1096,In_950,In_713);
nor U1097 (N_1097,In_97,In_14);
nor U1098 (N_1098,In_999,In_472);
nand U1099 (N_1099,In_187,In_190);
and U1100 (N_1100,In_1323,In_740);
or U1101 (N_1101,In_711,In_1358);
or U1102 (N_1102,In_1395,In_1181);
nor U1103 (N_1103,In_789,In_478);
and U1104 (N_1104,In_1360,In_293);
and U1105 (N_1105,In_646,In_792);
or U1106 (N_1106,In_260,In_351);
xor U1107 (N_1107,In_570,In_1340);
and U1108 (N_1108,In_894,In_636);
nand U1109 (N_1109,In_1429,In_1409);
or U1110 (N_1110,In_1154,In_417);
nand U1111 (N_1111,In_685,In_459);
and U1112 (N_1112,In_1037,In_1052);
nand U1113 (N_1113,In_855,In_268);
and U1114 (N_1114,In_247,In_501);
or U1115 (N_1115,In_1012,In_424);
or U1116 (N_1116,In_1488,In_870);
nand U1117 (N_1117,In_879,In_875);
nand U1118 (N_1118,In_149,In_817);
and U1119 (N_1119,In_343,In_1497);
nor U1120 (N_1120,In_830,In_1423);
nor U1121 (N_1121,In_466,In_805);
xnor U1122 (N_1122,In_1259,In_1074);
or U1123 (N_1123,In_864,In_1493);
nand U1124 (N_1124,In_498,In_1012);
nand U1125 (N_1125,In_1073,In_1176);
nand U1126 (N_1126,In_1125,In_1346);
or U1127 (N_1127,In_278,In_407);
nand U1128 (N_1128,In_1076,In_753);
and U1129 (N_1129,In_1322,In_623);
and U1130 (N_1130,In_974,In_14);
xnor U1131 (N_1131,In_92,In_1026);
or U1132 (N_1132,In_790,In_1246);
nor U1133 (N_1133,In_803,In_1116);
or U1134 (N_1134,In_1339,In_1000);
nand U1135 (N_1135,In_183,In_952);
and U1136 (N_1136,In_17,In_1282);
and U1137 (N_1137,In_365,In_455);
nor U1138 (N_1138,In_1347,In_951);
or U1139 (N_1139,In_1498,In_1056);
and U1140 (N_1140,In_1401,In_355);
or U1141 (N_1141,In_502,In_389);
and U1142 (N_1142,In_299,In_605);
and U1143 (N_1143,In_396,In_295);
or U1144 (N_1144,In_1486,In_96);
or U1145 (N_1145,In_882,In_124);
nand U1146 (N_1146,In_762,In_1356);
nor U1147 (N_1147,In_434,In_133);
xor U1148 (N_1148,In_1479,In_22);
and U1149 (N_1149,In_371,In_84);
or U1150 (N_1150,In_653,In_1080);
nand U1151 (N_1151,In_1386,In_248);
or U1152 (N_1152,In_985,In_1221);
and U1153 (N_1153,In_101,In_971);
and U1154 (N_1154,In_55,In_376);
nand U1155 (N_1155,In_805,In_170);
nor U1156 (N_1156,In_62,In_78);
nor U1157 (N_1157,In_312,In_582);
nand U1158 (N_1158,In_167,In_1062);
nand U1159 (N_1159,In_487,In_519);
xor U1160 (N_1160,In_33,In_876);
or U1161 (N_1161,In_146,In_359);
and U1162 (N_1162,In_824,In_1382);
nand U1163 (N_1163,In_274,In_1460);
nor U1164 (N_1164,In_262,In_1312);
nor U1165 (N_1165,In_1446,In_848);
or U1166 (N_1166,In_480,In_815);
or U1167 (N_1167,In_46,In_1330);
and U1168 (N_1168,In_87,In_1356);
or U1169 (N_1169,In_1196,In_762);
nor U1170 (N_1170,In_153,In_656);
or U1171 (N_1171,In_56,In_664);
nand U1172 (N_1172,In_1383,In_940);
nand U1173 (N_1173,In_1233,In_157);
nand U1174 (N_1174,In_659,In_1086);
nor U1175 (N_1175,In_904,In_285);
nand U1176 (N_1176,In_957,In_683);
nand U1177 (N_1177,In_1251,In_771);
and U1178 (N_1178,In_410,In_746);
nand U1179 (N_1179,In_1461,In_249);
nor U1180 (N_1180,In_1076,In_532);
xnor U1181 (N_1181,In_1234,In_1111);
and U1182 (N_1182,In_1430,In_1079);
nor U1183 (N_1183,In_1039,In_713);
nand U1184 (N_1184,In_888,In_556);
and U1185 (N_1185,In_684,In_467);
xor U1186 (N_1186,In_1271,In_420);
xnor U1187 (N_1187,In_1191,In_439);
nand U1188 (N_1188,In_428,In_946);
nand U1189 (N_1189,In_291,In_1092);
and U1190 (N_1190,In_86,In_222);
nor U1191 (N_1191,In_564,In_314);
xnor U1192 (N_1192,In_789,In_422);
nor U1193 (N_1193,In_355,In_634);
and U1194 (N_1194,In_1120,In_776);
and U1195 (N_1195,In_1221,In_844);
nand U1196 (N_1196,In_1221,In_81);
and U1197 (N_1197,In_869,In_681);
and U1198 (N_1198,In_712,In_604);
nor U1199 (N_1199,In_759,In_875);
nor U1200 (N_1200,In_188,In_266);
nor U1201 (N_1201,In_1074,In_257);
xor U1202 (N_1202,In_240,In_1325);
and U1203 (N_1203,In_887,In_736);
and U1204 (N_1204,In_398,In_767);
or U1205 (N_1205,In_1032,In_168);
and U1206 (N_1206,In_678,In_250);
and U1207 (N_1207,In_502,In_140);
xnor U1208 (N_1208,In_141,In_305);
and U1209 (N_1209,In_1341,In_466);
nor U1210 (N_1210,In_1092,In_952);
nand U1211 (N_1211,In_708,In_238);
nor U1212 (N_1212,In_843,In_405);
nand U1213 (N_1213,In_255,In_477);
and U1214 (N_1214,In_1029,In_591);
and U1215 (N_1215,In_558,In_1419);
nand U1216 (N_1216,In_797,In_1109);
xnor U1217 (N_1217,In_432,In_547);
and U1218 (N_1218,In_438,In_86);
or U1219 (N_1219,In_1372,In_1437);
or U1220 (N_1220,In_1242,In_1001);
or U1221 (N_1221,In_224,In_629);
and U1222 (N_1222,In_498,In_1095);
nand U1223 (N_1223,In_1092,In_1442);
nor U1224 (N_1224,In_94,In_118);
nor U1225 (N_1225,In_887,In_1213);
nand U1226 (N_1226,In_1077,In_621);
and U1227 (N_1227,In_662,In_373);
or U1228 (N_1228,In_339,In_899);
and U1229 (N_1229,In_1402,In_130);
nand U1230 (N_1230,In_608,In_880);
nand U1231 (N_1231,In_1124,In_228);
and U1232 (N_1232,In_444,In_1118);
nor U1233 (N_1233,In_1117,In_10);
and U1234 (N_1234,In_1328,In_1110);
nand U1235 (N_1235,In_1324,In_740);
and U1236 (N_1236,In_957,In_1362);
nor U1237 (N_1237,In_692,In_1376);
and U1238 (N_1238,In_1430,In_293);
nor U1239 (N_1239,In_1398,In_1002);
or U1240 (N_1240,In_394,In_797);
or U1241 (N_1241,In_393,In_1031);
or U1242 (N_1242,In_1053,In_116);
nor U1243 (N_1243,In_1161,In_143);
and U1244 (N_1244,In_1093,In_796);
nand U1245 (N_1245,In_901,In_355);
nand U1246 (N_1246,In_1416,In_1354);
nand U1247 (N_1247,In_544,In_1304);
nand U1248 (N_1248,In_1498,In_812);
or U1249 (N_1249,In_1335,In_369);
and U1250 (N_1250,In_970,In_752);
or U1251 (N_1251,In_1497,In_293);
or U1252 (N_1252,In_51,In_466);
nand U1253 (N_1253,In_1,In_134);
nand U1254 (N_1254,In_1257,In_622);
nand U1255 (N_1255,In_1313,In_355);
nor U1256 (N_1256,In_813,In_109);
nand U1257 (N_1257,In_579,In_767);
nor U1258 (N_1258,In_938,In_1433);
nor U1259 (N_1259,In_1376,In_1184);
and U1260 (N_1260,In_667,In_615);
and U1261 (N_1261,In_52,In_162);
nor U1262 (N_1262,In_259,In_30);
xnor U1263 (N_1263,In_187,In_1241);
xor U1264 (N_1264,In_1412,In_781);
nor U1265 (N_1265,In_552,In_815);
nor U1266 (N_1266,In_888,In_531);
nor U1267 (N_1267,In_1327,In_700);
nor U1268 (N_1268,In_754,In_501);
and U1269 (N_1269,In_195,In_1289);
and U1270 (N_1270,In_62,In_858);
or U1271 (N_1271,In_960,In_531);
xnor U1272 (N_1272,In_544,In_753);
nand U1273 (N_1273,In_1339,In_251);
nand U1274 (N_1274,In_789,In_529);
or U1275 (N_1275,In_623,In_1157);
or U1276 (N_1276,In_257,In_1145);
nand U1277 (N_1277,In_1225,In_215);
and U1278 (N_1278,In_1412,In_1473);
or U1279 (N_1279,In_946,In_415);
and U1280 (N_1280,In_350,In_394);
xnor U1281 (N_1281,In_504,In_882);
or U1282 (N_1282,In_1496,In_958);
xor U1283 (N_1283,In_533,In_322);
nor U1284 (N_1284,In_1323,In_216);
nand U1285 (N_1285,In_723,In_535);
nand U1286 (N_1286,In_1215,In_254);
xor U1287 (N_1287,In_427,In_513);
and U1288 (N_1288,In_1243,In_1289);
nand U1289 (N_1289,In_387,In_935);
nor U1290 (N_1290,In_714,In_1004);
nor U1291 (N_1291,In_249,In_663);
nand U1292 (N_1292,In_276,In_849);
nand U1293 (N_1293,In_883,In_1020);
nand U1294 (N_1294,In_1118,In_1183);
nand U1295 (N_1295,In_786,In_1244);
xnor U1296 (N_1296,In_1415,In_222);
and U1297 (N_1297,In_489,In_1210);
or U1298 (N_1298,In_251,In_689);
nand U1299 (N_1299,In_268,In_46);
nor U1300 (N_1300,In_1075,In_1412);
xnor U1301 (N_1301,In_838,In_1159);
and U1302 (N_1302,In_264,In_517);
nor U1303 (N_1303,In_630,In_1182);
or U1304 (N_1304,In_424,In_1266);
and U1305 (N_1305,In_1476,In_354);
xor U1306 (N_1306,In_1210,In_851);
nor U1307 (N_1307,In_817,In_1160);
nand U1308 (N_1308,In_495,In_1284);
nand U1309 (N_1309,In_1015,In_1385);
or U1310 (N_1310,In_40,In_1274);
or U1311 (N_1311,In_1,In_533);
nand U1312 (N_1312,In_1422,In_616);
or U1313 (N_1313,In_879,In_327);
and U1314 (N_1314,In_164,In_680);
and U1315 (N_1315,In_1110,In_245);
nor U1316 (N_1316,In_686,In_210);
and U1317 (N_1317,In_1471,In_1188);
nand U1318 (N_1318,In_1260,In_1305);
nor U1319 (N_1319,In_736,In_713);
or U1320 (N_1320,In_728,In_863);
or U1321 (N_1321,In_431,In_669);
nand U1322 (N_1322,In_166,In_684);
and U1323 (N_1323,In_1416,In_456);
and U1324 (N_1324,In_626,In_344);
and U1325 (N_1325,In_1045,In_505);
or U1326 (N_1326,In_1245,In_1023);
or U1327 (N_1327,In_1395,In_573);
and U1328 (N_1328,In_1307,In_534);
nand U1329 (N_1329,In_1186,In_208);
and U1330 (N_1330,In_317,In_1036);
or U1331 (N_1331,In_1090,In_44);
and U1332 (N_1332,In_1483,In_81);
nor U1333 (N_1333,In_1357,In_1070);
nor U1334 (N_1334,In_184,In_1);
and U1335 (N_1335,In_645,In_86);
nor U1336 (N_1336,In_1237,In_179);
nand U1337 (N_1337,In_527,In_1431);
and U1338 (N_1338,In_737,In_458);
nor U1339 (N_1339,In_602,In_1479);
xnor U1340 (N_1340,In_435,In_84);
nor U1341 (N_1341,In_213,In_224);
nand U1342 (N_1342,In_1057,In_1211);
or U1343 (N_1343,In_1345,In_1312);
or U1344 (N_1344,In_10,In_898);
and U1345 (N_1345,In_373,In_140);
nor U1346 (N_1346,In_211,In_509);
nand U1347 (N_1347,In_1361,In_1373);
xor U1348 (N_1348,In_985,In_304);
and U1349 (N_1349,In_1012,In_959);
nand U1350 (N_1350,In_359,In_1126);
nand U1351 (N_1351,In_1073,In_1228);
and U1352 (N_1352,In_1388,In_1380);
and U1353 (N_1353,In_370,In_206);
and U1354 (N_1354,In_859,In_452);
nor U1355 (N_1355,In_229,In_541);
nor U1356 (N_1356,In_1486,In_1435);
and U1357 (N_1357,In_1148,In_477);
or U1358 (N_1358,In_1082,In_595);
and U1359 (N_1359,In_94,In_444);
nor U1360 (N_1360,In_865,In_336);
or U1361 (N_1361,In_485,In_1463);
xor U1362 (N_1362,In_456,In_100);
nand U1363 (N_1363,In_1430,In_1);
nand U1364 (N_1364,In_1413,In_1331);
nor U1365 (N_1365,In_1189,In_1416);
nor U1366 (N_1366,In_82,In_400);
or U1367 (N_1367,In_1442,In_268);
and U1368 (N_1368,In_781,In_1432);
and U1369 (N_1369,In_1413,In_189);
and U1370 (N_1370,In_1005,In_544);
and U1371 (N_1371,In_902,In_454);
nor U1372 (N_1372,In_788,In_1251);
and U1373 (N_1373,In_407,In_437);
nor U1374 (N_1374,In_1074,In_180);
nor U1375 (N_1375,In_1191,In_1402);
or U1376 (N_1376,In_1378,In_1351);
or U1377 (N_1377,In_898,In_1150);
xnor U1378 (N_1378,In_7,In_653);
nor U1379 (N_1379,In_1491,In_17);
nand U1380 (N_1380,In_1337,In_563);
nand U1381 (N_1381,In_102,In_843);
and U1382 (N_1382,In_359,In_752);
nand U1383 (N_1383,In_648,In_600);
or U1384 (N_1384,In_944,In_1081);
nor U1385 (N_1385,In_392,In_529);
nand U1386 (N_1386,In_605,In_1192);
nor U1387 (N_1387,In_1365,In_1272);
and U1388 (N_1388,In_637,In_984);
nor U1389 (N_1389,In_205,In_1477);
nand U1390 (N_1390,In_355,In_161);
or U1391 (N_1391,In_215,In_1200);
and U1392 (N_1392,In_357,In_1439);
and U1393 (N_1393,In_1434,In_1333);
nor U1394 (N_1394,In_1177,In_931);
or U1395 (N_1395,In_1224,In_233);
and U1396 (N_1396,In_513,In_673);
nand U1397 (N_1397,In_826,In_1379);
xor U1398 (N_1398,In_258,In_575);
or U1399 (N_1399,In_1205,In_698);
or U1400 (N_1400,In_1388,In_877);
or U1401 (N_1401,In_501,In_1325);
or U1402 (N_1402,In_371,In_645);
or U1403 (N_1403,In_863,In_1075);
nand U1404 (N_1404,In_785,In_914);
xnor U1405 (N_1405,In_544,In_188);
and U1406 (N_1406,In_12,In_1479);
nor U1407 (N_1407,In_814,In_331);
nor U1408 (N_1408,In_901,In_1250);
and U1409 (N_1409,In_1474,In_300);
nor U1410 (N_1410,In_937,In_765);
and U1411 (N_1411,In_950,In_187);
or U1412 (N_1412,In_1355,In_130);
nand U1413 (N_1413,In_712,In_814);
nand U1414 (N_1414,In_1193,In_902);
xor U1415 (N_1415,In_1128,In_838);
or U1416 (N_1416,In_422,In_443);
and U1417 (N_1417,In_494,In_514);
nor U1418 (N_1418,In_768,In_789);
or U1419 (N_1419,In_841,In_794);
nand U1420 (N_1420,In_906,In_240);
or U1421 (N_1421,In_146,In_1112);
nand U1422 (N_1422,In_1095,In_724);
nand U1423 (N_1423,In_771,In_799);
nand U1424 (N_1424,In_1453,In_1296);
and U1425 (N_1425,In_1046,In_1255);
nand U1426 (N_1426,In_982,In_1151);
nor U1427 (N_1427,In_232,In_1245);
or U1428 (N_1428,In_226,In_285);
and U1429 (N_1429,In_1146,In_164);
or U1430 (N_1430,In_276,In_258);
or U1431 (N_1431,In_198,In_725);
xor U1432 (N_1432,In_1077,In_1184);
nand U1433 (N_1433,In_894,In_386);
nand U1434 (N_1434,In_349,In_934);
or U1435 (N_1435,In_1496,In_698);
nor U1436 (N_1436,In_186,In_892);
and U1437 (N_1437,In_1232,In_113);
nand U1438 (N_1438,In_984,In_938);
and U1439 (N_1439,In_379,In_520);
nor U1440 (N_1440,In_1176,In_29);
and U1441 (N_1441,In_1219,In_819);
and U1442 (N_1442,In_723,In_599);
or U1443 (N_1443,In_405,In_1093);
nand U1444 (N_1444,In_1420,In_401);
nand U1445 (N_1445,In_1090,In_296);
or U1446 (N_1446,In_693,In_311);
nor U1447 (N_1447,In_331,In_914);
or U1448 (N_1448,In_929,In_1102);
or U1449 (N_1449,In_166,In_188);
nor U1450 (N_1450,In_1193,In_870);
or U1451 (N_1451,In_1162,In_313);
or U1452 (N_1452,In_2,In_1147);
nand U1453 (N_1453,In_1195,In_493);
and U1454 (N_1454,In_1192,In_161);
nor U1455 (N_1455,In_1451,In_1105);
and U1456 (N_1456,In_1052,In_230);
nand U1457 (N_1457,In_932,In_1093);
and U1458 (N_1458,In_227,In_1283);
nor U1459 (N_1459,In_1196,In_582);
nand U1460 (N_1460,In_120,In_1027);
or U1461 (N_1461,In_51,In_935);
nor U1462 (N_1462,In_1361,In_140);
and U1463 (N_1463,In_1350,In_400);
nor U1464 (N_1464,In_644,In_297);
and U1465 (N_1465,In_914,In_105);
nand U1466 (N_1466,In_1129,In_771);
nand U1467 (N_1467,In_57,In_97);
nor U1468 (N_1468,In_937,In_1237);
and U1469 (N_1469,In_832,In_634);
nor U1470 (N_1470,In_512,In_139);
and U1471 (N_1471,In_375,In_794);
or U1472 (N_1472,In_29,In_0);
nand U1473 (N_1473,In_63,In_1162);
nand U1474 (N_1474,In_831,In_99);
nor U1475 (N_1475,In_212,In_808);
and U1476 (N_1476,In_323,In_1);
nand U1477 (N_1477,In_929,In_62);
and U1478 (N_1478,In_508,In_21);
xor U1479 (N_1479,In_748,In_1406);
nand U1480 (N_1480,In_63,In_58);
xor U1481 (N_1481,In_494,In_844);
or U1482 (N_1482,In_1349,In_262);
nand U1483 (N_1483,In_952,In_1181);
nor U1484 (N_1484,In_679,In_1264);
and U1485 (N_1485,In_483,In_862);
xor U1486 (N_1486,In_1178,In_1008);
and U1487 (N_1487,In_833,In_1263);
and U1488 (N_1488,In_1432,In_534);
and U1489 (N_1489,In_205,In_1100);
nor U1490 (N_1490,In_594,In_1227);
nand U1491 (N_1491,In_8,In_124);
or U1492 (N_1492,In_1274,In_490);
xor U1493 (N_1493,In_532,In_246);
or U1494 (N_1494,In_1026,In_364);
and U1495 (N_1495,In_755,In_609);
nor U1496 (N_1496,In_166,In_995);
xnor U1497 (N_1497,In_1420,In_1185);
or U1498 (N_1498,In_600,In_447);
nand U1499 (N_1499,In_1288,In_697);
nand U1500 (N_1500,In_545,In_152);
and U1501 (N_1501,In_1438,In_666);
and U1502 (N_1502,In_30,In_54);
nand U1503 (N_1503,In_539,In_480);
or U1504 (N_1504,In_52,In_369);
or U1505 (N_1505,In_215,In_618);
and U1506 (N_1506,In_841,In_950);
nand U1507 (N_1507,In_235,In_676);
nor U1508 (N_1508,In_93,In_1322);
and U1509 (N_1509,In_79,In_488);
nand U1510 (N_1510,In_693,In_608);
nor U1511 (N_1511,In_1218,In_1448);
nand U1512 (N_1512,In_167,In_1127);
nand U1513 (N_1513,In_900,In_592);
nor U1514 (N_1514,In_282,In_898);
nand U1515 (N_1515,In_252,In_134);
and U1516 (N_1516,In_537,In_949);
xor U1517 (N_1517,In_355,In_798);
nor U1518 (N_1518,In_714,In_1175);
nor U1519 (N_1519,In_1301,In_650);
or U1520 (N_1520,In_28,In_33);
nand U1521 (N_1521,In_1479,In_289);
nand U1522 (N_1522,In_900,In_298);
nor U1523 (N_1523,In_1340,In_353);
nand U1524 (N_1524,In_738,In_698);
xor U1525 (N_1525,In_758,In_560);
or U1526 (N_1526,In_795,In_504);
and U1527 (N_1527,In_117,In_720);
or U1528 (N_1528,In_376,In_975);
and U1529 (N_1529,In_976,In_752);
or U1530 (N_1530,In_991,In_627);
nor U1531 (N_1531,In_1050,In_81);
or U1532 (N_1532,In_770,In_354);
or U1533 (N_1533,In_480,In_555);
or U1534 (N_1534,In_648,In_1267);
and U1535 (N_1535,In_1180,In_259);
nand U1536 (N_1536,In_747,In_107);
nand U1537 (N_1537,In_152,In_427);
nor U1538 (N_1538,In_1132,In_205);
and U1539 (N_1539,In_848,In_634);
and U1540 (N_1540,In_388,In_116);
and U1541 (N_1541,In_703,In_1293);
xor U1542 (N_1542,In_719,In_272);
nor U1543 (N_1543,In_185,In_1444);
nand U1544 (N_1544,In_502,In_681);
nor U1545 (N_1545,In_1163,In_1296);
and U1546 (N_1546,In_533,In_914);
or U1547 (N_1547,In_55,In_392);
nand U1548 (N_1548,In_767,In_201);
and U1549 (N_1549,In_534,In_144);
nand U1550 (N_1550,In_822,In_246);
or U1551 (N_1551,In_1375,In_1123);
nor U1552 (N_1552,In_414,In_255);
or U1553 (N_1553,In_113,In_28);
nor U1554 (N_1554,In_214,In_1349);
and U1555 (N_1555,In_357,In_442);
and U1556 (N_1556,In_431,In_329);
nand U1557 (N_1557,In_298,In_875);
or U1558 (N_1558,In_772,In_1378);
xor U1559 (N_1559,In_1209,In_485);
and U1560 (N_1560,In_602,In_758);
nor U1561 (N_1561,In_511,In_721);
or U1562 (N_1562,In_620,In_256);
xnor U1563 (N_1563,In_1060,In_809);
nand U1564 (N_1564,In_115,In_1074);
or U1565 (N_1565,In_460,In_697);
or U1566 (N_1566,In_1082,In_838);
and U1567 (N_1567,In_1230,In_1322);
nand U1568 (N_1568,In_1185,In_911);
nor U1569 (N_1569,In_1365,In_63);
nand U1570 (N_1570,In_987,In_671);
or U1571 (N_1571,In_310,In_1402);
nand U1572 (N_1572,In_180,In_760);
nand U1573 (N_1573,In_542,In_851);
nor U1574 (N_1574,In_845,In_191);
and U1575 (N_1575,In_976,In_1210);
or U1576 (N_1576,In_578,In_650);
nand U1577 (N_1577,In_355,In_1247);
or U1578 (N_1578,In_1361,In_1343);
nor U1579 (N_1579,In_833,In_859);
or U1580 (N_1580,In_336,In_1007);
nand U1581 (N_1581,In_1454,In_886);
nor U1582 (N_1582,In_1386,In_696);
or U1583 (N_1583,In_868,In_105);
or U1584 (N_1584,In_1030,In_217);
or U1585 (N_1585,In_1488,In_36);
nor U1586 (N_1586,In_843,In_45);
or U1587 (N_1587,In_283,In_1324);
nand U1588 (N_1588,In_731,In_1265);
and U1589 (N_1589,In_395,In_264);
xnor U1590 (N_1590,In_1333,In_365);
and U1591 (N_1591,In_494,In_937);
and U1592 (N_1592,In_54,In_686);
xnor U1593 (N_1593,In_168,In_298);
xor U1594 (N_1594,In_43,In_439);
and U1595 (N_1595,In_1158,In_51);
or U1596 (N_1596,In_984,In_439);
nor U1597 (N_1597,In_604,In_951);
nor U1598 (N_1598,In_122,In_643);
and U1599 (N_1599,In_442,In_606);
nand U1600 (N_1600,In_368,In_968);
or U1601 (N_1601,In_114,In_232);
nand U1602 (N_1602,In_1294,In_491);
or U1603 (N_1603,In_481,In_1113);
and U1604 (N_1604,In_383,In_1318);
or U1605 (N_1605,In_718,In_204);
nor U1606 (N_1606,In_73,In_378);
or U1607 (N_1607,In_896,In_492);
and U1608 (N_1608,In_1235,In_598);
nor U1609 (N_1609,In_529,In_1301);
nand U1610 (N_1610,In_255,In_860);
or U1611 (N_1611,In_505,In_318);
or U1612 (N_1612,In_54,In_1261);
nor U1613 (N_1613,In_654,In_313);
xor U1614 (N_1614,In_759,In_487);
or U1615 (N_1615,In_583,In_981);
xnor U1616 (N_1616,In_1344,In_799);
xor U1617 (N_1617,In_160,In_388);
nand U1618 (N_1618,In_509,In_693);
xor U1619 (N_1619,In_1010,In_702);
or U1620 (N_1620,In_663,In_1298);
or U1621 (N_1621,In_1136,In_1309);
and U1622 (N_1622,In_1466,In_963);
and U1623 (N_1623,In_808,In_192);
nor U1624 (N_1624,In_611,In_1405);
or U1625 (N_1625,In_190,In_793);
nor U1626 (N_1626,In_927,In_1016);
nor U1627 (N_1627,In_382,In_171);
and U1628 (N_1628,In_1221,In_339);
xor U1629 (N_1629,In_333,In_1271);
nand U1630 (N_1630,In_635,In_1154);
nor U1631 (N_1631,In_1013,In_164);
or U1632 (N_1632,In_652,In_60);
and U1633 (N_1633,In_157,In_584);
nor U1634 (N_1634,In_191,In_895);
nor U1635 (N_1635,In_810,In_425);
nand U1636 (N_1636,In_353,In_549);
and U1637 (N_1637,In_623,In_905);
nor U1638 (N_1638,In_246,In_171);
nor U1639 (N_1639,In_233,In_555);
or U1640 (N_1640,In_1483,In_1188);
or U1641 (N_1641,In_1031,In_1355);
xnor U1642 (N_1642,In_1316,In_943);
and U1643 (N_1643,In_1145,In_250);
xor U1644 (N_1644,In_1353,In_863);
and U1645 (N_1645,In_728,In_1280);
or U1646 (N_1646,In_460,In_583);
nand U1647 (N_1647,In_1256,In_267);
nor U1648 (N_1648,In_1162,In_1029);
and U1649 (N_1649,In_1055,In_538);
nor U1650 (N_1650,In_1467,In_1311);
and U1651 (N_1651,In_974,In_1074);
or U1652 (N_1652,In_1499,In_159);
nor U1653 (N_1653,In_1026,In_898);
nand U1654 (N_1654,In_1236,In_823);
and U1655 (N_1655,In_1198,In_1341);
and U1656 (N_1656,In_1443,In_1001);
and U1657 (N_1657,In_1351,In_623);
and U1658 (N_1658,In_662,In_1216);
xnor U1659 (N_1659,In_116,In_935);
xnor U1660 (N_1660,In_111,In_1324);
nor U1661 (N_1661,In_418,In_1466);
nand U1662 (N_1662,In_1433,In_1248);
nand U1663 (N_1663,In_940,In_1028);
or U1664 (N_1664,In_141,In_1055);
or U1665 (N_1665,In_1464,In_450);
or U1666 (N_1666,In_1472,In_44);
or U1667 (N_1667,In_287,In_1033);
nand U1668 (N_1668,In_1254,In_113);
and U1669 (N_1669,In_1017,In_1477);
and U1670 (N_1670,In_1235,In_250);
nor U1671 (N_1671,In_418,In_972);
nor U1672 (N_1672,In_714,In_187);
nor U1673 (N_1673,In_533,In_883);
or U1674 (N_1674,In_1385,In_1473);
and U1675 (N_1675,In_1155,In_1494);
and U1676 (N_1676,In_328,In_1189);
nand U1677 (N_1677,In_876,In_77);
or U1678 (N_1678,In_1375,In_516);
nor U1679 (N_1679,In_428,In_789);
and U1680 (N_1680,In_756,In_1205);
and U1681 (N_1681,In_724,In_1341);
and U1682 (N_1682,In_1095,In_149);
or U1683 (N_1683,In_505,In_712);
nand U1684 (N_1684,In_1433,In_859);
or U1685 (N_1685,In_468,In_1468);
and U1686 (N_1686,In_1497,In_1210);
and U1687 (N_1687,In_898,In_1224);
or U1688 (N_1688,In_675,In_769);
and U1689 (N_1689,In_509,In_1380);
nand U1690 (N_1690,In_985,In_235);
nor U1691 (N_1691,In_789,In_361);
or U1692 (N_1692,In_715,In_1030);
nor U1693 (N_1693,In_908,In_922);
nor U1694 (N_1694,In_216,In_377);
and U1695 (N_1695,In_928,In_946);
nor U1696 (N_1696,In_820,In_1417);
and U1697 (N_1697,In_733,In_850);
and U1698 (N_1698,In_1047,In_925);
or U1699 (N_1699,In_963,In_576);
nand U1700 (N_1700,In_1038,In_130);
nor U1701 (N_1701,In_536,In_1342);
and U1702 (N_1702,In_125,In_67);
nor U1703 (N_1703,In_1374,In_536);
or U1704 (N_1704,In_1256,In_1021);
nand U1705 (N_1705,In_666,In_3);
nand U1706 (N_1706,In_95,In_606);
nand U1707 (N_1707,In_61,In_416);
nand U1708 (N_1708,In_189,In_512);
or U1709 (N_1709,In_537,In_1088);
nand U1710 (N_1710,In_1232,In_1277);
nor U1711 (N_1711,In_587,In_503);
or U1712 (N_1712,In_1459,In_829);
and U1713 (N_1713,In_1011,In_700);
nand U1714 (N_1714,In_1252,In_768);
nor U1715 (N_1715,In_1165,In_912);
nor U1716 (N_1716,In_523,In_604);
and U1717 (N_1717,In_535,In_382);
or U1718 (N_1718,In_712,In_659);
and U1719 (N_1719,In_1343,In_761);
nand U1720 (N_1720,In_1121,In_211);
or U1721 (N_1721,In_511,In_1165);
or U1722 (N_1722,In_578,In_171);
and U1723 (N_1723,In_536,In_1012);
or U1724 (N_1724,In_32,In_710);
or U1725 (N_1725,In_1427,In_582);
or U1726 (N_1726,In_1139,In_1186);
nor U1727 (N_1727,In_1227,In_255);
xor U1728 (N_1728,In_106,In_14);
or U1729 (N_1729,In_1281,In_591);
and U1730 (N_1730,In_733,In_1384);
and U1731 (N_1731,In_674,In_1171);
and U1732 (N_1732,In_971,In_1206);
xnor U1733 (N_1733,In_1403,In_1074);
or U1734 (N_1734,In_1388,In_984);
or U1735 (N_1735,In_1279,In_59);
or U1736 (N_1736,In_125,In_943);
or U1737 (N_1737,In_1197,In_1216);
nor U1738 (N_1738,In_781,In_1358);
nor U1739 (N_1739,In_700,In_779);
or U1740 (N_1740,In_1071,In_338);
and U1741 (N_1741,In_1154,In_175);
and U1742 (N_1742,In_1087,In_771);
and U1743 (N_1743,In_1134,In_1151);
nor U1744 (N_1744,In_592,In_868);
or U1745 (N_1745,In_183,In_375);
xor U1746 (N_1746,In_956,In_321);
nor U1747 (N_1747,In_70,In_375);
or U1748 (N_1748,In_1237,In_255);
or U1749 (N_1749,In_613,In_902);
xor U1750 (N_1750,In_1244,In_8);
or U1751 (N_1751,In_68,In_542);
or U1752 (N_1752,In_1107,In_880);
xor U1753 (N_1753,In_49,In_423);
and U1754 (N_1754,In_875,In_1444);
nand U1755 (N_1755,In_507,In_1105);
nor U1756 (N_1756,In_712,In_809);
nor U1757 (N_1757,In_1196,In_739);
or U1758 (N_1758,In_935,In_1120);
nand U1759 (N_1759,In_284,In_135);
and U1760 (N_1760,In_723,In_27);
xor U1761 (N_1761,In_671,In_124);
or U1762 (N_1762,In_1109,In_178);
nand U1763 (N_1763,In_268,In_779);
nand U1764 (N_1764,In_674,In_1080);
or U1765 (N_1765,In_120,In_225);
nand U1766 (N_1766,In_1001,In_842);
nor U1767 (N_1767,In_1034,In_1240);
and U1768 (N_1768,In_270,In_1283);
and U1769 (N_1769,In_1348,In_1483);
and U1770 (N_1770,In_958,In_281);
or U1771 (N_1771,In_385,In_560);
xnor U1772 (N_1772,In_1168,In_1420);
or U1773 (N_1773,In_1267,In_559);
nor U1774 (N_1774,In_333,In_427);
nand U1775 (N_1775,In_845,In_1456);
nand U1776 (N_1776,In_1274,In_128);
or U1777 (N_1777,In_630,In_1211);
xor U1778 (N_1778,In_393,In_987);
nor U1779 (N_1779,In_238,In_650);
or U1780 (N_1780,In_926,In_958);
and U1781 (N_1781,In_504,In_1019);
xnor U1782 (N_1782,In_898,In_1202);
and U1783 (N_1783,In_1449,In_99);
nand U1784 (N_1784,In_1119,In_1418);
nor U1785 (N_1785,In_1027,In_1377);
nand U1786 (N_1786,In_201,In_1449);
nand U1787 (N_1787,In_998,In_1066);
or U1788 (N_1788,In_94,In_1488);
nor U1789 (N_1789,In_592,In_1246);
nand U1790 (N_1790,In_1444,In_284);
nor U1791 (N_1791,In_1134,In_549);
or U1792 (N_1792,In_25,In_283);
or U1793 (N_1793,In_954,In_810);
nand U1794 (N_1794,In_826,In_734);
nand U1795 (N_1795,In_344,In_660);
xor U1796 (N_1796,In_828,In_480);
and U1797 (N_1797,In_1341,In_892);
nand U1798 (N_1798,In_1381,In_1123);
xor U1799 (N_1799,In_741,In_1140);
nor U1800 (N_1800,In_1173,In_1039);
nor U1801 (N_1801,In_1237,In_403);
or U1802 (N_1802,In_627,In_980);
nand U1803 (N_1803,In_1069,In_586);
or U1804 (N_1804,In_487,In_777);
nor U1805 (N_1805,In_1011,In_98);
nor U1806 (N_1806,In_1297,In_1051);
nand U1807 (N_1807,In_1285,In_48);
or U1808 (N_1808,In_1084,In_1166);
and U1809 (N_1809,In_675,In_1070);
and U1810 (N_1810,In_1394,In_229);
and U1811 (N_1811,In_282,In_1045);
nor U1812 (N_1812,In_380,In_1246);
nor U1813 (N_1813,In_181,In_113);
nand U1814 (N_1814,In_895,In_832);
or U1815 (N_1815,In_832,In_293);
nand U1816 (N_1816,In_241,In_732);
or U1817 (N_1817,In_1171,In_1125);
nand U1818 (N_1818,In_900,In_1430);
nor U1819 (N_1819,In_600,In_521);
nand U1820 (N_1820,In_603,In_943);
nor U1821 (N_1821,In_417,In_495);
nor U1822 (N_1822,In_1053,In_1010);
or U1823 (N_1823,In_690,In_1466);
or U1824 (N_1824,In_359,In_336);
and U1825 (N_1825,In_1396,In_31);
xnor U1826 (N_1826,In_572,In_1378);
nand U1827 (N_1827,In_352,In_507);
nand U1828 (N_1828,In_671,In_933);
and U1829 (N_1829,In_1278,In_365);
nor U1830 (N_1830,In_66,In_157);
xnor U1831 (N_1831,In_988,In_130);
and U1832 (N_1832,In_1257,In_683);
or U1833 (N_1833,In_441,In_1027);
nor U1834 (N_1834,In_48,In_37);
or U1835 (N_1835,In_165,In_263);
and U1836 (N_1836,In_350,In_981);
and U1837 (N_1837,In_847,In_274);
or U1838 (N_1838,In_946,In_151);
or U1839 (N_1839,In_689,In_247);
or U1840 (N_1840,In_2,In_1149);
or U1841 (N_1841,In_231,In_292);
nand U1842 (N_1842,In_1416,In_1418);
or U1843 (N_1843,In_156,In_929);
and U1844 (N_1844,In_635,In_940);
nor U1845 (N_1845,In_593,In_379);
or U1846 (N_1846,In_1461,In_375);
nor U1847 (N_1847,In_854,In_382);
nor U1848 (N_1848,In_50,In_389);
xor U1849 (N_1849,In_1297,In_1227);
xnor U1850 (N_1850,In_95,In_1060);
xnor U1851 (N_1851,In_92,In_268);
nor U1852 (N_1852,In_1217,In_1182);
nor U1853 (N_1853,In_970,In_1074);
or U1854 (N_1854,In_1414,In_306);
or U1855 (N_1855,In_642,In_94);
and U1856 (N_1856,In_630,In_908);
nand U1857 (N_1857,In_1490,In_1376);
and U1858 (N_1858,In_398,In_1239);
nand U1859 (N_1859,In_331,In_283);
nand U1860 (N_1860,In_997,In_913);
or U1861 (N_1861,In_302,In_1402);
nand U1862 (N_1862,In_894,In_1090);
and U1863 (N_1863,In_954,In_1372);
nand U1864 (N_1864,In_88,In_440);
or U1865 (N_1865,In_876,In_1127);
nor U1866 (N_1866,In_915,In_1323);
or U1867 (N_1867,In_20,In_190);
and U1868 (N_1868,In_146,In_368);
nor U1869 (N_1869,In_928,In_1175);
nor U1870 (N_1870,In_633,In_17);
or U1871 (N_1871,In_923,In_173);
or U1872 (N_1872,In_145,In_899);
or U1873 (N_1873,In_1277,In_1005);
or U1874 (N_1874,In_258,In_890);
and U1875 (N_1875,In_1129,In_582);
nand U1876 (N_1876,In_297,In_45);
or U1877 (N_1877,In_840,In_446);
xor U1878 (N_1878,In_367,In_648);
or U1879 (N_1879,In_1274,In_19);
nand U1880 (N_1880,In_353,In_1370);
xor U1881 (N_1881,In_636,In_1333);
or U1882 (N_1882,In_750,In_819);
nor U1883 (N_1883,In_204,In_792);
and U1884 (N_1884,In_1011,In_153);
and U1885 (N_1885,In_1356,In_1192);
or U1886 (N_1886,In_355,In_1160);
nand U1887 (N_1887,In_775,In_432);
or U1888 (N_1888,In_790,In_578);
and U1889 (N_1889,In_16,In_1462);
nand U1890 (N_1890,In_720,In_151);
and U1891 (N_1891,In_424,In_676);
xnor U1892 (N_1892,In_238,In_787);
or U1893 (N_1893,In_1192,In_982);
and U1894 (N_1894,In_933,In_966);
or U1895 (N_1895,In_814,In_782);
nor U1896 (N_1896,In_986,In_139);
and U1897 (N_1897,In_116,In_478);
nor U1898 (N_1898,In_461,In_377);
nor U1899 (N_1899,In_1203,In_699);
nor U1900 (N_1900,In_1046,In_1365);
and U1901 (N_1901,In_218,In_1158);
nor U1902 (N_1902,In_41,In_1341);
xor U1903 (N_1903,In_630,In_681);
nand U1904 (N_1904,In_481,In_1340);
xor U1905 (N_1905,In_396,In_829);
nor U1906 (N_1906,In_804,In_591);
and U1907 (N_1907,In_834,In_978);
or U1908 (N_1908,In_536,In_418);
nor U1909 (N_1909,In_1071,In_1014);
or U1910 (N_1910,In_1096,In_155);
or U1911 (N_1911,In_1059,In_928);
xnor U1912 (N_1912,In_1157,In_1229);
xnor U1913 (N_1913,In_1131,In_641);
xnor U1914 (N_1914,In_218,In_21);
or U1915 (N_1915,In_1191,In_644);
xor U1916 (N_1916,In_82,In_850);
or U1917 (N_1917,In_87,In_733);
nand U1918 (N_1918,In_810,In_1090);
nor U1919 (N_1919,In_61,In_457);
and U1920 (N_1920,In_327,In_649);
nand U1921 (N_1921,In_863,In_868);
and U1922 (N_1922,In_1133,In_1318);
and U1923 (N_1923,In_1263,In_495);
or U1924 (N_1924,In_435,In_1288);
or U1925 (N_1925,In_452,In_941);
nor U1926 (N_1926,In_949,In_448);
nor U1927 (N_1927,In_1485,In_281);
or U1928 (N_1928,In_348,In_801);
nor U1929 (N_1929,In_111,In_1366);
nand U1930 (N_1930,In_772,In_623);
nor U1931 (N_1931,In_1359,In_1252);
nand U1932 (N_1932,In_726,In_677);
nor U1933 (N_1933,In_1329,In_749);
xnor U1934 (N_1934,In_105,In_1234);
nand U1935 (N_1935,In_454,In_456);
nor U1936 (N_1936,In_1375,In_933);
xor U1937 (N_1937,In_1087,In_1479);
or U1938 (N_1938,In_988,In_1379);
and U1939 (N_1939,In_295,In_1402);
or U1940 (N_1940,In_1199,In_1478);
and U1941 (N_1941,In_758,In_179);
nor U1942 (N_1942,In_1381,In_169);
and U1943 (N_1943,In_833,In_507);
nor U1944 (N_1944,In_551,In_1351);
nor U1945 (N_1945,In_606,In_663);
xor U1946 (N_1946,In_1433,In_116);
or U1947 (N_1947,In_1126,In_177);
nor U1948 (N_1948,In_457,In_1442);
and U1949 (N_1949,In_145,In_505);
and U1950 (N_1950,In_981,In_878);
and U1951 (N_1951,In_421,In_1391);
or U1952 (N_1952,In_1176,In_445);
and U1953 (N_1953,In_1482,In_396);
nand U1954 (N_1954,In_365,In_791);
xor U1955 (N_1955,In_1277,In_1359);
xor U1956 (N_1956,In_497,In_434);
xor U1957 (N_1957,In_1354,In_1100);
xor U1958 (N_1958,In_1210,In_260);
nand U1959 (N_1959,In_215,In_1460);
nor U1960 (N_1960,In_824,In_116);
or U1961 (N_1961,In_448,In_998);
nor U1962 (N_1962,In_903,In_27);
or U1963 (N_1963,In_1222,In_619);
and U1964 (N_1964,In_10,In_190);
and U1965 (N_1965,In_862,In_1166);
nor U1966 (N_1966,In_1235,In_1118);
and U1967 (N_1967,In_1213,In_510);
or U1968 (N_1968,In_44,In_271);
and U1969 (N_1969,In_385,In_107);
or U1970 (N_1970,In_722,In_973);
and U1971 (N_1971,In_564,In_1212);
and U1972 (N_1972,In_688,In_1164);
xnor U1973 (N_1973,In_308,In_561);
nor U1974 (N_1974,In_1248,In_1128);
and U1975 (N_1975,In_603,In_1147);
and U1976 (N_1976,In_284,In_1142);
nand U1977 (N_1977,In_615,In_172);
nor U1978 (N_1978,In_489,In_1149);
and U1979 (N_1979,In_1434,In_150);
nand U1980 (N_1980,In_133,In_887);
nor U1981 (N_1981,In_1383,In_1462);
nor U1982 (N_1982,In_563,In_1490);
xor U1983 (N_1983,In_888,In_467);
nand U1984 (N_1984,In_508,In_986);
nor U1985 (N_1985,In_740,In_1378);
or U1986 (N_1986,In_189,In_836);
or U1987 (N_1987,In_842,In_743);
and U1988 (N_1988,In_667,In_274);
and U1989 (N_1989,In_1357,In_15);
nor U1990 (N_1990,In_550,In_626);
nor U1991 (N_1991,In_1254,In_1338);
xnor U1992 (N_1992,In_608,In_621);
or U1993 (N_1993,In_1280,In_1480);
or U1994 (N_1994,In_602,In_202);
or U1995 (N_1995,In_156,In_1382);
nand U1996 (N_1996,In_780,In_377);
nor U1997 (N_1997,In_602,In_270);
or U1998 (N_1998,In_753,In_764);
or U1999 (N_1999,In_238,In_245);
nand U2000 (N_2000,In_1175,In_133);
or U2001 (N_2001,In_667,In_621);
xor U2002 (N_2002,In_328,In_801);
or U2003 (N_2003,In_49,In_665);
or U2004 (N_2004,In_1030,In_30);
or U2005 (N_2005,In_866,In_598);
and U2006 (N_2006,In_1328,In_414);
and U2007 (N_2007,In_9,In_559);
and U2008 (N_2008,In_769,In_231);
or U2009 (N_2009,In_438,In_598);
or U2010 (N_2010,In_1282,In_1457);
and U2011 (N_2011,In_1185,In_380);
nor U2012 (N_2012,In_187,In_987);
or U2013 (N_2013,In_938,In_703);
nor U2014 (N_2014,In_1082,In_212);
nor U2015 (N_2015,In_1053,In_813);
nand U2016 (N_2016,In_368,In_829);
or U2017 (N_2017,In_407,In_612);
nand U2018 (N_2018,In_774,In_222);
xor U2019 (N_2019,In_1258,In_365);
xnor U2020 (N_2020,In_1216,In_758);
nor U2021 (N_2021,In_783,In_618);
or U2022 (N_2022,In_1395,In_265);
and U2023 (N_2023,In_393,In_968);
xnor U2024 (N_2024,In_53,In_1114);
nand U2025 (N_2025,In_1392,In_1369);
nand U2026 (N_2026,In_736,In_902);
nand U2027 (N_2027,In_107,In_847);
nor U2028 (N_2028,In_1119,In_1000);
or U2029 (N_2029,In_1091,In_522);
or U2030 (N_2030,In_185,In_873);
and U2031 (N_2031,In_1255,In_31);
nor U2032 (N_2032,In_65,In_797);
nor U2033 (N_2033,In_532,In_724);
nor U2034 (N_2034,In_1147,In_117);
nand U2035 (N_2035,In_1166,In_793);
nor U2036 (N_2036,In_600,In_67);
xnor U2037 (N_2037,In_401,In_680);
xor U2038 (N_2038,In_143,In_1448);
xnor U2039 (N_2039,In_885,In_1215);
nor U2040 (N_2040,In_1497,In_455);
xor U2041 (N_2041,In_200,In_1229);
nor U2042 (N_2042,In_587,In_879);
nor U2043 (N_2043,In_178,In_1130);
nand U2044 (N_2044,In_563,In_324);
nand U2045 (N_2045,In_1059,In_822);
nor U2046 (N_2046,In_1004,In_776);
and U2047 (N_2047,In_1192,In_205);
nor U2048 (N_2048,In_1125,In_179);
nand U2049 (N_2049,In_916,In_557);
nand U2050 (N_2050,In_957,In_214);
nor U2051 (N_2051,In_160,In_1294);
and U2052 (N_2052,In_581,In_382);
xnor U2053 (N_2053,In_1362,In_436);
and U2054 (N_2054,In_1381,In_268);
and U2055 (N_2055,In_1227,In_568);
xor U2056 (N_2056,In_1244,In_891);
nand U2057 (N_2057,In_41,In_820);
nand U2058 (N_2058,In_327,In_49);
and U2059 (N_2059,In_578,In_320);
nor U2060 (N_2060,In_530,In_1174);
nor U2061 (N_2061,In_1004,In_392);
and U2062 (N_2062,In_509,In_708);
nand U2063 (N_2063,In_131,In_180);
nand U2064 (N_2064,In_994,In_619);
nor U2065 (N_2065,In_998,In_536);
nand U2066 (N_2066,In_1455,In_661);
nand U2067 (N_2067,In_1197,In_1267);
or U2068 (N_2068,In_304,In_339);
nor U2069 (N_2069,In_174,In_4);
or U2070 (N_2070,In_379,In_993);
xor U2071 (N_2071,In_126,In_489);
and U2072 (N_2072,In_1429,In_1333);
and U2073 (N_2073,In_753,In_981);
nand U2074 (N_2074,In_673,In_1136);
or U2075 (N_2075,In_1490,In_1036);
xnor U2076 (N_2076,In_1297,In_1225);
nor U2077 (N_2077,In_695,In_1135);
or U2078 (N_2078,In_1300,In_647);
nor U2079 (N_2079,In_1317,In_102);
or U2080 (N_2080,In_1386,In_167);
or U2081 (N_2081,In_532,In_278);
nand U2082 (N_2082,In_37,In_1123);
and U2083 (N_2083,In_28,In_1047);
and U2084 (N_2084,In_696,In_1264);
or U2085 (N_2085,In_1100,In_1219);
and U2086 (N_2086,In_1080,In_146);
nand U2087 (N_2087,In_1417,In_234);
or U2088 (N_2088,In_356,In_629);
nor U2089 (N_2089,In_192,In_340);
nor U2090 (N_2090,In_1238,In_1460);
and U2091 (N_2091,In_1336,In_285);
and U2092 (N_2092,In_184,In_175);
nand U2093 (N_2093,In_459,In_1088);
nand U2094 (N_2094,In_36,In_1052);
nand U2095 (N_2095,In_134,In_876);
and U2096 (N_2096,In_929,In_608);
or U2097 (N_2097,In_1446,In_759);
xor U2098 (N_2098,In_257,In_19);
nor U2099 (N_2099,In_454,In_412);
nor U2100 (N_2100,In_1281,In_514);
and U2101 (N_2101,In_1499,In_37);
and U2102 (N_2102,In_91,In_793);
or U2103 (N_2103,In_8,In_1283);
and U2104 (N_2104,In_668,In_308);
or U2105 (N_2105,In_354,In_1320);
nand U2106 (N_2106,In_415,In_646);
or U2107 (N_2107,In_156,In_738);
and U2108 (N_2108,In_385,In_1425);
nand U2109 (N_2109,In_366,In_988);
nand U2110 (N_2110,In_1479,In_749);
nand U2111 (N_2111,In_188,In_86);
and U2112 (N_2112,In_459,In_1356);
nor U2113 (N_2113,In_1084,In_507);
nor U2114 (N_2114,In_1230,In_1212);
nand U2115 (N_2115,In_242,In_647);
or U2116 (N_2116,In_348,In_999);
and U2117 (N_2117,In_941,In_1157);
xor U2118 (N_2118,In_892,In_69);
and U2119 (N_2119,In_378,In_1368);
or U2120 (N_2120,In_244,In_1126);
nand U2121 (N_2121,In_521,In_1392);
nand U2122 (N_2122,In_1213,In_174);
and U2123 (N_2123,In_823,In_1209);
and U2124 (N_2124,In_90,In_625);
nand U2125 (N_2125,In_158,In_1462);
nor U2126 (N_2126,In_1440,In_1401);
or U2127 (N_2127,In_715,In_1213);
xnor U2128 (N_2128,In_1358,In_1097);
or U2129 (N_2129,In_1169,In_180);
and U2130 (N_2130,In_1010,In_1127);
or U2131 (N_2131,In_469,In_1242);
xor U2132 (N_2132,In_1002,In_948);
nor U2133 (N_2133,In_456,In_429);
and U2134 (N_2134,In_309,In_301);
or U2135 (N_2135,In_20,In_137);
or U2136 (N_2136,In_1397,In_520);
and U2137 (N_2137,In_1223,In_351);
or U2138 (N_2138,In_438,In_832);
nand U2139 (N_2139,In_1351,In_932);
or U2140 (N_2140,In_323,In_404);
and U2141 (N_2141,In_5,In_564);
nand U2142 (N_2142,In_736,In_320);
nor U2143 (N_2143,In_1393,In_1198);
nand U2144 (N_2144,In_554,In_723);
nand U2145 (N_2145,In_819,In_1297);
nor U2146 (N_2146,In_715,In_918);
nor U2147 (N_2147,In_887,In_588);
and U2148 (N_2148,In_224,In_664);
or U2149 (N_2149,In_660,In_609);
and U2150 (N_2150,In_1214,In_271);
and U2151 (N_2151,In_561,In_321);
xor U2152 (N_2152,In_184,In_317);
nor U2153 (N_2153,In_982,In_289);
nand U2154 (N_2154,In_876,In_24);
or U2155 (N_2155,In_265,In_360);
and U2156 (N_2156,In_426,In_834);
and U2157 (N_2157,In_690,In_14);
nor U2158 (N_2158,In_506,In_696);
nand U2159 (N_2159,In_989,In_990);
xor U2160 (N_2160,In_1356,In_258);
and U2161 (N_2161,In_582,In_1200);
nand U2162 (N_2162,In_987,In_579);
nor U2163 (N_2163,In_1473,In_353);
xor U2164 (N_2164,In_795,In_631);
and U2165 (N_2165,In_800,In_45);
nand U2166 (N_2166,In_995,In_794);
or U2167 (N_2167,In_966,In_293);
nand U2168 (N_2168,In_1433,In_1330);
or U2169 (N_2169,In_1122,In_602);
or U2170 (N_2170,In_703,In_595);
xor U2171 (N_2171,In_748,In_1252);
xor U2172 (N_2172,In_900,In_407);
or U2173 (N_2173,In_1080,In_652);
xnor U2174 (N_2174,In_831,In_740);
and U2175 (N_2175,In_1238,In_742);
nand U2176 (N_2176,In_859,In_1194);
nand U2177 (N_2177,In_670,In_456);
or U2178 (N_2178,In_199,In_1024);
or U2179 (N_2179,In_153,In_886);
or U2180 (N_2180,In_1153,In_84);
xor U2181 (N_2181,In_639,In_855);
and U2182 (N_2182,In_1172,In_837);
and U2183 (N_2183,In_270,In_285);
nand U2184 (N_2184,In_1011,In_694);
and U2185 (N_2185,In_1473,In_300);
or U2186 (N_2186,In_1092,In_458);
xor U2187 (N_2187,In_308,In_484);
and U2188 (N_2188,In_627,In_741);
nand U2189 (N_2189,In_1064,In_737);
nor U2190 (N_2190,In_133,In_730);
and U2191 (N_2191,In_26,In_340);
nand U2192 (N_2192,In_561,In_486);
and U2193 (N_2193,In_1337,In_349);
and U2194 (N_2194,In_249,In_1474);
nand U2195 (N_2195,In_652,In_364);
and U2196 (N_2196,In_698,In_500);
nand U2197 (N_2197,In_588,In_822);
nand U2198 (N_2198,In_1446,In_1465);
nor U2199 (N_2199,In_96,In_576);
and U2200 (N_2200,In_978,In_1272);
or U2201 (N_2201,In_1015,In_844);
nand U2202 (N_2202,In_617,In_1022);
or U2203 (N_2203,In_966,In_460);
or U2204 (N_2204,In_495,In_1221);
nor U2205 (N_2205,In_294,In_685);
nor U2206 (N_2206,In_429,In_762);
and U2207 (N_2207,In_1368,In_1456);
nor U2208 (N_2208,In_682,In_769);
nor U2209 (N_2209,In_972,In_407);
and U2210 (N_2210,In_1351,In_1074);
nor U2211 (N_2211,In_314,In_726);
and U2212 (N_2212,In_633,In_1118);
or U2213 (N_2213,In_1424,In_46);
nand U2214 (N_2214,In_101,In_678);
nor U2215 (N_2215,In_169,In_1171);
or U2216 (N_2216,In_72,In_887);
and U2217 (N_2217,In_155,In_593);
and U2218 (N_2218,In_318,In_75);
and U2219 (N_2219,In_92,In_1232);
or U2220 (N_2220,In_1280,In_800);
and U2221 (N_2221,In_819,In_508);
or U2222 (N_2222,In_139,In_1394);
xnor U2223 (N_2223,In_1387,In_1288);
and U2224 (N_2224,In_734,In_740);
and U2225 (N_2225,In_1075,In_954);
and U2226 (N_2226,In_191,In_92);
or U2227 (N_2227,In_555,In_450);
nor U2228 (N_2228,In_366,In_979);
and U2229 (N_2229,In_124,In_714);
nor U2230 (N_2230,In_1098,In_1343);
nand U2231 (N_2231,In_442,In_174);
and U2232 (N_2232,In_167,In_325);
nand U2233 (N_2233,In_1064,In_700);
nor U2234 (N_2234,In_171,In_489);
and U2235 (N_2235,In_1137,In_366);
nor U2236 (N_2236,In_307,In_512);
xor U2237 (N_2237,In_603,In_78);
or U2238 (N_2238,In_598,In_159);
or U2239 (N_2239,In_275,In_554);
or U2240 (N_2240,In_1239,In_1355);
nand U2241 (N_2241,In_114,In_481);
xor U2242 (N_2242,In_458,In_901);
nand U2243 (N_2243,In_1417,In_1362);
and U2244 (N_2244,In_138,In_19);
and U2245 (N_2245,In_1101,In_836);
nand U2246 (N_2246,In_519,In_1436);
and U2247 (N_2247,In_1358,In_670);
or U2248 (N_2248,In_627,In_463);
xor U2249 (N_2249,In_1374,In_772);
and U2250 (N_2250,In_857,In_757);
or U2251 (N_2251,In_661,In_796);
nor U2252 (N_2252,In_930,In_564);
and U2253 (N_2253,In_835,In_645);
nor U2254 (N_2254,In_426,In_660);
or U2255 (N_2255,In_553,In_1127);
nor U2256 (N_2256,In_203,In_1488);
and U2257 (N_2257,In_644,In_838);
or U2258 (N_2258,In_179,In_874);
nand U2259 (N_2259,In_400,In_202);
or U2260 (N_2260,In_371,In_432);
nor U2261 (N_2261,In_1209,In_1404);
or U2262 (N_2262,In_774,In_63);
or U2263 (N_2263,In_938,In_386);
and U2264 (N_2264,In_506,In_997);
nor U2265 (N_2265,In_668,In_1247);
nand U2266 (N_2266,In_305,In_230);
xnor U2267 (N_2267,In_791,In_1216);
and U2268 (N_2268,In_39,In_1480);
and U2269 (N_2269,In_14,In_192);
xor U2270 (N_2270,In_1000,In_1002);
nand U2271 (N_2271,In_1102,In_115);
nand U2272 (N_2272,In_721,In_936);
nor U2273 (N_2273,In_1300,In_1133);
and U2274 (N_2274,In_416,In_1180);
nor U2275 (N_2275,In_308,In_418);
or U2276 (N_2276,In_1206,In_727);
nand U2277 (N_2277,In_1480,In_980);
nand U2278 (N_2278,In_154,In_1167);
or U2279 (N_2279,In_313,In_199);
nand U2280 (N_2280,In_261,In_355);
and U2281 (N_2281,In_603,In_1247);
nand U2282 (N_2282,In_689,In_883);
or U2283 (N_2283,In_422,In_713);
and U2284 (N_2284,In_845,In_781);
or U2285 (N_2285,In_880,In_710);
and U2286 (N_2286,In_915,In_191);
nor U2287 (N_2287,In_983,In_41);
and U2288 (N_2288,In_461,In_561);
nand U2289 (N_2289,In_1019,In_1200);
nor U2290 (N_2290,In_478,In_785);
nor U2291 (N_2291,In_270,In_547);
nand U2292 (N_2292,In_191,In_1355);
or U2293 (N_2293,In_488,In_170);
nor U2294 (N_2294,In_725,In_568);
nor U2295 (N_2295,In_672,In_289);
nor U2296 (N_2296,In_440,In_66);
or U2297 (N_2297,In_721,In_1218);
nand U2298 (N_2298,In_25,In_274);
or U2299 (N_2299,In_756,In_773);
and U2300 (N_2300,In_1397,In_1481);
nor U2301 (N_2301,In_13,In_369);
and U2302 (N_2302,In_1385,In_764);
nand U2303 (N_2303,In_1148,In_67);
and U2304 (N_2304,In_951,In_844);
or U2305 (N_2305,In_613,In_166);
or U2306 (N_2306,In_143,In_17);
nand U2307 (N_2307,In_489,In_1355);
nand U2308 (N_2308,In_1150,In_398);
or U2309 (N_2309,In_1081,In_766);
nand U2310 (N_2310,In_1027,In_957);
nor U2311 (N_2311,In_214,In_243);
and U2312 (N_2312,In_1212,In_1214);
and U2313 (N_2313,In_850,In_800);
nand U2314 (N_2314,In_893,In_526);
nand U2315 (N_2315,In_434,In_1020);
nand U2316 (N_2316,In_1191,In_307);
and U2317 (N_2317,In_1081,In_820);
nand U2318 (N_2318,In_595,In_165);
nor U2319 (N_2319,In_320,In_1375);
and U2320 (N_2320,In_370,In_572);
xor U2321 (N_2321,In_1007,In_1166);
xnor U2322 (N_2322,In_601,In_501);
and U2323 (N_2323,In_798,In_787);
xnor U2324 (N_2324,In_606,In_1117);
or U2325 (N_2325,In_681,In_792);
or U2326 (N_2326,In_747,In_482);
and U2327 (N_2327,In_419,In_181);
xnor U2328 (N_2328,In_726,In_920);
and U2329 (N_2329,In_1048,In_699);
or U2330 (N_2330,In_1179,In_617);
and U2331 (N_2331,In_465,In_541);
nand U2332 (N_2332,In_88,In_1308);
and U2333 (N_2333,In_548,In_390);
xnor U2334 (N_2334,In_1021,In_262);
nor U2335 (N_2335,In_621,In_744);
and U2336 (N_2336,In_1112,In_840);
nand U2337 (N_2337,In_351,In_1285);
nand U2338 (N_2338,In_871,In_1161);
nand U2339 (N_2339,In_509,In_193);
or U2340 (N_2340,In_217,In_1058);
or U2341 (N_2341,In_195,In_543);
nor U2342 (N_2342,In_921,In_738);
nor U2343 (N_2343,In_1207,In_1257);
or U2344 (N_2344,In_190,In_664);
and U2345 (N_2345,In_480,In_81);
nand U2346 (N_2346,In_594,In_1354);
or U2347 (N_2347,In_550,In_1479);
or U2348 (N_2348,In_1422,In_548);
nand U2349 (N_2349,In_817,In_1199);
nand U2350 (N_2350,In_1457,In_114);
or U2351 (N_2351,In_772,In_1022);
nor U2352 (N_2352,In_1215,In_1374);
or U2353 (N_2353,In_85,In_1130);
and U2354 (N_2354,In_559,In_337);
nor U2355 (N_2355,In_1475,In_1330);
nor U2356 (N_2356,In_703,In_1319);
nand U2357 (N_2357,In_1223,In_544);
and U2358 (N_2358,In_217,In_892);
and U2359 (N_2359,In_1414,In_8);
or U2360 (N_2360,In_541,In_380);
or U2361 (N_2361,In_569,In_557);
or U2362 (N_2362,In_107,In_1264);
nor U2363 (N_2363,In_751,In_453);
xor U2364 (N_2364,In_528,In_202);
nor U2365 (N_2365,In_1094,In_149);
nor U2366 (N_2366,In_703,In_1060);
xor U2367 (N_2367,In_231,In_766);
or U2368 (N_2368,In_25,In_648);
xor U2369 (N_2369,In_234,In_767);
or U2370 (N_2370,In_366,In_1419);
nand U2371 (N_2371,In_183,In_1030);
nand U2372 (N_2372,In_729,In_984);
nor U2373 (N_2373,In_691,In_1197);
or U2374 (N_2374,In_5,In_1384);
nand U2375 (N_2375,In_1386,In_83);
nand U2376 (N_2376,In_1012,In_1072);
nand U2377 (N_2377,In_399,In_476);
nor U2378 (N_2378,In_1051,In_540);
and U2379 (N_2379,In_740,In_960);
and U2380 (N_2380,In_791,In_431);
nor U2381 (N_2381,In_272,In_196);
xnor U2382 (N_2382,In_256,In_698);
nand U2383 (N_2383,In_13,In_977);
or U2384 (N_2384,In_422,In_1444);
or U2385 (N_2385,In_1279,In_1103);
nor U2386 (N_2386,In_1332,In_1079);
nor U2387 (N_2387,In_481,In_358);
and U2388 (N_2388,In_1300,In_21);
or U2389 (N_2389,In_1208,In_943);
xnor U2390 (N_2390,In_884,In_36);
nor U2391 (N_2391,In_784,In_498);
nor U2392 (N_2392,In_267,In_1383);
and U2393 (N_2393,In_627,In_1291);
nand U2394 (N_2394,In_1360,In_297);
or U2395 (N_2395,In_1183,In_923);
xnor U2396 (N_2396,In_759,In_651);
nor U2397 (N_2397,In_83,In_583);
xor U2398 (N_2398,In_1207,In_1049);
and U2399 (N_2399,In_950,In_514);
and U2400 (N_2400,In_430,In_1118);
and U2401 (N_2401,In_1014,In_3);
and U2402 (N_2402,In_643,In_235);
nor U2403 (N_2403,In_142,In_1374);
nor U2404 (N_2404,In_1152,In_864);
or U2405 (N_2405,In_1430,In_297);
nand U2406 (N_2406,In_332,In_119);
and U2407 (N_2407,In_1217,In_814);
or U2408 (N_2408,In_299,In_801);
or U2409 (N_2409,In_398,In_1319);
xnor U2410 (N_2410,In_1106,In_670);
xor U2411 (N_2411,In_668,In_709);
nand U2412 (N_2412,In_511,In_974);
or U2413 (N_2413,In_478,In_1436);
and U2414 (N_2414,In_685,In_1085);
and U2415 (N_2415,In_1116,In_957);
and U2416 (N_2416,In_219,In_1425);
or U2417 (N_2417,In_198,In_1304);
nor U2418 (N_2418,In_1461,In_1071);
nor U2419 (N_2419,In_21,In_1307);
nor U2420 (N_2420,In_44,In_803);
or U2421 (N_2421,In_1062,In_978);
nor U2422 (N_2422,In_1401,In_530);
nand U2423 (N_2423,In_70,In_698);
and U2424 (N_2424,In_432,In_443);
and U2425 (N_2425,In_995,In_752);
xor U2426 (N_2426,In_128,In_1173);
nand U2427 (N_2427,In_422,In_1233);
nor U2428 (N_2428,In_546,In_1449);
xnor U2429 (N_2429,In_668,In_1177);
xnor U2430 (N_2430,In_1447,In_143);
or U2431 (N_2431,In_550,In_280);
xor U2432 (N_2432,In_144,In_1382);
or U2433 (N_2433,In_1041,In_640);
and U2434 (N_2434,In_403,In_653);
or U2435 (N_2435,In_1469,In_665);
nor U2436 (N_2436,In_39,In_40);
or U2437 (N_2437,In_332,In_1238);
and U2438 (N_2438,In_1366,In_955);
and U2439 (N_2439,In_1498,In_1249);
nand U2440 (N_2440,In_244,In_994);
and U2441 (N_2441,In_376,In_573);
nor U2442 (N_2442,In_373,In_361);
and U2443 (N_2443,In_1294,In_1363);
nor U2444 (N_2444,In_468,In_1483);
and U2445 (N_2445,In_1331,In_645);
xor U2446 (N_2446,In_977,In_1202);
or U2447 (N_2447,In_1061,In_948);
nand U2448 (N_2448,In_114,In_928);
xor U2449 (N_2449,In_1111,In_238);
or U2450 (N_2450,In_600,In_1393);
and U2451 (N_2451,In_1098,In_1);
xnor U2452 (N_2452,In_1055,In_1028);
nor U2453 (N_2453,In_432,In_916);
and U2454 (N_2454,In_527,In_783);
and U2455 (N_2455,In_1207,In_303);
and U2456 (N_2456,In_376,In_1159);
nor U2457 (N_2457,In_1024,In_34);
nand U2458 (N_2458,In_831,In_937);
xor U2459 (N_2459,In_298,In_1064);
xor U2460 (N_2460,In_1225,In_633);
and U2461 (N_2461,In_1361,In_877);
nand U2462 (N_2462,In_974,In_1202);
and U2463 (N_2463,In_663,In_220);
nand U2464 (N_2464,In_983,In_489);
nand U2465 (N_2465,In_1393,In_1159);
or U2466 (N_2466,In_312,In_452);
nor U2467 (N_2467,In_721,In_328);
and U2468 (N_2468,In_303,In_117);
nand U2469 (N_2469,In_394,In_58);
xor U2470 (N_2470,In_0,In_1280);
and U2471 (N_2471,In_314,In_530);
nand U2472 (N_2472,In_736,In_897);
nand U2473 (N_2473,In_401,In_694);
and U2474 (N_2474,In_528,In_1143);
and U2475 (N_2475,In_893,In_258);
and U2476 (N_2476,In_311,In_1061);
and U2477 (N_2477,In_218,In_912);
and U2478 (N_2478,In_37,In_1197);
nor U2479 (N_2479,In_858,In_1040);
or U2480 (N_2480,In_1010,In_834);
nor U2481 (N_2481,In_1439,In_595);
or U2482 (N_2482,In_1239,In_744);
nor U2483 (N_2483,In_1428,In_339);
nand U2484 (N_2484,In_300,In_373);
nand U2485 (N_2485,In_653,In_1350);
nand U2486 (N_2486,In_334,In_1058);
nand U2487 (N_2487,In_355,In_582);
nand U2488 (N_2488,In_378,In_1039);
xor U2489 (N_2489,In_170,In_250);
nand U2490 (N_2490,In_532,In_89);
and U2491 (N_2491,In_42,In_1463);
or U2492 (N_2492,In_1042,In_1170);
nand U2493 (N_2493,In_1277,In_492);
nor U2494 (N_2494,In_774,In_574);
or U2495 (N_2495,In_457,In_271);
and U2496 (N_2496,In_1066,In_749);
nand U2497 (N_2497,In_988,In_1323);
or U2498 (N_2498,In_1345,In_291);
and U2499 (N_2499,In_1347,In_565);
nand U2500 (N_2500,In_825,In_782);
or U2501 (N_2501,In_553,In_605);
nand U2502 (N_2502,In_21,In_943);
nand U2503 (N_2503,In_426,In_1187);
or U2504 (N_2504,In_1464,In_1186);
nor U2505 (N_2505,In_528,In_1227);
xor U2506 (N_2506,In_1212,In_372);
and U2507 (N_2507,In_1420,In_875);
and U2508 (N_2508,In_287,In_1415);
or U2509 (N_2509,In_1198,In_249);
and U2510 (N_2510,In_1270,In_1047);
or U2511 (N_2511,In_527,In_1049);
xnor U2512 (N_2512,In_1291,In_1316);
nor U2513 (N_2513,In_881,In_1166);
nand U2514 (N_2514,In_899,In_1079);
nand U2515 (N_2515,In_192,In_231);
nand U2516 (N_2516,In_584,In_788);
and U2517 (N_2517,In_882,In_632);
nand U2518 (N_2518,In_564,In_122);
and U2519 (N_2519,In_494,In_810);
or U2520 (N_2520,In_515,In_348);
and U2521 (N_2521,In_1018,In_1333);
xor U2522 (N_2522,In_377,In_1318);
or U2523 (N_2523,In_819,In_295);
nand U2524 (N_2524,In_105,In_364);
nor U2525 (N_2525,In_913,In_262);
xnor U2526 (N_2526,In_464,In_345);
and U2527 (N_2527,In_465,In_817);
nor U2528 (N_2528,In_737,In_1463);
and U2529 (N_2529,In_28,In_910);
or U2530 (N_2530,In_796,In_1032);
xnor U2531 (N_2531,In_1026,In_1067);
nor U2532 (N_2532,In_1334,In_82);
nand U2533 (N_2533,In_493,In_1088);
nand U2534 (N_2534,In_674,In_1335);
or U2535 (N_2535,In_418,In_1117);
nor U2536 (N_2536,In_272,In_378);
or U2537 (N_2537,In_1346,In_1321);
or U2538 (N_2538,In_752,In_451);
nor U2539 (N_2539,In_502,In_522);
and U2540 (N_2540,In_277,In_32);
and U2541 (N_2541,In_192,In_1005);
nor U2542 (N_2542,In_962,In_425);
and U2543 (N_2543,In_65,In_970);
or U2544 (N_2544,In_928,In_1040);
nor U2545 (N_2545,In_1044,In_1170);
nor U2546 (N_2546,In_522,In_1197);
nor U2547 (N_2547,In_67,In_779);
and U2548 (N_2548,In_742,In_269);
and U2549 (N_2549,In_375,In_202);
or U2550 (N_2550,In_377,In_690);
nand U2551 (N_2551,In_400,In_1338);
nor U2552 (N_2552,In_240,In_39);
and U2553 (N_2553,In_104,In_1434);
nand U2554 (N_2554,In_1305,In_1363);
nor U2555 (N_2555,In_1146,In_48);
nand U2556 (N_2556,In_388,In_860);
xnor U2557 (N_2557,In_689,In_1417);
nor U2558 (N_2558,In_983,In_1046);
and U2559 (N_2559,In_39,In_1350);
or U2560 (N_2560,In_1152,In_250);
and U2561 (N_2561,In_114,In_856);
and U2562 (N_2562,In_1010,In_1371);
and U2563 (N_2563,In_481,In_804);
nor U2564 (N_2564,In_1082,In_1040);
or U2565 (N_2565,In_1330,In_1292);
nor U2566 (N_2566,In_1040,In_354);
nand U2567 (N_2567,In_651,In_36);
or U2568 (N_2568,In_698,In_1348);
and U2569 (N_2569,In_722,In_400);
and U2570 (N_2570,In_670,In_400);
or U2571 (N_2571,In_1232,In_706);
and U2572 (N_2572,In_385,In_967);
and U2573 (N_2573,In_892,In_1159);
xnor U2574 (N_2574,In_1228,In_1414);
and U2575 (N_2575,In_588,In_1309);
or U2576 (N_2576,In_1141,In_467);
xor U2577 (N_2577,In_422,In_460);
or U2578 (N_2578,In_293,In_1442);
or U2579 (N_2579,In_574,In_40);
or U2580 (N_2580,In_347,In_844);
or U2581 (N_2581,In_1095,In_477);
nand U2582 (N_2582,In_1405,In_1491);
and U2583 (N_2583,In_840,In_315);
or U2584 (N_2584,In_951,In_1451);
and U2585 (N_2585,In_971,In_887);
nand U2586 (N_2586,In_866,In_652);
or U2587 (N_2587,In_1196,In_1192);
and U2588 (N_2588,In_1230,In_379);
or U2589 (N_2589,In_1298,In_1185);
and U2590 (N_2590,In_859,In_1416);
nand U2591 (N_2591,In_1315,In_1022);
xnor U2592 (N_2592,In_1027,In_1357);
xor U2593 (N_2593,In_628,In_1373);
xor U2594 (N_2594,In_52,In_948);
nor U2595 (N_2595,In_1476,In_1046);
or U2596 (N_2596,In_506,In_677);
nand U2597 (N_2597,In_868,In_16);
and U2598 (N_2598,In_1098,In_462);
nand U2599 (N_2599,In_782,In_9);
or U2600 (N_2600,In_676,In_1306);
nor U2601 (N_2601,In_1111,In_210);
nand U2602 (N_2602,In_1291,In_678);
and U2603 (N_2603,In_560,In_1153);
and U2604 (N_2604,In_171,In_23);
nand U2605 (N_2605,In_811,In_517);
nand U2606 (N_2606,In_270,In_1447);
and U2607 (N_2607,In_376,In_1295);
nor U2608 (N_2608,In_341,In_168);
and U2609 (N_2609,In_794,In_1326);
nor U2610 (N_2610,In_913,In_260);
and U2611 (N_2611,In_92,In_919);
nand U2612 (N_2612,In_411,In_587);
nand U2613 (N_2613,In_1097,In_106);
or U2614 (N_2614,In_1049,In_217);
and U2615 (N_2615,In_798,In_665);
nor U2616 (N_2616,In_708,In_1155);
nand U2617 (N_2617,In_1001,In_977);
and U2618 (N_2618,In_776,In_1285);
nand U2619 (N_2619,In_283,In_252);
and U2620 (N_2620,In_1271,In_698);
nand U2621 (N_2621,In_721,In_326);
or U2622 (N_2622,In_359,In_684);
or U2623 (N_2623,In_397,In_1104);
xnor U2624 (N_2624,In_256,In_986);
nor U2625 (N_2625,In_727,In_589);
nand U2626 (N_2626,In_685,In_1354);
nor U2627 (N_2627,In_636,In_903);
nor U2628 (N_2628,In_667,In_214);
nor U2629 (N_2629,In_1248,In_909);
nand U2630 (N_2630,In_235,In_1219);
and U2631 (N_2631,In_1433,In_1468);
or U2632 (N_2632,In_1262,In_1165);
nor U2633 (N_2633,In_1204,In_1110);
and U2634 (N_2634,In_1209,In_1211);
or U2635 (N_2635,In_1313,In_152);
or U2636 (N_2636,In_115,In_1442);
nor U2637 (N_2637,In_1379,In_168);
and U2638 (N_2638,In_1198,In_536);
or U2639 (N_2639,In_518,In_1361);
xor U2640 (N_2640,In_1145,In_414);
or U2641 (N_2641,In_323,In_1322);
nand U2642 (N_2642,In_1115,In_3);
xnor U2643 (N_2643,In_1172,In_1456);
or U2644 (N_2644,In_999,In_287);
and U2645 (N_2645,In_454,In_759);
and U2646 (N_2646,In_178,In_950);
nand U2647 (N_2647,In_334,In_711);
or U2648 (N_2648,In_239,In_421);
or U2649 (N_2649,In_747,In_12);
nand U2650 (N_2650,In_195,In_1128);
and U2651 (N_2651,In_344,In_1240);
and U2652 (N_2652,In_878,In_1306);
nand U2653 (N_2653,In_268,In_1257);
nor U2654 (N_2654,In_414,In_345);
and U2655 (N_2655,In_676,In_1284);
nor U2656 (N_2656,In_853,In_524);
and U2657 (N_2657,In_1238,In_72);
or U2658 (N_2658,In_101,In_29);
and U2659 (N_2659,In_494,In_894);
xor U2660 (N_2660,In_988,In_21);
or U2661 (N_2661,In_589,In_700);
nor U2662 (N_2662,In_1201,In_174);
or U2663 (N_2663,In_828,In_530);
nor U2664 (N_2664,In_1110,In_1198);
xor U2665 (N_2665,In_857,In_1286);
or U2666 (N_2666,In_423,In_1128);
xor U2667 (N_2667,In_495,In_525);
or U2668 (N_2668,In_37,In_336);
and U2669 (N_2669,In_580,In_451);
nor U2670 (N_2670,In_1314,In_148);
nand U2671 (N_2671,In_950,In_587);
nor U2672 (N_2672,In_539,In_529);
or U2673 (N_2673,In_697,In_479);
or U2674 (N_2674,In_411,In_69);
or U2675 (N_2675,In_979,In_513);
nand U2676 (N_2676,In_717,In_1023);
nand U2677 (N_2677,In_816,In_727);
nand U2678 (N_2678,In_302,In_1134);
nor U2679 (N_2679,In_101,In_151);
or U2680 (N_2680,In_511,In_728);
or U2681 (N_2681,In_19,In_178);
and U2682 (N_2682,In_854,In_936);
nand U2683 (N_2683,In_570,In_1308);
nor U2684 (N_2684,In_60,In_1220);
nand U2685 (N_2685,In_1065,In_537);
or U2686 (N_2686,In_117,In_1391);
xor U2687 (N_2687,In_621,In_54);
nor U2688 (N_2688,In_633,In_112);
or U2689 (N_2689,In_1345,In_295);
nor U2690 (N_2690,In_689,In_1118);
nor U2691 (N_2691,In_809,In_53);
nand U2692 (N_2692,In_1110,In_486);
or U2693 (N_2693,In_1344,In_36);
nand U2694 (N_2694,In_681,In_1182);
nand U2695 (N_2695,In_773,In_38);
nor U2696 (N_2696,In_165,In_41);
nor U2697 (N_2697,In_820,In_36);
and U2698 (N_2698,In_888,In_1197);
and U2699 (N_2699,In_429,In_159);
nor U2700 (N_2700,In_1132,In_412);
nand U2701 (N_2701,In_107,In_240);
xor U2702 (N_2702,In_263,In_62);
nand U2703 (N_2703,In_229,In_555);
nor U2704 (N_2704,In_824,In_524);
and U2705 (N_2705,In_1132,In_991);
or U2706 (N_2706,In_672,In_307);
nand U2707 (N_2707,In_831,In_441);
and U2708 (N_2708,In_1175,In_602);
and U2709 (N_2709,In_709,In_1268);
nor U2710 (N_2710,In_502,In_694);
xnor U2711 (N_2711,In_1200,In_60);
nand U2712 (N_2712,In_454,In_56);
and U2713 (N_2713,In_901,In_1163);
or U2714 (N_2714,In_1100,In_684);
nor U2715 (N_2715,In_1421,In_824);
nand U2716 (N_2716,In_18,In_1054);
nand U2717 (N_2717,In_90,In_334);
nand U2718 (N_2718,In_1033,In_1478);
or U2719 (N_2719,In_670,In_1451);
nor U2720 (N_2720,In_802,In_80);
and U2721 (N_2721,In_1158,In_1149);
xor U2722 (N_2722,In_751,In_907);
nand U2723 (N_2723,In_1371,In_121);
or U2724 (N_2724,In_1440,In_1069);
nor U2725 (N_2725,In_1068,In_155);
or U2726 (N_2726,In_632,In_772);
nor U2727 (N_2727,In_1144,In_1228);
nor U2728 (N_2728,In_218,In_285);
and U2729 (N_2729,In_493,In_1086);
xnor U2730 (N_2730,In_531,In_600);
xor U2731 (N_2731,In_1270,In_1267);
and U2732 (N_2732,In_195,In_1108);
nand U2733 (N_2733,In_470,In_1404);
nor U2734 (N_2734,In_1034,In_668);
nand U2735 (N_2735,In_451,In_611);
or U2736 (N_2736,In_806,In_516);
and U2737 (N_2737,In_253,In_245);
nand U2738 (N_2738,In_543,In_183);
or U2739 (N_2739,In_769,In_992);
nor U2740 (N_2740,In_810,In_841);
or U2741 (N_2741,In_48,In_648);
or U2742 (N_2742,In_951,In_155);
or U2743 (N_2743,In_551,In_1054);
and U2744 (N_2744,In_1347,In_1208);
nand U2745 (N_2745,In_779,In_646);
nand U2746 (N_2746,In_31,In_314);
and U2747 (N_2747,In_975,In_884);
and U2748 (N_2748,In_274,In_42);
and U2749 (N_2749,In_653,In_1030);
or U2750 (N_2750,In_1199,In_0);
nor U2751 (N_2751,In_1309,In_1019);
nor U2752 (N_2752,In_243,In_911);
nand U2753 (N_2753,In_241,In_117);
nand U2754 (N_2754,In_755,In_1273);
and U2755 (N_2755,In_713,In_85);
and U2756 (N_2756,In_579,In_1205);
nand U2757 (N_2757,In_1378,In_449);
nor U2758 (N_2758,In_506,In_443);
and U2759 (N_2759,In_1368,In_4);
nand U2760 (N_2760,In_976,In_728);
nand U2761 (N_2761,In_88,In_502);
nor U2762 (N_2762,In_1248,In_969);
xor U2763 (N_2763,In_278,In_1205);
nand U2764 (N_2764,In_898,In_1315);
or U2765 (N_2765,In_178,In_132);
nand U2766 (N_2766,In_160,In_231);
or U2767 (N_2767,In_1196,In_1210);
nand U2768 (N_2768,In_227,In_958);
nor U2769 (N_2769,In_1315,In_1228);
nand U2770 (N_2770,In_1467,In_1280);
xnor U2771 (N_2771,In_517,In_133);
nand U2772 (N_2772,In_1320,In_946);
and U2773 (N_2773,In_55,In_334);
xor U2774 (N_2774,In_560,In_938);
or U2775 (N_2775,In_1359,In_163);
and U2776 (N_2776,In_335,In_138);
or U2777 (N_2777,In_996,In_474);
nand U2778 (N_2778,In_1321,In_39);
or U2779 (N_2779,In_654,In_514);
or U2780 (N_2780,In_1264,In_1055);
xnor U2781 (N_2781,In_497,In_216);
nand U2782 (N_2782,In_5,In_1487);
and U2783 (N_2783,In_1118,In_948);
nand U2784 (N_2784,In_386,In_991);
or U2785 (N_2785,In_1476,In_135);
nor U2786 (N_2786,In_1382,In_170);
xnor U2787 (N_2787,In_1018,In_752);
nand U2788 (N_2788,In_1379,In_1122);
xor U2789 (N_2789,In_1143,In_650);
or U2790 (N_2790,In_78,In_182);
and U2791 (N_2791,In_1404,In_211);
and U2792 (N_2792,In_295,In_1207);
xnor U2793 (N_2793,In_968,In_1145);
xnor U2794 (N_2794,In_621,In_1158);
nor U2795 (N_2795,In_83,In_149);
xnor U2796 (N_2796,In_1215,In_270);
and U2797 (N_2797,In_1154,In_516);
or U2798 (N_2798,In_780,In_1120);
nand U2799 (N_2799,In_586,In_969);
or U2800 (N_2800,In_585,In_5);
and U2801 (N_2801,In_1363,In_1166);
and U2802 (N_2802,In_106,In_1013);
nand U2803 (N_2803,In_351,In_562);
and U2804 (N_2804,In_714,In_437);
nand U2805 (N_2805,In_1363,In_1008);
nand U2806 (N_2806,In_928,In_817);
and U2807 (N_2807,In_1005,In_1458);
nand U2808 (N_2808,In_1088,In_1063);
nand U2809 (N_2809,In_670,In_506);
or U2810 (N_2810,In_1160,In_958);
nand U2811 (N_2811,In_551,In_755);
nand U2812 (N_2812,In_874,In_1431);
nand U2813 (N_2813,In_197,In_31);
nand U2814 (N_2814,In_250,In_341);
or U2815 (N_2815,In_209,In_1144);
and U2816 (N_2816,In_1328,In_1306);
and U2817 (N_2817,In_1008,In_670);
or U2818 (N_2818,In_1328,In_73);
nand U2819 (N_2819,In_811,In_949);
nand U2820 (N_2820,In_874,In_387);
nor U2821 (N_2821,In_324,In_390);
and U2822 (N_2822,In_1331,In_1016);
and U2823 (N_2823,In_602,In_2);
nand U2824 (N_2824,In_543,In_610);
nor U2825 (N_2825,In_937,In_1268);
or U2826 (N_2826,In_706,In_312);
and U2827 (N_2827,In_426,In_919);
nor U2828 (N_2828,In_14,In_172);
and U2829 (N_2829,In_409,In_1153);
nor U2830 (N_2830,In_1064,In_797);
nand U2831 (N_2831,In_769,In_13);
or U2832 (N_2832,In_1452,In_1344);
or U2833 (N_2833,In_1466,In_844);
and U2834 (N_2834,In_365,In_612);
and U2835 (N_2835,In_1177,In_393);
or U2836 (N_2836,In_779,In_259);
or U2837 (N_2837,In_371,In_1148);
nor U2838 (N_2838,In_630,In_1128);
and U2839 (N_2839,In_1424,In_912);
nor U2840 (N_2840,In_606,In_1024);
and U2841 (N_2841,In_700,In_237);
and U2842 (N_2842,In_303,In_103);
xor U2843 (N_2843,In_216,In_462);
or U2844 (N_2844,In_609,In_898);
or U2845 (N_2845,In_1218,In_1280);
nor U2846 (N_2846,In_402,In_510);
nand U2847 (N_2847,In_581,In_1277);
nor U2848 (N_2848,In_809,In_416);
xor U2849 (N_2849,In_1201,In_1376);
nand U2850 (N_2850,In_867,In_800);
xnor U2851 (N_2851,In_1152,In_1300);
and U2852 (N_2852,In_579,In_1099);
nor U2853 (N_2853,In_987,In_1271);
nor U2854 (N_2854,In_889,In_535);
and U2855 (N_2855,In_817,In_860);
and U2856 (N_2856,In_996,In_306);
nor U2857 (N_2857,In_1469,In_947);
nor U2858 (N_2858,In_852,In_697);
and U2859 (N_2859,In_1126,In_977);
nand U2860 (N_2860,In_1052,In_1088);
nor U2861 (N_2861,In_676,In_148);
or U2862 (N_2862,In_915,In_601);
or U2863 (N_2863,In_535,In_1269);
nand U2864 (N_2864,In_34,In_1151);
nand U2865 (N_2865,In_846,In_356);
nand U2866 (N_2866,In_299,In_320);
nor U2867 (N_2867,In_288,In_422);
nand U2868 (N_2868,In_761,In_318);
and U2869 (N_2869,In_1420,In_116);
or U2870 (N_2870,In_784,In_1375);
nor U2871 (N_2871,In_273,In_1009);
nor U2872 (N_2872,In_362,In_224);
and U2873 (N_2873,In_684,In_1366);
and U2874 (N_2874,In_46,In_271);
nand U2875 (N_2875,In_1004,In_734);
nand U2876 (N_2876,In_557,In_781);
and U2877 (N_2877,In_624,In_263);
and U2878 (N_2878,In_589,In_731);
nand U2879 (N_2879,In_436,In_11);
or U2880 (N_2880,In_1422,In_371);
xnor U2881 (N_2881,In_850,In_1406);
or U2882 (N_2882,In_1326,In_159);
or U2883 (N_2883,In_1153,In_532);
and U2884 (N_2884,In_1347,In_827);
xnor U2885 (N_2885,In_74,In_1083);
nor U2886 (N_2886,In_1498,In_979);
nor U2887 (N_2887,In_1014,In_796);
nand U2888 (N_2888,In_350,In_1189);
or U2889 (N_2889,In_1282,In_1478);
or U2890 (N_2890,In_1305,In_144);
nor U2891 (N_2891,In_1212,In_363);
nor U2892 (N_2892,In_1228,In_1003);
nor U2893 (N_2893,In_1306,In_315);
xnor U2894 (N_2894,In_1170,In_227);
nand U2895 (N_2895,In_1221,In_524);
and U2896 (N_2896,In_1134,In_684);
or U2897 (N_2897,In_568,In_801);
nand U2898 (N_2898,In_775,In_1206);
and U2899 (N_2899,In_622,In_424);
or U2900 (N_2900,In_1422,In_400);
nor U2901 (N_2901,In_1234,In_531);
nor U2902 (N_2902,In_50,In_167);
xnor U2903 (N_2903,In_448,In_908);
or U2904 (N_2904,In_1300,In_689);
and U2905 (N_2905,In_526,In_762);
nand U2906 (N_2906,In_495,In_346);
and U2907 (N_2907,In_892,In_1054);
nand U2908 (N_2908,In_603,In_332);
nor U2909 (N_2909,In_92,In_956);
nand U2910 (N_2910,In_606,In_697);
nor U2911 (N_2911,In_480,In_651);
nor U2912 (N_2912,In_124,In_762);
nor U2913 (N_2913,In_911,In_934);
or U2914 (N_2914,In_1228,In_1300);
nand U2915 (N_2915,In_1007,In_1479);
and U2916 (N_2916,In_708,In_1354);
nor U2917 (N_2917,In_1149,In_1437);
or U2918 (N_2918,In_709,In_1360);
and U2919 (N_2919,In_698,In_1180);
nor U2920 (N_2920,In_579,In_765);
or U2921 (N_2921,In_1471,In_1378);
nor U2922 (N_2922,In_1006,In_256);
and U2923 (N_2923,In_237,In_1004);
and U2924 (N_2924,In_23,In_1210);
nand U2925 (N_2925,In_317,In_287);
and U2926 (N_2926,In_833,In_1021);
nand U2927 (N_2927,In_1446,In_1345);
and U2928 (N_2928,In_1421,In_870);
nor U2929 (N_2929,In_1355,In_1326);
or U2930 (N_2930,In_862,In_808);
and U2931 (N_2931,In_87,In_148);
or U2932 (N_2932,In_1093,In_231);
nor U2933 (N_2933,In_155,In_313);
nor U2934 (N_2934,In_994,In_446);
xor U2935 (N_2935,In_896,In_915);
and U2936 (N_2936,In_767,In_424);
nand U2937 (N_2937,In_1091,In_39);
or U2938 (N_2938,In_427,In_218);
xor U2939 (N_2939,In_1213,In_522);
nor U2940 (N_2940,In_884,In_1003);
nor U2941 (N_2941,In_25,In_37);
nor U2942 (N_2942,In_632,In_927);
or U2943 (N_2943,In_67,In_208);
and U2944 (N_2944,In_758,In_528);
or U2945 (N_2945,In_426,In_763);
and U2946 (N_2946,In_614,In_84);
nand U2947 (N_2947,In_113,In_264);
xnor U2948 (N_2948,In_859,In_1413);
and U2949 (N_2949,In_138,In_592);
nor U2950 (N_2950,In_795,In_1176);
nor U2951 (N_2951,In_617,In_111);
or U2952 (N_2952,In_683,In_500);
or U2953 (N_2953,In_412,In_892);
xnor U2954 (N_2954,In_1495,In_160);
nand U2955 (N_2955,In_1074,In_365);
nand U2956 (N_2956,In_182,In_1082);
nand U2957 (N_2957,In_1448,In_383);
nor U2958 (N_2958,In_1143,In_573);
or U2959 (N_2959,In_1467,In_389);
xnor U2960 (N_2960,In_892,In_420);
nor U2961 (N_2961,In_1317,In_364);
xor U2962 (N_2962,In_661,In_1019);
nand U2963 (N_2963,In_1006,In_515);
nor U2964 (N_2964,In_32,In_196);
nor U2965 (N_2965,In_38,In_101);
and U2966 (N_2966,In_67,In_752);
nand U2967 (N_2967,In_955,In_1171);
or U2968 (N_2968,In_370,In_275);
or U2969 (N_2969,In_1270,In_563);
or U2970 (N_2970,In_433,In_297);
and U2971 (N_2971,In_57,In_225);
nor U2972 (N_2972,In_1085,In_782);
nor U2973 (N_2973,In_1023,In_615);
and U2974 (N_2974,In_1486,In_625);
nand U2975 (N_2975,In_321,In_1112);
and U2976 (N_2976,In_103,In_399);
xnor U2977 (N_2977,In_1108,In_1460);
and U2978 (N_2978,In_1299,In_167);
or U2979 (N_2979,In_1423,In_1186);
nor U2980 (N_2980,In_133,In_1159);
and U2981 (N_2981,In_339,In_1042);
nand U2982 (N_2982,In_467,In_1398);
or U2983 (N_2983,In_893,In_919);
and U2984 (N_2984,In_183,In_814);
nand U2985 (N_2985,In_162,In_619);
and U2986 (N_2986,In_972,In_453);
and U2987 (N_2987,In_1235,In_1363);
nor U2988 (N_2988,In_1241,In_773);
or U2989 (N_2989,In_759,In_64);
nor U2990 (N_2990,In_487,In_25);
or U2991 (N_2991,In_523,In_1246);
nand U2992 (N_2992,In_362,In_1436);
nor U2993 (N_2993,In_955,In_169);
xnor U2994 (N_2994,In_768,In_715);
and U2995 (N_2995,In_848,In_305);
and U2996 (N_2996,In_1442,In_882);
or U2997 (N_2997,In_12,In_240);
or U2998 (N_2998,In_913,In_1179);
nand U2999 (N_2999,In_1156,In_64);
and U3000 (N_3000,N_1162,N_742);
nand U3001 (N_3001,N_1490,N_199);
nand U3002 (N_3002,N_1718,N_2125);
or U3003 (N_3003,N_1966,N_1370);
and U3004 (N_3004,N_498,N_1601);
nor U3005 (N_3005,N_2577,N_2860);
or U3006 (N_3006,N_258,N_2554);
nor U3007 (N_3007,N_1137,N_1158);
and U3008 (N_3008,N_226,N_1526);
nor U3009 (N_3009,N_1856,N_56);
and U3010 (N_3010,N_1083,N_906);
and U3011 (N_3011,N_704,N_64);
xor U3012 (N_3012,N_1928,N_329);
nand U3013 (N_3013,N_1198,N_2164);
or U3014 (N_3014,N_1330,N_1834);
and U3015 (N_3015,N_438,N_2962);
nand U3016 (N_3016,N_2438,N_124);
and U3017 (N_3017,N_2705,N_2160);
xnor U3018 (N_3018,N_1958,N_2474);
and U3019 (N_3019,N_2206,N_1295);
nor U3020 (N_3020,N_2730,N_545);
or U3021 (N_3021,N_1345,N_730);
and U3022 (N_3022,N_17,N_988);
and U3023 (N_3023,N_1393,N_2139);
or U3024 (N_3024,N_2996,N_1402);
nor U3025 (N_3025,N_2159,N_1418);
xnor U3026 (N_3026,N_844,N_1863);
and U3027 (N_3027,N_2243,N_1236);
nand U3028 (N_3028,N_2685,N_965);
nand U3029 (N_3029,N_1914,N_2901);
nor U3030 (N_3030,N_721,N_1964);
nor U3031 (N_3031,N_2064,N_1397);
nor U3032 (N_3032,N_2426,N_436);
nand U3033 (N_3033,N_1617,N_785);
and U3034 (N_3034,N_2497,N_2609);
xor U3035 (N_3035,N_2382,N_2462);
xor U3036 (N_3036,N_1380,N_584);
nor U3037 (N_3037,N_2496,N_29);
and U3038 (N_3038,N_1484,N_2407);
and U3039 (N_3039,N_1520,N_84);
or U3040 (N_3040,N_1460,N_132);
or U3041 (N_3041,N_2072,N_678);
xnor U3042 (N_3042,N_1637,N_1682);
nand U3043 (N_3043,N_2572,N_107);
nor U3044 (N_3044,N_2356,N_2930);
or U3045 (N_3045,N_578,N_316);
and U3046 (N_3046,N_2748,N_1759);
and U3047 (N_3047,N_2334,N_1245);
nand U3048 (N_3048,N_2921,N_1736);
nor U3049 (N_3049,N_2693,N_1780);
nor U3050 (N_3050,N_1716,N_1726);
and U3051 (N_3051,N_298,N_2684);
or U3052 (N_3052,N_1364,N_2044);
nand U3053 (N_3053,N_2217,N_2654);
or U3054 (N_3054,N_469,N_2936);
or U3055 (N_3055,N_1949,N_1085);
xor U3056 (N_3056,N_2415,N_273);
and U3057 (N_3057,N_1668,N_2652);
nor U3058 (N_3058,N_2276,N_1240);
nand U3059 (N_3059,N_1891,N_2491);
or U3060 (N_3060,N_2175,N_2897);
and U3061 (N_3061,N_1292,N_2545);
and U3062 (N_3062,N_1803,N_2723);
nor U3063 (N_3063,N_1406,N_2547);
nor U3064 (N_3064,N_1093,N_45);
or U3065 (N_3065,N_253,N_1416);
or U3066 (N_3066,N_2953,N_708);
or U3067 (N_3067,N_1235,N_143);
nand U3068 (N_3068,N_523,N_604);
and U3069 (N_3069,N_1183,N_2863);
xor U3070 (N_3070,N_2477,N_1409);
nand U3071 (N_3071,N_2784,N_1392);
and U3072 (N_3072,N_2190,N_2445);
or U3073 (N_3073,N_1150,N_950);
or U3074 (N_3074,N_1355,N_145);
and U3075 (N_3075,N_1514,N_1212);
nor U3076 (N_3076,N_2738,N_512);
nor U3077 (N_3077,N_2137,N_1979);
and U3078 (N_3078,N_840,N_2218);
or U3079 (N_3079,N_756,N_2941);
or U3080 (N_3080,N_2511,N_789);
nor U3081 (N_3081,N_2879,N_1388);
nor U3082 (N_3082,N_1847,N_419);
or U3083 (N_3083,N_2963,N_414);
and U3084 (N_3084,N_1200,N_1133);
nand U3085 (N_3085,N_1519,N_2914);
nand U3086 (N_3086,N_1322,N_2655);
nand U3087 (N_3087,N_234,N_1850);
and U3088 (N_3088,N_1268,N_1907);
nand U3089 (N_3089,N_717,N_1925);
and U3090 (N_3090,N_2246,N_1144);
nor U3091 (N_3091,N_1291,N_562);
or U3092 (N_3092,N_2856,N_2595);
nand U3093 (N_3093,N_1404,N_311);
and U3094 (N_3094,N_1366,N_1115);
and U3095 (N_3095,N_1274,N_1211);
or U3096 (N_3096,N_2665,N_751);
or U3097 (N_3097,N_247,N_2024);
nand U3098 (N_3098,N_2455,N_916);
nor U3099 (N_3099,N_2877,N_698);
nor U3100 (N_3100,N_763,N_2145);
nor U3101 (N_3101,N_2295,N_215);
or U3102 (N_3102,N_640,N_392);
and U3103 (N_3103,N_860,N_799);
nand U3104 (N_3104,N_2297,N_1511);
or U3105 (N_3105,N_2339,N_144);
nand U3106 (N_3106,N_172,N_75);
nand U3107 (N_3107,N_2363,N_2308);
nand U3108 (N_3108,N_1636,N_672);
or U3109 (N_3109,N_82,N_1510);
or U3110 (N_3110,N_2107,N_384);
and U3111 (N_3111,N_2696,N_2481);
nor U3112 (N_3112,N_2593,N_125);
nor U3113 (N_3113,N_2326,N_1614);
nand U3114 (N_3114,N_126,N_1230);
nor U3115 (N_3115,N_2759,N_2940);
nand U3116 (N_3116,N_520,N_798);
and U3117 (N_3117,N_286,N_1571);
or U3118 (N_3118,N_2031,N_855);
nand U3119 (N_3119,N_1646,N_301);
nand U3120 (N_3120,N_2893,N_1018);
and U3121 (N_3121,N_1023,N_1662);
xor U3122 (N_3122,N_1982,N_2235);
nand U3123 (N_3123,N_2776,N_2765);
xor U3124 (N_3124,N_1942,N_2550);
or U3125 (N_3125,N_170,N_1604);
and U3126 (N_3126,N_1440,N_2868);
or U3127 (N_3127,N_2883,N_1621);
or U3128 (N_3128,N_1879,N_448);
nand U3129 (N_3129,N_493,N_2488);
or U3130 (N_3130,N_2985,N_2715);
nand U3131 (N_3131,N_2974,N_2752);
and U3132 (N_3132,N_2196,N_2848);
and U3133 (N_3133,N_2179,N_423);
and U3134 (N_3134,N_1499,N_1913);
xor U3135 (N_3135,N_1170,N_1715);
and U3136 (N_3136,N_1990,N_2116);
nor U3137 (N_3137,N_2420,N_1316);
or U3138 (N_3138,N_150,N_2878);
or U3139 (N_3139,N_591,N_1528);
nand U3140 (N_3140,N_2251,N_1625);
nand U3141 (N_3141,N_1559,N_995);
and U3142 (N_3142,N_2074,N_446);
nor U3143 (N_3143,N_961,N_984);
nor U3144 (N_3144,N_325,N_675);
and U3145 (N_3145,N_2129,N_2626);
and U3146 (N_3146,N_2512,N_921);
or U3147 (N_3147,N_1785,N_1313);
nor U3148 (N_3148,N_1497,N_676);
xor U3149 (N_3149,N_2051,N_1727);
nand U3150 (N_3150,N_1870,N_412);
and U3151 (N_3151,N_1813,N_1975);
or U3152 (N_3152,N_1744,N_935);
nand U3153 (N_3153,N_2305,N_1096);
and U3154 (N_3154,N_34,N_2845);
or U3155 (N_3155,N_2908,N_1581);
nand U3156 (N_3156,N_1831,N_1037);
and U3157 (N_3157,N_2011,N_352);
and U3158 (N_3158,N_1413,N_1858);
nor U3159 (N_3159,N_868,N_1420);
nor U3160 (N_3160,N_979,N_2102);
nand U3161 (N_3161,N_2084,N_910);
or U3162 (N_3162,N_2726,N_2358);
nand U3163 (N_3163,N_953,N_2714);
and U3164 (N_3164,N_38,N_758);
and U3165 (N_3165,N_1303,N_2866);
nand U3166 (N_3166,N_1052,N_2795);
xnor U3167 (N_3167,N_2742,N_2805);
nor U3168 (N_3168,N_1675,N_831);
or U3169 (N_3169,N_1441,N_408);
nand U3170 (N_3170,N_440,N_1740);
xor U3171 (N_3171,N_175,N_2144);
and U3172 (N_3172,N_2884,N_2046);
and U3173 (N_3173,N_1560,N_944);
or U3174 (N_3174,N_942,N_36);
and U3175 (N_3175,N_1221,N_123);
nor U3176 (N_3176,N_926,N_5);
nor U3177 (N_3177,N_715,N_1408);
xor U3178 (N_3178,N_2029,N_195);
nand U3179 (N_3179,N_333,N_1729);
xor U3180 (N_3180,N_713,N_573);
nor U3181 (N_3181,N_1157,N_154);
nor U3182 (N_3182,N_1830,N_236);
nand U3183 (N_3183,N_1061,N_1905);
nor U3184 (N_3184,N_239,N_687);
and U3185 (N_3185,N_1709,N_92);
or U3186 (N_3186,N_2777,N_1011);
nand U3187 (N_3187,N_2331,N_1635);
or U3188 (N_3188,N_572,N_769);
or U3189 (N_3189,N_393,N_2118);
nand U3190 (N_3190,N_1687,N_2484);
nor U3191 (N_3191,N_2403,N_2416);
xor U3192 (N_3192,N_2707,N_560);
or U3193 (N_3193,N_473,N_1771);
or U3194 (N_3194,N_96,N_2376);
or U3195 (N_3195,N_1118,N_608);
and U3196 (N_3196,N_1871,N_937);
nor U3197 (N_3197,N_2855,N_1633);
and U3198 (N_3198,N_1993,N_2058);
or U3199 (N_3199,N_2119,N_2389);
xor U3200 (N_3200,N_1462,N_1634);
or U3201 (N_3201,N_1283,N_2008);
nand U3202 (N_3202,N_2713,N_57);
nor U3203 (N_3203,N_2092,N_699);
and U3204 (N_3204,N_1032,N_1590);
xnor U3205 (N_3205,N_2952,N_33);
and U3206 (N_3206,N_692,N_256);
nor U3207 (N_3207,N_2161,N_1923);
and U3208 (N_3208,N_52,N_1678);
xnor U3209 (N_3209,N_2030,N_19);
and U3210 (N_3210,N_207,N_2561);
and U3211 (N_3211,N_960,N_2034);
xnor U3212 (N_3212,N_390,N_167);
nor U3213 (N_3213,N_1181,N_67);
or U3214 (N_3214,N_2183,N_1917);
nor U3215 (N_3215,N_86,N_2386);
xnor U3216 (N_3216,N_2712,N_260);
nor U3217 (N_3217,N_735,N_2900);
or U3218 (N_3218,N_1950,N_1430);
and U3219 (N_3219,N_1789,N_1794);
and U3220 (N_3220,N_2103,N_2247);
xor U3221 (N_3221,N_1491,N_1541);
and U3222 (N_3222,N_2988,N_2898);
nand U3223 (N_3223,N_962,N_1896);
or U3224 (N_3224,N_579,N_2719);
nor U3225 (N_3225,N_2458,N_596);
and U3226 (N_3226,N_196,N_1063);
nor U3227 (N_3227,N_1278,N_2956);
and U3228 (N_3228,N_53,N_1171);
and U3229 (N_3229,N_212,N_775);
nand U3230 (N_3230,N_1049,N_654);
and U3231 (N_3231,N_1802,N_2661);
nand U3232 (N_3232,N_2429,N_1584);
and U3233 (N_3233,N_2670,N_2019);
or U3234 (N_3234,N_2569,N_1536);
or U3235 (N_3235,N_2439,N_1351);
nor U3236 (N_3236,N_569,N_720);
nand U3237 (N_3237,N_1114,N_1358);
and U3238 (N_3238,N_623,N_865);
nand U3239 (N_3239,N_2039,N_2352);
xnor U3240 (N_3240,N_2230,N_2068);
or U3241 (N_3241,N_753,N_1807);
and U3242 (N_3242,N_2851,N_1013);
nor U3243 (N_3243,N_2583,N_2443);
nor U3244 (N_3244,N_1901,N_1963);
nand U3245 (N_3245,N_2923,N_1795);
nor U3246 (N_3246,N_2066,N_2506);
and U3247 (N_3247,N_1055,N_757);
and U3248 (N_3248,N_2990,N_872);
and U3249 (N_3249,N_1693,N_112);
and U3250 (N_3250,N_1009,N_221);
nand U3251 (N_3251,N_537,N_893);
nor U3252 (N_3252,N_1097,N_1199);
or U3253 (N_3253,N_547,N_1855);
or U3254 (N_3254,N_1369,N_718);
or U3255 (N_3255,N_2708,N_2410);
nor U3256 (N_3256,N_80,N_214);
or U3257 (N_3257,N_851,N_1338);
nand U3258 (N_3258,N_1868,N_435);
and U3259 (N_3259,N_94,N_2345);
or U3260 (N_3260,N_1225,N_1796);
and U3261 (N_3261,N_1340,N_561);
nor U3262 (N_3262,N_341,N_543);
nor U3263 (N_3263,N_875,N_1110);
or U3264 (N_3264,N_1640,N_488);
nor U3265 (N_3265,N_565,N_1786);
nor U3266 (N_3266,N_1247,N_531);
nor U3267 (N_3267,N_454,N_922);
nand U3268 (N_3268,N_2819,N_1655);
or U3269 (N_3269,N_402,N_1453);
nor U3270 (N_3270,N_2490,N_2181);
nor U3271 (N_3271,N_1327,N_1166);
nor U3272 (N_3272,N_2966,N_140);
or U3273 (N_3273,N_1600,N_2886);
nor U3274 (N_3274,N_1732,N_2498);
and U3275 (N_3275,N_2465,N_2934);
nand U3276 (N_3276,N_2405,N_1220);
xnor U3277 (N_3277,N_2870,N_306);
or U3278 (N_3278,N_2724,N_2560);
and U3279 (N_3279,N_2005,N_429);
and U3280 (N_3280,N_817,N_670);
and U3281 (N_3281,N_585,N_2434);
nand U3282 (N_3282,N_650,N_2680);
or U3283 (N_3283,N_540,N_554);
and U3284 (N_3284,N_71,N_729);
nand U3285 (N_3285,N_1749,N_2057);
nor U3286 (N_3286,N_2409,N_2796);
or U3287 (N_3287,N_2228,N_193);
nor U3288 (N_3288,N_2307,N_2278);
xnor U3289 (N_3289,N_857,N_2913);
nand U3290 (N_3290,N_2902,N_2033);
and U3291 (N_3291,N_2596,N_85);
and U3292 (N_3292,N_895,N_1232);
nand U3293 (N_3293,N_1937,N_2277);
and U3294 (N_3294,N_828,N_567);
nand U3295 (N_3295,N_2843,N_1981);
nand U3296 (N_3296,N_1007,N_2542);
xor U3297 (N_3297,N_2747,N_609);
xnor U3298 (N_3298,N_1643,N_280);
nor U3299 (N_3299,N_2323,N_237);
and U3300 (N_3300,N_109,N_1546);
or U3301 (N_3301,N_2585,N_778);
xnor U3302 (N_3302,N_497,N_2301);
nand U3303 (N_3303,N_511,N_1681);
or U3304 (N_3304,N_340,N_141);
nor U3305 (N_3305,N_1696,N_1332);
or U3306 (N_3306,N_2385,N_856);
or U3307 (N_3307,N_399,N_2229);
and U3308 (N_3308,N_2091,N_2803);
nand U3309 (N_3309,N_1639,N_2353);
and U3310 (N_3310,N_2627,N_2601);
nand U3311 (N_3311,N_658,N_1280);
nor U3312 (N_3312,N_2060,N_1348);
nor U3313 (N_3313,N_2146,N_1573);
nand U3314 (N_3314,N_1429,N_1034);
nor U3315 (N_3315,N_225,N_1217);
or U3316 (N_3316,N_701,N_1534);
or U3317 (N_3317,N_946,N_1141);
or U3318 (N_3318,N_1906,N_1275);
nand U3319 (N_3319,N_2516,N_1618);
and U3320 (N_3320,N_1190,N_2998);
and U3321 (N_3321,N_1523,N_956);
nor U3322 (N_3322,N_2578,N_2349);
nor U3323 (N_3323,N_2694,N_295);
nor U3324 (N_3324,N_2037,N_1872);
nand U3325 (N_3325,N_2249,N_466);
or U3326 (N_3326,N_1261,N_359);
nand U3327 (N_3327,N_1102,N_1058);
nand U3328 (N_3328,N_2523,N_1310);
or U3329 (N_3329,N_2254,N_2156);
nand U3330 (N_3330,N_2522,N_2291);
nor U3331 (N_3331,N_1371,N_2800);
xor U3332 (N_3332,N_2790,N_2720);
xnor U3333 (N_3333,N_1821,N_2813);
nor U3334 (N_3334,N_2987,N_2613);
xor U3335 (N_3335,N_1059,N_736);
nand U3336 (N_3336,N_791,N_1112);
xnor U3337 (N_3337,N_426,N_93);
or U3338 (N_3338,N_1281,N_651);
nand U3339 (N_3339,N_890,N_2929);
and U3340 (N_3340,N_2273,N_289);
nand U3341 (N_3341,N_344,N_951);
nand U3342 (N_3342,N_1638,N_2574);
xor U3343 (N_3343,N_1259,N_931);
and U3344 (N_3344,N_504,N_1615);
nand U3345 (N_3345,N_1983,N_1583);
and U3346 (N_3346,N_2381,N_2967);
xnor U3347 (N_3347,N_1778,N_2185);
nand U3348 (N_3348,N_1515,N_2279);
or U3349 (N_3349,N_157,N_528);
nand U3350 (N_3350,N_1131,N_2098);
nand U3351 (N_3351,N_164,N_1999);
and U3352 (N_3352,N_1944,N_113);
nand U3353 (N_3353,N_982,N_2924);
nand U3354 (N_3354,N_575,N_1686);
nand U3355 (N_3355,N_2906,N_387);
or U3356 (N_3356,N_2262,N_1734);
and U3357 (N_3357,N_1974,N_376);
nor U3358 (N_3358,N_2544,N_550);
nor U3359 (N_3359,N_770,N_2062);
and U3360 (N_3360,N_278,N_747);
nor U3361 (N_3361,N_1658,N_1237);
or U3362 (N_3362,N_2088,N_1837);
nor U3363 (N_3363,N_1854,N_2781);
nand U3364 (N_3364,N_10,N_1126);
and U3365 (N_3365,N_1829,N_2061);
and U3366 (N_3366,N_2832,N_471);
nor U3367 (N_3367,N_1006,N_2165);
xnor U3368 (N_3368,N_1781,N_1597);
nand U3369 (N_3369,N_2359,N_1273);
nand U3370 (N_3370,N_2556,N_2109);
xnor U3371 (N_3371,N_76,N_1187);
nor U3372 (N_3372,N_2433,N_546);
or U3373 (N_3373,N_2440,N_1970);
nor U3374 (N_3374,N_858,N_1412);
nor U3375 (N_3375,N_2683,N_2508);
and U3376 (N_3376,N_739,N_55);
nand U3377 (N_3377,N_318,N_274);
or U3378 (N_3378,N_2823,N_1605);
and U3379 (N_3379,N_495,N_1205);
or U3380 (N_3380,N_1521,N_940);
nand U3381 (N_3381,N_1619,N_40);
nor U3382 (N_3382,N_914,N_2399);
nand U3383 (N_3383,N_2903,N_1216);
or U3384 (N_3384,N_1522,N_1334);
nand U3385 (N_3385,N_2581,N_2499);
or U3386 (N_3386,N_2620,N_2396);
nand U3387 (N_3387,N_2451,N_1739);
nand U3388 (N_3388,N_1793,N_1611);
nor U3389 (N_3389,N_548,N_305);
nand U3390 (N_3390,N_2728,N_1869);
and U3391 (N_3391,N_79,N_2018);
and U3392 (N_3392,N_1790,N_200);
nor U3393 (N_3393,N_122,N_1288);
nand U3394 (N_3394,N_1773,N_1218);
nand U3395 (N_3395,N_35,N_1326);
and U3396 (N_3396,N_2945,N_1717);
nand U3397 (N_3397,N_502,N_2362);
and U3398 (N_3398,N_13,N_31);
and U3399 (N_3399,N_3,N_566);
or U3400 (N_3400,N_1004,N_886);
nand U3401 (N_3401,N_2199,N_771);
or U3402 (N_3402,N_2208,N_1231);
or U3403 (N_3403,N_2347,N_2397);
nor U3404 (N_3404,N_1098,N_353);
nand U3405 (N_3405,N_1040,N_1161);
nor U3406 (N_3406,N_227,N_1298);
nand U3407 (N_3407,N_2285,N_1381);
or U3408 (N_3408,N_2435,N_2106);
nor U3409 (N_3409,N_168,N_980);
xnor U3410 (N_3410,N_2983,N_2384);
or U3411 (N_3411,N_517,N_1654);
nor U3412 (N_3412,N_1548,N_184);
nor U3413 (N_3413,N_1095,N_1804);
or U3414 (N_3414,N_1179,N_2398);
xor U3415 (N_3415,N_722,N_49);
or U3416 (N_3416,N_1062,N_1357);
nor U3417 (N_3417,N_131,N_1939);
and U3418 (N_3418,N_1951,N_1279);
nor U3419 (N_3419,N_2425,N_328);
and U3420 (N_3420,N_625,N_1254);
and U3421 (N_3421,N_1223,N_58);
nand U3422 (N_3422,N_1751,N_2794);
nor U3423 (N_3423,N_2772,N_902);
nand U3424 (N_3424,N_2422,N_2839);
nor U3425 (N_3425,N_1196,N_2639);
nor U3426 (N_3426,N_1912,N_2290);
nand U3427 (N_3427,N_660,N_2180);
nand U3428 (N_3428,N_2338,N_1346);
xor U3429 (N_3429,N_242,N_282);
and U3430 (N_3430,N_2272,N_1512);
or U3431 (N_3431,N_1285,N_405);
xnor U3432 (N_3432,N_2552,N_1700);
or U3433 (N_3433,N_2073,N_1244);
xnor U3434 (N_3434,N_1185,N_1173);
or U3435 (N_3435,N_1620,N_2575);
and U3436 (N_3436,N_2688,N_2566);
or U3437 (N_3437,N_267,N_1991);
or U3438 (N_3438,N_1073,N_1588);
xnor U3439 (N_3439,N_920,N_2178);
nor U3440 (N_3440,N_1943,N_2241);
or U3441 (N_3441,N_66,N_2123);
nand U3442 (N_3442,N_1020,N_1501);
or U3443 (N_3443,N_647,N_41);
xnor U3444 (N_3444,N_37,N_1030);
nand U3445 (N_3445,N_830,N_1438);
nand U3446 (N_3446,N_1764,N_137);
nor U3447 (N_3447,N_2989,N_1561);
and U3448 (N_3448,N_643,N_2486);
or U3449 (N_3449,N_2920,N_2911);
nor U3450 (N_3450,N_2871,N_2402);
and U3451 (N_3451,N_494,N_661);
and U3452 (N_3452,N_873,N_706);
or U3453 (N_3453,N_2799,N_1496);
nor U3454 (N_3454,N_483,N_2657);
nor U3455 (N_3455,N_2427,N_1945);
and U3456 (N_3456,N_1823,N_1962);
and U3457 (N_3457,N_1562,N_1125);
xnor U3458 (N_3458,N_255,N_1887);
xor U3459 (N_3459,N_2604,N_2938);
or U3460 (N_3460,N_1551,N_1524);
nor U3461 (N_3461,N_1743,N_509);
or U3462 (N_3462,N_1057,N_2943);
and U3463 (N_3463,N_188,N_1466);
or U3464 (N_3464,N_2751,N_68);
nand U3465 (N_3465,N_2762,N_26);
xor U3466 (N_3466,N_2841,N_1566);
nand U3467 (N_3467,N_663,N_1146);
nor U3468 (N_3468,N_1390,N_2853);
or U3469 (N_3469,N_1971,N_978);
nor U3470 (N_3470,N_1432,N_680);
nand U3471 (N_3471,N_2148,N_2815);
and U3472 (N_3472,N_2460,N_2954);
and U3473 (N_3473,N_2617,N_635);
xnor U3474 (N_3474,N_1209,N_2136);
and U3475 (N_3475,N_2450,N_321);
or U3476 (N_3476,N_2047,N_194);
and U3477 (N_3477,N_1184,N_1297);
nor U3478 (N_3478,N_2905,N_2417);
nor U3479 (N_3479,N_2108,N_848);
nor U3480 (N_3480,N_2341,N_598);
or U3481 (N_3481,N_1155,N_1877);
nand U3482 (N_3482,N_2226,N_2210);
and U3483 (N_3483,N_339,N_2172);
and U3484 (N_3484,N_603,N_406);
nor U3485 (N_3485,N_541,N_2764);
nor U3486 (N_3486,N_2335,N_683);
or U3487 (N_3487,N_958,N_1650);
nor U3488 (N_3488,N_2492,N_571);
and U3489 (N_3489,N_1094,N_2252);
or U3490 (N_3490,N_2198,N_476);
nand U3491 (N_3491,N_1493,N_2534);
or U3492 (N_3492,N_1627,N_134);
and U3493 (N_3493,N_1296,N_283);
nor U3494 (N_3494,N_2850,N_2942);
xor U3495 (N_3495,N_2782,N_2946);
nor U3496 (N_3496,N_192,N_269);
nand U3497 (N_3497,N_1109,N_1219);
nand U3498 (N_3498,N_1111,N_642);
nand U3499 (N_3499,N_667,N_2155);
nor U3500 (N_3500,N_524,N_244);
nand U3501 (N_3501,N_444,N_1665);
or U3502 (N_3502,N_2027,N_1661);
nor U3503 (N_3503,N_2961,N_1210);
or U3504 (N_3504,N_2802,N_2695);
and U3505 (N_3505,N_433,N_2101);
and U3506 (N_3506,N_2546,N_320);
nand U3507 (N_3507,N_1898,N_556);
nand U3508 (N_3508,N_1735,N_767);
nand U3509 (N_3509,N_2393,N_1256);
or U3510 (N_3510,N_2662,N_424);
nor U3511 (N_3511,N_1533,N_2641);
nand U3512 (N_3512,N_811,N_2527);
or U3513 (N_3513,N_1748,N_766);
xor U3514 (N_3514,N_1135,N_1207);
or U3515 (N_3515,N_2111,N_1653);
nand U3516 (N_3516,N_2315,N_932);
nor U3517 (N_3517,N_2937,N_1578);
or U3518 (N_3518,N_1888,N_1488);
nor U3519 (N_3519,N_702,N_1315);
nor U3520 (N_3520,N_404,N_304);
and U3521 (N_3521,N_781,N_847);
nand U3522 (N_3522,N_1459,N_748);
xnor U3523 (N_3523,N_518,N_2570);
xor U3524 (N_3524,N_2735,N_59);
nand U3525 (N_3525,N_1903,N_293);
or U3526 (N_3526,N_2126,N_266);
nand U3527 (N_3527,N_871,N_1988);
nor U3528 (N_3528,N_2763,N_50);
nor U3529 (N_3529,N_1349,N_161);
nor U3530 (N_3530,N_1956,N_2756);
nand U3531 (N_3531,N_2224,N_2182);
nand U3532 (N_3532,N_11,N_1206);
nand U3533 (N_3533,N_2994,N_128);
xor U3534 (N_3534,N_970,N_538);
xor U3535 (N_3535,N_411,N_587);
or U3536 (N_3536,N_162,N_1629);
nor U3537 (N_3537,N_2227,N_1363);
or U3538 (N_3538,N_1142,N_2158);
nor U3539 (N_3539,N_1431,N_2242);
and U3540 (N_3540,N_1042,N_468);
and U3541 (N_3541,N_1824,N_1091);
nor U3542 (N_3542,N_398,N_2538);
and U3543 (N_3543,N_792,N_1263);
nand U3544 (N_3544,N_182,N_619);
or U3545 (N_3545,N_189,N_2292);
and U3546 (N_3546,N_1399,N_208);
or U3547 (N_3547,N_2672,N_534);
and U3548 (N_3548,N_1882,N_138);
nand U3549 (N_3549,N_2328,N_1239);
nor U3550 (N_3550,N_659,N_1730);
nor U3551 (N_3551,N_2562,N_947);
and U3552 (N_3552,N_1421,N_467);
and U3553 (N_3553,N_2493,N_2130);
nor U3554 (N_3554,N_1513,N_2207);
and U3555 (N_3555,N_501,N_1189);
nand U3556 (N_3556,N_2112,N_1996);
nand U3557 (N_3557,N_300,N_2360);
xor U3558 (N_3558,N_1516,N_1737);
or U3559 (N_3559,N_2015,N_2167);
nand U3560 (N_3560,N_1132,N_1382);
nor U3561 (N_3561,N_370,N_749);
nand U3562 (N_3562,N_510,N_2645);
and U3563 (N_3563,N_582,N_1755);
and U3564 (N_3564,N_637,N_268);
or U3565 (N_3565,N_2869,N_2115);
or U3566 (N_3566,N_516,N_1105);
and U3567 (N_3567,N_768,N_2430);
nand U3568 (N_3568,N_2528,N_927);
or U3569 (N_3569,N_2052,N_1352);
xor U3570 (N_3570,N_2134,N_1269);
nand U3571 (N_3571,N_2471,N_1457);
nand U3572 (N_3572,N_733,N_290);
or U3573 (N_3573,N_1014,N_797);
xnor U3574 (N_3574,N_2927,N_1164);
nor U3575 (N_3575,N_2375,N_1801);
nor U3576 (N_3576,N_485,N_2599);
or U3577 (N_3577,N_1531,N_1586);
or U3578 (N_3578,N_793,N_2202);
or U3579 (N_3579,N_2255,N_2);
xnor U3580 (N_3580,N_809,N_1257);
nand U3581 (N_3581,N_1645,N_2899);
or U3582 (N_3582,N_1379,N_1973);
nand U3583 (N_3583,N_1998,N_460);
nor U3584 (N_3584,N_458,N_1079);
nor U3585 (N_3585,N_2007,N_2821);
and U3586 (N_3586,N_1733,N_2020);
nor U3587 (N_3587,N_933,N_1902);
nor U3588 (N_3588,N_1707,N_1663);
nand U3589 (N_3589,N_2689,N_2459);
or U3590 (N_3590,N_478,N_1087);
and U3591 (N_3591,N_1405,N_250);
or U3592 (N_3592,N_417,N_252);
or U3593 (N_3593,N_2737,N_2313);
and U3594 (N_3594,N_1433,N_780);
and U3595 (N_3595,N_1849,N_1194);
xnor U3596 (N_3596,N_2096,N_2298);
nand U3597 (N_3597,N_570,N_2056);
xnor U3598 (N_3598,N_1479,N_1019);
or U3599 (N_3599,N_1160,N_2690);
nand U3600 (N_3600,N_665,N_2441);
nor U3601 (N_3601,N_1766,N_677);
or U3602 (N_3602,N_1815,N_2969);
or U3603 (N_3603,N_2530,N_764);
nor U3604 (N_3604,N_1926,N_1651);
nor U3605 (N_3605,N_1746,N_2122);
and U3606 (N_3606,N_1319,N_1783);
xnor U3607 (N_3607,N_1168,N_2656);
nand U3608 (N_3608,N_2633,N_1626);
or U3609 (N_3609,N_65,N_500);
and U3610 (N_3610,N_2186,N_2069);
nand U3611 (N_3611,N_377,N_2885);
or U3612 (N_3612,N_784,N_1814);
or U3613 (N_3613,N_1770,N_977);
and U3614 (N_3614,N_2976,N_1836);
nor U3615 (N_3615,N_1471,N_312);
and U3616 (N_3616,N_1550,N_1241);
and U3617 (N_3617,N_2734,N_2383);
and U3618 (N_3618,N_714,N_1074);
xor U3619 (N_3619,N_574,N_1434);
and U3620 (N_3620,N_2344,N_662);
or U3621 (N_3621,N_990,N_1706);
xor U3622 (N_3622,N_32,N_1776);
nor U3623 (N_3623,N_2959,N_118);
and U3624 (N_3624,N_308,N_2892);
nand U3625 (N_3625,N_241,N_1046);
nand U3626 (N_3626,N_2846,N_2124);
nand U3627 (N_3627,N_2622,N_2874);
xor U3628 (N_3628,N_2808,N_2234);
and U3629 (N_3629,N_1557,N_203);
nor U3630 (N_3630,N_612,N_2761);
or U3631 (N_3631,N_2065,N_1139);
nand U3632 (N_3632,N_2548,N_2679);
or U3633 (N_3633,N_2391,N_2275);
and U3634 (N_3634,N_2812,N_1482);
or U3635 (N_3635,N_2316,N_1564);
nand U3636 (N_3636,N_2706,N_381);
xnor U3637 (N_3637,N_2204,N_2944);
and U3638 (N_3638,N_2423,N_2563);
nand U3639 (N_3639,N_1152,N_754);
or U3640 (N_3640,N_2834,N_1692);
and U3641 (N_3641,N_2283,N_2248);
and U3642 (N_3642,N_1047,N_823);
or U3643 (N_3643,N_2909,N_669);
nor U3644 (N_3644,N_1810,N_2553);
nand U3645 (N_3645,N_1676,N_394);
and U3646 (N_3646,N_2718,N_705);
nand U3647 (N_3647,N_452,N_2428);
or U3648 (N_3648,N_2237,N_2269);
or U3649 (N_3649,N_1563,N_2076);
and U3650 (N_3650,N_2378,N_1690);
nor U3651 (N_3651,N_2184,N_1517);
and U3652 (N_3652,N_2873,N_586);
nand U3653 (N_3653,N_2932,N_2801);
or U3654 (N_3654,N_323,N_2950);
or U3655 (N_3655,N_2984,N_2935);
xor U3656 (N_3656,N_592,N_197);
or U3657 (N_3657,N_2002,N_2502);
or U3658 (N_3658,N_1485,N_557);
or U3659 (N_3659,N_1857,N_639);
xnor U3660 (N_3660,N_1022,N_966);
and U3661 (N_3661,N_2537,N_14);
or U3662 (N_3662,N_2503,N_27);
nor U3663 (N_3663,N_1948,N_296);
or U3664 (N_3664,N_568,N_492);
nor U3665 (N_3665,N_284,N_1897);
nand U3666 (N_3666,N_2281,N_461);
or U3667 (N_3667,N_100,N_1116);
nand U3668 (N_3668,N_2094,N_119);
and U3669 (N_3669,N_1884,N_455);
or U3670 (N_3670,N_684,N_2867);
nor U3671 (N_3671,N_1267,N_2300);
and U3672 (N_3672,N_1969,N_1612);
or U3673 (N_3673,N_2082,N_2887);
and U3674 (N_3674,N_2806,N_331);
or U3675 (N_3675,N_463,N_2826);
or U3676 (N_3676,N_803,N_259);
and U3677 (N_3677,N_20,N_1572);
and U3678 (N_3678,N_1698,N_576);
xor U3679 (N_3679,N_1243,N_2452);
or U3680 (N_3680,N_1848,N_102);
nand U3681 (N_3681,N_2973,N_2529);
or U3682 (N_3682,N_2624,N_450);
or U3683 (N_3683,N_1908,N_810);
nor U3684 (N_3684,N_2787,N_117);
and U3685 (N_3685,N_481,N_1163);
nor U3686 (N_3686,N_807,N_991);
or U3687 (N_3687,N_2271,N_505);
nand U3688 (N_3688,N_445,N_1);
xor U3689 (N_3689,N_833,N_1922);
nor U3690 (N_3690,N_2844,N_1053);
xnor U3691 (N_3691,N_1741,N_2931);
nor U3692 (N_3692,N_1747,N_439);
and U3693 (N_3693,N_879,N_2692);
or U3694 (N_3694,N_542,N_712);
nor U3695 (N_3695,N_1224,N_1145);
or U3696 (N_3696,N_1762,N_2740);
and U3697 (N_3697,N_159,N_521);
nand U3698 (N_3698,N_2203,N_2727);
or U3699 (N_3699,N_919,N_2631);
nand U3700 (N_3700,N_209,N_700);
nand U3701 (N_3701,N_388,N_580);
or U3702 (N_3702,N_2982,N_1555);
nor U3703 (N_3703,N_317,N_2260);
and U3704 (N_3704,N_2205,N_2745);
and U3705 (N_3705,N_2191,N_999);
xnor U3706 (N_3706,N_1321,N_2238);
nor U3707 (N_3707,N_2779,N_2947);
and U3708 (N_3708,N_2667,N_607);
or U3709 (N_3709,N_2053,N_2223);
and U3710 (N_3710,N_87,N_903);
or U3711 (N_3711,N_1075,N_465);
or U3712 (N_3712,N_1464,N_1753);
or U3713 (N_3713,N_1486,N_89);
nand U3714 (N_3714,N_302,N_2837);
nand U3715 (N_3715,N_54,N_2749);
or U3716 (N_3716,N_2699,N_2259);
nand U3717 (N_3717,N_401,N_2280);
nor U3718 (N_3718,N_183,N_1909);
nand U3719 (N_3719,N_1029,N_1656);
nor U3720 (N_3720,N_1016,N_563);
and U3721 (N_3721,N_90,N_2721);
nand U3722 (N_3722,N_2371,N_2589);
xor U3723 (N_3723,N_1311,N_179);
or U3724 (N_3724,N_349,N_622);
and U3725 (N_3725,N_2614,N_696);
nand U3726 (N_3726,N_1820,N_1191);
or U3727 (N_3727,N_2852,N_1043);
xnor U3728 (N_3728,N_2032,N_23);
nor U3729 (N_3729,N_422,N_2580);
nor U3730 (N_3730,N_2559,N_2392);
or U3731 (N_3731,N_1251,N_2067);
nor U3732 (N_3732,N_2505,N_1156);
nor U3733 (N_3733,N_176,N_1875);
and U3734 (N_3734,N_1918,N_1389);
or U3735 (N_3735,N_2588,N_1108);
and U3736 (N_3736,N_822,N_2309);
nand U3737 (N_3737,N_457,N_2977);
nor U3738 (N_3738,N_1738,N_2193);
and U3739 (N_3739,N_1294,N_1475);
nor U3740 (N_3740,N_148,N_2390);
or U3741 (N_3741,N_326,N_83);
and U3742 (N_3742,N_2453,N_6);
and U3743 (N_3743,N_1450,N_992);
nand U3744 (N_3744,N_2016,N_1414);
nor U3745 (N_3745,N_955,N_549);
and U3746 (N_3746,N_1000,N_2395);
xnor U3747 (N_3747,N_887,N_2475);
or U3748 (N_3748,N_2840,N_1881);
xnor U3749 (N_3749,N_2619,N_1265);
or U3750 (N_3750,N_1264,N_2467);
nor U3751 (N_3751,N_1808,N_1929);
or U3752 (N_3752,N_795,N_351);
nand U3753 (N_3753,N_1589,N_1201);
nor U3754 (N_3754,N_2642,N_1543);
nand U3755 (N_3755,N_1289,N_297);
and U3756 (N_3756,N_153,N_1777);
nand U3757 (N_3757,N_975,N_2682);
xor U3758 (N_3758,N_915,N_2095);
nor U3759 (N_3759,N_1575,N_1331);
nand U3760 (N_3760,N_1299,N_174);
nand U3761 (N_3761,N_491,N_1356);
and U3762 (N_3762,N_552,N_2608);
nand U3763 (N_3763,N_2267,N_826);
or U3764 (N_3764,N_2986,N_1775);
nor U3765 (N_3765,N_2501,N_832);
nor U3766 (N_3766,N_1008,N_2539);
or U3767 (N_3767,N_447,N_685);
xnor U3768 (N_3768,N_898,N_152);
and U3769 (N_3769,N_850,N_2814);
xor U3770 (N_3770,N_1697,N_649);
xor U3771 (N_3771,N_2000,N_2050);
nor U3772 (N_3772,N_652,N_2894);
nand U3773 (N_3773,N_9,N_1695);
nor U3774 (N_3774,N_1124,N_913);
nand U3775 (N_3775,N_1606,N_1532);
and U3776 (N_3776,N_39,N_279);
nand U3777 (N_3777,N_1644,N_1978);
xnor U3778 (N_3778,N_2702,N_802);
nand U3779 (N_3779,N_2200,N_121);
and U3780 (N_3780,N_1307,N_1660);
or U3781 (N_3781,N_2507,N_655);
nand U3782 (N_3782,N_2804,N_930);
nor U3783 (N_3783,N_235,N_1934);
or U3784 (N_3784,N_1012,N_1477);
nand U3785 (N_3785,N_1616,N_146);
and U3786 (N_3786,N_2461,N_2369);
nand U3787 (N_3787,N_1128,N_2322);
and U3788 (N_3788,N_2817,N_1468);
xnor U3789 (N_3789,N_2582,N_883);
nor U3790 (N_3790,N_127,N_1980);
and U3791 (N_3791,N_1731,N_2912);
nand U3792 (N_3792,N_682,N_2141);
nor U3793 (N_3793,N_434,N_307);
xor U3794 (N_3794,N_46,N_882);
xnor U3795 (N_3795,N_1048,N_908);
and U3796 (N_3796,N_294,N_1300);
and U3797 (N_3797,N_2083,N_994);
and U3798 (N_3798,N_2859,N_1866);
and U3799 (N_3799,N_210,N_2444);
or U3800 (N_3800,N_18,N_1435);
nand U3801 (N_3801,N_1323,N_2303);
or U3802 (N_3802,N_613,N_690);
nand U3803 (N_3803,N_1503,N_985);
xor U3804 (N_3804,N_1500,N_213);
nand U3805 (N_3805,N_2128,N_1826);
nand U3806 (N_3806,N_261,N_2306);
and U3807 (N_3807,N_1286,N_2087);
and U3808 (N_3808,N_1386,N_1809);
and U3809 (N_3809,N_1472,N_2535);
or U3810 (N_3810,N_1649,N_2263);
nand U3811 (N_3811,N_61,N_849);
nor U3812 (N_3812,N_248,N_859);
nand U3813 (N_3813,N_1467,N_12);
and U3814 (N_3814,N_2611,N_324);
or U3815 (N_3815,N_2099,N_2660);
or U3816 (N_3816,N_2177,N_1920);
xnor U3817 (N_3817,N_2605,N_368);
nand U3818 (N_3818,N_618,N_299);
or U3819 (N_3819,N_2127,N_732);
or U3820 (N_3820,N_2287,N_2521);
xor U3821 (N_3821,N_2992,N_2414);
or U3822 (N_3822,N_2437,N_820);
nor U3823 (N_3823,N_2980,N_1084);
or U3824 (N_3824,N_1587,N_160);
nor U3825 (N_3825,N_1214,N_892);
nor U3826 (N_3826,N_1915,N_2621);
nor U3827 (N_3827,N_2187,N_1229);
or U3828 (N_3828,N_1933,N_2698);
and U3829 (N_3829,N_2669,N_1805);
or U3830 (N_3830,N_877,N_726);
or U3831 (N_3831,N_2648,N_2602);
xnor U3832 (N_3832,N_2090,N_503);
and U3833 (N_3833,N_2540,N_1582);
nand U3834 (N_3834,N_1143,N_335);
nand U3835 (N_3835,N_876,N_2310);
and U3836 (N_3836,N_1745,N_2549);
or U3837 (N_3837,N_139,N_846);
and U3838 (N_3838,N_1919,N_2035);
nand U3839 (N_3839,N_1835,N_1121);
or U3840 (N_3840,N_1417,N_379);
nand U3841 (N_3841,N_313,N_2791);
and U3842 (N_3842,N_2215,N_553);
and U3843 (N_3843,N_350,N_2373);
nor U3844 (N_3844,N_532,N_2028);
or U3845 (N_3845,N_1784,N_2836);
or U3846 (N_3846,N_1504,N_421);
or U3847 (N_3847,N_2573,N_2600);
xnor U3848 (N_3848,N_755,N_2675);
or U3849 (N_3849,N_2077,N_551);
nor U3850 (N_3850,N_2531,N_1342);
and U3851 (N_3851,N_1470,N_354);
nor U3852 (N_3852,N_2006,N_2968);
or U3853 (N_3853,N_2997,N_1343);
and U3854 (N_3854,N_645,N_2716);
nand U3855 (N_3855,N_973,N_1258);
or U3856 (N_3856,N_2377,N_2649);
xnor U3857 (N_3857,N_2054,N_2350);
nor U3858 (N_3858,N_614,N_1400);
nand U3859 (N_3859,N_976,N_1233);
and U3860 (N_3860,N_477,N_1117);
or U3861 (N_3861,N_1941,N_1480);
and U3862 (N_3862,N_2551,N_2413);
and U3863 (N_3863,N_2849,N_2818);
or U3864 (N_3864,N_2701,N_616);
nand U3865 (N_3865,N_2770,N_581);
nand U3866 (N_3866,N_644,N_1262);
nor U3867 (N_3867,N_1101,N_1542);
nor U3868 (N_3868,N_211,N_1750);
or U3869 (N_3869,N_2081,N_1701);
xor U3870 (N_3870,N_1249,N_774);
nor U3871 (N_3871,N_2769,N_2012);
or U3872 (N_3872,N_70,N_2634);
or U3873 (N_3873,N_2256,N_285);
nand U3874 (N_3874,N_389,N_420);
nor U3875 (N_3875,N_1672,N_864);
or U3876 (N_3876,N_1594,N_2296);
or U3877 (N_3877,N_1277,N_1689);
nand U3878 (N_3878,N_4,N_1576);
nand U3879 (N_3879,N_2114,N_506);
and U3880 (N_3880,N_1679,N_812);
and U3881 (N_3881,N_2919,N_2658);
nand U3882 (N_3882,N_413,N_1069);
and U3883 (N_3883,N_1498,N_1724);
xor U3884 (N_3884,N_2213,N_1238);
nor U3885 (N_3885,N_963,N_1728);
nand U3886 (N_3886,N_595,N_1648);
nand U3887 (N_3887,N_1066,N_1362);
nand U3888 (N_3888,N_691,N_251);
nand U3889 (N_3889,N_2615,N_437);
nand U3890 (N_3890,N_1924,N_602);
nand U3891 (N_3891,N_1328,N_1415);
nand U3892 (N_3892,N_1193,N_818);
nor U3893 (N_3893,N_1916,N_843);
or U3894 (N_3894,N_838,N_2003);
nand U3895 (N_3895,N_829,N_2995);
nor U3896 (N_3896,N_1845,N_1361);
and U3897 (N_3897,N_1647,N_1792);
xnor U3898 (N_3898,N_2780,N_315);
and U3899 (N_3899,N_2816,N_1642);
xnor U3900 (N_3900,N_441,N_464);
nor U3901 (N_3901,N_15,N_2495);
nor U3902 (N_3902,N_385,N_836);
or U3903 (N_3903,N_1911,N_231);
or U3904 (N_3904,N_2673,N_611);
nor U3905 (N_3905,N_287,N_114);
nor U3906 (N_3906,N_1752,N_2933);
and U3907 (N_3907,N_474,N_2270);
nand U3908 (N_3908,N_219,N_1407);
or U3909 (N_3909,N_2021,N_741);
and U3910 (N_3910,N_240,N_801);
and U3911 (N_3911,N_361,N_484);
or U3912 (N_3912,N_1886,N_348);
and U3913 (N_3913,N_1591,N_369);
nand U3914 (N_3914,N_1921,N_2925);
or U3915 (N_3915,N_1828,N_1383);
xor U3916 (N_3916,N_1284,N_535);
nor U3917 (N_3917,N_1403,N_1422);
nor U3918 (N_3918,N_1904,N_508);
and U3919 (N_3919,N_1302,N_2348);
xnor U3920 (N_3920,N_1782,N_1172);
or U3921 (N_3921,N_1123,N_2265);
nor U3922 (N_3922,N_2864,N_765);
and U3923 (N_3923,N_2999,N_185);
or U3924 (N_3924,N_2623,N_1452);
xor U3925 (N_3925,N_1451,N_929);
and U3926 (N_3926,N_1977,N_777);
and U3927 (N_3927,N_2266,N_2710);
and U3928 (N_3928,N_2357,N_2895);
and U3929 (N_3929,N_983,N_2771);
and U3930 (N_3930,N_1799,N_2250);
nand U3931 (N_3931,N_2736,N_2643);
nor U3932 (N_3932,N_479,N_1624);
or U3933 (N_3933,N_2201,N_395);
xor U3934 (N_3934,N_2807,N_2153);
and U3935 (N_3935,N_2404,N_1613);
or U3936 (N_3936,N_2518,N_1178);
nand U3937 (N_3937,N_7,N_1350);
nand U3938 (N_3938,N_264,N_2333);
and U3939 (N_3939,N_2463,N_664);
xnor U3940 (N_3940,N_2590,N_246);
nor U3941 (N_3941,N_1553,N_1127);
or U3942 (N_3942,N_813,N_786);
and U3943 (N_3943,N_2922,N_2711);
xnor U3944 (N_3944,N_1378,N_834);
or U3945 (N_3945,N_1842,N_907);
or U3946 (N_3946,N_1843,N_2587);
or U3947 (N_3947,N_1396,N_514);
and U3948 (N_3948,N_1165,N_941);
and U3949 (N_3949,N_2120,N_2147);
nor U3950 (N_3950,N_1953,N_1537);
and U3951 (N_3951,N_2519,N_694);
and U3952 (N_3952,N_272,N_1078);
nand U3953 (N_3953,N_1761,N_2677);
xor U3954 (N_3954,N_668,N_889);
and U3955 (N_3955,N_2876,N_2557);
or U3956 (N_3956,N_1186,N_1540);
and U3957 (N_3957,N_2327,N_81);
and U3958 (N_3958,N_2697,N_1341);
and U3959 (N_3959,N_2097,N_1041);
nor U3960 (N_3960,N_2355,N_1569);
nand U3961 (N_3961,N_2616,N_2110);
nand U3962 (N_3962,N_1044,N_271);
nor U3963 (N_3963,N_2571,N_2678);
nor U3964 (N_3964,N_1304,N_2664);
xor U3965 (N_3965,N_2676,N_1684);
nand U3966 (N_3966,N_489,N_2163);
and U3967 (N_3967,N_1365,N_1505);
nand U3968 (N_3968,N_1670,N_2632);
and U3969 (N_3969,N_2717,N_1202);
or U3970 (N_3970,N_222,N_986);
xor U3971 (N_3971,N_1188,N_688);
and U3972 (N_3972,N_519,N_594);
nor U3973 (N_3973,N_2978,N_224);
xor U3974 (N_3974,N_202,N_2040);
nand U3975 (N_3975,N_1154,N_852);
or U3976 (N_3976,N_1445,N_2013);
nand U3977 (N_3977,N_1354,N_338);
and U3978 (N_3978,N_2133,N_116);
xor U3979 (N_3979,N_24,N_2387);
or U3980 (N_3980,N_2786,N_1215);
and U3981 (N_3981,N_2483,N_854);
nor U3982 (N_3982,N_794,N_2152);
and U3983 (N_3983,N_2351,N_314);
nor U3984 (N_3984,N_597,N_249);
and U3985 (N_3985,N_136,N_187);
nor U3986 (N_3986,N_2955,N_2189);
or U3987 (N_3987,N_657,N_2264);
nand U3988 (N_3988,N_1250,N_1757);
nor U3989 (N_3989,N_1552,N_2317);
xnor U3990 (N_3990,N_2070,N_2644);
nor U3991 (N_3991,N_1767,N_1702);
nor U3992 (N_3992,N_2558,N_2567);
nor U3993 (N_3993,N_345,N_1140);
nand U3994 (N_3994,N_709,N_1610);
and U3995 (N_3995,N_151,N_638);
nand U3996 (N_3996,N_1494,N_1657);
and U3997 (N_3997,N_590,N_2342);
nor U3998 (N_3998,N_362,N_710);
or U3999 (N_3999,N_1242,N_2991);
and U4000 (N_4000,N_2150,N_228);
xor U4001 (N_4001,N_2907,N_2767);
xor U4002 (N_4002,N_762,N_2768);
nor U4003 (N_4003,N_257,N_206);
xor U4004 (N_4004,N_583,N_1122);
and U4005 (N_4005,N_391,N_2022);
nor U4006 (N_4006,N_2774,N_1035);
and U4007 (N_4007,N_1255,N_1038);
and U4008 (N_4008,N_1159,N_111);
nor U4009 (N_4009,N_825,N_48);
nand U4010 (N_4010,N_745,N_104);
nor U4011 (N_4011,N_1426,N_1175);
and U4012 (N_4012,N_1986,N_288);
nor U4013 (N_4013,N_1428,N_1987);
xnor U4014 (N_4014,N_1103,N_158);
nand U4015 (N_4015,N_2478,N_934);
nor U4016 (N_4016,N_1456,N_969);
xor U4017 (N_4017,N_2100,N_1174);
and U4018 (N_4018,N_2949,N_1469);
or U4019 (N_4019,N_1742,N_432);
and U4020 (N_4020,N_1652,N_2691);
nand U4021 (N_4021,N_2374,N_1293);
nor U4022 (N_4022,N_2890,N_723);
nor U4023 (N_4023,N_773,N_149);
and U4024 (N_4024,N_2209,N_870);
nor U4025 (N_4025,N_1927,N_1398);
or U4026 (N_4026,N_1609,N_2466);
and U4027 (N_4027,N_1711,N_761);
and U4028 (N_4028,N_1579,N_1228);
or U4029 (N_4029,N_1623,N_2071);
nand U4030 (N_4030,N_291,N_91);
and U4031 (N_4031,N_1253,N_2394);
or U4032 (N_4032,N_1846,N_1632);
and U4033 (N_4033,N_2861,N_470);
xnor U4034 (N_4034,N_346,N_396);
nor U4035 (N_4035,N_2221,N_2651);
nor U4036 (N_4036,N_522,N_1153);
nand U4037 (N_4037,N_1580,N_880);
and U4038 (N_4038,N_2023,N_2085);
nand U4039 (N_4039,N_1001,N_73);
or U4040 (N_4040,N_2625,N_2473);
nand U4041 (N_4041,N_2343,N_407);
nand U4042 (N_4042,N_2411,N_2282);
nand U4043 (N_4043,N_1028,N_1222);
and U4044 (N_4044,N_2001,N_44);
and U4045 (N_4045,N_2827,N_2036);
and U4046 (N_4046,N_342,N_2793);
or U4047 (N_4047,N_1106,N_593);
nand U4048 (N_4048,N_805,N_2610);
nor U4049 (N_4049,N_954,N_806);
and U4050 (N_4050,N_2811,N_1547);
and U4051 (N_4051,N_1051,N_2513);
or U4052 (N_4052,N_425,N_2526);
or U4053 (N_4053,N_409,N_130);
xor U4054 (N_4054,N_909,N_1703);
nand U4055 (N_4055,N_2958,N_1463);
xnor U4056 (N_4056,N_841,N_674);
or U4057 (N_4057,N_2891,N_1825);
or U4058 (N_4058,N_1502,N_2299);
nor U4059 (N_4059,N_430,N_539);
nand U4060 (N_4060,N_1841,N_343);
or U4061 (N_4061,N_2400,N_2231);
nand U4062 (N_4062,N_2872,N_2681);
or U4063 (N_4063,N_874,N_2480);
nand U4064 (N_4064,N_1900,N_442);
nor U4065 (N_4065,N_2687,N_1791);
and U4066 (N_4066,N_2367,N_2055);
nand U4067 (N_4067,N_746,N_169);
or U4068 (N_4068,N_1895,N_686);
nand U4069 (N_4069,N_1086,N_1454);
nor U4070 (N_4070,N_1772,N_2703);
or U4071 (N_4071,N_456,N_1465);
or U4072 (N_4072,N_1266,N_1967);
nor U4073 (N_4073,N_1481,N_77);
nand U4074 (N_4074,N_403,N_2750);
nand U4075 (N_4075,N_1938,N_853);
nor U4076 (N_4076,N_1585,N_808);
nor U4077 (N_4077,N_617,N_1539);
nor U4078 (N_4078,N_51,N_1455);
nand U4079 (N_4079,N_2783,N_1411);
or U4080 (N_4080,N_2536,N_972);
or U4081 (N_4081,N_2157,N_2195);
nand U4082 (N_4082,N_711,N_1060);
nor U4083 (N_4083,N_230,N_303);
nand U4084 (N_4084,N_1324,N_1359);
nand U4085 (N_4085,N_2532,N_1439);
xnor U4086 (N_4086,N_2059,N_1671);
nor U4087 (N_4087,N_1935,N_1071);
and U4088 (N_4088,N_1177,N_1151);
or U4089 (N_4089,N_2166,N_2131);
and U4090 (N_4090,N_1961,N_2089);
and U4091 (N_4091,N_1930,N_1787);
and U4092 (N_4092,N_47,N_416);
and U4093 (N_4093,N_2431,N_2979);
nand U4094 (N_4094,N_1005,N_2364);
nor U4095 (N_4095,N_371,N_2135);
and U4096 (N_4096,N_630,N_2142);
or U4097 (N_4097,N_1271,N_1368);
and U4098 (N_4098,N_2543,N_1025);
and U4099 (N_4099,N_2079,N_1873);
and U4100 (N_4100,N_2132,N_1387);
nor U4101 (N_4101,N_1932,N_2151);
or U4102 (N_4102,N_1596,N_1976);
nor U4103 (N_4103,N_30,N_968);
or U4104 (N_4104,N_559,N_2668);
or U4105 (N_4105,N_1673,N_866);
nor U4106 (N_4106,N_1290,N_719);
and U4107 (N_4107,N_2659,N_367);
or U4108 (N_4108,N_1002,N_2026);
and U4109 (N_4109,N_987,N_1816);
nand U4110 (N_4110,N_787,N_2312);
nand U4111 (N_4111,N_120,N_1148);
or U4112 (N_4112,N_2324,N_380);
nand U4113 (N_4113,N_653,N_1883);
or U4114 (N_4114,N_1960,N_1473);
nand U4115 (N_4115,N_1308,N_821);
nor U4116 (N_4116,N_2380,N_2565);
nand U4117 (N_4117,N_2038,N_69);
nand U4118 (N_4118,N_782,N_1822);
nand U4119 (N_4119,N_2379,N_891);
xnor U4120 (N_4120,N_410,N_2320);
nor U4121 (N_4121,N_319,N_378);
and U4122 (N_4122,N_2041,N_779);
nor U4123 (N_4123,N_1444,N_2862);
xnor U4124 (N_4124,N_220,N_2766);
nand U4125 (N_4125,N_626,N_1722);
nor U4126 (N_4126,N_2635,N_8);
nand U4127 (N_4127,N_2169,N_2825);
nand U4128 (N_4128,N_1862,N_1138);
nor U4129 (N_4129,N_1839,N_2258);
nor U4130 (N_4130,N_2500,N_178);
nor U4131 (N_4131,N_1518,N_918);
and U4132 (N_4132,N_1840,N_2754);
or U4133 (N_4133,N_1779,N_1373);
xor U4134 (N_4134,N_2630,N_1844);
and U4135 (N_4135,N_656,N_372);
or U4136 (N_4136,N_911,N_2857);
nand U4137 (N_4137,N_1899,N_815);
nor U4138 (N_4138,N_198,N_1130);
xor U4139 (N_4139,N_1437,N_2882);
nand U4140 (N_4140,N_917,N_462);
nand U4141 (N_4141,N_1089,N_1800);
nand U4142 (N_4142,N_1819,N_2964);
nor U4143 (N_4143,N_2579,N_888);
and U4144 (N_4144,N_2043,N_731);
xor U4145 (N_4145,N_2858,N_1599);
or U4146 (N_4146,N_904,N_636);
xnor U4147 (N_4147,N_964,N_99);
xor U4148 (N_4148,N_1714,N_1424);
nand U4149 (N_4149,N_2154,N_186);
nand U4150 (N_4150,N_2321,N_2773);
nand U4151 (N_4151,N_1100,N_1788);
or U4152 (N_4152,N_544,N_627);
nor U4153 (N_4153,N_1446,N_2524);
and U4154 (N_4154,N_624,N_472);
nand U4155 (N_4155,N_2928,N_2336);
nor U4156 (N_4156,N_254,N_2926);
nand U4157 (N_4157,N_2510,N_386);
xor U4158 (N_4158,N_744,N_60);
nor U4159 (N_4159,N_1527,N_1270);
xor U4160 (N_4160,N_2304,N_1203);
nor U4161 (N_4161,N_337,N_2758);
nand U4162 (N_4162,N_1003,N_1442);
or U4163 (N_4163,N_1134,N_1720);
nand U4164 (N_4164,N_1309,N_205);
nor U4165 (N_4165,N_2330,N_606);
and U4166 (N_4166,N_2319,N_233);
or U4167 (N_4167,N_1774,N_1448);
nand U4168 (N_4168,N_740,N_1688);
and U4169 (N_4169,N_2366,N_482);
nor U4170 (N_4170,N_621,N_232);
and U4171 (N_4171,N_374,N_695);
and U4172 (N_4172,N_1833,N_1710);
xnor U4173 (N_4173,N_1147,N_2671);
nor U4174 (N_4174,N_2093,N_981);
nand U4175 (N_4175,N_1995,N_218);
nor U4176 (N_4176,N_536,N_1910);
and U4177 (N_4177,N_2245,N_2401);
nor U4178 (N_4178,N_974,N_1817);
nand U4179 (N_4179,N_1507,N_1992);
and U4180 (N_4180,N_156,N_2010);
nor U4181 (N_4181,N_2586,N_1487);
or U4182 (N_4182,N_2948,N_115);
nand U4183 (N_4183,N_496,N_1593);
nor U4184 (N_4184,N_2514,N_1985);
nand U4185 (N_4185,N_1853,N_2972);
or U4186 (N_4186,N_400,N_737);
nor U4187 (N_4187,N_276,N_2446);
or U4188 (N_4188,N_837,N_1478);
nor U4189 (N_4189,N_2798,N_2286);
xnor U4190 (N_4190,N_1631,N_2173);
nand U4191 (N_4191,N_601,N_177);
nor U4192 (N_4192,N_1458,N_459);
nand U4193 (N_4193,N_1474,N_2214);
or U4194 (N_4194,N_310,N_1385);
nor U4195 (N_4195,N_1890,N_2368);
and U4196 (N_4196,N_1641,N_1180);
or U4197 (N_4197,N_72,N_1713);
or U4198 (N_4198,N_1376,N_216);
and U4199 (N_4199,N_1374,N_641);
nand U4200 (N_4200,N_2960,N_1072);
nor U4201 (N_4201,N_1204,N_2457);
or U4202 (N_4202,N_2957,N_480);
or U4203 (N_4203,N_217,N_129);
nor U4204 (N_4204,N_861,N_703);
nand U4205 (N_4205,N_924,N_1092);
nand U4206 (N_4206,N_790,N_1335);
and U4207 (N_4207,N_671,N_336);
nor U4208 (N_4208,N_2372,N_78);
nand U4209 (N_4209,N_1192,N_2722);
nor U4210 (N_4210,N_2340,N_2830);
nand U4211 (N_4211,N_1182,N_365);
and U4212 (N_4212,N_2468,N_2318);
or U4213 (N_4213,N_1509,N_2489);
or U4214 (N_4214,N_2294,N_1874);
nand U4215 (N_4215,N_486,N_1955);
nand U4216 (N_4216,N_1492,N_648);
nand U4217 (N_4217,N_2917,N_800);
xor U4218 (N_4218,N_1113,N_2576);
and U4219 (N_4219,N_1602,N_1282);
or U4220 (N_4220,N_88,N_2479);
nor U4221 (N_4221,N_1622,N_1360);
and U4222 (N_4222,N_2447,N_2476);
nor U4223 (N_4223,N_2219,N_555);
nor U4224 (N_4224,N_1694,N_1033);
and U4225 (N_4225,N_2739,N_1015);
or U4226 (N_4226,N_1968,N_1026);
and U4227 (N_4227,N_1305,N_2346);
and U4228 (N_4228,N_397,N_1952);
or U4229 (N_4229,N_166,N_330);
and U4230 (N_4230,N_2448,N_1325);
nor U4231 (N_4231,N_1461,N_165);
or U4232 (N_4232,N_530,N_171);
and U4233 (N_4233,N_1940,N_998);
nand U4234 (N_4234,N_728,N_1427);
nand U4235 (N_4235,N_679,N_2365);
or U4236 (N_4236,N_1260,N_1077);
and U4237 (N_4237,N_631,N_2753);
and U4238 (N_4238,N_2140,N_1489);
and U4239 (N_4239,N_2881,N_1530);
or U4240 (N_4240,N_2048,N_1090);
nor U4241 (N_4241,N_1954,N_1659);
nor U4242 (N_4242,N_1677,N_2638);
nor U4243 (N_4243,N_673,N_896);
and U4244 (N_4244,N_347,N_1574);
xor U4245 (N_4245,N_842,N_936);
or U4246 (N_4246,N_816,N_1337);
or U4247 (N_4247,N_2731,N_599);
nand U4248 (N_4248,N_2785,N_418);
xnor U4249 (N_4249,N_43,N_190);
and U4250 (N_4250,N_2314,N_1957);
or U4251 (N_4251,N_1021,N_2419);
nor U4252 (N_4252,N_2888,N_449);
nand U4253 (N_4253,N_1375,N_1447);
nand U4254 (N_4254,N_1538,N_1476);
nor U4255 (N_4255,N_1508,N_1568);
nor U4256 (N_4256,N_610,N_427);
and U4257 (N_4257,N_1056,N_1721);
nand U4258 (N_4258,N_750,N_2854);
nor U4259 (N_4259,N_1525,N_2192);
nor U4260 (N_4260,N_135,N_1558);
or U4261 (N_4261,N_2332,N_957);
nand U4262 (N_4262,N_1607,N_0);
and U4263 (N_4263,N_2653,N_2149);
and U4264 (N_4264,N_1867,N_363);
nand U4265 (N_4265,N_2971,N_1989);
nor U4266 (N_4266,N_912,N_360);
nor U4267 (N_4267,N_1878,N_2618);
or U4268 (N_4268,N_1754,N_2775);
or U4269 (N_4269,N_1965,N_2686);
nand U4270 (N_4270,N_2225,N_2469);
or U4271 (N_4271,N_1067,N_1685);
or U4272 (N_4272,N_693,N_1010);
or U4273 (N_4273,N_2810,N_1213);
or U4274 (N_4274,N_2700,N_1149);
nand U4275 (N_4275,N_899,N_2865);
nor U4276 (N_4276,N_1410,N_1674);
xor U4277 (N_4277,N_1885,N_716);
nor U4278 (N_4278,N_1333,N_2746);
nand U4279 (N_4279,N_2725,N_2449);
xor U4280 (N_4280,N_2138,N_1936);
xor U4281 (N_4281,N_788,N_2835);
nor U4282 (N_4282,N_600,N_2211);
or U4283 (N_4283,N_2822,N_1797);
or U4284 (N_4284,N_634,N_2729);
xor U4285 (N_4285,N_971,N_707);
xor U4286 (N_4286,N_2168,N_2412);
nand U4287 (N_4287,N_2117,N_1425);
or U4288 (N_4288,N_443,N_2325);
and U4289 (N_4289,N_364,N_2612);
nand U4290 (N_4290,N_2555,N_1120);
or U4291 (N_4291,N_2421,N_943);
nand U4292 (N_4292,N_1495,N_862);
nor U4293 (N_4293,N_2080,N_796);
nor U4294 (N_4294,N_1246,N_1931);
and U4295 (N_4295,N_2406,N_1669);
or U4296 (N_4296,N_1119,N_2354);
and U4297 (N_4297,N_451,N_2533);
and U4298 (N_4298,N_564,N_2515);
xnor U4299 (N_4299,N_1666,N_1947);
or U4300 (N_4300,N_2792,N_1136);
nor U4301 (N_4301,N_355,N_173);
nand U4302 (N_4302,N_1336,N_2904);
and U4303 (N_4303,N_1024,N_1959);
nand U4304 (N_4304,N_428,N_1031);
xnor U4305 (N_4305,N_1317,N_1045);
nor U4306 (N_4306,N_2176,N_22);
and U4307 (N_4307,N_375,N_1070);
nand U4308 (N_4308,N_2268,N_2162);
and U4309 (N_4309,N_2442,N_1318);
nand U4310 (N_4310,N_74,N_1806);
nand U4311 (N_4311,N_2591,N_2257);
nand U4312 (N_4312,N_382,N_1017);
or U4313 (N_4313,N_106,N_1227);
nor U4314 (N_4314,N_689,N_2025);
nand U4315 (N_4315,N_1545,N_783);
or U4316 (N_4316,N_2487,N_1068);
or U4317 (N_4317,N_1039,N_281);
nor U4318 (N_4318,N_776,N_1765);
nand U4319 (N_4319,N_925,N_2646);
and U4320 (N_4320,N_270,N_1197);
and U4321 (N_4321,N_620,N_697);
nand U4322 (N_4322,N_1860,N_110);
nor U4323 (N_4323,N_2329,N_2981);
or U4324 (N_4324,N_1598,N_238);
nor U4325 (N_4325,N_2009,N_2674);
nor U4326 (N_4326,N_2284,N_2910);
or U4327 (N_4327,N_772,N_490);
nor U4328 (N_4328,N_989,N_204);
nor U4329 (N_4329,N_2788,N_2472);
nand U4330 (N_4330,N_1081,N_2889);
nor U4331 (N_4331,N_615,N_1827);
nand U4332 (N_4332,N_1852,N_1195);
nand U4333 (N_4333,N_1608,N_2220);
and U4334 (N_4334,N_533,N_1344);
and U4335 (N_4335,N_1861,N_133);
nor U4336 (N_4336,N_1395,N_526);
nor U4337 (N_4337,N_181,N_1339);
or U4338 (N_4338,N_666,N_605);
or U4339 (N_4339,N_1567,N_2014);
nor U4340 (N_4340,N_2829,N_1312);
nor U4341 (N_4341,N_1248,N_1436);
or U4342 (N_4342,N_1064,N_2732);
and U4343 (N_4343,N_558,N_1723);
or U4344 (N_4344,N_1699,N_1865);
nor U4345 (N_4345,N_633,N_2004);
nor U4346 (N_4346,N_2105,N_1169);
and U4347 (N_4347,N_1301,N_2636);
and U4348 (N_4348,N_1314,N_967);
nor U4349 (N_4349,N_2918,N_1367);
and U4350 (N_4350,N_2831,N_2454);
nor U4351 (N_4351,N_265,N_2171);
nand U4352 (N_4352,N_1864,N_357);
nand U4353 (N_4353,N_2504,N_2063);
xnor U4354 (N_4354,N_1565,N_180);
xnor U4355 (N_4355,N_949,N_1946);
or U4356 (N_4356,N_201,N_939);
and U4357 (N_4357,N_2289,N_2741);
nand U4358 (N_4358,N_1818,N_245);
xnor U4359 (N_4359,N_1592,N_727);
nor U4360 (N_4360,N_2302,N_1483);
and U4361 (N_4361,N_2017,N_1234);
and U4362 (N_4362,N_2993,N_1176);
or U4363 (N_4363,N_1889,N_881);
or U4364 (N_4364,N_1104,N_1630);
and U4365 (N_4365,N_2470,N_1306);
or U4366 (N_4366,N_2789,N_1577);
nand U4367 (N_4367,N_1384,N_1719);
xor U4368 (N_4368,N_2594,N_2525);
and U4369 (N_4369,N_2240,N_948);
or U4370 (N_4370,N_1276,N_839);
or U4371 (N_4371,N_1760,N_1226);
nor U4372 (N_4372,N_1997,N_2509);
or U4373 (N_4373,N_147,N_2456);
nor U4374 (N_4374,N_952,N_2432);
nor U4375 (N_4375,N_2261,N_191);
and U4376 (N_4376,N_835,N_1811);
xor U4377 (N_4377,N_2045,N_752);
and U4378 (N_4378,N_2666,N_358);
and U4379 (N_4379,N_529,N_1054);
and U4380 (N_4380,N_1347,N_2485);
nor U4381 (N_4381,N_1252,N_2233);
xnor U4382 (N_4382,N_275,N_2916);
nand U4383 (N_4383,N_928,N_2606);
nand U4384 (N_4384,N_2075,N_819);
or U4385 (N_4385,N_2603,N_804);
nand U4386 (N_4386,N_1705,N_743);
nor U4387 (N_4387,N_2424,N_103);
nand U4388 (N_4388,N_98,N_2170);
or U4389 (N_4389,N_1570,N_2915);
or U4390 (N_4390,N_2778,N_2197);
or U4391 (N_4391,N_2042,N_2970);
or U4392 (N_4392,N_262,N_1549);
nor U4393 (N_4393,N_2143,N_1372);
xor U4394 (N_4394,N_525,N_101);
nor U4395 (N_4395,N_487,N_2174);
and U4396 (N_4396,N_2880,N_2274);
nand U4397 (N_4397,N_884,N_2388);
nand U4398 (N_4398,N_2086,N_996);
and U4399 (N_4399,N_2293,N_2875);
nor U4400 (N_4400,N_1394,N_1683);
nand U4401 (N_4401,N_2188,N_1099);
nand U4402 (N_4402,N_2828,N_959);
and U4403 (N_4403,N_1812,N_2078);
nand U4404 (N_4404,N_142,N_1984);
nor U4405 (N_4405,N_2436,N_905);
nor U4406 (N_4406,N_327,N_2408);
nor U4407 (N_4407,N_1320,N_2744);
nand U4408 (N_4408,N_334,N_993);
nand U4409 (N_4409,N_507,N_2592);
and U4410 (N_4410,N_2568,N_885);
and U4411 (N_4411,N_95,N_814);
nand U4412 (N_4412,N_356,N_97);
or U4413 (N_4413,N_475,N_2896);
nor U4414 (N_4414,N_2965,N_1712);
nand U4415 (N_4415,N_1076,N_2311);
or U4416 (N_4416,N_2838,N_2640);
nor U4417 (N_4417,N_1768,N_28);
or U4418 (N_4418,N_1027,N_453);
or U4419 (N_4419,N_1756,N_108);
nand U4420 (N_4420,N_2418,N_1680);
and U4421 (N_4421,N_62,N_827);
and U4422 (N_4422,N_2824,N_2517);
nand U4423 (N_4423,N_383,N_897);
and U4424 (N_4424,N_1876,N_725);
or U4425 (N_4425,N_2236,N_760);
xnor U4426 (N_4426,N_63,N_894);
xnor U4427 (N_4427,N_163,N_945);
nor U4428 (N_4428,N_2520,N_1556);
or U4429 (N_4429,N_2113,N_513);
nor U4430 (N_4430,N_1443,N_2847);
nor U4431 (N_4431,N_1391,N_1419);
or U4432 (N_4432,N_2797,N_1036);
and U4433 (N_4433,N_2833,N_2628);
nor U4434 (N_4434,N_2494,N_2541);
nand U4435 (N_4435,N_431,N_2733);
nand U4436 (N_4436,N_2216,N_2755);
nand U4437 (N_4437,N_42,N_900);
xor U4438 (N_4438,N_1758,N_2704);
or U4439 (N_4439,N_632,N_2598);
or U4440 (N_4440,N_1667,N_21);
nor U4441 (N_4441,N_16,N_499);
and U4442 (N_4442,N_1603,N_1535);
and U4443 (N_4443,N_2212,N_1704);
nand U4444 (N_4444,N_1080,N_681);
xor U4445 (N_4445,N_1065,N_1880);
nand U4446 (N_4446,N_1529,N_2121);
nor U4447 (N_4447,N_1107,N_292);
nand U4448 (N_4448,N_1894,N_923);
nor U4449 (N_4449,N_2647,N_527);
and U4450 (N_4450,N_2650,N_2607);
nand U4451 (N_4451,N_2809,N_1892);
xnor U4452 (N_4452,N_2482,N_263);
or U4453 (N_4453,N_901,N_2464);
or U4454 (N_4454,N_2820,N_1769);
and U4455 (N_4455,N_2194,N_2370);
nand U4456 (N_4456,N_1506,N_1859);
nor U4457 (N_4457,N_2584,N_1691);
xnor U4458 (N_4458,N_2564,N_845);
nand U4459 (N_4459,N_2757,N_2049);
xnor U4460 (N_4460,N_1329,N_734);
xor U4461 (N_4461,N_2253,N_2709);
and U4462 (N_4462,N_1595,N_1050);
or U4463 (N_4463,N_2951,N_366);
nor U4464 (N_4464,N_1851,N_628);
nor U4465 (N_4465,N_1088,N_1129);
and U4466 (N_4466,N_1994,N_1287);
and U4467 (N_4467,N_1628,N_938);
and U4468 (N_4468,N_25,N_2222);
nor U4469 (N_4469,N_2239,N_223);
or U4470 (N_4470,N_2743,N_2760);
nor U4471 (N_4471,N_867,N_277);
or U4472 (N_4472,N_243,N_724);
xnor U4473 (N_4473,N_588,N_1544);
xor U4474 (N_4474,N_1377,N_332);
or U4475 (N_4475,N_1082,N_1763);
nor U4476 (N_4476,N_2975,N_2232);
nand U4477 (N_4477,N_1272,N_824);
nand U4478 (N_4478,N_646,N_1664);
nor U4479 (N_4479,N_2939,N_105);
or U4480 (N_4480,N_878,N_759);
nand U4481 (N_4481,N_1423,N_869);
nor U4482 (N_4482,N_2637,N_863);
and U4483 (N_4483,N_738,N_2361);
and U4484 (N_4484,N_1798,N_1725);
nand U4485 (N_4485,N_2842,N_2104);
and U4486 (N_4486,N_229,N_2629);
nand U4487 (N_4487,N_2244,N_997);
or U4488 (N_4488,N_373,N_415);
nand U4489 (N_4489,N_1972,N_1167);
xnor U4490 (N_4490,N_155,N_1708);
xnor U4491 (N_4491,N_2288,N_1449);
nand U4492 (N_4492,N_1353,N_322);
nand U4493 (N_4493,N_1401,N_1893);
and U4494 (N_4494,N_309,N_629);
nor U4495 (N_4495,N_1208,N_1832);
or U4496 (N_4496,N_1838,N_515);
nand U4497 (N_4497,N_2663,N_1554);
nand U4498 (N_4498,N_577,N_2597);
or U4499 (N_4499,N_2337,N_589);
nand U4500 (N_4500,N_1891,N_2798);
xnor U4501 (N_4501,N_2852,N_2113);
nor U4502 (N_4502,N_2507,N_1786);
and U4503 (N_4503,N_1036,N_205);
nor U4504 (N_4504,N_526,N_2890);
nand U4505 (N_4505,N_2350,N_865);
and U4506 (N_4506,N_1639,N_1252);
nand U4507 (N_4507,N_2869,N_1712);
or U4508 (N_4508,N_2722,N_1972);
or U4509 (N_4509,N_2399,N_2381);
and U4510 (N_4510,N_2622,N_1666);
nor U4511 (N_4511,N_0,N_1155);
nor U4512 (N_4512,N_237,N_2148);
and U4513 (N_4513,N_1419,N_2677);
xnor U4514 (N_4514,N_2056,N_2811);
nand U4515 (N_4515,N_2174,N_511);
nor U4516 (N_4516,N_2637,N_677);
nor U4517 (N_4517,N_262,N_1902);
or U4518 (N_4518,N_2669,N_1722);
nor U4519 (N_4519,N_2013,N_420);
nor U4520 (N_4520,N_1997,N_702);
and U4521 (N_4521,N_1518,N_1113);
nor U4522 (N_4522,N_2099,N_1675);
or U4523 (N_4523,N_1164,N_2710);
nand U4524 (N_4524,N_1903,N_2143);
xor U4525 (N_4525,N_1211,N_2204);
or U4526 (N_4526,N_2635,N_2036);
or U4527 (N_4527,N_1278,N_1534);
or U4528 (N_4528,N_654,N_2041);
nor U4529 (N_4529,N_525,N_2886);
nor U4530 (N_4530,N_640,N_536);
nor U4531 (N_4531,N_1995,N_792);
or U4532 (N_4532,N_2852,N_2762);
and U4533 (N_4533,N_1518,N_799);
xnor U4534 (N_4534,N_43,N_1480);
or U4535 (N_4535,N_1023,N_2377);
nand U4536 (N_4536,N_1549,N_1893);
nor U4537 (N_4537,N_224,N_2577);
or U4538 (N_4538,N_1980,N_2071);
nor U4539 (N_4539,N_1213,N_2168);
nor U4540 (N_4540,N_197,N_764);
or U4541 (N_4541,N_2474,N_2439);
and U4542 (N_4542,N_630,N_2063);
nor U4543 (N_4543,N_933,N_1538);
and U4544 (N_4544,N_2214,N_2906);
nor U4545 (N_4545,N_18,N_2943);
nand U4546 (N_4546,N_1765,N_1230);
or U4547 (N_4547,N_2011,N_1283);
or U4548 (N_4548,N_1627,N_674);
nand U4549 (N_4549,N_757,N_2040);
nor U4550 (N_4550,N_1000,N_2049);
or U4551 (N_4551,N_984,N_1036);
xnor U4552 (N_4552,N_967,N_932);
and U4553 (N_4553,N_446,N_2176);
and U4554 (N_4554,N_1765,N_917);
and U4555 (N_4555,N_1379,N_2736);
nor U4556 (N_4556,N_910,N_182);
and U4557 (N_4557,N_283,N_2192);
or U4558 (N_4558,N_1540,N_1299);
or U4559 (N_4559,N_2893,N_1815);
xnor U4560 (N_4560,N_236,N_2055);
and U4561 (N_4561,N_66,N_1140);
nand U4562 (N_4562,N_1668,N_798);
xor U4563 (N_4563,N_1617,N_136);
and U4564 (N_4564,N_1259,N_1879);
nor U4565 (N_4565,N_556,N_1677);
or U4566 (N_4566,N_2783,N_1032);
or U4567 (N_4567,N_1073,N_2325);
nor U4568 (N_4568,N_811,N_280);
nand U4569 (N_4569,N_650,N_1318);
nor U4570 (N_4570,N_1321,N_2309);
or U4571 (N_4571,N_535,N_2522);
nand U4572 (N_4572,N_1858,N_2926);
or U4573 (N_4573,N_1225,N_1989);
nor U4574 (N_4574,N_1010,N_1197);
nor U4575 (N_4575,N_1000,N_1058);
or U4576 (N_4576,N_2160,N_918);
nand U4577 (N_4577,N_325,N_2429);
nand U4578 (N_4578,N_2607,N_2616);
or U4579 (N_4579,N_2632,N_1204);
or U4580 (N_4580,N_1248,N_478);
nor U4581 (N_4581,N_735,N_2335);
and U4582 (N_4582,N_1349,N_1291);
and U4583 (N_4583,N_952,N_2291);
xnor U4584 (N_4584,N_2802,N_827);
nand U4585 (N_4585,N_2582,N_1744);
nor U4586 (N_4586,N_1519,N_2056);
and U4587 (N_4587,N_2995,N_1155);
nor U4588 (N_4588,N_819,N_1371);
nand U4589 (N_4589,N_962,N_822);
nand U4590 (N_4590,N_1690,N_943);
and U4591 (N_4591,N_2861,N_2174);
or U4592 (N_4592,N_1990,N_2096);
nand U4593 (N_4593,N_519,N_859);
or U4594 (N_4594,N_1002,N_364);
xnor U4595 (N_4595,N_699,N_70);
nor U4596 (N_4596,N_1268,N_2173);
nand U4597 (N_4597,N_330,N_874);
xor U4598 (N_4598,N_2002,N_2709);
nand U4599 (N_4599,N_1580,N_724);
nor U4600 (N_4600,N_170,N_328);
and U4601 (N_4601,N_482,N_2244);
xnor U4602 (N_4602,N_593,N_2865);
nor U4603 (N_4603,N_347,N_2557);
nor U4604 (N_4604,N_2518,N_2738);
nand U4605 (N_4605,N_1090,N_431);
nor U4606 (N_4606,N_2870,N_1020);
and U4607 (N_4607,N_514,N_1856);
or U4608 (N_4608,N_2902,N_2182);
nand U4609 (N_4609,N_1485,N_140);
nor U4610 (N_4610,N_1178,N_2237);
nor U4611 (N_4611,N_1708,N_379);
and U4612 (N_4612,N_2191,N_1056);
and U4613 (N_4613,N_2433,N_2028);
nand U4614 (N_4614,N_1199,N_2907);
and U4615 (N_4615,N_2192,N_1312);
or U4616 (N_4616,N_1351,N_526);
and U4617 (N_4617,N_2627,N_2111);
nor U4618 (N_4618,N_2753,N_1185);
nand U4619 (N_4619,N_2862,N_415);
nand U4620 (N_4620,N_77,N_1723);
and U4621 (N_4621,N_1531,N_2607);
nor U4622 (N_4622,N_2160,N_1939);
nor U4623 (N_4623,N_312,N_990);
nand U4624 (N_4624,N_1058,N_2357);
and U4625 (N_4625,N_620,N_153);
and U4626 (N_4626,N_510,N_224);
xnor U4627 (N_4627,N_563,N_2053);
nand U4628 (N_4628,N_253,N_445);
or U4629 (N_4629,N_560,N_213);
or U4630 (N_4630,N_1105,N_2380);
and U4631 (N_4631,N_2684,N_156);
nor U4632 (N_4632,N_1634,N_2485);
xnor U4633 (N_4633,N_2907,N_890);
nand U4634 (N_4634,N_15,N_2551);
or U4635 (N_4635,N_2864,N_45);
nand U4636 (N_4636,N_1052,N_212);
or U4637 (N_4637,N_1372,N_1177);
nor U4638 (N_4638,N_905,N_1149);
and U4639 (N_4639,N_1721,N_2580);
and U4640 (N_4640,N_461,N_2869);
xnor U4641 (N_4641,N_524,N_1819);
and U4642 (N_4642,N_228,N_871);
nand U4643 (N_4643,N_1250,N_1635);
and U4644 (N_4644,N_1730,N_1699);
and U4645 (N_4645,N_1050,N_2278);
or U4646 (N_4646,N_131,N_919);
or U4647 (N_4647,N_130,N_350);
nor U4648 (N_4648,N_1957,N_2841);
nand U4649 (N_4649,N_2503,N_1800);
or U4650 (N_4650,N_1214,N_2959);
or U4651 (N_4651,N_1923,N_2020);
or U4652 (N_4652,N_2899,N_2580);
or U4653 (N_4653,N_2631,N_205);
nand U4654 (N_4654,N_2910,N_2802);
nand U4655 (N_4655,N_1065,N_2523);
and U4656 (N_4656,N_2087,N_1354);
nand U4657 (N_4657,N_1054,N_1560);
and U4658 (N_4658,N_2210,N_119);
nor U4659 (N_4659,N_754,N_2175);
and U4660 (N_4660,N_2354,N_366);
nor U4661 (N_4661,N_432,N_422);
and U4662 (N_4662,N_1976,N_851);
or U4663 (N_4663,N_1783,N_428);
and U4664 (N_4664,N_709,N_2735);
or U4665 (N_4665,N_324,N_788);
or U4666 (N_4666,N_1504,N_2567);
and U4667 (N_4667,N_1996,N_2017);
or U4668 (N_4668,N_2045,N_700);
or U4669 (N_4669,N_2761,N_780);
nor U4670 (N_4670,N_181,N_680);
and U4671 (N_4671,N_2241,N_2816);
or U4672 (N_4672,N_1931,N_1585);
or U4673 (N_4673,N_1626,N_1327);
nor U4674 (N_4674,N_1922,N_1738);
and U4675 (N_4675,N_2573,N_1108);
or U4676 (N_4676,N_92,N_2368);
and U4677 (N_4677,N_780,N_918);
and U4678 (N_4678,N_707,N_1918);
and U4679 (N_4679,N_2690,N_48);
xnor U4680 (N_4680,N_1724,N_448);
nor U4681 (N_4681,N_458,N_250);
and U4682 (N_4682,N_760,N_1311);
or U4683 (N_4683,N_363,N_1988);
or U4684 (N_4684,N_2711,N_2576);
nand U4685 (N_4685,N_243,N_1595);
or U4686 (N_4686,N_2420,N_2617);
nand U4687 (N_4687,N_1011,N_2615);
nand U4688 (N_4688,N_1608,N_2175);
nand U4689 (N_4689,N_2002,N_1060);
nor U4690 (N_4690,N_2522,N_590);
or U4691 (N_4691,N_977,N_2160);
or U4692 (N_4692,N_696,N_1938);
nand U4693 (N_4693,N_1526,N_1813);
nand U4694 (N_4694,N_1264,N_2492);
nor U4695 (N_4695,N_2627,N_2968);
nand U4696 (N_4696,N_200,N_62);
nor U4697 (N_4697,N_2533,N_858);
or U4698 (N_4698,N_2479,N_2399);
nor U4699 (N_4699,N_1563,N_6);
nand U4700 (N_4700,N_632,N_700);
nand U4701 (N_4701,N_245,N_1836);
nor U4702 (N_4702,N_2949,N_2907);
nand U4703 (N_4703,N_1381,N_2628);
nor U4704 (N_4704,N_1244,N_2126);
and U4705 (N_4705,N_588,N_874);
or U4706 (N_4706,N_2002,N_2868);
and U4707 (N_4707,N_2289,N_2077);
or U4708 (N_4708,N_2515,N_1796);
nand U4709 (N_4709,N_2150,N_2257);
nor U4710 (N_4710,N_1003,N_1190);
nor U4711 (N_4711,N_810,N_1556);
or U4712 (N_4712,N_2028,N_2106);
nand U4713 (N_4713,N_2389,N_1003);
or U4714 (N_4714,N_2404,N_180);
or U4715 (N_4715,N_1879,N_1892);
nor U4716 (N_4716,N_2156,N_574);
nand U4717 (N_4717,N_2835,N_278);
nor U4718 (N_4718,N_1165,N_77);
xor U4719 (N_4719,N_369,N_309);
nor U4720 (N_4720,N_1992,N_269);
xnor U4721 (N_4721,N_2749,N_2286);
and U4722 (N_4722,N_366,N_1263);
and U4723 (N_4723,N_1788,N_344);
nand U4724 (N_4724,N_2569,N_1473);
nand U4725 (N_4725,N_2953,N_1310);
xnor U4726 (N_4726,N_71,N_2033);
or U4727 (N_4727,N_1404,N_1328);
nor U4728 (N_4728,N_183,N_1272);
xor U4729 (N_4729,N_2474,N_195);
nor U4730 (N_4730,N_576,N_2682);
nor U4731 (N_4731,N_1985,N_1417);
nand U4732 (N_4732,N_2499,N_726);
and U4733 (N_4733,N_1308,N_2320);
xnor U4734 (N_4734,N_2844,N_1587);
or U4735 (N_4735,N_2715,N_887);
nor U4736 (N_4736,N_2649,N_1876);
or U4737 (N_4737,N_606,N_2940);
nand U4738 (N_4738,N_267,N_258);
xnor U4739 (N_4739,N_1460,N_1628);
xnor U4740 (N_4740,N_2898,N_178);
nand U4741 (N_4741,N_2201,N_2508);
or U4742 (N_4742,N_856,N_2154);
xnor U4743 (N_4743,N_1900,N_2918);
nor U4744 (N_4744,N_2725,N_1425);
xnor U4745 (N_4745,N_1626,N_2690);
nand U4746 (N_4746,N_366,N_1674);
or U4747 (N_4747,N_1187,N_142);
nand U4748 (N_4748,N_1727,N_22);
or U4749 (N_4749,N_2049,N_1314);
nand U4750 (N_4750,N_1952,N_90);
or U4751 (N_4751,N_823,N_1287);
and U4752 (N_4752,N_488,N_2708);
and U4753 (N_4753,N_1703,N_284);
nor U4754 (N_4754,N_463,N_2595);
nand U4755 (N_4755,N_2666,N_1860);
and U4756 (N_4756,N_1756,N_1016);
nor U4757 (N_4757,N_904,N_2287);
or U4758 (N_4758,N_2744,N_1366);
nor U4759 (N_4759,N_2997,N_868);
or U4760 (N_4760,N_2984,N_1111);
nand U4761 (N_4761,N_2652,N_754);
and U4762 (N_4762,N_2362,N_2969);
nand U4763 (N_4763,N_433,N_1695);
and U4764 (N_4764,N_1840,N_405);
and U4765 (N_4765,N_204,N_1021);
nor U4766 (N_4766,N_2718,N_1863);
and U4767 (N_4767,N_653,N_1981);
or U4768 (N_4768,N_1623,N_1148);
or U4769 (N_4769,N_2599,N_2871);
and U4770 (N_4770,N_2771,N_102);
nand U4771 (N_4771,N_1922,N_1443);
nor U4772 (N_4772,N_2198,N_755);
nor U4773 (N_4773,N_143,N_2944);
nor U4774 (N_4774,N_1532,N_2007);
nor U4775 (N_4775,N_1313,N_2533);
and U4776 (N_4776,N_2676,N_1701);
and U4777 (N_4777,N_2900,N_2045);
nor U4778 (N_4778,N_2603,N_87);
nor U4779 (N_4779,N_292,N_2629);
nand U4780 (N_4780,N_314,N_548);
and U4781 (N_4781,N_1392,N_1556);
nor U4782 (N_4782,N_1069,N_927);
xor U4783 (N_4783,N_1255,N_744);
nand U4784 (N_4784,N_1193,N_2567);
xor U4785 (N_4785,N_1702,N_1600);
nor U4786 (N_4786,N_2471,N_1320);
nor U4787 (N_4787,N_381,N_1003);
or U4788 (N_4788,N_757,N_300);
or U4789 (N_4789,N_433,N_2144);
nor U4790 (N_4790,N_786,N_859);
or U4791 (N_4791,N_1005,N_1308);
xnor U4792 (N_4792,N_2490,N_2987);
nor U4793 (N_4793,N_2633,N_2354);
or U4794 (N_4794,N_1114,N_2107);
nor U4795 (N_4795,N_408,N_2053);
or U4796 (N_4796,N_2976,N_2049);
nor U4797 (N_4797,N_200,N_585);
nor U4798 (N_4798,N_616,N_2563);
or U4799 (N_4799,N_501,N_134);
nand U4800 (N_4800,N_2789,N_1867);
nor U4801 (N_4801,N_738,N_894);
xnor U4802 (N_4802,N_1742,N_959);
and U4803 (N_4803,N_505,N_1164);
or U4804 (N_4804,N_1674,N_2337);
xor U4805 (N_4805,N_2204,N_434);
xnor U4806 (N_4806,N_2085,N_1418);
and U4807 (N_4807,N_651,N_343);
nand U4808 (N_4808,N_989,N_2470);
nand U4809 (N_4809,N_1734,N_2186);
and U4810 (N_4810,N_256,N_1360);
or U4811 (N_4811,N_1607,N_138);
nand U4812 (N_4812,N_1545,N_1274);
nand U4813 (N_4813,N_763,N_1049);
xnor U4814 (N_4814,N_1902,N_22);
nand U4815 (N_4815,N_812,N_1651);
and U4816 (N_4816,N_2669,N_203);
nand U4817 (N_4817,N_898,N_2430);
or U4818 (N_4818,N_1765,N_2995);
nor U4819 (N_4819,N_541,N_2093);
and U4820 (N_4820,N_2566,N_1573);
and U4821 (N_4821,N_2873,N_2868);
xor U4822 (N_4822,N_2410,N_1859);
nor U4823 (N_4823,N_530,N_468);
and U4824 (N_4824,N_74,N_1839);
nor U4825 (N_4825,N_1395,N_2516);
and U4826 (N_4826,N_2537,N_1747);
nor U4827 (N_4827,N_2501,N_1954);
nor U4828 (N_4828,N_1802,N_2625);
or U4829 (N_4829,N_383,N_314);
nor U4830 (N_4830,N_620,N_1727);
nand U4831 (N_4831,N_1611,N_600);
and U4832 (N_4832,N_2869,N_127);
xnor U4833 (N_4833,N_2899,N_2285);
nor U4834 (N_4834,N_1628,N_2653);
nand U4835 (N_4835,N_70,N_2271);
and U4836 (N_4836,N_1766,N_2150);
and U4837 (N_4837,N_1603,N_1776);
nor U4838 (N_4838,N_1482,N_694);
nor U4839 (N_4839,N_1917,N_2167);
nor U4840 (N_4840,N_1479,N_529);
nand U4841 (N_4841,N_1041,N_88);
nor U4842 (N_4842,N_2627,N_1767);
nor U4843 (N_4843,N_2269,N_1710);
nand U4844 (N_4844,N_542,N_2741);
or U4845 (N_4845,N_1439,N_29);
or U4846 (N_4846,N_87,N_1944);
nand U4847 (N_4847,N_2518,N_1348);
and U4848 (N_4848,N_1547,N_2956);
nand U4849 (N_4849,N_894,N_1312);
or U4850 (N_4850,N_1926,N_2706);
nor U4851 (N_4851,N_2957,N_1434);
nand U4852 (N_4852,N_2424,N_183);
and U4853 (N_4853,N_2457,N_2686);
xor U4854 (N_4854,N_73,N_2705);
or U4855 (N_4855,N_8,N_528);
nand U4856 (N_4856,N_2283,N_2807);
or U4857 (N_4857,N_241,N_2731);
xor U4858 (N_4858,N_2625,N_1102);
nand U4859 (N_4859,N_2036,N_194);
and U4860 (N_4860,N_608,N_579);
nand U4861 (N_4861,N_2089,N_1134);
nor U4862 (N_4862,N_1767,N_2582);
nand U4863 (N_4863,N_83,N_2430);
and U4864 (N_4864,N_1270,N_1559);
or U4865 (N_4865,N_1666,N_1067);
and U4866 (N_4866,N_1353,N_1967);
or U4867 (N_4867,N_2296,N_2946);
nor U4868 (N_4868,N_1257,N_198);
and U4869 (N_4869,N_2501,N_1151);
nor U4870 (N_4870,N_1522,N_1383);
nand U4871 (N_4871,N_1224,N_610);
nand U4872 (N_4872,N_263,N_2658);
nand U4873 (N_4873,N_918,N_1088);
and U4874 (N_4874,N_2584,N_1682);
and U4875 (N_4875,N_2467,N_2563);
and U4876 (N_4876,N_2729,N_1140);
nor U4877 (N_4877,N_221,N_436);
nor U4878 (N_4878,N_2590,N_1805);
xnor U4879 (N_4879,N_868,N_2755);
nor U4880 (N_4880,N_2952,N_1337);
or U4881 (N_4881,N_100,N_745);
and U4882 (N_4882,N_940,N_2718);
and U4883 (N_4883,N_2260,N_2096);
or U4884 (N_4884,N_1800,N_414);
and U4885 (N_4885,N_2656,N_702);
nand U4886 (N_4886,N_2262,N_2008);
or U4887 (N_4887,N_1808,N_1210);
xnor U4888 (N_4888,N_1997,N_996);
nor U4889 (N_4889,N_2439,N_2182);
or U4890 (N_4890,N_2480,N_1787);
nor U4891 (N_4891,N_1255,N_1585);
xnor U4892 (N_4892,N_829,N_1298);
and U4893 (N_4893,N_565,N_1702);
nand U4894 (N_4894,N_2978,N_1996);
and U4895 (N_4895,N_346,N_2856);
nand U4896 (N_4896,N_1004,N_38);
nor U4897 (N_4897,N_803,N_1689);
or U4898 (N_4898,N_2790,N_2064);
nand U4899 (N_4899,N_647,N_731);
nor U4900 (N_4900,N_1836,N_2347);
and U4901 (N_4901,N_1921,N_44);
or U4902 (N_4902,N_2296,N_2652);
and U4903 (N_4903,N_2352,N_2848);
or U4904 (N_4904,N_1950,N_333);
and U4905 (N_4905,N_1865,N_680);
nor U4906 (N_4906,N_273,N_2256);
or U4907 (N_4907,N_2442,N_1390);
xnor U4908 (N_4908,N_2880,N_945);
and U4909 (N_4909,N_396,N_2466);
nor U4910 (N_4910,N_1571,N_2061);
xnor U4911 (N_4911,N_2425,N_2142);
nor U4912 (N_4912,N_1189,N_395);
and U4913 (N_4913,N_2755,N_1397);
nand U4914 (N_4914,N_1616,N_2696);
xnor U4915 (N_4915,N_82,N_943);
or U4916 (N_4916,N_2467,N_754);
or U4917 (N_4917,N_1077,N_1905);
nand U4918 (N_4918,N_952,N_1440);
nand U4919 (N_4919,N_428,N_2234);
nand U4920 (N_4920,N_2714,N_1563);
nor U4921 (N_4921,N_2573,N_1950);
nand U4922 (N_4922,N_988,N_927);
and U4923 (N_4923,N_2129,N_1667);
nand U4924 (N_4924,N_1512,N_2135);
nor U4925 (N_4925,N_1828,N_2042);
nand U4926 (N_4926,N_1803,N_1410);
nor U4927 (N_4927,N_393,N_2149);
and U4928 (N_4928,N_1466,N_2462);
and U4929 (N_4929,N_1348,N_2955);
nand U4930 (N_4930,N_1403,N_2792);
and U4931 (N_4931,N_1231,N_1661);
or U4932 (N_4932,N_423,N_803);
or U4933 (N_4933,N_1781,N_2165);
and U4934 (N_4934,N_1822,N_2719);
nand U4935 (N_4935,N_1371,N_2135);
or U4936 (N_4936,N_122,N_1240);
nor U4937 (N_4937,N_1947,N_2958);
nand U4938 (N_4938,N_979,N_2460);
nor U4939 (N_4939,N_215,N_2466);
and U4940 (N_4940,N_1784,N_1690);
nand U4941 (N_4941,N_1272,N_613);
xnor U4942 (N_4942,N_2292,N_12);
or U4943 (N_4943,N_1897,N_1511);
and U4944 (N_4944,N_2929,N_712);
nand U4945 (N_4945,N_1113,N_1347);
nor U4946 (N_4946,N_194,N_1514);
nor U4947 (N_4947,N_2839,N_833);
and U4948 (N_4948,N_2386,N_1725);
and U4949 (N_4949,N_1533,N_1772);
or U4950 (N_4950,N_2566,N_2378);
and U4951 (N_4951,N_1539,N_1476);
nor U4952 (N_4952,N_733,N_1794);
nand U4953 (N_4953,N_384,N_909);
or U4954 (N_4954,N_2159,N_1487);
and U4955 (N_4955,N_1249,N_735);
and U4956 (N_4956,N_2825,N_2976);
or U4957 (N_4957,N_1001,N_2438);
or U4958 (N_4958,N_39,N_2058);
nand U4959 (N_4959,N_590,N_50);
nand U4960 (N_4960,N_2851,N_2116);
nor U4961 (N_4961,N_1335,N_1350);
or U4962 (N_4962,N_2905,N_1427);
nand U4963 (N_4963,N_2662,N_1660);
nand U4964 (N_4964,N_2955,N_125);
nor U4965 (N_4965,N_1565,N_935);
and U4966 (N_4966,N_404,N_924);
nand U4967 (N_4967,N_819,N_1569);
and U4968 (N_4968,N_2997,N_2237);
or U4969 (N_4969,N_1636,N_1881);
or U4970 (N_4970,N_1219,N_2655);
nand U4971 (N_4971,N_729,N_2342);
and U4972 (N_4972,N_2176,N_330);
xor U4973 (N_4973,N_82,N_2836);
or U4974 (N_4974,N_1141,N_726);
or U4975 (N_4975,N_2544,N_471);
and U4976 (N_4976,N_2423,N_2440);
or U4977 (N_4977,N_1502,N_1495);
nor U4978 (N_4978,N_1910,N_2536);
and U4979 (N_4979,N_1686,N_2448);
and U4980 (N_4980,N_666,N_811);
nor U4981 (N_4981,N_1901,N_334);
and U4982 (N_4982,N_2479,N_869);
and U4983 (N_4983,N_1653,N_1142);
or U4984 (N_4984,N_616,N_2961);
xnor U4985 (N_4985,N_1385,N_163);
or U4986 (N_4986,N_2664,N_255);
nor U4987 (N_4987,N_1398,N_620);
and U4988 (N_4988,N_1065,N_1267);
or U4989 (N_4989,N_711,N_889);
xor U4990 (N_4990,N_436,N_116);
xnor U4991 (N_4991,N_2810,N_549);
nor U4992 (N_4992,N_973,N_270);
nand U4993 (N_4993,N_234,N_436);
or U4994 (N_4994,N_1376,N_902);
nor U4995 (N_4995,N_624,N_2632);
nor U4996 (N_4996,N_1693,N_1417);
nand U4997 (N_4997,N_2632,N_165);
nand U4998 (N_4998,N_2773,N_774);
nand U4999 (N_4999,N_2742,N_1842);
xnor U5000 (N_5000,N_1232,N_1529);
or U5001 (N_5001,N_1807,N_929);
or U5002 (N_5002,N_2099,N_1415);
nor U5003 (N_5003,N_648,N_1625);
nand U5004 (N_5004,N_2634,N_2054);
xor U5005 (N_5005,N_560,N_442);
nand U5006 (N_5006,N_1733,N_2915);
and U5007 (N_5007,N_940,N_493);
and U5008 (N_5008,N_1040,N_2762);
nor U5009 (N_5009,N_2440,N_497);
and U5010 (N_5010,N_997,N_2288);
and U5011 (N_5011,N_2066,N_2371);
xnor U5012 (N_5012,N_151,N_1740);
or U5013 (N_5013,N_270,N_1086);
and U5014 (N_5014,N_1620,N_365);
xnor U5015 (N_5015,N_1609,N_1073);
xor U5016 (N_5016,N_1664,N_619);
or U5017 (N_5017,N_256,N_983);
nand U5018 (N_5018,N_1761,N_2518);
and U5019 (N_5019,N_2034,N_2916);
and U5020 (N_5020,N_836,N_2608);
nor U5021 (N_5021,N_1928,N_1213);
nor U5022 (N_5022,N_506,N_686);
or U5023 (N_5023,N_660,N_2281);
nor U5024 (N_5024,N_2608,N_264);
and U5025 (N_5025,N_1563,N_2229);
nor U5026 (N_5026,N_311,N_966);
and U5027 (N_5027,N_48,N_2285);
and U5028 (N_5028,N_2633,N_2265);
and U5029 (N_5029,N_2237,N_1558);
nor U5030 (N_5030,N_878,N_115);
nand U5031 (N_5031,N_2473,N_2328);
nor U5032 (N_5032,N_1557,N_1048);
nor U5033 (N_5033,N_1791,N_329);
nor U5034 (N_5034,N_132,N_1925);
nor U5035 (N_5035,N_2419,N_49);
or U5036 (N_5036,N_2064,N_2907);
or U5037 (N_5037,N_2004,N_1031);
nor U5038 (N_5038,N_2320,N_1140);
or U5039 (N_5039,N_1520,N_256);
or U5040 (N_5040,N_2381,N_949);
nand U5041 (N_5041,N_1963,N_2080);
nor U5042 (N_5042,N_1237,N_2132);
xor U5043 (N_5043,N_2881,N_1337);
nand U5044 (N_5044,N_1399,N_273);
nor U5045 (N_5045,N_2105,N_2536);
or U5046 (N_5046,N_1498,N_2611);
and U5047 (N_5047,N_591,N_2239);
nand U5048 (N_5048,N_2665,N_2768);
or U5049 (N_5049,N_1158,N_2094);
or U5050 (N_5050,N_1588,N_2260);
nor U5051 (N_5051,N_2426,N_2104);
nor U5052 (N_5052,N_2565,N_924);
or U5053 (N_5053,N_186,N_1098);
xor U5054 (N_5054,N_1345,N_1795);
nor U5055 (N_5055,N_2208,N_2818);
or U5056 (N_5056,N_126,N_2469);
and U5057 (N_5057,N_1966,N_2804);
and U5058 (N_5058,N_1028,N_277);
nor U5059 (N_5059,N_2021,N_1565);
or U5060 (N_5060,N_2543,N_1696);
nand U5061 (N_5061,N_258,N_850);
or U5062 (N_5062,N_362,N_374);
and U5063 (N_5063,N_1316,N_2322);
or U5064 (N_5064,N_2990,N_1654);
nand U5065 (N_5065,N_2733,N_2354);
nor U5066 (N_5066,N_2073,N_197);
or U5067 (N_5067,N_1522,N_885);
nand U5068 (N_5068,N_850,N_12);
and U5069 (N_5069,N_355,N_2524);
nor U5070 (N_5070,N_370,N_578);
nor U5071 (N_5071,N_1007,N_818);
nand U5072 (N_5072,N_696,N_1476);
and U5073 (N_5073,N_2617,N_2456);
and U5074 (N_5074,N_695,N_1178);
nor U5075 (N_5075,N_668,N_2913);
and U5076 (N_5076,N_823,N_700);
nor U5077 (N_5077,N_2307,N_96);
and U5078 (N_5078,N_1170,N_364);
or U5079 (N_5079,N_954,N_1989);
and U5080 (N_5080,N_1213,N_673);
nor U5081 (N_5081,N_1407,N_2385);
nand U5082 (N_5082,N_2044,N_396);
nand U5083 (N_5083,N_539,N_214);
nand U5084 (N_5084,N_2366,N_2277);
xnor U5085 (N_5085,N_2801,N_1884);
xnor U5086 (N_5086,N_1707,N_1703);
or U5087 (N_5087,N_1024,N_212);
and U5088 (N_5088,N_726,N_174);
and U5089 (N_5089,N_2792,N_1441);
xor U5090 (N_5090,N_1596,N_1558);
nand U5091 (N_5091,N_1727,N_1451);
and U5092 (N_5092,N_206,N_1815);
nor U5093 (N_5093,N_1451,N_914);
or U5094 (N_5094,N_1120,N_196);
nand U5095 (N_5095,N_1551,N_523);
or U5096 (N_5096,N_2058,N_439);
xnor U5097 (N_5097,N_697,N_458);
nand U5098 (N_5098,N_369,N_1082);
nand U5099 (N_5099,N_765,N_1251);
nand U5100 (N_5100,N_2092,N_1731);
nor U5101 (N_5101,N_854,N_1605);
nor U5102 (N_5102,N_2584,N_1186);
and U5103 (N_5103,N_2812,N_693);
and U5104 (N_5104,N_250,N_344);
and U5105 (N_5105,N_1896,N_2417);
and U5106 (N_5106,N_53,N_1804);
nor U5107 (N_5107,N_1977,N_961);
or U5108 (N_5108,N_2862,N_2112);
nand U5109 (N_5109,N_571,N_1679);
nand U5110 (N_5110,N_2250,N_1911);
or U5111 (N_5111,N_2550,N_2410);
or U5112 (N_5112,N_2199,N_2605);
nand U5113 (N_5113,N_2695,N_2812);
nor U5114 (N_5114,N_2713,N_942);
or U5115 (N_5115,N_1191,N_2948);
and U5116 (N_5116,N_674,N_2139);
and U5117 (N_5117,N_1769,N_568);
nor U5118 (N_5118,N_2097,N_2154);
nor U5119 (N_5119,N_2401,N_2845);
nand U5120 (N_5120,N_70,N_2057);
nor U5121 (N_5121,N_793,N_2713);
or U5122 (N_5122,N_36,N_1725);
and U5123 (N_5123,N_2280,N_41);
or U5124 (N_5124,N_2595,N_460);
nand U5125 (N_5125,N_1147,N_2021);
nand U5126 (N_5126,N_2510,N_1857);
nand U5127 (N_5127,N_2664,N_1057);
xor U5128 (N_5128,N_934,N_1683);
and U5129 (N_5129,N_655,N_1048);
and U5130 (N_5130,N_937,N_1813);
xor U5131 (N_5131,N_2088,N_283);
or U5132 (N_5132,N_2791,N_2453);
or U5133 (N_5133,N_156,N_157);
and U5134 (N_5134,N_1232,N_1261);
or U5135 (N_5135,N_251,N_1165);
and U5136 (N_5136,N_1500,N_292);
nor U5137 (N_5137,N_1583,N_2442);
nand U5138 (N_5138,N_2905,N_2829);
or U5139 (N_5139,N_1543,N_2737);
or U5140 (N_5140,N_515,N_329);
xor U5141 (N_5141,N_1888,N_1716);
and U5142 (N_5142,N_722,N_1842);
xor U5143 (N_5143,N_1117,N_258);
xor U5144 (N_5144,N_2965,N_808);
nand U5145 (N_5145,N_2488,N_2356);
and U5146 (N_5146,N_766,N_271);
and U5147 (N_5147,N_1728,N_1295);
and U5148 (N_5148,N_1823,N_1714);
nor U5149 (N_5149,N_1911,N_2052);
nand U5150 (N_5150,N_1026,N_1740);
and U5151 (N_5151,N_1279,N_1205);
or U5152 (N_5152,N_2012,N_1279);
or U5153 (N_5153,N_2176,N_683);
and U5154 (N_5154,N_420,N_1626);
or U5155 (N_5155,N_1677,N_454);
xnor U5156 (N_5156,N_2485,N_656);
and U5157 (N_5157,N_1394,N_2425);
nand U5158 (N_5158,N_602,N_1117);
xnor U5159 (N_5159,N_583,N_2113);
xnor U5160 (N_5160,N_2674,N_615);
xor U5161 (N_5161,N_1790,N_2205);
or U5162 (N_5162,N_391,N_2468);
nand U5163 (N_5163,N_1476,N_1004);
nand U5164 (N_5164,N_756,N_544);
or U5165 (N_5165,N_2348,N_1537);
nand U5166 (N_5166,N_2447,N_2254);
and U5167 (N_5167,N_1736,N_811);
and U5168 (N_5168,N_1502,N_1094);
nor U5169 (N_5169,N_1886,N_288);
and U5170 (N_5170,N_1564,N_1514);
and U5171 (N_5171,N_1693,N_969);
and U5172 (N_5172,N_721,N_2473);
nand U5173 (N_5173,N_1761,N_2272);
nor U5174 (N_5174,N_1968,N_2994);
nand U5175 (N_5175,N_901,N_64);
and U5176 (N_5176,N_2182,N_2035);
nand U5177 (N_5177,N_2124,N_2999);
and U5178 (N_5178,N_1206,N_2372);
or U5179 (N_5179,N_1981,N_1950);
or U5180 (N_5180,N_2668,N_579);
nand U5181 (N_5181,N_1849,N_2311);
and U5182 (N_5182,N_310,N_1826);
and U5183 (N_5183,N_1505,N_1148);
and U5184 (N_5184,N_2255,N_1809);
and U5185 (N_5185,N_2401,N_1924);
or U5186 (N_5186,N_239,N_2760);
or U5187 (N_5187,N_1062,N_518);
nand U5188 (N_5188,N_1088,N_396);
nor U5189 (N_5189,N_1893,N_679);
nand U5190 (N_5190,N_1260,N_594);
and U5191 (N_5191,N_674,N_2560);
nor U5192 (N_5192,N_1644,N_2485);
nor U5193 (N_5193,N_269,N_2330);
or U5194 (N_5194,N_569,N_72);
or U5195 (N_5195,N_1518,N_558);
nor U5196 (N_5196,N_1808,N_1431);
nor U5197 (N_5197,N_2666,N_189);
nand U5198 (N_5198,N_2256,N_581);
and U5199 (N_5199,N_1631,N_609);
and U5200 (N_5200,N_584,N_2278);
or U5201 (N_5201,N_910,N_246);
or U5202 (N_5202,N_1672,N_2697);
nand U5203 (N_5203,N_1115,N_965);
nand U5204 (N_5204,N_2576,N_1868);
nand U5205 (N_5205,N_1069,N_1969);
nand U5206 (N_5206,N_1463,N_1004);
nor U5207 (N_5207,N_1177,N_2699);
and U5208 (N_5208,N_934,N_1384);
and U5209 (N_5209,N_915,N_1752);
or U5210 (N_5210,N_2314,N_969);
nand U5211 (N_5211,N_392,N_120);
nand U5212 (N_5212,N_1098,N_2740);
or U5213 (N_5213,N_2009,N_1412);
nand U5214 (N_5214,N_2837,N_2269);
nand U5215 (N_5215,N_2336,N_1117);
nor U5216 (N_5216,N_2259,N_210);
nor U5217 (N_5217,N_2797,N_2248);
nand U5218 (N_5218,N_2648,N_2528);
or U5219 (N_5219,N_2062,N_2365);
xor U5220 (N_5220,N_2598,N_2384);
or U5221 (N_5221,N_2945,N_179);
or U5222 (N_5222,N_684,N_1185);
nor U5223 (N_5223,N_2392,N_2370);
nand U5224 (N_5224,N_514,N_2688);
nor U5225 (N_5225,N_1290,N_1168);
or U5226 (N_5226,N_2202,N_1368);
nor U5227 (N_5227,N_1041,N_2356);
or U5228 (N_5228,N_1272,N_2552);
nor U5229 (N_5229,N_2882,N_585);
xor U5230 (N_5230,N_2261,N_2109);
nor U5231 (N_5231,N_1634,N_1667);
or U5232 (N_5232,N_60,N_1957);
nor U5233 (N_5233,N_1885,N_1562);
or U5234 (N_5234,N_73,N_791);
xnor U5235 (N_5235,N_2752,N_2261);
or U5236 (N_5236,N_1909,N_1675);
or U5237 (N_5237,N_813,N_2289);
and U5238 (N_5238,N_391,N_2922);
xnor U5239 (N_5239,N_203,N_1756);
and U5240 (N_5240,N_1466,N_1130);
nor U5241 (N_5241,N_2990,N_1557);
or U5242 (N_5242,N_2700,N_1411);
nor U5243 (N_5243,N_1185,N_1065);
nor U5244 (N_5244,N_1279,N_1727);
and U5245 (N_5245,N_1500,N_1205);
nand U5246 (N_5246,N_1671,N_2197);
and U5247 (N_5247,N_312,N_477);
xor U5248 (N_5248,N_600,N_2813);
and U5249 (N_5249,N_1747,N_2089);
or U5250 (N_5250,N_844,N_2288);
nor U5251 (N_5251,N_2198,N_2649);
nor U5252 (N_5252,N_661,N_958);
nor U5253 (N_5253,N_2087,N_963);
nand U5254 (N_5254,N_1888,N_917);
and U5255 (N_5255,N_1475,N_1125);
xnor U5256 (N_5256,N_602,N_499);
nand U5257 (N_5257,N_1639,N_307);
nand U5258 (N_5258,N_1496,N_786);
and U5259 (N_5259,N_2488,N_1995);
nand U5260 (N_5260,N_2222,N_1342);
nand U5261 (N_5261,N_1866,N_408);
nor U5262 (N_5262,N_2905,N_2906);
nand U5263 (N_5263,N_1034,N_400);
xnor U5264 (N_5264,N_1336,N_2331);
and U5265 (N_5265,N_2360,N_155);
xnor U5266 (N_5266,N_1892,N_350);
nor U5267 (N_5267,N_1073,N_2430);
nor U5268 (N_5268,N_438,N_2039);
nand U5269 (N_5269,N_2512,N_2358);
or U5270 (N_5270,N_507,N_1548);
or U5271 (N_5271,N_2680,N_1894);
nand U5272 (N_5272,N_2347,N_748);
nor U5273 (N_5273,N_1984,N_844);
nor U5274 (N_5274,N_977,N_2945);
nor U5275 (N_5275,N_391,N_2159);
nor U5276 (N_5276,N_2913,N_1808);
nand U5277 (N_5277,N_381,N_640);
or U5278 (N_5278,N_2439,N_256);
nor U5279 (N_5279,N_473,N_1856);
nand U5280 (N_5280,N_1115,N_403);
nand U5281 (N_5281,N_938,N_1035);
nand U5282 (N_5282,N_2196,N_1478);
nor U5283 (N_5283,N_234,N_1245);
or U5284 (N_5284,N_789,N_2611);
or U5285 (N_5285,N_70,N_411);
and U5286 (N_5286,N_2377,N_1085);
or U5287 (N_5287,N_1059,N_280);
xnor U5288 (N_5288,N_63,N_945);
xnor U5289 (N_5289,N_1494,N_1366);
nor U5290 (N_5290,N_750,N_551);
nand U5291 (N_5291,N_1447,N_169);
or U5292 (N_5292,N_2971,N_1180);
nand U5293 (N_5293,N_2769,N_1164);
and U5294 (N_5294,N_2998,N_2567);
or U5295 (N_5295,N_2668,N_2182);
nor U5296 (N_5296,N_2390,N_1761);
nor U5297 (N_5297,N_1555,N_672);
nand U5298 (N_5298,N_781,N_2935);
nor U5299 (N_5299,N_1265,N_2291);
or U5300 (N_5300,N_2371,N_811);
nand U5301 (N_5301,N_2575,N_2672);
or U5302 (N_5302,N_137,N_1694);
or U5303 (N_5303,N_242,N_1857);
nor U5304 (N_5304,N_2366,N_1009);
xnor U5305 (N_5305,N_1084,N_2219);
nor U5306 (N_5306,N_2960,N_2866);
nor U5307 (N_5307,N_1213,N_1212);
nor U5308 (N_5308,N_1128,N_2309);
or U5309 (N_5309,N_1353,N_1211);
xnor U5310 (N_5310,N_1656,N_1659);
nor U5311 (N_5311,N_2190,N_2736);
xnor U5312 (N_5312,N_443,N_308);
nand U5313 (N_5313,N_1144,N_1824);
or U5314 (N_5314,N_579,N_1212);
nand U5315 (N_5315,N_2183,N_2476);
or U5316 (N_5316,N_2991,N_277);
nor U5317 (N_5317,N_2933,N_1847);
nand U5318 (N_5318,N_1920,N_1648);
and U5319 (N_5319,N_1551,N_1995);
or U5320 (N_5320,N_2489,N_1098);
and U5321 (N_5321,N_587,N_2526);
or U5322 (N_5322,N_1819,N_259);
nor U5323 (N_5323,N_47,N_1022);
nand U5324 (N_5324,N_325,N_2883);
and U5325 (N_5325,N_1146,N_872);
or U5326 (N_5326,N_104,N_2909);
nor U5327 (N_5327,N_1007,N_2613);
or U5328 (N_5328,N_459,N_2931);
nor U5329 (N_5329,N_1731,N_98);
or U5330 (N_5330,N_1076,N_1456);
and U5331 (N_5331,N_1777,N_2262);
nor U5332 (N_5332,N_1700,N_2333);
nand U5333 (N_5333,N_342,N_1069);
xnor U5334 (N_5334,N_299,N_933);
or U5335 (N_5335,N_45,N_1652);
nand U5336 (N_5336,N_1069,N_792);
nand U5337 (N_5337,N_1465,N_1039);
nand U5338 (N_5338,N_1592,N_1565);
and U5339 (N_5339,N_851,N_2922);
nand U5340 (N_5340,N_61,N_1775);
nor U5341 (N_5341,N_2843,N_1931);
nand U5342 (N_5342,N_1994,N_1449);
nand U5343 (N_5343,N_2503,N_1516);
nor U5344 (N_5344,N_2058,N_531);
nand U5345 (N_5345,N_2305,N_2308);
nand U5346 (N_5346,N_2402,N_2150);
nor U5347 (N_5347,N_698,N_531);
nor U5348 (N_5348,N_1542,N_707);
or U5349 (N_5349,N_2277,N_167);
nor U5350 (N_5350,N_2313,N_172);
nor U5351 (N_5351,N_686,N_625);
nor U5352 (N_5352,N_34,N_1919);
or U5353 (N_5353,N_2997,N_590);
xor U5354 (N_5354,N_2650,N_1637);
nor U5355 (N_5355,N_2224,N_2323);
xor U5356 (N_5356,N_614,N_962);
or U5357 (N_5357,N_1249,N_2429);
and U5358 (N_5358,N_2029,N_639);
and U5359 (N_5359,N_1907,N_1207);
xor U5360 (N_5360,N_2275,N_2376);
or U5361 (N_5361,N_113,N_1694);
nor U5362 (N_5362,N_1618,N_2152);
nand U5363 (N_5363,N_171,N_1296);
nand U5364 (N_5364,N_1045,N_1826);
and U5365 (N_5365,N_212,N_1467);
or U5366 (N_5366,N_1154,N_271);
and U5367 (N_5367,N_1966,N_267);
nand U5368 (N_5368,N_2390,N_2986);
nor U5369 (N_5369,N_597,N_1608);
or U5370 (N_5370,N_275,N_2300);
or U5371 (N_5371,N_1237,N_1891);
and U5372 (N_5372,N_2573,N_902);
xnor U5373 (N_5373,N_2791,N_714);
nand U5374 (N_5374,N_179,N_1630);
nor U5375 (N_5375,N_2382,N_515);
or U5376 (N_5376,N_1902,N_2397);
or U5377 (N_5377,N_1281,N_2095);
or U5378 (N_5378,N_2175,N_2684);
nor U5379 (N_5379,N_125,N_799);
and U5380 (N_5380,N_2112,N_378);
xor U5381 (N_5381,N_1270,N_2725);
nor U5382 (N_5382,N_1526,N_2564);
nand U5383 (N_5383,N_2309,N_121);
and U5384 (N_5384,N_1945,N_1638);
nand U5385 (N_5385,N_961,N_650);
and U5386 (N_5386,N_1153,N_2578);
xnor U5387 (N_5387,N_2055,N_1213);
nand U5388 (N_5388,N_2921,N_2692);
nor U5389 (N_5389,N_55,N_757);
nor U5390 (N_5390,N_2035,N_156);
and U5391 (N_5391,N_2031,N_1785);
and U5392 (N_5392,N_2773,N_2053);
nand U5393 (N_5393,N_684,N_1644);
or U5394 (N_5394,N_1832,N_702);
nand U5395 (N_5395,N_2285,N_2151);
nand U5396 (N_5396,N_529,N_386);
nor U5397 (N_5397,N_922,N_1550);
or U5398 (N_5398,N_1901,N_1470);
nand U5399 (N_5399,N_1681,N_596);
nand U5400 (N_5400,N_2637,N_2293);
or U5401 (N_5401,N_1605,N_2571);
nor U5402 (N_5402,N_1384,N_1163);
and U5403 (N_5403,N_269,N_1228);
and U5404 (N_5404,N_1841,N_1381);
nand U5405 (N_5405,N_2931,N_1928);
nand U5406 (N_5406,N_2969,N_124);
nand U5407 (N_5407,N_2003,N_703);
nor U5408 (N_5408,N_1772,N_2700);
nor U5409 (N_5409,N_2780,N_243);
xor U5410 (N_5410,N_2563,N_611);
and U5411 (N_5411,N_2510,N_1498);
nand U5412 (N_5412,N_2643,N_2562);
and U5413 (N_5413,N_2604,N_2081);
nand U5414 (N_5414,N_608,N_672);
nor U5415 (N_5415,N_2600,N_546);
or U5416 (N_5416,N_410,N_1410);
nor U5417 (N_5417,N_863,N_1006);
or U5418 (N_5418,N_1620,N_1217);
nand U5419 (N_5419,N_1134,N_786);
or U5420 (N_5420,N_535,N_1316);
nand U5421 (N_5421,N_559,N_197);
and U5422 (N_5422,N_1158,N_2293);
nand U5423 (N_5423,N_808,N_533);
or U5424 (N_5424,N_1023,N_2368);
xor U5425 (N_5425,N_749,N_2185);
and U5426 (N_5426,N_2108,N_1626);
and U5427 (N_5427,N_1453,N_481);
and U5428 (N_5428,N_2237,N_781);
nand U5429 (N_5429,N_533,N_481);
nand U5430 (N_5430,N_1750,N_659);
nand U5431 (N_5431,N_2613,N_26);
and U5432 (N_5432,N_1878,N_515);
nand U5433 (N_5433,N_2751,N_2134);
and U5434 (N_5434,N_2335,N_1488);
and U5435 (N_5435,N_585,N_68);
or U5436 (N_5436,N_2445,N_2934);
nor U5437 (N_5437,N_514,N_2508);
or U5438 (N_5438,N_86,N_1049);
or U5439 (N_5439,N_1759,N_2055);
and U5440 (N_5440,N_252,N_176);
nor U5441 (N_5441,N_463,N_2082);
nand U5442 (N_5442,N_1148,N_1958);
nand U5443 (N_5443,N_1783,N_1597);
nor U5444 (N_5444,N_1681,N_35);
and U5445 (N_5445,N_1626,N_2980);
nand U5446 (N_5446,N_2038,N_412);
or U5447 (N_5447,N_2457,N_715);
xnor U5448 (N_5448,N_1904,N_1861);
nor U5449 (N_5449,N_1416,N_1911);
nor U5450 (N_5450,N_2329,N_298);
nor U5451 (N_5451,N_1338,N_1992);
nor U5452 (N_5452,N_1024,N_2189);
and U5453 (N_5453,N_1229,N_2289);
nand U5454 (N_5454,N_2244,N_1089);
and U5455 (N_5455,N_559,N_1010);
nand U5456 (N_5456,N_2664,N_2233);
or U5457 (N_5457,N_2755,N_1854);
or U5458 (N_5458,N_1156,N_1476);
xor U5459 (N_5459,N_2416,N_38);
or U5460 (N_5460,N_2636,N_806);
or U5461 (N_5461,N_1203,N_480);
xnor U5462 (N_5462,N_2407,N_1176);
nor U5463 (N_5463,N_525,N_1631);
xnor U5464 (N_5464,N_2270,N_1236);
xor U5465 (N_5465,N_1451,N_2467);
and U5466 (N_5466,N_1238,N_1869);
or U5467 (N_5467,N_309,N_2781);
nand U5468 (N_5468,N_2328,N_359);
xnor U5469 (N_5469,N_1340,N_2267);
or U5470 (N_5470,N_719,N_1952);
nor U5471 (N_5471,N_245,N_278);
nor U5472 (N_5472,N_2682,N_1808);
nand U5473 (N_5473,N_980,N_492);
nor U5474 (N_5474,N_1691,N_318);
nor U5475 (N_5475,N_1916,N_2836);
or U5476 (N_5476,N_294,N_1486);
nand U5477 (N_5477,N_811,N_2626);
or U5478 (N_5478,N_646,N_155);
and U5479 (N_5479,N_111,N_2625);
nor U5480 (N_5480,N_1639,N_594);
and U5481 (N_5481,N_1748,N_2934);
nor U5482 (N_5482,N_1270,N_2843);
nor U5483 (N_5483,N_1601,N_597);
and U5484 (N_5484,N_67,N_831);
nand U5485 (N_5485,N_2621,N_31);
nor U5486 (N_5486,N_1735,N_1412);
nor U5487 (N_5487,N_292,N_1999);
nand U5488 (N_5488,N_1613,N_1233);
nand U5489 (N_5489,N_1623,N_1765);
xnor U5490 (N_5490,N_327,N_2405);
nor U5491 (N_5491,N_2874,N_1591);
nor U5492 (N_5492,N_1520,N_911);
nand U5493 (N_5493,N_285,N_2944);
nor U5494 (N_5494,N_2399,N_2912);
xor U5495 (N_5495,N_200,N_249);
nand U5496 (N_5496,N_106,N_1488);
or U5497 (N_5497,N_1894,N_51);
nand U5498 (N_5498,N_1774,N_481);
nor U5499 (N_5499,N_644,N_2511);
nand U5500 (N_5500,N_1925,N_2423);
and U5501 (N_5501,N_10,N_772);
or U5502 (N_5502,N_1075,N_308);
nor U5503 (N_5503,N_1480,N_2372);
and U5504 (N_5504,N_2272,N_1683);
and U5505 (N_5505,N_220,N_1358);
nand U5506 (N_5506,N_82,N_918);
nor U5507 (N_5507,N_1411,N_62);
or U5508 (N_5508,N_1088,N_2953);
and U5509 (N_5509,N_1436,N_870);
and U5510 (N_5510,N_1933,N_2911);
nand U5511 (N_5511,N_1693,N_1234);
nand U5512 (N_5512,N_1767,N_2043);
or U5513 (N_5513,N_1297,N_2025);
or U5514 (N_5514,N_2756,N_22);
nor U5515 (N_5515,N_903,N_2155);
xor U5516 (N_5516,N_2882,N_478);
or U5517 (N_5517,N_1234,N_2977);
nor U5518 (N_5518,N_918,N_666);
nor U5519 (N_5519,N_2551,N_1132);
or U5520 (N_5520,N_2444,N_1818);
nand U5521 (N_5521,N_2438,N_2467);
nand U5522 (N_5522,N_2512,N_2653);
nand U5523 (N_5523,N_1838,N_2823);
nor U5524 (N_5524,N_2207,N_2716);
nor U5525 (N_5525,N_2169,N_629);
or U5526 (N_5526,N_2404,N_1242);
xnor U5527 (N_5527,N_2938,N_1222);
or U5528 (N_5528,N_2924,N_1415);
or U5529 (N_5529,N_2009,N_127);
nor U5530 (N_5530,N_1636,N_1720);
nand U5531 (N_5531,N_472,N_690);
or U5532 (N_5532,N_1191,N_795);
and U5533 (N_5533,N_587,N_79);
xor U5534 (N_5534,N_270,N_2109);
nor U5535 (N_5535,N_465,N_621);
xor U5536 (N_5536,N_1759,N_2471);
or U5537 (N_5537,N_911,N_1207);
nor U5538 (N_5538,N_344,N_301);
nor U5539 (N_5539,N_2394,N_1896);
nand U5540 (N_5540,N_1122,N_2856);
or U5541 (N_5541,N_956,N_2480);
nand U5542 (N_5542,N_2661,N_272);
nor U5543 (N_5543,N_2283,N_2314);
or U5544 (N_5544,N_598,N_2411);
and U5545 (N_5545,N_724,N_1839);
nand U5546 (N_5546,N_833,N_1816);
nor U5547 (N_5547,N_1687,N_453);
nor U5548 (N_5548,N_2054,N_1075);
and U5549 (N_5549,N_181,N_997);
nor U5550 (N_5550,N_1204,N_657);
nor U5551 (N_5551,N_811,N_994);
nor U5552 (N_5552,N_1540,N_2126);
or U5553 (N_5553,N_805,N_1929);
nor U5554 (N_5554,N_2486,N_2458);
or U5555 (N_5555,N_2612,N_1276);
and U5556 (N_5556,N_797,N_257);
and U5557 (N_5557,N_509,N_1260);
nor U5558 (N_5558,N_2288,N_2803);
or U5559 (N_5559,N_2662,N_158);
nor U5560 (N_5560,N_193,N_1706);
or U5561 (N_5561,N_2997,N_2262);
or U5562 (N_5562,N_1720,N_1140);
nand U5563 (N_5563,N_2180,N_55);
or U5564 (N_5564,N_2704,N_2899);
or U5565 (N_5565,N_2478,N_2637);
and U5566 (N_5566,N_1047,N_371);
nor U5567 (N_5567,N_2961,N_436);
or U5568 (N_5568,N_1053,N_2596);
or U5569 (N_5569,N_631,N_925);
and U5570 (N_5570,N_1324,N_2553);
and U5571 (N_5571,N_1914,N_226);
and U5572 (N_5572,N_1844,N_1443);
nand U5573 (N_5573,N_149,N_108);
and U5574 (N_5574,N_125,N_855);
nand U5575 (N_5575,N_861,N_1599);
xor U5576 (N_5576,N_2232,N_2476);
nor U5577 (N_5577,N_772,N_2154);
and U5578 (N_5578,N_91,N_2102);
nor U5579 (N_5579,N_1967,N_251);
nand U5580 (N_5580,N_849,N_220);
and U5581 (N_5581,N_338,N_1307);
or U5582 (N_5582,N_1516,N_1208);
nand U5583 (N_5583,N_2520,N_2421);
xnor U5584 (N_5584,N_1583,N_2113);
or U5585 (N_5585,N_745,N_1442);
and U5586 (N_5586,N_2621,N_2629);
and U5587 (N_5587,N_882,N_2121);
nor U5588 (N_5588,N_278,N_373);
nor U5589 (N_5589,N_1537,N_1386);
and U5590 (N_5590,N_2837,N_693);
or U5591 (N_5591,N_1588,N_2851);
nand U5592 (N_5592,N_1986,N_643);
and U5593 (N_5593,N_2371,N_2090);
and U5594 (N_5594,N_693,N_457);
or U5595 (N_5595,N_2518,N_1601);
xor U5596 (N_5596,N_706,N_2778);
nor U5597 (N_5597,N_265,N_10);
and U5598 (N_5598,N_2111,N_1489);
or U5599 (N_5599,N_770,N_1573);
nor U5600 (N_5600,N_2349,N_1555);
nor U5601 (N_5601,N_911,N_682);
or U5602 (N_5602,N_2743,N_212);
nand U5603 (N_5603,N_1678,N_1282);
or U5604 (N_5604,N_690,N_666);
nand U5605 (N_5605,N_2481,N_319);
nor U5606 (N_5606,N_1250,N_803);
and U5607 (N_5607,N_1154,N_1679);
or U5608 (N_5608,N_290,N_421);
or U5609 (N_5609,N_1638,N_1677);
nor U5610 (N_5610,N_1255,N_80);
nor U5611 (N_5611,N_2375,N_1574);
and U5612 (N_5612,N_2786,N_921);
nor U5613 (N_5613,N_2045,N_2416);
or U5614 (N_5614,N_3,N_1837);
or U5615 (N_5615,N_311,N_2096);
or U5616 (N_5616,N_749,N_2086);
nand U5617 (N_5617,N_686,N_1708);
xor U5618 (N_5618,N_892,N_1727);
nand U5619 (N_5619,N_2587,N_1135);
or U5620 (N_5620,N_1597,N_161);
nand U5621 (N_5621,N_172,N_1609);
nor U5622 (N_5622,N_364,N_1411);
and U5623 (N_5623,N_224,N_292);
nor U5624 (N_5624,N_109,N_1358);
and U5625 (N_5625,N_668,N_2847);
nand U5626 (N_5626,N_1210,N_242);
and U5627 (N_5627,N_1131,N_2495);
nand U5628 (N_5628,N_2979,N_247);
nand U5629 (N_5629,N_1669,N_2044);
nor U5630 (N_5630,N_2573,N_120);
xnor U5631 (N_5631,N_1395,N_2992);
and U5632 (N_5632,N_1529,N_736);
nor U5633 (N_5633,N_1476,N_1819);
nor U5634 (N_5634,N_1405,N_1387);
or U5635 (N_5635,N_2866,N_2785);
nor U5636 (N_5636,N_172,N_881);
nor U5637 (N_5637,N_2377,N_1189);
and U5638 (N_5638,N_2398,N_98);
or U5639 (N_5639,N_949,N_833);
or U5640 (N_5640,N_2267,N_1803);
nor U5641 (N_5641,N_17,N_89);
or U5642 (N_5642,N_2861,N_2265);
and U5643 (N_5643,N_2010,N_624);
and U5644 (N_5644,N_144,N_301);
or U5645 (N_5645,N_2693,N_2311);
nor U5646 (N_5646,N_2733,N_2683);
or U5647 (N_5647,N_2374,N_2837);
xor U5648 (N_5648,N_1075,N_41);
or U5649 (N_5649,N_2624,N_2792);
and U5650 (N_5650,N_1249,N_1144);
nor U5651 (N_5651,N_1466,N_2262);
or U5652 (N_5652,N_930,N_1741);
nor U5653 (N_5653,N_417,N_2660);
nand U5654 (N_5654,N_1362,N_1928);
or U5655 (N_5655,N_544,N_2257);
and U5656 (N_5656,N_1194,N_1414);
nand U5657 (N_5657,N_2866,N_2882);
nor U5658 (N_5658,N_2792,N_2299);
and U5659 (N_5659,N_520,N_1475);
nor U5660 (N_5660,N_850,N_1807);
xnor U5661 (N_5661,N_1613,N_404);
nand U5662 (N_5662,N_56,N_193);
xor U5663 (N_5663,N_887,N_732);
xor U5664 (N_5664,N_1608,N_1678);
nand U5665 (N_5665,N_2338,N_2249);
nand U5666 (N_5666,N_1617,N_692);
and U5667 (N_5667,N_2064,N_1305);
nand U5668 (N_5668,N_246,N_1330);
and U5669 (N_5669,N_75,N_1607);
or U5670 (N_5670,N_303,N_2110);
nand U5671 (N_5671,N_1656,N_2734);
nor U5672 (N_5672,N_1107,N_2684);
nor U5673 (N_5673,N_1159,N_1717);
and U5674 (N_5674,N_1359,N_1680);
nor U5675 (N_5675,N_550,N_493);
and U5676 (N_5676,N_1430,N_1375);
nor U5677 (N_5677,N_1269,N_2151);
nand U5678 (N_5678,N_2799,N_1797);
and U5679 (N_5679,N_2204,N_1435);
xor U5680 (N_5680,N_320,N_2921);
nand U5681 (N_5681,N_2223,N_936);
and U5682 (N_5682,N_1300,N_1148);
nor U5683 (N_5683,N_1226,N_2376);
nand U5684 (N_5684,N_2835,N_2614);
and U5685 (N_5685,N_1089,N_1355);
nand U5686 (N_5686,N_377,N_1646);
nor U5687 (N_5687,N_866,N_1871);
nand U5688 (N_5688,N_1026,N_1507);
nand U5689 (N_5689,N_2783,N_2954);
and U5690 (N_5690,N_2849,N_1159);
or U5691 (N_5691,N_2152,N_2103);
or U5692 (N_5692,N_1412,N_473);
xor U5693 (N_5693,N_1955,N_1885);
or U5694 (N_5694,N_682,N_1673);
or U5695 (N_5695,N_2315,N_1039);
and U5696 (N_5696,N_387,N_1061);
nand U5697 (N_5697,N_2561,N_252);
xnor U5698 (N_5698,N_1494,N_351);
and U5699 (N_5699,N_2325,N_2640);
and U5700 (N_5700,N_2369,N_460);
xor U5701 (N_5701,N_3,N_784);
and U5702 (N_5702,N_1511,N_2601);
nand U5703 (N_5703,N_828,N_599);
nand U5704 (N_5704,N_1381,N_299);
nor U5705 (N_5705,N_2307,N_2628);
nand U5706 (N_5706,N_2044,N_2916);
nor U5707 (N_5707,N_222,N_1425);
nand U5708 (N_5708,N_2426,N_1793);
and U5709 (N_5709,N_2673,N_1402);
nor U5710 (N_5710,N_1340,N_647);
or U5711 (N_5711,N_1528,N_1563);
nand U5712 (N_5712,N_1871,N_1458);
and U5713 (N_5713,N_2050,N_2870);
and U5714 (N_5714,N_2313,N_333);
nor U5715 (N_5715,N_711,N_2324);
or U5716 (N_5716,N_2800,N_656);
or U5717 (N_5717,N_1480,N_2420);
or U5718 (N_5718,N_1651,N_1390);
nand U5719 (N_5719,N_772,N_2894);
and U5720 (N_5720,N_113,N_2449);
and U5721 (N_5721,N_1076,N_2004);
or U5722 (N_5722,N_963,N_1655);
or U5723 (N_5723,N_1164,N_578);
xor U5724 (N_5724,N_610,N_1282);
or U5725 (N_5725,N_1182,N_1576);
nor U5726 (N_5726,N_188,N_1151);
nor U5727 (N_5727,N_2959,N_174);
or U5728 (N_5728,N_1892,N_2528);
nor U5729 (N_5729,N_462,N_2066);
nand U5730 (N_5730,N_665,N_1322);
and U5731 (N_5731,N_614,N_699);
and U5732 (N_5732,N_2128,N_1312);
and U5733 (N_5733,N_411,N_2198);
nor U5734 (N_5734,N_943,N_1678);
and U5735 (N_5735,N_1831,N_866);
nand U5736 (N_5736,N_239,N_1741);
or U5737 (N_5737,N_2860,N_1639);
and U5738 (N_5738,N_1791,N_849);
nor U5739 (N_5739,N_699,N_2714);
nor U5740 (N_5740,N_1118,N_1037);
nor U5741 (N_5741,N_2532,N_312);
nand U5742 (N_5742,N_1963,N_2308);
nand U5743 (N_5743,N_2382,N_1514);
or U5744 (N_5744,N_1902,N_795);
nor U5745 (N_5745,N_2920,N_1727);
nand U5746 (N_5746,N_592,N_1836);
and U5747 (N_5747,N_2608,N_2194);
nor U5748 (N_5748,N_1643,N_991);
or U5749 (N_5749,N_1618,N_919);
nand U5750 (N_5750,N_2490,N_619);
xor U5751 (N_5751,N_1965,N_970);
xor U5752 (N_5752,N_878,N_807);
nor U5753 (N_5753,N_2053,N_2687);
and U5754 (N_5754,N_2320,N_2214);
nor U5755 (N_5755,N_794,N_1096);
and U5756 (N_5756,N_15,N_2268);
and U5757 (N_5757,N_2881,N_299);
xor U5758 (N_5758,N_640,N_1390);
and U5759 (N_5759,N_2784,N_225);
xnor U5760 (N_5760,N_897,N_1696);
nor U5761 (N_5761,N_1987,N_1137);
and U5762 (N_5762,N_509,N_350);
nor U5763 (N_5763,N_2101,N_2217);
and U5764 (N_5764,N_597,N_823);
nor U5765 (N_5765,N_1982,N_1617);
nor U5766 (N_5766,N_1084,N_2522);
nand U5767 (N_5767,N_50,N_2948);
xor U5768 (N_5768,N_169,N_2357);
nand U5769 (N_5769,N_39,N_655);
nor U5770 (N_5770,N_1062,N_637);
nor U5771 (N_5771,N_1711,N_1728);
or U5772 (N_5772,N_1629,N_453);
nand U5773 (N_5773,N_1855,N_432);
nor U5774 (N_5774,N_33,N_2039);
xnor U5775 (N_5775,N_372,N_2599);
or U5776 (N_5776,N_1593,N_2001);
or U5777 (N_5777,N_32,N_1227);
and U5778 (N_5778,N_749,N_2400);
nor U5779 (N_5779,N_1314,N_1788);
and U5780 (N_5780,N_1854,N_175);
nand U5781 (N_5781,N_268,N_1177);
xor U5782 (N_5782,N_330,N_2883);
or U5783 (N_5783,N_618,N_1868);
and U5784 (N_5784,N_1705,N_1738);
and U5785 (N_5785,N_1343,N_1886);
nand U5786 (N_5786,N_962,N_2420);
and U5787 (N_5787,N_2387,N_2148);
nand U5788 (N_5788,N_931,N_167);
and U5789 (N_5789,N_763,N_764);
and U5790 (N_5790,N_123,N_1086);
or U5791 (N_5791,N_1120,N_230);
nor U5792 (N_5792,N_2523,N_2989);
and U5793 (N_5793,N_700,N_754);
and U5794 (N_5794,N_2031,N_2676);
nor U5795 (N_5795,N_2065,N_1586);
nor U5796 (N_5796,N_485,N_1233);
nor U5797 (N_5797,N_426,N_2982);
nor U5798 (N_5798,N_1360,N_106);
xnor U5799 (N_5799,N_1436,N_1066);
or U5800 (N_5800,N_1625,N_2219);
and U5801 (N_5801,N_2260,N_628);
nand U5802 (N_5802,N_54,N_53);
and U5803 (N_5803,N_1732,N_698);
nor U5804 (N_5804,N_198,N_52);
nand U5805 (N_5805,N_1091,N_1751);
or U5806 (N_5806,N_829,N_583);
xor U5807 (N_5807,N_1033,N_2724);
nor U5808 (N_5808,N_459,N_656);
nor U5809 (N_5809,N_2724,N_230);
or U5810 (N_5810,N_754,N_2423);
nor U5811 (N_5811,N_1610,N_1987);
and U5812 (N_5812,N_874,N_343);
or U5813 (N_5813,N_2072,N_1153);
nor U5814 (N_5814,N_682,N_2232);
and U5815 (N_5815,N_1746,N_619);
nor U5816 (N_5816,N_1459,N_335);
and U5817 (N_5817,N_2788,N_289);
nand U5818 (N_5818,N_2416,N_923);
or U5819 (N_5819,N_1328,N_927);
nand U5820 (N_5820,N_2792,N_2457);
nand U5821 (N_5821,N_1686,N_2859);
nand U5822 (N_5822,N_586,N_2293);
and U5823 (N_5823,N_1760,N_1656);
nor U5824 (N_5824,N_2995,N_1142);
nand U5825 (N_5825,N_487,N_225);
nand U5826 (N_5826,N_2885,N_2330);
nand U5827 (N_5827,N_316,N_1982);
nor U5828 (N_5828,N_1330,N_45);
or U5829 (N_5829,N_677,N_2601);
and U5830 (N_5830,N_79,N_300);
or U5831 (N_5831,N_418,N_1144);
nand U5832 (N_5832,N_1939,N_2976);
nor U5833 (N_5833,N_2050,N_707);
nand U5834 (N_5834,N_2407,N_1246);
and U5835 (N_5835,N_2195,N_412);
nand U5836 (N_5836,N_1684,N_2161);
and U5837 (N_5837,N_2832,N_1853);
xnor U5838 (N_5838,N_1179,N_544);
nand U5839 (N_5839,N_2932,N_1731);
xnor U5840 (N_5840,N_1255,N_782);
xor U5841 (N_5841,N_1547,N_605);
nand U5842 (N_5842,N_550,N_2153);
or U5843 (N_5843,N_1407,N_2205);
nand U5844 (N_5844,N_602,N_2159);
nor U5845 (N_5845,N_1600,N_2109);
nor U5846 (N_5846,N_2725,N_854);
nand U5847 (N_5847,N_2098,N_2104);
and U5848 (N_5848,N_135,N_1145);
xnor U5849 (N_5849,N_1741,N_2917);
nor U5850 (N_5850,N_267,N_852);
nor U5851 (N_5851,N_82,N_838);
xor U5852 (N_5852,N_1137,N_1546);
and U5853 (N_5853,N_1828,N_791);
nand U5854 (N_5854,N_1399,N_635);
or U5855 (N_5855,N_660,N_461);
or U5856 (N_5856,N_1271,N_1216);
xor U5857 (N_5857,N_433,N_1864);
or U5858 (N_5858,N_1768,N_20);
nor U5859 (N_5859,N_320,N_756);
or U5860 (N_5860,N_2680,N_1689);
nand U5861 (N_5861,N_2150,N_1522);
or U5862 (N_5862,N_1055,N_1046);
nand U5863 (N_5863,N_2513,N_494);
and U5864 (N_5864,N_826,N_1733);
or U5865 (N_5865,N_2407,N_1146);
nor U5866 (N_5866,N_2549,N_1410);
or U5867 (N_5867,N_1752,N_1251);
or U5868 (N_5868,N_1466,N_2978);
nand U5869 (N_5869,N_2196,N_1381);
and U5870 (N_5870,N_1524,N_2058);
nor U5871 (N_5871,N_1296,N_2192);
or U5872 (N_5872,N_1335,N_64);
nand U5873 (N_5873,N_610,N_2712);
or U5874 (N_5874,N_54,N_2831);
and U5875 (N_5875,N_2064,N_2678);
and U5876 (N_5876,N_962,N_2413);
nand U5877 (N_5877,N_2160,N_1833);
or U5878 (N_5878,N_827,N_1967);
or U5879 (N_5879,N_1104,N_2241);
or U5880 (N_5880,N_349,N_290);
or U5881 (N_5881,N_1405,N_2027);
nand U5882 (N_5882,N_2331,N_2678);
nor U5883 (N_5883,N_663,N_2310);
and U5884 (N_5884,N_543,N_2130);
or U5885 (N_5885,N_38,N_577);
nor U5886 (N_5886,N_522,N_2951);
nand U5887 (N_5887,N_1861,N_2468);
nor U5888 (N_5888,N_834,N_1914);
or U5889 (N_5889,N_682,N_1200);
and U5890 (N_5890,N_2892,N_2843);
or U5891 (N_5891,N_968,N_2693);
nand U5892 (N_5892,N_722,N_1125);
nor U5893 (N_5893,N_2422,N_2886);
nor U5894 (N_5894,N_2250,N_2969);
and U5895 (N_5895,N_2411,N_615);
or U5896 (N_5896,N_1692,N_1909);
nor U5897 (N_5897,N_1579,N_177);
and U5898 (N_5898,N_1775,N_279);
and U5899 (N_5899,N_2848,N_601);
or U5900 (N_5900,N_2619,N_790);
nor U5901 (N_5901,N_2123,N_2697);
or U5902 (N_5902,N_2601,N_593);
nand U5903 (N_5903,N_2544,N_2794);
and U5904 (N_5904,N_2507,N_2172);
or U5905 (N_5905,N_813,N_915);
nand U5906 (N_5906,N_1221,N_627);
nand U5907 (N_5907,N_2751,N_2897);
xor U5908 (N_5908,N_1005,N_361);
nand U5909 (N_5909,N_2199,N_1472);
or U5910 (N_5910,N_963,N_1865);
and U5911 (N_5911,N_641,N_883);
nor U5912 (N_5912,N_1858,N_1655);
or U5913 (N_5913,N_2574,N_1317);
nor U5914 (N_5914,N_1122,N_2470);
xor U5915 (N_5915,N_52,N_1584);
nor U5916 (N_5916,N_2448,N_2794);
nor U5917 (N_5917,N_672,N_158);
and U5918 (N_5918,N_612,N_72);
and U5919 (N_5919,N_1277,N_2183);
and U5920 (N_5920,N_889,N_2501);
nor U5921 (N_5921,N_486,N_2827);
nand U5922 (N_5922,N_483,N_2117);
nor U5923 (N_5923,N_1807,N_2147);
nand U5924 (N_5924,N_2553,N_2661);
nor U5925 (N_5925,N_662,N_2208);
or U5926 (N_5926,N_156,N_1386);
or U5927 (N_5927,N_658,N_813);
nor U5928 (N_5928,N_2527,N_2382);
and U5929 (N_5929,N_262,N_2389);
and U5930 (N_5930,N_1673,N_399);
and U5931 (N_5931,N_665,N_2911);
or U5932 (N_5932,N_1550,N_762);
or U5933 (N_5933,N_2554,N_1559);
nor U5934 (N_5934,N_1725,N_1022);
nand U5935 (N_5935,N_2447,N_367);
or U5936 (N_5936,N_1275,N_2172);
and U5937 (N_5937,N_133,N_1215);
nand U5938 (N_5938,N_1113,N_1579);
nand U5939 (N_5939,N_711,N_2168);
nand U5940 (N_5940,N_751,N_2844);
nand U5941 (N_5941,N_354,N_1942);
and U5942 (N_5942,N_518,N_208);
nand U5943 (N_5943,N_2352,N_2016);
xnor U5944 (N_5944,N_2309,N_157);
nor U5945 (N_5945,N_190,N_2059);
and U5946 (N_5946,N_2016,N_1634);
and U5947 (N_5947,N_2625,N_1618);
or U5948 (N_5948,N_992,N_1052);
nor U5949 (N_5949,N_2907,N_1167);
and U5950 (N_5950,N_2757,N_2964);
xnor U5951 (N_5951,N_326,N_2340);
or U5952 (N_5952,N_840,N_2835);
nand U5953 (N_5953,N_2230,N_909);
and U5954 (N_5954,N_2296,N_570);
nor U5955 (N_5955,N_2108,N_2323);
nor U5956 (N_5956,N_1969,N_2703);
nor U5957 (N_5957,N_692,N_909);
and U5958 (N_5958,N_990,N_2142);
nor U5959 (N_5959,N_340,N_2895);
nand U5960 (N_5960,N_2253,N_876);
nand U5961 (N_5961,N_2385,N_2327);
or U5962 (N_5962,N_481,N_2020);
nor U5963 (N_5963,N_2394,N_270);
or U5964 (N_5964,N_1727,N_1553);
and U5965 (N_5965,N_923,N_69);
nand U5966 (N_5966,N_224,N_2959);
and U5967 (N_5967,N_1260,N_806);
and U5968 (N_5968,N_1206,N_1381);
xnor U5969 (N_5969,N_544,N_1280);
xnor U5970 (N_5970,N_1809,N_2476);
or U5971 (N_5971,N_483,N_2629);
nand U5972 (N_5972,N_409,N_1326);
and U5973 (N_5973,N_896,N_2571);
and U5974 (N_5974,N_669,N_2490);
or U5975 (N_5975,N_2288,N_2529);
nand U5976 (N_5976,N_2713,N_529);
xor U5977 (N_5977,N_80,N_1026);
nor U5978 (N_5978,N_271,N_462);
nand U5979 (N_5979,N_1134,N_1567);
or U5980 (N_5980,N_1464,N_2797);
and U5981 (N_5981,N_1377,N_958);
nand U5982 (N_5982,N_262,N_512);
nand U5983 (N_5983,N_1193,N_66);
and U5984 (N_5984,N_989,N_2128);
and U5985 (N_5985,N_817,N_1243);
nand U5986 (N_5986,N_1210,N_686);
and U5987 (N_5987,N_823,N_1372);
nor U5988 (N_5988,N_2196,N_1790);
or U5989 (N_5989,N_1751,N_2084);
and U5990 (N_5990,N_285,N_2224);
and U5991 (N_5991,N_1398,N_1299);
or U5992 (N_5992,N_1228,N_1434);
xnor U5993 (N_5993,N_1937,N_1250);
and U5994 (N_5994,N_56,N_2119);
nor U5995 (N_5995,N_2034,N_842);
nand U5996 (N_5996,N_1324,N_2664);
and U5997 (N_5997,N_2699,N_609);
nor U5998 (N_5998,N_407,N_933);
nor U5999 (N_5999,N_2930,N_1381);
and U6000 (N_6000,N_4474,N_3304);
or U6001 (N_6001,N_3441,N_5830);
nor U6002 (N_6002,N_3348,N_5617);
nor U6003 (N_6003,N_3804,N_4435);
or U6004 (N_6004,N_5360,N_3813);
nand U6005 (N_6005,N_5253,N_5128);
or U6006 (N_6006,N_4295,N_3614);
or U6007 (N_6007,N_3930,N_4483);
nand U6008 (N_6008,N_5153,N_4487);
and U6009 (N_6009,N_3091,N_3186);
nor U6010 (N_6010,N_3648,N_3159);
and U6011 (N_6011,N_4739,N_4714);
and U6012 (N_6012,N_5117,N_3965);
and U6013 (N_6013,N_5505,N_5653);
or U6014 (N_6014,N_4137,N_5004);
or U6015 (N_6015,N_5196,N_4785);
nor U6016 (N_6016,N_4448,N_4783);
nand U6017 (N_6017,N_4215,N_5036);
or U6018 (N_6018,N_5813,N_3279);
nor U6019 (N_6019,N_3633,N_4471);
xnor U6020 (N_6020,N_4498,N_3995);
or U6021 (N_6021,N_4050,N_5557);
nand U6022 (N_6022,N_5787,N_4475);
or U6023 (N_6023,N_3410,N_5393);
nand U6024 (N_6024,N_3577,N_5355);
nand U6025 (N_6025,N_5510,N_3966);
or U6026 (N_6026,N_3696,N_4259);
and U6027 (N_6027,N_4890,N_4712);
nand U6028 (N_6028,N_3097,N_5678);
xor U6029 (N_6029,N_5046,N_4367);
nor U6030 (N_6030,N_5127,N_4465);
or U6031 (N_6031,N_4132,N_3613);
nor U6032 (N_6032,N_4624,N_5332);
or U6033 (N_6033,N_4638,N_5189);
and U6034 (N_6034,N_5842,N_5151);
nand U6035 (N_6035,N_5862,N_4901);
nor U6036 (N_6036,N_4514,N_3865);
and U6037 (N_6037,N_4942,N_3043);
or U6038 (N_6038,N_3503,N_4679);
or U6039 (N_6039,N_5186,N_3058);
and U6040 (N_6040,N_4711,N_3364);
nand U6041 (N_6041,N_4315,N_5331);
nor U6042 (N_6042,N_4470,N_5583);
nand U6043 (N_6043,N_4781,N_3877);
and U6044 (N_6044,N_4303,N_4113);
and U6045 (N_6045,N_3333,N_4366);
nor U6046 (N_6046,N_4911,N_4799);
and U6047 (N_6047,N_5069,N_4904);
nand U6048 (N_6048,N_4128,N_5758);
nand U6049 (N_6049,N_3164,N_4899);
nor U6050 (N_6050,N_5742,N_3079);
or U6051 (N_6051,N_4539,N_5042);
nor U6052 (N_6052,N_3303,N_5792);
nand U6053 (N_6053,N_5957,N_4531);
or U6054 (N_6054,N_3690,N_3431);
nand U6055 (N_6055,N_5696,N_3928);
and U6056 (N_6056,N_5750,N_4232);
nand U6057 (N_6057,N_5741,N_5118);
or U6058 (N_6058,N_5348,N_4306);
nand U6059 (N_6059,N_4895,N_3429);
nor U6060 (N_6060,N_5287,N_3669);
xnor U6061 (N_6061,N_5943,N_3171);
or U6062 (N_6062,N_3347,N_3387);
and U6063 (N_6063,N_4385,N_4505);
nand U6064 (N_6064,N_5652,N_3760);
and U6065 (N_6065,N_3045,N_3775);
xor U6066 (N_6066,N_3184,N_3548);
nor U6067 (N_6067,N_4497,N_4844);
and U6068 (N_6068,N_5575,N_4089);
nand U6069 (N_6069,N_4064,N_4863);
nor U6070 (N_6070,N_5412,N_3415);
nor U6071 (N_6071,N_5834,N_3353);
xor U6072 (N_6072,N_5887,N_3562);
or U6073 (N_6073,N_3601,N_5686);
nor U6074 (N_6074,N_5033,N_5804);
or U6075 (N_6075,N_5316,N_5717);
or U6076 (N_6076,N_3893,N_3898);
and U6077 (N_6077,N_5755,N_5642);
and U6078 (N_6078,N_3486,N_4707);
nand U6079 (N_6079,N_3419,N_3454);
nand U6080 (N_6080,N_4380,N_5718);
and U6081 (N_6081,N_4496,N_5247);
or U6082 (N_6082,N_3863,N_4946);
nor U6083 (N_6083,N_3367,N_4187);
xor U6084 (N_6084,N_5725,N_5070);
nor U6085 (N_6085,N_3909,N_3497);
xnor U6086 (N_6086,N_3447,N_4406);
nand U6087 (N_6087,N_5109,N_5697);
nand U6088 (N_6088,N_4544,N_5278);
nor U6089 (N_6089,N_5378,N_4851);
nor U6090 (N_6090,N_4114,N_5384);
nor U6091 (N_6091,N_4750,N_3942);
nand U6092 (N_6092,N_5727,N_5936);
nor U6093 (N_6093,N_4323,N_4481);
nor U6094 (N_6094,N_4980,N_3940);
or U6095 (N_6095,N_5322,N_5567);
and U6096 (N_6096,N_5212,N_3978);
or U6097 (N_6097,N_5334,N_5876);
nand U6098 (N_6098,N_4680,N_4871);
or U6099 (N_6099,N_3744,N_3133);
nand U6100 (N_6100,N_5641,N_5220);
nand U6101 (N_6101,N_3708,N_4825);
and U6102 (N_6102,N_5207,N_4964);
nor U6103 (N_6103,N_3688,N_5720);
nand U6104 (N_6104,N_5132,N_3076);
nor U6105 (N_6105,N_4422,N_4099);
nand U6106 (N_6106,N_4070,N_3717);
xnor U6107 (N_6107,N_3626,N_3567);
or U6108 (N_6108,N_3011,N_4381);
or U6109 (N_6109,N_3163,N_4744);
or U6110 (N_6110,N_3662,N_5194);
nand U6111 (N_6111,N_5131,N_5877);
and U6112 (N_6112,N_3561,N_5781);
and U6113 (N_6113,N_4637,N_4996);
or U6114 (N_6114,N_4670,N_4379);
or U6115 (N_6115,N_5875,N_4408);
or U6116 (N_6116,N_4865,N_4704);
xnor U6117 (N_6117,N_3212,N_3014);
nand U6118 (N_6118,N_4566,N_5238);
or U6119 (N_6119,N_3802,N_5704);
or U6120 (N_6120,N_4508,N_5476);
and U6121 (N_6121,N_4725,N_5722);
nor U6122 (N_6122,N_5739,N_4433);
or U6123 (N_6123,N_3094,N_3983);
nand U6124 (N_6124,N_3559,N_5285);
and U6125 (N_6125,N_3388,N_5255);
nand U6126 (N_6126,N_3224,N_4226);
nor U6127 (N_6127,N_4374,N_3569);
nor U6128 (N_6128,N_3025,N_4488);
nor U6129 (N_6129,N_5065,N_3709);
or U6130 (N_6130,N_4960,N_4933);
xor U6131 (N_6131,N_5283,N_4296);
or U6132 (N_6132,N_5863,N_4082);
nand U6133 (N_6133,N_5607,N_5568);
and U6134 (N_6134,N_5462,N_5942);
or U6135 (N_6135,N_5879,N_3738);
xnor U6136 (N_6136,N_5346,N_4741);
nor U6137 (N_6137,N_4956,N_3330);
nand U6138 (N_6138,N_5410,N_5856);
and U6139 (N_6139,N_5888,N_4558);
nand U6140 (N_6140,N_3193,N_4390);
nand U6141 (N_6141,N_4044,N_3361);
and U6142 (N_6142,N_3927,N_3439);
or U6143 (N_6143,N_4004,N_5363);
or U6144 (N_6144,N_3147,N_4138);
nor U6145 (N_6145,N_3836,N_4131);
and U6146 (N_6146,N_4772,N_5963);
and U6147 (N_6147,N_5602,N_5681);
nor U6148 (N_6148,N_4127,N_5313);
and U6149 (N_6149,N_3023,N_4611);
and U6150 (N_6150,N_3882,N_4063);
or U6151 (N_6151,N_5839,N_5330);
nor U6152 (N_6152,N_4376,N_4605);
nand U6153 (N_6153,N_5992,N_5689);
and U6154 (N_6154,N_4009,N_4349);
nor U6155 (N_6155,N_4212,N_5794);
and U6156 (N_6156,N_5265,N_3903);
and U6157 (N_6157,N_5647,N_5685);
nand U6158 (N_6158,N_4421,N_3313);
or U6159 (N_6159,N_4446,N_4631);
nor U6160 (N_6160,N_3950,N_3967);
or U6161 (N_6161,N_5587,N_4789);
xnor U6162 (N_6162,N_4565,N_4934);
or U6163 (N_6163,N_5045,N_3495);
or U6164 (N_6164,N_5983,N_3945);
xor U6165 (N_6165,N_5236,N_3956);
nor U6166 (N_6166,N_4540,N_4582);
nor U6167 (N_6167,N_3484,N_3565);
nor U6168 (N_6168,N_5625,N_3739);
xor U6169 (N_6169,N_3203,N_5086);
xor U6170 (N_6170,N_5053,N_5616);
xor U6171 (N_6171,N_5063,N_5408);
nor U6172 (N_6172,N_3753,N_3478);
or U6173 (N_6173,N_4104,N_3161);
and U6174 (N_6174,N_3496,N_5555);
and U6175 (N_6175,N_4142,N_4849);
or U6176 (N_6176,N_5754,N_3434);
nand U6177 (N_6177,N_4102,N_5397);
or U6178 (N_6178,N_4165,N_4231);
and U6179 (N_6179,N_5209,N_5262);
nand U6180 (N_6180,N_4860,N_4893);
and U6181 (N_6181,N_5039,N_5263);
nand U6182 (N_6182,N_4333,N_4067);
xnor U6183 (N_6183,N_4297,N_4793);
nand U6184 (N_6184,N_3047,N_4814);
xor U6185 (N_6185,N_3911,N_5179);
or U6186 (N_6186,N_4676,N_5048);
or U6187 (N_6187,N_4427,N_3336);
or U6188 (N_6188,N_4503,N_4103);
or U6189 (N_6189,N_3174,N_5318);
nand U6190 (N_6190,N_3078,N_3343);
nand U6191 (N_6191,N_3964,N_5541);
and U6192 (N_6192,N_4669,N_4019);
nor U6193 (N_6193,N_5810,N_5841);
or U6194 (N_6194,N_5141,N_4346);
and U6195 (N_6195,N_4199,N_4755);
nand U6196 (N_6196,N_5517,N_4155);
nand U6197 (N_6197,N_4800,N_4641);
or U6198 (N_6198,N_4843,N_4920);
and U6199 (N_6199,N_3469,N_5581);
and U6200 (N_6200,N_4726,N_3056);
nor U6201 (N_6201,N_4154,N_3460);
or U6202 (N_6202,N_4358,N_3425);
nor U6203 (N_6203,N_5747,N_3102);
nor U6204 (N_6204,N_5225,N_4902);
nand U6205 (N_6205,N_5114,N_3449);
xor U6206 (N_6206,N_3229,N_5231);
and U6207 (N_6207,N_3187,N_5105);
nor U6208 (N_6208,N_3602,N_5799);
or U6209 (N_6209,N_3675,N_3947);
or U6210 (N_6210,N_3477,N_4411);
nand U6211 (N_6211,N_3828,N_4207);
xor U6212 (N_6212,N_5950,N_3665);
or U6213 (N_6213,N_5564,N_4889);
nand U6214 (N_6214,N_5767,N_3618);
and U6215 (N_6215,N_4667,N_5972);
and U6216 (N_6216,N_4754,N_3612);
nor U6217 (N_6217,N_4083,N_5480);
xor U6218 (N_6218,N_4938,N_3914);
nand U6219 (N_6219,N_4047,N_4925);
and U6220 (N_6220,N_5562,N_4198);
or U6221 (N_6221,N_3158,N_3374);
xor U6222 (N_6222,N_4491,N_5622);
nor U6223 (N_6223,N_5143,N_4195);
or U6224 (N_6224,N_3743,N_5391);
nand U6225 (N_6225,N_3890,N_4357);
or U6226 (N_6226,N_4947,N_3100);
xor U6227 (N_6227,N_4106,N_3924);
or U6228 (N_6228,N_3116,N_4819);
nand U6229 (N_6229,N_5650,N_4576);
and U6230 (N_6230,N_5561,N_3906);
and U6231 (N_6231,N_5107,N_5292);
xnor U6232 (N_6232,N_5599,N_5379);
and U6233 (N_6233,N_4213,N_3029);
and U6234 (N_6234,N_3476,N_4857);
and U6235 (N_6235,N_3634,N_4500);
nand U6236 (N_6236,N_3329,N_5244);
and U6237 (N_6237,N_5481,N_4268);
nand U6238 (N_6238,N_4484,N_4413);
nor U6239 (N_6239,N_5094,N_3571);
and U6240 (N_6240,N_4175,N_3642);
or U6241 (N_6241,N_3302,N_5882);
nand U6242 (N_6242,N_5276,N_5881);
or U6243 (N_6243,N_5901,N_5190);
nand U6244 (N_6244,N_4324,N_5509);
or U6245 (N_6245,N_3574,N_3166);
and U6246 (N_6246,N_4763,N_4267);
and U6247 (N_6247,N_3710,N_4469);
nand U6248 (N_6248,N_5277,N_5203);
nor U6249 (N_6249,N_4482,N_4093);
and U6250 (N_6250,N_5089,N_4197);
or U6251 (N_6251,N_3766,N_4629);
and U6252 (N_6252,N_5612,N_4405);
nor U6253 (N_6253,N_5266,N_5826);
or U6254 (N_6254,N_5026,N_3283);
and U6255 (N_6255,N_5608,N_4094);
nor U6256 (N_6256,N_4630,N_4943);
and U6257 (N_6257,N_3630,N_5748);
or U6258 (N_6258,N_4628,N_3385);
or U6259 (N_6259,N_3500,N_3472);
xor U6260 (N_6260,N_3941,N_3923);
or U6261 (N_6261,N_4869,N_3190);
nor U6262 (N_6262,N_3705,N_3922);
or U6263 (N_6263,N_4115,N_5746);
or U6264 (N_6264,N_4988,N_4150);
or U6265 (N_6265,N_3145,N_3216);
and U6266 (N_6266,N_3383,N_3122);
nand U6267 (N_6267,N_3134,N_5445);
or U6268 (N_6268,N_3993,N_3197);
nand U6269 (N_6269,N_3232,N_4972);
and U6270 (N_6270,N_3480,N_3272);
nand U6271 (N_6271,N_4332,N_5252);
nor U6272 (N_6272,N_5496,N_3342);
nand U6273 (N_6273,N_3390,N_5631);
nor U6274 (N_6274,N_3632,N_4662);
nand U6275 (N_6275,N_5431,N_3889);
and U6276 (N_6276,N_5035,N_4135);
nor U6277 (N_6277,N_3270,N_5520);
and U6278 (N_6278,N_3711,N_4745);
nor U6279 (N_6279,N_5645,N_5289);
or U6280 (N_6280,N_4770,N_3445);
nor U6281 (N_6281,N_5310,N_3511);
or U6282 (N_6282,N_4782,N_4610);
and U6283 (N_6283,N_5728,N_5020);
or U6284 (N_6284,N_4157,N_3243);
and U6285 (N_6285,N_4329,N_3057);
nand U6286 (N_6286,N_5084,N_4583);
and U6287 (N_6287,N_3022,N_5846);
nor U6288 (N_6288,N_5494,N_5890);
or U6289 (N_6289,N_5451,N_4042);
and U6290 (N_6290,N_5130,N_5405);
or U6291 (N_6291,N_3671,N_5155);
xor U6292 (N_6292,N_4119,N_4509);
and U6293 (N_6293,N_4798,N_4459);
nor U6294 (N_6294,N_3845,N_3332);
nor U6295 (N_6295,N_4118,N_3211);
nor U6296 (N_6296,N_3098,N_4519);
nor U6297 (N_6297,N_5695,N_3370);
or U6298 (N_6298,N_3532,N_5730);
xor U6299 (N_6299,N_4824,N_5140);
or U6300 (N_6300,N_5521,N_5549);
and U6301 (N_6301,N_4437,N_5396);
nand U6302 (N_6302,N_3829,N_5623);
or U6303 (N_6303,N_3595,N_3801);
or U6304 (N_6304,N_3809,N_5579);
nand U6305 (N_6305,N_3412,N_5757);
and U6306 (N_6306,N_3653,N_4919);
nand U6307 (N_6307,N_4037,N_4997);
nand U6308 (N_6308,N_4600,N_3432);
nand U6309 (N_6309,N_3200,N_3723);
and U6310 (N_6310,N_4139,N_4816);
nor U6311 (N_6311,N_5734,N_5492);
nor U6312 (N_6312,N_4233,N_5914);
or U6313 (N_6313,N_3408,N_5210);
and U6314 (N_6314,N_4691,N_3470);
nand U6315 (N_6315,N_3868,N_4905);
nor U6316 (N_6316,N_4318,N_5110);
and U6317 (N_6317,N_3312,N_4794);
nor U6318 (N_6318,N_3202,N_4204);
nor U6319 (N_6319,N_5336,N_5670);
or U6320 (N_6320,N_3162,N_5075);
or U6321 (N_6321,N_4144,N_5947);
and U6322 (N_6322,N_5241,N_5347);
nor U6323 (N_6323,N_3101,N_3720);
and U6324 (N_6324,N_3126,N_4697);
or U6325 (N_6325,N_5796,N_3450);
nor U6326 (N_6326,N_4924,N_5638);
and U6327 (N_6327,N_4426,N_4034);
and U6328 (N_6328,N_4492,N_4856);
xor U6329 (N_6329,N_5774,N_3583);
nor U6330 (N_6330,N_4549,N_3958);
nand U6331 (N_6331,N_5539,N_5953);
and U6332 (N_6332,N_5303,N_5368);
and U6333 (N_6333,N_5420,N_4577);
and U6334 (N_6334,N_5937,N_5604);
nor U6335 (N_6335,N_5426,N_3615);
and U6336 (N_6336,N_3522,N_4211);
nand U6337 (N_6337,N_5603,N_4249);
nor U6338 (N_6338,N_5495,N_5392);
and U6339 (N_6339,N_5924,N_4216);
nor U6340 (N_6340,N_4423,N_5300);
nor U6341 (N_6341,N_5074,N_3714);
and U6342 (N_6342,N_3253,N_3780);
nor U6343 (N_6343,N_4049,N_5161);
or U6344 (N_6344,N_3555,N_3680);
or U6345 (N_6345,N_4952,N_3859);
or U6346 (N_6346,N_3579,N_5949);
or U6347 (N_6347,N_3526,N_4161);
or U6348 (N_6348,N_4971,N_3027);
or U6349 (N_6349,N_5524,N_3443);
or U6350 (N_6350,N_5955,N_5665);
nor U6351 (N_6351,N_4591,N_4732);
or U6352 (N_6352,N_4285,N_5580);
or U6353 (N_6353,N_4693,N_5129);
or U6354 (N_6354,N_3015,N_4903);
nor U6355 (N_6355,N_5227,N_4340);
nand U6356 (N_6356,N_5951,N_3871);
or U6357 (N_6357,N_4181,N_3883);
nor U6358 (N_6358,N_3436,N_5658);
or U6359 (N_6359,N_3654,N_4708);
nor U6360 (N_6360,N_4359,N_4145);
and U6361 (N_6361,N_5553,N_4317);
nor U6362 (N_6362,N_3123,N_3799);
nand U6363 (N_6363,N_4438,N_5744);
or U6364 (N_6364,N_5025,N_5546);
and U6365 (N_6365,N_4927,N_4253);
nor U6366 (N_6366,N_5167,N_4649);
or U6367 (N_6367,N_3108,N_4271);
or U6368 (N_6368,N_4516,N_4289);
nor U6369 (N_6369,N_5797,N_3844);
or U6370 (N_6370,N_5596,N_3619);
or U6371 (N_6371,N_3345,N_4372);
and U6372 (N_6372,N_5789,N_5526);
xnor U6373 (N_6373,N_4573,N_3598);
or U6374 (N_6374,N_3444,N_3386);
nor U6375 (N_6375,N_3538,N_5011);
nor U6376 (N_6376,N_5133,N_4721);
and U6377 (N_6377,N_5569,N_3936);
or U6378 (N_6378,N_4767,N_4056);
or U6379 (N_6379,N_4524,N_5712);
and U6380 (N_6380,N_3407,N_5613);
nand U6381 (N_6381,N_3248,N_3349);
nand U6382 (N_6382,N_3886,N_5905);
nand U6383 (N_6383,N_4717,N_5869);
nand U6384 (N_6384,N_4547,N_4014);
nor U6385 (N_6385,N_3510,N_5113);
nor U6386 (N_6386,N_5068,N_3787);
nor U6387 (N_6387,N_3918,N_5700);
nor U6388 (N_6388,N_4961,N_3933);
or U6389 (N_6389,N_5447,N_4986);
nand U6390 (N_6390,N_3404,N_4888);
and U6391 (N_6391,N_3069,N_5441);
nor U6392 (N_6392,N_3119,N_3892);
xor U6393 (N_6393,N_3396,N_4148);
nor U6394 (N_6394,N_4822,N_5424);
or U6395 (N_6395,N_4153,N_5605);
and U6396 (N_6396,N_4829,N_3221);
nor U6397 (N_6397,N_4360,N_3533);
xor U6398 (N_6398,N_4586,N_4223);
nor U6399 (N_6399,N_5199,N_4559);
nand U6400 (N_6400,N_4238,N_4832);
or U6401 (N_6401,N_5552,N_4894);
nand U6402 (N_6402,N_5958,N_4040);
or U6403 (N_6403,N_5464,N_3490);
or U6404 (N_6404,N_3725,N_3352);
nor U6405 (N_6405,N_3563,N_4926);
nor U6406 (N_6406,N_5907,N_3136);
xnor U6407 (N_6407,N_5537,N_5073);
nor U6408 (N_6408,N_4369,N_4339);
xor U6409 (N_6409,N_3769,N_5077);
and U6410 (N_6410,N_4328,N_3188);
or U6411 (N_6411,N_3062,N_5425);
and U6412 (N_6412,N_4736,N_4476);
nor U6413 (N_6413,N_3120,N_3132);
nand U6414 (N_6414,N_4293,N_3849);
nor U6415 (N_6415,N_5216,N_3453);
nand U6416 (N_6416,N_5427,N_3660);
or U6417 (N_6417,N_5661,N_5899);
or U6418 (N_6418,N_3597,N_5988);
and U6419 (N_6419,N_4337,N_4092);
xor U6420 (N_6420,N_3182,N_4257);
nor U6421 (N_6421,N_3808,N_3647);
nor U6422 (N_6422,N_5691,N_5801);
or U6423 (N_6423,N_4111,N_4244);
xnor U6424 (N_6424,N_4478,N_4298);
nor U6425 (N_6425,N_5382,N_4310);
and U6426 (N_6426,N_5687,N_5506);
nor U6427 (N_6427,N_5482,N_4853);
nor U6428 (N_6428,N_5745,N_5099);
nor U6429 (N_6429,N_4391,N_3999);
nand U6430 (N_6430,N_5578,N_5032);
and U6431 (N_6431,N_3196,N_3381);
or U6432 (N_6432,N_3734,N_4201);
and U6433 (N_6433,N_5007,N_5267);
or U6434 (N_6434,N_5594,N_5223);
nand U6435 (N_6435,N_3296,N_4765);
nor U6436 (N_6436,N_3281,N_5651);
xor U6437 (N_6437,N_5002,N_3695);
nor U6438 (N_6438,N_4909,N_4395);
and U6439 (N_6439,N_4490,N_3273);
and U6440 (N_6440,N_5508,N_4615);
nand U6441 (N_6441,N_5772,N_5814);
or U6442 (N_6442,N_4659,N_4959);
xnor U6443 (N_6443,N_3608,N_3875);
and U6444 (N_6444,N_4931,N_5184);
and U6445 (N_6445,N_3327,N_4156);
and U6446 (N_6446,N_5591,N_3540);
or U6447 (N_6447,N_3001,N_4341);
nand U6448 (N_6448,N_3085,N_5761);
and U6449 (N_6449,N_5023,N_4344);
or U6450 (N_6450,N_3254,N_3834);
nand U6451 (N_6451,N_4862,N_3527);
nand U6452 (N_6452,N_3068,N_5824);
nor U6453 (N_6453,N_4068,N_3240);
xor U6454 (N_6454,N_3019,N_4643);
or U6455 (N_6455,N_3682,N_5369);
or U6456 (N_6456,N_3316,N_5335);
nand U6457 (N_6457,N_5430,N_3721);
nand U6458 (N_6458,N_4999,N_5442);
nand U6459 (N_6459,N_4906,N_4363);
nand U6460 (N_6460,N_4425,N_3908);
or U6461 (N_6461,N_5654,N_3806);
nor U6462 (N_6462,N_5078,N_3587);
nor U6463 (N_6463,N_4236,N_4694);
nor U6464 (N_6464,N_4400,N_4720);
nand U6465 (N_6465,N_3811,N_5095);
nand U6466 (N_6466,N_3237,N_4907);
nor U6467 (N_6467,N_3409,N_4731);
nand U6468 (N_6468,N_5635,N_5915);
nand U6469 (N_6469,N_5843,N_3797);
nand U6470 (N_6470,N_3896,N_3090);
nand U6471 (N_6471,N_4075,N_3915);
and U6472 (N_6472,N_5922,N_4684);
nor U6473 (N_6473,N_3290,N_4321);
or U6474 (N_6474,N_5453,N_3997);
nand U6475 (N_6475,N_5903,N_4970);
and U6476 (N_6476,N_4787,N_5411);
and U6477 (N_6477,N_5719,N_4878);
and U6478 (N_6478,N_4748,N_5386);
nor U6479 (N_6479,N_3866,N_5636);
nor U6480 (N_6480,N_3139,N_5059);
and U6481 (N_6481,N_3640,N_5294);
nor U6482 (N_6482,N_5698,N_4668);
or U6483 (N_6483,N_5067,N_4414);
nor U6484 (N_6484,N_4619,N_4866);
xor U6485 (N_6485,N_4022,N_4282);
or U6486 (N_6486,N_4815,N_3902);
nand U6487 (N_6487,N_3009,N_4673);
and U6488 (N_6488,N_4561,N_4170);
and U6489 (N_6489,N_5543,N_5204);
xnor U6490 (N_6490,N_5234,N_5174);
nand U6491 (N_6491,N_3021,N_3391);
xor U6492 (N_6492,N_5780,N_3543);
nand U6493 (N_6493,N_4283,N_3050);
and U6494 (N_6494,N_4277,N_3125);
nand U6495 (N_6495,N_4290,N_5560);
nor U6496 (N_6496,N_3039,N_5080);
nor U6497 (N_6497,N_5864,N_3716);
nor U6498 (N_6498,N_4859,N_3641);
or U6499 (N_6499,N_5768,N_3261);
and U6500 (N_6500,N_3250,N_4564);
nor U6501 (N_6501,N_3402,N_5434);
nand U6502 (N_6502,N_3814,N_3437);
xnor U6503 (N_6503,N_5173,N_3389);
and U6504 (N_6504,N_4912,N_4982);
or U6505 (N_6505,N_4002,N_4718);
or U6506 (N_6506,N_5554,N_4046);
nand U6507 (N_6507,N_4795,N_5548);
and U6508 (N_6508,N_4035,N_5971);
nor U6509 (N_6509,N_4831,N_3362);
nor U6510 (N_6510,N_5043,N_3670);
and U6511 (N_6511,N_3698,N_4008);
xor U6512 (N_6512,N_3268,N_5333);
nor U6513 (N_6513,N_4203,N_3028);
or U6514 (N_6514,N_5666,N_4003);
or U6515 (N_6515,N_4287,N_5597);
and U6516 (N_6516,N_3643,N_3646);
nor U6517 (N_6517,N_5868,N_5051);
and U6518 (N_6518,N_4685,N_5667);
or U6519 (N_6519,N_5443,N_3610);
and U6520 (N_6520,N_4041,N_3718);
nand U6521 (N_6521,N_4458,N_4214);
and U6522 (N_6522,N_5230,N_4243);
or U6523 (N_6523,N_4171,N_3502);
or U6524 (N_6524,N_5126,N_3117);
nand U6525 (N_6525,N_3118,N_3722);
and U6526 (N_6526,N_5469,N_3244);
or U6527 (N_6527,N_4634,N_5872);
and U6528 (N_6528,N_5454,N_4626);
xnor U6529 (N_6529,N_4827,N_3550);
nand U6530 (N_6530,N_3631,N_5802);
nand U6531 (N_6531,N_3524,N_5101);
nor U6532 (N_6532,N_4644,N_4929);
and U6533 (N_6533,N_5291,N_4117);
or U6534 (N_6534,N_4987,N_4266);
nor U6535 (N_6535,N_3623,N_3777);
nand U6536 (N_6536,N_4584,N_4526);
or U6537 (N_6537,N_4167,N_5836);
nor U6538 (N_6538,N_5372,N_4601);
and U6539 (N_6539,N_3588,N_4780);
or U6540 (N_6540,N_5980,N_3063);
nand U6541 (N_6541,N_4695,N_4246);
nor U6542 (N_6542,N_3099,N_4724);
and U6543 (N_6543,N_5782,N_3843);
xnor U6544 (N_6544,N_5900,N_4292);
or U6545 (N_6545,N_4826,N_5488);
nor U6546 (N_6546,N_5895,N_5640);
and U6547 (N_6547,N_5996,N_5528);
nand U6548 (N_6548,N_4045,N_3399);
or U6549 (N_6549,N_5182,N_4535);
nor U6550 (N_6550,N_4939,N_4219);
or U6551 (N_6551,N_4702,N_3241);
or U6552 (N_6552,N_5460,N_5307);
or U6553 (N_6553,N_3937,N_5465);
nor U6554 (N_6554,N_4896,N_4051);
and U6555 (N_6555,N_4055,N_3276);
nand U6556 (N_6556,N_5222,N_3054);
and U6557 (N_6557,N_3128,N_4221);
nor U6558 (N_6558,N_3397,N_3573);
nor U6559 (N_6559,N_3005,N_3673);
nand U6560 (N_6560,N_3895,N_5925);
xnor U6561 (N_6561,N_4120,N_3055);
or U6562 (N_6562,N_4834,N_5643);
nand U6563 (N_6563,N_3649,N_5500);
nand U6564 (N_6564,N_3269,N_5884);
and U6565 (N_6565,N_3585,N_5713);
or U6566 (N_6566,N_4842,N_5848);
nand U6567 (N_6567,N_4602,N_3984);
nor U6568 (N_6568,N_4749,N_3521);
nand U6569 (N_6569,N_3850,N_4313);
or U6570 (N_6570,N_3061,N_5817);
and U6571 (N_6571,N_5891,N_5437);
nand U6572 (N_6572,N_5703,N_5735);
or U6573 (N_6573,N_3406,N_4963);
nor U6574 (N_6574,N_5243,N_4312);
or U6575 (N_6575,N_4716,N_4122);
nor U6576 (N_6576,N_5245,N_3427);
nand U6577 (N_6577,N_4820,N_3030);
or U6578 (N_6578,N_4553,N_4527);
or U6579 (N_6579,N_4095,N_4791);
nor U6580 (N_6580,N_4090,N_5964);
and U6581 (N_6581,N_3838,N_5851);
and U6582 (N_6582,N_3037,N_5233);
xnor U6583 (N_6583,N_4882,N_3700);
and U6584 (N_6584,N_4116,N_4151);
nor U6585 (N_6585,N_5047,N_4998);
nand U6586 (N_6586,N_3201,N_4241);
and U6587 (N_6587,N_4392,N_5908);
or U6588 (N_6588,N_5979,N_3291);
nand U6589 (N_6589,N_5450,N_4053);
nand U6590 (N_6590,N_3735,N_5058);
xnor U6591 (N_6591,N_5913,N_3205);
nand U6592 (N_6592,N_4623,N_3259);
or U6593 (N_6593,N_4883,N_5999);
nor U6594 (N_6594,N_4764,N_5064);
xnor U6595 (N_6595,N_5191,N_5987);
nand U6596 (N_6596,N_4345,N_5152);
or U6597 (N_6597,N_3059,N_5281);
nand U6598 (N_6598,N_3463,N_5022);
xor U6599 (N_6599,N_5028,N_3236);
and U6600 (N_6600,N_3572,N_4812);
nand U6601 (N_6601,N_4133,N_3731);
or U6602 (N_6602,N_4548,N_5024);
xor U6603 (N_6603,N_5590,N_4830);
nor U6604 (N_6604,N_5166,N_4675);
xor U6605 (N_6605,N_5135,N_3204);
nor U6606 (N_6606,N_5504,N_5984);
nor U6607 (N_6607,N_3403,N_3853);
nand U6608 (N_6608,N_4280,N_3916);
xnor U6609 (N_6609,N_4202,N_4880);
nand U6610 (N_6610,N_5345,N_5898);
and U6611 (N_6611,N_5620,N_3963);
or U6612 (N_6612,N_5847,N_4525);
or U6613 (N_6613,N_3894,N_5974);
nand U6614 (N_6614,N_3144,N_3925);
xor U6615 (N_6615,N_5235,N_4778);
or U6616 (N_6616,N_4706,N_3242);
and U6617 (N_6617,N_3366,N_3376);
and U6618 (N_6618,N_5349,N_3249);
or U6619 (N_6619,N_5271,N_4627);
nand U6620 (N_6620,N_3135,N_3073);
nor U6621 (N_6621,N_4958,N_3324);
nand U6622 (N_6622,N_3976,N_4529);
or U6623 (N_6623,N_5100,N_4384);
xor U6624 (N_6624,N_3727,N_5072);
or U6625 (N_6625,N_5928,N_4424);
and U6626 (N_6626,N_4461,N_3537);
nand U6627 (N_6627,N_4587,N_4788);
nor U6628 (N_6628,N_5493,N_3635);
or U6629 (N_6629,N_4773,N_3339);
and U6630 (N_6630,N_5994,N_3611);
nand U6631 (N_6631,N_5498,N_5502);
nand U6632 (N_6632,N_5675,N_4072);
or U6633 (N_6633,N_5513,N_3346);
nor U6634 (N_6634,N_3095,N_5455);
and U6635 (N_6635,N_3932,N_5816);
nor U6636 (N_6636,N_3002,N_4674);
or U6637 (N_6637,N_5061,N_4797);
nor U6638 (N_6638,N_3786,N_3740);
xnor U6639 (N_6639,N_5282,N_3757);
nand U6640 (N_6640,N_4511,N_3818);
or U6641 (N_6641,N_5822,N_5296);
nand U6642 (N_6642,N_4242,N_5315);
or U6643 (N_6643,N_3901,N_3382);
nand U6644 (N_6644,N_5993,N_4079);
or U6645 (N_6645,N_5340,N_3552);
and U6646 (N_6646,N_3358,N_5736);
and U6647 (N_6647,N_4356,N_3493);
nor U6648 (N_6648,N_4228,N_5663);
nor U6649 (N_6649,N_4149,N_3617);
nand U6650 (N_6650,N_4071,N_5589);
or U6651 (N_6651,N_4364,N_3515);
nand U6652 (N_6652,N_5395,N_3729);
nand U6653 (N_6653,N_3862,N_4723);
and U6654 (N_6654,N_4984,N_4010);
or U6655 (N_6655,N_5407,N_5337);
or U6656 (N_6656,N_4088,N_3114);
nor U6657 (N_6657,N_5503,N_3426);
or U6658 (N_6658,N_4599,N_5142);
or U6659 (N_6659,N_3309,N_4451);
nor U6660 (N_6660,N_3354,N_3481);
or U6661 (N_6661,N_3560,N_3951);
and U6662 (N_6662,N_3888,N_5610);
or U6663 (N_6663,N_5812,N_4838);
and U6664 (N_6664,N_4568,N_5705);
nand U6665 (N_6665,N_3170,N_4900);
or U6666 (N_6666,N_3065,N_3049);
nand U6667 (N_6667,N_4809,N_4538);
nor U6668 (N_6668,N_4362,N_3067);
nor U6669 (N_6669,N_5614,N_5962);
nor U6670 (N_6670,N_5121,N_3487);
nand U6671 (N_6671,N_5793,N_4993);
nor U6672 (N_6672,N_5096,N_3935);
and U6673 (N_6673,N_5585,N_4463);
nor U6674 (N_6674,N_5601,N_4528);
nand U6675 (N_6675,N_3299,N_4658);
and U6676 (N_6676,N_4368,N_5637);
nor U6677 (N_6677,N_3684,N_3713);
nand U6678 (N_6678,N_4330,N_4311);
and U6679 (N_6679,N_3507,N_3322);
and U6680 (N_6680,N_5260,N_5342);
or U6681 (N_6681,N_5224,N_5997);
or U6682 (N_6682,N_5400,N_3060);
nand U6683 (N_6683,N_4689,N_4141);
nor U6684 (N_6684,N_5297,N_5860);
or U6685 (N_6685,N_4976,N_5619);
nor U6686 (N_6686,N_4172,N_4123);
and U6687 (N_6687,N_4743,N_3208);
nand U6688 (N_6688,N_4234,N_5102);
nand U6689 (N_6689,N_4733,N_4567);
nor U6690 (N_6690,N_4940,N_3266);
and U6691 (N_6691,N_5423,N_3689);
xnor U6692 (N_6692,N_4060,N_3827);
nor U6693 (N_6693,N_3131,N_5732);
and U6694 (N_6694,N_4682,N_3467);
or U6695 (N_6695,N_3977,N_4639);
nor U6696 (N_6696,N_5467,N_5966);
and U6697 (N_6697,N_4664,N_4728);
and U6698 (N_6698,N_5786,N_5572);
or U6699 (N_6699,N_4261,N_3151);
nand U6700 (N_6700,N_3031,N_5677);
nand U6701 (N_6701,N_4715,N_3938);
nand U6702 (N_6702,N_4126,N_3629);
nand U6703 (N_6703,N_4562,N_3194);
xnor U6704 (N_6704,N_5375,N_3985);
nor U6705 (N_6705,N_4608,N_4342);
and U6706 (N_6706,N_5009,N_3275);
nand U6707 (N_6707,N_3880,N_3255);
or U6708 (N_6708,N_3774,N_3536);
nor U6709 (N_6709,N_3466,N_3413);
or U6710 (N_6710,N_3474,N_5081);
nor U6711 (N_6711,N_4351,N_4386);
nand U6712 (N_6712,N_4479,N_3295);
nor U6713 (N_6713,N_5005,N_5684);
or U6714 (N_6714,N_4032,N_3082);
nor U6715 (N_6715,N_4817,N_3007);
xor U6716 (N_6716,N_5960,N_4760);
and U6717 (N_6717,N_3899,N_3016);
and U6718 (N_6718,N_5574,N_4325);
or U6719 (N_6719,N_5894,N_5169);
nand U6720 (N_6720,N_5298,N_5859);
nand U6721 (N_6721,N_4823,N_4560);
nand U6722 (N_6722,N_3953,N_5674);
and U6723 (N_6723,N_5724,N_4278);
or U6724 (N_6724,N_3788,N_5563);
nand U6725 (N_6725,N_3231,N_5374);
nor U6726 (N_6726,N_3328,N_4158);
nor U6727 (N_6727,N_3081,N_4404);
and U6728 (N_6728,N_5791,N_3726);
nor U6729 (N_6729,N_4352,N_3473);
nand U6730 (N_6730,N_4436,N_3046);
nand U6731 (N_6731,N_5321,N_3907);
and U6732 (N_6732,N_3994,N_3351);
nand U6733 (N_6733,N_3305,N_3115);
xor U6734 (N_6734,N_4164,N_4688);
nor U6735 (N_6735,N_3857,N_4872);
and U6736 (N_6736,N_5989,N_3075);
nor U6737 (N_6737,N_4178,N_4365);
xnor U6738 (N_6738,N_3957,N_5406);
nor U6739 (N_6739,N_3807,N_3285);
and U6740 (N_6740,N_3796,N_3488);
nor U6741 (N_6741,N_5246,N_3594);
or U6742 (N_6742,N_4722,N_3017);
nand U6743 (N_6743,N_4916,N_3955);
nand U6744 (N_6744,N_4005,N_5515);
nor U6745 (N_6745,N_5835,N_3040);
xor U6746 (N_6746,N_4076,N_4239);
and U6747 (N_6747,N_3564,N_4255);
nand U6748 (N_6748,N_3692,N_5381);
nand U6749 (N_6749,N_5354,N_4746);
or U6750 (N_6750,N_5112,N_4416);
or U6751 (N_6751,N_3180,N_4620);
nor U6752 (N_6752,N_4007,N_3812);
nor U6753 (N_6753,N_3794,N_4687);
nand U6754 (N_6754,N_5093,N_3599);
and U6755 (N_6755,N_4054,N_5219);
nand U6756 (N_6756,N_3112,N_3181);
and U6757 (N_6757,N_5329,N_4806);
nor U6758 (N_6758,N_3724,N_3842);
and U6759 (N_6759,N_4846,N_5180);
and U6760 (N_6760,N_5798,N_3767);
or U6761 (N_6761,N_4810,N_3707);
nor U6762 (N_6762,N_5125,N_3912);
and U6763 (N_6763,N_4429,N_4700);
or U6764 (N_6764,N_4389,N_3321);
nand U6765 (N_6765,N_3761,N_5150);
and U6766 (N_6766,N_5147,N_4836);
or U6767 (N_6767,N_4452,N_3841);
and U6768 (N_6768,N_5249,N_3756);
and U6769 (N_6769,N_4985,N_3331);
and U6770 (N_6770,N_3247,N_3092);
nand U6771 (N_6771,N_4013,N_3485);
nand U6772 (N_6772,N_5968,N_4813);
nor U6773 (N_6773,N_5145,N_4876);
nand U6774 (N_6774,N_4407,N_5470);
and U6775 (N_6775,N_5108,N_5759);
or U6776 (N_6776,N_5201,N_3124);
or U6777 (N_6777,N_4552,N_3300);
nor U6778 (N_6778,N_4751,N_4403);
nand U6779 (N_6779,N_5738,N_4402);
nand U6780 (N_6780,N_3080,N_3297);
nor U6781 (N_6781,N_4967,N_3755);
or U6782 (N_6782,N_5522,N_3053);
and U6783 (N_6783,N_4245,N_3551);
or U6784 (N_6784,N_3651,N_3719);
nor U6785 (N_6785,N_3596,N_4730);
nand U6786 (N_6786,N_3152,N_4124);
nand U6787 (N_6787,N_5031,N_3459);
or U6788 (N_6788,N_5491,N_4672);
and U6789 (N_6789,N_4240,N_5006);
xor U6790 (N_6790,N_3699,N_5702);
and U6791 (N_6791,N_5646,N_4314);
nor U6792 (N_6792,N_5995,N_3858);
nand U6793 (N_6793,N_4543,N_5618);
nor U6794 (N_6794,N_3783,N_5422);
or U6795 (N_6795,N_4734,N_3954);
nor U6796 (N_6796,N_3973,N_4533);
nor U6797 (N_6797,N_3371,N_3314);
or U6798 (N_6798,N_3072,N_3130);
or U6799 (N_6799,N_3970,N_4401);
and U6800 (N_6800,N_4162,N_3962);
xor U6801 (N_6801,N_5328,N_5000);
nor U6802 (N_6802,N_4174,N_5343);
and U6803 (N_6803,N_5935,N_4603);
or U6804 (N_6804,N_5633,N_5595);
and U6805 (N_6805,N_4058,N_3512);
nor U6806 (N_6806,N_4353,N_5760);
or U6807 (N_6807,N_5308,N_5485);
nor U6808 (N_6808,N_5394,N_3990);
nand U6809 (N_6809,N_3674,N_3636);
or U6810 (N_6810,N_3793,N_5319);
or U6811 (N_6811,N_3420,N_5258);
nor U6812 (N_6812,N_5671,N_3852);
nand U6813 (N_6813,N_5934,N_5611);
or U6814 (N_6814,N_4444,N_5501);
or U6815 (N_6815,N_5821,N_5897);
or U6816 (N_6816,N_4941,N_5530);
nor U6817 (N_6817,N_3917,N_5088);
and U6818 (N_6818,N_3637,N_4833);
nor U6819 (N_6819,N_3639,N_3568);
nand U6820 (N_6820,N_5961,N_3991);
nand U6821 (N_6821,N_4468,N_3509);
xor U6822 (N_6822,N_3341,N_3982);
xnor U6823 (N_6823,N_4855,N_3442);
or U6824 (N_6824,N_3547,N_5708);
or U6825 (N_6825,N_5056,N_3987);
and U6826 (N_6826,N_4130,N_4247);
nor U6827 (N_6827,N_5208,N_4000);
nor U6828 (N_6828,N_5967,N_5162);
nand U6829 (N_6829,N_4237,N_4821);
and U6830 (N_6830,N_4192,N_5158);
nand U6831 (N_6831,N_3810,N_3759);
or U6832 (N_6832,N_4086,N_5170);
and U6833 (N_6833,N_4371,N_4805);
and U6834 (N_6834,N_4309,N_4229);
nor U6835 (N_6835,N_5906,N_3430);
or U6836 (N_6836,N_3252,N_4563);
and U6837 (N_6837,N_5272,N_3603);
xor U6838 (N_6838,N_5311,N_5683);
or U6839 (N_6839,N_3137,N_4129);
xor U6840 (N_6840,N_4864,N_5930);
and U6841 (N_6841,N_5911,N_4647);
nand U6842 (N_6842,N_4579,N_5417);
nand U6843 (N_6843,N_3292,N_5634);
or U6844 (N_6844,N_3554,N_5550);
nand U6845 (N_6845,N_5752,N_4713);
and U6846 (N_6846,N_3627,N_4604);
xor U6847 (N_6847,N_4264,N_3944);
and U6848 (N_6848,N_4021,N_4930);
nor U6849 (N_6849,N_4966,N_5518);
or U6850 (N_6850,N_5662,N_5783);
or U6851 (N_6851,N_5449,N_3464);
nor U6852 (N_6852,N_3066,N_4614);
nand U6853 (N_6853,N_4350,N_5404);
nor U6854 (N_6854,N_4877,N_4607);
xnor U6855 (N_6855,N_5998,N_4196);
and U6856 (N_6856,N_3975,N_4854);
or U6857 (N_6857,N_3621,N_4908);
and U6858 (N_6858,N_5582,N_3319);
nor U6859 (N_6859,N_3189,N_3479);
nor U6860 (N_6860,N_5729,N_3772);
or U6861 (N_6861,N_4661,N_3969);
nor U6862 (N_6862,N_3881,N_4656);
nand U6863 (N_6863,N_5163,N_5965);
nand U6864 (N_6864,N_5669,N_4254);
xnor U6865 (N_6865,N_4968,N_3870);
nand U6866 (N_6866,N_3913,N_4737);
nor U6867 (N_6867,N_3293,N_3746);
nor U6868 (N_6868,N_3657,N_3215);
nor U6869 (N_6869,N_3529,N_5175);
nand U6870 (N_6870,N_4183,N_4510);
and U6871 (N_6871,N_4512,N_3032);
nor U6872 (N_6872,N_4439,N_4443);
and U6873 (N_6873,N_4522,N_4858);
nand U6874 (N_6874,N_5027,N_3105);
nor U6875 (N_6875,N_4098,N_5098);
or U6876 (N_6876,N_4031,N_3148);
nor U6877 (N_6877,N_3736,N_5558);
and U6878 (N_6878,N_4185,N_3199);
and U6879 (N_6879,N_5439,N_3752);
or U6880 (N_6880,N_3921,N_4875);
and U6881 (N_6881,N_3157,N_5545);
xnor U6882 (N_6882,N_3233,N_4802);
and U6883 (N_6883,N_3676,N_3645);
nor U6884 (N_6884,N_3169,N_3377);
and U6885 (N_6885,N_4235,N_4493);
or U6886 (N_6886,N_5833,N_3513);
and U6887 (N_6887,N_5301,N_3686);
nor U6888 (N_6888,N_5861,N_5398);
or U6889 (N_6889,N_4030,N_4260);
and U6890 (N_6890,N_3048,N_5116);
nand U6891 (N_6891,N_4250,N_3790);
nor U6892 (N_6892,N_4521,N_4294);
or U6893 (N_6893,N_4059,N_4758);
and U6894 (N_6894,N_5598,N_5044);
xor U6895 (N_6895,N_5715,N_4194);
xnor U6896 (N_6896,N_3245,N_5171);
or U6897 (N_6897,N_5370,N_5682);
or U6898 (N_6898,N_5838,N_4632);
and U6899 (N_6899,N_4735,N_4375);
or U6900 (N_6900,N_5531,N_3878);
nand U6901 (N_6901,N_3856,N_4709);
or U6902 (N_6902,N_5490,N_4593);
nor U6903 (N_6903,N_5673,N_5221);
or U6904 (N_6904,N_5777,N_5037);
nor U6905 (N_6905,N_3861,N_3867);
nand U6906 (N_6906,N_4393,N_3142);
nand U6907 (N_6907,N_4975,N_4065);
and U6908 (N_6908,N_5519,N_5192);
and U6909 (N_6909,N_5664,N_4480);
and U6910 (N_6910,N_5885,N_4272);
and U6911 (N_6911,N_3535,N_4640);
or U6912 (N_6912,N_4269,N_4343);
nor U6913 (N_6913,N_3620,N_5534);
or U6914 (N_6914,N_3771,N_4663);
or U6915 (N_6915,N_3026,N_3694);
or U6916 (N_6916,N_5976,N_5106);
nor U6917 (N_6917,N_5559,N_5655);
nand U6918 (N_6918,N_4263,N_3873);
and U6919 (N_6919,N_3262,N_4069);
and U6920 (N_6920,N_4033,N_4850);
and U6921 (N_6921,N_5479,N_4949);
nand U6922 (N_6922,N_4974,N_3557);
and U6923 (N_6923,N_4808,N_5389);
or U6924 (N_6924,N_5753,N_5867);
nor U6925 (N_6925,N_4387,N_5969);
and U6926 (N_6926,N_4665,N_5639);
or U6927 (N_6927,N_5181,N_3517);
or U6928 (N_6928,N_4948,N_5218);
nor U6929 (N_6929,N_3219,N_5021);
nor U6930 (N_6930,N_4043,N_5806);
and U6931 (N_6931,N_5344,N_3475);
nand U6932 (N_6932,N_5889,N_3989);
or U6933 (N_6933,N_4520,N_4378);
and U6934 (N_6934,N_3822,N_5377);
nand U6935 (N_6935,N_4026,N_5440);
nand U6936 (N_6936,N_4331,N_4884);
nor U6937 (N_6937,N_5312,N_5933);
or U6938 (N_6938,N_5256,N_4462);
and U6939 (N_6939,N_5090,N_4180);
nor U6940 (N_6940,N_4636,N_5248);
xor U6941 (N_6941,N_3156,N_3624);
or U6942 (N_6942,N_5401,N_4084);
nand U6943 (N_6943,N_3363,N_5385);
nand U6944 (N_6944,N_5356,N_5164);
nor U6945 (N_6945,N_4506,N_3121);
xor U6946 (N_6946,N_5588,N_5438);
nor U6947 (N_6947,N_4621,N_4081);
nor U6948 (N_6948,N_3392,N_5714);
nand U6949 (N_6949,N_5991,N_4224);
or U6950 (N_6950,N_4029,N_3667);
nand U6951 (N_6951,N_4140,N_3763);
xor U6952 (N_6952,N_4570,N_5837);
or U6953 (N_6953,N_4517,N_5275);
nor U6954 (N_6954,N_3228,N_4556);
or U6955 (N_6955,N_4307,N_5946);
nand U6956 (N_6956,N_4983,N_4284);
nor U6957 (N_6957,N_3778,N_3747);
nand U6958 (N_6958,N_3566,N_4146);
or U6959 (N_6959,N_4048,N_5931);
or U6960 (N_6960,N_4348,N_4645);
and U6961 (N_6961,N_3424,N_5874);
nor U6962 (N_6962,N_4210,N_3910);
nand U6963 (N_6963,N_3298,N_3703);
nor U6964 (N_6964,N_5413,N_5399);
and U6965 (N_6965,N_4409,N_5062);
nand U6966 (N_6966,N_4777,N_5909);
or U6967 (N_6967,N_5415,N_3832);
or U6968 (N_6968,N_4052,N_5341);
nor U6969 (N_6969,N_4222,N_5878);
nor U6970 (N_6970,N_5892,N_4848);
nand U6971 (N_6971,N_3284,N_5693);
and U6972 (N_6972,N_4523,N_4580);
and U6973 (N_6973,N_5124,N_3691);
nor U6974 (N_6974,N_5366,N_5030);
and U6975 (N_6975,N_5019,N_3528);
nand U6976 (N_6976,N_4017,N_4101);
nor U6977 (N_6977,N_3089,N_4594);
or U6978 (N_6978,N_5029,N_4464);
nand U6979 (N_6979,N_3416,N_3225);
or U6980 (N_6980,N_4486,N_3570);
nand U6981 (N_6981,N_3592,N_3175);
and U6982 (N_6982,N_4546,N_5535);
and U6983 (N_6983,N_5820,N_3210);
or U6984 (N_6984,N_5250,N_5115);
or U6985 (N_6985,N_4950,N_3821);
nor U6986 (N_6986,N_5433,N_3824);
nor U6987 (N_6987,N_4495,N_3310);
xor U6988 (N_6988,N_3960,N_5273);
and U6989 (N_6989,N_4449,N_3414);
and U6990 (N_6990,N_5376,N_3356);
nor U6991 (N_6991,N_3350,N_5226);
nand U6992 (N_6992,N_4555,N_5293);
nor U6993 (N_6993,N_4163,N_5435);
nand U6994 (N_6994,N_3584,N_4622);
or U6995 (N_6995,N_5049,N_5040);
nand U6996 (N_6996,N_5251,N_5159);
xor U6997 (N_6997,N_5621,N_4651);
nand U6998 (N_6998,N_3678,N_5008);
and U6999 (N_6999,N_4179,N_4973);
nor U7000 (N_7000,N_5097,N_3036);
or U7001 (N_7001,N_4779,N_4338);
nand U7002 (N_7002,N_4766,N_5137);
or U7003 (N_7003,N_5380,N_5764);
nor U7004 (N_7004,N_5978,N_3482);
and U7005 (N_7005,N_3446,N_3934);
and U7006 (N_7006,N_5193,N_5352);
or U7007 (N_7007,N_3179,N_5823);
nor U7008 (N_7008,N_3679,N_3192);
and U7009 (N_7009,N_4166,N_4441);
nor U7010 (N_7010,N_3320,N_3287);
nand U7011 (N_7011,N_5593,N_4678);
or U7012 (N_7012,N_4756,N_4397);
and U7013 (N_7013,N_4554,N_3433);
nand U7014 (N_7014,N_3939,N_4928);
or U7015 (N_7015,N_4217,N_5123);
and U7016 (N_7016,N_3876,N_5525);
and U7017 (N_7017,N_5657,N_3107);
nor U7018 (N_7018,N_5168,N_5279);
nor U7019 (N_7019,N_4472,N_5778);
nor U7020 (N_7020,N_4914,N_4710);
or U7021 (N_7021,N_4177,N_4038);
nand U7022 (N_7022,N_3018,N_5185);
nor U7023 (N_7023,N_3664,N_4792);
nor U7024 (N_7024,N_4502,N_5104);
or U7025 (N_7025,N_4018,N_5409);
xor U7026 (N_7026,N_5938,N_3622);
nor U7027 (N_7027,N_4074,N_3325);
or U7028 (N_7028,N_5710,N_5855);
and U7029 (N_7029,N_5790,N_3360);
nor U7030 (N_7030,N_4828,N_5232);
or U7031 (N_7031,N_5428,N_4440);
nor U7032 (N_7032,N_3558,N_5350);
nor U7033 (N_7033,N_4419,N_4450);
or U7034 (N_7034,N_5079,N_5770);
xor U7035 (N_7035,N_4159,N_4377);
nor U7036 (N_7036,N_5929,N_5338);
nor U7037 (N_7037,N_5034,N_3864);
nand U7038 (N_7038,N_5286,N_5432);
nand U7039 (N_7039,N_3534,N_3968);
nand U7040 (N_7040,N_4686,N_4025);
nand U7041 (N_7041,N_3417,N_3625);
and U7042 (N_7042,N_3600,N_4590);
or U7043 (N_7043,N_5091,N_5448);
or U7044 (N_7044,N_5270,N_5357);
xor U7045 (N_7045,N_4299,N_5828);
and U7046 (N_7046,N_4989,N_5214);
nand U7047 (N_7047,N_3421,N_3220);
or U7048 (N_7048,N_4301,N_5831);
nor U7049 (N_7049,N_4173,N_5648);
and U7050 (N_7050,N_3776,N_3141);
or U7051 (N_7051,N_4189,N_4589);
and U7052 (N_7052,N_4399,N_4220);
nor U7053 (N_7053,N_4936,N_4609);
and U7054 (N_7054,N_4109,N_4616);
nand U7055 (N_7055,N_3504,N_4873);
nand U7056 (N_7056,N_3457,N_3972);
xnor U7057 (N_7057,N_4541,N_5852);
nor U7058 (N_7058,N_5134,N_4080);
nand U7059 (N_7059,N_4592,N_3748);
nor U7060 (N_7060,N_3223,N_5416);
nand U7061 (N_7061,N_3505,N_5540);
xnor U7062 (N_7062,N_4990,N_5472);
and U7063 (N_7063,N_5707,N_3384);
or U7064 (N_7064,N_4913,N_5306);
or U7065 (N_7065,N_4308,N_4537);
xnor U7066 (N_7066,N_3150,N_5197);
xor U7067 (N_7067,N_4447,N_5723);
nand U7068 (N_7068,N_4091,N_3663);
nor U7069 (N_7069,N_4288,N_5688);
and U7070 (N_7070,N_4176,N_3086);
nor U7071 (N_7071,N_4248,N_4612);
nand U7072 (N_7072,N_4747,N_4922);
nor U7073 (N_7073,N_3825,N_4394);
or U7074 (N_7074,N_5762,N_3926);
or U7075 (N_7075,N_5551,N_3754);
nand U7076 (N_7076,N_5880,N_5630);
or U7077 (N_7077,N_4191,N_3277);
nand U7078 (N_7078,N_5694,N_3264);
xnor U7079 (N_7079,N_5444,N_4057);
or U7080 (N_7080,N_4276,N_3606);
and U7081 (N_7081,N_5458,N_3762);
nor U7082 (N_7082,N_3749,N_5948);
and U7083 (N_7083,N_3628,N_5146);
or U7084 (N_7084,N_4606,N_5259);
and U7085 (N_7085,N_4020,N_4501);
nor U7086 (N_7086,N_3607,N_4078);
nor U7087 (N_7087,N_4494,N_4420);
and U7088 (N_7088,N_5353,N_3823);
and U7089 (N_7089,N_3267,N_3143);
nor U7090 (N_7090,N_4388,N_5295);
and U7091 (N_7091,N_3742,N_4769);
nor U7092 (N_7092,N_5018,N_5456);
nor U7093 (N_7093,N_4208,N_4729);
nand U7094 (N_7094,N_5944,N_4892);
xor U7095 (N_7095,N_3751,N_3656);
nor U7096 (N_7096,N_3855,N_4683);
or U7097 (N_7097,N_5054,N_5156);
nor U7098 (N_7098,N_5527,N_5038);
or U7099 (N_7099,N_4273,N_3311);
nor U7100 (N_7100,N_4028,N_3218);
xnor U7101 (N_7101,N_3946,N_3365);
and U7102 (N_7102,N_3638,N_4910);
and U7103 (N_7103,N_5436,N_5302);
and U7104 (N_7104,N_5566,N_4218);
nor U7105 (N_7105,N_5371,N_3318);
or U7106 (N_7106,N_5711,N_3207);
nor U7107 (N_7107,N_3435,N_3974);
xor U7108 (N_7108,N_3715,N_4633);
and U7109 (N_7109,N_3140,N_3096);
and U7110 (N_7110,N_3544,N_3815);
nor U7111 (N_7111,N_5362,N_3238);
xor U7112 (N_7112,N_4428,N_5873);
xnor U7113 (N_7113,N_5896,N_4327);
xor U7114 (N_7114,N_4977,N_4648);
nand U7115 (N_7115,N_3173,N_5484);
or U7116 (N_7116,N_4701,N_5087);
nand U7117 (N_7117,N_3819,N_3519);
nand U7118 (N_7118,N_3869,N_3539);
or U7119 (N_7119,N_3020,N_5419);
xnor U7120 (N_7120,N_3185,N_3492);
nor U7121 (N_7121,N_5756,N_5921);
and U7122 (N_7122,N_5187,N_3542);
nor U7123 (N_7123,N_5940,N_3306);
nor U7124 (N_7124,N_3042,N_3440);
and U7125 (N_7125,N_3024,N_3034);
nand U7126 (N_7126,N_4485,N_3178);
and U7127 (N_7127,N_5668,N_5309);
and U7128 (N_7128,N_5870,N_3395);
nand U7129 (N_7129,N_3372,N_5268);
and U7130 (N_7130,N_3609,N_3981);
nor U7131 (N_7131,N_5576,N_3217);
nor U7132 (N_7132,N_5871,N_3499);
xnor U7133 (N_7133,N_3741,N_4696);
or U7134 (N_7134,N_5536,N_4571);
nand U7135 (N_7135,N_5367,N_4200);
nand U7136 (N_7136,N_4110,N_4108);
and U7137 (N_7137,N_4417,N_4937);
nor U7138 (N_7138,N_3837,N_4642);
nand U7139 (N_7139,N_3087,N_3176);
nand U7140 (N_7140,N_5383,N_4677);
nand U7141 (N_7141,N_3462,N_5157);
nor U7142 (N_7142,N_4134,N_4456);
xor U7143 (N_7143,N_4867,N_5982);
nor U7144 (N_7144,N_4981,N_5466);
nor U7145 (N_7145,N_5012,N_3701);
and U7146 (N_7146,N_3206,N_5941);
or U7147 (N_7147,N_4477,N_3833);
and U7148 (N_7148,N_5532,N_4136);
nor U7149 (N_7149,N_5916,N_5499);
or U7150 (N_7150,N_5092,N_5177);
and U7151 (N_7151,N_5477,N_5066);
xnor U7152 (N_7152,N_3846,N_5468);
xnor U7153 (N_7153,N_3959,N_3498);
nor U7154 (N_7154,N_3491,N_4354);
nor U7155 (N_7155,N_5952,N_3451);
nor U7156 (N_7156,N_4991,N_3658);
and U7157 (N_7157,N_5237,N_3344);
xor U7158 (N_7158,N_5148,N_5421);
nor U7159 (N_7159,N_5825,N_4935);
and U7160 (N_7160,N_4625,N_3737);
nor U7161 (N_7161,N_5544,N_3008);
xnor U7162 (N_7162,N_5910,N_4945);
nor U7163 (N_7163,N_3110,N_4671);
and U7164 (N_7164,N_4881,N_4898);
nor U7165 (N_7165,N_5547,N_4291);
xor U7166 (N_7166,N_3929,N_5478);
and U7167 (N_7167,N_5850,N_4125);
nand U7168 (N_7168,N_3368,N_5866);
and U7169 (N_7169,N_4107,N_3093);
nor U7170 (N_7170,N_4335,N_4801);
nand U7171 (N_7171,N_4454,N_4542);
and U7172 (N_7172,N_4473,N_5473);
and U7173 (N_7173,N_4837,N_4699);
or U7174 (N_7174,N_3728,N_5538);
and U7175 (N_7175,N_5206,N_5149);
nand U7176 (N_7176,N_5314,N_4969);
nor U7177 (N_7177,N_5785,N_4066);
and U7178 (N_7178,N_3988,N_3549);
or U7179 (N_7179,N_3172,N_4530);
nand U7180 (N_7180,N_5533,N_4445);
or U7181 (N_7181,N_3785,N_3820);
nor U7182 (N_7182,N_3071,N_3582);
xnor U7183 (N_7183,N_3545,N_5917);
nand U7184 (N_7184,N_5959,N_5138);
or U7185 (N_7185,N_3308,N_5103);
nand U7186 (N_7186,N_4262,N_4784);
or U7187 (N_7187,N_4811,N_5886);
nand U7188 (N_7188,N_3884,N_3251);
and U7189 (N_7189,N_3301,N_4251);
and U7190 (N_7190,N_5701,N_5358);
or U7191 (N_7191,N_4100,N_4839);
and U7192 (N_7192,N_3227,N_3803);
nor U7193 (N_7193,N_3038,N_5365);
nand U7194 (N_7194,N_3234,N_4418);
and U7195 (N_7195,N_5805,N_3213);
nor U7196 (N_7196,N_4762,N_5200);
nand U7197 (N_7197,N_4705,N_4617);
or U7198 (N_7198,N_5586,N_4759);
nor U7199 (N_7199,N_5676,N_5299);
xnor U7200 (N_7200,N_3074,N_5463);
nor U7201 (N_7201,N_5632,N_5773);
and U7202 (N_7202,N_3393,N_3733);
or U7203 (N_7203,N_3616,N_5609);
nand U7204 (N_7204,N_3782,N_3380);
nor U7205 (N_7205,N_3681,N_4534);
and U7206 (N_7206,N_5165,N_4891);
or U7207 (N_7207,N_4206,N_5679);
xnor U7208 (N_7208,N_5854,N_3265);
xor U7209 (N_7209,N_3452,N_4897);
nand U7210 (N_7210,N_3773,N_3155);
or U7211 (N_7211,N_3004,N_5359);
nor U7212 (N_7212,N_3465,N_3214);
or U7213 (N_7213,N_3035,N_3541);
or U7214 (N_7214,N_3650,N_5015);
or U7215 (N_7215,N_4944,N_4396);
nor U7216 (N_7216,N_3872,N_3851);
xor U7217 (N_7217,N_5716,N_3083);
nand U7218 (N_7218,N_3111,N_5195);
and U7219 (N_7219,N_3438,N_3084);
and U7220 (N_7220,N_5858,N_3672);
and U7221 (N_7221,N_5692,N_3448);
and U7222 (N_7222,N_3874,N_5403);
and U7223 (N_7223,N_5726,N_5202);
nor U7224 (N_7224,N_4227,N_4457);
nor U7225 (N_7225,N_3520,N_5659);
or U7226 (N_7226,N_3590,N_4979);
xnor U7227 (N_7227,N_3289,N_4790);
nor U7228 (N_7228,N_3980,N_5973);
or U7229 (N_7229,N_4225,N_3661);
or U7230 (N_7230,N_5217,N_3138);
or U7231 (N_7231,N_4557,N_4302);
nand U7232 (N_7232,N_5776,N_5624);
nand U7233 (N_7233,N_3897,N_4169);
and U7234 (N_7234,N_5475,N_3257);
nor U7235 (N_7235,N_3357,N_4096);
xnor U7236 (N_7236,N_4738,N_3996);
nand U7237 (N_7237,N_4655,N_4646);
and U7238 (N_7238,N_3246,N_5014);
nand U7239 (N_7239,N_5050,N_3887);
nand U7240 (N_7240,N_3687,N_3394);
and U7241 (N_7241,N_5136,N_4432);
and U7242 (N_7242,N_4011,N_3816);
or U7243 (N_7243,N_4807,N_3576);
nor U7244 (N_7244,N_5809,N_4690);
and U7245 (N_7245,N_5429,N_4001);
or U7246 (N_7246,N_5242,N_3113);
and U7247 (N_7247,N_4666,N_3168);
nand U7248 (N_7248,N_3581,N_5784);
and U7249 (N_7249,N_3593,N_5956);
nand U7250 (N_7250,N_4467,N_3589);
xor U7251 (N_7251,N_3798,N_3943);
and U7252 (N_7252,N_5172,N_4992);
or U7253 (N_7253,N_4885,N_5228);
nand U7254 (N_7254,N_3167,N_3064);
nor U7255 (N_7255,N_3854,N_4410);
or U7256 (N_7256,N_3000,N_4168);
nand U7257 (N_7257,N_3077,N_4847);
and U7258 (N_7258,N_5288,N_3398);
xor U7259 (N_7259,N_3373,N_5055);
nand U7260 (N_7260,N_3531,N_5154);
nor U7261 (N_7261,N_3239,N_4265);
and U7262 (N_7262,N_4258,N_4077);
and U7263 (N_7263,N_5945,N_3456);
nand U7264 (N_7264,N_5489,N_5213);
or U7265 (N_7265,N_3805,N_3523);
nor U7266 (N_7266,N_3768,N_4160);
or U7267 (N_7267,N_4719,N_3260);
xnor U7268 (N_7268,N_3506,N_5457);
or U7269 (N_7269,N_4776,N_4887);
and U7270 (N_7270,N_5819,N_3986);
or U7271 (N_7271,N_4281,N_5542);
and U7272 (N_7272,N_5926,N_3088);
and U7273 (N_7273,N_4923,N_4036);
and U7274 (N_7274,N_5769,N_3256);
nor U7275 (N_7275,N_3146,N_3704);
nand U7276 (N_7276,N_5883,N_3732);
and U7277 (N_7277,N_5388,N_5390);
nand U7278 (N_7278,N_4740,N_3800);
or U7279 (N_7279,N_5269,N_5514);
and U7280 (N_7280,N_4886,N_3033);
nor U7281 (N_7281,N_3697,N_5990);
nand U7282 (N_7282,N_5083,N_4256);
nor U7283 (N_7283,N_4681,N_5085);
nand U7284 (N_7284,N_3546,N_3428);
xnor U7285 (N_7285,N_3952,N_5807);
nor U7286 (N_7286,N_3458,N_5800);
and U7287 (N_7287,N_3400,N_3840);
or U7288 (N_7288,N_5229,N_4015);
or U7289 (N_7289,N_5672,N_3553);
or U7290 (N_7290,N_5529,N_5324);
and U7291 (N_7291,N_5254,N_4039);
nand U7292 (N_7292,N_5261,N_4962);
or U7293 (N_7293,N_4774,N_5918);
nor U7294 (N_7294,N_5615,N_4105);
nand U7295 (N_7295,N_5461,N_4193);
nand U7296 (N_7296,N_3337,N_5111);
or U7297 (N_7297,N_3745,N_4692);
xnor U7298 (N_7298,N_4650,N_3961);
or U7299 (N_7299,N_4398,N_4804);
or U7300 (N_7300,N_5840,N_5927);
nor U7301 (N_7301,N_3685,N_5751);
and U7302 (N_7302,N_5857,N_5733);
nand U7303 (N_7303,N_3765,N_4087);
nor U7304 (N_7304,N_5902,N_3784);
nor U7305 (N_7305,N_5139,N_4550);
nor U7306 (N_7306,N_5119,N_4430);
and U7307 (N_7307,N_3817,N_5556);
or U7308 (N_7308,N_5264,N_4818);
nor U7309 (N_7309,N_3764,N_3683);
or U7310 (N_7310,N_4319,N_3580);
nand U7311 (N_7311,N_5985,N_3044);
or U7312 (N_7312,N_4932,N_4917);
and U7313 (N_7313,N_3258,N_3006);
and U7314 (N_7314,N_4957,N_4322);
and U7315 (N_7315,N_3971,N_4953);
nand U7316 (N_7316,N_5516,N_4578);
or U7317 (N_7317,N_5644,N_5986);
nor U7318 (N_7318,N_4507,N_5364);
and U7319 (N_7319,N_5144,N_4954);
nor U7320 (N_7320,N_5471,N_4771);
nor U7321 (N_7321,N_3666,N_4978);
or U7322 (N_7322,N_3010,N_3750);
nand U7323 (N_7323,N_5122,N_3920);
or U7324 (N_7324,N_4874,N_3847);
nand U7325 (N_7325,N_4252,N_5327);
nand U7326 (N_7326,N_3198,N_3315);
and U7327 (N_7327,N_3153,N_3791);
nand U7328 (N_7328,N_4188,N_5721);
or U7329 (N_7329,N_3326,N_3423);
and U7330 (N_7330,N_4286,N_3411);
nand U7331 (N_7331,N_5361,N_5731);
or U7332 (N_7332,N_5280,N_4761);
or U7333 (N_7333,N_5351,N_3789);
and U7334 (N_7334,N_3177,N_3422);
and U7335 (N_7335,N_3012,N_3652);
nand U7336 (N_7336,N_4027,N_3127);
xor U7337 (N_7337,N_3103,N_4618);
or U7338 (N_7338,N_3835,N_3379);
and U7339 (N_7339,N_3455,N_5626);
xor U7340 (N_7340,N_5570,N_4489);
nand U7341 (N_7341,N_4742,N_4598);
and U7342 (N_7342,N_4861,N_5629);
nand U7343 (N_7343,N_3052,N_4434);
and U7344 (N_7344,N_4147,N_3195);
or U7345 (N_7345,N_5459,N_4965);
xnor U7346 (N_7346,N_5240,N_3677);
or U7347 (N_7347,N_3106,N_4355);
and U7348 (N_7348,N_4532,N_3604);
or U7349 (N_7349,N_5511,N_4652);
and U7350 (N_7350,N_4453,N_3905);
nor U7351 (N_7351,N_5818,N_5446);
and U7352 (N_7352,N_3949,N_3525);
nor U7353 (N_7353,N_4499,N_3702);
xnor U7354 (N_7354,N_5920,N_3530);
nand U7355 (N_7355,N_3826,N_4588);
nand U7356 (N_7356,N_3288,N_5649);
nand U7357 (N_7357,N_4515,N_4518);
nor U7358 (N_7358,N_4383,N_4994);
and U7359 (N_7359,N_5680,N_5656);
or U7360 (N_7360,N_4143,N_3323);
nand U7361 (N_7361,N_5832,N_3340);
and U7362 (N_7362,N_5763,N_3471);
nor U7363 (N_7363,N_3770,N_4205);
nor U7364 (N_7364,N_5290,N_3659);
nand U7365 (N_7365,N_5853,N_4504);
nand U7366 (N_7366,N_3294,N_5057);
xnor U7367 (N_7367,N_4868,N_3461);
nor U7368 (N_7368,N_3605,N_4786);
nand U7369 (N_7369,N_5326,N_5178);
or U7370 (N_7370,N_5660,N_5211);
xnor U7371 (N_7371,N_5977,N_5690);
nand U7372 (N_7372,N_5845,N_5829);
and U7373 (N_7373,N_4840,N_3831);
and U7374 (N_7374,N_5017,N_3278);
and U7375 (N_7375,N_4752,N_3668);
or U7376 (N_7376,N_3516,N_5573);
and U7377 (N_7377,N_4657,N_3165);
or U7378 (N_7378,N_4006,N_5827);
and U7379 (N_7379,N_4575,N_3271);
or U7380 (N_7380,N_4727,N_5060);
nand U7381 (N_7381,N_3282,N_3931);
nand U7382 (N_7382,N_5970,N_3235);
nor U7383 (N_7383,N_4835,N_4768);
and U7384 (N_7384,N_5198,N_4190);
or U7385 (N_7385,N_3885,N_5766);
nor U7386 (N_7386,N_5414,N_5176);
or U7387 (N_7387,N_4121,N_4545);
xnor U7388 (N_7388,N_3369,N_4326);
nor U7389 (N_7389,N_5765,N_3712);
or U7390 (N_7390,N_4182,N_5010);
nor U7391 (N_7391,N_3070,N_3578);
or U7392 (N_7392,N_3795,N_3109);
or U7393 (N_7393,N_3830,N_3514);
or U7394 (N_7394,N_3003,N_4412);
and U7395 (N_7395,N_3979,N_4361);
nor U7396 (N_7396,N_3338,N_4597);
and U7397 (N_7397,N_3191,N_4654);
xnor U7398 (N_7398,N_4581,N_3508);
or U7399 (N_7399,N_4574,N_4061);
xnor U7400 (N_7400,N_3706,N_5627);
or U7401 (N_7401,N_5699,N_5923);
or U7402 (N_7402,N_5788,N_4951);
nor U7403 (N_7403,N_4382,N_5071);
xnor U7404 (N_7404,N_4596,N_5808);
xor U7405 (N_7405,N_5628,N_3418);
xor U7406 (N_7406,N_5592,N_3586);
and U7407 (N_7407,N_5709,N_4870);
nand U7408 (N_7408,N_3948,N_5487);
nand U7409 (N_7409,N_3591,N_3183);
nor U7410 (N_7410,N_5041,N_5584);
or U7411 (N_7411,N_5284,N_5507);
xnor U7412 (N_7412,N_3154,N_4016);
and U7413 (N_7413,N_3280,N_4536);
and U7414 (N_7414,N_3919,N_4300);
or U7415 (N_7415,N_3839,N_3401);
nand U7416 (N_7416,N_4062,N_5571);
or U7417 (N_7417,N_5402,N_5849);
nor U7418 (N_7418,N_5600,N_4921);
nor U7419 (N_7419,N_4304,N_3317);
or U7420 (N_7420,N_3483,N_3263);
nor U7421 (N_7421,N_5016,N_4073);
and U7422 (N_7422,N_4460,N_4653);
or U7423 (N_7423,N_3149,N_5483);
nor U7424 (N_7424,N_3758,N_5795);
nor U7425 (N_7425,N_3375,N_5497);
and U7426 (N_7426,N_4275,N_3104);
and U7427 (N_7427,N_5771,N_5160);
xnor U7428 (N_7428,N_5486,N_5257);
or U7429 (N_7429,N_3779,N_3230);
nor U7430 (N_7430,N_5815,N_5239);
and U7431 (N_7431,N_4085,N_5474);
nor U7432 (N_7432,N_3998,N_5418);
or U7433 (N_7433,N_5811,N_5904);
and U7434 (N_7434,N_3013,N_3556);
nand U7435 (N_7435,N_3781,N_3693);
nand U7436 (N_7436,N_5274,N_5954);
nor U7437 (N_7437,N_3222,N_3274);
and U7438 (N_7438,N_4635,N_5082);
xnor U7439 (N_7439,N_3286,N_3501);
nor U7440 (N_7440,N_4698,N_5565);
nor U7441 (N_7441,N_3860,N_3355);
xor U7442 (N_7442,N_4334,N_5339);
nand U7443 (N_7443,N_5001,N_5013);
and U7444 (N_7444,N_4551,N_4595);
or U7445 (N_7445,N_3489,N_5215);
nand U7446 (N_7446,N_3518,N_4112);
nand U7447 (N_7447,N_4024,N_5188);
nor U7448 (N_7448,N_4320,N_5373);
xnor U7449 (N_7449,N_5305,N_5052);
nand U7450 (N_7450,N_4775,N_4613);
nand U7451 (N_7451,N_4569,N_3792);
nor U7452 (N_7452,N_3335,N_5325);
nor U7453 (N_7453,N_4955,N_5183);
and U7454 (N_7454,N_5452,N_5706);
or U7455 (N_7455,N_4918,N_3468);
nor U7456 (N_7456,N_3334,N_5304);
or U7457 (N_7457,N_3307,N_5523);
xnor U7458 (N_7458,N_5932,N_4316);
nor U7459 (N_7459,N_3879,N_5606);
nand U7460 (N_7460,N_5775,N_5323);
nor U7461 (N_7461,N_4572,N_4023);
or U7462 (N_7462,N_4431,N_4466);
nand U7463 (N_7463,N_4852,N_4995);
xnor U7464 (N_7464,N_3160,N_3900);
or U7465 (N_7465,N_4753,N_3359);
nor U7466 (N_7466,N_3494,N_3226);
or U7467 (N_7467,N_3904,N_5981);
nand U7468 (N_7468,N_4703,N_4186);
and U7469 (N_7469,N_4796,N_4845);
nand U7470 (N_7470,N_3041,N_4415);
nand U7471 (N_7471,N_3848,N_4585);
and U7472 (N_7472,N_3992,N_4279);
xor U7473 (N_7473,N_5205,N_3730);
or U7474 (N_7474,N_5939,N_3655);
or U7475 (N_7475,N_4012,N_4336);
or U7476 (N_7476,N_5803,N_3129);
or U7477 (N_7477,N_3051,N_5512);
or U7478 (N_7478,N_4915,N_5749);
or U7479 (N_7479,N_5743,N_5779);
or U7480 (N_7480,N_3405,N_5577);
xor U7481 (N_7481,N_5919,N_5076);
nand U7482 (N_7482,N_4270,N_3891);
or U7483 (N_7483,N_3644,N_5975);
nor U7484 (N_7484,N_4841,N_5387);
nor U7485 (N_7485,N_5893,N_4513);
or U7486 (N_7486,N_5912,N_5320);
and U7487 (N_7487,N_5865,N_4152);
and U7488 (N_7488,N_4455,N_3209);
xor U7489 (N_7489,N_4305,N_4209);
nor U7490 (N_7490,N_4230,N_4757);
xnor U7491 (N_7491,N_4097,N_5740);
and U7492 (N_7492,N_4373,N_3575);
xnor U7493 (N_7493,N_4184,N_4274);
nand U7494 (N_7494,N_4347,N_4660);
or U7495 (N_7495,N_5844,N_3378);
nor U7496 (N_7496,N_4879,N_5120);
or U7497 (N_7497,N_5317,N_5737);
or U7498 (N_7498,N_4370,N_4442);
and U7499 (N_7499,N_5003,N_4803);
and U7500 (N_7500,N_5232,N_5030);
nor U7501 (N_7501,N_3394,N_4715);
xnor U7502 (N_7502,N_5074,N_4217);
and U7503 (N_7503,N_4921,N_5842);
and U7504 (N_7504,N_3631,N_4310);
and U7505 (N_7505,N_3948,N_3782);
nor U7506 (N_7506,N_5645,N_4358);
nand U7507 (N_7507,N_3406,N_5435);
and U7508 (N_7508,N_5301,N_3785);
nand U7509 (N_7509,N_3615,N_3741);
nand U7510 (N_7510,N_3421,N_4541);
nor U7511 (N_7511,N_4760,N_3117);
or U7512 (N_7512,N_5319,N_4215);
and U7513 (N_7513,N_4732,N_5900);
nor U7514 (N_7514,N_5015,N_4056);
nand U7515 (N_7515,N_3693,N_4864);
or U7516 (N_7516,N_5802,N_5058);
nand U7517 (N_7517,N_3867,N_3951);
or U7518 (N_7518,N_3228,N_4908);
nand U7519 (N_7519,N_5497,N_4936);
and U7520 (N_7520,N_5763,N_5693);
nor U7521 (N_7521,N_4544,N_3397);
nand U7522 (N_7522,N_4358,N_4080);
nand U7523 (N_7523,N_3911,N_4002);
or U7524 (N_7524,N_5229,N_4927);
nor U7525 (N_7525,N_4471,N_5211);
nor U7526 (N_7526,N_5661,N_5026);
and U7527 (N_7527,N_5415,N_3295);
nor U7528 (N_7528,N_4267,N_5320);
nor U7529 (N_7529,N_4967,N_5513);
nand U7530 (N_7530,N_3297,N_4615);
and U7531 (N_7531,N_3269,N_3728);
nand U7532 (N_7532,N_4495,N_4925);
nor U7533 (N_7533,N_4064,N_3959);
nor U7534 (N_7534,N_3354,N_4727);
nor U7535 (N_7535,N_5187,N_4697);
and U7536 (N_7536,N_3284,N_5290);
and U7537 (N_7537,N_5700,N_5514);
nand U7538 (N_7538,N_5251,N_5833);
nor U7539 (N_7539,N_3409,N_4490);
nand U7540 (N_7540,N_4594,N_3053);
and U7541 (N_7541,N_3378,N_5741);
nand U7542 (N_7542,N_3759,N_3634);
nor U7543 (N_7543,N_3750,N_5350);
and U7544 (N_7544,N_4427,N_3105);
and U7545 (N_7545,N_5545,N_5127);
nand U7546 (N_7546,N_3585,N_4887);
and U7547 (N_7547,N_3131,N_3987);
nand U7548 (N_7548,N_5812,N_3365);
nor U7549 (N_7549,N_4776,N_5861);
nor U7550 (N_7550,N_4674,N_3677);
and U7551 (N_7551,N_4116,N_5166);
or U7552 (N_7552,N_5072,N_4264);
nand U7553 (N_7553,N_3777,N_3418);
nand U7554 (N_7554,N_3279,N_3974);
xor U7555 (N_7555,N_5621,N_4255);
nor U7556 (N_7556,N_4339,N_3388);
xnor U7557 (N_7557,N_4834,N_4502);
or U7558 (N_7558,N_4709,N_5889);
and U7559 (N_7559,N_5267,N_4844);
xnor U7560 (N_7560,N_4172,N_5743);
nor U7561 (N_7561,N_4540,N_4636);
nor U7562 (N_7562,N_4079,N_5913);
nand U7563 (N_7563,N_5304,N_4081);
or U7564 (N_7564,N_3876,N_4562);
nor U7565 (N_7565,N_4206,N_3077);
or U7566 (N_7566,N_3948,N_3310);
xor U7567 (N_7567,N_4863,N_3979);
or U7568 (N_7568,N_5916,N_3453);
nand U7569 (N_7569,N_4182,N_5021);
xnor U7570 (N_7570,N_4967,N_3442);
nor U7571 (N_7571,N_4444,N_5945);
nor U7572 (N_7572,N_4121,N_5838);
nand U7573 (N_7573,N_4960,N_3938);
or U7574 (N_7574,N_4431,N_3065);
or U7575 (N_7575,N_3351,N_5951);
and U7576 (N_7576,N_3252,N_5495);
and U7577 (N_7577,N_5441,N_4620);
and U7578 (N_7578,N_4095,N_5033);
xnor U7579 (N_7579,N_3112,N_3042);
and U7580 (N_7580,N_3151,N_5441);
nor U7581 (N_7581,N_5461,N_4665);
nor U7582 (N_7582,N_3672,N_3644);
or U7583 (N_7583,N_4489,N_4229);
or U7584 (N_7584,N_5647,N_4902);
and U7585 (N_7585,N_3716,N_3929);
nor U7586 (N_7586,N_5167,N_3220);
nor U7587 (N_7587,N_3402,N_5840);
and U7588 (N_7588,N_3272,N_4935);
nand U7589 (N_7589,N_3068,N_3225);
and U7590 (N_7590,N_5752,N_5573);
nor U7591 (N_7591,N_5640,N_3668);
or U7592 (N_7592,N_3757,N_4514);
nand U7593 (N_7593,N_5681,N_3976);
xnor U7594 (N_7594,N_3059,N_4472);
or U7595 (N_7595,N_3672,N_5459);
and U7596 (N_7596,N_4471,N_5441);
and U7597 (N_7597,N_4532,N_5257);
and U7598 (N_7598,N_4884,N_4797);
or U7599 (N_7599,N_4992,N_3287);
or U7600 (N_7600,N_3820,N_3121);
and U7601 (N_7601,N_5930,N_4408);
nand U7602 (N_7602,N_4122,N_5391);
and U7603 (N_7603,N_3555,N_5618);
nand U7604 (N_7604,N_3290,N_3681);
or U7605 (N_7605,N_5429,N_4382);
nand U7606 (N_7606,N_5106,N_4321);
or U7607 (N_7607,N_4815,N_5507);
and U7608 (N_7608,N_3837,N_4768);
or U7609 (N_7609,N_3522,N_5215);
nand U7610 (N_7610,N_4071,N_5694);
nor U7611 (N_7611,N_4920,N_3855);
or U7612 (N_7612,N_3343,N_5448);
or U7613 (N_7613,N_4446,N_3855);
and U7614 (N_7614,N_5886,N_4454);
nand U7615 (N_7615,N_3164,N_4207);
or U7616 (N_7616,N_4573,N_4713);
xor U7617 (N_7617,N_5976,N_5238);
nor U7618 (N_7618,N_4893,N_5477);
nand U7619 (N_7619,N_5818,N_5559);
and U7620 (N_7620,N_4301,N_4724);
and U7621 (N_7621,N_5071,N_3115);
nand U7622 (N_7622,N_5374,N_4829);
nor U7623 (N_7623,N_4318,N_4742);
nand U7624 (N_7624,N_3205,N_4047);
nor U7625 (N_7625,N_5166,N_3929);
and U7626 (N_7626,N_3088,N_5177);
xnor U7627 (N_7627,N_4603,N_3933);
or U7628 (N_7628,N_4889,N_4777);
or U7629 (N_7629,N_5783,N_4898);
nand U7630 (N_7630,N_5900,N_4193);
and U7631 (N_7631,N_5460,N_3294);
nand U7632 (N_7632,N_4976,N_3350);
and U7633 (N_7633,N_3369,N_3628);
or U7634 (N_7634,N_5143,N_4025);
and U7635 (N_7635,N_4048,N_4801);
xnor U7636 (N_7636,N_4377,N_3709);
or U7637 (N_7637,N_4474,N_4135);
nor U7638 (N_7638,N_5358,N_4933);
and U7639 (N_7639,N_5491,N_4515);
xor U7640 (N_7640,N_3813,N_5792);
and U7641 (N_7641,N_4395,N_4496);
nand U7642 (N_7642,N_5992,N_4445);
nor U7643 (N_7643,N_5139,N_4483);
xor U7644 (N_7644,N_5790,N_5077);
nand U7645 (N_7645,N_4119,N_5256);
nand U7646 (N_7646,N_3925,N_5239);
nor U7647 (N_7647,N_4454,N_4129);
nor U7648 (N_7648,N_3725,N_3281);
or U7649 (N_7649,N_3877,N_3979);
or U7650 (N_7650,N_5364,N_3323);
nor U7651 (N_7651,N_5728,N_3938);
nand U7652 (N_7652,N_3863,N_3205);
and U7653 (N_7653,N_5865,N_4862);
or U7654 (N_7654,N_4894,N_5161);
nand U7655 (N_7655,N_4951,N_3456);
nor U7656 (N_7656,N_4169,N_4902);
xor U7657 (N_7657,N_3397,N_3197);
and U7658 (N_7658,N_3809,N_5294);
nand U7659 (N_7659,N_3537,N_5096);
nor U7660 (N_7660,N_3083,N_3147);
nor U7661 (N_7661,N_4212,N_4706);
xor U7662 (N_7662,N_5298,N_3644);
and U7663 (N_7663,N_5444,N_5670);
or U7664 (N_7664,N_4412,N_5765);
xor U7665 (N_7665,N_5426,N_3014);
xnor U7666 (N_7666,N_3733,N_3090);
and U7667 (N_7667,N_4066,N_4595);
nor U7668 (N_7668,N_3676,N_5025);
and U7669 (N_7669,N_4823,N_4845);
or U7670 (N_7670,N_5380,N_4118);
nor U7671 (N_7671,N_3480,N_5962);
or U7672 (N_7672,N_3083,N_5372);
or U7673 (N_7673,N_4541,N_4706);
xnor U7674 (N_7674,N_4579,N_3054);
and U7675 (N_7675,N_5147,N_5010);
and U7676 (N_7676,N_3874,N_5503);
or U7677 (N_7677,N_5868,N_5183);
nor U7678 (N_7678,N_5529,N_3581);
nor U7679 (N_7679,N_3831,N_4565);
nor U7680 (N_7680,N_5029,N_4668);
xor U7681 (N_7681,N_3918,N_5865);
and U7682 (N_7682,N_4222,N_5315);
and U7683 (N_7683,N_5992,N_4076);
or U7684 (N_7684,N_4269,N_5857);
nand U7685 (N_7685,N_5075,N_3560);
or U7686 (N_7686,N_3554,N_5700);
nand U7687 (N_7687,N_3110,N_3266);
nand U7688 (N_7688,N_5069,N_4736);
or U7689 (N_7689,N_3380,N_4749);
nor U7690 (N_7690,N_5165,N_5130);
and U7691 (N_7691,N_5570,N_5681);
nor U7692 (N_7692,N_3910,N_5914);
and U7693 (N_7693,N_3225,N_5404);
or U7694 (N_7694,N_4414,N_4544);
nor U7695 (N_7695,N_3122,N_4173);
and U7696 (N_7696,N_4603,N_4099);
and U7697 (N_7697,N_4564,N_5663);
or U7698 (N_7698,N_3556,N_5089);
xnor U7699 (N_7699,N_5381,N_3962);
nand U7700 (N_7700,N_5624,N_3189);
nor U7701 (N_7701,N_5585,N_3851);
or U7702 (N_7702,N_5476,N_4062);
nand U7703 (N_7703,N_5128,N_4040);
nor U7704 (N_7704,N_3313,N_4144);
nor U7705 (N_7705,N_5283,N_3398);
nand U7706 (N_7706,N_3800,N_3754);
nand U7707 (N_7707,N_5542,N_3926);
nand U7708 (N_7708,N_4534,N_4444);
or U7709 (N_7709,N_3310,N_5047);
and U7710 (N_7710,N_3547,N_3536);
and U7711 (N_7711,N_3493,N_4838);
nor U7712 (N_7712,N_3332,N_5071);
xnor U7713 (N_7713,N_5148,N_3285);
nor U7714 (N_7714,N_5863,N_4744);
nor U7715 (N_7715,N_4100,N_5853);
and U7716 (N_7716,N_3773,N_5591);
xnor U7717 (N_7717,N_4995,N_4694);
and U7718 (N_7718,N_5910,N_5649);
and U7719 (N_7719,N_5410,N_4689);
or U7720 (N_7720,N_4742,N_5227);
nor U7721 (N_7721,N_3893,N_4444);
xor U7722 (N_7722,N_3747,N_5928);
or U7723 (N_7723,N_5005,N_3697);
nand U7724 (N_7724,N_4706,N_4254);
and U7725 (N_7725,N_5595,N_3784);
nand U7726 (N_7726,N_5497,N_3259);
nor U7727 (N_7727,N_3356,N_4160);
nand U7728 (N_7728,N_5341,N_5468);
nor U7729 (N_7729,N_5476,N_3722);
or U7730 (N_7730,N_5702,N_4527);
nor U7731 (N_7731,N_4544,N_5974);
nor U7732 (N_7732,N_4472,N_5653);
or U7733 (N_7733,N_4316,N_5526);
nand U7734 (N_7734,N_3867,N_3276);
or U7735 (N_7735,N_5064,N_3185);
nand U7736 (N_7736,N_5425,N_5313);
or U7737 (N_7737,N_4963,N_5072);
nor U7738 (N_7738,N_5568,N_3211);
xor U7739 (N_7739,N_4873,N_4205);
nor U7740 (N_7740,N_4644,N_3633);
and U7741 (N_7741,N_5663,N_3875);
nor U7742 (N_7742,N_4982,N_3585);
nor U7743 (N_7743,N_4506,N_5444);
nor U7744 (N_7744,N_4130,N_5903);
nor U7745 (N_7745,N_3460,N_5678);
nor U7746 (N_7746,N_4682,N_3166);
and U7747 (N_7747,N_5015,N_3001);
and U7748 (N_7748,N_4572,N_5719);
or U7749 (N_7749,N_5529,N_3186);
nor U7750 (N_7750,N_4302,N_4239);
and U7751 (N_7751,N_3885,N_4112);
or U7752 (N_7752,N_5580,N_3777);
nand U7753 (N_7753,N_4150,N_4091);
and U7754 (N_7754,N_5152,N_3520);
xor U7755 (N_7755,N_4231,N_5151);
nor U7756 (N_7756,N_4733,N_5224);
nand U7757 (N_7757,N_3419,N_5347);
or U7758 (N_7758,N_4649,N_3952);
and U7759 (N_7759,N_4925,N_4437);
or U7760 (N_7760,N_3509,N_4422);
nor U7761 (N_7761,N_3656,N_5643);
and U7762 (N_7762,N_4475,N_5389);
xnor U7763 (N_7763,N_3953,N_4343);
xnor U7764 (N_7764,N_5560,N_4203);
xor U7765 (N_7765,N_4258,N_3662);
and U7766 (N_7766,N_4527,N_4011);
nand U7767 (N_7767,N_4126,N_4293);
or U7768 (N_7768,N_3719,N_3794);
or U7769 (N_7769,N_4086,N_4332);
or U7770 (N_7770,N_5846,N_4963);
xor U7771 (N_7771,N_5976,N_3271);
and U7772 (N_7772,N_4500,N_3795);
nand U7773 (N_7773,N_3026,N_3474);
nor U7774 (N_7774,N_5755,N_5389);
and U7775 (N_7775,N_5248,N_4654);
or U7776 (N_7776,N_4041,N_4902);
xor U7777 (N_7777,N_4534,N_5603);
nor U7778 (N_7778,N_3756,N_4638);
or U7779 (N_7779,N_3211,N_3719);
and U7780 (N_7780,N_3386,N_4694);
nand U7781 (N_7781,N_3079,N_4949);
or U7782 (N_7782,N_4427,N_4684);
and U7783 (N_7783,N_4892,N_4633);
nand U7784 (N_7784,N_3478,N_3111);
or U7785 (N_7785,N_5717,N_3839);
nor U7786 (N_7786,N_3265,N_5200);
nor U7787 (N_7787,N_3288,N_4931);
or U7788 (N_7788,N_5698,N_5525);
nor U7789 (N_7789,N_5028,N_3575);
nand U7790 (N_7790,N_4776,N_3364);
or U7791 (N_7791,N_5840,N_3849);
or U7792 (N_7792,N_5043,N_3956);
xnor U7793 (N_7793,N_4654,N_3397);
or U7794 (N_7794,N_3966,N_3661);
or U7795 (N_7795,N_3228,N_4440);
nor U7796 (N_7796,N_4909,N_4882);
nand U7797 (N_7797,N_3671,N_4639);
or U7798 (N_7798,N_3818,N_4034);
or U7799 (N_7799,N_5705,N_5357);
or U7800 (N_7800,N_4267,N_4984);
nor U7801 (N_7801,N_3420,N_3724);
and U7802 (N_7802,N_5775,N_4933);
or U7803 (N_7803,N_3941,N_4123);
nand U7804 (N_7804,N_5792,N_5496);
nor U7805 (N_7805,N_5696,N_4293);
and U7806 (N_7806,N_4068,N_3670);
and U7807 (N_7807,N_5476,N_5065);
and U7808 (N_7808,N_4990,N_4504);
nor U7809 (N_7809,N_5755,N_5970);
and U7810 (N_7810,N_4264,N_3805);
xor U7811 (N_7811,N_5586,N_5042);
xnor U7812 (N_7812,N_5573,N_4784);
and U7813 (N_7813,N_5732,N_3282);
nor U7814 (N_7814,N_5778,N_4646);
nand U7815 (N_7815,N_4585,N_4858);
nand U7816 (N_7816,N_3334,N_4705);
nor U7817 (N_7817,N_5831,N_5795);
or U7818 (N_7818,N_3031,N_5529);
nor U7819 (N_7819,N_3733,N_3710);
or U7820 (N_7820,N_3868,N_4899);
or U7821 (N_7821,N_3503,N_4644);
nor U7822 (N_7822,N_4042,N_4191);
nor U7823 (N_7823,N_3955,N_5993);
and U7824 (N_7824,N_5084,N_4134);
and U7825 (N_7825,N_4857,N_5117);
nand U7826 (N_7826,N_4206,N_4534);
nor U7827 (N_7827,N_4608,N_3436);
and U7828 (N_7828,N_5470,N_5552);
or U7829 (N_7829,N_3650,N_4965);
or U7830 (N_7830,N_3549,N_5655);
nor U7831 (N_7831,N_4769,N_3572);
xnor U7832 (N_7832,N_5860,N_5816);
or U7833 (N_7833,N_5726,N_4209);
nor U7834 (N_7834,N_5842,N_5917);
and U7835 (N_7835,N_5416,N_3077);
and U7836 (N_7836,N_3593,N_4407);
and U7837 (N_7837,N_4770,N_4386);
xor U7838 (N_7838,N_4873,N_3192);
and U7839 (N_7839,N_3620,N_4448);
or U7840 (N_7840,N_5606,N_5445);
nand U7841 (N_7841,N_4323,N_3296);
nor U7842 (N_7842,N_3981,N_3789);
or U7843 (N_7843,N_4678,N_3715);
and U7844 (N_7844,N_3516,N_5404);
or U7845 (N_7845,N_5417,N_4450);
and U7846 (N_7846,N_3269,N_3130);
nor U7847 (N_7847,N_3993,N_5050);
nand U7848 (N_7848,N_3777,N_5142);
nor U7849 (N_7849,N_4102,N_3102);
or U7850 (N_7850,N_3363,N_3883);
xor U7851 (N_7851,N_5149,N_5401);
or U7852 (N_7852,N_5022,N_4193);
and U7853 (N_7853,N_3921,N_4038);
nor U7854 (N_7854,N_3163,N_5310);
nor U7855 (N_7855,N_5341,N_4269);
nand U7856 (N_7856,N_5658,N_4918);
nand U7857 (N_7857,N_4032,N_4987);
and U7858 (N_7858,N_4894,N_4810);
xor U7859 (N_7859,N_5405,N_5676);
or U7860 (N_7860,N_3422,N_3796);
nand U7861 (N_7861,N_5261,N_5602);
nand U7862 (N_7862,N_5217,N_5615);
nor U7863 (N_7863,N_3381,N_4640);
or U7864 (N_7864,N_5974,N_4921);
nor U7865 (N_7865,N_3747,N_3201);
and U7866 (N_7866,N_4931,N_4768);
nand U7867 (N_7867,N_4482,N_5690);
xor U7868 (N_7868,N_3909,N_4423);
or U7869 (N_7869,N_5464,N_5813);
nor U7870 (N_7870,N_3633,N_4722);
nand U7871 (N_7871,N_5149,N_4990);
nand U7872 (N_7872,N_4382,N_5304);
and U7873 (N_7873,N_5626,N_4711);
and U7874 (N_7874,N_4803,N_4155);
xnor U7875 (N_7875,N_4165,N_4113);
and U7876 (N_7876,N_5111,N_3816);
nor U7877 (N_7877,N_3467,N_5857);
or U7878 (N_7878,N_5964,N_4128);
nor U7879 (N_7879,N_5425,N_3837);
nand U7880 (N_7880,N_3211,N_5562);
xor U7881 (N_7881,N_3615,N_3172);
or U7882 (N_7882,N_5819,N_4389);
or U7883 (N_7883,N_5557,N_4506);
or U7884 (N_7884,N_5053,N_5823);
or U7885 (N_7885,N_5109,N_5694);
or U7886 (N_7886,N_4207,N_3265);
nor U7887 (N_7887,N_5954,N_3848);
and U7888 (N_7888,N_4020,N_5229);
or U7889 (N_7889,N_4024,N_5076);
and U7890 (N_7890,N_5117,N_5954);
or U7891 (N_7891,N_5854,N_4291);
nor U7892 (N_7892,N_5143,N_3531);
xnor U7893 (N_7893,N_5095,N_5317);
or U7894 (N_7894,N_3461,N_5433);
nand U7895 (N_7895,N_5285,N_4761);
nor U7896 (N_7896,N_5745,N_3680);
and U7897 (N_7897,N_5941,N_5612);
or U7898 (N_7898,N_4996,N_4098);
and U7899 (N_7899,N_5260,N_3475);
nand U7900 (N_7900,N_5077,N_3828);
or U7901 (N_7901,N_5179,N_4834);
or U7902 (N_7902,N_4592,N_3249);
or U7903 (N_7903,N_4765,N_3499);
nor U7904 (N_7904,N_5079,N_4098);
xor U7905 (N_7905,N_3228,N_3000);
or U7906 (N_7906,N_4703,N_5634);
and U7907 (N_7907,N_5436,N_5256);
and U7908 (N_7908,N_3555,N_5803);
and U7909 (N_7909,N_3788,N_5944);
nand U7910 (N_7910,N_4929,N_4276);
and U7911 (N_7911,N_5831,N_4497);
nand U7912 (N_7912,N_4526,N_3888);
xnor U7913 (N_7913,N_5230,N_4689);
nand U7914 (N_7914,N_5702,N_3615);
nor U7915 (N_7915,N_5943,N_4780);
or U7916 (N_7916,N_3200,N_3275);
nand U7917 (N_7917,N_3146,N_4774);
nor U7918 (N_7918,N_4803,N_4645);
nor U7919 (N_7919,N_3221,N_5651);
nand U7920 (N_7920,N_4727,N_3452);
and U7921 (N_7921,N_4748,N_5078);
nor U7922 (N_7922,N_5844,N_3418);
or U7923 (N_7923,N_5990,N_3726);
and U7924 (N_7924,N_4847,N_4942);
and U7925 (N_7925,N_4579,N_3830);
and U7926 (N_7926,N_3234,N_3599);
or U7927 (N_7927,N_4811,N_3298);
nor U7928 (N_7928,N_3716,N_4938);
nor U7929 (N_7929,N_5744,N_3822);
or U7930 (N_7930,N_3433,N_5716);
and U7931 (N_7931,N_4370,N_5515);
or U7932 (N_7932,N_4066,N_5254);
nor U7933 (N_7933,N_5053,N_3384);
nor U7934 (N_7934,N_5800,N_4535);
or U7935 (N_7935,N_5015,N_3119);
nor U7936 (N_7936,N_3525,N_5348);
nand U7937 (N_7937,N_3293,N_4490);
nor U7938 (N_7938,N_3024,N_3570);
and U7939 (N_7939,N_5409,N_5730);
xor U7940 (N_7940,N_3854,N_5689);
nand U7941 (N_7941,N_5952,N_5002);
or U7942 (N_7942,N_5952,N_5186);
or U7943 (N_7943,N_3513,N_4778);
or U7944 (N_7944,N_4547,N_5990);
and U7945 (N_7945,N_5067,N_5288);
and U7946 (N_7946,N_3043,N_4780);
nand U7947 (N_7947,N_3633,N_4885);
or U7948 (N_7948,N_5680,N_4274);
nand U7949 (N_7949,N_4603,N_3058);
nand U7950 (N_7950,N_5287,N_4884);
or U7951 (N_7951,N_4737,N_3692);
nor U7952 (N_7952,N_5437,N_4734);
nand U7953 (N_7953,N_5848,N_5116);
nor U7954 (N_7954,N_5981,N_3617);
nor U7955 (N_7955,N_5542,N_5432);
nand U7956 (N_7956,N_4772,N_5966);
or U7957 (N_7957,N_4172,N_3290);
nor U7958 (N_7958,N_4253,N_3576);
nand U7959 (N_7959,N_5719,N_3205);
and U7960 (N_7960,N_5594,N_5596);
or U7961 (N_7961,N_3458,N_3793);
and U7962 (N_7962,N_4961,N_3713);
and U7963 (N_7963,N_4974,N_5345);
nor U7964 (N_7964,N_5048,N_3829);
or U7965 (N_7965,N_4922,N_4155);
and U7966 (N_7966,N_5591,N_3571);
nor U7967 (N_7967,N_5835,N_3378);
or U7968 (N_7968,N_3938,N_3347);
nand U7969 (N_7969,N_4891,N_3703);
nand U7970 (N_7970,N_5369,N_3620);
or U7971 (N_7971,N_5922,N_4245);
nor U7972 (N_7972,N_5323,N_3955);
and U7973 (N_7973,N_5777,N_4669);
xnor U7974 (N_7974,N_4510,N_3297);
nand U7975 (N_7975,N_4288,N_4191);
or U7976 (N_7976,N_3443,N_3386);
and U7977 (N_7977,N_5029,N_5595);
and U7978 (N_7978,N_4083,N_4691);
nor U7979 (N_7979,N_5626,N_5400);
xnor U7980 (N_7980,N_3383,N_4059);
nand U7981 (N_7981,N_3985,N_4544);
nor U7982 (N_7982,N_5914,N_5598);
or U7983 (N_7983,N_3248,N_3683);
nand U7984 (N_7984,N_3327,N_5007);
nor U7985 (N_7985,N_4530,N_5872);
and U7986 (N_7986,N_3128,N_4964);
nand U7987 (N_7987,N_3752,N_5805);
nor U7988 (N_7988,N_4982,N_4500);
nand U7989 (N_7989,N_4101,N_4138);
nor U7990 (N_7990,N_3686,N_5093);
and U7991 (N_7991,N_5538,N_3595);
nand U7992 (N_7992,N_4594,N_5153);
or U7993 (N_7993,N_3356,N_5484);
nand U7994 (N_7994,N_3901,N_3071);
xnor U7995 (N_7995,N_3239,N_4498);
nand U7996 (N_7996,N_5465,N_3027);
nand U7997 (N_7997,N_4890,N_3612);
nand U7998 (N_7998,N_3666,N_5350);
or U7999 (N_7999,N_4197,N_3648);
nor U8000 (N_8000,N_4484,N_4648);
nor U8001 (N_8001,N_5708,N_3271);
nand U8002 (N_8002,N_3180,N_5161);
or U8003 (N_8003,N_5807,N_3320);
xnor U8004 (N_8004,N_5477,N_4850);
or U8005 (N_8005,N_4423,N_3062);
or U8006 (N_8006,N_5521,N_5780);
nor U8007 (N_8007,N_5436,N_3092);
and U8008 (N_8008,N_5977,N_5542);
or U8009 (N_8009,N_4235,N_4445);
and U8010 (N_8010,N_4023,N_4755);
nor U8011 (N_8011,N_5724,N_4176);
or U8012 (N_8012,N_3889,N_3898);
and U8013 (N_8013,N_5958,N_5353);
or U8014 (N_8014,N_5723,N_3613);
xor U8015 (N_8015,N_5584,N_3443);
nand U8016 (N_8016,N_4764,N_4356);
xor U8017 (N_8017,N_4687,N_4337);
and U8018 (N_8018,N_4085,N_5038);
nor U8019 (N_8019,N_3037,N_5537);
nand U8020 (N_8020,N_4906,N_5059);
nor U8021 (N_8021,N_5081,N_4266);
nand U8022 (N_8022,N_5771,N_3108);
or U8023 (N_8023,N_5080,N_5038);
xnor U8024 (N_8024,N_5614,N_5496);
nor U8025 (N_8025,N_3191,N_3006);
or U8026 (N_8026,N_3570,N_5729);
and U8027 (N_8027,N_5102,N_4626);
or U8028 (N_8028,N_4476,N_5925);
and U8029 (N_8029,N_4513,N_5239);
nand U8030 (N_8030,N_5488,N_3684);
or U8031 (N_8031,N_5470,N_4301);
or U8032 (N_8032,N_3721,N_5609);
or U8033 (N_8033,N_4701,N_5590);
and U8034 (N_8034,N_5787,N_5800);
nand U8035 (N_8035,N_3644,N_3484);
xnor U8036 (N_8036,N_5238,N_5453);
xnor U8037 (N_8037,N_4897,N_3123);
nor U8038 (N_8038,N_4130,N_5320);
nand U8039 (N_8039,N_3028,N_4488);
and U8040 (N_8040,N_4746,N_3912);
and U8041 (N_8041,N_4028,N_4233);
xnor U8042 (N_8042,N_5417,N_3501);
and U8043 (N_8043,N_3319,N_4806);
or U8044 (N_8044,N_3635,N_3729);
and U8045 (N_8045,N_4119,N_5165);
nor U8046 (N_8046,N_5579,N_4993);
or U8047 (N_8047,N_4696,N_4782);
or U8048 (N_8048,N_4991,N_3120);
nor U8049 (N_8049,N_3625,N_5920);
nor U8050 (N_8050,N_3191,N_5906);
xor U8051 (N_8051,N_5616,N_3985);
and U8052 (N_8052,N_3755,N_3285);
nor U8053 (N_8053,N_5333,N_3646);
nor U8054 (N_8054,N_3223,N_3966);
or U8055 (N_8055,N_4082,N_4481);
nor U8056 (N_8056,N_3970,N_5859);
and U8057 (N_8057,N_3902,N_4525);
and U8058 (N_8058,N_5895,N_4442);
or U8059 (N_8059,N_4173,N_3665);
nand U8060 (N_8060,N_3463,N_5444);
nor U8061 (N_8061,N_4360,N_3658);
nor U8062 (N_8062,N_4577,N_5995);
nand U8063 (N_8063,N_5006,N_3262);
or U8064 (N_8064,N_4987,N_3414);
nand U8065 (N_8065,N_3096,N_4498);
and U8066 (N_8066,N_3317,N_5716);
nand U8067 (N_8067,N_5795,N_3566);
and U8068 (N_8068,N_3989,N_5618);
nor U8069 (N_8069,N_4601,N_5503);
nand U8070 (N_8070,N_5132,N_3089);
nor U8071 (N_8071,N_5537,N_5928);
nand U8072 (N_8072,N_3863,N_3549);
nand U8073 (N_8073,N_3554,N_4931);
or U8074 (N_8074,N_5249,N_4397);
and U8075 (N_8075,N_5102,N_4666);
nand U8076 (N_8076,N_3057,N_3605);
xor U8077 (N_8077,N_4108,N_4286);
and U8078 (N_8078,N_3504,N_4830);
nand U8079 (N_8079,N_5290,N_5854);
or U8080 (N_8080,N_3357,N_3099);
nor U8081 (N_8081,N_3213,N_3160);
nand U8082 (N_8082,N_5610,N_3250);
nand U8083 (N_8083,N_4741,N_5480);
and U8084 (N_8084,N_4155,N_4732);
or U8085 (N_8085,N_4616,N_5347);
nor U8086 (N_8086,N_5677,N_4231);
nand U8087 (N_8087,N_5944,N_4357);
nand U8088 (N_8088,N_5745,N_4537);
and U8089 (N_8089,N_3561,N_5221);
and U8090 (N_8090,N_5690,N_3074);
or U8091 (N_8091,N_4008,N_3097);
nor U8092 (N_8092,N_4775,N_4954);
or U8093 (N_8093,N_3264,N_4024);
nor U8094 (N_8094,N_5289,N_3450);
nand U8095 (N_8095,N_5311,N_3176);
or U8096 (N_8096,N_3003,N_5140);
xor U8097 (N_8097,N_4611,N_3363);
or U8098 (N_8098,N_5508,N_4621);
nand U8099 (N_8099,N_4002,N_3408);
nand U8100 (N_8100,N_5239,N_3832);
nor U8101 (N_8101,N_5437,N_5004);
or U8102 (N_8102,N_4824,N_3067);
nand U8103 (N_8103,N_5877,N_3974);
nor U8104 (N_8104,N_4729,N_3834);
nand U8105 (N_8105,N_3625,N_4047);
nand U8106 (N_8106,N_4307,N_5495);
or U8107 (N_8107,N_5049,N_3747);
nand U8108 (N_8108,N_3120,N_4184);
nand U8109 (N_8109,N_4006,N_3644);
and U8110 (N_8110,N_5870,N_3902);
nand U8111 (N_8111,N_3093,N_5138);
xor U8112 (N_8112,N_4340,N_5190);
nand U8113 (N_8113,N_4438,N_4049);
or U8114 (N_8114,N_3676,N_4725);
xnor U8115 (N_8115,N_5421,N_4335);
nand U8116 (N_8116,N_4686,N_3986);
and U8117 (N_8117,N_5850,N_3887);
nor U8118 (N_8118,N_5632,N_3948);
or U8119 (N_8119,N_5482,N_5929);
nand U8120 (N_8120,N_4523,N_3119);
nor U8121 (N_8121,N_3558,N_3641);
nor U8122 (N_8122,N_3271,N_5521);
and U8123 (N_8123,N_4398,N_4014);
nand U8124 (N_8124,N_4441,N_3310);
or U8125 (N_8125,N_5496,N_4852);
xnor U8126 (N_8126,N_3363,N_3210);
nand U8127 (N_8127,N_5066,N_4795);
nor U8128 (N_8128,N_4462,N_4057);
xor U8129 (N_8129,N_4868,N_3843);
nor U8130 (N_8130,N_5330,N_4389);
and U8131 (N_8131,N_5238,N_5770);
and U8132 (N_8132,N_3777,N_3373);
or U8133 (N_8133,N_4151,N_5139);
and U8134 (N_8134,N_3021,N_3096);
nand U8135 (N_8135,N_3452,N_5230);
nor U8136 (N_8136,N_4129,N_5509);
or U8137 (N_8137,N_4968,N_3323);
nand U8138 (N_8138,N_5034,N_3053);
and U8139 (N_8139,N_4035,N_5092);
xor U8140 (N_8140,N_5438,N_3582);
nand U8141 (N_8141,N_3018,N_5090);
and U8142 (N_8142,N_3221,N_4367);
nor U8143 (N_8143,N_5946,N_4000);
and U8144 (N_8144,N_4451,N_3867);
and U8145 (N_8145,N_5037,N_5971);
nor U8146 (N_8146,N_4603,N_3690);
xor U8147 (N_8147,N_4896,N_5759);
and U8148 (N_8148,N_4405,N_3062);
xor U8149 (N_8149,N_5440,N_4702);
nand U8150 (N_8150,N_4055,N_4369);
or U8151 (N_8151,N_4774,N_3145);
nand U8152 (N_8152,N_5535,N_5853);
nor U8153 (N_8153,N_3727,N_4144);
nand U8154 (N_8154,N_4323,N_4794);
and U8155 (N_8155,N_5596,N_5253);
nor U8156 (N_8156,N_5434,N_3236);
or U8157 (N_8157,N_4491,N_3976);
nand U8158 (N_8158,N_4380,N_5797);
nand U8159 (N_8159,N_5678,N_4070);
or U8160 (N_8160,N_3134,N_3067);
nor U8161 (N_8161,N_4629,N_5281);
nor U8162 (N_8162,N_4387,N_4856);
or U8163 (N_8163,N_3131,N_4090);
nand U8164 (N_8164,N_4083,N_3898);
xnor U8165 (N_8165,N_4623,N_4964);
nand U8166 (N_8166,N_5486,N_3104);
nor U8167 (N_8167,N_5904,N_3529);
nand U8168 (N_8168,N_3706,N_5267);
and U8169 (N_8169,N_4071,N_5412);
xnor U8170 (N_8170,N_4013,N_3138);
or U8171 (N_8171,N_4449,N_5119);
or U8172 (N_8172,N_3960,N_3014);
and U8173 (N_8173,N_4413,N_4724);
nand U8174 (N_8174,N_3640,N_5775);
and U8175 (N_8175,N_3327,N_5485);
nor U8176 (N_8176,N_5047,N_4287);
or U8177 (N_8177,N_3898,N_3249);
nor U8178 (N_8178,N_5444,N_4137);
nand U8179 (N_8179,N_4936,N_4317);
or U8180 (N_8180,N_5035,N_3711);
xnor U8181 (N_8181,N_3048,N_4239);
and U8182 (N_8182,N_5947,N_4960);
and U8183 (N_8183,N_4820,N_4835);
or U8184 (N_8184,N_3831,N_5277);
and U8185 (N_8185,N_3543,N_5243);
and U8186 (N_8186,N_5038,N_5010);
or U8187 (N_8187,N_5716,N_3694);
or U8188 (N_8188,N_3548,N_5456);
and U8189 (N_8189,N_3613,N_4261);
or U8190 (N_8190,N_5676,N_3252);
xnor U8191 (N_8191,N_4136,N_4649);
and U8192 (N_8192,N_4847,N_3661);
or U8193 (N_8193,N_4950,N_5876);
or U8194 (N_8194,N_4353,N_3243);
nor U8195 (N_8195,N_5227,N_3939);
or U8196 (N_8196,N_3149,N_4317);
or U8197 (N_8197,N_4759,N_4640);
and U8198 (N_8198,N_4235,N_4830);
or U8199 (N_8199,N_3355,N_3841);
nand U8200 (N_8200,N_4245,N_4006);
or U8201 (N_8201,N_5870,N_4657);
or U8202 (N_8202,N_4346,N_3457);
nor U8203 (N_8203,N_3750,N_3205);
or U8204 (N_8204,N_3890,N_3593);
or U8205 (N_8205,N_4213,N_5679);
or U8206 (N_8206,N_4729,N_3588);
nand U8207 (N_8207,N_3230,N_4570);
or U8208 (N_8208,N_3098,N_3323);
xnor U8209 (N_8209,N_3662,N_5399);
nor U8210 (N_8210,N_3132,N_3097);
or U8211 (N_8211,N_4941,N_5187);
nand U8212 (N_8212,N_4966,N_4461);
xor U8213 (N_8213,N_4200,N_5341);
or U8214 (N_8214,N_3960,N_5599);
nor U8215 (N_8215,N_3929,N_5761);
nor U8216 (N_8216,N_3299,N_4147);
or U8217 (N_8217,N_5970,N_3553);
nor U8218 (N_8218,N_5933,N_5803);
nand U8219 (N_8219,N_5589,N_5081);
and U8220 (N_8220,N_4707,N_3615);
nand U8221 (N_8221,N_4753,N_4450);
nor U8222 (N_8222,N_3054,N_5405);
nor U8223 (N_8223,N_5525,N_5805);
or U8224 (N_8224,N_3834,N_5472);
and U8225 (N_8225,N_3870,N_5127);
nor U8226 (N_8226,N_4313,N_5075);
or U8227 (N_8227,N_5251,N_4660);
nand U8228 (N_8228,N_4626,N_4220);
nor U8229 (N_8229,N_4101,N_4695);
nand U8230 (N_8230,N_3654,N_3149);
nand U8231 (N_8231,N_3240,N_4763);
or U8232 (N_8232,N_3692,N_3245);
nor U8233 (N_8233,N_4464,N_3682);
or U8234 (N_8234,N_4608,N_5743);
and U8235 (N_8235,N_3492,N_5724);
and U8236 (N_8236,N_5446,N_5366);
and U8237 (N_8237,N_4847,N_5792);
nand U8238 (N_8238,N_5565,N_3260);
and U8239 (N_8239,N_4083,N_5784);
nor U8240 (N_8240,N_5449,N_5235);
and U8241 (N_8241,N_3403,N_5643);
xnor U8242 (N_8242,N_4282,N_3417);
xor U8243 (N_8243,N_3011,N_5243);
nand U8244 (N_8244,N_3769,N_5503);
and U8245 (N_8245,N_4389,N_4417);
and U8246 (N_8246,N_5033,N_3228);
and U8247 (N_8247,N_5795,N_3950);
or U8248 (N_8248,N_4661,N_3483);
nor U8249 (N_8249,N_3964,N_4106);
xnor U8250 (N_8250,N_3327,N_5915);
nand U8251 (N_8251,N_5776,N_5567);
and U8252 (N_8252,N_5221,N_4706);
or U8253 (N_8253,N_5137,N_5143);
and U8254 (N_8254,N_4693,N_3403);
and U8255 (N_8255,N_3681,N_5151);
nand U8256 (N_8256,N_4688,N_5879);
nand U8257 (N_8257,N_5620,N_4240);
and U8258 (N_8258,N_5926,N_4658);
and U8259 (N_8259,N_3179,N_5216);
nand U8260 (N_8260,N_3388,N_4402);
nor U8261 (N_8261,N_5501,N_5893);
and U8262 (N_8262,N_3466,N_4060);
and U8263 (N_8263,N_4733,N_4448);
nand U8264 (N_8264,N_3354,N_4706);
nand U8265 (N_8265,N_4544,N_5557);
nor U8266 (N_8266,N_3801,N_5900);
nand U8267 (N_8267,N_4367,N_5200);
xor U8268 (N_8268,N_3911,N_5164);
and U8269 (N_8269,N_4012,N_4130);
and U8270 (N_8270,N_5125,N_3579);
xor U8271 (N_8271,N_5178,N_4891);
and U8272 (N_8272,N_3962,N_5014);
nor U8273 (N_8273,N_3445,N_5741);
nor U8274 (N_8274,N_4208,N_3405);
nand U8275 (N_8275,N_3779,N_5450);
or U8276 (N_8276,N_5208,N_4080);
nor U8277 (N_8277,N_5317,N_3398);
or U8278 (N_8278,N_4492,N_5350);
and U8279 (N_8279,N_5498,N_5819);
or U8280 (N_8280,N_5593,N_5035);
and U8281 (N_8281,N_4010,N_3236);
nand U8282 (N_8282,N_5515,N_5252);
or U8283 (N_8283,N_5820,N_3260);
and U8284 (N_8284,N_4725,N_3296);
or U8285 (N_8285,N_3713,N_4026);
nor U8286 (N_8286,N_4340,N_5722);
nor U8287 (N_8287,N_5841,N_4507);
or U8288 (N_8288,N_5581,N_3229);
nor U8289 (N_8289,N_3001,N_4881);
nand U8290 (N_8290,N_3505,N_3259);
nand U8291 (N_8291,N_5761,N_5742);
nand U8292 (N_8292,N_4790,N_5286);
and U8293 (N_8293,N_4861,N_3531);
nand U8294 (N_8294,N_4676,N_5494);
and U8295 (N_8295,N_4237,N_4868);
xnor U8296 (N_8296,N_5934,N_5386);
nand U8297 (N_8297,N_3165,N_4224);
and U8298 (N_8298,N_4726,N_4398);
or U8299 (N_8299,N_3414,N_5014);
nand U8300 (N_8300,N_4883,N_3010);
or U8301 (N_8301,N_5995,N_4999);
nand U8302 (N_8302,N_3375,N_3968);
nor U8303 (N_8303,N_3264,N_4971);
or U8304 (N_8304,N_4366,N_3731);
nand U8305 (N_8305,N_4576,N_3611);
nand U8306 (N_8306,N_5422,N_4694);
nand U8307 (N_8307,N_4080,N_3574);
or U8308 (N_8308,N_5630,N_5799);
xnor U8309 (N_8309,N_4529,N_3142);
nand U8310 (N_8310,N_5817,N_5682);
or U8311 (N_8311,N_3784,N_4266);
nor U8312 (N_8312,N_5225,N_3429);
and U8313 (N_8313,N_4518,N_5582);
and U8314 (N_8314,N_3487,N_4257);
nor U8315 (N_8315,N_5855,N_3068);
or U8316 (N_8316,N_3422,N_4516);
or U8317 (N_8317,N_3571,N_5756);
and U8318 (N_8318,N_4679,N_3862);
nor U8319 (N_8319,N_4672,N_3323);
or U8320 (N_8320,N_4725,N_5960);
and U8321 (N_8321,N_5106,N_4243);
xor U8322 (N_8322,N_3188,N_5455);
nor U8323 (N_8323,N_4411,N_4949);
nor U8324 (N_8324,N_5089,N_4902);
xnor U8325 (N_8325,N_3855,N_4309);
nor U8326 (N_8326,N_5461,N_5582);
and U8327 (N_8327,N_4550,N_3978);
and U8328 (N_8328,N_4930,N_5962);
or U8329 (N_8329,N_5915,N_5844);
nand U8330 (N_8330,N_5668,N_3817);
nand U8331 (N_8331,N_3998,N_4019);
nor U8332 (N_8332,N_3869,N_3133);
nor U8333 (N_8333,N_5146,N_4725);
nand U8334 (N_8334,N_3729,N_5915);
xnor U8335 (N_8335,N_5762,N_3440);
nor U8336 (N_8336,N_3552,N_3162);
nand U8337 (N_8337,N_5122,N_4048);
nand U8338 (N_8338,N_4427,N_3989);
nor U8339 (N_8339,N_3074,N_4036);
nor U8340 (N_8340,N_5657,N_3468);
nor U8341 (N_8341,N_3883,N_5291);
nor U8342 (N_8342,N_5331,N_5382);
nand U8343 (N_8343,N_5794,N_5803);
and U8344 (N_8344,N_3271,N_4739);
nor U8345 (N_8345,N_4256,N_5613);
nor U8346 (N_8346,N_4194,N_3998);
and U8347 (N_8347,N_5491,N_4371);
nand U8348 (N_8348,N_4375,N_5893);
nor U8349 (N_8349,N_5231,N_3548);
nor U8350 (N_8350,N_3467,N_5989);
nand U8351 (N_8351,N_3923,N_4251);
nand U8352 (N_8352,N_3922,N_4561);
and U8353 (N_8353,N_5044,N_3274);
and U8354 (N_8354,N_3169,N_4937);
and U8355 (N_8355,N_5996,N_5637);
nand U8356 (N_8356,N_4112,N_3958);
or U8357 (N_8357,N_3545,N_3028);
and U8358 (N_8358,N_4406,N_5775);
and U8359 (N_8359,N_3679,N_5043);
and U8360 (N_8360,N_4132,N_4423);
nor U8361 (N_8361,N_5253,N_5211);
or U8362 (N_8362,N_5275,N_5538);
nor U8363 (N_8363,N_4151,N_5075);
and U8364 (N_8364,N_5594,N_4758);
or U8365 (N_8365,N_3549,N_5309);
or U8366 (N_8366,N_3382,N_3296);
and U8367 (N_8367,N_5258,N_4576);
nand U8368 (N_8368,N_3615,N_3319);
and U8369 (N_8369,N_3249,N_4567);
nor U8370 (N_8370,N_5608,N_5707);
nor U8371 (N_8371,N_4958,N_3608);
nor U8372 (N_8372,N_5142,N_5258);
nor U8373 (N_8373,N_3475,N_4268);
nor U8374 (N_8374,N_4154,N_5412);
nand U8375 (N_8375,N_5865,N_4216);
nand U8376 (N_8376,N_3194,N_5179);
nor U8377 (N_8377,N_3185,N_3902);
nor U8378 (N_8378,N_3190,N_3373);
nor U8379 (N_8379,N_3663,N_3424);
nand U8380 (N_8380,N_5579,N_3342);
nor U8381 (N_8381,N_5677,N_3573);
nor U8382 (N_8382,N_4356,N_3875);
and U8383 (N_8383,N_4789,N_5018);
nand U8384 (N_8384,N_3789,N_5360);
and U8385 (N_8385,N_5738,N_4198);
nand U8386 (N_8386,N_3893,N_5958);
or U8387 (N_8387,N_3282,N_4918);
xnor U8388 (N_8388,N_4187,N_3116);
xnor U8389 (N_8389,N_3384,N_3312);
or U8390 (N_8390,N_5684,N_4077);
and U8391 (N_8391,N_3822,N_5695);
or U8392 (N_8392,N_4705,N_5425);
nor U8393 (N_8393,N_3371,N_4528);
nand U8394 (N_8394,N_3243,N_4180);
nor U8395 (N_8395,N_3869,N_4924);
nor U8396 (N_8396,N_3831,N_4867);
nand U8397 (N_8397,N_5228,N_5095);
nand U8398 (N_8398,N_4571,N_3339);
or U8399 (N_8399,N_4126,N_5162);
xnor U8400 (N_8400,N_4722,N_4670);
nand U8401 (N_8401,N_3449,N_3249);
nor U8402 (N_8402,N_5702,N_4981);
nand U8403 (N_8403,N_4786,N_4050);
and U8404 (N_8404,N_5215,N_3918);
or U8405 (N_8405,N_3012,N_3898);
nor U8406 (N_8406,N_5931,N_4265);
or U8407 (N_8407,N_3788,N_4828);
nand U8408 (N_8408,N_4457,N_4724);
xnor U8409 (N_8409,N_5777,N_5392);
nor U8410 (N_8410,N_5475,N_3518);
or U8411 (N_8411,N_4968,N_4517);
and U8412 (N_8412,N_4618,N_3345);
nor U8413 (N_8413,N_5233,N_5435);
and U8414 (N_8414,N_3323,N_5766);
nor U8415 (N_8415,N_3957,N_4371);
nor U8416 (N_8416,N_4738,N_3615);
and U8417 (N_8417,N_3922,N_5752);
nand U8418 (N_8418,N_4447,N_5274);
nand U8419 (N_8419,N_3739,N_5616);
nor U8420 (N_8420,N_3749,N_5656);
nand U8421 (N_8421,N_5718,N_3877);
and U8422 (N_8422,N_5500,N_3303);
nor U8423 (N_8423,N_4837,N_5735);
and U8424 (N_8424,N_5946,N_4117);
nand U8425 (N_8425,N_3212,N_4986);
nand U8426 (N_8426,N_3909,N_3260);
and U8427 (N_8427,N_4304,N_3062);
nand U8428 (N_8428,N_3081,N_3241);
xnor U8429 (N_8429,N_3723,N_4284);
and U8430 (N_8430,N_3235,N_4291);
nor U8431 (N_8431,N_5676,N_3320);
and U8432 (N_8432,N_5000,N_3037);
nor U8433 (N_8433,N_3468,N_5912);
nand U8434 (N_8434,N_5904,N_5215);
nor U8435 (N_8435,N_5838,N_4172);
nand U8436 (N_8436,N_3082,N_5117);
xnor U8437 (N_8437,N_4824,N_4113);
nand U8438 (N_8438,N_3418,N_5848);
or U8439 (N_8439,N_5304,N_3781);
nor U8440 (N_8440,N_5261,N_3106);
or U8441 (N_8441,N_3320,N_5475);
and U8442 (N_8442,N_3767,N_4376);
or U8443 (N_8443,N_3515,N_3398);
or U8444 (N_8444,N_4990,N_5767);
nand U8445 (N_8445,N_5384,N_5819);
xnor U8446 (N_8446,N_3644,N_4864);
and U8447 (N_8447,N_5601,N_3362);
xnor U8448 (N_8448,N_3729,N_5547);
or U8449 (N_8449,N_5237,N_5413);
nor U8450 (N_8450,N_4570,N_5267);
nor U8451 (N_8451,N_3832,N_5082);
or U8452 (N_8452,N_4278,N_4757);
xor U8453 (N_8453,N_5919,N_3205);
or U8454 (N_8454,N_4782,N_4278);
nor U8455 (N_8455,N_4037,N_3506);
or U8456 (N_8456,N_3050,N_5600);
and U8457 (N_8457,N_4494,N_4053);
nand U8458 (N_8458,N_5051,N_3462);
nor U8459 (N_8459,N_5176,N_5234);
xnor U8460 (N_8460,N_3439,N_4270);
nand U8461 (N_8461,N_3730,N_5788);
or U8462 (N_8462,N_3520,N_5778);
nand U8463 (N_8463,N_3673,N_5311);
or U8464 (N_8464,N_3549,N_4850);
xnor U8465 (N_8465,N_5877,N_5809);
or U8466 (N_8466,N_5553,N_4377);
and U8467 (N_8467,N_3574,N_4990);
and U8468 (N_8468,N_3260,N_3195);
or U8469 (N_8469,N_4666,N_3545);
and U8470 (N_8470,N_3359,N_3707);
and U8471 (N_8471,N_3004,N_5872);
nand U8472 (N_8472,N_5781,N_3380);
nor U8473 (N_8473,N_3196,N_3211);
nand U8474 (N_8474,N_3298,N_4008);
nor U8475 (N_8475,N_5365,N_4955);
nand U8476 (N_8476,N_3013,N_4223);
or U8477 (N_8477,N_4064,N_5718);
nand U8478 (N_8478,N_4094,N_5903);
and U8479 (N_8479,N_3558,N_5742);
and U8480 (N_8480,N_5794,N_4789);
or U8481 (N_8481,N_5060,N_5541);
and U8482 (N_8482,N_4088,N_4245);
or U8483 (N_8483,N_3074,N_3580);
or U8484 (N_8484,N_4688,N_4235);
or U8485 (N_8485,N_5247,N_5529);
nor U8486 (N_8486,N_4231,N_5276);
xor U8487 (N_8487,N_3844,N_4976);
or U8488 (N_8488,N_3610,N_5202);
nor U8489 (N_8489,N_4298,N_3398);
nand U8490 (N_8490,N_3915,N_3035);
nor U8491 (N_8491,N_5639,N_3185);
xnor U8492 (N_8492,N_4325,N_5839);
and U8493 (N_8493,N_4328,N_4684);
or U8494 (N_8494,N_5307,N_3764);
or U8495 (N_8495,N_4811,N_5053);
or U8496 (N_8496,N_3217,N_4781);
and U8497 (N_8497,N_3743,N_5479);
or U8498 (N_8498,N_4017,N_5368);
nand U8499 (N_8499,N_5916,N_5882);
or U8500 (N_8500,N_5991,N_4327);
nor U8501 (N_8501,N_3231,N_4035);
nor U8502 (N_8502,N_4805,N_5053);
nand U8503 (N_8503,N_4226,N_3185);
xor U8504 (N_8504,N_3375,N_5208);
nand U8505 (N_8505,N_3396,N_3111);
or U8506 (N_8506,N_5263,N_3716);
nand U8507 (N_8507,N_3464,N_4020);
xnor U8508 (N_8508,N_3618,N_5524);
nor U8509 (N_8509,N_4322,N_5605);
or U8510 (N_8510,N_5641,N_5126);
xnor U8511 (N_8511,N_3757,N_3805);
and U8512 (N_8512,N_3912,N_4091);
nand U8513 (N_8513,N_3039,N_3982);
nand U8514 (N_8514,N_5781,N_3652);
nand U8515 (N_8515,N_4791,N_3470);
or U8516 (N_8516,N_4984,N_3572);
and U8517 (N_8517,N_5791,N_5007);
nor U8518 (N_8518,N_5513,N_4673);
nand U8519 (N_8519,N_3590,N_3276);
nand U8520 (N_8520,N_3931,N_4503);
nor U8521 (N_8521,N_3017,N_5000);
nand U8522 (N_8522,N_5204,N_3440);
nor U8523 (N_8523,N_4092,N_3930);
xor U8524 (N_8524,N_4609,N_5413);
nand U8525 (N_8525,N_5664,N_4370);
and U8526 (N_8526,N_4225,N_5463);
or U8527 (N_8527,N_4261,N_3800);
nor U8528 (N_8528,N_5734,N_5242);
and U8529 (N_8529,N_3687,N_5846);
nand U8530 (N_8530,N_4388,N_5849);
nand U8531 (N_8531,N_5993,N_5216);
xor U8532 (N_8532,N_4653,N_3997);
and U8533 (N_8533,N_4326,N_3538);
or U8534 (N_8534,N_4383,N_4450);
and U8535 (N_8535,N_5597,N_5327);
nor U8536 (N_8536,N_4037,N_3644);
and U8537 (N_8537,N_4839,N_3285);
nor U8538 (N_8538,N_3613,N_3832);
nand U8539 (N_8539,N_3028,N_4570);
nor U8540 (N_8540,N_5378,N_3251);
nor U8541 (N_8541,N_4681,N_5725);
and U8542 (N_8542,N_5966,N_5567);
nor U8543 (N_8543,N_3068,N_4880);
and U8544 (N_8544,N_3732,N_4062);
xnor U8545 (N_8545,N_5060,N_3522);
and U8546 (N_8546,N_4278,N_3286);
and U8547 (N_8547,N_4061,N_4943);
xnor U8548 (N_8548,N_5512,N_5364);
nand U8549 (N_8549,N_3371,N_5661);
xor U8550 (N_8550,N_4138,N_4862);
nand U8551 (N_8551,N_4743,N_5098);
nand U8552 (N_8552,N_3579,N_4483);
or U8553 (N_8553,N_4135,N_4303);
and U8554 (N_8554,N_4484,N_3586);
nor U8555 (N_8555,N_4445,N_5218);
or U8556 (N_8556,N_5720,N_3620);
nand U8557 (N_8557,N_3949,N_3810);
and U8558 (N_8558,N_3550,N_5956);
nand U8559 (N_8559,N_5545,N_5018);
or U8560 (N_8560,N_5697,N_4055);
xor U8561 (N_8561,N_4943,N_3191);
or U8562 (N_8562,N_4603,N_5483);
nor U8563 (N_8563,N_5155,N_5756);
nand U8564 (N_8564,N_5461,N_5876);
and U8565 (N_8565,N_5281,N_4593);
nand U8566 (N_8566,N_3305,N_4782);
nand U8567 (N_8567,N_4983,N_3901);
nor U8568 (N_8568,N_4447,N_3579);
and U8569 (N_8569,N_3247,N_3584);
and U8570 (N_8570,N_5241,N_3537);
nand U8571 (N_8571,N_5669,N_5702);
and U8572 (N_8572,N_5496,N_5232);
and U8573 (N_8573,N_4063,N_3591);
nand U8574 (N_8574,N_4607,N_5719);
nand U8575 (N_8575,N_5751,N_3867);
nand U8576 (N_8576,N_5346,N_3712);
nand U8577 (N_8577,N_5391,N_4321);
or U8578 (N_8578,N_3122,N_3739);
and U8579 (N_8579,N_5501,N_5261);
nand U8580 (N_8580,N_3009,N_4030);
and U8581 (N_8581,N_4186,N_5978);
nor U8582 (N_8582,N_5795,N_5551);
nor U8583 (N_8583,N_5034,N_4660);
nor U8584 (N_8584,N_4163,N_3899);
nand U8585 (N_8585,N_3522,N_4043);
or U8586 (N_8586,N_3908,N_5600);
or U8587 (N_8587,N_3682,N_5132);
and U8588 (N_8588,N_4551,N_5599);
and U8589 (N_8589,N_4029,N_5123);
nor U8590 (N_8590,N_4129,N_3891);
nand U8591 (N_8591,N_3166,N_3074);
nor U8592 (N_8592,N_4466,N_4546);
xnor U8593 (N_8593,N_5229,N_5381);
and U8594 (N_8594,N_4176,N_5225);
and U8595 (N_8595,N_4242,N_3151);
and U8596 (N_8596,N_5975,N_4238);
nor U8597 (N_8597,N_5884,N_5500);
and U8598 (N_8598,N_4958,N_3417);
or U8599 (N_8599,N_4289,N_4985);
or U8600 (N_8600,N_3013,N_3291);
xnor U8601 (N_8601,N_4207,N_3599);
or U8602 (N_8602,N_3112,N_3868);
nand U8603 (N_8603,N_5142,N_5475);
and U8604 (N_8604,N_5387,N_4890);
nor U8605 (N_8605,N_4755,N_4696);
or U8606 (N_8606,N_5562,N_3616);
or U8607 (N_8607,N_3726,N_3085);
nand U8608 (N_8608,N_5377,N_5791);
nand U8609 (N_8609,N_4856,N_4563);
xor U8610 (N_8610,N_4452,N_5185);
or U8611 (N_8611,N_3364,N_3003);
or U8612 (N_8612,N_5500,N_5774);
nor U8613 (N_8613,N_5111,N_3829);
or U8614 (N_8614,N_4573,N_3182);
and U8615 (N_8615,N_3196,N_3429);
or U8616 (N_8616,N_3390,N_5530);
nor U8617 (N_8617,N_4910,N_4808);
or U8618 (N_8618,N_4768,N_4619);
or U8619 (N_8619,N_3243,N_4961);
and U8620 (N_8620,N_4224,N_5205);
nor U8621 (N_8621,N_5779,N_5976);
nand U8622 (N_8622,N_3789,N_4447);
or U8623 (N_8623,N_5396,N_3191);
nor U8624 (N_8624,N_3635,N_3445);
and U8625 (N_8625,N_3073,N_4956);
or U8626 (N_8626,N_3516,N_4523);
xor U8627 (N_8627,N_5584,N_5886);
or U8628 (N_8628,N_4789,N_5300);
and U8629 (N_8629,N_5754,N_4224);
and U8630 (N_8630,N_3244,N_3534);
and U8631 (N_8631,N_3552,N_4968);
or U8632 (N_8632,N_3793,N_3502);
or U8633 (N_8633,N_4463,N_3404);
and U8634 (N_8634,N_3972,N_5126);
nor U8635 (N_8635,N_3794,N_5362);
and U8636 (N_8636,N_3390,N_5698);
or U8637 (N_8637,N_5773,N_4809);
nand U8638 (N_8638,N_4622,N_3017);
or U8639 (N_8639,N_3947,N_3586);
nor U8640 (N_8640,N_3675,N_3205);
and U8641 (N_8641,N_3463,N_5647);
and U8642 (N_8642,N_3368,N_3288);
xor U8643 (N_8643,N_5643,N_5836);
and U8644 (N_8644,N_4888,N_3869);
and U8645 (N_8645,N_3062,N_5183);
nand U8646 (N_8646,N_3084,N_5106);
nand U8647 (N_8647,N_4952,N_3775);
nor U8648 (N_8648,N_5387,N_3995);
nor U8649 (N_8649,N_5258,N_3551);
and U8650 (N_8650,N_4609,N_3519);
or U8651 (N_8651,N_5242,N_4268);
or U8652 (N_8652,N_5032,N_4007);
nand U8653 (N_8653,N_3571,N_3561);
nand U8654 (N_8654,N_4600,N_4937);
nand U8655 (N_8655,N_5441,N_5568);
nand U8656 (N_8656,N_5023,N_4278);
or U8657 (N_8657,N_3913,N_3798);
nor U8658 (N_8658,N_5523,N_5151);
nor U8659 (N_8659,N_3511,N_4171);
or U8660 (N_8660,N_5649,N_4564);
and U8661 (N_8661,N_5347,N_5101);
nand U8662 (N_8662,N_4650,N_3589);
nor U8663 (N_8663,N_3738,N_5973);
or U8664 (N_8664,N_3013,N_5864);
or U8665 (N_8665,N_4772,N_4609);
nand U8666 (N_8666,N_5961,N_5578);
nor U8667 (N_8667,N_5562,N_5122);
xor U8668 (N_8668,N_3148,N_5643);
and U8669 (N_8669,N_3512,N_5897);
or U8670 (N_8670,N_4061,N_3934);
and U8671 (N_8671,N_3703,N_3794);
nand U8672 (N_8672,N_3578,N_4524);
or U8673 (N_8673,N_4228,N_4485);
nor U8674 (N_8674,N_3077,N_5174);
or U8675 (N_8675,N_4864,N_5077);
nor U8676 (N_8676,N_3970,N_4692);
and U8677 (N_8677,N_4834,N_5810);
xor U8678 (N_8678,N_4452,N_4498);
nand U8679 (N_8679,N_5851,N_3408);
and U8680 (N_8680,N_4619,N_5382);
nand U8681 (N_8681,N_5656,N_5581);
nor U8682 (N_8682,N_5999,N_4736);
nand U8683 (N_8683,N_4510,N_3708);
and U8684 (N_8684,N_3524,N_3209);
or U8685 (N_8685,N_4386,N_5978);
nand U8686 (N_8686,N_4039,N_3986);
and U8687 (N_8687,N_3094,N_4801);
and U8688 (N_8688,N_5314,N_4940);
nand U8689 (N_8689,N_4872,N_5576);
nor U8690 (N_8690,N_3871,N_5046);
xnor U8691 (N_8691,N_4335,N_5439);
or U8692 (N_8692,N_4172,N_3839);
nand U8693 (N_8693,N_4136,N_5268);
or U8694 (N_8694,N_5924,N_4869);
and U8695 (N_8695,N_4369,N_4540);
nor U8696 (N_8696,N_5052,N_4277);
nand U8697 (N_8697,N_3325,N_3256);
xnor U8698 (N_8698,N_5059,N_4625);
xnor U8699 (N_8699,N_5461,N_3005);
nor U8700 (N_8700,N_4208,N_5794);
and U8701 (N_8701,N_3148,N_3046);
or U8702 (N_8702,N_5640,N_4080);
and U8703 (N_8703,N_3798,N_5738);
xor U8704 (N_8704,N_3241,N_4512);
and U8705 (N_8705,N_3277,N_3956);
nand U8706 (N_8706,N_3047,N_5235);
nand U8707 (N_8707,N_5907,N_3729);
nor U8708 (N_8708,N_3883,N_3493);
nor U8709 (N_8709,N_3767,N_3318);
or U8710 (N_8710,N_4738,N_3987);
and U8711 (N_8711,N_5738,N_5395);
and U8712 (N_8712,N_5174,N_3943);
nor U8713 (N_8713,N_5019,N_3388);
nor U8714 (N_8714,N_5741,N_4269);
nand U8715 (N_8715,N_5903,N_4114);
and U8716 (N_8716,N_4102,N_5240);
and U8717 (N_8717,N_5577,N_4902);
or U8718 (N_8718,N_5715,N_4981);
or U8719 (N_8719,N_5500,N_5340);
xnor U8720 (N_8720,N_5583,N_4929);
nor U8721 (N_8721,N_5198,N_4678);
and U8722 (N_8722,N_5451,N_4274);
nor U8723 (N_8723,N_3655,N_4292);
xor U8724 (N_8724,N_3720,N_5258);
nand U8725 (N_8725,N_4542,N_4534);
or U8726 (N_8726,N_3221,N_4003);
and U8727 (N_8727,N_5002,N_4181);
or U8728 (N_8728,N_5925,N_5926);
nor U8729 (N_8729,N_4935,N_4888);
xnor U8730 (N_8730,N_3426,N_3986);
or U8731 (N_8731,N_4967,N_3246);
and U8732 (N_8732,N_3301,N_3024);
nand U8733 (N_8733,N_3415,N_4318);
or U8734 (N_8734,N_4467,N_5717);
or U8735 (N_8735,N_5999,N_4557);
and U8736 (N_8736,N_3647,N_5792);
or U8737 (N_8737,N_5590,N_4752);
xnor U8738 (N_8738,N_5406,N_5229);
or U8739 (N_8739,N_4047,N_3955);
nor U8740 (N_8740,N_4492,N_4592);
or U8741 (N_8741,N_3745,N_5976);
nor U8742 (N_8742,N_5016,N_4411);
nor U8743 (N_8743,N_3831,N_5560);
xor U8744 (N_8744,N_5439,N_3250);
and U8745 (N_8745,N_3818,N_4769);
nor U8746 (N_8746,N_4318,N_5491);
nand U8747 (N_8747,N_5535,N_5824);
nor U8748 (N_8748,N_5644,N_5385);
and U8749 (N_8749,N_3194,N_5938);
or U8750 (N_8750,N_5770,N_4830);
nand U8751 (N_8751,N_3402,N_5574);
nand U8752 (N_8752,N_3659,N_4702);
or U8753 (N_8753,N_3843,N_4136);
or U8754 (N_8754,N_5066,N_3398);
xor U8755 (N_8755,N_3516,N_3618);
xnor U8756 (N_8756,N_4505,N_3542);
or U8757 (N_8757,N_3939,N_5723);
or U8758 (N_8758,N_4809,N_3565);
and U8759 (N_8759,N_5894,N_4440);
nand U8760 (N_8760,N_4307,N_3210);
nor U8761 (N_8761,N_5101,N_5480);
nand U8762 (N_8762,N_3517,N_5385);
or U8763 (N_8763,N_3983,N_5208);
xnor U8764 (N_8764,N_5936,N_4970);
nand U8765 (N_8765,N_5801,N_3333);
or U8766 (N_8766,N_5552,N_3372);
nand U8767 (N_8767,N_3787,N_5515);
xor U8768 (N_8768,N_5827,N_3503);
nand U8769 (N_8769,N_4411,N_4546);
nand U8770 (N_8770,N_4139,N_5771);
nand U8771 (N_8771,N_4445,N_3351);
or U8772 (N_8772,N_4000,N_3382);
nor U8773 (N_8773,N_3035,N_5310);
nand U8774 (N_8774,N_5499,N_4036);
nor U8775 (N_8775,N_3640,N_5280);
or U8776 (N_8776,N_5215,N_4920);
nor U8777 (N_8777,N_3263,N_4085);
nand U8778 (N_8778,N_5536,N_4892);
xnor U8779 (N_8779,N_5614,N_5084);
nand U8780 (N_8780,N_3022,N_3804);
or U8781 (N_8781,N_5941,N_3984);
nor U8782 (N_8782,N_4110,N_3084);
or U8783 (N_8783,N_4411,N_5296);
nor U8784 (N_8784,N_5518,N_5669);
xnor U8785 (N_8785,N_4121,N_4399);
nor U8786 (N_8786,N_3085,N_5406);
and U8787 (N_8787,N_3135,N_3838);
nand U8788 (N_8788,N_3273,N_3761);
or U8789 (N_8789,N_4163,N_5343);
and U8790 (N_8790,N_3215,N_5240);
or U8791 (N_8791,N_5454,N_4263);
xor U8792 (N_8792,N_4554,N_3398);
or U8793 (N_8793,N_4444,N_4512);
nor U8794 (N_8794,N_3753,N_5311);
and U8795 (N_8795,N_5490,N_5735);
and U8796 (N_8796,N_5147,N_4425);
or U8797 (N_8797,N_5303,N_4025);
nor U8798 (N_8798,N_4173,N_5477);
nand U8799 (N_8799,N_5310,N_3803);
nand U8800 (N_8800,N_5756,N_3326);
nand U8801 (N_8801,N_3559,N_3347);
and U8802 (N_8802,N_4439,N_4048);
nand U8803 (N_8803,N_5692,N_5420);
and U8804 (N_8804,N_5345,N_5215);
nor U8805 (N_8805,N_4200,N_3492);
or U8806 (N_8806,N_3178,N_3149);
and U8807 (N_8807,N_3750,N_4116);
nor U8808 (N_8808,N_5685,N_5492);
nand U8809 (N_8809,N_4305,N_3444);
or U8810 (N_8810,N_5389,N_5817);
xor U8811 (N_8811,N_3928,N_4400);
and U8812 (N_8812,N_5169,N_4421);
or U8813 (N_8813,N_3045,N_5104);
and U8814 (N_8814,N_4098,N_3996);
nand U8815 (N_8815,N_4578,N_4276);
nor U8816 (N_8816,N_3142,N_4894);
and U8817 (N_8817,N_4007,N_5609);
or U8818 (N_8818,N_3708,N_3260);
nand U8819 (N_8819,N_5434,N_5796);
nor U8820 (N_8820,N_4635,N_5096);
nor U8821 (N_8821,N_4263,N_5394);
or U8822 (N_8822,N_3156,N_5007);
and U8823 (N_8823,N_5080,N_3911);
or U8824 (N_8824,N_3108,N_5373);
nor U8825 (N_8825,N_4740,N_3082);
or U8826 (N_8826,N_3859,N_5229);
nor U8827 (N_8827,N_4212,N_5294);
nor U8828 (N_8828,N_5336,N_4284);
xor U8829 (N_8829,N_4564,N_4962);
and U8830 (N_8830,N_4523,N_3149);
or U8831 (N_8831,N_5241,N_3358);
xor U8832 (N_8832,N_3557,N_5250);
or U8833 (N_8833,N_5111,N_3504);
nand U8834 (N_8834,N_5277,N_5749);
xnor U8835 (N_8835,N_3437,N_4424);
or U8836 (N_8836,N_5720,N_4235);
and U8837 (N_8837,N_4791,N_3757);
nor U8838 (N_8838,N_4486,N_4113);
nor U8839 (N_8839,N_5084,N_3629);
nand U8840 (N_8840,N_5590,N_3962);
and U8841 (N_8841,N_3643,N_4126);
and U8842 (N_8842,N_5981,N_5755);
nor U8843 (N_8843,N_3876,N_5795);
and U8844 (N_8844,N_5132,N_4674);
nor U8845 (N_8845,N_4293,N_5361);
nand U8846 (N_8846,N_3955,N_5180);
or U8847 (N_8847,N_5137,N_4460);
or U8848 (N_8848,N_3997,N_4992);
nand U8849 (N_8849,N_3636,N_5732);
or U8850 (N_8850,N_3037,N_5952);
nand U8851 (N_8851,N_5831,N_4878);
or U8852 (N_8852,N_4530,N_5782);
or U8853 (N_8853,N_4763,N_3258);
nor U8854 (N_8854,N_4792,N_5752);
nor U8855 (N_8855,N_4456,N_4158);
nor U8856 (N_8856,N_3250,N_3754);
and U8857 (N_8857,N_4517,N_5273);
and U8858 (N_8858,N_5352,N_4205);
nor U8859 (N_8859,N_3316,N_4918);
and U8860 (N_8860,N_3271,N_5963);
nor U8861 (N_8861,N_3088,N_4806);
nor U8862 (N_8862,N_5670,N_4125);
and U8863 (N_8863,N_3384,N_4234);
or U8864 (N_8864,N_5759,N_3816);
nand U8865 (N_8865,N_5757,N_5351);
or U8866 (N_8866,N_5263,N_3361);
nand U8867 (N_8867,N_3968,N_3791);
and U8868 (N_8868,N_3549,N_4616);
nor U8869 (N_8869,N_3601,N_3055);
nand U8870 (N_8870,N_4296,N_5677);
or U8871 (N_8871,N_5692,N_5053);
or U8872 (N_8872,N_4973,N_4063);
and U8873 (N_8873,N_5801,N_3485);
nor U8874 (N_8874,N_5831,N_4437);
and U8875 (N_8875,N_4591,N_3224);
xor U8876 (N_8876,N_5585,N_4148);
or U8877 (N_8877,N_5026,N_3198);
nor U8878 (N_8878,N_3963,N_3159);
nand U8879 (N_8879,N_4174,N_5997);
or U8880 (N_8880,N_5822,N_4389);
nor U8881 (N_8881,N_4943,N_5997);
nand U8882 (N_8882,N_5467,N_5669);
and U8883 (N_8883,N_3149,N_4647);
nand U8884 (N_8884,N_4532,N_5961);
xnor U8885 (N_8885,N_3260,N_5901);
and U8886 (N_8886,N_4143,N_3977);
or U8887 (N_8887,N_3187,N_3428);
nand U8888 (N_8888,N_3508,N_5120);
or U8889 (N_8889,N_5353,N_5220);
or U8890 (N_8890,N_3981,N_4835);
or U8891 (N_8891,N_5482,N_3618);
and U8892 (N_8892,N_4422,N_3017);
nand U8893 (N_8893,N_4110,N_5561);
nand U8894 (N_8894,N_4881,N_3579);
nand U8895 (N_8895,N_5952,N_4539);
nor U8896 (N_8896,N_3176,N_3256);
nor U8897 (N_8897,N_4968,N_3776);
xor U8898 (N_8898,N_4410,N_5172);
and U8899 (N_8899,N_5163,N_5954);
nand U8900 (N_8900,N_5887,N_4966);
xnor U8901 (N_8901,N_5337,N_3918);
nand U8902 (N_8902,N_5403,N_3023);
or U8903 (N_8903,N_3560,N_4791);
nor U8904 (N_8904,N_5101,N_3889);
or U8905 (N_8905,N_5287,N_3386);
nor U8906 (N_8906,N_3975,N_3247);
or U8907 (N_8907,N_5489,N_5942);
and U8908 (N_8908,N_5356,N_5908);
or U8909 (N_8909,N_3385,N_3620);
nor U8910 (N_8910,N_3054,N_3482);
xor U8911 (N_8911,N_5125,N_3927);
or U8912 (N_8912,N_3923,N_5349);
and U8913 (N_8913,N_5419,N_3483);
or U8914 (N_8914,N_5701,N_5366);
and U8915 (N_8915,N_5287,N_5763);
nand U8916 (N_8916,N_4350,N_4157);
nand U8917 (N_8917,N_4054,N_3723);
nand U8918 (N_8918,N_4696,N_5340);
nand U8919 (N_8919,N_3953,N_3997);
xor U8920 (N_8920,N_5732,N_4310);
and U8921 (N_8921,N_4617,N_4419);
nor U8922 (N_8922,N_4507,N_4999);
xor U8923 (N_8923,N_3569,N_4058);
or U8924 (N_8924,N_3264,N_3800);
or U8925 (N_8925,N_5710,N_3357);
xor U8926 (N_8926,N_5357,N_5347);
or U8927 (N_8927,N_5343,N_5068);
nor U8928 (N_8928,N_4554,N_3137);
and U8929 (N_8929,N_3524,N_3277);
nand U8930 (N_8930,N_3004,N_3474);
or U8931 (N_8931,N_3302,N_3079);
xor U8932 (N_8932,N_5831,N_4285);
xor U8933 (N_8933,N_4799,N_3162);
xnor U8934 (N_8934,N_3673,N_4288);
nor U8935 (N_8935,N_5724,N_5676);
nor U8936 (N_8936,N_3426,N_4754);
and U8937 (N_8937,N_4001,N_3103);
and U8938 (N_8938,N_5320,N_4754);
nor U8939 (N_8939,N_5101,N_4550);
and U8940 (N_8940,N_3212,N_5341);
nand U8941 (N_8941,N_5537,N_5742);
nand U8942 (N_8942,N_3826,N_3075);
nand U8943 (N_8943,N_4964,N_3978);
nor U8944 (N_8944,N_4915,N_3175);
and U8945 (N_8945,N_5867,N_4098);
and U8946 (N_8946,N_5246,N_3637);
xor U8947 (N_8947,N_5058,N_5131);
nand U8948 (N_8948,N_4014,N_4924);
or U8949 (N_8949,N_4410,N_4191);
or U8950 (N_8950,N_4546,N_3761);
nor U8951 (N_8951,N_5812,N_4700);
xor U8952 (N_8952,N_4812,N_3081);
nand U8953 (N_8953,N_5202,N_5953);
and U8954 (N_8954,N_5710,N_3772);
or U8955 (N_8955,N_5649,N_4925);
or U8956 (N_8956,N_4830,N_5057);
nor U8957 (N_8957,N_5067,N_5385);
and U8958 (N_8958,N_5992,N_3644);
nor U8959 (N_8959,N_3041,N_3421);
and U8960 (N_8960,N_4738,N_5470);
xnor U8961 (N_8961,N_4806,N_4181);
or U8962 (N_8962,N_5582,N_5415);
or U8963 (N_8963,N_4155,N_5840);
or U8964 (N_8964,N_4265,N_5225);
nor U8965 (N_8965,N_3072,N_3915);
and U8966 (N_8966,N_3546,N_4736);
or U8967 (N_8967,N_5019,N_5670);
or U8968 (N_8968,N_4637,N_4240);
nand U8969 (N_8969,N_3537,N_4200);
or U8970 (N_8970,N_3616,N_5687);
nand U8971 (N_8971,N_5733,N_4577);
nand U8972 (N_8972,N_5049,N_3991);
nor U8973 (N_8973,N_4961,N_3642);
nand U8974 (N_8974,N_3063,N_5413);
nor U8975 (N_8975,N_4939,N_4374);
nor U8976 (N_8976,N_5233,N_4793);
nand U8977 (N_8977,N_5079,N_4597);
and U8978 (N_8978,N_5676,N_5325);
and U8979 (N_8979,N_3545,N_5176);
nor U8980 (N_8980,N_5741,N_4699);
nor U8981 (N_8981,N_3479,N_5676);
nor U8982 (N_8982,N_4635,N_4310);
nor U8983 (N_8983,N_5486,N_3627);
or U8984 (N_8984,N_3915,N_3358);
and U8985 (N_8985,N_3650,N_4807);
nor U8986 (N_8986,N_3272,N_3558);
and U8987 (N_8987,N_4231,N_5471);
or U8988 (N_8988,N_5976,N_5077);
or U8989 (N_8989,N_3641,N_3716);
and U8990 (N_8990,N_3596,N_3965);
or U8991 (N_8991,N_3523,N_3613);
or U8992 (N_8992,N_3589,N_5500);
nor U8993 (N_8993,N_3380,N_4359);
or U8994 (N_8994,N_3626,N_5662);
or U8995 (N_8995,N_3831,N_3208);
nand U8996 (N_8996,N_5235,N_3233);
and U8997 (N_8997,N_5859,N_4823);
and U8998 (N_8998,N_4942,N_3325);
or U8999 (N_8999,N_4524,N_3476);
or U9000 (N_9000,N_6826,N_6373);
xnor U9001 (N_9001,N_6994,N_7813);
nand U9002 (N_9002,N_6509,N_8519);
nand U9003 (N_9003,N_7402,N_7706);
nand U9004 (N_9004,N_8471,N_8634);
nor U9005 (N_9005,N_7640,N_6828);
and U9006 (N_9006,N_7908,N_7188);
nor U9007 (N_9007,N_7973,N_6011);
and U9008 (N_9008,N_8762,N_7148);
and U9009 (N_9009,N_6553,N_7222);
nor U9010 (N_9010,N_8728,N_8518);
nor U9011 (N_9011,N_7626,N_6411);
nor U9012 (N_9012,N_8100,N_8124);
and U9013 (N_9013,N_7763,N_7038);
and U9014 (N_9014,N_8313,N_7975);
or U9015 (N_9015,N_7514,N_8995);
nand U9016 (N_9016,N_6135,N_8337);
or U9017 (N_9017,N_8073,N_6948);
nand U9018 (N_9018,N_8635,N_8404);
nor U9019 (N_9019,N_6380,N_6143);
xnor U9020 (N_9020,N_8132,N_7823);
nand U9021 (N_9021,N_8600,N_8269);
nor U9022 (N_9022,N_7886,N_8862);
or U9023 (N_9023,N_8060,N_8240);
nand U9024 (N_9024,N_8914,N_8382);
and U9025 (N_9025,N_7010,N_7515);
xnor U9026 (N_9026,N_7866,N_7169);
nand U9027 (N_9027,N_7898,N_8553);
nand U9028 (N_9028,N_6110,N_7360);
or U9029 (N_9029,N_6600,N_6378);
nor U9030 (N_9030,N_6657,N_8890);
and U9031 (N_9031,N_7569,N_6158);
nor U9032 (N_9032,N_6480,N_6671);
and U9033 (N_9033,N_8896,N_6598);
nor U9034 (N_9034,N_7059,N_6286);
nand U9035 (N_9035,N_6140,N_6257);
nor U9036 (N_9036,N_6961,N_6099);
or U9037 (N_9037,N_7998,N_8733);
nor U9038 (N_9038,N_7115,N_6415);
xnor U9039 (N_9039,N_8984,N_8388);
and U9040 (N_9040,N_6796,N_8602);
xor U9041 (N_9041,N_6417,N_7372);
nor U9042 (N_9042,N_6637,N_8442);
nor U9043 (N_9043,N_7939,N_7433);
nor U9044 (N_9044,N_7214,N_6429);
nand U9045 (N_9045,N_8145,N_7534);
nor U9046 (N_9046,N_8411,N_6683);
or U9047 (N_9047,N_6303,N_6245);
nand U9048 (N_9048,N_6564,N_7604);
nor U9049 (N_9049,N_6336,N_8129);
nor U9050 (N_9050,N_7272,N_6879);
nand U9051 (N_9051,N_8689,N_6269);
and U9052 (N_9052,N_7710,N_8090);
xor U9053 (N_9053,N_7841,N_6547);
nor U9054 (N_9054,N_8034,N_8538);
and U9055 (N_9055,N_6096,N_6439);
nor U9056 (N_9056,N_6492,N_8247);
and U9057 (N_9057,N_8118,N_6399);
or U9058 (N_9058,N_7957,N_7619);
and U9059 (N_9059,N_6333,N_6406);
nor U9060 (N_9060,N_6473,N_6891);
and U9061 (N_9061,N_8649,N_6074);
nand U9062 (N_9062,N_7458,N_6702);
nand U9063 (N_9063,N_8112,N_6706);
and U9064 (N_9064,N_6493,N_8128);
xor U9065 (N_9065,N_7613,N_6832);
nor U9066 (N_9066,N_6265,N_8727);
nand U9067 (N_9067,N_6460,N_6264);
and U9068 (N_9068,N_7774,N_8378);
nand U9069 (N_9069,N_7137,N_7971);
nand U9070 (N_9070,N_7002,N_8005);
or U9071 (N_9071,N_6347,N_8393);
nor U9072 (N_9072,N_6216,N_7996);
nor U9073 (N_9073,N_8324,N_6240);
or U9074 (N_9074,N_8398,N_7063);
nor U9075 (N_9075,N_6113,N_6023);
xor U9076 (N_9076,N_8966,N_6782);
nor U9077 (N_9077,N_7902,N_7885);
nand U9078 (N_9078,N_7437,N_8929);
nand U9079 (N_9079,N_6822,N_7098);
or U9080 (N_9080,N_7209,N_6328);
and U9081 (N_9081,N_8250,N_8109);
or U9082 (N_9082,N_6050,N_6164);
nand U9083 (N_9083,N_7788,N_6990);
or U9084 (N_9084,N_7199,N_8924);
nor U9085 (N_9085,N_8584,N_6072);
and U9086 (N_9086,N_6563,N_6424);
xnor U9087 (N_9087,N_6397,N_6794);
or U9088 (N_9088,N_8195,N_7612);
xnor U9089 (N_9089,N_7691,N_6668);
or U9090 (N_9090,N_7698,N_6019);
nor U9091 (N_9091,N_8556,N_7171);
nand U9092 (N_9092,N_8040,N_6066);
and U9093 (N_9093,N_8791,N_7665);
or U9094 (N_9094,N_8687,N_8930);
nand U9095 (N_9095,N_8991,N_6043);
nand U9096 (N_9096,N_6645,N_8714);
nand U9097 (N_9097,N_6490,N_6345);
nor U9098 (N_9098,N_8350,N_6958);
nor U9099 (N_9099,N_6881,N_6360);
or U9100 (N_9100,N_8940,N_7662);
nor U9101 (N_9101,N_7532,N_8778);
or U9102 (N_9102,N_7088,N_7268);
and U9103 (N_9103,N_8598,N_7663);
or U9104 (N_9104,N_7307,N_6992);
and U9105 (N_9105,N_6778,N_7332);
or U9106 (N_9106,N_8773,N_6758);
and U9107 (N_9107,N_7164,N_6418);
and U9108 (N_9108,N_8945,N_6372);
or U9109 (N_9109,N_8867,N_6403);
or U9110 (N_9110,N_7993,N_8531);
nor U9111 (N_9111,N_6849,N_6747);
and U9112 (N_9112,N_7543,N_7771);
or U9113 (N_9113,N_8296,N_6398);
nand U9114 (N_9114,N_7225,N_6394);
or U9115 (N_9115,N_6151,N_7986);
xor U9116 (N_9116,N_8986,N_6389);
nand U9117 (N_9117,N_6463,N_7039);
or U9118 (N_9118,N_8744,N_6582);
nand U9119 (N_9119,N_6540,N_7487);
nand U9120 (N_9120,N_6344,N_8459);
or U9121 (N_9121,N_8190,N_7347);
and U9122 (N_9122,N_8879,N_6251);
and U9123 (N_9123,N_6478,N_8506);
and U9124 (N_9124,N_6745,N_6369);
nand U9125 (N_9125,N_8285,N_7364);
nand U9126 (N_9126,N_8780,N_8811);
nor U9127 (N_9127,N_7995,N_7477);
or U9128 (N_9128,N_6341,N_7353);
nand U9129 (N_9129,N_7557,N_6890);
nand U9130 (N_9130,N_6972,N_6756);
or U9131 (N_9131,N_6400,N_7559);
nor U9132 (N_9132,N_6425,N_6712);
and U9133 (N_9133,N_8782,N_7976);
or U9134 (N_9134,N_8505,N_6029);
xnor U9135 (N_9135,N_6438,N_7451);
and U9136 (N_9136,N_8310,N_7285);
and U9137 (N_9137,N_7684,N_7349);
nor U9138 (N_9138,N_8770,N_7642);
nand U9139 (N_9139,N_8814,N_7843);
nor U9140 (N_9140,N_7439,N_7562);
nor U9141 (N_9141,N_7953,N_8695);
nand U9142 (N_9142,N_8209,N_6759);
or U9143 (N_9143,N_6532,N_7201);
nand U9144 (N_9144,N_7611,N_8069);
or U9145 (N_9145,N_6453,N_7988);
or U9146 (N_9146,N_6988,N_7831);
nor U9147 (N_9147,N_7297,N_8655);
or U9148 (N_9148,N_6277,N_8332);
or U9149 (N_9149,N_7978,N_6451);
nand U9150 (N_9150,N_8444,N_7262);
and U9151 (N_9151,N_7019,N_8044);
and U9152 (N_9152,N_6193,N_7119);
nor U9153 (N_9153,N_6491,N_7577);
nor U9154 (N_9154,N_7983,N_7529);
and U9155 (N_9155,N_7591,N_8164);
and U9156 (N_9156,N_7936,N_6833);
or U9157 (N_9157,N_6725,N_8371);
and U9158 (N_9158,N_6648,N_7354);
nand U9159 (N_9159,N_8148,N_6496);
nor U9160 (N_9160,N_6044,N_6253);
and U9161 (N_9161,N_7784,N_7455);
or U9162 (N_9162,N_8723,N_7609);
nor U9163 (N_9163,N_8386,N_6984);
and U9164 (N_9164,N_8882,N_7549);
nand U9165 (N_9165,N_7842,N_7153);
nor U9166 (N_9166,N_8274,N_8622);
xnor U9167 (N_9167,N_6577,N_8554);
and U9168 (N_9168,N_8970,N_6755);
nand U9169 (N_9169,N_6610,N_6635);
or U9170 (N_9170,N_8732,N_8877);
or U9171 (N_9171,N_8140,N_8189);
and U9172 (N_9172,N_6789,N_6586);
or U9173 (N_9173,N_7342,N_6457);
or U9174 (N_9174,N_8070,N_8900);
nor U9175 (N_9175,N_8088,N_7634);
nand U9176 (N_9176,N_8604,N_6230);
nand U9177 (N_9177,N_8126,N_7748);
nand U9178 (N_9178,N_7617,N_6868);
nor U9179 (N_9179,N_7463,N_8827);
nand U9180 (N_9180,N_8059,N_8690);
nand U9181 (N_9181,N_7783,N_7900);
and U9182 (N_9182,N_7368,N_6944);
nand U9183 (N_9183,N_7413,N_6060);
and U9184 (N_9184,N_8054,N_7099);
and U9185 (N_9185,N_6089,N_6293);
and U9186 (N_9186,N_6521,N_8299);
or U9187 (N_9187,N_8955,N_6827);
and U9188 (N_9188,N_6481,N_7053);
or U9189 (N_9189,N_6073,N_8328);
nand U9190 (N_9190,N_8683,N_8819);
and U9191 (N_9191,N_7992,N_6168);
nor U9192 (N_9192,N_6996,N_8353);
nand U9193 (N_9193,N_8482,N_6325);
nand U9194 (N_9194,N_6276,N_6780);
nand U9195 (N_9195,N_6621,N_6618);
or U9196 (N_9196,N_7257,N_6811);
or U9197 (N_9197,N_6641,N_7418);
or U9198 (N_9198,N_8658,N_7440);
or U9199 (N_9199,N_7065,N_8641);
nor U9200 (N_9200,N_6969,N_7274);
nor U9201 (N_9201,N_6874,N_6410);
nand U9202 (N_9202,N_7263,N_6539);
nor U9203 (N_9203,N_7178,N_6844);
or U9204 (N_9204,N_8866,N_7001);
and U9205 (N_9205,N_8605,N_7825);
nor U9206 (N_9206,N_6973,N_6554);
or U9207 (N_9207,N_6578,N_7804);
nand U9208 (N_9208,N_7448,N_6664);
nand U9209 (N_9209,N_6906,N_8460);
nand U9210 (N_9210,N_8872,N_7300);
and U9211 (N_9211,N_8495,N_8917);
or U9212 (N_9212,N_7812,N_6526);
and U9213 (N_9213,N_8636,N_7105);
and U9214 (N_9214,N_6602,N_6383);
nand U9215 (N_9215,N_7072,N_6153);
and U9216 (N_9216,N_7074,N_7614);
or U9217 (N_9217,N_7339,N_6538);
xor U9218 (N_9218,N_7674,N_8254);
and U9219 (N_9219,N_8102,N_7068);
nand U9220 (N_9220,N_6674,N_7984);
and U9221 (N_9221,N_8113,N_7003);
nor U9222 (N_9222,N_8461,N_8138);
xnor U9223 (N_9223,N_8028,N_6957);
and U9224 (N_9224,N_8300,N_6359);
nor U9225 (N_9225,N_7311,N_6639);
xor U9226 (N_9226,N_6144,N_7530);
nand U9227 (N_9227,N_8893,N_7140);
nor U9228 (N_9228,N_8847,N_7722);
or U9229 (N_9229,N_8338,N_7453);
nand U9230 (N_9230,N_8185,N_6880);
or U9231 (N_9231,N_6051,N_8842);
and U9232 (N_9232,N_8215,N_6772);
and U9233 (N_9233,N_7282,N_6090);
nor U9234 (N_9234,N_7382,N_7505);
nor U9235 (N_9235,N_6260,N_7426);
nand U9236 (N_9236,N_8628,N_7527);
nand U9237 (N_9237,N_6129,N_7159);
and U9238 (N_9238,N_6024,N_8419);
and U9239 (N_9239,N_7991,N_8654);
or U9240 (N_9240,N_7821,N_8038);
and U9241 (N_9241,N_8142,N_8524);
or U9242 (N_9242,N_6018,N_6791);
or U9243 (N_9243,N_6413,N_7276);
nand U9244 (N_9244,N_8513,N_6565);
nor U9245 (N_9245,N_8965,N_8078);
xnor U9246 (N_9246,N_8171,N_6786);
or U9247 (N_9247,N_8772,N_6715);
xor U9248 (N_9248,N_7791,N_6280);
xor U9249 (N_9249,N_6771,N_7671);
or U9250 (N_9250,N_8389,N_6670);
and U9251 (N_9251,N_6177,N_7264);
nor U9252 (N_9252,N_8640,N_8267);
or U9253 (N_9253,N_7132,N_7482);
nor U9254 (N_9254,N_6788,N_8368);
xnor U9255 (N_9255,N_6839,N_6311);
or U9256 (N_9256,N_7570,N_6160);
and U9257 (N_9257,N_6427,N_8183);
nor U9258 (N_9258,N_7919,N_7914);
xnor U9259 (N_9259,N_6430,N_6302);
or U9260 (N_9260,N_8938,N_8103);
and U9261 (N_9261,N_7938,N_7600);
nand U9262 (N_9262,N_6693,N_6506);
nand U9263 (N_9263,N_7025,N_8918);
and U9264 (N_9264,N_7203,N_8743);
or U9265 (N_9265,N_6749,N_7305);
or U9266 (N_9266,N_7678,N_6797);
and U9267 (N_9267,N_7785,N_8273);
nand U9268 (N_9268,N_8431,N_7888);
or U9269 (N_9269,N_8362,N_7348);
and U9270 (N_9270,N_8472,N_6834);
and U9271 (N_9271,N_6825,N_7330);
xnor U9272 (N_9272,N_7740,N_7582);
and U9273 (N_9273,N_7669,N_8599);
or U9274 (N_9274,N_7909,N_7755);
nand U9275 (N_9275,N_8321,N_7251);
nand U9276 (N_9276,N_8627,N_6631);
or U9277 (N_9277,N_6675,N_6897);
or U9278 (N_9278,N_8899,N_7492);
and U9279 (N_9279,N_8509,N_7365);
nand U9280 (N_9280,N_6142,N_8826);
nand U9281 (N_9281,N_7808,N_6013);
nand U9282 (N_9282,N_6139,N_8191);
and U9283 (N_9283,N_6332,N_7352);
or U9284 (N_9284,N_6542,N_6807);
and U9285 (N_9285,N_7762,N_6301);
or U9286 (N_9286,N_8391,N_7138);
nor U9287 (N_9287,N_6465,N_8530);
nand U9288 (N_9288,N_6649,N_8318);
nand U9289 (N_9289,N_7583,N_6154);
nand U9290 (N_9290,N_7700,N_7447);
nor U9291 (N_9291,N_6213,N_7345);
and U9292 (N_9292,N_8905,N_7344);
nand U9293 (N_9293,N_8061,N_6132);
or U9294 (N_9294,N_6545,N_7692);
xor U9295 (N_9295,N_8445,N_8475);
or U9296 (N_9296,N_7799,N_7457);
or U9297 (N_9297,N_8990,N_7014);
nand U9298 (N_9298,N_8216,N_7660);
nand U9299 (N_9299,N_7571,N_8558);
nand U9300 (N_9300,N_7632,N_7797);
nor U9301 (N_9301,N_8305,N_7040);
and U9302 (N_9302,N_7717,N_7685);
or U9303 (N_9303,N_8740,N_8993);
nor U9304 (N_9304,N_6767,N_8768);
nor U9305 (N_9305,N_8960,N_7573);
or U9306 (N_9306,N_7228,N_7008);
nor U9307 (N_9307,N_6587,N_7699);
and U9308 (N_9308,N_6981,N_8776);
or U9309 (N_9309,N_8895,N_6560);
nor U9310 (N_9310,N_6754,N_6779);
and U9311 (N_9311,N_7175,N_8700);
nor U9312 (N_9312,N_8571,N_7446);
nor U9313 (N_9313,N_8210,N_6556);
or U9314 (N_9314,N_8994,N_8241);
nand U9315 (N_9315,N_8117,N_7884);
nand U9316 (N_9316,N_7240,N_6067);
nor U9317 (N_9317,N_7630,N_6209);
and U9318 (N_9318,N_7542,N_7800);
nor U9319 (N_9319,N_8053,N_6845);
xor U9320 (N_9320,N_7256,N_8972);
and U9321 (N_9321,N_8565,N_8498);
nor U9322 (N_9322,N_7107,N_6616);
nand U9323 (N_9323,N_7517,N_8718);
and U9324 (N_9324,N_7045,N_8479);
and U9325 (N_9325,N_7377,N_8111);
xnor U9326 (N_9326,N_6573,N_6040);
or U9327 (N_9327,N_8522,N_8001);
and U9328 (N_9328,N_8345,N_8792);
and U9329 (N_9329,N_7046,N_6781);
xor U9330 (N_9330,N_7949,N_8165);
or U9331 (N_9331,N_7122,N_7955);
xnor U9332 (N_9332,N_8949,N_6030);
nor U9333 (N_9333,N_8464,N_6580);
nor U9334 (N_9334,N_7716,N_7450);
and U9335 (N_9335,N_7395,N_8094);
and U9336 (N_9336,N_7292,N_6255);
nor U9337 (N_9337,N_7320,N_8741);
or U9338 (N_9338,N_6235,N_8335);
or U9339 (N_9339,N_7473,N_8228);
nor U9340 (N_9340,N_7719,N_8065);
and U9341 (N_9341,N_7754,N_8594);
and U9342 (N_9342,N_8192,N_6862);
or U9343 (N_9343,N_8499,N_7681);
nand U9344 (N_9344,N_8815,N_7479);
nor U9345 (N_9345,N_8286,N_7895);
and U9346 (N_9346,N_7567,N_8010);
nand U9347 (N_9347,N_6047,N_7597);
or U9348 (N_9348,N_8726,N_6515);
xor U9349 (N_9349,N_6307,N_8717);
nand U9350 (N_9350,N_8797,N_7255);
and U9351 (N_9351,N_7288,N_8450);
xnor U9352 (N_9352,N_8760,N_8429);
nor U9353 (N_9353,N_6707,N_6180);
or U9354 (N_9354,N_6713,N_7221);
or U9355 (N_9355,N_8962,N_7430);
or U9356 (N_9356,N_8119,N_8774);
nor U9357 (N_9357,N_8333,N_7967);
nor U9358 (N_9358,N_7772,N_7598);
and U9359 (N_9359,N_8055,N_6133);
or U9360 (N_9360,N_8226,N_7932);
and U9361 (N_9361,N_7789,N_7390);
or U9362 (N_9362,N_7781,N_6724);
nand U9363 (N_9363,N_7087,N_8468);
xnor U9364 (N_9364,N_8178,N_6677);
xnor U9365 (N_9365,N_8014,N_8643);
nand U9366 (N_9366,N_8426,N_7215);
xor U9367 (N_9367,N_6364,N_6581);
and U9368 (N_9368,N_8786,N_6250);
xnor U9369 (N_9369,N_6229,N_8330);
nor U9370 (N_9370,N_7085,N_8301);
or U9371 (N_9371,N_7403,N_6290);
or U9372 (N_9372,N_7849,N_7015);
and U9373 (N_9373,N_6872,N_6278);
nor U9374 (N_9374,N_6842,N_6365);
nor U9375 (N_9375,N_6982,N_7623);
or U9376 (N_9376,N_7337,N_7468);
nor U9377 (N_9377,N_7855,N_6798);
xor U9378 (N_9378,N_6126,N_6527);
or U9379 (N_9379,N_8294,N_8159);
nand U9380 (N_9380,N_7398,N_6533);
nor U9381 (N_9381,N_8436,N_7911);
nor U9382 (N_9382,N_8810,N_8123);
or U9383 (N_9383,N_7928,N_8146);
or U9384 (N_9384,N_6294,N_7050);
xor U9385 (N_9385,N_8818,N_8707);
or U9386 (N_9386,N_7874,N_6026);
nand U9387 (N_9387,N_8455,N_8572);
and U9388 (N_9388,N_7205,N_6721);
nor U9389 (N_9389,N_6226,N_8985);
or U9390 (N_9390,N_8315,N_7007);
nand U9391 (N_9391,N_6784,N_6672);
and U9392 (N_9392,N_8618,N_8162);
or U9393 (N_9393,N_8730,N_7679);
nor U9394 (N_9394,N_7411,N_8910);
or U9395 (N_9395,N_7047,N_7476);
nand U9396 (N_9396,N_7868,N_6628);
nor U9397 (N_9397,N_8856,N_6599);
and U9398 (N_9398,N_8981,N_8617);
nand U9399 (N_9399,N_7250,N_7284);
or U9400 (N_9400,N_7193,N_6007);
and U9401 (N_9401,N_8526,N_8002);
and U9402 (N_9402,N_7904,N_8409);
nor U9403 (N_9403,N_6274,N_6196);
nor U9404 (N_9404,N_8638,N_6912);
nor U9405 (N_9405,N_6021,N_6225);
xor U9406 (N_9406,N_8339,N_7017);
nor U9407 (N_9407,N_7013,N_7226);
nor U9408 (N_9408,N_8812,N_6927);
nor U9409 (N_9409,N_8457,N_6951);
or U9410 (N_9410,N_6738,N_6039);
or U9411 (N_9411,N_7497,N_7139);
xor U9412 (N_9412,N_8068,N_7081);
or U9413 (N_9413,N_8104,N_7507);
nor U9414 (N_9414,N_7810,N_7705);
nand U9415 (N_9415,N_7668,N_8578);
nand U9416 (N_9416,N_7645,N_8430);
nor U9417 (N_9417,N_6472,N_6009);
nand U9418 (N_9418,N_6873,N_7478);
nor U9419 (N_9419,N_8947,N_8153);
or U9420 (N_9420,N_6660,N_6312);
nor U9421 (N_9421,N_7295,N_7142);
nand U9422 (N_9422,N_6076,N_6661);
and U9423 (N_9423,N_6134,N_7982);
and U9424 (N_9424,N_6687,N_8682);
xor U9425 (N_9425,N_7596,N_8753);
nor U9426 (N_9426,N_6368,N_6183);
or U9427 (N_9427,N_8322,N_8201);
or U9428 (N_9428,N_7826,N_8934);
nand U9429 (N_9429,N_7231,N_8595);
and U9430 (N_9430,N_6867,N_6805);
nor U9431 (N_9431,N_7229,N_7715);
nand U9432 (N_9432,N_6646,N_7218);
and U9433 (N_9433,N_6654,N_8514);
nor U9434 (N_9434,N_7946,N_8708);
nand U9435 (N_9435,N_7100,N_6002);
and U9436 (N_9436,N_6450,N_8729);
xor U9437 (N_9437,N_8257,N_6469);
nor U9438 (N_9438,N_7879,N_7920);
nor U9439 (N_9439,N_7179,N_7802);
nor U9440 (N_9440,N_8375,N_8894);
and U9441 (N_9441,N_6314,N_7877);
and U9442 (N_9442,N_7702,N_6501);
nor U9443 (N_9443,N_8706,N_8395);
and U9444 (N_9444,N_7279,N_7861);
nor U9445 (N_9445,N_7011,N_7381);
and U9446 (N_9446,N_6367,N_7243);
nor U9447 (N_9447,N_8624,N_8897);
nand U9448 (N_9448,N_7406,N_8306);
or U9449 (N_9449,N_6928,N_6095);
nand U9450 (N_9450,N_8451,N_6017);
nand U9451 (N_9451,N_7371,N_6052);
or U9452 (N_9452,N_7303,N_8343);
xor U9453 (N_9453,N_7067,N_8453);
nor U9454 (N_9454,N_7157,N_7156);
nand U9455 (N_9455,N_7659,N_8838);
and U9456 (N_9456,N_8570,N_7767);
or U9457 (N_9457,N_6281,N_8280);
or U9458 (N_9458,N_8648,N_8549);
nor U9459 (N_9459,N_7499,N_7872);
or U9460 (N_9460,N_8837,N_8891);
and U9461 (N_9461,N_6182,N_8406);
nand U9462 (N_9462,N_8828,N_6178);
xor U9463 (N_9463,N_8211,N_7780);
and U9464 (N_9464,N_6933,N_6461);
nor U9465 (N_9465,N_8434,N_8881);
or U9466 (N_9466,N_7027,N_7325);
or U9467 (N_9467,N_8408,N_7431);
or U9468 (N_9468,N_6696,N_6423);
xor U9469 (N_9469,N_8067,N_8466);
and U9470 (N_9470,N_6138,N_7123);
or U9471 (N_9471,N_8912,N_7220);
and U9472 (N_9472,N_8268,N_6776);
and U9473 (N_9473,N_6171,N_7362);
nor U9474 (N_9474,N_8456,N_6513);
or U9475 (N_9475,N_7464,N_6351);
or U9476 (N_9476,N_6861,N_8660);
nand U9477 (N_9477,N_6227,N_8417);
xor U9478 (N_9478,N_6316,N_8504);
nor U9479 (N_9479,N_6219,N_8120);
or U9480 (N_9480,N_8546,N_7601);
xor U9481 (N_9481,N_6519,N_8331);
xor U9482 (N_9482,N_8295,N_6100);
xnor U9483 (N_9483,N_7210,N_8166);
and U9484 (N_9484,N_8204,N_6381);
nand U9485 (N_9485,N_6847,N_7846);
nand U9486 (N_9486,N_8223,N_6233);
and U9487 (N_9487,N_8081,N_6016);
nor U9488 (N_9488,N_7061,N_7836);
nand U9489 (N_9489,N_6486,N_8720);
or U9490 (N_9490,N_7648,N_6773);
nor U9491 (N_9491,N_8405,N_6606);
and U9492 (N_9492,N_6348,N_7397);
nor U9493 (N_9493,N_6596,N_7432);
or U9494 (N_9494,N_6184,N_8903);
nor U9495 (N_9495,N_6733,N_8415);
nor U9496 (N_9496,N_6543,N_6470);
or U9497 (N_9497,N_8224,N_7707);
nor U9498 (N_9498,N_6447,N_8243);
xnor U9499 (N_9499,N_7945,N_8016);
nand U9500 (N_9500,N_8959,N_6889);
or U9501 (N_9501,N_8801,N_6387);
nand U9502 (N_9502,N_8520,N_6701);
xor U9503 (N_9503,N_7091,N_7615);
or U9504 (N_9504,N_8625,N_8251);
nand U9505 (N_9505,N_6393,N_6605);
nor U9506 (N_9506,N_8264,N_7181);
nor U9507 (N_9507,N_8359,N_6262);
and U9508 (N_9508,N_6541,N_7894);
or U9509 (N_9509,N_6795,N_7576);
or U9510 (N_9510,N_7064,N_8478);
or U9511 (N_9511,N_6830,N_6165);
nor U9512 (N_9512,N_8252,N_6420);
nor U9513 (N_9513,N_8502,N_8781);
xnor U9514 (N_9514,N_8788,N_6967);
nor U9515 (N_9515,N_8134,N_8921);
or U9516 (N_9516,N_6119,N_8785);
nor U9517 (N_9517,N_8033,N_6850);
nand U9518 (N_9518,N_7927,N_8587);
and U9519 (N_9519,N_6238,N_6291);
or U9520 (N_9520,N_6703,N_7837);
xor U9521 (N_9521,N_7298,N_6597);
nand U9522 (N_9522,N_7486,N_6918);
nor U9523 (N_9523,N_8686,N_6729);
nand U9524 (N_9524,N_8176,N_8662);
or U9525 (N_9525,N_8106,N_8566);
xor U9526 (N_9526,N_7321,N_6576);
nor U9527 (N_9527,N_8663,N_6753);
or U9528 (N_9528,N_6419,N_6114);
or U9529 (N_9529,N_6934,N_7805);
or U9530 (N_9530,N_8369,N_6188);
or U9531 (N_9531,N_6719,N_7934);
and U9532 (N_9532,N_8020,N_7388);
nand U9533 (N_9533,N_7990,N_8425);
nor U9534 (N_9534,N_6609,N_7422);
nand U9535 (N_9535,N_6892,N_6131);
xor U9536 (N_9536,N_8401,N_7962);
or U9537 (N_9537,N_8883,N_7631);
xnor U9538 (N_9538,N_6181,N_8168);
nand U9539 (N_9539,N_7815,N_7541);
xor U9540 (N_9540,N_7128,N_6108);
or U9541 (N_9541,N_8194,N_7380);
nor U9542 (N_9542,N_8379,N_7524);
and U9543 (N_9543,N_7196,N_7151);
nor U9544 (N_9544,N_6484,N_8590);
or U9545 (N_9545,N_6710,N_8681);
and U9546 (N_9546,N_8535,N_8376);
nor U9547 (N_9547,N_8446,N_6520);
or U9548 (N_9548,N_7558,N_8977);
nor U9549 (N_9549,N_8458,N_8657);
xor U9550 (N_9550,N_6000,N_7343);
and U9551 (N_9551,N_8018,N_8050);
nand U9552 (N_9552,N_6483,N_8370);
nor U9553 (N_9553,N_6816,N_6487);
or U9554 (N_9554,N_6416,N_7523);
xnor U9555 (N_9555,N_6062,N_7049);
and U9556 (N_9556,N_8927,N_7933);
or U9557 (N_9557,N_8854,N_8680);
or U9558 (N_9558,N_8563,N_7317);
xnor U9559 (N_9559,N_7034,N_7723);
nor U9560 (N_9560,N_7625,N_7273);
or U9561 (N_9561,N_7646,N_8481);
or U9562 (N_9562,N_8586,N_6723);
and U9563 (N_9563,N_6726,N_8501);
and U9564 (N_9564,N_8323,N_7009);
nand U9565 (N_9565,N_7190,N_6157);
nor U9566 (N_9566,N_7520,N_6187);
or U9567 (N_9567,N_7794,N_8787);
xnor U9568 (N_9568,N_6801,N_8885);
and U9569 (N_9569,N_8500,N_8941);
and U9570 (N_9570,N_7587,N_8886);
or U9571 (N_9571,N_8676,N_7807);
or U9572 (N_9572,N_7456,N_7749);
and U9573 (N_9573,N_7313,N_7490);
and U9574 (N_9574,N_7018,N_6571);
nand U9575 (N_9575,N_7436,N_7732);
nor U9576 (N_9576,N_8992,N_8579);
and U9577 (N_9577,N_6127,N_7761);
or U9578 (N_9578,N_6048,N_7160);
and U9579 (N_9579,N_8646,N_7795);
or U9580 (N_9580,N_7816,N_7667);
nand U9581 (N_9581,N_6976,N_8645);
nand U9582 (N_9582,N_8898,N_8329);
or U9583 (N_9583,N_6075,N_6684);
and U9584 (N_9584,N_6764,N_8996);
nand U9585 (N_9585,N_8077,N_7247);
or U9586 (N_9586,N_7232,N_8821);
nand U9587 (N_9587,N_8341,N_8552);
and U9588 (N_9588,N_8281,N_6446);
or U9589 (N_9589,N_8462,N_7219);
or U9590 (N_9590,N_8585,N_7471);
nor U9591 (N_9591,N_8048,N_7333);
and U9592 (N_9592,N_7714,N_7032);
nor U9593 (N_9593,N_8203,N_7083);
or U9594 (N_9594,N_6103,N_6929);
nor U9595 (N_9595,N_6570,N_8354);
xor U9596 (N_9596,N_7921,N_6421);
xnor U9597 (N_9597,N_6653,N_8161);
xnor U9598 (N_9598,N_8152,N_8151);
and U9599 (N_9599,N_8248,N_7369);
or U9600 (N_9600,N_7580,N_6167);
nand U9601 (N_9601,N_6846,N_8626);
or U9602 (N_9602,N_7848,N_7206);
or U9603 (N_9603,N_7924,N_7270);
and U9604 (N_9604,N_8913,N_6231);
or U9605 (N_9605,N_6949,N_6819);
nand U9606 (N_9606,N_8080,N_7359);
nand U9607 (N_9607,N_8410,N_8693);
and U9608 (N_9608,N_6297,N_7400);
nand U9609 (N_9609,N_7314,N_7086);
and U9610 (N_9610,N_7496,N_6191);
and U9611 (N_9611,N_7312,N_6436);
and U9612 (N_9612,N_8397,N_7420);
and U9613 (N_9613,N_6681,N_8017);
or U9614 (N_9614,N_6741,N_7860);
or U9615 (N_9615,N_8197,N_6594);
nor U9616 (N_9616,N_8569,N_6877);
nand U9617 (N_9617,N_8998,N_8619);
or U9618 (N_9618,N_7026,N_7494);
and U9619 (N_9619,N_8364,N_7189);
or U9620 (N_9620,N_7806,N_6775);
or U9621 (N_9621,N_8936,N_6595);
nor U9622 (N_9622,N_6569,N_6623);
nor U9623 (N_9623,N_8260,N_6201);
nand U9624 (N_9624,N_6613,N_6611);
or U9625 (N_9625,N_8283,N_6377);
or U9626 (N_9626,N_7787,N_8611);
nor U9627 (N_9627,N_6237,N_7969);
and U9628 (N_9628,N_7720,N_8057);
or U9629 (N_9629,N_6329,N_6901);
and U9630 (N_9630,N_8661,N_6149);
nor U9631 (N_9631,N_7726,N_7966);
or U9632 (N_9632,N_8463,N_7563);
and U9633 (N_9633,N_6498,N_7833);
nor U9634 (N_9634,N_8266,N_6592);
and U9635 (N_9635,N_6882,N_7711);
xnor U9636 (N_9636,N_6783,N_8534);
xnor U9637 (N_9637,N_6964,N_6306);
xnor U9638 (N_9638,N_8629,N_8544);
nand U9639 (N_9639,N_7111,N_7417);
and U9640 (N_9640,N_7734,N_8022);
nand U9641 (N_9641,N_7235,N_6966);
nand U9642 (N_9642,N_7438,N_8710);
nor U9643 (N_9643,N_8794,N_8607);
nor U9644 (N_9644,N_6477,N_8314);
and U9645 (N_9645,N_8620,N_8857);
and U9646 (N_9646,N_8336,N_8521);
or U9647 (N_9647,N_7980,N_6829);
xnor U9648 (N_9648,N_7759,N_6162);
nand U9649 (N_9649,N_8973,N_6583);
nand U9650 (N_9650,N_6198,N_6370);
or U9651 (N_9651,N_7427,N_7410);
nor U9652 (N_9652,N_7603,N_7859);
nand U9653 (N_9653,N_6840,N_7082);
nor U9654 (N_9654,N_8089,N_7452);
nand U9655 (N_9655,N_8659,N_7124);
and U9656 (N_9656,N_6769,N_8476);
and U9657 (N_9657,N_7134,N_7666);
or U9658 (N_9658,N_6955,N_6268);
and U9659 (N_9659,N_7637,N_6025);
xnor U9660 (N_9660,N_6871,N_6020);
and U9661 (N_9661,N_7442,N_8000);
or U9662 (N_9662,N_8909,N_7271);
or U9663 (N_9663,N_6197,N_6272);
xor U9664 (N_9664,N_6082,N_7186);
and U9665 (N_9665,N_7737,N_6989);
nor U9666 (N_9666,N_7483,N_7518);
or U9667 (N_9667,N_7237,N_7819);
and U9668 (N_9668,N_6042,N_6505);
nand U9669 (N_9669,N_6078,N_6118);
xnor U9670 (N_9670,N_7244,N_8623);
or U9671 (N_9671,N_7607,N_8056);
nand U9672 (N_9672,N_8288,N_6682);
xor U9673 (N_9673,N_6507,N_6292);
and U9674 (N_9674,N_8865,N_6210);
nand U9675 (N_9675,N_8489,N_7878);
nor U9676 (N_9676,N_7550,N_6993);
and U9677 (N_9677,N_7488,N_7197);
nor U9678 (N_9678,N_7504,N_8465);
nor U9679 (N_9679,N_7760,N_7224);
nand U9680 (N_9680,N_7907,N_7172);
nand U9681 (N_9681,N_7168,N_8853);
or U9682 (N_9682,N_7419,N_7260);
nor U9683 (N_9683,N_6983,N_6659);
and U9684 (N_9684,N_7324,N_6222);
and U9685 (N_9685,N_8596,N_7449);
nand U9686 (N_9686,N_8360,N_6402);
nor U9687 (N_9687,N_6603,N_6362);
or U9688 (N_9688,N_7592,N_8219);
and U9689 (N_9689,N_6689,N_6471);
nor U9690 (N_9690,N_6211,N_8447);
or U9691 (N_9691,N_7624,N_7042);
or U9692 (N_9692,N_7242,N_7952);
or U9693 (N_9693,N_8779,N_6985);
nand U9694 (N_9694,N_8235,N_6189);
or U9695 (N_9695,N_8492,N_7917);
and U9696 (N_9696,N_6953,N_7656);
nand U9697 (N_9697,N_7703,N_6517);
nand U9698 (N_9698,N_6221,N_6705);
xor U9699 (N_9699,N_6761,N_7522);
nor U9700 (N_9700,N_8177,N_7283);
nor U9701 (N_9701,N_8817,N_6917);
nor U9702 (N_9702,N_7346,N_7318);
or U9703 (N_9703,N_8754,N_8180);
and U9704 (N_9704,N_6987,N_6342);
nand U9705 (N_9705,N_6650,N_8906);
and U9706 (N_9706,N_6806,N_8023);
nor U9707 (N_9707,N_6932,N_6058);
nand U9708 (N_9708,N_8541,N_7840);
nand U9709 (N_9709,N_8403,N_7249);
and U9710 (N_9710,N_8796,N_8043);
nor U9711 (N_9711,N_6105,N_6503);
nand U9712 (N_9712,N_8806,N_6939);
and U9713 (N_9713,N_6680,N_6568);
nor U9714 (N_9714,N_6008,N_7756);
or U9715 (N_9715,N_8508,N_7408);
nand U9716 (N_9716,N_7310,N_8297);
or U9717 (N_9717,N_8349,N_6145);
or U9718 (N_9718,N_6056,N_8931);
or U9719 (N_9719,N_6220,N_7416);
and U9720 (N_9720,N_6914,N_6950);
or U9721 (N_9721,N_7141,N_8125);
nand U9722 (N_9722,N_8769,N_8046);
xnor U9723 (N_9723,N_6137,N_6435);
xor U9724 (N_9724,N_7863,N_6730);
or U9725 (N_9725,N_8452,N_8422);
and U9726 (N_9726,N_6731,N_8948);
or U9727 (N_9727,N_6375,N_8577);
nor U9728 (N_9728,N_6656,N_7602);
or U9729 (N_9729,N_6284,N_6334);
nand U9730 (N_9730,N_8275,N_7254);
and U9731 (N_9731,N_8483,N_7443);
or U9732 (N_9732,N_7429,N_7004);
or U9733 (N_9733,N_6619,N_8831);
and U9734 (N_9734,N_6169,N_8597);
or U9735 (N_9735,N_8935,N_6121);
nand U9736 (N_9736,N_6875,N_8848);
xnor U9737 (N_9737,N_7336,N_8845);
or U9738 (N_9738,N_8039,N_6147);
and U9739 (N_9739,N_8008,N_8214);
nor U9740 (N_9740,N_6647,N_8363);
or U9741 (N_9741,N_7185,N_8908);
or U9742 (N_9742,N_8540,N_8007);
or U9743 (N_9743,N_6848,N_7338);
or U9744 (N_9744,N_7639,N_6101);
or U9745 (N_9745,N_7999,N_6324);
or U9746 (N_9746,N_7052,N_6808);
or U9747 (N_9747,N_6512,N_8258);
nor U9748 (N_9748,N_7994,N_8383);
or U9749 (N_9749,N_6589,N_7012);
or U9750 (N_9750,N_6414,N_8380);
or U9751 (N_9751,N_6243,N_6557);
xor U9752 (N_9752,N_7204,N_7947);
or U9753 (N_9753,N_7745,N_8188);
xnor U9754 (N_9754,N_6321,N_6727);
xor U9755 (N_9755,N_8807,N_8207);
nand U9756 (N_9756,N_6155,N_8734);
and U9757 (N_9757,N_8816,N_7769);
nand U9758 (N_9758,N_7248,N_7554);
or U9759 (N_9759,N_6548,N_7509);
nor U9760 (N_9760,N_6179,N_6686);
or U9761 (N_9761,N_6550,N_6117);
nor U9762 (N_9762,N_8702,N_6045);
nor U9763 (N_9763,N_6124,N_8911);
or U9764 (N_9764,N_7981,N_7491);
or U9765 (N_9765,N_8737,N_7404);
nor U9766 (N_9766,N_8344,N_7744);
or U9767 (N_9767,N_6979,N_6028);
nand U9768 (N_9768,N_7078,N_7590);
and U9769 (N_9769,N_7117,N_8198);
nor U9770 (N_9770,N_7356,N_6335);
nor U9771 (N_9771,N_8820,N_7977);
nor U9772 (N_9772,N_8366,N_7658);
or U9773 (N_9773,N_7227,N_8603);
nor U9774 (N_9774,N_7709,N_7423);
nand U9775 (N_9775,N_6217,N_8775);
nand U9776 (N_9776,N_6970,N_6037);
nand U9777 (N_9777,N_8440,N_8650);
nand U9778 (N_9778,N_7472,N_8713);
or U9779 (N_9779,N_6720,N_8863);
or U9780 (N_9780,N_8983,N_8644);
nand U9781 (N_9781,N_8488,N_7299);
xnor U9782 (N_9782,N_7682,N_7041);
nand U9783 (N_9783,N_7641,N_8511);
nand U9784 (N_9784,N_6261,N_6669);
nor U9785 (N_9785,N_7057,N_6391);
nand U9786 (N_9786,N_7536,N_8668);
or U9787 (N_9787,N_8218,N_8631);
nand U9788 (N_9788,N_8532,N_8888);
nand U9789 (N_9789,N_7858,N_6440);
xor U9790 (N_9790,N_8637,N_7818);
nor U9791 (N_9791,N_6817,N_6622);
nor U9792 (N_9792,N_7513,N_6327);
and U9793 (N_9793,N_8545,N_8527);
or U9794 (N_9794,N_6968,N_7835);
nor U9795 (N_9795,N_7670,N_7407);
nand U9796 (N_9796,N_7421,N_8833);
and U9797 (N_9797,N_6485,N_6883);
or U9798 (N_9798,N_7652,N_7853);
or U9799 (N_9799,N_6838,N_6482);
nand U9800 (N_9800,N_8255,N_7944);
nor U9801 (N_9801,N_7323,N_7512);
nand U9802 (N_9802,N_6965,N_7043);
and U9803 (N_9803,N_8232,N_8503);
nor U9804 (N_9804,N_7876,N_8355);
and U9805 (N_9805,N_8688,N_8227);
or U9806 (N_9806,N_7830,N_8844);
xor U9807 (N_9807,N_7158,N_6566);
or U9808 (N_9808,N_7475,N_7379);
or U9809 (N_9809,N_8536,N_8108);
and U9810 (N_9810,N_7136,N_6591);
xor U9811 (N_9811,N_6338,N_8158);
nor U9812 (N_9812,N_8427,N_8841);
xnor U9813 (N_9813,N_6748,N_8167);
nor U9814 (N_9814,N_8099,N_7718);
or U9815 (N_9815,N_6309,N_7561);
xor U9816 (N_9816,N_6163,N_6185);
nand U9817 (N_9817,N_6555,N_7170);
and U9818 (N_9818,N_6607,N_6094);
nand U9819 (N_9819,N_8282,N_6464);
nor U9820 (N_9820,N_8202,N_7922);
nand U9821 (N_9821,N_7958,N_7687);
nand U9822 (N_9822,N_7076,N_8035);
nor U9823 (N_9823,N_6940,N_8957);
or U9824 (N_9824,N_8238,N_6186);
or U9825 (N_9825,N_6615,N_7104);
or U9826 (N_9826,N_8222,N_6841);
nor U9827 (N_9827,N_6258,N_8087);
and U9828 (N_9828,N_6223,N_6022);
and U9829 (N_9829,N_6765,N_6629);
and U9830 (N_9830,N_6404,N_6954);
or U9831 (N_9831,N_7540,N_7101);
xor U9832 (N_9832,N_6510,N_8829);
nand U9833 (N_9833,N_8952,N_7202);
or U9834 (N_9834,N_8428,N_8261);
nor U9835 (N_9835,N_7112,N_8205);
xnor U9836 (N_9836,N_8832,N_7016);
nor U9837 (N_9837,N_8259,N_7655);
or U9838 (N_9838,N_7943,N_8652);
nand U9839 (N_9839,N_7803,N_8790);
xnor U9840 (N_9840,N_6159,N_8346);
or U9841 (N_9841,N_6433,N_8154);
nor U9842 (N_9842,N_8843,N_7764);
nor U9843 (N_9843,N_6299,N_8813);
xnor U9844 (N_9844,N_6374,N_6575);
and U9845 (N_9845,N_8220,N_6128);
nand U9846 (N_9846,N_8086,N_7935);
nor U9847 (N_9847,N_8855,N_7233);
nor U9848 (N_9848,N_8149,N_7080);
nand U9849 (N_9849,N_6991,N_7383);
nand U9850 (N_9850,N_6350,N_6640);
nand U9851 (N_9851,N_7163,N_7890);
and U9852 (N_9852,N_7126,N_8616);
and U9853 (N_9853,N_7108,N_8562);
and U9854 (N_9854,N_7278,N_6270);
and U9855 (N_9855,N_6612,N_8019);
nand U9856 (N_9856,N_6012,N_6561);
or U9857 (N_9857,N_6034,N_8042);
and U9858 (N_9858,N_7686,N_7538);
nand U9859 (N_9859,N_8182,N_8671);
nand U9860 (N_9860,N_7396,N_7972);
nor U9861 (N_9861,N_7566,N_8115);
xor U9862 (N_9862,N_8699,N_8961);
or U9863 (N_9863,N_7374,N_7241);
and U9864 (N_9864,N_6971,N_7963);
xnor U9865 (N_9865,N_7951,N_7184);
or U9866 (N_9866,N_7696,N_7852);
nand U9867 (N_9867,N_7930,N_6437);
nand U9868 (N_9868,N_7578,N_8064);
nor U9869 (N_9869,N_6763,N_7883);
nor U9870 (N_9870,N_8105,N_7618);
nand U9871 (N_9871,N_7079,N_7291);
nand U9872 (N_9872,N_6980,N_6886);
and U9873 (N_9873,N_7636,N_7073);
nand U9874 (N_9874,N_8083,N_8606);
nand U9875 (N_9875,N_7741,N_8387);
and U9876 (N_9876,N_8764,N_6921);
or U9877 (N_9877,N_8340,N_6087);
or U9878 (N_9878,N_7265,N_6035);
nor U9879 (N_9879,N_6700,N_7150);
xor U9880 (N_9880,N_6915,N_6909);
or U9881 (N_9881,N_7824,N_8568);
nand U9882 (N_9882,N_7941,N_6624);
and U9883 (N_9883,N_7370,N_8875);
or U9884 (N_9884,N_6053,N_6069);
and U9885 (N_9885,N_7146,N_8348);
and U9886 (N_9886,N_7508,N_6813);
nand U9887 (N_9887,N_8139,N_6106);
xnor U9888 (N_9888,N_7326,N_8750);
nor U9889 (N_9889,N_8925,N_8696);
nor U9890 (N_9890,N_6843,N_6382);
and U9891 (N_9891,N_7985,N_8424);
and U9892 (N_9892,N_6176,N_8759);
and U9893 (N_9893,N_7610,N_8263);
nand U9894 (N_9894,N_7102,N_6320);
or U9895 (N_9895,N_6232,N_8878);
and U9896 (N_9896,N_6636,N_8011);
nand U9897 (N_9897,N_8292,N_6409);
nor U9898 (N_9898,N_7664,N_7820);
nor U9899 (N_9899,N_8916,N_7832);
and U9900 (N_9900,N_7873,N_8200);
nand U9901 (N_9901,N_6212,N_8311);
or U9902 (N_9902,N_6036,N_8385);
nand U9903 (N_9903,N_7912,N_8722);
and U9904 (N_9904,N_7177,N_6064);
nand U9905 (N_9905,N_7090,N_6289);
or U9906 (N_9906,N_8474,N_7739);
and U9907 (N_9907,N_6102,N_8800);
nand U9908 (N_9908,N_8958,N_6952);
and U9909 (N_9909,N_8071,N_8851);
and U9910 (N_9910,N_6098,N_8901);
and U9911 (N_9911,N_7187,N_7062);
nand U9912 (N_9912,N_8861,N_6931);
nand U9913 (N_9913,N_7495,N_8999);
and U9914 (N_9914,N_8547,N_8485);
nand U9915 (N_9915,N_6228,N_6899);
nor U9916 (N_9916,N_7267,N_7964);
nor U9917 (N_9917,N_8186,N_8963);
or U9918 (N_9918,N_6537,N_7746);
or U9919 (N_9919,N_8156,N_7731);
and U9920 (N_9920,N_8516,N_6919);
nor U9921 (N_9921,N_8029,N_6319);
and U9922 (N_9922,N_6234,N_7394);
and U9923 (N_9923,N_8763,N_7208);
nand U9924 (N_9924,N_7127,N_8742);
nor U9925 (N_9925,N_7650,N_6444);
nand U9926 (N_9926,N_8614,N_7093);
or U9927 (N_9927,N_6714,N_8172);
nand U9928 (N_9928,N_8757,N_8229);
nor U9929 (N_9929,N_6263,N_7474);
or U9930 (N_9930,N_6885,N_7680);
nand U9931 (N_9931,N_7643,N_6945);
nor U9932 (N_9932,N_8213,N_8490);
and U9933 (N_9933,N_7954,N_6079);
or U9934 (N_9934,N_6642,N_7531);
or U9935 (N_9935,N_6014,N_8868);
nand U9936 (N_9936,N_8272,N_6080);
nand U9937 (N_9937,N_6790,N_8756);
nand U9938 (N_9938,N_8798,N_7552);
xnor U9939 (N_9939,N_6960,N_6910);
nor U9940 (N_9940,N_7546,N_7965);
nand U9941 (N_9941,N_7882,N_8358);
or U9942 (N_9942,N_7355,N_8978);
xnor U9943 (N_9943,N_7399,N_7621);
nor U9944 (N_9944,N_6448,N_7690);
and U9945 (N_9945,N_7850,N_8666);
nand U9946 (N_9946,N_8199,N_7871);
and U9947 (N_9947,N_7412,N_7077);
and U9948 (N_9948,N_8588,N_7281);
nand U9949 (N_9949,N_8746,N_7351);
nand U9950 (N_9950,N_7286,N_7828);
nor U9951 (N_9951,N_6913,N_6445);
nand U9952 (N_9952,N_6173,N_6494);
nand U9953 (N_9953,N_6405,N_6065);
nand U9954 (N_9954,N_7516,N_8956);
and U9955 (N_9955,N_8928,N_7051);
nand U9956 (N_9956,N_8473,N_8615);
nand U9957 (N_9957,N_7280,N_8850);
and U9958 (N_9958,N_7875,N_8075);
and U9959 (N_9959,N_6937,N_8761);
nand U9960 (N_9960,N_6799,N_6476);
or U9961 (N_9961,N_7441,N_6665);
and U9962 (N_9962,N_8433,N_7776);
nor U9963 (N_9963,N_6695,N_6911);
or U9964 (N_9964,N_8095,N_8384);
xor U9965 (N_9965,N_8555,N_7329);
nor U9966 (N_9966,N_8823,N_6716);
nor U9967 (N_9967,N_7236,N_7688);
nand U9968 (N_9968,N_8943,N_6865);
and U9969 (N_9969,N_7786,N_8846);
nand U9970 (N_9970,N_7387,N_8564);
or U9971 (N_9971,N_8157,N_7887);
xnor U9972 (N_9972,N_8225,N_8236);
or U9973 (N_9973,N_6963,N_7968);
xnor U9974 (N_9974,N_8725,N_6259);
nor U9975 (N_9975,N_8396,N_8487);
or U9976 (N_9976,N_8298,N_7989);
nand U9977 (N_9977,N_7584,N_7750);
and U9978 (N_9978,N_8470,N_6315);
or U9979 (N_9979,N_8003,N_7701);
or U9980 (N_9980,N_7096,N_8208);
or U9981 (N_9981,N_7036,N_7173);
and U9982 (N_9982,N_8361,N_6544);
xnor U9983 (N_9983,N_6704,N_7510);
xnor U9984 (N_9984,N_6643,N_6617);
or U9985 (N_9985,N_7620,N_8880);
nand U9986 (N_9986,N_8206,N_6658);
and U9987 (N_9987,N_6999,N_6567);
nand U9988 (N_9988,N_6086,N_6247);
nand U9989 (N_9989,N_7589,N_8735);
nand U9990 (N_9990,N_6739,N_6376);
nor U9991 (N_9991,N_6267,N_8976);
nand U9992 (N_9992,N_6531,N_7956);
and U9993 (N_9993,N_8193,N_7376);
and U9994 (N_9994,N_6562,N_6524);
or U9995 (N_9995,N_6236,N_7304);
or U9996 (N_9996,N_6904,N_7870);
nand U9997 (N_9997,N_8352,N_7809);
nor U9998 (N_9998,N_7845,N_8144);
nand U9999 (N_9999,N_8291,N_7544);
nor U10000 (N_10000,N_7428,N_8234);
and U10001 (N_10001,N_6692,N_8278);
and U10002 (N_10002,N_8130,N_8656);
nor U10003 (N_10003,N_7230,N_6762);
nand U10004 (N_10004,N_6454,N_8024);
nor U10005 (N_10005,N_6287,N_6802);
nand U10006 (N_10006,N_6195,N_7200);
nand U10007 (N_10007,N_7735,N_6459);
or U10008 (N_10008,N_8356,N_8533);
nor U10009 (N_10009,N_8642,N_6588);
nand U10010 (N_10010,N_6136,N_6863);
and U10011 (N_10011,N_7950,N_7023);
and U10012 (N_10012,N_7661,N_8155);
and U10013 (N_10013,N_7075,N_6054);
or U10014 (N_10014,N_7979,N_8542);
nand U10015 (N_10015,N_7331,N_7521);
nor U10016 (N_10016,N_6943,N_8673);
and U10017 (N_10017,N_7653,N_6271);
or U10018 (N_10018,N_6431,N_7217);
or U10019 (N_10019,N_7462,N_6441);
nor U10020 (N_10020,N_7252,N_6893);
nor U10021 (N_10021,N_7363,N_6331);
or U10022 (N_10022,N_8771,N_6836);
nand U10023 (N_10023,N_8937,N_6511);
nor U10024 (N_10024,N_7765,N_7758);
or U10025 (N_10025,N_6218,N_7366);
and U10026 (N_10026,N_6735,N_6734);
or U10027 (N_10027,N_8835,N_6768);
nor U10028 (N_10028,N_7915,N_6241);
and U10029 (N_10029,N_6528,N_7502);
and U10030 (N_10030,N_6462,N_7071);
and U10031 (N_10031,N_7889,N_6285);
nand U10032 (N_10032,N_8284,N_6254);
nor U10033 (N_10033,N_7425,N_6673);
or U10034 (N_10034,N_6662,N_8308);
or U10035 (N_10035,N_8304,N_8969);
nor U10036 (N_10036,N_7535,N_6941);
xnor U10037 (N_10037,N_8493,N_6884);
and U10038 (N_10038,N_7926,N_8932);
nor U10039 (N_10039,N_7216,N_7867);
nand U10040 (N_10040,N_8122,N_6685);
nand U10041 (N_10041,N_7253,N_7213);
nand U10042 (N_10042,N_7094,N_6516);
nor U10043 (N_10043,N_7195,N_8887);
and U10044 (N_10044,N_7606,N_8027);
xnor U10045 (N_10045,N_8143,N_7161);
and U10046 (N_10046,N_8041,N_7556);
or U10047 (N_10047,N_7869,N_6083);
nor U10048 (N_10048,N_6085,N_7959);
nand U10049 (N_10049,N_7044,N_6412);
and U10050 (N_10050,N_8443,N_8685);
nor U10051 (N_10051,N_6666,N_8684);
nand U10052 (N_10052,N_7925,N_7058);
or U10053 (N_10053,N_8031,N_8237);
nor U10054 (N_10054,N_6027,N_8030);
and U10055 (N_10055,N_7827,N_8859);
nor U10056 (N_10056,N_6489,N_8559);
xor U10057 (N_10057,N_6559,N_6866);
and U10058 (N_10058,N_8719,N_7916);
or U10059 (N_10059,N_7367,N_8712);
nor U10060 (N_10060,N_7595,N_7095);
nor U10061 (N_10061,N_6458,N_8494);
nand U10062 (N_10062,N_7116,N_7757);
or U10063 (N_10063,N_7306,N_7327);
nor U10064 (N_10064,N_8173,N_7378);
or U10065 (N_10065,N_6804,N_7155);
or U10066 (N_10066,N_6860,N_7358);
nor U10067 (N_10067,N_8449,N_7269);
xor U10068 (N_10068,N_6888,N_7713);
nor U10069 (N_10069,N_6522,N_6353);
and U10070 (N_10070,N_6152,N_7777);
or U10071 (N_10071,N_8988,N_7593);
nor U10072 (N_10072,N_6455,N_7793);
nand U10073 (N_10073,N_8692,N_7545);
nand U10074 (N_10074,N_8231,N_6708);
or U10075 (N_10075,N_6426,N_7191);
and U10076 (N_10076,N_7048,N_7258);
or U10077 (N_10077,N_6003,N_8062);
nor U10078 (N_10078,N_6722,N_6608);
nor U10079 (N_10079,N_8989,N_7555);
or U10080 (N_10080,N_8334,N_6878);
or U10081 (N_10081,N_6063,N_8047);
xnor U10082 (N_10082,N_7547,N_8864);
and U10083 (N_10083,N_8432,N_6760);
and U10084 (N_10084,N_7753,N_7695);
nand U10085 (N_10085,N_8849,N_8307);
xnor U10086 (N_10086,N_7724,N_8953);
or U10087 (N_10087,N_7498,N_8748);
and U10088 (N_10088,N_6777,N_7751);
or U10089 (N_10089,N_6855,N_6366);
nand U10090 (N_10090,N_8802,N_6787);
or U10091 (N_10091,N_6500,N_6766);
nand U10092 (N_10092,N_8101,N_7865);
nand U10093 (N_10093,N_7683,N_6579);
nor U10094 (N_10094,N_6442,N_7180);
or U10095 (N_10095,N_6273,N_7145);
or U10096 (N_10096,N_8608,N_8647);
and U10097 (N_10097,N_7469,N_7415);
and U10098 (N_10098,N_8630,N_7622);
nand U10099 (N_10099,N_6456,N_6298);
xnor U10100 (N_10100,N_7633,N_6208);
or U10101 (N_10101,N_7162,N_8469);
or U10102 (N_10102,N_8964,N_7266);
nand U10103 (N_10103,N_7373,N_6318);
xor U10104 (N_10104,N_7743,N_6752);
xor U10105 (N_10105,N_8244,N_8051);
nand U10106 (N_10106,N_8576,N_8347);
or U10107 (N_10107,N_8789,N_6033);
or U10108 (N_10108,N_8435,N_6148);
nor U10109 (N_10109,N_7712,N_6343);
or U10110 (N_10110,N_7629,N_6895);
nand U10111 (N_10111,N_7572,N_6711);
xor U10112 (N_10112,N_6474,N_8233);
xnor U10113 (N_10113,N_8747,N_8830);
or U10114 (N_10114,N_8110,N_7798);
or U10115 (N_10115,N_8583,N_8058);
xnor U10116 (N_10116,N_7752,N_6920);
nor U10117 (N_10117,N_8694,N_8317);
and U10118 (N_10118,N_6150,N_7290);
xnor U10119 (N_10119,N_6585,N_6690);
nand U10120 (N_10120,N_6352,N_7704);
nor U10121 (N_10121,N_7461,N_7484);
nand U10122 (N_10122,N_8276,N_8179);
xor U10123 (N_10123,N_8967,N_8834);
and U10124 (N_10124,N_8092,N_7092);
or U10125 (N_10125,N_6978,N_6115);
and U10126 (N_10126,N_6032,N_7149);
nand U10127 (N_10127,N_6864,N_7654);
and U10128 (N_10128,N_8009,N_6468);
and U10129 (N_10129,N_8079,N_8150);
or U10130 (N_10130,N_8793,N_7166);
nor U10131 (N_10131,N_6962,N_8365);
nor U10132 (N_10132,N_6288,N_6998);
xor U10133 (N_10133,N_7060,N_6574);
and U10134 (N_10134,N_7728,N_6627);
and U10135 (N_10135,N_6974,N_6869);
and U10136 (N_10136,N_7768,N_6923);
or U10137 (N_10137,N_8975,N_8621);
nor U10138 (N_10138,N_6310,N_6534);
and U10139 (N_10139,N_7133,N_8181);
and U10140 (N_10140,N_6634,N_8968);
or U10141 (N_10141,N_7896,N_6823);
nand U10142 (N_10142,N_8672,N_7792);
xnor U10143 (N_10143,N_7942,N_7485);
nand U10144 (N_10144,N_6572,N_6887);
nor U10145 (N_10145,N_6837,N_8799);
nor U10146 (N_10146,N_8351,N_6361);
and U10147 (N_10147,N_6815,N_6750);
and U10148 (N_10148,N_6549,N_6728);
nor U10149 (N_10149,N_8860,N_6732);
or U10150 (N_10150,N_7147,N_8098);
nor U10151 (N_10151,N_7773,N_8072);
or U10152 (N_10152,N_7341,N_6497);
nor U10153 (N_10153,N_7207,N_7480);
nor U10154 (N_10154,N_8004,N_7811);
nand U10155 (N_10155,N_8745,N_7721);
nor U10156 (N_10156,N_6107,N_6206);
nand U10157 (N_10157,N_6061,N_8320);
or U10158 (N_10158,N_7708,N_7778);
nor U10159 (N_10159,N_6279,N_8437);
nand U10160 (N_10160,N_8902,N_7361);
nor U10161 (N_10161,N_8926,N_8697);
and U10162 (N_10162,N_8822,N_8013);
xor U10163 (N_10163,N_6239,N_6479);
nand U10164 (N_10164,N_7322,N_7829);
nor U10165 (N_10165,N_8312,N_6038);
and U10166 (N_10166,N_7031,N_8904);
nand U10167 (N_10167,N_6785,N_8270);
nand U10168 (N_10168,N_7030,N_7401);
and U10169 (N_10169,N_6488,N_7651);
or U10170 (N_10170,N_8480,N_7445);
nand U10171 (N_10171,N_7644,N_7350);
nor U10172 (N_10172,N_7635,N_6853);
or U10173 (N_10173,N_7961,N_7537);
xnor U10174 (N_10174,N_6630,N_8441);
nor U10175 (N_10175,N_7259,N_6900);
and U10176 (N_10176,N_6907,N_6200);
nor U10177 (N_10177,N_7176,N_6614);
nor U10178 (N_10178,N_7647,N_6626);
nor U10179 (N_10179,N_6407,N_8982);
nor U10180 (N_10180,N_8784,N_7302);
nand U10181 (N_10181,N_7392,N_7937);
and U10182 (N_10182,N_7301,N_8160);
nor U10183 (N_10183,N_8184,N_8438);
xor U10184 (N_10184,N_8922,N_8892);
and U10185 (N_10185,N_6203,N_6390);
nor U10186 (N_10186,N_8357,N_6379);
or U10187 (N_10187,N_6246,N_8074);
nor U10188 (N_10188,N_6283,N_6166);
and U10189 (N_10189,N_6175,N_6266);
or U10190 (N_10190,N_6986,N_8783);
nor U10191 (N_10191,N_6903,N_7131);
nand U10192 (N_10192,N_7564,N_6851);
nand U10193 (N_10193,N_8613,N_6432);
nand U10194 (N_10194,N_6308,N_7605);
and U10195 (N_10195,N_6688,N_8551);
nand U10196 (N_10196,N_6995,N_6092);
nand U10197 (N_10197,N_7905,N_7736);
nand U10198 (N_10198,N_6395,N_7862);
and U10199 (N_10199,N_8950,N_6275);
nor U10200 (N_10200,N_8612,N_6282);
nor U10201 (N_10201,N_8669,N_8127);
nand U10202 (N_10202,N_6824,N_8085);
nand U10203 (N_10203,N_8082,N_7125);
nor U10204 (N_10204,N_6590,N_6215);
xor U10205 (N_10205,N_7308,N_8486);
nor U10206 (N_10206,N_7328,N_8711);
nor U10207 (N_10207,N_8691,N_6475);
or U10208 (N_10208,N_7796,N_6125);
nor U10209 (N_10209,N_6141,N_8795);
and U10210 (N_10210,N_8303,N_8407);
and U10211 (N_10211,N_8242,N_8560);
or U10212 (N_10212,N_8015,N_6349);
nand U10213 (N_10213,N_7066,N_6194);
nor U10214 (N_10214,N_8751,N_6905);
xor U10215 (N_10215,N_6525,N_6248);
and U10216 (N_10216,N_7024,N_6922);
and U10217 (N_10217,N_7847,N_8840);
and U10218 (N_10218,N_7817,N_8169);
nor U10219 (N_10219,N_6004,N_6363);
nor U10220 (N_10220,N_6330,N_6935);
or U10221 (N_10221,N_7560,N_8575);
nor U10222 (N_10222,N_8609,N_6857);
nand U10223 (N_10223,N_7309,N_8245);
and U10224 (N_10224,N_7393,N_8187);
nand U10225 (N_10225,N_8670,N_8497);
nand U10226 (N_10226,N_8870,N_7192);
nor U10227 (N_10227,N_8824,N_7689);
or U10228 (N_10228,N_6358,N_8639);
nor U10229 (N_10229,N_8664,N_8239);
nor U10230 (N_10230,N_6975,N_6691);
nand U10231 (N_10231,N_7470,N_6041);
or U10232 (N_10232,N_6757,N_7675);
xnor U10233 (N_10233,N_7565,N_8665);
and U10234 (N_10234,N_7006,N_6831);
or U10235 (N_10235,N_6084,N_6408);
and U10236 (N_10236,N_6856,N_8889);
and U10237 (N_10237,N_7568,N_7435);
or U10238 (N_10238,N_6678,N_8884);
and U10239 (N_10239,N_6392,N_8302);
and U10240 (N_10240,N_6109,N_6357);
or U10241 (N_10241,N_7649,N_8876);
nand U10242 (N_10242,N_6535,N_8874);
and U10243 (N_10243,N_7118,N_6322);
xnor U10244 (N_10244,N_6852,N_6536);
xor U10245 (N_10245,N_7697,N_8858);
nand U10246 (N_10246,N_7834,N_8701);
and U10247 (N_10247,N_6130,N_7386);
nand U10248 (N_10248,N_6385,N_6809);
and U10249 (N_10249,N_6091,N_7500);
or U10250 (N_10250,N_7738,N_7528);
nand U10251 (N_10251,N_6947,N_6304);
and U10252 (N_10252,N_7627,N_7857);
nor U10253 (N_10253,N_7676,N_8523);
and U10254 (N_10254,N_6214,N_7375);
and U10255 (N_10255,N_8593,N_8373);
xor U10256 (N_10256,N_7384,N_8279);
nand U10257 (N_10257,N_6792,N_7022);
and U10258 (N_10258,N_7144,N_6977);
or U10259 (N_10259,N_8971,N_6604);
nand U10260 (N_10260,N_6926,N_8758);
and U10261 (N_10261,N_8667,N_8249);
nor U10262 (N_10262,N_7779,N_8400);
and U10263 (N_10263,N_6055,N_8491);
and U10264 (N_10264,N_7020,N_6046);
nor U10265 (N_10265,N_7335,N_8093);
nor U10266 (N_10266,N_6925,N_7296);
nor U10267 (N_10267,N_7501,N_8246);
nor U10268 (N_10268,N_6010,N_8253);
and U10269 (N_10269,N_8804,N_7782);
xnor U10270 (N_10270,N_7897,N_8412);
nand U10271 (N_10271,N_8651,N_8709);
nand U10272 (N_10272,N_7579,N_6508);
and U10273 (N_10273,N_8374,N_7113);
and U10274 (N_10274,N_8037,N_8749);
nand U10275 (N_10275,N_8423,N_6644);
nand U10276 (N_10276,N_7454,N_6354);
or U10277 (N_10277,N_7822,N_7056);
and U10278 (N_10278,N_7864,N_6898);
nand U10279 (N_10279,N_8289,N_8731);
or U10280 (N_10280,N_7334,N_6821);
nand U10281 (N_10281,N_6499,N_7586);
nor U10282 (N_10282,N_6699,N_7770);
and U10283 (N_10283,N_8946,N_6252);
and U10284 (N_10284,N_6633,N_7103);
xor U10285 (N_10285,N_8515,N_8097);
or U10286 (N_10286,N_6156,N_8951);
nor U10287 (N_10287,N_8325,N_7551);
and U10288 (N_10288,N_6300,N_8413);
or U10289 (N_10289,N_8724,N_8477);
and U10290 (N_10290,N_7110,N_8517);
xnor U10291 (N_10291,N_8512,N_8942);
xnor U10292 (N_10292,N_7923,N_8114);
and U10293 (N_10293,N_8025,N_6466);
and U10294 (N_10294,N_6396,N_6296);
or U10295 (N_10295,N_8265,N_6946);
nand U10296 (N_10296,N_6104,N_7340);
nor U10297 (N_10297,N_8256,N_6694);
xnor U10298 (N_10298,N_7525,N_7899);
or U10299 (N_10299,N_8084,N_8230);
nor U10300 (N_10300,N_7608,N_8163);
and U10301 (N_10301,N_8414,N_6601);
nand U10302 (N_10302,N_8342,N_8107);
xor U10303 (N_10303,N_7638,N_7114);
nor U10304 (N_10304,N_6244,N_7594);
or U10305 (N_10305,N_8421,N_6744);
xor U10306 (N_10306,N_6504,N_8096);
and U10307 (N_10307,N_6774,N_8752);
xnor U10308 (N_10308,N_6146,N_6326);
or U10309 (N_10309,N_8212,N_8805);
and U10310 (N_10310,N_7037,N_6207);
and U10311 (N_10311,N_6558,N_6529);
or U10312 (N_10312,N_6057,N_6518);
nor U10313 (N_10313,N_7409,N_6122);
nand U10314 (N_10314,N_6709,N_7245);
or U10315 (N_10315,N_8420,N_8923);
nand U10316 (N_10316,N_7021,N_6422);
nor U10317 (N_10317,N_7997,N_6112);
or U10318 (N_10318,N_7109,N_8919);
or U10319 (N_10319,N_7880,N_7533);
xnor U10320 (N_10320,N_6679,N_6202);
nand U10321 (N_10321,N_7130,N_6097);
or U10322 (N_10322,N_7238,N_7844);
nor U10323 (N_10323,N_8997,N_6346);
and U10324 (N_10324,N_8803,N_7467);
and U10325 (N_10325,N_6523,N_7391);
or U10326 (N_10326,N_8217,N_6224);
and U10327 (N_10327,N_8418,N_7672);
xnor U10328 (N_10328,N_6916,N_8052);
and U10329 (N_10329,N_7548,N_7790);
nor U10330 (N_10330,N_6717,N_6800);
and U10331 (N_10331,N_6093,N_7574);
or U10332 (N_10332,N_7506,N_8980);
and U10333 (N_10333,N_8675,N_8539);
or U10334 (N_10334,N_6355,N_7677);
nor U10335 (N_10335,N_8316,N_8021);
nand U10336 (N_10336,N_6313,N_6356);
and U10337 (N_10337,N_7234,N_6199);
and U10338 (N_10338,N_8032,N_8582);
nand U10339 (N_10339,N_6059,N_8496);
nor U10340 (N_10340,N_6434,N_7465);
and U10341 (N_10341,N_7212,N_6249);
xor U10342 (N_10342,N_8561,N_8767);
and U10343 (N_10343,N_8581,N_7434);
and U10344 (N_10344,N_6593,N_7553);
nand U10345 (N_10345,N_7588,N_7405);
and U10346 (N_10346,N_8290,N_6031);
or U10347 (N_10347,N_7673,N_7511);
or U10348 (N_10348,N_6305,N_7585);
xor U10349 (N_10349,N_7575,N_6663);
and U10350 (N_10350,N_7198,N_8589);
nor U10351 (N_10351,N_8915,N_6111);
nand U10352 (N_10352,N_7730,N_6172);
xnor U10353 (N_10353,N_6502,N_7121);
nand U10354 (N_10354,N_7775,N_7174);
nor U10355 (N_10355,N_6770,N_7503);
xnor U10356 (N_10356,N_6452,N_8739);
xor U10357 (N_10357,N_8869,N_8293);
or U10358 (N_10358,N_6428,N_8979);
and U10359 (N_10359,N_7913,N_6170);
or U10360 (N_10360,N_8045,N_7519);
nor U10361 (N_10361,N_7903,N_8766);
nor U10362 (N_10362,N_6751,N_6120);
and U10363 (N_10363,N_8871,N_6081);
xor U10364 (N_10364,N_8939,N_7028);
nand U10365 (N_10365,N_6814,N_6495);
or U10366 (N_10366,N_6204,N_8221);
or U10367 (N_10367,N_8381,N_8416);
or U10368 (N_10368,N_7143,N_6068);
or U10369 (N_10369,N_6997,N_6015);
nor U10370 (N_10370,N_7694,N_6001);
and U10371 (N_10371,N_6443,N_6908);
and U10372 (N_10372,N_7460,N_7287);
and U10373 (N_10373,N_8825,N_7319);
or U10374 (N_10374,N_7881,N_8907);
nor U10375 (N_10375,N_8287,N_8170);
nor U10376 (N_10376,N_8954,N_8704);
and U10377 (N_10377,N_7974,N_8454);
or U10378 (N_10378,N_8448,N_7918);
or U10379 (N_10379,N_6339,N_8610);
nand U10380 (N_10380,N_6902,N_8698);
nand U10381 (N_10381,N_6896,N_7929);
or U10382 (N_10382,N_6551,N_6697);
nand U10383 (N_10383,N_8399,N_8839);
nor U10384 (N_10384,N_7891,N_8136);
xnor U10385 (N_10385,N_8309,N_7424);
nor U10386 (N_10386,N_7906,N_6530);
nand U10387 (N_10387,N_7106,N_7489);
or U10388 (N_10388,N_6340,N_8131);
and U10389 (N_10389,N_8439,N_6718);
nand U10390 (N_10390,N_7084,N_6116);
or U10391 (N_10391,N_7729,N_7970);
and U10392 (N_10392,N_6386,N_8543);
nor U10393 (N_10393,N_7033,N_8653);
and U10394 (N_10394,N_8319,N_7581);
nand U10395 (N_10395,N_7165,N_6742);
and U10396 (N_10396,N_7315,N_8592);
and U10397 (N_10397,N_7657,N_6514);
and U10398 (N_10398,N_6835,N_7466);
nor U10399 (N_10399,N_6956,N_6938);
and U10400 (N_10400,N_6812,N_8528);
or U10401 (N_10401,N_6077,N_8873);
nor U10402 (N_10402,N_7733,N_8933);
or U10403 (N_10403,N_7385,N_7000);
nand U10404 (N_10404,N_8141,N_8601);
or U10405 (N_10405,N_8484,N_6924);
nor U10406 (N_10406,N_7293,N_6818);
nand U10407 (N_10407,N_6295,N_6384);
or U10408 (N_10408,N_7183,N_7182);
nor U10409 (N_10409,N_6876,N_8550);
nor U10410 (N_10410,N_6467,N_7289);
and U10411 (N_10411,N_8557,N_6070);
nand U10412 (N_10412,N_7246,N_8525);
xor U10413 (N_10413,N_8091,N_7294);
nor U10414 (N_10414,N_7277,N_6371);
nor U10415 (N_10415,N_7070,N_6256);
nor U10416 (N_10416,N_7893,N_8147);
and U10417 (N_10417,N_8076,N_8402);
nor U10418 (N_10418,N_7316,N_7910);
nor U10419 (N_10419,N_6858,N_7940);
or U10420 (N_10420,N_8116,N_8377);
nor U10421 (N_10421,N_7693,N_8716);
nand U10422 (N_10422,N_7444,N_7029);
and U10423 (N_10423,N_8327,N_8174);
nor U10424 (N_10424,N_6820,N_6655);
nor U10425 (N_10425,N_6870,N_8394);
nand U10426 (N_10426,N_8135,N_7261);
nor U10427 (N_10427,N_6652,N_7089);
nand U10428 (N_10428,N_6192,N_6620);
nand U10429 (N_10429,N_7526,N_7055);
nand U10430 (N_10430,N_7459,N_6736);
nand U10431 (N_10431,N_7097,N_7389);
xor U10432 (N_10432,N_6942,N_8277);
or U10433 (N_10433,N_7948,N_8574);
nor U10434 (N_10434,N_7481,N_6632);
nand U10435 (N_10435,N_7766,N_7814);
nand U10436 (N_10436,N_8262,N_7211);
and U10437 (N_10437,N_7960,N_8326);
nand U10438 (N_10438,N_7747,N_6959);
or U10439 (N_10439,N_7152,N_6936);
nor U10440 (N_10440,N_6123,N_8175);
nor U10441 (N_10441,N_7120,N_8944);
nor U10442 (N_10442,N_7005,N_8567);
nand U10443 (N_10443,N_6071,N_8507);
or U10444 (N_10444,N_7599,N_8133);
xnor U10445 (N_10445,N_8196,N_6854);
and U10446 (N_10446,N_6698,N_8765);
nand U10447 (N_10447,N_6323,N_6388);
and U10448 (N_10448,N_8063,N_6638);
and U10449 (N_10449,N_8755,N_8121);
nand U10450 (N_10450,N_7838,N_6894);
nor U10451 (N_10451,N_7901,N_7854);
nor U10452 (N_10452,N_8632,N_6190);
nand U10453 (N_10453,N_8674,N_7892);
nor U10454 (N_10454,N_6667,N_6859);
nor U10455 (N_10455,N_6242,N_8049);
nand U10456 (N_10456,N_7035,N_7856);
or U10457 (N_10457,N_8721,N_7742);
and U10458 (N_10458,N_8633,N_6810);
nor U10459 (N_10459,N_8920,N_8736);
nand U10460 (N_10460,N_8036,N_8580);
or U10461 (N_10461,N_8026,N_7851);
nor U10462 (N_10462,N_8066,N_8738);
nand U10463 (N_10463,N_7725,N_7414);
nor U10464 (N_10464,N_8006,N_6930);
nor U10465 (N_10465,N_6005,N_7135);
and U10466 (N_10466,N_7539,N_7628);
or U10467 (N_10467,N_6174,N_7616);
nor U10468 (N_10468,N_8367,N_6743);
and U10469 (N_10469,N_7727,N_8777);
and U10470 (N_10470,N_8510,N_6737);
nor U10471 (N_10471,N_7801,N_6552);
nor U10472 (N_10472,N_6161,N_7275);
and U10473 (N_10473,N_8705,N_8390);
and U10474 (N_10474,N_7987,N_6317);
and U10475 (N_10475,N_6746,N_8808);
nand U10476 (N_10476,N_6401,N_7493);
nor U10477 (N_10477,N_6088,N_8271);
nand U10478 (N_10478,N_6625,N_8392);
or U10479 (N_10479,N_7931,N_7223);
and U10480 (N_10480,N_8677,N_6546);
xnor U10481 (N_10481,N_7154,N_6449);
nor U10482 (N_10482,N_6049,N_6803);
nand U10483 (N_10483,N_8467,N_8836);
nor U10484 (N_10484,N_8809,N_8679);
nor U10485 (N_10485,N_8548,N_8974);
nand U10486 (N_10486,N_8012,N_8537);
nor U10487 (N_10487,N_8372,N_7129);
or U10488 (N_10488,N_7839,N_7239);
or U10489 (N_10489,N_6651,N_8591);
or U10490 (N_10490,N_8852,N_8678);
or U10491 (N_10491,N_6793,N_7069);
nand U10492 (N_10492,N_8703,N_8137);
nand U10493 (N_10493,N_8529,N_6006);
or U10494 (N_10494,N_8987,N_7357);
nand U10495 (N_10495,N_8573,N_7054);
nand U10496 (N_10496,N_6584,N_6676);
nor U10497 (N_10497,N_8715,N_7167);
or U10498 (N_10498,N_6740,N_7194);
nand U10499 (N_10499,N_6337,N_6205);
nand U10500 (N_10500,N_8974,N_8938);
xnor U10501 (N_10501,N_8019,N_6840);
and U10502 (N_10502,N_8843,N_8745);
or U10503 (N_10503,N_8292,N_7024);
nand U10504 (N_10504,N_6019,N_8196);
nor U10505 (N_10505,N_6126,N_8701);
and U10506 (N_10506,N_6240,N_7204);
and U10507 (N_10507,N_6791,N_8098);
nand U10508 (N_10508,N_7568,N_8021);
and U10509 (N_10509,N_8521,N_7545);
xor U10510 (N_10510,N_6632,N_6291);
or U10511 (N_10511,N_8387,N_6735);
and U10512 (N_10512,N_7096,N_7222);
nand U10513 (N_10513,N_7024,N_6360);
or U10514 (N_10514,N_7570,N_6905);
nand U10515 (N_10515,N_7106,N_7364);
or U10516 (N_10516,N_6533,N_7477);
nand U10517 (N_10517,N_8338,N_6604);
xnor U10518 (N_10518,N_6888,N_6023);
or U10519 (N_10519,N_8856,N_7058);
and U10520 (N_10520,N_8539,N_6482);
nand U10521 (N_10521,N_7419,N_7994);
or U10522 (N_10522,N_6325,N_8968);
nor U10523 (N_10523,N_6295,N_6794);
or U10524 (N_10524,N_8960,N_8094);
and U10525 (N_10525,N_8335,N_6636);
nand U10526 (N_10526,N_6407,N_7123);
nor U10527 (N_10527,N_7896,N_6971);
and U10528 (N_10528,N_8194,N_6407);
or U10529 (N_10529,N_7377,N_7676);
nand U10530 (N_10530,N_7939,N_6184);
xnor U10531 (N_10531,N_7988,N_7006);
and U10532 (N_10532,N_7663,N_6394);
nand U10533 (N_10533,N_6721,N_7589);
xnor U10534 (N_10534,N_6209,N_6041);
nor U10535 (N_10535,N_6057,N_7999);
nor U10536 (N_10536,N_6004,N_7534);
or U10537 (N_10537,N_8323,N_8833);
nor U10538 (N_10538,N_7226,N_8605);
and U10539 (N_10539,N_7214,N_7226);
nand U10540 (N_10540,N_7451,N_8830);
xnor U10541 (N_10541,N_7427,N_8193);
and U10542 (N_10542,N_6586,N_6308);
xor U10543 (N_10543,N_8077,N_7119);
nand U10544 (N_10544,N_8399,N_8967);
nor U10545 (N_10545,N_8917,N_7015);
or U10546 (N_10546,N_7600,N_8894);
nand U10547 (N_10547,N_6451,N_7077);
nor U10548 (N_10548,N_6207,N_7193);
and U10549 (N_10549,N_6484,N_8233);
nand U10550 (N_10550,N_7813,N_6629);
nor U10551 (N_10551,N_6738,N_6598);
nand U10552 (N_10552,N_7325,N_7355);
xnor U10553 (N_10553,N_6797,N_6120);
and U10554 (N_10554,N_7620,N_8511);
nand U10555 (N_10555,N_7691,N_7085);
and U10556 (N_10556,N_6279,N_7195);
or U10557 (N_10557,N_8554,N_8161);
or U10558 (N_10558,N_7382,N_7646);
xor U10559 (N_10559,N_6639,N_7993);
nor U10560 (N_10560,N_8798,N_8206);
nor U10561 (N_10561,N_7374,N_7646);
and U10562 (N_10562,N_6298,N_8099);
nor U10563 (N_10563,N_7876,N_7476);
nand U10564 (N_10564,N_6049,N_6889);
nor U10565 (N_10565,N_6229,N_8379);
nand U10566 (N_10566,N_8107,N_8408);
nand U10567 (N_10567,N_8685,N_7300);
xor U10568 (N_10568,N_6849,N_8640);
and U10569 (N_10569,N_8846,N_7476);
xor U10570 (N_10570,N_8271,N_6600);
and U10571 (N_10571,N_8205,N_8497);
nor U10572 (N_10572,N_8424,N_6971);
nor U10573 (N_10573,N_6968,N_7454);
nand U10574 (N_10574,N_6388,N_8628);
and U10575 (N_10575,N_7187,N_7001);
and U10576 (N_10576,N_6281,N_6282);
nand U10577 (N_10577,N_8034,N_8459);
nand U10578 (N_10578,N_8041,N_8099);
or U10579 (N_10579,N_8081,N_6256);
or U10580 (N_10580,N_6855,N_8381);
nor U10581 (N_10581,N_6623,N_7737);
nand U10582 (N_10582,N_7498,N_7236);
and U10583 (N_10583,N_6086,N_8535);
and U10584 (N_10584,N_7347,N_8995);
nand U10585 (N_10585,N_6297,N_7372);
or U10586 (N_10586,N_8735,N_6526);
and U10587 (N_10587,N_6040,N_8661);
nor U10588 (N_10588,N_7779,N_8054);
nor U10589 (N_10589,N_8392,N_7581);
and U10590 (N_10590,N_8091,N_8828);
xnor U10591 (N_10591,N_6183,N_7681);
and U10592 (N_10592,N_8967,N_8510);
nand U10593 (N_10593,N_8942,N_7307);
or U10594 (N_10594,N_7775,N_7447);
or U10595 (N_10595,N_7268,N_8493);
and U10596 (N_10596,N_7955,N_8371);
and U10597 (N_10597,N_6327,N_6512);
nor U10598 (N_10598,N_8748,N_8132);
or U10599 (N_10599,N_6714,N_7134);
and U10600 (N_10600,N_7602,N_7884);
nor U10601 (N_10601,N_6698,N_8780);
nor U10602 (N_10602,N_6397,N_6290);
or U10603 (N_10603,N_6346,N_6003);
nor U10604 (N_10604,N_7096,N_8346);
nor U10605 (N_10605,N_7302,N_6046);
nand U10606 (N_10606,N_7585,N_7410);
nor U10607 (N_10607,N_8822,N_6974);
nor U10608 (N_10608,N_6934,N_6025);
nor U10609 (N_10609,N_6804,N_8954);
nor U10610 (N_10610,N_8085,N_6373);
or U10611 (N_10611,N_7350,N_6004);
and U10612 (N_10612,N_7999,N_7802);
nor U10613 (N_10613,N_7052,N_6163);
nor U10614 (N_10614,N_7003,N_7973);
or U10615 (N_10615,N_7810,N_8052);
and U10616 (N_10616,N_8733,N_7949);
and U10617 (N_10617,N_7525,N_7181);
nor U10618 (N_10618,N_8473,N_7163);
xor U10619 (N_10619,N_6363,N_8819);
and U10620 (N_10620,N_6532,N_6884);
nor U10621 (N_10621,N_6011,N_7370);
nor U10622 (N_10622,N_8710,N_8812);
nand U10623 (N_10623,N_8680,N_7231);
nand U10624 (N_10624,N_8681,N_8314);
xnor U10625 (N_10625,N_6794,N_6426);
or U10626 (N_10626,N_7826,N_7418);
nor U10627 (N_10627,N_7327,N_8467);
nor U10628 (N_10628,N_6035,N_6086);
or U10629 (N_10629,N_8446,N_8428);
nand U10630 (N_10630,N_8798,N_6969);
or U10631 (N_10631,N_7904,N_8165);
nor U10632 (N_10632,N_8184,N_6272);
nand U10633 (N_10633,N_6341,N_6859);
nand U10634 (N_10634,N_7417,N_8345);
or U10635 (N_10635,N_8059,N_7485);
nand U10636 (N_10636,N_7328,N_6625);
xnor U10637 (N_10637,N_8409,N_6260);
nor U10638 (N_10638,N_8768,N_6242);
nor U10639 (N_10639,N_7887,N_8262);
nor U10640 (N_10640,N_8340,N_8782);
nand U10641 (N_10641,N_8776,N_7876);
nor U10642 (N_10642,N_7798,N_8446);
xor U10643 (N_10643,N_7654,N_8579);
nor U10644 (N_10644,N_6501,N_6916);
or U10645 (N_10645,N_6547,N_7706);
or U10646 (N_10646,N_7573,N_7523);
or U10647 (N_10647,N_6369,N_8127);
xor U10648 (N_10648,N_6763,N_7740);
nor U10649 (N_10649,N_7280,N_7936);
and U10650 (N_10650,N_8163,N_7651);
nor U10651 (N_10651,N_7703,N_8454);
nor U10652 (N_10652,N_8557,N_8499);
nand U10653 (N_10653,N_8807,N_7356);
nor U10654 (N_10654,N_8325,N_8944);
nand U10655 (N_10655,N_7297,N_7894);
nor U10656 (N_10656,N_7858,N_8588);
nand U10657 (N_10657,N_6288,N_7449);
nand U10658 (N_10658,N_8499,N_8366);
nand U10659 (N_10659,N_7049,N_7173);
nor U10660 (N_10660,N_7510,N_6116);
nand U10661 (N_10661,N_6907,N_7210);
and U10662 (N_10662,N_7752,N_8993);
nand U10663 (N_10663,N_8717,N_8104);
and U10664 (N_10664,N_7720,N_8487);
or U10665 (N_10665,N_7444,N_8281);
nor U10666 (N_10666,N_7649,N_7217);
nor U10667 (N_10667,N_6010,N_7945);
xor U10668 (N_10668,N_6321,N_7752);
nor U10669 (N_10669,N_7152,N_6604);
nand U10670 (N_10670,N_7209,N_6296);
xnor U10671 (N_10671,N_7883,N_8342);
nand U10672 (N_10672,N_6969,N_6598);
and U10673 (N_10673,N_7016,N_6242);
or U10674 (N_10674,N_6813,N_6117);
nor U10675 (N_10675,N_6381,N_7049);
nand U10676 (N_10676,N_6021,N_7651);
xor U10677 (N_10677,N_8666,N_8704);
nand U10678 (N_10678,N_7551,N_6740);
and U10679 (N_10679,N_6325,N_7177);
and U10680 (N_10680,N_6230,N_7978);
nor U10681 (N_10681,N_7288,N_7465);
nand U10682 (N_10682,N_8340,N_7185);
and U10683 (N_10683,N_7220,N_6321);
nand U10684 (N_10684,N_6789,N_8280);
nor U10685 (N_10685,N_6714,N_6845);
and U10686 (N_10686,N_7183,N_6578);
nor U10687 (N_10687,N_7853,N_8607);
nand U10688 (N_10688,N_8426,N_8810);
or U10689 (N_10689,N_7929,N_6331);
nand U10690 (N_10690,N_7368,N_6537);
or U10691 (N_10691,N_8819,N_7267);
or U10692 (N_10692,N_6822,N_7644);
and U10693 (N_10693,N_7580,N_6909);
xor U10694 (N_10694,N_7313,N_6579);
xnor U10695 (N_10695,N_7705,N_8203);
nand U10696 (N_10696,N_8314,N_7891);
nor U10697 (N_10697,N_7538,N_6049);
and U10698 (N_10698,N_8737,N_7045);
or U10699 (N_10699,N_7118,N_7378);
nand U10700 (N_10700,N_8130,N_6695);
or U10701 (N_10701,N_6251,N_7004);
xnor U10702 (N_10702,N_6885,N_8192);
xor U10703 (N_10703,N_7795,N_7123);
nand U10704 (N_10704,N_7279,N_6575);
or U10705 (N_10705,N_6216,N_7929);
and U10706 (N_10706,N_8084,N_6507);
nand U10707 (N_10707,N_6443,N_6429);
or U10708 (N_10708,N_6940,N_8557);
xnor U10709 (N_10709,N_8193,N_8512);
nand U10710 (N_10710,N_6191,N_7335);
and U10711 (N_10711,N_8707,N_8028);
xor U10712 (N_10712,N_6325,N_7706);
and U10713 (N_10713,N_7346,N_6149);
and U10714 (N_10714,N_7538,N_8627);
nand U10715 (N_10715,N_6215,N_7132);
nor U10716 (N_10716,N_6664,N_8642);
nor U10717 (N_10717,N_7416,N_6467);
or U10718 (N_10718,N_8441,N_6179);
or U10719 (N_10719,N_6508,N_8871);
and U10720 (N_10720,N_8955,N_8679);
nand U10721 (N_10721,N_7167,N_6818);
nand U10722 (N_10722,N_6598,N_6918);
nor U10723 (N_10723,N_6855,N_6644);
and U10724 (N_10724,N_6937,N_8006);
nor U10725 (N_10725,N_7317,N_7520);
nand U10726 (N_10726,N_6337,N_6832);
or U10727 (N_10727,N_8510,N_6454);
and U10728 (N_10728,N_6975,N_7597);
or U10729 (N_10729,N_8474,N_7803);
nand U10730 (N_10730,N_7530,N_7549);
nor U10731 (N_10731,N_6235,N_7380);
and U10732 (N_10732,N_6676,N_6486);
xor U10733 (N_10733,N_7051,N_7823);
nand U10734 (N_10734,N_7408,N_8227);
and U10735 (N_10735,N_8077,N_7073);
nor U10736 (N_10736,N_8638,N_6162);
and U10737 (N_10737,N_7436,N_8655);
and U10738 (N_10738,N_8182,N_6726);
nor U10739 (N_10739,N_6069,N_7500);
nand U10740 (N_10740,N_6940,N_7006);
nand U10741 (N_10741,N_8484,N_6778);
or U10742 (N_10742,N_8288,N_8703);
xor U10743 (N_10743,N_6741,N_7150);
nand U10744 (N_10744,N_8887,N_7650);
or U10745 (N_10745,N_6407,N_8431);
nor U10746 (N_10746,N_6994,N_6118);
and U10747 (N_10747,N_7061,N_7575);
nor U10748 (N_10748,N_8267,N_6557);
nor U10749 (N_10749,N_8066,N_7486);
nor U10750 (N_10750,N_8058,N_6374);
nand U10751 (N_10751,N_6949,N_8526);
or U10752 (N_10752,N_6680,N_7127);
nand U10753 (N_10753,N_8131,N_7000);
nor U10754 (N_10754,N_7636,N_6553);
nand U10755 (N_10755,N_8924,N_8845);
and U10756 (N_10756,N_6406,N_6382);
xor U10757 (N_10757,N_8158,N_8016);
or U10758 (N_10758,N_8251,N_7177);
nand U10759 (N_10759,N_6688,N_8536);
and U10760 (N_10760,N_8710,N_7616);
and U10761 (N_10761,N_8805,N_8988);
or U10762 (N_10762,N_7911,N_7302);
or U10763 (N_10763,N_7027,N_7302);
and U10764 (N_10764,N_7008,N_6985);
and U10765 (N_10765,N_8204,N_7774);
or U10766 (N_10766,N_8904,N_6775);
nand U10767 (N_10767,N_6312,N_6670);
nand U10768 (N_10768,N_7579,N_6433);
and U10769 (N_10769,N_6595,N_7709);
or U10770 (N_10770,N_6798,N_7960);
and U10771 (N_10771,N_8397,N_6688);
nor U10772 (N_10772,N_6190,N_8065);
and U10773 (N_10773,N_7933,N_8942);
nor U10774 (N_10774,N_7672,N_7750);
and U10775 (N_10775,N_6595,N_7397);
nand U10776 (N_10776,N_7387,N_6995);
and U10777 (N_10777,N_6738,N_6534);
nor U10778 (N_10778,N_8410,N_6606);
nand U10779 (N_10779,N_6895,N_6202);
nand U10780 (N_10780,N_8776,N_8036);
xor U10781 (N_10781,N_8502,N_6844);
or U10782 (N_10782,N_6526,N_8346);
or U10783 (N_10783,N_6961,N_7981);
or U10784 (N_10784,N_7764,N_6205);
nor U10785 (N_10785,N_8108,N_8382);
and U10786 (N_10786,N_8585,N_8862);
nor U10787 (N_10787,N_7070,N_8296);
and U10788 (N_10788,N_8829,N_6828);
nand U10789 (N_10789,N_8376,N_8019);
or U10790 (N_10790,N_8272,N_8313);
nand U10791 (N_10791,N_8688,N_8265);
nand U10792 (N_10792,N_7469,N_7454);
and U10793 (N_10793,N_8530,N_7858);
nand U10794 (N_10794,N_6248,N_6016);
or U10795 (N_10795,N_7428,N_6678);
or U10796 (N_10796,N_8258,N_6778);
nor U10797 (N_10797,N_8308,N_6682);
nor U10798 (N_10798,N_8384,N_6709);
nor U10799 (N_10799,N_7631,N_6748);
nand U10800 (N_10800,N_6179,N_8558);
nor U10801 (N_10801,N_8160,N_7937);
and U10802 (N_10802,N_6377,N_6903);
xnor U10803 (N_10803,N_6806,N_6836);
nand U10804 (N_10804,N_6802,N_7981);
nand U10805 (N_10805,N_7923,N_6428);
nand U10806 (N_10806,N_8709,N_7331);
and U10807 (N_10807,N_6344,N_7183);
or U10808 (N_10808,N_6428,N_8494);
and U10809 (N_10809,N_6930,N_6484);
and U10810 (N_10810,N_7402,N_6999);
or U10811 (N_10811,N_7321,N_8174);
nand U10812 (N_10812,N_8362,N_7692);
and U10813 (N_10813,N_8940,N_7449);
nand U10814 (N_10814,N_6905,N_7438);
nand U10815 (N_10815,N_8412,N_8243);
and U10816 (N_10816,N_6619,N_6445);
or U10817 (N_10817,N_8804,N_7211);
and U10818 (N_10818,N_6708,N_6014);
nor U10819 (N_10819,N_7142,N_8406);
nor U10820 (N_10820,N_7341,N_8372);
nand U10821 (N_10821,N_8182,N_6983);
nand U10822 (N_10822,N_8482,N_7051);
and U10823 (N_10823,N_7061,N_7211);
nor U10824 (N_10824,N_8772,N_7172);
nor U10825 (N_10825,N_6750,N_7371);
and U10826 (N_10826,N_7324,N_7316);
xnor U10827 (N_10827,N_6460,N_8383);
and U10828 (N_10828,N_8723,N_8614);
nand U10829 (N_10829,N_8761,N_7529);
or U10830 (N_10830,N_7358,N_8222);
nand U10831 (N_10831,N_7041,N_7937);
and U10832 (N_10832,N_7502,N_8095);
or U10833 (N_10833,N_7727,N_8463);
nand U10834 (N_10834,N_8864,N_8894);
xnor U10835 (N_10835,N_8799,N_7291);
nand U10836 (N_10836,N_8745,N_6501);
nand U10837 (N_10837,N_6304,N_8906);
xor U10838 (N_10838,N_7538,N_8747);
xnor U10839 (N_10839,N_8917,N_8765);
xor U10840 (N_10840,N_6499,N_8726);
and U10841 (N_10841,N_6055,N_6395);
xor U10842 (N_10842,N_8981,N_6764);
and U10843 (N_10843,N_8005,N_7069);
and U10844 (N_10844,N_6288,N_8338);
nor U10845 (N_10845,N_8673,N_7874);
nand U10846 (N_10846,N_6212,N_8119);
nand U10847 (N_10847,N_7725,N_7254);
or U10848 (N_10848,N_7334,N_6257);
nor U10849 (N_10849,N_6523,N_8799);
or U10850 (N_10850,N_8533,N_7322);
nor U10851 (N_10851,N_7724,N_7506);
or U10852 (N_10852,N_6546,N_8601);
nor U10853 (N_10853,N_7156,N_7112);
or U10854 (N_10854,N_7504,N_7233);
or U10855 (N_10855,N_7831,N_8963);
or U10856 (N_10856,N_8147,N_6272);
nor U10857 (N_10857,N_6994,N_8469);
nand U10858 (N_10858,N_6353,N_6112);
or U10859 (N_10859,N_7972,N_8085);
nor U10860 (N_10860,N_7903,N_8290);
nand U10861 (N_10861,N_8122,N_6357);
or U10862 (N_10862,N_6804,N_6430);
nand U10863 (N_10863,N_6967,N_8989);
and U10864 (N_10864,N_6078,N_8304);
or U10865 (N_10865,N_6734,N_8598);
xor U10866 (N_10866,N_7587,N_6438);
and U10867 (N_10867,N_6100,N_7715);
nor U10868 (N_10868,N_6663,N_6561);
nand U10869 (N_10869,N_8080,N_8716);
nand U10870 (N_10870,N_7624,N_7292);
nand U10871 (N_10871,N_8177,N_8978);
and U10872 (N_10872,N_7234,N_6970);
xor U10873 (N_10873,N_8956,N_8790);
and U10874 (N_10874,N_8794,N_8415);
nor U10875 (N_10875,N_7077,N_8711);
nand U10876 (N_10876,N_8427,N_8017);
nor U10877 (N_10877,N_7919,N_7846);
nand U10878 (N_10878,N_6379,N_6350);
or U10879 (N_10879,N_7237,N_6342);
or U10880 (N_10880,N_6842,N_6567);
nand U10881 (N_10881,N_7263,N_7917);
and U10882 (N_10882,N_7595,N_7826);
nand U10883 (N_10883,N_8268,N_8256);
xnor U10884 (N_10884,N_7769,N_8288);
nand U10885 (N_10885,N_6763,N_6297);
nand U10886 (N_10886,N_6244,N_7370);
nor U10887 (N_10887,N_6522,N_6702);
or U10888 (N_10888,N_7498,N_6912);
nor U10889 (N_10889,N_6652,N_8340);
and U10890 (N_10890,N_6778,N_7179);
nor U10891 (N_10891,N_7270,N_8344);
and U10892 (N_10892,N_8898,N_8301);
and U10893 (N_10893,N_6440,N_6308);
or U10894 (N_10894,N_7346,N_6468);
nand U10895 (N_10895,N_8975,N_8138);
nand U10896 (N_10896,N_6908,N_8900);
nand U10897 (N_10897,N_7969,N_6173);
and U10898 (N_10898,N_8638,N_6463);
nor U10899 (N_10899,N_6712,N_6893);
and U10900 (N_10900,N_7083,N_8259);
nand U10901 (N_10901,N_6255,N_7034);
or U10902 (N_10902,N_6918,N_7615);
or U10903 (N_10903,N_6637,N_7611);
nor U10904 (N_10904,N_7225,N_7791);
xnor U10905 (N_10905,N_7444,N_6000);
nand U10906 (N_10906,N_6610,N_8843);
nor U10907 (N_10907,N_8726,N_6494);
nor U10908 (N_10908,N_7787,N_8738);
nand U10909 (N_10909,N_6111,N_6495);
or U10910 (N_10910,N_6390,N_7333);
xnor U10911 (N_10911,N_8483,N_7825);
nor U10912 (N_10912,N_6183,N_8792);
nor U10913 (N_10913,N_7888,N_6134);
nor U10914 (N_10914,N_8459,N_7694);
nor U10915 (N_10915,N_7967,N_8081);
and U10916 (N_10916,N_7946,N_8787);
or U10917 (N_10917,N_6365,N_7421);
nor U10918 (N_10918,N_8061,N_8135);
nand U10919 (N_10919,N_7299,N_8348);
nand U10920 (N_10920,N_8667,N_8292);
nand U10921 (N_10921,N_6553,N_6115);
and U10922 (N_10922,N_7275,N_6726);
or U10923 (N_10923,N_6786,N_7542);
or U10924 (N_10924,N_8356,N_8240);
nand U10925 (N_10925,N_8993,N_7474);
nor U10926 (N_10926,N_7357,N_6852);
or U10927 (N_10927,N_7195,N_7329);
or U10928 (N_10928,N_7910,N_6828);
nor U10929 (N_10929,N_7363,N_6837);
nand U10930 (N_10930,N_7595,N_8995);
xor U10931 (N_10931,N_8996,N_6557);
nand U10932 (N_10932,N_7031,N_6504);
nor U10933 (N_10933,N_6296,N_7069);
nor U10934 (N_10934,N_7745,N_6503);
nand U10935 (N_10935,N_6834,N_6385);
nand U10936 (N_10936,N_8852,N_8305);
or U10937 (N_10937,N_8200,N_6565);
nand U10938 (N_10938,N_7206,N_8821);
nand U10939 (N_10939,N_6827,N_8644);
and U10940 (N_10940,N_8294,N_7184);
nand U10941 (N_10941,N_7650,N_8519);
nand U10942 (N_10942,N_6196,N_6761);
nand U10943 (N_10943,N_8395,N_8339);
or U10944 (N_10944,N_6623,N_6039);
nor U10945 (N_10945,N_7302,N_7980);
and U10946 (N_10946,N_7269,N_8098);
nor U10947 (N_10947,N_7558,N_8996);
xor U10948 (N_10948,N_8749,N_6241);
and U10949 (N_10949,N_6551,N_6725);
nand U10950 (N_10950,N_6296,N_7576);
or U10951 (N_10951,N_8930,N_8545);
or U10952 (N_10952,N_6525,N_7651);
xor U10953 (N_10953,N_6928,N_6455);
or U10954 (N_10954,N_8142,N_6432);
or U10955 (N_10955,N_7534,N_8378);
xnor U10956 (N_10956,N_8246,N_8288);
nor U10957 (N_10957,N_7104,N_8015);
or U10958 (N_10958,N_7653,N_8908);
nand U10959 (N_10959,N_8448,N_6871);
nand U10960 (N_10960,N_8357,N_8193);
and U10961 (N_10961,N_7903,N_6497);
or U10962 (N_10962,N_7299,N_8663);
nor U10963 (N_10963,N_7267,N_8253);
nand U10964 (N_10964,N_6967,N_7847);
or U10965 (N_10965,N_8377,N_7917);
nor U10966 (N_10966,N_8604,N_8102);
or U10967 (N_10967,N_6691,N_6009);
nor U10968 (N_10968,N_8452,N_6900);
nand U10969 (N_10969,N_6258,N_6382);
and U10970 (N_10970,N_7811,N_8233);
nor U10971 (N_10971,N_8858,N_7741);
nand U10972 (N_10972,N_6517,N_8128);
nor U10973 (N_10973,N_8521,N_8178);
xnor U10974 (N_10974,N_7299,N_7360);
nand U10975 (N_10975,N_6015,N_8723);
nor U10976 (N_10976,N_8055,N_8445);
nand U10977 (N_10977,N_8432,N_7635);
nor U10978 (N_10978,N_7282,N_8206);
nor U10979 (N_10979,N_7566,N_8146);
nor U10980 (N_10980,N_6784,N_6988);
or U10981 (N_10981,N_8103,N_8586);
or U10982 (N_10982,N_8512,N_8925);
nor U10983 (N_10983,N_7817,N_7262);
or U10984 (N_10984,N_7629,N_6605);
and U10985 (N_10985,N_6562,N_7157);
and U10986 (N_10986,N_7727,N_6031);
and U10987 (N_10987,N_8660,N_8376);
nor U10988 (N_10988,N_7712,N_6749);
nand U10989 (N_10989,N_7519,N_7107);
and U10990 (N_10990,N_7786,N_7430);
xnor U10991 (N_10991,N_7729,N_8686);
nor U10992 (N_10992,N_8512,N_8594);
nor U10993 (N_10993,N_6397,N_7510);
nand U10994 (N_10994,N_6580,N_6394);
or U10995 (N_10995,N_6733,N_7189);
nor U10996 (N_10996,N_7220,N_6057);
or U10997 (N_10997,N_6797,N_7294);
xnor U10998 (N_10998,N_7576,N_8347);
and U10999 (N_10999,N_7097,N_8064);
nor U11000 (N_11000,N_6572,N_8389);
xor U11001 (N_11001,N_8882,N_8286);
nand U11002 (N_11002,N_8331,N_6466);
or U11003 (N_11003,N_8135,N_7049);
nand U11004 (N_11004,N_8871,N_7090);
and U11005 (N_11005,N_6099,N_7559);
or U11006 (N_11006,N_8876,N_6631);
nand U11007 (N_11007,N_7682,N_6150);
nor U11008 (N_11008,N_7959,N_7545);
nand U11009 (N_11009,N_8181,N_6554);
or U11010 (N_11010,N_7260,N_8267);
or U11011 (N_11011,N_6788,N_6070);
nand U11012 (N_11012,N_7869,N_6834);
and U11013 (N_11013,N_7170,N_8166);
and U11014 (N_11014,N_7075,N_6290);
and U11015 (N_11015,N_8851,N_8166);
and U11016 (N_11016,N_8781,N_7902);
and U11017 (N_11017,N_8471,N_7433);
and U11018 (N_11018,N_6461,N_7513);
or U11019 (N_11019,N_7360,N_6531);
nand U11020 (N_11020,N_6209,N_8248);
xnor U11021 (N_11021,N_7257,N_6606);
nand U11022 (N_11022,N_6844,N_8621);
and U11023 (N_11023,N_6473,N_8136);
nor U11024 (N_11024,N_6073,N_8214);
or U11025 (N_11025,N_7362,N_7116);
and U11026 (N_11026,N_6431,N_8528);
nand U11027 (N_11027,N_6150,N_6383);
or U11028 (N_11028,N_6429,N_6593);
nor U11029 (N_11029,N_7996,N_6798);
xnor U11030 (N_11030,N_6153,N_6146);
nor U11031 (N_11031,N_7694,N_8810);
xor U11032 (N_11032,N_6794,N_6237);
and U11033 (N_11033,N_6992,N_8185);
or U11034 (N_11034,N_7408,N_7728);
and U11035 (N_11035,N_8596,N_6947);
and U11036 (N_11036,N_8755,N_6164);
nor U11037 (N_11037,N_6417,N_6639);
or U11038 (N_11038,N_8729,N_7981);
or U11039 (N_11039,N_6739,N_6125);
nand U11040 (N_11040,N_8542,N_7681);
nand U11041 (N_11041,N_7149,N_8641);
or U11042 (N_11042,N_6157,N_6835);
and U11043 (N_11043,N_6169,N_7062);
and U11044 (N_11044,N_6755,N_7185);
or U11045 (N_11045,N_8273,N_7042);
or U11046 (N_11046,N_8868,N_7858);
xor U11047 (N_11047,N_6254,N_6899);
or U11048 (N_11048,N_8321,N_6158);
nand U11049 (N_11049,N_6101,N_7629);
or U11050 (N_11050,N_8977,N_8237);
and U11051 (N_11051,N_7878,N_6526);
nand U11052 (N_11052,N_6564,N_7022);
and U11053 (N_11053,N_8120,N_7226);
nand U11054 (N_11054,N_7843,N_6210);
and U11055 (N_11055,N_6991,N_7585);
nor U11056 (N_11056,N_8742,N_7422);
xnor U11057 (N_11057,N_7049,N_7208);
and U11058 (N_11058,N_8371,N_7747);
nor U11059 (N_11059,N_8719,N_7846);
and U11060 (N_11060,N_8956,N_6861);
nor U11061 (N_11061,N_8061,N_8915);
or U11062 (N_11062,N_7956,N_8624);
nand U11063 (N_11063,N_8744,N_7868);
nor U11064 (N_11064,N_8897,N_7930);
xnor U11065 (N_11065,N_6295,N_6051);
nand U11066 (N_11066,N_7949,N_8314);
nor U11067 (N_11067,N_6685,N_7434);
and U11068 (N_11068,N_6158,N_7360);
or U11069 (N_11069,N_7564,N_6599);
nor U11070 (N_11070,N_6828,N_8719);
nor U11071 (N_11071,N_7980,N_6513);
xnor U11072 (N_11072,N_8247,N_7344);
and U11073 (N_11073,N_6279,N_6164);
nor U11074 (N_11074,N_6673,N_6586);
or U11075 (N_11075,N_6778,N_6983);
or U11076 (N_11076,N_6314,N_8456);
nand U11077 (N_11077,N_7076,N_7227);
or U11078 (N_11078,N_8408,N_7510);
xor U11079 (N_11079,N_7698,N_6443);
and U11080 (N_11080,N_8758,N_7118);
or U11081 (N_11081,N_7810,N_7877);
nor U11082 (N_11082,N_8469,N_7746);
nor U11083 (N_11083,N_8966,N_8875);
or U11084 (N_11084,N_7780,N_6236);
and U11085 (N_11085,N_8140,N_7247);
xor U11086 (N_11086,N_8385,N_6310);
nor U11087 (N_11087,N_7468,N_6356);
and U11088 (N_11088,N_7567,N_8636);
xor U11089 (N_11089,N_7461,N_6712);
nor U11090 (N_11090,N_8565,N_7879);
nand U11091 (N_11091,N_8365,N_7694);
and U11092 (N_11092,N_8643,N_8143);
nand U11093 (N_11093,N_8850,N_8347);
and U11094 (N_11094,N_7468,N_7668);
and U11095 (N_11095,N_6331,N_8297);
nor U11096 (N_11096,N_8751,N_8737);
xor U11097 (N_11097,N_7018,N_8550);
nand U11098 (N_11098,N_6206,N_7424);
and U11099 (N_11099,N_7420,N_7718);
nor U11100 (N_11100,N_8377,N_7513);
nand U11101 (N_11101,N_7322,N_7723);
nor U11102 (N_11102,N_6432,N_7811);
nor U11103 (N_11103,N_6166,N_8493);
nor U11104 (N_11104,N_8464,N_7598);
nand U11105 (N_11105,N_6934,N_6076);
or U11106 (N_11106,N_6590,N_6094);
nor U11107 (N_11107,N_7082,N_7778);
nor U11108 (N_11108,N_6787,N_7623);
and U11109 (N_11109,N_7575,N_7433);
and U11110 (N_11110,N_6953,N_6772);
nand U11111 (N_11111,N_8930,N_6000);
xnor U11112 (N_11112,N_6653,N_8582);
nand U11113 (N_11113,N_7684,N_7118);
or U11114 (N_11114,N_8894,N_6209);
nor U11115 (N_11115,N_8910,N_7510);
nand U11116 (N_11116,N_7997,N_6180);
nor U11117 (N_11117,N_7694,N_7756);
xnor U11118 (N_11118,N_6464,N_6863);
nor U11119 (N_11119,N_7965,N_7423);
and U11120 (N_11120,N_8899,N_6528);
xnor U11121 (N_11121,N_6845,N_7128);
and U11122 (N_11122,N_6418,N_7270);
and U11123 (N_11123,N_8336,N_6835);
xor U11124 (N_11124,N_6724,N_8885);
and U11125 (N_11125,N_6706,N_7289);
and U11126 (N_11126,N_6276,N_8603);
nor U11127 (N_11127,N_7211,N_7069);
or U11128 (N_11128,N_8287,N_8617);
xor U11129 (N_11129,N_7906,N_8733);
or U11130 (N_11130,N_8665,N_7839);
and U11131 (N_11131,N_8302,N_7405);
or U11132 (N_11132,N_6822,N_7366);
or U11133 (N_11133,N_7896,N_6385);
and U11134 (N_11134,N_7683,N_7090);
nor U11135 (N_11135,N_6464,N_8058);
nor U11136 (N_11136,N_8275,N_7103);
nand U11137 (N_11137,N_6851,N_8791);
and U11138 (N_11138,N_6721,N_7397);
or U11139 (N_11139,N_7927,N_7064);
and U11140 (N_11140,N_8055,N_6627);
nand U11141 (N_11141,N_7994,N_8144);
nor U11142 (N_11142,N_6295,N_6533);
nand U11143 (N_11143,N_7019,N_6342);
nand U11144 (N_11144,N_6279,N_7961);
nor U11145 (N_11145,N_8215,N_7255);
xnor U11146 (N_11146,N_8636,N_6979);
nand U11147 (N_11147,N_8567,N_8631);
nand U11148 (N_11148,N_7922,N_7679);
and U11149 (N_11149,N_8827,N_7064);
nor U11150 (N_11150,N_7258,N_8201);
and U11151 (N_11151,N_8492,N_8351);
or U11152 (N_11152,N_8788,N_8331);
xor U11153 (N_11153,N_6958,N_7059);
nand U11154 (N_11154,N_8626,N_7168);
nor U11155 (N_11155,N_6561,N_8571);
nand U11156 (N_11156,N_7407,N_7808);
and U11157 (N_11157,N_7099,N_8488);
or U11158 (N_11158,N_7711,N_8685);
nand U11159 (N_11159,N_8355,N_6144);
and U11160 (N_11160,N_7485,N_8298);
xor U11161 (N_11161,N_8931,N_8512);
or U11162 (N_11162,N_8280,N_6354);
nor U11163 (N_11163,N_7648,N_8190);
and U11164 (N_11164,N_7013,N_6366);
xnor U11165 (N_11165,N_6937,N_7340);
nand U11166 (N_11166,N_6705,N_7648);
and U11167 (N_11167,N_6780,N_6665);
and U11168 (N_11168,N_6166,N_7844);
or U11169 (N_11169,N_6195,N_6326);
and U11170 (N_11170,N_8481,N_6658);
xnor U11171 (N_11171,N_7797,N_7354);
nand U11172 (N_11172,N_6086,N_7481);
and U11173 (N_11173,N_7783,N_7137);
nor U11174 (N_11174,N_7965,N_7757);
nand U11175 (N_11175,N_7305,N_8828);
and U11176 (N_11176,N_6858,N_7939);
or U11177 (N_11177,N_8270,N_8236);
and U11178 (N_11178,N_6811,N_6868);
or U11179 (N_11179,N_6948,N_8138);
xor U11180 (N_11180,N_7651,N_6906);
and U11181 (N_11181,N_8570,N_6511);
or U11182 (N_11182,N_8063,N_7540);
nand U11183 (N_11183,N_7217,N_7308);
or U11184 (N_11184,N_7806,N_6354);
and U11185 (N_11185,N_8452,N_8528);
nand U11186 (N_11186,N_6334,N_7046);
nor U11187 (N_11187,N_7758,N_6600);
nand U11188 (N_11188,N_6909,N_6602);
xnor U11189 (N_11189,N_8290,N_7066);
nand U11190 (N_11190,N_8021,N_8497);
and U11191 (N_11191,N_8336,N_7868);
or U11192 (N_11192,N_6248,N_7721);
nor U11193 (N_11193,N_7849,N_6310);
and U11194 (N_11194,N_6944,N_8036);
and U11195 (N_11195,N_7505,N_6016);
or U11196 (N_11196,N_8263,N_7531);
xor U11197 (N_11197,N_6092,N_8483);
nand U11198 (N_11198,N_7846,N_8080);
xnor U11199 (N_11199,N_6252,N_7249);
and U11200 (N_11200,N_8101,N_8955);
nand U11201 (N_11201,N_6782,N_7938);
nor U11202 (N_11202,N_7590,N_8100);
nand U11203 (N_11203,N_8367,N_6494);
nand U11204 (N_11204,N_7390,N_6846);
nor U11205 (N_11205,N_7202,N_7834);
nor U11206 (N_11206,N_6534,N_8092);
nand U11207 (N_11207,N_6566,N_8565);
nor U11208 (N_11208,N_6653,N_8763);
nand U11209 (N_11209,N_7999,N_7455);
or U11210 (N_11210,N_7234,N_8619);
and U11211 (N_11211,N_8681,N_8952);
nor U11212 (N_11212,N_6781,N_8612);
or U11213 (N_11213,N_6489,N_8949);
nor U11214 (N_11214,N_6759,N_8411);
or U11215 (N_11215,N_6360,N_8145);
and U11216 (N_11216,N_8728,N_6741);
and U11217 (N_11217,N_6602,N_6328);
nand U11218 (N_11218,N_6913,N_6431);
or U11219 (N_11219,N_7423,N_6421);
xnor U11220 (N_11220,N_7923,N_8410);
or U11221 (N_11221,N_6565,N_6376);
nand U11222 (N_11222,N_8630,N_8667);
nand U11223 (N_11223,N_6601,N_8519);
and U11224 (N_11224,N_7288,N_6656);
nor U11225 (N_11225,N_6242,N_7502);
nor U11226 (N_11226,N_6959,N_8167);
and U11227 (N_11227,N_6125,N_8763);
nand U11228 (N_11228,N_6049,N_8586);
and U11229 (N_11229,N_6929,N_7629);
nand U11230 (N_11230,N_8031,N_6286);
or U11231 (N_11231,N_8763,N_7789);
and U11232 (N_11232,N_7352,N_7102);
and U11233 (N_11233,N_6815,N_6338);
nand U11234 (N_11234,N_6059,N_8330);
or U11235 (N_11235,N_6903,N_6239);
nor U11236 (N_11236,N_7697,N_6232);
nor U11237 (N_11237,N_8038,N_7710);
or U11238 (N_11238,N_8247,N_6038);
nand U11239 (N_11239,N_6093,N_8286);
nand U11240 (N_11240,N_7553,N_6042);
or U11241 (N_11241,N_7174,N_7374);
nor U11242 (N_11242,N_6612,N_7328);
nor U11243 (N_11243,N_8457,N_8973);
and U11244 (N_11244,N_8693,N_8265);
nor U11245 (N_11245,N_7223,N_8510);
or U11246 (N_11246,N_7830,N_7998);
nor U11247 (N_11247,N_8315,N_8353);
or U11248 (N_11248,N_6578,N_7944);
nor U11249 (N_11249,N_6274,N_6684);
and U11250 (N_11250,N_8119,N_6275);
nand U11251 (N_11251,N_8923,N_8045);
and U11252 (N_11252,N_8807,N_8356);
or U11253 (N_11253,N_7454,N_6716);
or U11254 (N_11254,N_7188,N_6134);
or U11255 (N_11255,N_6406,N_6284);
and U11256 (N_11256,N_7439,N_6137);
or U11257 (N_11257,N_7559,N_8734);
or U11258 (N_11258,N_6870,N_6651);
nor U11259 (N_11259,N_7770,N_8828);
nand U11260 (N_11260,N_6364,N_7766);
nor U11261 (N_11261,N_8155,N_7458);
nor U11262 (N_11262,N_7299,N_7592);
nand U11263 (N_11263,N_6229,N_8966);
nand U11264 (N_11264,N_6689,N_7932);
and U11265 (N_11265,N_7288,N_7555);
or U11266 (N_11266,N_8692,N_8417);
and U11267 (N_11267,N_6438,N_8935);
nand U11268 (N_11268,N_7563,N_6591);
nor U11269 (N_11269,N_6577,N_6506);
nor U11270 (N_11270,N_7503,N_7109);
nor U11271 (N_11271,N_6176,N_6322);
nor U11272 (N_11272,N_8487,N_8370);
or U11273 (N_11273,N_7459,N_6948);
or U11274 (N_11274,N_7170,N_6633);
and U11275 (N_11275,N_7409,N_7024);
and U11276 (N_11276,N_6823,N_8983);
xor U11277 (N_11277,N_7501,N_7194);
or U11278 (N_11278,N_7632,N_7185);
and U11279 (N_11279,N_6596,N_6229);
or U11280 (N_11280,N_6727,N_7399);
and U11281 (N_11281,N_7853,N_8882);
or U11282 (N_11282,N_6625,N_7177);
or U11283 (N_11283,N_8287,N_6088);
nand U11284 (N_11284,N_7745,N_8465);
nor U11285 (N_11285,N_8759,N_6665);
nand U11286 (N_11286,N_8602,N_7569);
nor U11287 (N_11287,N_8803,N_7890);
nor U11288 (N_11288,N_8272,N_8651);
and U11289 (N_11289,N_7338,N_8243);
nand U11290 (N_11290,N_6016,N_6011);
nor U11291 (N_11291,N_8306,N_8128);
nand U11292 (N_11292,N_6330,N_7738);
nand U11293 (N_11293,N_7638,N_6192);
and U11294 (N_11294,N_8282,N_7342);
nor U11295 (N_11295,N_8516,N_7230);
or U11296 (N_11296,N_6370,N_8911);
and U11297 (N_11297,N_7476,N_6219);
and U11298 (N_11298,N_6534,N_7251);
nor U11299 (N_11299,N_6504,N_8018);
or U11300 (N_11300,N_7906,N_6906);
nand U11301 (N_11301,N_8045,N_6200);
or U11302 (N_11302,N_6019,N_7096);
nor U11303 (N_11303,N_7379,N_6912);
nand U11304 (N_11304,N_8085,N_6673);
and U11305 (N_11305,N_6237,N_7184);
or U11306 (N_11306,N_7962,N_6665);
or U11307 (N_11307,N_6990,N_7150);
nor U11308 (N_11308,N_8607,N_6845);
nor U11309 (N_11309,N_8828,N_6490);
and U11310 (N_11310,N_7345,N_8933);
nand U11311 (N_11311,N_8692,N_7787);
and U11312 (N_11312,N_7495,N_7043);
nor U11313 (N_11313,N_7259,N_7229);
and U11314 (N_11314,N_7076,N_6639);
nor U11315 (N_11315,N_6540,N_7943);
xor U11316 (N_11316,N_8588,N_6810);
and U11317 (N_11317,N_7848,N_7961);
or U11318 (N_11318,N_8769,N_6631);
and U11319 (N_11319,N_8508,N_8673);
nor U11320 (N_11320,N_8191,N_8199);
or U11321 (N_11321,N_7099,N_6270);
xor U11322 (N_11322,N_7162,N_8306);
or U11323 (N_11323,N_8618,N_7781);
nand U11324 (N_11324,N_6264,N_7529);
nor U11325 (N_11325,N_7902,N_7104);
and U11326 (N_11326,N_8256,N_6976);
and U11327 (N_11327,N_8562,N_8174);
and U11328 (N_11328,N_6049,N_8877);
nor U11329 (N_11329,N_8328,N_7269);
or U11330 (N_11330,N_8262,N_8060);
and U11331 (N_11331,N_7460,N_6471);
xnor U11332 (N_11332,N_7746,N_6569);
nand U11333 (N_11333,N_6686,N_7840);
nor U11334 (N_11334,N_6827,N_6514);
nand U11335 (N_11335,N_7799,N_8058);
nand U11336 (N_11336,N_6036,N_6847);
nand U11337 (N_11337,N_7437,N_6431);
xor U11338 (N_11338,N_6890,N_8264);
xor U11339 (N_11339,N_6933,N_8784);
nor U11340 (N_11340,N_6591,N_7400);
or U11341 (N_11341,N_6349,N_8691);
nor U11342 (N_11342,N_8784,N_6369);
or U11343 (N_11343,N_8964,N_6711);
or U11344 (N_11344,N_7811,N_6763);
or U11345 (N_11345,N_6740,N_6601);
and U11346 (N_11346,N_6569,N_7226);
nor U11347 (N_11347,N_7646,N_8378);
nor U11348 (N_11348,N_7768,N_6024);
nand U11349 (N_11349,N_6110,N_6297);
nand U11350 (N_11350,N_8292,N_8555);
nor U11351 (N_11351,N_6829,N_8673);
and U11352 (N_11352,N_8560,N_7142);
nor U11353 (N_11353,N_8105,N_6847);
and U11354 (N_11354,N_8325,N_8843);
nor U11355 (N_11355,N_8146,N_8296);
nor U11356 (N_11356,N_8372,N_7194);
or U11357 (N_11357,N_6529,N_6905);
or U11358 (N_11358,N_6175,N_7935);
xnor U11359 (N_11359,N_7600,N_6333);
xor U11360 (N_11360,N_7040,N_6409);
or U11361 (N_11361,N_6547,N_6053);
or U11362 (N_11362,N_7103,N_7393);
or U11363 (N_11363,N_6087,N_8530);
and U11364 (N_11364,N_6644,N_7184);
nand U11365 (N_11365,N_6254,N_6817);
nor U11366 (N_11366,N_8983,N_8150);
or U11367 (N_11367,N_7562,N_7339);
or U11368 (N_11368,N_8257,N_8705);
nand U11369 (N_11369,N_7063,N_6125);
xor U11370 (N_11370,N_8189,N_8464);
or U11371 (N_11371,N_6294,N_7486);
or U11372 (N_11372,N_7787,N_6952);
nor U11373 (N_11373,N_6194,N_7643);
and U11374 (N_11374,N_8000,N_7372);
nor U11375 (N_11375,N_6872,N_6115);
nand U11376 (N_11376,N_7333,N_6739);
nand U11377 (N_11377,N_6402,N_7579);
and U11378 (N_11378,N_6219,N_7701);
and U11379 (N_11379,N_7532,N_7473);
nor U11380 (N_11380,N_6105,N_7744);
or U11381 (N_11381,N_7776,N_7140);
nor U11382 (N_11382,N_7604,N_8079);
or U11383 (N_11383,N_7753,N_7049);
or U11384 (N_11384,N_8469,N_6074);
and U11385 (N_11385,N_7279,N_8907);
or U11386 (N_11386,N_6598,N_6375);
or U11387 (N_11387,N_8610,N_7957);
nand U11388 (N_11388,N_8113,N_6864);
or U11389 (N_11389,N_7345,N_7567);
nor U11390 (N_11390,N_8086,N_6900);
and U11391 (N_11391,N_7161,N_8158);
xor U11392 (N_11392,N_8182,N_7466);
and U11393 (N_11393,N_8033,N_8447);
xnor U11394 (N_11394,N_6161,N_8719);
nor U11395 (N_11395,N_8773,N_8322);
nor U11396 (N_11396,N_7589,N_7048);
nor U11397 (N_11397,N_7841,N_7715);
nor U11398 (N_11398,N_6834,N_7148);
nand U11399 (N_11399,N_7390,N_8181);
nor U11400 (N_11400,N_8375,N_6309);
and U11401 (N_11401,N_6525,N_7295);
and U11402 (N_11402,N_8117,N_7392);
nand U11403 (N_11403,N_6302,N_7069);
or U11404 (N_11404,N_6783,N_7142);
nor U11405 (N_11405,N_7221,N_8933);
and U11406 (N_11406,N_7380,N_8104);
and U11407 (N_11407,N_6381,N_7331);
xor U11408 (N_11408,N_6988,N_6453);
nor U11409 (N_11409,N_6952,N_7770);
nand U11410 (N_11410,N_8235,N_7992);
or U11411 (N_11411,N_7809,N_6973);
and U11412 (N_11412,N_8469,N_7604);
xor U11413 (N_11413,N_8039,N_7034);
and U11414 (N_11414,N_6222,N_7239);
nand U11415 (N_11415,N_6363,N_6574);
xor U11416 (N_11416,N_6060,N_6349);
or U11417 (N_11417,N_8730,N_6760);
and U11418 (N_11418,N_6384,N_6067);
and U11419 (N_11419,N_7828,N_6812);
nor U11420 (N_11420,N_6623,N_7378);
and U11421 (N_11421,N_7084,N_7489);
nor U11422 (N_11422,N_6682,N_8214);
or U11423 (N_11423,N_7755,N_7365);
xnor U11424 (N_11424,N_7933,N_6929);
and U11425 (N_11425,N_7722,N_6936);
nand U11426 (N_11426,N_8920,N_7041);
xor U11427 (N_11427,N_8835,N_6431);
and U11428 (N_11428,N_8386,N_8989);
nand U11429 (N_11429,N_6996,N_6062);
and U11430 (N_11430,N_8234,N_8438);
nor U11431 (N_11431,N_6718,N_6533);
or U11432 (N_11432,N_6518,N_8264);
and U11433 (N_11433,N_8728,N_8634);
or U11434 (N_11434,N_8172,N_7419);
nand U11435 (N_11435,N_7289,N_7437);
nand U11436 (N_11436,N_6023,N_6778);
and U11437 (N_11437,N_8674,N_7338);
nand U11438 (N_11438,N_6086,N_7759);
and U11439 (N_11439,N_7915,N_8743);
xor U11440 (N_11440,N_6463,N_7547);
xor U11441 (N_11441,N_7782,N_7695);
and U11442 (N_11442,N_8925,N_8240);
and U11443 (N_11443,N_8807,N_8399);
nor U11444 (N_11444,N_6378,N_8063);
nor U11445 (N_11445,N_8312,N_6244);
nand U11446 (N_11446,N_6315,N_6959);
and U11447 (N_11447,N_8585,N_8071);
or U11448 (N_11448,N_8019,N_7268);
and U11449 (N_11449,N_6461,N_8614);
nor U11450 (N_11450,N_7081,N_7777);
nand U11451 (N_11451,N_6459,N_7061);
nand U11452 (N_11452,N_8567,N_7139);
or U11453 (N_11453,N_6199,N_6808);
or U11454 (N_11454,N_8603,N_8796);
or U11455 (N_11455,N_7708,N_8769);
nand U11456 (N_11456,N_6767,N_6966);
nor U11457 (N_11457,N_7725,N_6778);
xnor U11458 (N_11458,N_8967,N_8264);
and U11459 (N_11459,N_8542,N_7335);
nand U11460 (N_11460,N_6223,N_7516);
and U11461 (N_11461,N_7813,N_8080);
nor U11462 (N_11462,N_7017,N_6348);
nand U11463 (N_11463,N_8839,N_7324);
xor U11464 (N_11464,N_6293,N_6592);
nand U11465 (N_11465,N_7445,N_8241);
xor U11466 (N_11466,N_8875,N_6200);
and U11467 (N_11467,N_6052,N_8414);
and U11468 (N_11468,N_6014,N_7899);
nand U11469 (N_11469,N_8361,N_7594);
nand U11470 (N_11470,N_7657,N_8864);
xnor U11471 (N_11471,N_8613,N_8410);
and U11472 (N_11472,N_6709,N_7635);
nand U11473 (N_11473,N_7653,N_6501);
nor U11474 (N_11474,N_6560,N_6946);
nand U11475 (N_11475,N_8789,N_8107);
nor U11476 (N_11476,N_7466,N_8707);
xnor U11477 (N_11477,N_6427,N_6974);
nand U11478 (N_11478,N_6719,N_6417);
or U11479 (N_11479,N_8485,N_7828);
nand U11480 (N_11480,N_6265,N_6517);
and U11481 (N_11481,N_7852,N_8756);
or U11482 (N_11482,N_6136,N_6579);
and U11483 (N_11483,N_8302,N_6016);
and U11484 (N_11484,N_6815,N_6929);
and U11485 (N_11485,N_6143,N_8130);
nand U11486 (N_11486,N_7339,N_8861);
nand U11487 (N_11487,N_7765,N_6263);
xor U11488 (N_11488,N_7396,N_7891);
nor U11489 (N_11489,N_6947,N_6056);
xor U11490 (N_11490,N_6332,N_7809);
nor U11491 (N_11491,N_6564,N_6143);
xnor U11492 (N_11492,N_6742,N_7312);
xnor U11493 (N_11493,N_6726,N_6319);
and U11494 (N_11494,N_6984,N_8808);
or U11495 (N_11495,N_8127,N_6004);
and U11496 (N_11496,N_8364,N_6712);
or U11497 (N_11497,N_7944,N_8776);
nand U11498 (N_11498,N_6464,N_6924);
and U11499 (N_11499,N_6662,N_6398);
or U11500 (N_11500,N_6278,N_8109);
nand U11501 (N_11501,N_7288,N_8093);
or U11502 (N_11502,N_7326,N_6936);
and U11503 (N_11503,N_6003,N_6970);
or U11504 (N_11504,N_8467,N_8881);
nand U11505 (N_11505,N_6517,N_7262);
or U11506 (N_11506,N_8326,N_8045);
or U11507 (N_11507,N_6147,N_8261);
nand U11508 (N_11508,N_8754,N_6092);
nand U11509 (N_11509,N_7663,N_7830);
nor U11510 (N_11510,N_7415,N_7949);
and U11511 (N_11511,N_7786,N_6430);
nand U11512 (N_11512,N_7260,N_6397);
xor U11513 (N_11513,N_8055,N_8017);
nand U11514 (N_11514,N_7920,N_8465);
xor U11515 (N_11515,N_7296,N_7180);
and U11516 (N_11516,N_8207,N_6914);
nor U11517 (N_11517,N_7627,N_7837);
nand U11518 (N_11518,N_7935,N_8804);
and U11519 (N_11519,N_8005,N_8421);
or U11520 (N_11520,N_7002,N_7270);
nand U11521 (N_11521,N_6572,N_6680);
nand U11522 (N_11522,N_7907,N_6002);
or U11523 (N_11523,N_6829,N_7364);
xor U11524 (N_11524,N_6671,N_6650);
or U11525 (N_11525,N_8200,N_7171);
and U11526 (N_11526,N_8168,N_8528);
and U11527 (N_11527,N_6655,N_8068);
xor U11528 (N_11528,N_8768,N_7964);
or U11529 (N_11529,N_7773,N_6204);
xor U11530 (N_11530,N_8137,N_8119);
or U11531 (N_11531,N_8231,N_8977);
and U11532 (N_11532,N_7746,N_7895);
and U11533 (N_11533,N_8639,N_6231);
nand U11534 (N_11534,N_6790,N_7926);
and U11535 (N_11535,N_8597,N_8216);
and U11536 (N_11536,N_8866,N_8357);
and U11537 (N_11537,N_8192,N_8341);
nor U11538 (N_11538,N_7060,N_7487);
nor U11539 (N_11539,N_6608,N_6348);
nor U11540 (N_11540,N_7951,N_6605);
nor U11541 (N_11541,N_7131,N_8848);
nand U11542 (N_11542,N_8022,N_6737);
or U11543 (N_11543,N_6828,N_6369);
nand U11544 (N_11544,N_8497,N_7575);
and U11545 (N_11545,N_6385,N_7753);
or U11546 (N_11546,N_6185,N_6417);
or U11547 (N_11547,N_6664,N_7711);
xnor U11548 (N_11548,N_8412,N_6245);
xnor U11549 (N_11549,N_8088,N_7549);
and U11550 (N_11550,N_7426,N_8346);
and U11551 (N_11551,N_6604,N_7669);
nand U11552 (N_11552,N_6008,N_6751);
xor U11553 (N_11553,N_6219,N_6441);
or U11554 (N_11554,N_6482,N_8583);
or U11555 (N_11555,N_7914,N_8840);
nand U11556 (N_11556,N_8735,N_7078);
xnor U11557 (N_11557,N_6858,N_7656);
and U11558 (N_11558,N_6109,N_6876);
nor U11559 (N_11559,N_6534,N_6131);
xnor U11560 (N_11560,N_6872,N_7338);
or U11561 (N_11561,N_7658,N_6093);
nor U11562 (N_11562,N_8561,N_6333);
and U11563 (N_11563,N_6143,N_7795);
xnor U11564 (N_11564,N_6800,N_6207);
and U11565 (N_11565,N_7549,N_6773);
nor U11566 (N_11566,N_7376,N_6985);
or U11567 (N_11567,N_6886,N_8853);
or U11568 (N_11568,N_8378,N_8598);
nor U11569 (N_11569,N_6973,N_7495);
nor U11570 (N_11570,N_6942,N_6795);
and U11571 (N_11571,N_6912,N_6432);
xor U11572 (N_11572,N_6933,N_6741);
nand U11573 (N_11573,N_8874,N_6977);
nor U11574 (N_11574,N_8427,N_8253);
or U11575 (N_11575,N_8019,N_7190);
nand U11576 (N_11576,N_6501,N_6374);
or U11577 (N_11577,N_7211,N_6146);
xnor U11578 (N_11578,N_7316,N_6367);
and U11579 (N_11579,N_8346,N_6353);
and U11580 (N_11580,N_8350,N_7834);
xnor U11581 (N_11581,N_6274,N_6722);
xnor U11582 (N_11582,N_7623,N_7381);
nor U11583 (N_11583,N_8529,N_7837);
or U11584 (N_11584,N_6048,N_7243);
or U11585 (N_11585,N_6788,N_6418);
nand U11586 (N_11586,N_6092,N_6134);
or U11587 (N_11587,N_6462,N_8876);
or U11588 (N_11588,N_7742,N_8154);
or U11589 (N_11589,N_8139,N_7382);
xnor U11590 (N_11590,N_7955,N_6679);
or U11591 (N_11591,N_6791,N_6875);
and U11592 (N_11592,N_6555,N_7965);
and U11593 (N_11593,N_6337,N_7790);
nand U11594 (N_11594,N_7334,N_8980);
and U11595 (N_11595,N_8465,N_8733);
or U11596 (N_11596,N_6948,N_6866);
and U11597 (N_11597,N_8548,N_8454);
or U11598 (N_11598,N_8607,N_8514);
nand U11599 (N_11599,N_7360,N_7285);
or U11600 (N_11600,N_8584,N_6346);
nand U11601 (N_11601,N_7596,N_7311);
and U11602 (N_11602,N_8454,N_8266);
xnor U11603 (N_11603,N_7623,N_7222);
and U11604 (N_11604,N_7351,N_7702);
and U11605 (N_11605,N_8319,N_8036);
and U11606 (N_11606,N_7897,N_7301);
or U11607 (N_11607,N_6633,N_7957);
and U11608 (N_11608,N_7364,N_6223);
and U11609 (N_11609,N_7621,N_8567);
or U11610 (N_11610,N_8478,N_7734);
xnor U11611 (N_11611,N_8957,N_6536);
nand U11612 (N_11612,N_6645,N_6340);
xor U11613 (N_11613,N_8648,N_7387);
and U11614 (N_11614,N_6656,N_7476);
and U11615 (N_11615,N_6740,N_6817);
and U11616 (N_11616,N_8436,N_6738);
and U11617 (N_11617,N_8587,N_6293);
or U11618 (N_11618,N_6624,N_6313);
nor U11619 (N_11619,N_8772,N_8507);
and U11620 (N_11620,N_8195,N_7480);
nor U11621 (N_11621,N_8695,N_7522);
or U11622 (N_11622,N_7084,N_6161);
or U11623 (N_11623,N_7268,N_8856);
or U11624 (N_11624,N_6947,N_6217);
xnor U11625 (N_11625,N_6359,N_6976);
nand U11626 (N_11626,N_8066,N_7988);
nand U11627 (N_11627,N_8520,N_6074);
xnor U11628 (N_11628,N_6705,N_8093);
nand U11629 (N_11629,N_7546,N_8534);
or U11630 (N_11630,N_7507,N_6295);
xnor U11631 (N_11631,N_8838,N_7914);
nor U11632 (N_11632,N_8386,N_8357);
or U11633 (N_11633,N_8573,N_7178);
or U11634 (N_11634,N_8755,N_8018);
or U11635 (N_11635,N_8471,N_7746);
or U11636 (N_11636,N_8776,N_8229);
or U11637 (N_11637,N_7224,N_8462);
or U11638 (N_11638,N_7625,N_8273);
xor U11639 (N_11639,N_8992,N_8244);
and U11640 (N_11640,N_8648,N_7934);
nand U11641 (N_11641,N_7239,N_7716);
xnor U11642 (N_11642,N_6203,N_7429);
xnor U11643 (N_11643,N_8720,N_6595);
nor U11644 (N_11644,N_6445,N_8503);
nand U11645 (N_11645,N_8849,N_6745);
nor U11646 (N_11646,N_7213,N_7876);
nor U11647 (N_11647,N_6561,N_8219);
nand U11648 (N_11648,N_7323,N_7810);
nor U11649 (N_11649,N_6431,N_8352);
nor U11650 (N_11650,N_8859,N_8653);
nor U11651 (N_11651,N_7673,N_7393);
and U11652 (N_11652,N_8864,N_6000);
nand U11653 (N_11653,N_6663,N_8623);
or U11654 (N_11654,N_6138,N_7709);
and U11655 (N_11655,N_6735,N_7468);
xor U11656 (N_11656,N_8871,N_7014);
and U11657 (N_11657,N_7112,N_7487);
and U11658 (N_11658,N_6113,N_7753);
nand U11659 (N_11659,N_7361,N_6625);
and U11660 (N_11660,N_8812,N_8366);
and U11661 (N_11661,N_8824,N_8406);
nor U11662 (N_11662,N_8026,N_7146);
or U11663 (N_11663,N_7259,N_8561);
nand U11664 (N_11664,N_8859,N_6650);
xor U11665 (N_11665,N_7764,N_7753);
nand U11666 (N_11666,N_7447,N_8539);
nor U11667 (N_11667,N_7512,N_6697);
nor U11668 (N_11668,N_6645,N_8214);
nor U11669 (N_11669,N_6706,N_6001);
nor U11670 (N_11670,N_7521,N_8740);
xor U11671 (N_11671,N_7079,N_7353);
and U11672 (N_11672,N_8495,N_8693);
nor U11673 (N_11673,N_8430,N_6693);
and U11674 (N_11674,N_7810,N_8124);
nand U11675 (N_11675,N_7193,N_6915);
or U11676 (N_11676,N_6562,N_6978);
nand U11677 (N_11677,N_6159,N_7352);
nor U11678 (N_11678,N_7136,N_8248);
xnor U11679 (N_11679,N_7576,N_7927);
and U11680 (N_11680,N_7096,N_8274);
nor U11681 (N_11681,N_8868,N_6118);
xor U11682 (N_11682,N_8041,N_8854);
nand U11683 (N_11683,N_7589,N_8891);
and U11684 (N_11684,N_7283,N_6249);
and U11685 (N_11685,N_6845,N_6486);
nor U11686 (N_11686,N_7214,N_7299);
or U11687 (N_11687,N_7948,N_6365);
nor U11688 (N_11688,N_8953,N_6254);
nand U11689 (N_11689,N_6633,N_6707);
nor U11690 (N_11690,N_6819,N_6765);
nand U11691 (N_11691,N_8126,N_8728);
nor U11692 (N_11692,N_8934,N_7657);
or U11693 (N_11693,N_7198,N_7410);
and U11694 (N_11694,N_6746,N_8054);
nor U11695 (N_11695,N_8876,N_8885);
nor U11696 (N_11696,N_7332,N_8166);
or U11697 (N_11697,N_7256,N_6119);
nor U11698 (N_11698,N_6093,N_8268);
and U11699 (N_11699,N_8747,N_7811);
or U11700 (N_11700,N_8668,N_6081);
or U11701 (N_11701,N_8957,N_7849);
nor U11702 (N_11702,N_8978,N_8122);
and U11703 (N_11703,N_6914,N_7743);
nor U11704 (N_11704,N_6647,N_8049);
nand U11705 (N_11705,N_6190,N_6737);
and U11706 (N_11706,N_6903,N_7440);
nor U11707 (N_11707,N_7492,N_8539);
or U11708 (N_11708,N_8646,N_7900);
xor U11709 (N_11709,N_6483,N_8074);
nor U11710 (N_11710,N_7806,N_8109);
or U11711 (N_11711,N_8896,N_8736);
or U11712 (N_11712,N_7241,N_6812);
xnor U11713 (N_11713,N_6287,N_8632);
nor U11714 (N_11714,N_6075,N_8836);
and U11715 (N_11715,N_6371,N_7500);
nand U11716 (N_11716,N_6431,N_6226);
nor U11717 (N_11717,N_7013,N_8836);
nor U11718 (N_11718,N_7599,N_7342);
xor U11719 (N_11719,N_7125,N_7677);
and U11720 (N_11720,N_8432,N_8100);
nand U11721 (N_11721,N_8877,N_7247);
nor U11722 (N_11722,N_8529,N_7517);
nand U11723 (N_11723,N_7570,N_7337);
nand U11724 (N_11724,N_6310,N_6934);
or U11725 (N_11725,N_8183,N_6475);
nor U11726 (N_11726,N_7172,N_6316);
nor U11727 (N_11727,N_6253,N_6215);
and U11728 (N_11728,N_7081,N_6977);
or U11729 (N_11729,N_8620,N_6403);
nor U11730 (N_11730,N_6893,N_7910);
nor U11731 (N_11731,N_7088,N_8572);
nor U11732 (N_11732,N_7821,N_7185);
xor U11733 (N_11733,N_6782,N_7522);
xnor U11734 (N_11734,N_8764,N_6231);
nor U11735 (N_11735,N_7105,N_7108);
nand U11736 (N_11736,N_7194,N_6742);
and U11737 (N_11737,N_8855,N_6377);
xnor U11738 (N_11738,N_8260,N_8376);
and U11739 (N_11739,N_7017,N_6330);
xnor U11740 (N_11740,N_6981,N_6386);
xor U11741 (N_11741,N_7450,N_6274);
and U11742 (N_11742,N_7599,N_6864);
or U11743 (N_11743,N_8773,N_6702);
and U11744 (N_11744,N_8658,N_8836);
or U11745 (N_11745,N_8786,N_7823);
nor U11746 (N_11746,N_6882,N_7326);
nor U11747 (N_11747,N_6515,N_6427);
nand U11748 (N_11748,N_7165,N_6687);
xor U11749 (N_11749,N_8773,N_8231);
nor U11750 (N_11750,N_8049,N_7490);
nand U11751 (N_11751,N_6092,N_6771);
xnor U11752 (N_11752,N_6810,N_6012);
or U11753 (N_11753,N_6122,N_7420);
nand U11754 (N_11754,N_8788,N_6243);
nand U11755 (N_11755,N_8392,N_8942);
xor U11756 (N_11756,N_7821,N_7929);
and U11757 (N_11757,N_7441,N_6262);
or U11758 (N_11758,N_8062,N_6625);
nor U11759 (N_11759,N_7487,N_7260);
nor U11760 (N_11760,N_7744,N_7160);
nand U11761 (N_11761,N_7675,N_7055);
nand U11762 (N_11762,N_8027,N_7645);
xor U11763 (N_11763,N_6192,N_8856);
nor U11764 (N_11764,N_6468,N_7264);
nand U11765 (N_11765,N_8562,N_7340);
or U11766 (N_11766,N_8222,N_6120);
nand U11767 (N_11767,N_7562,N_6099);
and U11768 (N_11768,N_7716,N_6363);
nor U11769 (N_11769,N_7828,N_7019);
or U11770 (N_11770,N_7877,N_8981);
or U11771 (N_11771,N_8946,N_7988);
nor U11772 (N_11772,N_6431,N_7554);
nand U11773 (N_11773,N_8527,N_8849);
xor U11774 (N_11774,N_6669,N_8178);
nand U11775 (N_11775,N_6327,N_7702);
and U11776 (N_11776,N_6464,N_8872);
and U11777 (N_11777,N_6720,N_7332);
nor U11778 (N_11778,N_6617,N_8992);
nand U11779 (N_11779,N_6317,N_8472);
nand U11780 (N_11780,N_8648,N_6345);
nor U11781 (N_11781,N_8156,N_6900);
or U11782 (N_11782,N_6308,N_8314);
nand U11783 (N_11783,N_6557,N_7245);
nor U11784 (N_11784,N_8510,N_7663);
or U11785 (N_11785,N_8286,N_7905);
and U11786 (N_11786,N_8469,N_7298);
nor U11787 (N_11787,N_6773,N_8322);
and U11788 (N_11788,N_6666,N_8092);
or U11789 (N_11789,N_6099,N_7089);
or U11790 (N_11790,N_8613,N_8617);
or U11791 (N_11791,N_7656,N_6126);
or U11792 (N_11792,N_6968,N_8916);
and U11793 (N_11793,N_7125,N_7325);
nand U11794 (N_11794,N_8878,N_6560);
and U11795 (N_11795,N_7407,N_8131);
nand U11796 (N_11796,N_8032,N_7734);
nand U11797 (N_11797,N_8322,N_6746);
or U11798 (N_11798,N_7151,N_7097);
nor U11799 (N_11799,N_7237,N_8997);
xnor U11800 (N_11800,N_7277,N_8256);
nand U11801 (N_11801,N_6380,N_6435);
and U11802 (N_11802,N_6508,N_6029);
or U11803 (N_11803,N_8220,N_7409);
nor U11804 (N_11804,N_6005,N_8553);
nand U11805 (N_11805,N_8279,N_7132);
and U11806 (N_11806,N_6257,N_7057);
or U11807 (N_11807,N_8443,N_6005);
nor U11808 (N_11808,N_6603,N_7503);
and U11809 (N_11809,N_7406,N_7774);
and U11810 (N_11810,N_8379,N_7455);
nand U11811 (N_11811,N_8120,N_6088);
and U11812 (N_11812,N_8105,N_8529);
or U11813 (N_11813,N_6401,N_8548);
or U11814 (N_11814,N_6082,N_7069);
or U11815 (N_11815,N_8399,N_7856);
xor U11816 (N_11816,N_6781,N_6272);
nor U11817 (N_11817,N_6312,N_7710);
nand U11818 (N_11818,N_7207,N_8192);
nand U11819 (N_11819,N_8456,N_6215);
and U11820 (N_11820,N_7389,N_7713);
or U11821 (N_11821,N_8179,N_8165);
nor U11822 (N_11822,N_8947,N_8472);
and U11823 (N_11823,N_8088,N_7807);
nor U11824 (N_11824,N_8130,N_7377);
and U11825 (N_11825,N_6483,N_6443);
nand U11826 (N_11826,N_7854,N_7295);
or U11827 (N_11827,N_8876,N_7822);
nor U11828 (N_11828,N_8592,N_7545);
nand U11829 (N_11829,N_6371,N_8098);
and U11830 (N_11830,N_8446,N_8991);
and U11831 (N_11831,N_8145,N_8414);
or U11832 (N_11832,N_8321,N_8039);
or U11833 (N_11833,N_6507,N_7391);
nand U11834 (N_11834,N_7415,N_7288);
nor U11835 (N_11835,N_8952,N_7853);
nor U11836 (N_11836,N_8198,N_8913);
nor U11837 (N_11837,N_6798,N_8948);
nor U11838 (N_11838,N_7090,N_7933);
nand U11839 (N_11839,N_6075,N_8499);
and U11840 (N_11840,N_6171,N_6297);
xnor U11841 (N_11841,N_8349,N_8654);
nand U11842 (N_11842,N_8827,N_6871);
or U11843 (N_11843,N_6429,N_6340);
nor U11844 (N_11844,N_7944,N_7210);
nor U11845 (N_11845,N_7114,N_6246);
or U11846 (N_11846,N_6767,N_8410);
or U11847 (N_11847,N_8969,N_7835);
nor U11848 (N_11848,N_7017,N_7214);
or U11849 (N_11849,N_8681,N_7070);
nor U11850 (N_11850,N_6375,N_6870);
xnor U11851 (N_11851,N_8981,N_6451);
xnor U11852 (N_11852,N_7744,N_6974);
nor U11853 (N_11853,N_7328,N_6545);
nand U11854 (N_11854,N_8844,N_8333);
and U11855 (N_11855,N_8921,N_7676);
and U11856 (N_11856,N_8445,N_6140);
or U11857 (N_11857,N_7289,N_6459);
nand U11858 (N_11858,N_6437,N_8074);
and U11859 (N_11859,N_8465,N_6361);
nand U11860 (N_11860,N_6769,N_6425);
and U11861 (N_11861,N_8165,N_8232);
xor U11862 (N_11862,N_8879,N_8989);
xor U11863 (N_11863,N_8639,N_8451);
and U11864 (N_11864,N_7249,N_7773);
xnor U11865 (N_11865,N_6316,N_7665);
and U11866 (N_11866,N_8883,N_6381);
and U11867 (N_11867,N_6537,N_8663);
nand U11868 (N_11868,N_6174,N_7463);
and U11869 (N_11869,N_8949,N_7890);
or U11870 (N_11870,N_6267,N_6688);
xnor U11871 (N_11871,N_6186,N_7282);
nand U11872 (N_11872,N_7694,N_8366);
nand U11873 (N_11873,N_6515,N_7883);
or U11874 (N_11874,N_6558,N_7147);
nand U11875 (N_11875,N_8018,N_8566);
and U11876 (N_11876,N_7159,N_7126);
and U11877 (N_11877,N_8466,N_7504);
or U11878 (N_11878,N_7094,N_6029);
nand U11879 (N_11879,N_8476,N_7036);
xnor U11880 (N_11880,N_7418,N_8905);
or U11881 (N_11881,N_6323,N_7809);
xnor U11882 (N_11882,N_8271,N_7870);
nor U11883 (N_11883,N_8109,N_7718);
or U11884 (N_11884,N_8127,N_6071);
nor U11885 (N_11885,N_8185,N_8370);
nor U11886 (N_11886,N_7448,N_6460);
and U11887 (N_11887,N_7502,N_7274);
nor U11888 (N_11888,N_7632,N_8044);
nand U11889 (N_11889,N_6640,N_8459);
and U11890 (N_11890,N_8119,N_6165);
or U11891 (N_11891,N_8624,N_7630);
or U11892 (N_11892,N_7412,N_7550);
nand U11893 (N_11893,N_7783,N_6301);
and U11894 (N_11894,N_8563,N_7356);
nand U11895 (N_11895,N_8252,N_7015);
nor U11896 (N_11896,N_6415,N_7832);
nor U11897 (N_11897,N_7302,N_7635);
nor U11898 (N_11898,N_7012,N_6641);
nand U11899 (N_11899,N_8149,N_8687);
nand U11900 (N_11900,N_6974,N_7666);
nor U11901 (N_11901,N_8204,N_6818);
or U11902 (N_11902,N_6521,N_6099);
or U11903 (N_11903,N_7893,N_7821);
xnor U11904 (N_11904,N_8288,N_6846);
or U11905 (N_11905,N_6701,N_6261);
and U11906 (N_11906,N_8968,N_8452);
nand U11907 (N_11907,N_8723,N_6719);
nor U11908 (N_11908,N_8928,N_7662);
nand U11909 (N_11909,N_8316,N_7433);
nor U11910 (N_11910,N_7817,N_6298);
or U11911 (N_11911,N_7276,N_7481);
nand U11912 (N_11912,N_6615,N_8418);
xnor U11913 (N_11913,N_7891,N_6401);
or U11914 (N_11914,N_7891,N_7958);
xor U11915 (N_11915,N_7339,N_7214);
or U11916 (N_11916,N_6839,N_8514);
and U11917 (N_11917,N_8821,N_6234);
nor U11918 (N_11918,N_8297,N_8767);
nor U11919 (N_11919,N_6496,N_6366);
and U11920 (N_11920,N_8211,N_8769);
nor U11921 (N_11921,N_8214,N_6496);
nand U11922 (N_11922,N_7216,N_6205);
and U11923 (N_11923,N_6404,N_7927);
nand U11924 (N_11924,N_8377,N_8472);
or U11925 (N_11925,N_8395,N_8948);
or U11926 (N_11926,N_7484,N_7289);
nand U11927 (N_11927,N_6479,N_8828);
nor U11928 (N_11928,N_8688,N_8872);
and U11929 (N_11929,N_6115,N_8739);
nand U11930 (N_11930,N_6684,N_7362);
or U11931 (N_11931,N_7672,N_7864);
nor U11932 (N_11932,N_6713,N_6015);
nor U11933 (N_11933,N_6442,N_8943);
nand U11934 (N_11934,N_7319,N_7419);
nand U11935 (N_11935,N_6111,N_8816);
nor U11936 (N_11936,N_6335,N_7125);
and U11937 (N_11937,N_6610,N_7005);
or U11938 (N_11938,N_6492,N_7515);
nand U11939 (N_11939,N_8756,N_7940);
nand U11940 (N_11940,N_8188,N_8606);
and U11941 (N_11941,N_8364,N_7207);
nor U11942 (N_11942,N_8624,N_7252);
or U11943 (N_11943,N_8192,N_7550);
nor U11944 (N_11944,N_8350,N_7295);
nor U11945 (N_11945,N_7925,N_8518);
and U11946 (N_11946,N_6488,N_7324);
and U11947 (N_11947,N_8190,N_7856);
and U11948 (N_11948,N_7190,N_8735);
or U11949 (N_11949,N_7631,N_8999);
or U11950 (N_11950,N_6856,N_7002);
nand U11951 (N_11951,N_8833,N_7187);
or U11952 (N_11952,N_8948,N_8482);
nand U11953 (N_11953,N_7230,N_6921);
and U11954 (N_11954,N_6334,N_8885);
or U11955 (N_11955,N_7681,N_6412);
nor U11956 (N_11956,N_7280,N_6659);
nand U11957 (N_11957,N_8171,N_7629);
nor U11958 (N_11958,N_6088,N_6894);
or U11959 (N_11959,N_6694,N_7362);
nand U11960 (N_11960,N_7542,N_7479);
and U11961 (N_11961,N_7990,N_6862);
or U11962 (N_11962,N_7430,N_7393);
nor U11963 (N_11963,N_7588,N_7555);
nor U11964 (N_11964,N_7574,N_7296);
or U11965 (N_11965,N_7255,N_7198);
nor U11966 (N_11966,N_8370,N_7013);
nand U11967 (N_11967,N_7250,N_8721);
nor U11968 (N_11968,N_7754,N_8457);
xnor U11969 (N_11969,N_6019,N_7109);
xnor U11970 (N_11970,N_6097,N_7378);
nor U11971 (N_11971,N_6483,N_8818);
xnor U11972 (N_11972,N_8041,N_8713);
nand U11973 (N_11973,N_7932,N_6624);
xnor U11974 (N_11974,N_8645,N_8814);
or U11975 (N_11975,N_8084,N_8740);
or U11976 (N_11976,N_8659,N_8756);
nand U11977 (N_11977,N_7791,N_8835);
nand U11978 (N_11978,N_6645,N_8550);
and U11979 (N_11979,N_8912,N_6289);
nand U11980 (N_11980,N_8443,N_8563);
nor U11981 (N_11981,N_8224,N_8409);
and U11982 (N_11982,N_6262,N_7604);
or U11983 (N_11983,N_7131,N_8678);
or U11984 (N_11984,N_7114,N_6532);
nor U11985 (N_11985,N_8685,N_7787);
nor U11986 (N_11986,N_7976,N_8315);
nor U11987 (N_11987,N_8856,N_8849);
and U11988 (N_11988,N_8154,N_7933);
or U11989 (N_11989,N_6480,N_8451);
or U11990 (N_11990,N_6316,N_6500);
xnor U11991 (N_11991,N_6877,N_7832);
or U11992 (N_11992,N_8017,N_7700);
and U11993 (N_11993,N_6894,N_8004);
nand U11994 (N_11994,N_7665,N_6686);
xor U11995 (N_11995,N_6581,N_8593);
xor U11996 (N_11996,N_8765,N_6170);
xor U11997 (N_11997,N_6213,N_8283);
nor U11998 (N_11998,N_6690,N_7714);
or U11999 (N_11999,N_8428,N_7792);
nand U12000 (N_12000,N_11136,N_10888);
and U12001 (N_12001,N_11090,N_9434);
and U12002 (N_12002,N_10406,N_10466);
nor U12003 (N_12003,N_9508,N_10164);
nor U12004 (N_12004,N_9295,N_10831);
or U12005 (N_12005,N_10154,N_10349);
xnor U12006 (N_12006,N_9461,N_11309);
nand U12007 (N_12007,N_11927,N_11495);
nor U12008 (N_12008,N_11909,N_10423);
and U12009 (N_12009,N_10446,N_9006);
nand U12010 (N_12010,N_9813,N_10573);
nor U12011 (N_12011,N_10306,N_9377);
or U12012 (N_12012,N_9633,N_11230);
and U12013 (N_12013,N_11558,N_11698);
or U12014 (N_12014,N_10759,N_9334);
nor U12015 (N_12015,N_10510,N_10687);
or U12016 (N_12016,N_11995,N_11506);
nor U12017 (N_12017,N_11490,N_11646);
or U12018 (N_12018,N_11680,N_10812);
nand U12019 (N_12019,N_10585,N_10444);
nor U12020 (N_12020,N_10201,N_10369);
and U12021 (N_12021,N_9060,N_9206);
nor U12022 (N_12022,N_10742,N_11221);
and U12023 (N_12023,N_9689,N_10161);
nand U12024 (N_12024,N_10608,N_11417);
nand U12025 (N_12025,N_9964,N_11205);
xnor U12026 (N_12026,N_10377,N_11633);
or U12027 (N_12027,N_11093,N_9845);
nand U12028 (N_12028,N_9766,N_10101);
and U12029 (N_12029,N_10633,N_11589);
or U12030 (N_12030,N_9404,N_10326);
or U12031 (N_12031,N_10331,N_9979);
nor U12032 (N_12032,N_10422,N_11605);
nand U12033 (N_12033,N_10179,N_11365);
xnor U12034 (N_12034,N_10288,N_11721);
xnor U12035 (N_12035,N_10231,N_10594);
nor U12036 (N_12036,N_11815,N_11241);
or U12037 (N_12037,N_9215,N_11638);
nor U12038 (N_12038,N_11117,N_10930);
nand U12039 (N_12039,N_10503,N_10455);
or U12040 (N_12040,N_11869,N_10250);
and U12041 (N_12041,N_11462,N_10419);
nand U12042 (N_12042,N_9237,N_9024);
xnor U12043 (N_12043,N_9363,N_10114);
or U12044 (N_12044,N_10512,N_10843);
nor U12045 (N_12045,N_10227,N_10667);
nand U12046 (N_12046,N_10702,N_9829);
and U12047 (N_12047,N_10652,N_10277);
nand U12048 (N_12048,N_9509,N_10710);
and U12049 (N_12049,N_11277,N_9165);
or U12050 (N_12050,N_9659,N_10621);
xnor U12051 (N_12051,N_10494,N_10690);
nand U12052 (N_12052,N_10435,N_10097);
and U12053 (N_12053,N_9588,N_10243);
nand U12054 (N_12054,N_9546,N_10000);
nor U12055 (N_12055,N_11655,N_11162);
nand U12056 (N_12056,N_11038,N_11678);
or U12057 (N_12057,N_9208,N_11318);
or U12058 (N_12058,N_9186,N_10966);
nor U12059 (N_12059,N_9634,N_9138);
nand U12060 (N_12060,N_11897,N_9765);
or U12061 (N_12061,N_10875,N_9364);
nand U12062 (N_12062,N_11240,N_9784);
nand U12063 (N_12063,N_11586,N_10357);
or U12064 (N_12064,N_10763,N_10488);
and U12065 (N_12065,N_10789,N_10213);
xnor U12066 (N_12066,N_9817,N_11046);
nand U12067 (N_12067,N_11849,N_9419);
and U12068 (N_12068,N_9867,N_9712);
and U12069 (N_12069,N_10911,N_9886);
xnor U12070 (N_12070,N_10170,N_10801);
nor U12071 (N_12071,N_11665,N_9604);
nor U12072 (N_12072,N_9852,N_10611);
and U12073 (N_12073,N_9063,N_11320);
nor U12074 (N_12074,N_11986,N_9737);
nand U12075 (N_12075,N_11756,N_10432);
nand U12076 (N_12076,N_10299,N_9500);
or U12077 (N_12077,N_10136,N_11306);
or U12078 (N_12078,N_10648,N_11775);
or U12079 (N_12079,N_9221,N_11045);
and U12080 (N_12080,N_11793,N_11015);
and U12081 (N_12081,N_9438,N_9350);
or U12082 (N_12082,N_10134,N_9565);
or U12083 (N_12083,N_9247,N_10159);
or U12084 (N_12084,N_11585,N_9644);
nor U12085 (N_12085,N_10175,N_10739);
and U12086 (N_12086,N_9581,N_9281);
and U12087 (N_12087,N_11673,N_11156);
or U12088 (N_12088,N_11911,N_9714);
nand U12089 (N_12089,N_11774,N_10701);
and U12090 (N_12090,N_10901,N_11514);
nand U12091 (N_12091,N_10713,N_9445);
nor U12092 (N_12092,N_11223,N_11693);
nor U12093 (N_12093,N_9055,N_9536);
and U12094 (N_12094,N_11537,N_9615);
and U12095 (N_12095,N_11200,N_10669);
nand U12096 (N_12096,N_11860,N_9043);
and U12097 (N_12097,N_11974,N_10246);
nor U12098 (N_12098,N_11294,N_9749);
nand U12099 (N_12099,N_9609,N_10990);
or U12100 (N_12100,N_11456,N_11054);
and U12101 (N_12101,N_10087,N_11044);
nand U12102 (N_12102,N_10526,N_10784);
nand U12103 (N_12103,N_10963,N_11316);
and U12104 (N_12104,N_9480,N_10183);
nand U12105 (N_12105,N_11194,N_11727);
xnor U12106 (N_12106,N_11268,N_9132);
xnor U12107 (N_12107,N_10511,N_11557);
nand U12108 (N_12108,N_10076,N_10480);
nand U12109 (N_12109,N_11576,N_11718);
nor U12110 (N_12110,N_10502,N_11875);
xor U12111 (N_12111,N_9803,N_9345);
nor U12112 (N_12112,N_11000,N_11145);
nor U12113 (N_12113,N_11746,N_9007);
xnor U12114 (N_12114,N_10853,N_11349);
nand U12115 (N_12115,N_10320,N_11425);
nand U12116 (N_12116,N_11778,N_10430);
nor U12117 (N_12117,N_11254,N_10009);
nand U12118 (N_12118,N_9718,N_11766);
xor U12119 (N_12119,N_9904,N_9820);
nor U12120 (N_12120,N_9870,N_10174);
nor U12121 (N_12121,N_9413,N_9527);
or U12122 (N_12122,N_9433,N_9080);
and U12123 (N_12123,N_10537,N_11578);
nor U12124 (N_12124,N_9516,N_11299);
nand U12125 (N_12125,N_9750,N_11526);
nor U12126 (N_12126,N_9626,N_11352);
nor U12127 (N_12127,N_10577,N_10785);
nand U12128 (N_12128,N_9321,N_10885);
nand U12129 (N_12129,N_9760,N_9680);
nor U12130 (N_12130,N_11532,N_10313);
nor U12131 (N_12131,N_10260,N_9592);
nand U12132 (N_12132,N_11438,N_9287);
and U12133 (N_12133,N_9403,N_9435);
or U12134 (N_12134,N_10465,N_9798);
and U12135 (N_12135,N_9943,N_11226);
nand U12136 (N_12136,N_11256,N_10664);
nor U12137 (N_12137,N_11658,N_9601);
nand U12138 (N_12138,N_10947,N_9910);
or U12139 (N_12139,N_10576,N_10056);
nor U12140 (N_12140,N_11685,N_9915);
xor U12141 (N_12141,N_10152,N_11469);
or U12142 (N_12142,N_11828,N_11253);
nand U12143 (N_12143,N_9235,N_9518);
and U12144 (N_12144,N_10881,N_11197);
and U12145 (N_12145,N_11065,N_10807);
xor U12146 (N_12146,N_10327,N_11811);
nor U12147 (N_12147,N_10783,N_11584);
nand U12148 (N_12148,N_11672,N_9980);
nand U12149 (N_12149,N_11058,N_10962);
nor U12150 (N_12150,N_11062,N_11668);
or U12151 (N_12151,N_10378,N_9047);
nor U12152 (N_12152,N_9486,N_10704);
or U12153 (N_12153,N_10469,N_11824);
xor U12154 (N_12154,N_11708,N_10192);
and U12155 (N_12155,N_10113,N_9594);
nor U12156 (N_12156,N_9258,N_10300);
and U12157 (N_12157,N_11738,N_9761);
nor U12158 (N_12158,N_11273,N_11423);
xor U12159 (N_12159,N_9828,N_11939);
xnor U12160 (N_12160,N_10632,N_9277);
nor U12161 (N_12161,N_10041,N_11606);
xnor U12162 (N_12162,N_9203,N_11189);
and U12163 (N_12163,N_10979,N_9802);
nor U12164 (N_12164,N_10043,N_9094);
and U12165 (N_12165,N_11217,N_9387);
xnor U12166 (N_12166,N_9078,N_9693);
and U12167 (N_12167,N_9576,N_11813);
or U12168 (N_12168,N_11920,N_11224);
xor U12169 (N_12169,N_10513,N_9073);
nand U12170 (N_12170,N_11488,N_10971);
and U12171 (N_12171,N_9757,N_9201);
nor U12172 (N_12172,N_11982,N_9960);
nor U12173 (N_12173,N_9847,N_9999);
or U12174 (N_12174,N_9264,N_10359);
or U12175 (N_12175,N_10827,N_9416);
or U12176 (N_12176,N_11998,N_9959);
nand U12177 (N_12177,N_11235,N_11888);
and U12178 (N_12178,N_9195,N_11702);
and U12179 (N_12179,N_10994,N_11288);
or U12180 (N_12180,N_10298,N_10761);
or U12181 (N_12181,N_10956,N_10119);
or U12182 (N_12182,N_11692,N_9294);
nand U12183 (N_12183,N_9139,N_10597);
nand U12184 (N_12184,N_9587,N_9523);
or U12185 (N_12185,N_11843,N_9283);
nor U12186 (N_12186,N_11512,N_11321);
nor U12187 (N_12187,N_10737,N_10389);
and U12188 (N_12188,N_11025,N_11696);
nor U12189 (N_12189,N_11945,N_11121);
nor U12190 (N_12190,N_11402,N_10999);
and U12191 (N_12191,N_9234,N_10339);
nor U12192 (N_12192,N_10766,N_9112);
or U12193 (N_12193,N_9009,N_11498);
nor U12194 (N_12194,N_10651,N_9674);
or U12195 (N_12195,N_9973,N_11150);
nor U12196 (N_12196,N_10137,N_10323);
nor U12197 (N_12197,N_10004,N_9935);
and U12198 (N_12198,N_11543,N_10336);
xnor U12199 (N_12199,N_9767,N_11039);
nand U12200 (N_12200,N_10055,N_11616);
and U12201 (N_12201,N_9746,N_11794);
or U12202 (N_12202,N_10301,N_9412);
and U12203 (N_12203,N_9570,N_11475);
nor U12204 (N_12204,N_9679,N_11394);
or U12205 (N_12205,N_10772,N_10005);
or U12206 (N_12206,N_10547,N_11211);
and U12207 (N_12207,N_9431,N_9781);
nor U12208 (N_12208,N_11149,N_10057);
and U12209 (N_12209,N_11750,N_11639);
or U12210 (N_12210,N_9015,N_11878);
and U12211 (N_12211,N_9447,N_10413);
nor U12212 (N_12212,N_9957,N_10539);
nor U12213 (N_12213,N_9695,N_9968);
and U12214 (N_12214,N_10553,N_10256);
or U12215 (N_12215,N_10921,N_9066);
or U12216 (N_12216,N_9386,N_11546);
nor U12217 (N_12217,N_9623,N_10626);
xnor U12218 (N_12218,N_11356,N_11393);
and U12219 (N_12219,N_10160,N_9183);
and U12220 (N_12220,N_10517,N_9284);
nor U12221 (N_12221,N_9612,N_10720);
and U12222 (N_12222,N_9134,N_9149);
and U12223 (N_12223,N_10204,N_10031);
and U12224 (N_12224,N_11745,N_9918);
nor U12225 (N_12225,N_9809,N_10282);
xnor U12226 (N_12226,N_9953,N_11534);
and U12227 (N_12227,N_10965,N_9544);
nand U12228 (N_12228,N_9929,N_11023);
xor U12229 (N_12229,N_11967,N_9896);
nand U12230 (N_12230,N_11631,N_9358);
or U12231 (N_12231,N_11964,N_10582);
nand U12232 (N_12232,N_11019,N_10679);
and U12233 (N_12233,N_10987,N_10694);
or U12234 (N_12234,N_10437,N_9879);
or U12235 (N_12235,N_10036,N_11012);
nor U12236 (N_12236,N_9975,N_10833);
nand U12237 (N_12237,N_10916,N_10066);
nor U12238 (N_12238,N_11547,N_9299);
or U12239 (N_12239,N_9522,N_11414);
nand U12240 (N_12240,N_9502,N_10354);
nor U12241 (N_12241,N_11077,N_11755);
and U12242 (N_12242,N_9173,N_9187);
nand U12243 (N_12243,N_10989,N_11050);
nand U12244 (N_12244,N_10844,N_9494);
and U12245 (N_12245,N_9641,N_9102);
and U12246 (N_12246,N_11380,N_10208);
and U12247 (N_12247,N_9426,N_11583);
nor U12248 (N_12248,N_11400,N_9843);
nand U12249 (N_12249,N_10123,N_9451);
and U12250 (N_12250,N_11762,N_10670);
or U12251 (N_12251,N_9214,N_9161);
xnor U12252 (N_12252,N_11119,N_10474);
nand U12253 (N_12253,N_10310,N_9643);
xor U12254 (N_12254,N_11203,N_9270);
and U12255 (N_12255,N_10586,N_11823);
or U12256 (N_12256,N_9467,N_11401);
nor U12257 (N_12257,N_10024,N_11305);
and U12258 (N_12258,N_9468,N_10823);
xor U12259 (N_12259,N_10862,N_11190);
or U12260 (N_12260,N_10025,N_10361);
and U12261 (N_12261,N_11097,N_9000);
or U12262 (N_12262,N_10187,N_11724);
or U12263 (N_12263,N_11752,N_11113);
nor U12264 (N_12264,N_11800,N_10333);
or U12265 (N_12265,N_11617,N_10949);
or U12266 (N_12266,N_9901,N_9764);
nor U12267 (N_12267,N_10438,N_11291);
or U12268 (N_12268,N_10809,N_11720);
nand U12269 (N_12269,N_11931,N_9337);
nand U12270 (N_12270,N_9137,N_10360);
nor U12271 (N_12271,N_10490,N_10666);
and U12272 (N_12272,N_10214,N_9889);
nor U12273 (N_12273,N_9857,N_11722);
nor U12274 (N_12274,N_9156,N_9956);
nor U12275 (N_12275,N_9023,N_9231);
nor U12276 (N_12276,N_9150,N_10578);
nand U12277 (N_12277,N_9101,N_10481);
nor U12278 (N_12278,N_11049,N_10927);
and U12279 (N_12279,N_10840,N_10824);
xnor U12280 (N_12280,N_9926,N_11464);
and U12281 (N_12281,N_9721,N_11748);
xor U12282 (N_12282,N_9729,N_11178);
nand U12283 (N_12283,N_10748,N_10524);
nand U12284 (N_12284,N_10064,N_11921);
nand U12285 (N_12285,N_11016,N_9021);
xor U12286 (N_12286,N_9653,N_11031);
and U12287 (N_12287,N_9035,N_11980);
or U12288 (N_12288,N_9177,N_9728);
or U12289 (N_12289,N_10415,N_9367);
and U12290 (N_12290,N_9359,N_11844);
xnor U12291 (N_12291,N_9184,N_9204);
and U12292 (N_12292,N_11172,N_11949);
nor U12293 (N_12293,N_11670,N_11422);
nor U12294 (N_12294,N_9030,N_9562);
nand U12295 (N_12295,N_10506,N_10839);
nor U12296 (N_12296,N_9263,N_11675);
nor U12297 (N_12297,N_11701,N_10755);
or U12298 (N_12298,N_9538,N_10616);
nand U12299 (N_12299,N_11887,N_10902);
or U12300 (N_12300,N_10030,N_9940);
nor U12301 (N_12301,N_11202,N_11826);
and U12302 (N_12302,N_9928,N_10094);
nand U12303 (N_12303,N_10799,N_11032);
or U12304 (N_12304,N_11517,N_10290);
nor U12305 (N_12305,N_11327,N_9869);
nand U12306 (N_12306,N_9984,N_9315);
nand U12307 (N_12307,N_11504,N_11773);
nand U12308 (N_12308,N_11528,N_9630);
or U12309 (N_12309,N_10238,N_11222);
nand U12310 (N_12310,N_9361,N_10708);
nor U12311 (N_12311,N_11199,N_9564);
or U12312 (N_12312,N_10668,N_11102);
nand U12313 (N_12313,N_10443,N_9109);
or U12314 (N_12314,N_11161,N_10796);
nand U12315 (N_12315,N_10905,N_11733);
nand U12316 (N_12316,N_9533,N_11968);
nand U12317 (N_12317,N_9949,N_10428);
or U12318 (N_12318,N_11231,N_10135);
and U12319 (N_12319,N_11225,N_10634);
or U12320 (N_12320,N_9099,N_10845);
or U12321 (N_12321,N_10545,N_11419);
nor U12322 (N_12322,N_11886,N_9477);
and U12323 (N_12323,N_10653,N_11053);
and U12324 (N_12324,N_11148,N_10912);
nand U12325 (N_12325,N_10954,N_10983);
nor U12326 (N_12326,N_9121,N_11452);
or U12327 (N_12327,N_9937,N_11014);
and U12328 (N_12328,N_10207,N_10278);
or U12329 (N_12329,N_9266,N_11919);
and U12330 (N_12330,N_10138,N_9560);
nand U12331 (N_12331,N_11577,N_10491);
and U12332 (N_12332,N_9097,N_11783);
xor U12333 (N_12333,N_10734,N_9705);
nor U12334 (N_12334,N_10452,N_9970);
nor U12335 (N_12335,N_11866,N_9213);
or U12336 (N_12336,N_10731,N_11215);
and U12337 (N_12337,N_9571,N_11454);
or U12338 (N_12338,N_9662,N_11261);
nand U12339 (N_12339,N_9182,N_9541);
nor U12340 (N_12340,N_11287,N_11421);
or U12341 (N_12341,N_10681,N_11334);
nand U12342 (N_12342,N_11264,N_10082);
nand U12343 (N_12343,N_9563,N_11258);
and U12344 (N_12344,N_11064,N_9193);
nand U12345 (N_12345,N_11078,N_11619);
nor U12346 (N_12346,N_9976,N_10023);
nand U12347 (N_12347,N_11715,N_9569);
nor U12348 (N_12348,N_11624,N_9172);
or U12349 (N_12349,N_10341,N_11377);
nand U12350 (N_12350,N_11410,N_9810);
and U12351 (N_12351,N_9791,N_11924);
nor U12352 (N_12352,N_10928,N_9526);
or U12353 (N_12353,N_10944,N_10913);
or U12354 (N_12354,N_9224,N_11879);
nand U12355 (N_12355,N_9474,N_9397);
and U12356 (N_12356,N_10418,N_11867);
nor U12357 (N_12357,N_11188,N_10504);
nor U12358 (N_12358,N_10972,N_9582);
xnor U12359 (N_12359,N_10834,N_9342);
xnor U12360 (N_12360,N_9780,N_9042);
nor U12361 (N_12361,N_9566,N_10098);
and U12362 (N_12362,N_10528,N_9806);
nand U12363 (N_12363,N_9220,N_9585);
or U12364 (N_12364,N_10079,N_10588);
nor U12365 (N_12365,N_9069,N_11729);
and U12366 (N_12366,N_9049,N_11816);
nand U12367 (N_12367,N_10850,N_9561);
nand U12368 (N_12368,N_9200,N_11483);
nor U12369 (N_12369,N_10729,N_9994);
nand U12370 (N_12370,N_11135,N_11789);
nor U12371 (N_12371,N_11643,N_11232);
nand U12372 (N_12372,N_9027,N_11848);
and U12373 (N_12373,N_10293,N_10675);
nand U12374 (N_12374,N_11596,N_11247);
xnor U12375 (N_12375,N_9331,N_9925);
or U12376 (N_12376,N_9490,N_10691);
and U12377 (N_12377,N_11388,N_11020);
or U12378 (N_12378,N_10953,N_9759);
nand U12379 (N_12379,N_10316,N_10587);
or U12380 (N_12380,N_10693,N_11263);
nor U12381 (N_12381,N_11830,N_10699);
nor U12382 (N_12382,N_9991,N_11043);
nor U12383 (N_12383,N_11851,N_11168);
nand U12384 (N_12384,N_9301,N_10777);
nand U12385 (N_12385,N_10434,N_11105);
and U12386 (N_12386,N_11373,N_10399);
nor U12387 (N_12387,N_9180,N_10907);
nand U12388 (N_12388,N_10631,N_10206);
nor U12389 (N_12389,N_9921,N_11918);
and U12390 (N_12390,N_9464,N_9271);
nor U12391 (N_12391,N_9647,N_11216);
nand U12392 (N_12392,N_11366,N_10347);
xor U12393 (N_12393,N_11540,N_11341);
nor U12394 (N_12394,N_10685,N_9743);
and U12395 (N_12395,N_11257,N_11530);
and U12396 (N_12396,N_10890,N_9558);
and U12397 (N_12397,N_11991,N_11037);
xor U12398 (N_12398,N_9476,N_11218);
nand U12399 (N_12399,N_9550,N_9133);
or U12400 (N_12400,N_9788,N_11096);
and U12401 (N_12401,N_11458,N_11769);
nand U12402 (N_12402,N_9318,N_9954);
nand U12403 (N_12403,N_11677,N_9782);
or U12404 (N_12404,N_11611,N_10968);
nand U12405 (N_12405,N_10063,N_11627);
and U12406 (N_12406,N_9324,N_9497);
nand U12407 (N_12407,N_11346,N_11963);
nor U12408 (N_12408,N_10052,N_9371);
or U12409 (N_12409,N_11937,N_10975);
or U12410 (N_12410,N_11251,N_11048);
xnor U12411 (N_12411,N_10067,N_10939);
or U12412 (N_12412,N_10798,N_11703);
or U12413 (N_12413,N_9374,N_9924);
nor U12414 (N_12414,N_11590,N_9912);
xnor U12415 (N_12415,N_10220,N_10745);
and U12416 (N_12416,N_11331,N_10014);
nor U12417 (N_12417,N_10787,N_10746);
nor U12418 (N_12418,N_11040,N_10908);
or U12419 (N_12419,N_11889,N_11817);
or U12420 (N_12420,N_10920,N_11212);
or U12421 (N_12421,N_11772,N_10240);
or U12422 (N_12422,N_9650,N_11947);
and U12423 (N_12423,N_9091,N_9504);
and U12424 (N_12424,N_9362,N_11418);
nand U12425 (N_12425,N_9465,N_9545);
and U12426 (N_12426,N_9126,N_11694);
nand U12427 (N_12427,N_10924,N_10496);
nand U12428 (N_12428,N_10325,N_9864);
nor U12429 (N_12429,N_9740,N_10559);
or U12430 (N_12430,N_10458,N_9075);
or U12431 (N_12431,N_9265,N_11629);
and U12432 (N_12432,N_10350,N_10988);
and U12433 (N_12433,N_10897,N_11700);
nor U12434 (N_12434,N_11412,N_9107);
and U12435 (N_12435,N_9118,N_9082);
or U12436 (N_12436,N_10252,N_10049);
nor U12437 (N_12437,N_10472,N_9310);
or U12438 (N_12438,N_9116,N_10176);
nand U12439 (N_12439,N_10236,N_11420);
or U12440 (N_12440,N_11322,N_10895);
or U12441 (N_12441,N_10604,N_11953);
or U12442 (N_12442,N_11167,N_9160);
and U12443 (N_12443,N_10507,N_10516);
nor U12444 (N_12444,N_9162,N_9323);
nand U12445 (N_12445,N_10658,N_11818);
or U12446 (N_12446,N_11569,N_9900);
nand U12447 (N_12447,N_9036,N_10165);
or U12448 (N_12448,N_11147,N_10663);
and U12449 (N_12449,N_11736,N_11883);
nor U12450 (N_12450,N_11681,N_10925);
or U12451 (N_12451,N_10964,N_9863);
and U12452 (N_12452,N_11143,N_10473);
or U12453 (N_12453,N_11370,N_9100);
xnor U12454 (N_12454,N_11567,N_10348);
or U12455 (N_12455,N_11801,N_9530);
xnor U12456 (N_12456,N_9671,N_9878);
or U12457 (N_12457,N_10678,N_11940);
and U12458 (N_12458,N_9907,N_9690);
or U12459 (N_12459,N_10478,N_9409);
and U12460 (N_12460,N_9376,N_10188);
nor U12461 (N_12461,N_11507,N_10062);
or U12462 (N_12462,N_9232,N_11989);
xnor U12463 (N_12463,N_11302,N_10672);
or U12464 (N_12464,N_10811,N_11966);
nand U12465 (N_12465,N_11355,N_11245);
and U12466 (N_12466,N_9989,N_9894);
and U12467 (N_12467,N_11171,N_11146);
and U12468 (N_12468,N_9939,N_10442);
or U12469 (N_12469,N_11902,N_10728);
nand U12470 (N_12470,N_9632,N_11669);
nor U12471 (N_12471,N_10501,N_11609);
and U12472 (N_12472,N_10106,N_11771);
nand U12473 (N_12473,N_10941,N_10467);
and U12474 (N_12474,N_10574,N_11730);
and U12475 (N_12475,N_10977,N_11201);
or U12476 (N_12476,N_11396,N_10011);
nand U12477 (N_12477,N_10698,N_11613);
nand U12478 (N_12478,N_11381,N_11280);
or U12479 (N_12479,N_11725,N_11574);
and U12480 (N_12480,N_10695,N_10408);
nor U12481 (N_12481,N_9758,N_11267);
nor U12482 (N_12482,N_10806,N_10998);
and U12483 (N_12483,N_10561,N_11988);
or U12484 (N_12484,N_10791,N_11990);
or U12485 (N_12485,N_11865,N_11293);
or U12486 (N_12486,N_11485,N_10078);
nand U12487 (N_12487,N_9452,N_9484);
nor U12488 (N_12488,N_10117,N_11958);
nand U12489 (N_12489,N_10567,N_9236);
or U12490 (N_12490,N_11743,N_10686);
and U12491 (N_12491,N_9672,N_9510);
nand U12492 (N_12492,N_10622,N_10943);
nor U12493 (N_12493,N_10210,N_10371);
or U12494 (N_12494,N_11186,N_9077);
nor U12495 (N_12495,N_11834,N_9827);
and U12496 (N_12496,N_10358,N_11164);
nand U12497 (N_12497,N_10757,N_10525);
xor U12498 (N_12498,N_10398,N_9972);
and U12499 (N_12499,N_10550,N_10232);
xor U12500 (N_12500,N_11081,N_10656);
and U12501 (N_12501,N_11808,N_10792);
xnor U12502 (N_12502,N_9733,N_9072);
and U12503 (N_12503,N_9233,N_11151);
or U12504 (N_12504,N_10475,N_10786);
or U12505 (N_12505,N_10424,N_11060);
and U12506 (N_12506,N_10199,N_9168);
nor U12507 (N_12507,N_11581,N_11877);
nand U12508 (N_12508,N_9273,N_11279);
or U12509 (N_12509,N_9019,N_9747);
nand U12510 (N_12510,N_10281,N_10050);
and U12511 (N_12511,N_9227,N_9093);
xor U12512 (N_12512,N_10654,N_9010);
nand U12513 (N_12513,N_10286,N_10915);
or U12514 (N_12514,N_11601,N_10397);
nor U12515 (N_12515,N_10743,N_9763);
nor U12516 (N_12516,N_9145,N_10482);
and U12517 (N_12517,N_9017,N_11654);
nand U12518 (N_12518,N_11169,N_9482);
nor U12519 (N_12519,N_11130,N_10549);
nand U12520 (N_12520,N_9385,N_9574);
nor U12521 (N_12521,N_11531,N_9151);
or U12522 (N_12522,N_11470,N_9057);
nor U12523 (N_12523,N_10981,N_11285);
and U12524 (N_12524,N_11281,N_10131);
nor U12525 (N_12525,N_11403,N_9866);
nand U12526 (N_12526,N_9966,N_10416);
or U12527 (N_12527,N_10314,N_9785);
nand U12528 (N_12528,N_9534,N_11398);
nor U12529 (N_12529,N_9559,N_10219);
nand U12530 (N_12530,N_9614,N_10414);
or U12531 (N_12531,N_11604,N_10195);
and U12532 (N_12532,N_9381,N_9893);
and U12533 (N_12533,N_11447,N_9877);
xor U12534 (N_12534,N_10033,N_11229);
nor U12535 (N_12535,N_10145,N_10554);
and U12536 (N_12536,N_9218,N_9902);
and U12537 (N_12537,N_11636,N_10615);
and U12538 (N_12538,N_10900,N_11484);
nand U12539 (N_12539,N_11901,N_10519);
or U12540 (N_12540,N_9192,N_11656);
nor U12541 (N_12541,N_11128,N_9487);
or U12542 (N_12542,N_11379,N_9333);
nor U12543 (N_12543,N_9293,N_9871);
nand U12544 (N_12544,N_9142,N_10762);
nor U12545 (N_12545,N_9702,N_11067);
or U12546 (N_12546,N_10935,N_9613);
or U12547 (N_12547,N_9104,N_11747);
nand U12548 (N_12548,N_10610,N_10028);
or U12549 (N_12549,N_10551,N_10345);
and U12550 (N_12550,N_9444,N_10919);
and U12551 (N_12551,N_10262,N_10859);
xor U12552 (N_12552,N_11083,N_11466);
and U12553 (N_12553,N_9432,N_11519);
nand U12554 (N_12554,N_11820,N_11430);
nor U12555 (N_12555,N_11459,N_11024);
and U12556 (N_12556,N_10104,N_11846);
or U12557 (N_12557,N_10364,N_11976);
nand U12558 (N_12558,N_11282,N_11597);
nand U12559 (N_12559,N_9716,N_10641);
nand U12560 (N_12560,N_9521,N_10093);
nor U12561 (N_12561,N_9459,N_11363);
nand U12562 (N_12562,N_10508,N_11453);
nor U12563 (N_12563,N_10952,N_10863);
nand U12564 (N_12564,N_9996,N_10268);
nand U12565 (N_12565,N_9636,N_11560);
nor U12566 (N_12566,N_11413,N_10247);
nor U12567 (N_12567,N_10058,N_11325);
and U12568 (N_12568,N_9700,N_10027);
nand U12569 (N_12569,N_11870,N_10355);
xor U12570 (N_12570,N_9053,N_11929);
and U12571 (N_12571,N_10303,N_9478);
nand U12572 (N_12572,N_10019,N_11814);
nor U12573 (N_12573,N_11984,N_10662);
or U12574 (N_12574,N_9191,N_10317);
or U12575 (N_12575,N_10460,N_9699);
nor U12576 (N_12576,N_11330,N_10081);
nand U12577 (N_12577,N_11548,N_11116);
nor U12578 (N_12578,N_10400,N_10321);
and U12579 (N_12579,N_10189,N_9769);
nor U12580 (N_12580,N_11970,N_11835);
nand U12581 (N_12581,N_9732,N_10623);
nand U12582 (N_12582,N_11987,N_10100);
nand U12583 (N_12583,N_11767,N_10936);
and U12584 (N_12584,N_11347,N_9812);
nor U12585 (N_12585,N_10103,N_10861);
nand U12586 (N_12586,N_10039,N_9335);
or U12587 (N_12587,N_10102,N_11362);
nor U12588 (N_12588,N_9378,N_10163);
nand U12589 (N_12589,N_10448,N_9033);
nor U12590 (N_12590,N_11441,N_9537);
nand U12591 (N_12591,N_11776,N_10726);
nor U12592 (N_12592,N_9667,N_11803);
nor U12593 (N_12593,N_11115,N_9993);
nand U12594 (N_12594,N_9485,N_10957);
and U12595 (N_12595,N_11993,N_10296);
and U12596 (N_12596,N_10196,N_11489);
and U12597 (N_12597,N_9286,N_9624);
nor U12598 (N_12598,N_11354,N_9797);
xor U12599 (N_12599,N_9365,N_10835);
and U12600 (N_12600,N_11806,N_9288);
xor U12601 (N_12601,N_11994,N_11985);
or U12602 (N_12602,N_11195,N_11580);
xnor U12603 (N_12603,N_9774,N_10144);
nand U12604 (N_12604,N_9962,N_11943);
or U12605 (N_12605,N_11515,N_9197);
and U12606 (N_12606,N_10048,N_9410);
and U12607 (N_12607,N_10705,N_11753);
and U12608 (N_12608,N_9076,N_9638);
nor U12609 (N_12609,N_9606,N_9114);
xor U12610 (N_12610,N_10951,N_9440);
nand U12611 (N_12611,N_11018,N_11374);
nor U12612 (N_12612,N_10449,N_11163);
and U12613 (N_12613,N_11563,N_9519);
nand U12614 (N_12614,N_10439,N_11642);
nor U12615 (N_12615,N_10065,N_9839);
xor U12616 (N_12616,N_9255,N_9778);
nand U12617 (N_12617,N_10738,N_9637);
nor U12618 (N_12618,N_11444,N_11856);
nor U12619 (N_12619,N_9348,N_10808);
nand U12620 (N_12620,N_11822,N_10109);
nand U12621 (N_12621,N_9744,N_9997);
nor U12622 (N_12622,N_11706,N_9174);
and U12623 (N_12623,N_11908,N_11184);
nor U12624 (N_12624,N_10837,N_10878);
nor U12625 (N_12625,N_10006,N_11304);
and U12626 (N_12626,N_10090,N_11699);
nor U12627 (N_12627,N_11250,N_9454);
nand U12628 (N_12628,N_9395,N_11541);
nor U12629 (N_12629,N_10917,N_10118);
nand U12630 (N_12630,N_10780,N_11382);
nor U12631 (N_12631,N_11644,N_11898);
nor U12632 (N_12632,N_10429,N_9595);
or U12633 (N_12633,N_10499,N_11004);
and U12634 (N_12634,N_9936,N_9383);
and U12635 (N_12635,N_9020,N_10876);
and U12636 (N_12636,N_9289,N_9252);
nor U12637 (N_12637,N_9590,N_10521);
nor U12638 (N_12638,N_10883,N_10407);
or U12639 (N_12639,N_9430,N_10334);
or U12640 (N_12640,N_10946,N_9967);
and U12641 (N_12641,N_10869,N_10072);
nor U12642 (N_12642,N_11463,N_9396);
nand U12643 (N_12643,N_9488,N_10639);
or U12644 (N_12644,N_11620,N_10945);
and U12645 (N_12645,N_9144,N_10272);
nor U12646 (N_12646,N_11634,N_11858);
or U12647 (N_12647,N_11133,N_10733);
and U12648 (N_12648,N_9717,N_9158);
nand U12649 (N_12649,N_10569,N_9825);
nand U12650 (N_12650,N_9054,N_11948);
nor U12651 (N_12651,N_11290,N_9603);
and U12652 (N_12652,N_11274,N_11652);
nor U12653 (N_12653,N_11873,N_10451);
or U12654 (N_12654,N_9352,N_10291);
or U12655 (N_12655,N_11271,N_11003);
and U12656 (N_12656,N_11339,N_11390);
xnor U12657 (N_12657,N_11144,N_9875);
nand U12658 (N_12658,N_11785,N_10514);
and U12659 (N_12659,N_11348,N_10216);
and U12660 (N_12660,N_10541,N_10522);
nand U12661 (N_12661,N_11154,N_9838);
nor U12662 (N_12662,N_9115,N_10758);
and U12663 (N_12663,N_9489,N_9393);
and U12664 (N_12664,N_9556,N_9661);
nand U12665 (N_12665,N_9620,N_10760);
nand U12666 (N_12666,N_9762,N_11614);
or U12667 (N_12667,N_10411,N_9190);
xnor U12668 (N_12668,N_11034,N_9317);
nor U12669 (N_12669,N_10769,N_11451);
nor U12670 (N_12670,N_11595,N_10857);
nor U12671 (N_12671,N_11344,N_11335);
nand U12672 (N_12672,N_10707,N_11742);
and U12673 (N_12673,N_10259,N_11954);
nor U12674 (N_12674,N_11142,N_10828);
nand U12675 (N_12675,N_9261,N_9285);
nand U12676 (N_12676,N_10579,N_11001);
nor U12677 (N_12677,N_10089,N_10680);
and U12678 (N_12678,N_11448,N_10485);
and U12679 (N_12679,N_9658,N_9553);
or U12680 (N_12680,N_10035,N_11679);
nor U12681 (N_12681,N_10867,N_9955);
and U12682 (N_12682,N_9673,N_9471);
xnor U12683 (N_12683,N_11108,N_10985);
and U12684 (N_12684,N_11663,N_9723);
nor U12685 (N_12685,N_10382,N_9070);
nand U12686 (N_12686,N_9389,N_9514);
and U12687 (N_12687,N_10933,N_11942);
and U12688 (N_12688,N_9675,N_11357);
xnor U12689 (N_12689,N_11314,N_11805);
and U12690 (N_12690,N_11571,N_10233);
nor U12691 (N_12691,N_11496,N_9605);
and U12692 (N_12692,N_10271,N_10289);
and U12693 (N_12693,N_11503,N_9722);
and U12694 (N_12694,N_9640,N_9340);
and U12695 (N_12695,N_9039,N_10635);
nor U12696 (N_12696,N_11535,N_9952);
nor U12697 (N_12697,N_10459,N_9470);
xnor U12698 (N_12698,N_11751,N_9248);
nand U12699 (N_12699,N_11907,N_9617);
nor U12700 (N_12700,N_9290,N_9736);
or U12701 (N_12701,N_10873,N_11714);
and U12702 (N_12702,N_9988,N_11602);
or U12703 (N_12703,N_9463,N_11471);
nor U12704 (N_12704,N_9123,N_11599);
nor U12705 (N_12705,N_11885,N_10068);
or U12706 (N_12706,N_11732,N_9111);
or U12707 (N_12707,N_11092,N_11955);
nor U12708 (N_12708,N_11407,N_9815);
nand U12709 (N_12709,N_11582,N_11204);
xnor U12710 (N_12710,N_11109,N_11345);
nand U12711 (N_12711,N_9336,N_11234);
and U12712 (N_12712,N_9391,N_11704);
nand U12713 (N_12713,N_11155,N_9890);
xnor U12714 (N_12714,N_10147,N_9517);
nand U12715 (N_12715,N_9881,N_10304);
and U12716 (N_12716,N_11539,N_11415);
or U12717 (N_12717,N_9048,N_9824);
nor U12718 (N_12718,N_9141,N_9920);
nand U12719 (N_12719,N_10086,N_9425);
and U12720 (N_12720,N_10722,N_11180);
xnor U12721 (N_12721,N_11944,N_9741);
or U12722 (N_12722,N_11002,N_9280);
nand U12723 (N_12723,N_9032,N_10836);
nor U12724 (N_12724,N_10856,N_10805);
nand U12725 (N_12725,N_10584,N_11533);
or U12726 (N_12726,N_10228,N_9436);
nor U12727 (N_12727,N_10982,N_11522);
and U12728 (N_12728,N_11051,N_9849);
or U12729 (N_12729,N_11493,N_10692);
or U12730 (N_12730,N_10070,N_9995);
nor U12731 (N_12731,N_9472,N_9355);
nand U12732 (N_12732,N_10599,N_10822);
and U12733 (N_12733,N_10186,N_10126);
or U12734 (N_12734,N_9512,N_9105);
or U12735 (N_12735,N_9153,N_9243);
nor U12736 (N_12736,N_10122,N_11066);
nand U12737 (N_12737,N_11551,N_11006);
or U12738 (N_12738,N_11446,N_11837);
and U12739 (N_12739,N_10363,N_9460);
xor U12740 (N_12740,N_11635,N_11177);
nor U12741 (N_12741,N_10338,N_9079);
nand U12742 (N_12742,N_9302,N_9568);
xnor U12743 (N_12743,N_11249,N_9833);
and U12744 (N_12744,N_11612,N_10580);
nand U12745 (N_12745,N_9332,N_9368);
nor U12746 (N_12746,N_11749,N_10297);
and U12747 (N_12747,N_9745,N_9856);
nor U12748 (N_12748,N_11552,N_10770);
and U12749 (N_12749,N_9110,N_9373);
nand U12750 (N_12750,N_11784,N_9549);
or U12751 (N_12751,N_11479,N_10864);
and U12752 (N_12752,N_10084,N_11272);
xor U12753 (N_12753,N_9684,N_10454);
nand U12754 (N_12754,N_11284,N_9909);
nor U12755 (N_12755,N_10815,N_11465);
and U12756 (N_12756,N_9768,N_11467);
nor U12757 (N_12757,N_11477,N_10673);
xor U12758 (N_12758,N_9155,N_10716);
nand U12759 (N_12759,N_10849,N_9528);
or U12760 (N_12760,N_10609,N_9898);
nor U12761 (N_12761,N_10773,N_9171);
and U12762 (N_12762,N_9513,N_9730);
nor U12763 (N_12763,N_9085,N_10589);
nor U12764 (N_12764,N_11799,N_10396);
nor U12765 (N_12765,N_9064,N_9652);
or U12766 (N_12766,N_9992,N_11174);
xor U12767 (N_12767,N_10948,N_10542);
or U12768 (N_12768,N_10688,N_9305);
nor U12769 (N_12769,N_10788,N_11872);
or U12770 (N_12770,N_9616,N_10558);
nor U12771 (N_12771,N_9844,N_11079);
or U12772 (N_12772,N_10638,N_11857);
or U12773 (N_12773,N_11364,N_9279);
and U12774 (N_12774,N_9888,N_10969);
nor U12775 (N_12775,N_10555,N_10223);
nor U12776 (N_12776,N_11259,N_9254);
and U12777 (N_12777,N_9071,N_11946);
or U12778 (N_12778,N_9963,N_9356);
or U12779 (N_12779,N_11191,N_10595);
and U12780 (N_12780,N_9018,N_9351);
nand U12781 (N_12781,N_11492,N_9166);
nand U12782 (N_12782,N_11683,N_10158);
nand U12783 (N_12783,N_10315,N_10209);
nor U12784 (N_12784,N_10071,N_9578);
nand U12785 (N_12785,N_9202,N_11340);
and U12786 (N_12786,N_9858,N_10719);
nor U12787 (N_12787,N_10825,N_11214);
and U12788 (N_12788,N_9495,N_9353);
xnor U12789 (N_12789,N_11450,N_11810);
nand U12790 (N_12790,N_10776,N_10450);
or U12791 (N_12791,N_11052,N_10200);
xor U12792 (N_12792,N_9347,N_9783);
and U12793 (N_12793,N_10629,N_11874);
and U12794 (N_12794,N_9599,N_9026);
nor U12795 (N_12795,N_9003,N_9065);
and U12796 (N_12796,N_9591,N_10251);
and U12797 (N_12797,N_11482,N_9799);
nor U12798 (N_12798,N_9216,N_10660);
or U12799 (N_12799,N_9300,N_11198);
or U12800 (N_12800,N_10197,N_11792);
nand U12801 (N_12801,N_9986,N_10142);
nand U12802 (N_12802,N_11499,N_11972);
nand U12803 (N_12803,N_10978,N_9548);
nand U12804 (N_12804,N_10224,N_10248);
or U12805 (N_12805,N_9011,N_11579);
or U12806 (N_12806,N_11120,N_10092);
xnor U12807 (N_12807,N_11861,N_11328);
or U12808 (N_12808,N_10111,N_11709);
or U12809 (N_12809,N_11210,N_9709);
or U12810 (N_12810,N_10125,N_10721);
xnor U12811 (N_12811,N_11969,N_9291);
or U12812 (N_12812,N_11022,N_11426);
xnor U12813 (N_12813,N_10372,N_10128);
nor U12814 (N_12814,N_10735,N_10380);
and U12815 (N_12815,N_11333,N_11562);
nand U12816 (N_12816,N_11761,N_10229);
nand U12817 (N_12817,N_10124,N_11055);
or U12818 (N_12818,N_10976,N_10566);
nor U12819 (N_12819,N_11667,N_9725);
and U12820 (N_12820,N_11711,N_9095);
nand U12821 (N_12821,N_11520,N_9188);
or U12822 (N_12822,N_10343,N_11717);
or U12823 (N_12823,N_11941,N_11008);
nor U12824 (N_12824,N_9312,N_11068);
nand U12825 (N_12825,N_11862,N_10433);
nand U12826 (N_12826,N_10967,N_10795);
nor U12827 (N_12827,N_11840,N_11075);
nor U12828 (N_12828,N_10644,N_9724);
or U12829 (N_12829,N_9687,N_11593);
nand U12830 (N_12830,N_11977,N_9380);
xnor U12831 (N_12831,N_10425,N_10697);
or U12832 (N_12832,N_10095,N_11027);
xnor U12833 (N_12833,N_11244,N_9848);
and U12834 (N_12834,N_11397,N_10115);
and U12835 (N_12835,N_11085,N_10445);
and U12836 (N_12836,N_9639,N_11227);
nand U12837 (N_12837,N_10222,N_11592);
nand U12838 (N_12838,N_9390,N_9439);
nand U12839 (N_12839,N_9012,N_11623);
and U12840 (N_12840,N_10986,N_10520);
nand U12841 (N_12841,N_11416,N_9657);
or U12842 (N_12842,N_11565,N_11080);
nand U12843 (N_12843,N_10546,N_9755);
or U12844 (N_12844,N_10308,N_9914);
nor U12845 (N_12845,N_10752,N_9157);
nand U12846 (N_12846,N_10034,N_9748);
nand U12847 (N_12847,N_10591,N_10244);
nor U12848 (N_12848,N_11385,N_11372);
nor U12849 (N_12849,N_11550,N_11591);
and U12850 (N_12850,N_10492,N_9414);
and U12851 (N_12851,N_9084,N_10391);
nor U12852 (N_12852,N_11219,N_9163);
xor U12853 (N_12853,N_11734,N_11961);
nor U12854 (N_12854,N_9016,N_10696);
xnor U12855 (N_12855,N_9600,N_9808);
or U12856 (N_12856,N_10392,N_10468);
xnor U12857 (N_12857,N_9398,N_9692);
xnor U12858 (N_12858,N_9911,N_10129);
xnor U12859 (N_12859,N_11916,N_9441);
and U12860 (N_12860,N_10754,N_10793);
nand U12861 (N_12861,N_10961,N_9058);
and U12862 (N_12862,N_10854,N_11787);
xor U12863 (N_12863,N_11076,N_11138);
or U12864 (N_12864,N_11386,N_11192);
and U12865 (N_12865,N_9670,N_9618);
or U12866 (N_12866,N_11208,N_11206);
nand U12867 (N_12867,N_11183,N_9253);
and U12868 (N_12868,N_9836,N_11455);
nor U12869 (N_12869,N_10744,N_11938);
nand U12870 (N_12870,N_11074,N_11891);
and U12871 (N_12871,N_11114,N_9974);
and U12872 (N_12872,N_10486,N_11095);
and U12873 (N_12873,N_11782,N_9676);
nor U12874 (N_12874,N_10993,N_9103);
nor U12875 (N_12875,N_9554,N_10775);
xnor U12876 (N_12876,N_9306,N_10643);
nor U12877 (N_12877,N_10470,N_11645);
or U12878 (N_12878,N_11125,N_11278);
nor U12879 (N_12879,N_10995,N_9507);
and U12880 (N_12880,N_11021,N_11625);
or U12881 (N_12881,N_10960,N_10804);
nor U12882 (N_12882,N_9837,N_11494);
nor U12883 (N_12883,N_10198,N_9407);
and U12884 (N_12884,N_9442,N_9853);
or U12885 (N_12885,N_11193,N_11152);
or U12886 (N_12886,N_9152,N_10749);
or U12887 (N_12887,N_10689,N_11353);
nand U12888 (N_12888,N_11884,N_9719);
and U12889 (N_12889,N_11913,N_11276);
nand U12890 (N_12890,N_10649,N_10706);
nand U12891 (N_12891,N_9801,N_9916);
nand U12892 (N_12892,N_9207,N_10044);
nor U12893 (N_12893,N_9446,N_10088);
nand U12894 (N_12894,N_11359,N_9241);
nand U12895 (N_12895,N_10532,N_9242);
xor U12896 (N_12896,N_11486,N_9127);
and U12897 (N_12897,N_9415,N_9969);
or U12898 (N_12898,N_10401,N_9339);
and U12899 (N_12899,N_11481,N_10342);
and U12900 (N_12900,N_9932,N_11089);
and U12901 (N_12901,N_10712,N_10794);
xor U12902 (N_12902,N_9942,N_11196);
nor U12903 (N_12903,N_10818,N_11705);
xor U12904 (N_12904,N_10764,N_10462);
and U12905 (N_12905,N_11588,N_9462);
nand U12906 (N_12906,N_9790,N_9044);
nor U12907 (N_12907,N_10802,N_10753);
nor U12908 (N_12908,N_11185,N_9906);
or U12909 (N_12909,N_10565,N_9520);
nor U12910 (N_12910,N_10269,N_11181);
or U12911 (N_12911,N_9297,N_10013);
nand U12912 (N_12912,N_9119,N_9004);
and U12913 (N_12913,N_9682,N_9917);
or U12914 (N_12914,N_11659,N_11741);
xnor U12915 (N_12915,N_10955,N_11118);
and U12916 (N_12916,N_9779,N_11697);
xor U12917 (N_12917,N_11433,N_11917);
and U12918 (N_12918,N_10456,N_9681);
xor U12919 (N_12919,N_11236,N_10741);
nor U12920 (N_12920,N_11033,N_9543);
xnor U12921 (N_12921,N_9958,N_9742);
or U12922 (N_12922,N_9666,N_11707);
nand U12923 (N_12923,N_9816,N_10309);
nor U12924 (N_12924,N_11107,N_11853);
nor U12925 (N_12925,N_9739,N_11502);
xnor U12926 (N_12926,N_10007,N_10677);
nand U12927 (N_12927,N_9492,N_11157);
and U12928 (N_12928,N_11010,N_11744);
or U12929 (N_12929,N_11757,N_9535);
and U12930 (N_12930,N_11881,N_11900);
nand U12931 (N_12931,N_11461,N_11313);
nand U12932 (N_12932,N_11529,N_11832);
nand U12933 (N_12933,N_11575,N_10871);
and U12934 (N_12934,N_10046,N_10533);
nor U12935 (N_12935,N_11691,N_10646);
nor U12936 (N_12936,N_9394,N_11099);
xnor U12937 (N_12937,N_10108,N_10899);
or U12938 (N_12938,N_9313,N_11628);
nor U12939 (N_12939,N_9982,N_9882);
or U12940 (N_12940,N_10842,N_10538);
nand U12941 (N_12941,N_9642,N_9189);
nand U12942 (N_12942,N_9028,N_9344);
nor U12943 (N_12943,N_10426,N_10618);
nor U12944 (N_12944,N_11252,N_9402);
and U12945 (N_12945,N_11310,N_10318);
nor U12946 (N_12946,N_10617,N_10330);
and U12947 (N_12947,N_9421,N_10847);
nor U12948 (N_12948,N_10931,N_9777);
nor U12949 (N_12949,N_9683,N_9179);
or U12950 (N_12950,N_9800,N_11882);
nor U12951 (N_12951,N_10751,N_10150);
or U12952 (N_12952,N_11209,N_10385);
xor U12953 (N_12953,N_10335,N_9223);
nand U12954 (N_12954,N_9343,N_9014);
nand U12955 (N_12955,N_11587,N_9861);
nand U12956 (N_12956,N_9987,N_9892);
nor U12957 (N_12957,N_10218,N_10140);
xnor U12958 (N_12958,N_10740,N_9205);
nand U12959 (N_12959,N_10237,N_11760);
and U12960 (N_12960,N_11141,N_10280);
nand U12961 (N_12961,N_10860,N_11855);
and U12962 (N_12962,N_10324,N_11073);
or U12963 (N_12963,N_10906,N_9531);
and U12964 (N_12964,N_11570,N_11371);
or U12965 (N_12965,N_10221,N_11827);
xor U12966 (N_12966,N_10370,N_9278);
nand U12967 (N_12967,N_10181,N_10096);
or U12968 (N_12968,N_10768,N_11737);
and U12969 (N_12969,N_10016,N_10241);
nand U12970 (N_12970,N_10498,N_9677);
nor U12971 (N_12971,N_9456,N_10453);
or U12972 (N_12972,N_9025,N_10127);
nand U12973 (N_12973,N_9330,N_10774);
nand U12974 (N_12974,N_11660,N_9678);
and U12975 (N_12975,N_9098,N_11893);
and U12976 (N_12976,N_11553,N_9249);
and U12977 (N_12977,N_10929,N_10484);
and U12978 (N_12978,N_11600,N_9821);
nor U12979 (N_12979,N_10817,N_10767);
and U12980 (N_12980,N_11472,N_11790);
or U12981 (N_12981,N_11131,N_11427);
and U12982 (N_12982,N_9124,N_9840);
nor U12983 (N_12983,N_9927,N_10922);
xnor U12984 (N_12984,N_9304,N_11545);
or U12985 (N_12985,N_11649,N_10266);
nor U12986 (N_12986,N_11712,N_10390);
nand U12987 (N_12987,N_10420,N_10880);
xor U12988 (N_12988,N_9268,N_11432);
xnor U12989 (N_12989,N_9475,N_9140);
nor U12990 (N_12990,N_11262,N_10042);
and U12991 (N_12991,N_9899,N_9525);
nand U12992 (N_12992,N_9786,N_9664);
and U12993 (N_12993,N_11480,N_9884);
nand U12994 (N_12994,N_10910,N_9704);
and U12995 (N_12995,N_10037,N_10750);
nor U12996 (N_12996,N_10984,N_9185);
nor U12997 (N_12997,N_11406,N_11915);
and U12998 (N_12998,N_10601,N_9328);
nand U12999 (N_12999,N_10040,N_11332);
and U13000 (N_13000,N_10166,N_9473);
and U13001 (N_13001,N_11026,N_9931);
or U13002 (N_13002,N_11094,N_10141);
and U13003 (N_13003,N_11788,N_11925);
and U13004 (N_13004,N_11819,N_9668);
nand U13005 (N_13005,N_11573,N_9770);
nor U13006 (N_13006,N_10403,N_11098);
xor U13007 (N_13007,N_10463,N_9051);
nor U13008 (N_13008,N_11041,N_9625);
nor U13009 (N_13009,N_11686,N_11007);
xor U13010 (N_13010,N_11134,N_9257);
and U13011 (N_13011,N_10781,N_10973);
nor U13012 (N_13012,N_11005,N_9860);
and U13013 (N_13013,N_10018,N_11910);
and U13014 (N_13014,N_9651,N_9325);
or U13015 (N_13015,N_9129,N_11343);
nor U13016 (N_13016,N_11283,N_9081);
and U13017 (N_13017,N_11777,N_9735);
nor U13018 (N_13018,N_10598,N_9384);
or U13019 (N_13019,N_10500,N_11104);
xor U13020 (N_13020,N_11836,N_9822);
or U13021 (N_13021,N_9136,N_10120);
nor U13022 (N_13022,N_10202,N_9037);
and U13023 (N_13023,N_9417,N_11358);
nor U13024 (N_13024,N_11013,N_10540);
xnor U13025 (N_13025,N_11852,N_11295);
or U13026 (N_13026,N_11510,N_10886);
nor U13027 (N_13027,N_9872,N_11959);
and U13028 (N_13028,N_9830,N_9983);
or U13029 (N_13029,N_11880,N_9654);
nand U13030 (N_13030,N_10362,N_9181);
nand U13031 (N_13031,N_10627,N_10203);
or U13032 (N_13032,N_10008,N_10642);
nand U13033 (N_13033,N_9001,N_9309);
nand U13034 (N_13034,N_10245,N_10659);
and U13035 (N_13035,N_11260,N_9349);
or U13036 (N_13036,N_10417,N_9196);
nand U13037 (N_13037,N_10700,N_10155);
nor U13038 (N_13038,N_9320,N_9965);
or U13039 (N_13039,N_11384,N_10279);
or U13040 (N_13040,N_11726,N_11317);
or U13041 (N_13041,N_11139,N_11411);
or U13042 (N_13042,N_11246,N_11695);
nor U13043 (N_13043,N_10684,N_10841);
xnor U13044 (N_13044,N_11653,N_9948);
and U13045 (N_13045,N_10225,N_9013);
and U13046 (N_13046,N_9269,N_10329);
nor U13047 (N_13047,N_10374,N_9831);
nand U13048 (N_13048,N_10283,N_9922);
xnor U13049 (N_13049,N_11424,N_9212);
nand U13050 (N_13050,N_9859,N_10647);
or U13051 (N_13051,N_11367,N_11687);
nand U13052 (N_13052,N_9648,N_9583);
nand U13053 (N_13053,N_9038,N_9401);
or U13054 (N_13054,N_9131,N_10017);
or U13055 (N_13055,N_10628,N_9579);
nor U13056 (N_13056,N_9981,N_10471);
and U13057 (N_13057,N_11431,N_11030);
or U13058 (N_13058,N_9400,N_10254);
nor U13059 (N_13059,N_10645,N_9933);
xnor U13060 (N_13060,N_9663,N_11903);
nor U13061 (N_13061,N_11564,N_9370);
and U13062 (N_13062,N_10717,N_10022);
xnor U13063 (N_13063,N_10253,N_9178);
or U13064 (N_13064,N_10846,N_11360);
or U13065 (N_13065,N_9176,N_11768);
nor U13066 (N_13066,N_11640,N_10893);
and U13067 (N_13067,N_11508,N_10529);
or U13068 (N_13068,N_9496,N_11324);
or U13069 (N_13069,N_10572,N_11847);
nand U13070 (N_13070,N_10536,N_9796);
xnor U13071 (N_13071,N_9794,N_9850);
or U13072 (N_13072,N_10790,N_11648);
or U13073 (N_13073,N_9951,N_9219);
nor U13074 (N_13074,N_9589,N_11518);
nor U13075 (N_13075,N_9458,N_11266);
and U13076 (N_13076,N_10489,N_11904);
nor U13077 (N_13077,N_11057,N_9611);
nand U13078 (N_13078,N_9660,N_11674);
nor U13079 (N_13079,N_10714,N_11598);
nor U13080 (N_13080,N_10518,N_9619);
nor U13081 (N_13081,N_9135,N_10257);
and U13082 (N_13082,N_11009,N_11914);
or U13083 (N_13083,N_10234,N_9627);
xnor U13084 (N_13084,N_9275,N_9622);
nor U13085 (N_13085,N_11449,N_9873);
xor U13086 (N_13086,N_10436,N_10495);
and U13087 (N_13087,N_10172,N_11650);
nand U13088 (N_13088,N_10592,N_11500);
or U13089 (N_13089,N_9329,N_9267);
nand U13090 (N_13090,N_10381,N_11228);
xnor U13091 (N_13091,N_10275,N_11307);
or U13092 (N_13092,N_11072,N_10373);
nor U13093 (N_13093,N_11255,N_9005);
nand U13094 (N_13094,N_11626,N_10180);
nand U13095 (N_13095,N_11829,N_11166);
nor U13096 (N_13096,N_9819,N_10590);
or U13097 (N_13097,N_11689,N_9222);
nand U13098 (N_13098,N_10832,N_9399);
nor U13099 (N_13099,N_11796,N_10205);
and U13100 (N_13100,N_11056,N_10826);
nand U13101 (N_13101,N_11825,N_9046);
or U13102 (N_13102,N_11682,N_10012);
and U13103 (N_13103,N_10307,N_9481);
nand U13104 (N_13104,N_10080,N_10534);
nor U13105 (N_13105,N_10575,N_9707);
nand U13106 (N_13106,N_10715,N_11140);
or U13107 (N_13107,N_9646,N_10173);
nor U13108 (N_13108,N_9424,N_10059);
nor U13109 (N_13109,N_9703,N_11175);
nand U13110 (N_13110,N_11061,N_10509);
and U13111 (N_13111,N_11997,N_11275);
and U13112 (N_13112,N_11983,N_10858);
nor U13113 (N_13113,N_9804,N_11289);
or U13114 (N_13114,N_11664,N_10217);
and U13115 (N_13115,N_9210,N_11239);
nand U13116 (N_13116,N_10265,N_11965);
and U13117 (N_13117,N_11684,N_10367);
nand U13118 (N_13118,N_11437,N_10132);
or U13119 (N_13119,N_10724,N_10051);
nand U13120 (N_13120,N_11378,N_10980);
nand U13121 (N_13121,N_10896,N_9229);
and U13122 (N_13122,N_10614,N_10427);
and U13123 (N_13123,N_9074,N_10848);
and U13124 (N_13124,N_10620,N_10543);
nor U13125 (N_13125,N_9938,N_10612);
and U13126 (N_13126,N_11802,N_10606);
nor U13127 (N_13127,N_9607,N_11975);
or U13128 (N_13128,N_9338,N_10497);
or U13129 (N_13129,N_9298,N_10747);
nand U13130 (N_13130,N_10146,N_9260);
or U13131 (N_13131,N_11544,N_11671);
and U13132 (N_13132,N_9577,N_9388);
and U13133 (N_13133,N_11863,N_9408);
and U13134 (N_13134,N_10395,N_11501);
or U13135 (N_13135,N_11871,N_11127);
nor U13136 (N_13136,N_10074,N_11391);
nor U13137 (N_13137,N_9752,N_11895);
nor U13138 (N_13138,N_10855,N_9357);
and U13139 (N_13139,N_11713,N_9686);
xnor U13140 (N_13140,N_11735,N_10884);
nand U13141 (N_13141,N_9685,N_9148);
or U13142 (N_13142,N_11971,N_10909);
nor U13143 (N_13143,N_9466,N_9083);
nand U13144 (N_13144,N_11042,N_11511);
or U13145 (N_13145,N_9708,N_9341);
nand U13146 (N_13146,N_9567,N_11243);
and U13147 (N_13147,N_10273,N_11923);
nor U13148 (N_13148,N_11812,N_9327);
nor U13149 (N_13149,N_10110,N_11842);
nand U13150 (N_13150,N_11129,N_11460);
and U13151 (N_13151,N_11739,N_11082);
nand U13152 (N_13152,N_10340,N_11568);
and U13153 (N_13153,N_10581,N_10267);
and U13154 (N_13154,N_10851,N_9483);
and U13155 (N_13155,N_11662,N_9897);
and U13156 (N_13156,N_10958,N_11647);
nand U13157 (N_13157,N_11071,N_10657);
or U13158 (N_13158,N_10077,N_11538);
nand U13159 (N_13159,N_9052,N_10356);
xnor U13160 (N_13160,N_9891,N_10421);
and U13161 (N_13161,N_9542,N_10937);
nor U13162 (N_13162,N_11719,N_9040);
nor U13163 (N_13163,N_11922,N_9067);
and U13164 (N_13164,N_9846,N_11301);
or U13165 (N_13165,N_10830,N_10625);
nand U13166 (N_13166,N_11979,N_9120);
nand U13167 (N_13167,N_9696,N_11524);
nand U13168 (N_13168,N_9493,N_11439);
and U13169 (N_13169,N_11473,N_10630);
or U13170 (N_13170,N_9776,N_10069);
or U13171 (N_13171,N_9272,N_11160);
nand U13172 (N_13172,N_11409,N_10226);
and U13173 (N_13173,N_11536,N_10376);
nand U13174 (N_13174,N_11770,N_10311);
or U13175 (N_13175,N_11435,N_9108);
nor U13176 (N_13176,N_11238,N_9832);
nor U13177 (N_13177,N_11933,N_10346);
or U13178 (N_13178,N_10730,N_10194);
nor U13179 (N_13179,N_11621,N_11179);
xor U13180 (N_13180,N_11868,N_9669);
nor U13181 (N_13181,N_10779,N_9977);
nor U13182 (N_13182,N_11962,N_11176);
nand U13183 (N_13183,N_10261,N_10942);
and U13184 (N_13184,N_9437,N_9855);
nand U13185 (N_13185,N_10285,N_11070);
nand U13186 (N_13186,N_9710,N_9540);
and U13187 (N_13187,N_9754,N_11487);
nand U13188 (N_13188,N_9059,N_10613);
nand U13189 (N_13189,N_10365,N_9919);
or U13190 (N_13190,N_10464,N_10287);
and U13191 (N_13191,N_9727,N_9307);
nand U13192 (N_13192,N_10870,N_10997);
and U13193 (N_13193,N_11122,N_10255);
xnor U13194 (N_13194,N_11047,N_9555);
or U13195 (N_13195,N_9805,N_9945);
nand U13196 (N_13196,N_11934,N_9167);
nor U13197 (N_13197,N_11428,N_9086);
or U13198 (N_13198,N_11035,N_9154);
nand U13199 (N_13199,N_9694,N_9354);
and U13200 (N_13200,N_11286,N_11170);
xor U13201 (N_13201,N_11864,N_11069);
xor U13202 (N_13202,N_10029,N_10703);
nand U13203 (N_13203,N_11323,N_10483);
and U13204 (N_13204,N_9775,N_9818);
nor U13205 (N_13205,N_9096,N_9792);
or U13206 (N_13206,N_10725,N_9726);
and U13207 (N_13207,N_9125,N_11731);
and U13208 (N_13208,N_10650,N_10892);
nor U13209 (N_13209,N_11361,N_10637);
nor U13210 (N_13210,N_9649,N_11392);
nor U13211 (N_13211,N_9372,N_10292);
and U13212 (N_13212,N_11084,N_11797);
nor U13213 (N_13213,N_11566,N_10388);
or U13214 (N_13214,N_10923,N_10384);
or U13215 (N_13215,N_10351,N_9787);
and U13216 (N_13216,N_10178,N_9841);
nand U13217 (N_13217,N_9851,N_11248);
xnor U13218 (N_13218,N_9511,N_9772);
nor U13219 (N_13219,N_9311,N_9469);
and U13220 (N_13220,N_10157,N_11632);
and U13221 (N_13221,N_9876,N_11029);
or U13222 (N_13222,N_9411,N_11905);
xor U13223 (N_13223,N_11124,N_10153);
and U13224 (N_13224,N_10889,N_9913);
nand U13225 (N_13225,N_9369,N_10001);
or U13226 (N_13226,N_11112,N_11876);
nand U13227 (N_13227,N_9598,N_9610);
nor U13228 (N_13228,N_11594,N_11981);
xnor U13229 (N_13229,N_9056,N_9427);
nor U13230 (N_13230,N_11549,N_9418);
xor U13231 (N_13231,N_9584,N_11523);
nand U13232 (N_13232,N_11932,N_11207);
or U13233 (N_13233,N_11091,N_11651);
xor U13234 (N_13234,N_10479,N_9701);
nor U13235 (N_13235,N_11269,N_11126);
and U13236 (N_13236,N_9506,N_11395);
or U13237 (N_13237,N_10010,N_11957);
and U13238 (N_13238,N_10727,N_9698);
or U13239 (N_13239,N_9422,N_11996);
xnor U13240 (N_13240,N_10505,N_10162);
nor U13241 (N_13241,N_10624,N_10133);
and U13242 (N_13242,N_11992,N_9691);
nor U13243 (N_13243,N_11399,N_11912);
or U13244 (N_13244,N_11297,N_11928);
nand U13245 (N_13245,N_10903,N_9834);
nor U13246 (N_13246,N_11791,N_9406);
or U13247 (N_13247,N_9244,N_10991);
or U13248 (N_13248,N_9106,N_9557);
or U13249 (N_13249,N_9706,N_10940);
nor U13250 (N_13250,N_10312,N_10215);
xnor U13251 (N_13251,N_11930,N_10083);
and U13252 (N_13252,N_9375,N_11476);
and U13253 (N_13253,N_10368,N_9245);
nand U13254 (N_13254,N_9262,N_9602);
nand U13255 (N_13255,N_10061,N_9944);
and U13256 (N_13256,N_10829,N_10002);
xor U13257 (N_13257,N_11804,N_10112);
nand U13258 (N_13258,N_10143,N_10379);
xnor U13259 (N_13259,N_9250,N_9405);
or U13260 (N_13260,N_11086,N_11165);
or U13261 (N_13261,N_9256,N_10177);
or U13262 (N_13262,N_10073,N_9552);
and U13263 (N_13263,N_11728,N_11338);
or U13264 (N_13264,N_11892,N_11110);
or U13265 (N_13265,N_10778,N_11956);
nor U13266 (N_13266,N_10723,N_10319);
nand U13267 (N_13267,N_9420,N_10402);
nor U13268 (N_13268,N_10838,N_10332);
nor U13269 (N_13269,N_10718,N_10493);
nor U13270 (N_13270,N_10813,N_9239);
xnor U13271 (N_13271,N_10607,N_10531);
nand U13272 (N_13272,N_10600,N_9862);
nand U13273 (N_13273,N_9022,N_11375);
or U13274 (N_13274,N_11780,N_11509);
nor U13275 (N_13275,N_11821,N_9990);
and U13276 (N_13276,N_10548,N_10821);
and U13277 (N_13277,N_11443,N_9631);
xor U13278 (N_13278,N_9793,N_9128);
nor U13279 (N_13279,N_10593,N_11758);
and U13280 (N_13280,N_10328,N_10996);
nor U13281 (N_13281,N_11608,N_9947);
or U13282 (N_13282,N_11158,N_11723);
nand U13283 (N_13283,N_10107,N_10803);
or U13284 (N_13284,N_9211,N_11478);
nor U13285 (N_13285,N_11326,N_10249);
and U13286 (N_13286,N_9807,N_11559);
nor U13287 (N_13287,N_10169,N_10814);
nand U13288 (N_13288,N_10168,N_11442);
nand U13289 (N_13289,N_11063,N_9316);
nor U13290 (N_13290,N_11369,N_9379);
nand U13291 (N_13291,N_9240,N_11137);
and U13292 (N_13292,N_11688,N_10337);
and U13293 (N_13293,N_10476,N_9326);
nand U13294 (N_13294,N_10782,N_11754);
and U13295 (N_13295,N_9228,N_9199);
or U13296 (N_13296,N_11296,N_10563);
and U13297 (N_13297,N_9885,N_9194);
and U13298 (N_13298,N_10270,N_11087);
xnor U13299 (N_13299,N_11376,N_11187);
nand U13300 (N_13300,N_11950,N_10771);
or U13301 (N_13301,N_9175,N_9950);
nand U13302 (N_13302,N_10085,N_10053);
nor U13303 (N_13303,N_11637,N_9159);
nand U13304 (N_13304,N_10235,N_11434);
xor U13305 (N_13305,N_11342,N_9008);
or U13306 (N_13306,N_9573,N_11951);
and U13307 (N_13307,N_9259,N_10276);
and U13308 (N_13308,N_9503,N_10560);
and U13309 (N_13309,N_9629,N_10294);
nor U13310 (N_13310,N_10264,N_11292);
or U13311 (N_13311,N_9655,N_10879);
and U13312 (N_13312,N_10736,N_11265);
or U13313 (N_13313,N_9874,N_10557);
nand U13314 (N_13314,N_11572,N_11329);
nand U13315 (N_13315,N_10258,N_9880);
xnor U13316 (N_13316,N_11798,N_10523);
or U13317 (N_13317,N_10820,N_11839);
nand U13318 (N_13318,N_10852,N_11603);
xor U13319 (N_13319,N_11491,N_9572);
or U13320 (N_13320,N_11311,N_9498);
nor U13321 (N_13321,N_11106,N_9147);
xor U13322 (N_13322,N_9645,N_9089);
nor U13323 (N_13323,N_9961,N_11850);
or U13324 (N_13324,N_9450,N_10583);
nor U13325 (N_13325,N_11300,N_10038);
or U13326 (N_13326,N_11429,N_10305);
or U13327 (N_13327,N_10193,N_10060);
or U13328 (N_13328,N_10021,N_10387);
nor U13329 (N_13329,N_10105,N_10185);
nand U13330 (N_13330,N_11716,N_9087);
xor U13331 (N_13331,N_10149,N_9251);
nor U13332 (N_13332,N_10866,N_10571);
and U13333 (N_13333,N_9198,N_9529);
nor U13334 (N_13334,N_9209,N_11765);
xor U13335 (N_13335,N_9903,N_11561);
or U13336 (N_13336,N_10054,N_11436);
nor U13337 (N_13337,N_10116,N_9428);
and U13338 (N_13338,N_9971,N_9429);
nand U13339 (N_13339,N_10605,N_11556);
nand U13340 (N_13340,N_9088,N_11759);
nand U13341 (N_13341,N_9575,N_11666);
nor U13342 (N_13342,N_10020,N_10732);
or U13343 (N_13343,N_10655,N_11978);
nand U13344 (N_13344,N_10674,N_11935);
and U13345 (N_13345,N_11457,N_11710);
and U13346 (N_13346,N_10682,N_11764);
nor U13347 (N_13347,N_10891,N_9050);
and U13348 (N_13348,N_9296,N_10765);
and U13349 (N_13349,N_11906,N_11088);
nand U13350 (N_13350,N_11017,N_10904);
nor U13351 (N_13351,N_10619,N_9789);
or U13352 (N_13352,N_10819,N_9346);
nor U13353 (N_13353,N_9908,N_10393);
nor U13354 (N_13354,N_9169,N_11779);
xnor U13355 (N_13355,N_11103,N_11894);
and U13356 (N_13356,N_11368,N_10405);
nor U13357 (N_13357,N_9823,N_10544);
nand U13358 (N_13358,N_10383,N_11676);
and U13359 (N_13359,N_10934,N_10167);
or U13360 (N_13360,N_11315,N_9041);
xor U13361 (N_13361,N_10709,N_11312);
nand U13362 (N_13362,N_9226,N_9062);
nand U13363 (N_13363,N_11516,N_11153);
or U13364 (N_13364,N_10182,N_11220);
or U13365 (N_13365,N_11999,N_9505);
and U13366 (N_13366,N_11270,N_10353);
or U13367 (N_13367,N_10366,N_10568);
or U13368 (N_13368,N_10404,N_10603);
nor U13369 (N_13369,N_9449,N_10872);
or U13370 (N_13370,N_9031,N_11308);
and U13371 (N_13371,N_9002,N_11440);
or U13372 (N_13372,N_10184,N_10352);
nand U13373 (N_13373,N_11936,N_9597);
nor U13374 (N_13374,N_10477,N_9547);
and U13375 (N_13375,N_11298,N_9392);
and U13376 (N_13376,N_10556,N_11926);
xor U13377 (N_13377,N_11505,N_10487);
nand U13378 (N_13378,N_9934,N_9551);
and U13379 (N_13379,N_10868,N_11337);
nor U13380 (N_13380,N_10191,N_9443);
nand U13381 (N_13381,N_9319,N_11233);
or U13382 (N_13382,N_9314,N_11474);
nor U13383 (N_13383,N_11237,N_9308);
and U13384 (N_13384,N_9061,N_9887);
nor U13385 (N_13385,N_11173,N_9814);
xor U13386 (N_13386,N_9621,N_9985);
nor U13387 (N_13387,N_11896,N_11182);
or U13388 (N_13388,N_9322,N_10461);
and U13389 (N_13389,N_10914,N_10230);
or U13390 (N_13390,N_11336,N_10665);
and U13391 (N_13391,N_10640,N_9946);
nand U13392 (N_13392,N_9734,N_11101);
or U13393 (N_13393,N_9826,N_11445);
nor U13394 (N_13394,N_11389,N_9720);
nand U13395 (N_13395,N_10015,N_9713);
nor U13396 (N_13396,N_9423,N_10570);
and U13397 (N_13397,N_11404,N_10148);
or U13398 (N_13398,N_10440,N_10756);
or U13399 (N_13399,N_9276,N_11408);
nand U13400 (N_13400,N_9068,N_10562);
nand U13401 (N_13401,N_11554,N_9738);
or U13402 (N_13402,N_11011,N_11952);
or U13403 (N_13403,N_9865,N_10295);
or U13404 (N_13404,N_11350,N_9122);
xnor U13405 (N_13405,N_9455,N_10139);
nand U13406 (N_13406,N_10683,N_9756);
or U13407 (N_13407,N_10151,N_9771);
or U13408 (N_13408,N_10636,N_9753);
xor U13409 (N_13409,N_11468,N_10938);
and U13410 (N_13410,N_11525,N_10394);
and U13411 (N_13411,N_11622,N_10239);
and U13412 (N_13412,N_9453,N_9697);
and U13413 (N_13413,N_11960,N_11383);
or U13414 (N_13414,N_9515,N_10322);
nor U13415 (N_13415,N_10047,N_9905);
xor U13416 (N_13416,N_10130,N_10535);
xor U13417 (N_13417,N_11641,N_10661);
nor U13418 (N_13418,N_11690,N_10671);
or U13419 (N_13419,N_11497,N_10026);
and U13420 (N_13420,N_9842,N_9457);
nor U13421 (N_13421,N_10711,N_9580);
and U13422 (N_13422,N_9628,N_9225);
nand U13423 (N_13423,N_9688,N_10003);
xor U13424 (N_13424,N_11661,N_11630);
or U13425 (N_13425,N_11809,N_11610);
nor U13426 (N_13426,N_9499,N_9382);
and U13427 (N_13427,N_11890,N_11831);
and U13428 (N_13428,N_9635,N_11159);
or U13429 (N_13429,N_11028,N_10552);
nand U13430 (N_13430,N_10212,N_11854);
nand U13431 (N_13431,N_10877,N_9090);
nor U13432 (N_13432,N_10676,N_10409);
or U13433 (N_13433,N_11123,N_9029);
nand U13434 (N_13434,N_10032,N_9164);
nor U13435 (N_13435,N_9143,N_9795);
or U13436 (N_13436,N_9883,N_9117);
nor U13437 (N_13437,N_10797,N_11795);
or U13438 (N_13438,N_11845,N_10602);
and U13439 (N_13439,N_11899,N_9923);
or U13440 (N_13440,N_11618,N_9978);
nand U13441 (N_13441,N_9711,N_9282);
or U13442 (N_13442,N_10274,N_10410);
nand U13443 (N_13443,N_9608,N_9217);
xnor U13444 (N_13444,N_10874,N_10171);
and U13445 (N_13445,N_10375,N_11387);
nand U13446 (N_13446,N_11973,N_10284);
nand U13447 (N_13447,N_11555,N_11405);
nand U13448 (N_13448,N_9773,N_10344);
nand U13449 (N_13449,N_9246,N_11841);
or U13450 (N_13450,N_9130,N_9665);
and U13451 (N_13451,N_9491,N_10412);
and U13452 (N_13452,N_11527,N_9303);
or U13453 (N_13453,N_9092,N_11838);
and U13454 (N_13454,N_10865,N_10441);
nor U13455 (N_13455,N_10596,N_10099);
nor U13456 (N_13456,N_9586,N_10211);
xnor U13457 (N_13457,N_10045,N_11657);
and U13458 (N_13458,N_10816,N_11807);
xnor U13459 (N_13459,N_9113,N_10926);
nor U13460 (N_13460,N_9751,N_9539);
nor U13461 (N_13461,N_10564,N_9479);
and U13462 (N_13462,N_11059,N_9292);
nand U13463 (N_13463,N_9998,N_11100);
nor U13464 (N_13464,N_9593,N_11111);
or U13465 (N_13465,N_10918,N_9045);
nand U13466 (N_13466,N_10950,N_10530);
or U13467 (N_13467,N_9448,N_9715);
and U13468 (N_13468,N_9501,N_11763);
nor U13469 (N_13469,N_11859,N_11513);
or U13470 (N_13470,N_10898,N_9238);
or U13471 (N_13471,N_10431,N_10457);
nand U13472 (N_13472,N_9034,N_9366);
or U13473 (N_13473,N_9835,N_11319);
nand U13474 (N_13474,N_10932,N_9170);
or U13475 (N_13475,N_10527,N_11786);
nand U13476 (N_13476,N_9524,N_10121);
nand U13477 (N_13477,N_11607,N_9596);
or U13478 (N_13478,N_9941,N_10263);
or U13479 (N_13479,N_9532,N_11833);
nand U13480 (N_13480,N_9854,N_10800);
or U13481 (N_13481,N_9895,N_11615);
nand U13482 (N_13482,N_9230,N_11036);
nor U13483 (N_13483,N_10075,N_9146);
nand U13484 (N_13484,N_11242,N_11351);
nor U13485 (N_13485,N_9274,N_9731);
nor U13486 (N_13486,N_10882,N_10970);
nor U13487 (N_13487,N_11213,N_10974);
or U13488 (N_13488,N_10810,N_11781);
nor U13489 (N_13489,N_9868,N_9930);
nand U13490 (N_13490,N_11521,N_10894);
nand U13491 (N_13491,N_10302,N_9360);
or U13492 (N_13492,N_10992,N_10887);
nand U13493 (N_13493,N_11740,N_10242);
xnor U13494 (N_13494,N_10091,N_11132);
and U13495 (N_13495,N_10959,N_10386);
and U13496 (N_13496,N_10447,N_9656);
nor U13497 (N_13497,N_10156,N_11303);
or U13498 (N_13498,N_11542,N_9811);
xor U13499 (N_13499,N_10190,N_10515);
nand U13500 (N_13500,N_9043,N_9982);
nand U13501 (N_13501,N_10294,N_11757);
and U13502 (N_13502,N_9051,N_10247);
nand U13503 (N_13503,N_9353,N_11922);
nand U13504 (N_13504,N_11125,N_10439);
nand U13505 (N_13505,N_9123,N_9654);
xnor U13506 (N_13506,N_11721,N_10367);
nor U13507 (N_13507,N_11721,N_9458);
nor U13508 (N_13508,N_10125,N_9419);
and U13509 (N_13509,N_9758,N_9472);
nor U13510 (N_13510,N_10005,N_11941);
and U13511 (N_13511,N_9770,N_10855);
nand U13512 (N_13512,N_10333,N_11278);
nor U13513 (N_13513,N_10378,N_11427);
nand U13514 (N_13514,N_10172,N_9731);
and U13515 (N_13515,N_10172,N_10880);
and U13516 (N_13516,N_9838,N_9615);
xor U13517 (N_13517,N_10770,N_9704);
or U13518 (N_13518,N_11658,N_11385);
and U13519 (N_13519,N_10842,N_11235);
or U13520 (N_13520,N_9265,N_11476);
nor U13521 (N_13521,N_9118,N_11159);
xor U13522 (N_13522,N_9792,N_9977);
nand U13523 (N_13523,N_11681,N_9924);
or U13524 (N_13524,N_10855,N_10421);
nand U13525 (N_13525,N_11044,N_10583);
or U13526 (N_13526,N_10021,N_9562);
nor U13527 (N_13527,N_11917,N_9921);
nand U13528 (N_13528,N_10348,N_9229);
or U13529 (N_13529,N_10787,N_9947);
xnor U13530 (N_13530,N_9950,N_9906);
and U13531 (N_13531,N_10005,N_9196);
nor U13532 (N_13532,N_11532,N_10063);
or U13533 (N_13533,N_9798,N_9844);
and U13534 (N_13534,N_11266,N_11267);
or U13535 (N_13535,N_9333,N_11631);
or U13536 (N_13536,N_10153,N_11478);
nor U13537 (N_13537,N_9259,N_10701);
nand U13538 (N_13538,N_9922,N_10091);
xnor U13539 (N_13539,N_11511,N_11988);
or U13540 (N_13540,N_9190,N_10199);
and U13541 (N_13541,N_9284,N_10104);
and U13542 (N_13542,N_9721,N_10531);
or U13543 (N_13543,N_11319,N_10595);
or U13544 (N_13544,N_10692,N_11128);
and U13545 (N_13545,N_11235,N_9735);
nand U13546 (N_13546,N_11155,N_10974);
or U13547 (N_13547,N_9821,N_10628);
and U13548 (N_13548,N_11908,N_9526);
or U13549 (N_13549,N_10619,N_9223);
nand U13550 (N_13550,N_9994,N_9971);
and U13551 (N_13551,N_9387,N_9514);
nor U13552 (N_13552,N_11292,N_9048);
and U13553 (N_13553,N_10781,N_9857);
nor U13554 (N_13554,N_11611,N_9218);
and U13555 (N_13555,N_10186,N_10678);
or U13556 (N_13556,N_11311,N_10844);
and U13557 (N_13557,N_10060,N_9118);
and U13558 (N_13558,N_10590,N_11633);
and U13559 (N_13559,N_11057,N_9362);
nor U13560 (N_13560,N_9581,N_11380);
nor U13561 (N_13561,N_9792,N_9887);
nand U13562 (N_13562,N_10041,N_10402);
or U13563 (N_13563,N_9356,N_9585);
or U13564 (N_13564,N_9081,N_11141);
xor U13565 (N_13565,N_11285,N_11865);
nand U13566 (N_13566,N_9807,N_10139);
xnor U13567 (N_13567,N_11556,N_11896);
nand U13568 (N_13568,N_9299,N_10933);
and U13569 (N_13569,N_9797,N_11548);
nand U13570 (N_13570,N_9991,N_10215);
nand U13571 (N_13571,N_11502,N_9258);
and U13572 (N_13572,N_9116,N_10092);
nor U13573 (N_13573,N_9019,N_11469);
and U13574 (N_13574,N_9439,N_11746);
or U13575 (N_13575,N_10325,N_10869);
nand U13576 (N_13576,N_10742,N_10758);
nor U13577 (N_13577,N_9712,N_10894);
and U13578 (N_13578,N_9467,N_11703);
xnor U13579 (N_13579,N_10009,N_9573);
nor U13580 (N_13580,N_10386,N_10821);
nand U13581 (N_13581,N_10834,N_9079);
nand U13582 (N_13582,N_10991,N_10345);
nand U13583 (N_13583,N_9666,N_11967);
nor U13584 (N_13584,N_11087,N_9890);
nor U13585 (N_13585,N_11481,N_11371);
nor U13586 (N_13586,N_10906,N_11689);
or U13587 (N_13587,N_9932,N_11463);
or U13588 (N_13588,N_9526,N_9528);
nor U13589 (N_13589,N_11958,N_10611);
xnor U13590 (N_13590,N_10100,N_11657);
and U13591 (N_13591,N_9781,N_9819);
or U13592 (N_13592,N_10750,N_9991);
and U13593 (N_13593,N_10755,N_9269);
nand U13594 (N_13594,N_11733,N_9079);
or U13595 (N_13595,N_9803,N_10000);
or U13596 (N_13596,N_11724,N_10910);
or U13597 (N_13597,N_10425,N_9619);
or U13598 (N_13598,N_10645,N_9705);
and U13599 (N_13599,N_9929,N_11825);
nand U13600 (N_13600,N_9806,N_11830);
or U13601 (N_13601,N_9972,N_9979);
nor U13602 (N_13602,N_9321,N_11719);
xnor U13603 (N_13603,N_10056,N_10654);
xnor U13604 (N_13604,N_11189,N_9271);
nor U13605 (N_13605,N_11567,N_11471);
nand U13606 (N_13606,N_10843,N_11500);
xor U13607 (N_13607,N_9442,N_10808);
nand U13608 (N_13608,N_10634,N_11576);
nor U13609 (N_13609,N_9420,N_11295);
nand U13610 (N_13610,N_10964,N_11842);
nand U13611 (N_13611,N_9878,N_9831);
nor U13612 (N_13612,N_11486,N_11753);
or U13613 (N_13613,N_11108,N_10498);
nor U13614 (N_13614,N_9441,N_9460);
nand U13615 (N_13615,N_10837,N_11626);
xor U13616 (N_13616,N_10135,N_10618);
or U13617 (N_13617,N_11913,N_10315);
nor U13618 (N_13618,N_10350,N_10544);
or U13619 (N_13619,N_10097,N_11457);
nor U13620 (N_13620,N_10610,N_11214);
and U13621 (N_13621,N_9082,N_10415);
and U13622 (N_13622,N_9961,N_9035);
nor U13623 (N_13623,N_10574,N_9090);
xor U13624 (N_13624,N_9081,N_11906);
and U13625 (N_13625,N_11111,N_9570);
or U13626 (N_13626,N_10898,N_10039);
nand U13627 (N_13627,N_9901,N_9030);
or U13628 (N_13628,N_9809,N_10045);
xor U13629 (N_13629,N_11890,N_11841);
nor U13630 (N_13630,N_10162,N_10472);
xor U13631 (N_13631,N_9605,N_10372);
or U13632 (N_13632,N_9719,N_10677);
nand U13633 (N_13633,N_9317,N_10020);
or U13634 (N_13634,N_9257,N_10625);
and U13635 (N_13635,N_10800,N_9644);
or U13636 (N_13636,N_11292,N_9496);
nand U13637 (N_13637,N_9060,N_11033);
nor U13638 (N_13638,N_11384,N_11154);
xnor U13639 (N_13639,N_10620,N_11992);
nand U13640 (N_13640,N_11093,N_10794);
or U13641 (N_13641,N_9920,N_10780);
and U13642 (N_13642,N_9467,N_11903);
or U13643 (N_13643,N_9023,N_11048);
nand U13644 (N_13644,N_9719,N_10019);
or U13645 (N_13645,N_10487,N_9374);
nor U13646 (N_13646,N_11018,N_9385);
or U13647 (N_13647,N_11783,N_9495);
nand U13648 (N_13648,N_11990,N_9676);
nand U13649 (N_13649,N_10256,N_9557);
or U13650 (N_13650,N_10470,N_11298);
nand U13651 (N_13651,N_10616,N_10975);
nor U13652 (N_13652,N_9389,N_10666);
nand U13653 (N_13653,N_11163,N_11828);
xor U13654 (N_13654,N_10865,N_11553);
or U13655 (N_13655,N_10138,N_11857);
or U13656 (N_13656,N_9487,N_11812);
nor U13657 (N_13657,N_10879,N_10708);
nand U13658 (N_13658,N_11504,N_10366);
xnor U13659 (N_13659,N_11573,N_9417);
nor U13660 (N_13660,N_10327,N_9748);
nand U13661 (N_13661,N_11422,N_11806);
nand U13662 (N_13662,N_9050,N_9193);
xor U13663 (N_13663,N_11313,N_10740);
and U13664 (N_13664,N_10223,N_11710);
or U13665 (N_13665,N_11642,N_10992);
and U13666 (N_13666,N_10943,N_10691);
nor U13667 (N_13667,N_9056,N_11359);
nor U13668 (N_13668,N_9953,N_9600);
and U13669 (N_13669,N_10532,N_10452);
and U13670 (N_13670,N_10814,N_10084);
nor U13671 (N_13671,N_9917,N_10051);
or U13672 (N_13672,N_10099,N_10959);
xnor U13673 (N_13673,N_9704,N_10773);
nand U13674 (N_13674,N_9403,N_10942);
and U13675 (N_13675,N_10282,N_11968);
or U13676 (N_13676,N_11939,N_11617);
nor U13677 (N_13677,N_11337,N_9361);
nand U13678 (N_13678,N_9720,N_11274);
or U13679 (N_13679,N_9522,N_9460);
nor U13680 (N_13680,N_11148,N_10383);
and U13681 (N_13681,N_10971,N_10563);
and U13682 (N_13682,N_10274,N_11674);
xnor U13683 (N_13683,N_9365,N_10964);
or U13684 (N_13684,N_9926,N_11472);
or U13685 (N_13685,N_11924,N_9765);
nand U13686 (N_13686,N_9450,N_9988);
xor U13687 (N_13687,N_10070,N_11741);
nand U13688 (N_13688,N_11242,N_11887);
and U13689 (N_13689,N_10758,N_9826);
nand U13690 (N_13690,N_11155,N_11329);
nor U13691 (N_13691,N_11546,N_11493);
nor U13692 (N_13692,N_11057,N_10316);
nand U13693 (N_13693,N_9712,N_11663);
nor U13694 (N_13694,N_11597,N_10193);
nand U13695 (N_13695,N_11567,N_10845);
nor U13696 (N_13696,N_9972,N_11024);
nor U13697 (N_13697,N_11709,N_10291);
nand U13698 (N_13698,N_10113,N_9883);
nand U13699 (N_13699,N_11084,N_11414);
nand U13700 (N_13700,N_10409,N_10723);
nand U13701 (N_13701,N_11181,N_9374);
or U13702 (N_13702,N_10656,N_10990);
or U13703 (N_13703,N_9184,N_10062);
xnor U13704 (N_13704,N_10522,N_9762);
or U13705 (N_13705,N_9707,N_10864);
xor U13706 (N_13706,N_10719,N_9123);
xor U13707 (N_13707,N_10621,N_11921);
or U13708 (N_13708,N_11150,N_9587);
and U13709 (N_13709,N_9593,N_9054);
nor U13710 (N_13710,N_9893,N_9637);
or U13711 (N_13711,N_9383,N_9912);
or U13712 (N_13712,N_11824,N_11518);
nand U13713 (N_13713,N_10942,N_9363);
nor U13714 (N_13714,N_11745,N_9106);
nand U13715 (N_13715,N_9898,N_9957);
and U13716 (N_13716,N_9089,N_11534);
xor U13717 (N_13717,N_11520,N_10990);
or U13718 (N_13718,N_10552,N_10037);
xnor U13719 (N_13719,N_10278,N_9662);
nor U13720 (N_13720,N_9599,N_11875);
and U13721 (N_13721,N_10521,N_10006);
nand U13722 (N_13722,N_9892,N_9367);
or U13723 (N_13723,N_10891,N_9163);
nor U13724 (N_13724,N_11441,N_9024);
or U13725 (N_13725,N_11469,N_9084);
or U13726 (N_13726,N_11765,N_10629);
nor U13727 (N_13727,N_10368,N_9019);
xor U13728 (N_13728,N_9276,N_10323);
or U13729 (N_13729,N_10912,N_9594);
or U13730 (N_13730,N_11564,N_11498);
nand U13731 (N_13731,N_11330,N_10169);
or U13732 (N_13732,N_9339,N_10679);
nand U13733 (N_13733,N_10449,N_11421);
and U13734 (N_13734,N_9224,N_9300);
and U13735 (N_13735,N_11873,N_9614);
or U13736 (N_13736,N_10355,N_11465);
nand U13737 (N_13737,N_11886,N_11623);
nor U13738 (N_13738,N_11273,N_9587);
and U13739 (N_13739,N_11998,N_10398);
nand U13740 (N_13740,N_11146,N_10668);
nand U13741 (N_13741,N_11346,N_11993);
nor U13742 (N_13742,N_9591,N_9102);
nand U13743 (N_13743,N_11727,N_9012);
nor U13744 (N_13744,N_11571,N_9382);
nor U13745 (N_13745,N_9425,N_11335);
nand U13746 (N_13746,N_9284,N_11278);
nand U13747 (N_13747,N_11967,N_11413);
nand U13748 (N_13748,N_11906,N_9172);
or U13749 (N_13749,N_9991,N_9830);
nor U13750 (N_13750,N_9751,N_9968);
and U13751 (N_13751,N_9064,N_10978);
or U13752 (N_13752,N_11573,N_11348);
and U13753 (N_13753,N_9376,N_11616);
and U13754 (N_13754,N_9272,N_11597);
and U13755 (N_13755,N_9943,N_11838);
xnor U13756 (N_13756,N_9064,N_9013);
and U13757 (N_13757,N_11297,N_9930);
and U13758 (N_13758,N_11357,N_11514);
nand U13759 (N_13759,N_10230,N_9320);
xor U13760 (N_13760,N_10710,N_10808);
nor U13761 (N_13761,N_11946,N_9222);
or U13762 (N_13762,N_11432,N_9184);
nand U13763 (N_13763,N_11973,N_9622);
or U13764 (N_13764,N_11957,N_11854);
nand U13765 (N_13765,N_10408,N_10015);
nor U13766 (N_13766,N_9216,N_10336);
and U13767 (N_13767,N_10801,N_10258);
and U13768 (N_13768,N_10742,N_11970);
xor U13769 (N_13769,N_9151,N_10742);
and U13770 (N_13770,N_9321,N_9015);
xnor U13771 (N_13771,N_11552,N_11247);
nand U13772 (N_13772,N_11513,N_10295);
nor U13773 (N_13773,N_10600,N_11056);
or U13774 (N_13774,N_10941,N_9094);
nand U13775 (N_13775,N_10573,N_10630);
nor U13776 (N_13776,N_10824,N_10036);
nor U13777 (N_13777,N_11300,N_11703);
xnor U13778 (N_13778,N_10446,N_10872);
or U13779 (N_13779,N_11056,N_10722);
and U13780 (N_13780,N_9302,N_10017);
nor U13781 (N_13781,N_10325,N_10335);
or U13782 (N_13782,N_10481,N_10548);
and U13783 (N_13783,N_11874,N_11462);
nand U13784 (N_13784,N_11217,N_10147);
and U13785 (N_13785,N_9639,N_11809);
nand U13786 (N_13786,N_11966,N_9953);
and U13787 (N_13787,N_11267,N_11015);
and U13788 (N_13788,N_11460,N_10476);
nand U13789 (N_13789,N_11036,N_11190);
and U13790 (N_13790,N_10492,N_11568);
or U13791 (N_13791,N_10422,N_11396);
and U13792 (N_13792,N_11378,N_11534);
xor U13793 (N_13793,N_9821,N_9089);
and U13794 (N_13794,N_10278,N_9533);
nand U13795 (N_13795,N_9232,N_11529);
nor U13796 (N_13796,N_10270,N_10819);
nand U13797 (N_13797,N_9740,N_11748);
nand U13798 (N_13798,N_11026,N_10630);
xnor U13799 (N_13799,N_10495,N_10800);
or U13800 (N_13800,N_10483,N_9248);
nor U13801 (N_13801,N_11221,N_10272);
nor U13802 (N_13802,N_9641,N_11180);
and U13803 (N_13803,N_11447,N_11244);
and U13804 (N_13804,N_10470,N_11682);
or U13805 (N_13805,N_9564,N_11490);
or U13806 (N_13806,N_9683,N_10042);
nand U13807 (N_13807,N_10773,N_9461);
xor U13808 (N_13808,N_10367,N_11416);
or U13809 (N_13809,N_10448,N_11589);
or U13810 (N_13810,N_10770,N_9541);
or U13811 (N_13811,N_10997,N_11607);
nand U13812 (N_13812,N_11242,N_10565);
or U13813 (N_13813,N_11144,N_10350);
and U13814 (N_13814,N_11819,N_11536);
nand U13815 (N_13815,N_11947,N_9368);
nor U13816 (N_13816,N_10474,N_9118);
nand U13817 (N_13817,N_11138,N_11451);
nand U13818 (N_13818,N_9260,N_10377);
and U13819 (N_13819,N_9336,N_9538);
or U13820 (N_13820,N_11057,N_10927);
and U13821 (N_13821,N_10080,N_9662);
and U13822 (N_13822,N_9822,N_9861);
nor U13823 (N_13823,N_10380,N_10643);
or U13824 (N_13824,N_10088,N_11677);
or U13825 (N_13825,N_9192,N_11391);
or U13826 (N_13826,N_10592,N_11909);
and U13827 (N_13827,N_9874,N_10493);
and U13828 (N_13828,N_11790,N_11330);
nand U13829 (N_13829,N_11492,N_10533);
nand U13830 (N_13830,N_10565,N_10100);
nand U13831 (N_13831,N_9073,N_10992);
or U13832 (N_13832,N_9842,N_10849);
and U13833 (N_13833,N_11697,N_10085);
and U13834 (N_13834,N_9375,N_11932);
or U13835 (N_13835,N_9064,N_10620);
xnor U13836 (N_13836,N_9950,N_9593);
xnor U13837 (N_13837,N_9638,N_9502);
or U13838 (N_13838,N_11752,N_11324);
or U13839 (N_13839,N_9969,N_11277);
nor U13840 (N_13840,N_10801,N_11172);
nor U13841 (N_13841,N_11437,N_10020);
nor U13842 (N_13842,N_11100,N_10358);
nand U13843 (N_13843,N_9765,N_10433);
nand U13844 (N_13844,N_10938,N_10985);
nand U13845 (N_13845,N_10344,N_9199);
or U13846 (N_13846,N_11549,N_10738);
or U13847 (N_13847,N_10386,N_10435);
nand U13848 (N_13848,N_10202,N_9218);
and U13849 (N_13849,N_10007,N_10446);
and U13850 (N_13850,N_10877,N_11267);
or U13851 (N_13851,N_11317,N_9629);
or U13852 (N_13852,N_10982,N_11750);
and U13853 (N_13853,N_9401,N_9581);
nor U13854 (N_13854,N_9442,N_9660);
nand U13855 (N_13855,N_10979,N_10022);
and U13856 (N_13856,N_10085,N_10958);
xnor U13857 (N_13857,N_11694,N_10187);
or U13858 (N_13858,N_9255,N_11446);
and U13859 (N_13859,N_10982,N_9592);
xnor U13860 (N_13860,N_9647,N_11367);
and U13861 (N_13861,N_10246,N_11428);
and U13862 (N_13862,N_11620,N_10865);
xor U13863 (N_13863,N_10039,N_9886);
nand U13864 (N_13864,N_11292,N_11003);
and U13865 (N_13865,N_10934,N_11496);
nor U13866 (N_13866,N_9655,N_11726);
xnor U13867 (N_13867,N_11391,N_11477);
nor U13868 (N_13868,N_9437,N_11616);
nand U13869 (N_13869,N_11332,N_9605);
nor U13870 (N_13870,N_11100,N_11689);
nor U13871 (N_13871,N_10055,N_11310);
nand U13872 (N_13872,N_11185,N_9143);
nor U13873 (N_13873,N_9570,N_11283);
and U13874 (N_13874,N_9389,N_10862);
nand U13875 (N_13875,N_9391,N_11788);
or U13876 (N_13876,N_9205,N_10821);
and U13877 (N_13877,N_11195,N_9797);
or U13878 (N_13878,N_9032,N_10263);
or U13879 (N_13879,N_10102,N_9332);
nand U13880 (N_13880,N_11360,N_11973);
xnor U13881 (N_13881,N_9562,N_11457);
and U13882 (N_13882,N_11532,N_10504);
xnor U13883 (N_13883,N_10344,N_9793);
nor U13884 (N_13884,N_9630,N_11847);
xor U13885 (N_13885,N_9942,N_9204);
xor U13886 (N_13886,N_11657,N_11438);
nor U13887 (N_13887,N_10709,N_11054);
or U13888 (N_13888,N_11609,N_11713);
nand U13889 (N_13889,N_11756,N_10634);
nor U13890 (N_13890,N_10048,N_11891);
and U13891 (N_13891,N_9161,N_10672);
nor U13892 (N_13892,N_11926,N_9486);
nand U13893 (N_13893,N_9579,N_9537);
xnor U13894 (N_13894,N_9571,N_11558);
xor U13895 (N_13895,N_9764,N_9458);
xor U13896 (N_13896,N_11062,N_9229);
or U13897 (N_13897,N_11059,N_11510);
nand U13898 (N_13898,N_9019,N_11093);
or U13899 (N_13899,N_10408,N_10264);
xor U13900 (N_13900,N_11053,N_9051);
or U13901 (N_13901,N_9485,N_10800);
nor U13902 (N_13902,N_11168,N_10520);
or U13903 (N_13903,N_11532,N_10551);
nand U13904 (N_13904,N_9665,N_10815);
xnor U13905 (N_13905,N_9738,N_11272);
nor U13906 (N_13906,N_11978,N_9280);
or U13907 (N_13907,N_11219,N_10887);
nor U13908 (N_13908,N_11843,N_10758);
xnor U13909 (N_13909,N_11213,N_9779);
nand U13910 (N_13910,N_10210,N_11751);
xor U13911 (N_13911,N_10030,N_9545);
nand U13912 (N_13912,N_9136,N_9633);
or U13913 (N_13913,N_10165,N_11911);
and U13914 (N_13914,N_9480,N_10453);
nand U13915 (N_13915,N_11401,N_9472);
nor U13916 (N_13916,N_11692,N_9442);
or U13917 (N_13917,N_11587,N_9360);
nor U13918 (N_13918,N_11790,N_11913);
nor U13919 (N_13919,N_10307,N_9460);
or U13920 (N_13920,N_10851,N_9262);
nand U13921 (N_13921,N_10394,N_9641);
nand U13922 (N_13922,N_10830,N_10338);
xor U13923 (N_13923,N_9785,N_9376);
and U13924 (N_13924,N_10778,N_10031);
xnor U13925 (N_13925,N_10452,N_9696);
and U13926 (N_13926,N_9307,N_9550);
xor U13927 (N_13927,N_10121,N_10207);
nor U13928 (N_13928,N_10705,N_9729);
or U13929 (N_13929,N_9444,N_11223);
and U13930 (N_13930,N_10622,N_10693);
nor U13931 (N_13931,N_11576,N_9055);
nand U13932 (N_13932,N_11065,N_10567);
xnor U13933 (N_13933,N_11163,N_10592);
nor U13934 (N_13934,N_10025,N_9207);
nor U13935 (N_13935,N_10023,N_9614);
nor U13936 (N_13936,N_9906,N_10241);
nor U13937 (N_13937,N_10670,N_11780);
or U13938 (N_13938,N_9499,N_11978);
and U13939 (N_13939,N_10368,N_10466);
or U13940 (N_13940,N_10573,N_11089);
nor U13941 (N_13941,N_9840,N_9552);
nand U13942 (N_13942,N_9814,N_9858);
and U13943 (N_13943,N_10251,N_11995);
nand U13944 (N_13944,N_9953,N_9365);
or U13945 (N_13945,N_9759,N_9988);
nand U13946 (N_13946,N_9261,N_10410);
and U13947 (N_13947,N_9726,N_10268);
and U13948 (N_13948,N_9192,N_10353);
or U13949 (N_13949,N_9545,N_11005);
nand U13950 (N_13950,N_10649,N_10472);
xor U13951 (N_13951,N_9292,N_11155);
and U13952 (N_13952,N_11926,N_10992);
and U13953 (N_13953,N_10856,N_10291);
or U13954 (N_13954,N_9847,N_11854);
and U13955 (N_13955,N_11504,N_9436);
and U13956 (N_13956,N_11532,N_10553);
and U13957 (N_13957,N_11758,N_11461);
xor U13958 (N_13958,N_11942,N_10111);
nand U13959 (N_13959,N_10202,N_10552);
and U13960 (N_13960,N_9044,N_11205);
and U13961 (N_13961,N_9868,N_10559);
nor U13962 (N_13962,N_11129,N_9172);
nor U13963 (N_13963,N_9737,N_11055);
or U13964 (N_13964,N_11946,N_11840);
nand U13965 (N_13965,N_10431,N_10385);
nor U13966 (N_13966,N_10884,N_11388);
nor U13967 (N_13967,N_10446,N_10197);
and U13968 (N_13968,N_9025,N_9469);
and U13969 (N_13969,N_11056,N_10055);
nand U13970 (N_13970,N_10862,N_9894);
and U13971 (N_13971,N_11954,N_10443);
nor U13972 (N_13972,N_10403,N_10050);
or U13973 (N_13973,N_11381,N_11936);
nand U13974 (N_13974,N_9605,N_10858);
and U13975 (N_13975,N_11823,N_10661);
or U13976 (N_13976,N_10229,N_11601);
or U13977 (N_13977,N_10007,N_11526);
or U13978 (N_13978,N_9560,N_10946);
nand U13979 (N_13979,N_9058,N_10941);
and U13980 (N_13980,N_11088,N_9209);
nand U13981 (N_13981,N_9029,N_9099);
and U13982 (N_13982,N_11230,N_11718);
or U13983 (N_13983,N_10872,N_11679);
nor U13984 (N_13984,N_10273,N_11272);
and U13985 (N_13985,N_10098,N_9996);
and U13986 (N_13986,N_11951,N_9511);
nor U13987 (N_13987,N_11349,N_9988);
nor U13988 (N_13988,N_10090,N_10304);
or U13989 (N_13989,N_11132,N_10301);
nand U13990 (N_13990,N_10085,N_11126);
nor U13991 (N_13991,N_9469,N_9017);
nor U13992 (N_13992,N_10004,N_9708);
and U13993 (N_13993,N_10247,N_11870);
xor U13994 (N_13994,N_9869,N_9484);
and U13995 (N_13995,N_10501,N_10432);
nand U13996 (N_13996,N_10796,N_10753);
nor U13997 (N_13997,N_11494,N_9923);
nor U13998 (N_13998,N_9359,N_11422);
and U13999 (N_13999,N_9867,N_11898);
nor U14000 (N_14000,N_10651,N_10889);
nand U14001 (N_14001,N_9699,N_9457);
or U14002 (N_14002,N_11408,N_10499);
nor U14003 (N_14003,N_11414,N_10067);
nor U14004 (N_14004,N_10432,N_9174);
and U14005 (N_14005,N_10095,N_9787);
nor U14006 (N_14006,N_11328,N_9464);
nor U14007 (N_14007,N_9962,N_11755);
nor U14008 (N_14008,N_10747,N_9716);
nand U14009 (N_14009,N_11837,N_11168);
and U14010 (N_14010,N_11617,N_11703);
or U14011 (N_14011,N_11463,N_9468);
or U14012 (N_14012,N_9746,N_9749);
and U14013 (N_14013,N_10706,N_9576);
and U14014 (N_14014,N_9313,N_9272);
or U14015 (N_14015,N_9830,N_10429);
and U14016 (N_14016,N_11874,N_9789);
nand U14017 (N_14017,N_11979,N_11633);
nor U14018 (N_14018,N_10353,N_10703);
and U14019 (N_14019,N_9213,N_11126);
xnor U14020 (N_14020,N_10404,N_9265);
and U14021 (N_14021,N_10740,N_10830);
nor U14022 (N_14022,N_9717,N_11366);
nor U14023 (N_14023,N_11627,N_10715);
nand U14024 (N_14024,N_11464,N_11501);
and U14025 (N_14025,N_9510,N_10730);
nor U14026 (N_14026,N_10185,N_11832);
and U14027 (N_14027,N_11338,N_9090);
nor U14028 (N_14028,N_11819,N_10764);
nand U14029 (N_14029,N_10464,N_10726);
nand U14030 (N_14030,N_9879,N_10142);
and U14031 (N_14031,N_11634,N_10576);
xnor U14032 (N_14032,N_10572,N_10429);
or U14033 (N_14033,N_9537,N_10901);
and U14034 (N_14034,N_11264,N_9575);
or U14035 (N_14035,N_10817,N_10324);
nand U14036 (N_14036,N_10074,N_10927);
and U14037 (N_14037,N_11346,N_10943);
xor U14038 (N_14038,N_10044,N_11064);
nor U14039 (N_14039,N_10401,N_9767);
xor U14040 (N_14040,N_11127,N_9808);
nand U14041 (N_14041,N_11022,N_11900);
and U14042 (N_14042,N_9188,N_11970);
or U14043 (N_14043,N_9027,N_9337);
or U14044 (N_14044,N_9915,N_9805);
nand U14045 (N_14045,N_10328,N_11477);
nor U14046 (N_14046,N_11453,N_11074);
and U14047 (N_14047,N_11419,N_11307);
nor U14048 (N_14048,N_10345,N_11836);
or U14049 (N_14049,N_10418,N_10649);
xnor U14050 (N_14050,N_10853,N_10420);
and U14051 (N_14051,N_10105,N_10838);
and U14052 (N_14052,N_11192,N_9556);
nand U14053 (N_14053,N_11876,N_10509);
nand U14054 (N_14054,N_10290,N_10790);
nor U14055 (N_14055,N_11124,N_9652);
nand U14056 (N_14056,N_11519,N_10856);
nand U14057 (N_14057,N_11561,N_9964);
nor U14058 (N_14058,N_11738,N_10257);
nor U14059 (N_14059,N_10554,N_10783);
nand U14060 (N_14060,N_9021,N_9449);
xnor U14061 (N_14061,N_10607,N_9592);
nand U14062 (N_14062,N_11079,N_10078);
or U14063 (N_14063,N_10217,N_11994);
or U14064 (N_14064,N_9302,N_10316);
nor U14065 (N_14065,N_9867,N_11064);
nand U14066 (N_14066,N_11711,N_9184);
and U14067 (N_14067,N_11866,N_11916);
or U14068 (N_14068,N_9173,N_11443);
or U14069 (N_14069,N_10732,N_9139);
nor U14070 (N_14070,N_9861,N_9271);
xnor U14071 (N_14071,N_9621,N_11260);
nand U14072 (N_14072,N_9583,N_9444);
or U14073 (N_14073,N_9653,N_10941);
nor U14074 (N_14074,N_10036,N_10097);
and U14075 (N_14075,N_11128,N_11297);
nand U14076 (N_14076,N_11291,N_10141);
and U14077 (N_14077,N_11180,N_9610);
or U14078 (N_14078,N_9192,N_11893);
nand U14079 (N_14079,N_9357,N_11555);
xnor U14080 (N_14080,N_10437,N_11513);
nor U14081 (N_14081,N_9757,N_9932);
and U14082 (N_14082,N_9114,N_11057);
nor U14083 (N_14083,N_9749,N_10953);
and U14084 (N_14084,N_9486,N_11241);
nand U14085 (N_14085,N_11948,N_10314);
and U14086 (N_14086,N_10169,N_9164);
nand U14087 (N_14087,N_9979,N_9516);
or U14088 (N_14088,N_11685,N_9491);
or U14089 (N_14089,N_11051,N_10792);
nor U14090 (N_14090,N_11292,N_10814);
and U14091 (N_14091,N_9452,N_11129);
and U14092 (N_14092,N_11721,N_11212);
and U14093 (N_14093,N_10837,N_9952);
nor U14094 (N_14094,N_11171,N_10235);
nor U14095 (N_14095,N_9228,N_11662);
nand U14096 (N_14096,N_10177,N_9100);
or U14097 (N_14097,N_9053,N_11741);
xor U14098 (N_14098,N_9662,N_9374);
or U14099 (N_14099,N_10968,N_10296);
and U14100 (N_14100,N_9281,N_11074);
nand U14101 (N_14101,N_10579,N_10852);
nor U14102 (N_14102,N_10747,N_11230);
nand U14103 (N_14103,N_9990,N_11433);
and U14104 (N_14104,N_11203,N_10497);
nand U14105 (N_14105,N_9001,N_10540);
xor U14106 (N_14106,N_10627,N_9660);
nor U14107 (N_14107,N_10320,N_10937);
nor U14108 (N_14108,N_9510,N_10799);
or U14109 (N_14109,N_9083,N_9255);
or U14110 (N_14110,N_11208,N_11406);
or U14111 (N_14111,N_10360,N_9134);
nor U14112 (N_14112,N_10734,N_9965);
and U14113 (N_14113,N_11176,N_10442);
nand U14114 (N_14114,N_9932,N_10147);
or U14115 (N_14115,N_11091,N_11632);
or U14116 (N_14116,N_10612,N_9429);
nor U14117 (N_14117,N_9521,N_10385);
and U14118 (N_14118,N_11630,N_11489);
nand U14119 (N_14119,N_10472,N_9826);
nor U14120 (N_14120,N_10628,N_9391);
and U14121 (N_14121,N_10524,N_11117);
or U14122 (N_14122,N_10319,N_10861);
nor U14123 (N_14123,N_9395,N_11141);
xor U14124 (N_14124,N_11956,N_9696);
and U14125 (N_14125,N_9610,N_9961);
nand U14126 (N_14126,N_11056,N_10094);
and U14127 (N_14127,N_10325,N_11107);
nor U14128 (N_14128,N_11463,N_9120);
and U14129 (N_14129,N_10203,N_10201);
nor U14130 (N_14130,N_11543,N_10082);
and U14131 (N_14131,N_11431,N_10886);
or U14132 (N_14132,N_11415,N_10219);
nand U14133 (N_14133,N_11383,N_11948);
or U14134 (N_14134,N_9943,N_9892);
nand U14135 (N_14135,N_9553,N_9029);
nor U14136 (N_14136,N_11576,N_11424);
xor U14137 (N_14137,N_9662,N_10283);
or U14138 (N_14138,N_10368,N_11609);
and U14139 (N_14139,N_9886,N_10298);
nand U14140 (N_14140,N_9822,N_10421);
or U14141 (N_14141,N_11670,N_9715);
nand U14142 (N_14142,N_9828,N_10995);
or U14143 (N_14143,N_10857,N_11254);
nor U14144 (N_14144,N_10111,N_10328);
nand U14145 (N_14145,N_9323,N_11043);
and U14146 (N_14146,N_9941,N_11907);
and U14147 (N_14147,N_10301,N_9167);
or U14148 (N_14148,N_9750,N_10897);
nor U14149 (N_14149,N_10802,N_9936);
nor U14150 (N_14150,N_9527,N_11662);
or U14151 (N_14151,N_11387,N_10812);
and U14152 (N_14152,N_11398,N_10126);
or U14153 (N_14153,N_10748,N_10599);
or U14154 (N_14154,N_9898,N_9634);
or U14155 (N_14155,N_11603,N_10468);
and U14156 (N_14156,N_11513,N_10854);
or U14157 (N_14157,N_9765,N_11733);
or U14158 (N_14158,N_10465,N_10973);
nor U14159 (N_14159,N_9761,N_10653);
nand U14160 (N_14160,N_11813,N_11114);
and U14161 (N_14161,N_11924,N_11250);
and U14162 (N_14162,N_9747,N_11445);
nand U14163 (N_14163,N_11539,N_11366);
and U14164 (N_14164,N_9293,N_9884);
nand U14165 (N_14165,N_9061,N_10344);
or U14166 (N_14166,N_11673,N_9827);
nand U14167 (N_14167,N_10604,N_11978);
or U14168 (N_14168,N_10395,N_10177);
or U14169 (N_14169,N_10908,N_11916);
or U14170 (N_14170,N_9869,N_10377);
or U14171 (N_14171,N_11572,N_9501);
and U14172 (N_14172,N_10584,N_10015);
and U14173 (N_14173,N_11009,N_11114);
or U14174 (N_14174,N_11832,N_10723);
or U14175 (N_14175,N_10250,N_9106);
nor U14176 (N_14176,N_10986,N_11761);
and U14177 (N_14177,N_9531,N_9672);
nand U14178 (N_14178,N_11325,N_10453);
nand U14179 (N_14179,N_9192,N_10050);
and U14180 (N_14180,N_11662,N_10805);
nand U14181 (N_14181,N_9254,N_9548);
nand U14182 (N_14182,N_11372,N_9021);
nor U14183 (N_14183,N_10312,N_10523);
nor U14184 (N_14184,N_10328,N_9910);
and U14185 (N_14185,N_10717,N_11969);
xor U14186 (N_14186,N_11670,N_11130);
and U14187 (N_14187,N_11523,N_9070);
and U14188 (N_14188,N_11012,N_9950);
nand U14189 (N_14189,N_9527,N_11554);
xnor U14190 (N_14190,N_9275,N_9679);
xor U14191 (N_14191,N_11942,N_10918);
xnor U14192 (N_14192,N_11784,N_9397);
or U14193 (N_14193,N_10692,N_10061);
nand U14194 (N_14194,N_11530,N_9682);
and U14195 (N_14195,N_9590,N_10025);
nor U14196 (N_14196,N_9690,N_10572);
and U14197 (N_14197,N_10328,N_9291);
or U14198 (N_14198,N_10852,N_11599);
nor U14199 (N_14199,N_9045,N_11994);
xnor U14200 (N_14200,N_10761,N_11227);
nor U14201 (N_14201,N_11557,N_11873);
or U14202 (N_14202,N_10364,N_10432);
nand U14203 (N_14203,N_10650,N_9984);
and U14204 (N_14204,N_10313,N_10061);
and U14205 (N_14205,N_9657,N_10082);
or U14206 (N_14206,N_10843,N_10617);
nand U14207 (N_14207,N_9219,N_9198);
or U14208 (N_14208,N_9892,N_9330);
or U14209 (N_14209,N_11013,N_11748);
xor U14210 (N_14210,N_11444,N_10618);
or U14211 (N_14211,N_10187,N_9559);
nand U14212 (N_14212,N_9337,N_10055);
and U14213 (N_14213,N_10272,N_10078);
nand U14214 (N_14214,N_10411,N_11908);
nor U14215 (N_14215,N_10137,N_11910);
and U14216 (N_14216,N_11571,N_9235);
nand U14217 (N_14217,N_11164,N_11306);
nand U14218 (N_14218,N_9561,N_11309);
or U14219 (N_14219,N_11287,N_9299);
nand U14220 (N_14220,N_9673,N_10868);
xnor U14221 (N_14221,N_10953,N_9247);
nor U14222 (N_14222,N_9605,N_9570);
or U14223 (N_14223,N_11144,N_11205);
or U14224 (N_14224,N_10441,N_11681);
nand U14225 (N_14225,N_11727,N_10550);
nor U14226 (N_14226,N_10460,N_9330);
nand U14227 (N_14227,N_9585,N_9127);
or U14228 (N_14228,N_10831,N_11834);
nand U14229 (N_14229,N_10203,N_10947);
and U14230 (N_14230,N_11610,N_10065);
nor U14231 (N_14231,N_11669,N_9246);
and U14232 (N_14232,N_9788,N_9442);
nor U14233 (N_14233,N_11764,N_10833);
nand U14234 (N_14234,N_11568,N_10475);
and U14235 (N_14235,N_10384,N_11964);
or U14236 (N_14236,N_10889,N_11811);
or U14237 (N_14237,N_9636,N_11706);
or U14238 (N_14238,N_9158,N_10200);
or U14239 (N_14239,N_10956,N_9537);
and U14240 (N_14240,N_10054,N_9773);
nor U14241 (N_14241,N_11585,N_11698);
nor U14242 (N_14242,N_9554,N_9309);
or U14243 (N_14243,N_11607,N_11692);
or U14244 (N_14244,N_11197,N_9731);
and U14245 (N_14245,N_11729,N_10005);
nand U14246 (N_14246,N_10250,N_9634);
nor U14247 (N_14247,N_11848,N_11397);
nand U14248 (N_14248,N_10744,N_11840);
xor U14249 (N_14249,N_11897,N_11351);
xnor U14250 (N_14250,N_11014,N_10576);
nor U14251 (N_14251,N_10117,N_11781);
and U14252 (N_14252,N_11159,N_10019);
nor U14253 (N_14253,N_10728,N_9805);
xor U14254 (N_14254,N_10080,N_10937);
nand U14255 (N_14255,N_9083,N_11767);
nand U14256 (N_14256,N_9645,N_10086);
and U14257 (N_14257,N_9789,N_10136);
nand U14258 (N_14258,N_11351,N_11694);
nand U14259 (N_14259,N_9791,N_9434);
nor U14260 (N_14260,N_10113,N_10755);
nor U14261 (N_14261,N_9995,N_9142);
and U14262 (N_14262,N_9137,N_10678);
nor U14263 (N_14263,N_10160,N_11793);
nor U14264 (N_14264,N_9948,N_9957);
and U14265 (N_14265,N_11003,N_9884);
or U14266 (N_14266,N_11332,N_10500);
or U14267 (N_14267,N_11858,N_10796);
or U14268 (N_14268,N_10830,N_10018);
or U14269 (N_14269,N_10245,N_10428);
nor U14270 (N_14270,N_9168,N_9734);
or U14271 (N_14271,N_10351,N_10807);
and U14272 (N_14272,N_9839,N_10100);
xnor U14273 (N_14273,N_11177,N_10638);
or U14274 (N_14274,N_9858,N_9060);
nor U14275 (N_14275,N_10975,N_9574);
nand U14276 (N_14276,N_11594,N_10542);
nor U14277 (N_14277,N_11451,N_11415);
xnor U14278 (N_14278,N_9014,N_9605);
or U14279 (N_14279,N_11446,N_11233);
xnor U14280 (N_14280,N_10018,N_9182);
or U14281 (N_14281,N_10640,N_11073);
and U14282 (N_14282,N_11347,N_9052);
nand U14283 (N_14283,N_11543,N_10293);
and U14284 (N_14284,N_11844,N_10807);
or U14285 (N_14285,N_11255,N_9900);
xor U14286 (N_14286,N_9356,N_9708);
and U14287 (N_14287,N_11836,N_11426);
or U14288 (N_14288,N_10184,N_9275);
nand U14289 (N_14289,N_11967,N_11528);
nor U14290 (N_14290,N_9109,N_11177);
nand U14291 (N_14291,N_10398,N_11242);
xnor U14292 (N_14292,N_9546,N_9058);
or U14293 (N_14293,N_11390,N_9153);
and U14294 (N_14294,N_11223,N_11637);
nor U14295 (N_14295,N_9814,N_9884);
and U14296 (N_14296,N_9880,N_10177);
and U14297 (N_14297,N_11681,N_10395);
nor U14298 (N_14298,N_10864,N_11377);
nand U14299 (N_14299,N_11210,N_9060);
nand U14300 (N_14300,N_11892,N_11267);
or U14301 (N_14301,N_11026,N_10073);
nor U14302 (N_14302,N_9061,N_11622);
and U14303 (N_14303,N_10106,N_10860);
nand U14304 (N_14304,N_11000,N_10661);
nor U14305 (N_14305,N_9119,N_9606);
and U14306 (N_14306,N_11470,N_11647);
and U14307 (N_14307,N_10222,N_11853);
or U14308 (N_14308,N_10457,N_11867);
nand U14309 (N_14309,N_9247,N_10950);
nand U14310 (N_14310,N_11917,N_9948);
nand U14311 (N_14311,N_11928,N_11445);
or U14312 (N_14312,N_9164,N_9557);
xnor U14313 (N_14313,N_11421,N_9732);
nand U14314 (N_14314,N_11574,N_10646);
nand U14315 (N_14315,N_10318,N_10273);
nor U14316 (N_14316,N_10328,N_11381);
nand U14317 (N_14317,N_11139,N_11757);
or U14318 (N_14318,N_11878,N_11669);
nor U14319 (N_14319,N_9550,N_10896);
nand U14320 (N_14320,N_10279,N_10967);
nor U14321 (N_14321,N_9109,N_11776);
or U14322 (N_14322,N_11485,N_10906);
or U14323 (N_14323,N_9102,N_10210);
nand U14324 (N_14324,N_9369,N_11243);
xnor U14325 (N_14325,N_10414,N_10078);
or U14326 (N_14326,N_11094,N_10104);
nand U14327 (N_14327,N_9080,N_9991);
nor U14328 (N_14328,N_10243,N_10548);
and U14329 (N_14329,N_11639,N_9422);
or U14330 (N_14330,N_11891,N_9043);
nand U14331 (N_14331,N_10692,N_10330);
nand U14332 (N_14332,N_11488,N_10588);
and U14333 (N_14333,N_10955,N_9681);
nor U14334 (N_14334,N_10616,N_10106);
and U14335 (N_14335,N_11215,N_10950);
nand U14336 (N_14336,N_10308,N_10024);
nand U14337 (N_14337,N_11936,N_10500);
nor U14338 (N_14338,N_10507,N_11963);
nand U14339 (N_14339,N_10919,N_9073);
and U14340 (N_14340,N_11559,N_10488);
xor U14341 (N_14341,N_9331,N_11827);
and U14342 (N_14342,N_11498,N_9528);
xor U14343 (N_14343,N_9593,N_9845);
or U14344 (N_14344,N_10028,N_9371);
or U14345 (N_14345,N_11317,N_10652);
and U14346 (N_14346,N_11058,N_9188);
nand U14347 (N_14347,N_10575,N_10075);
xor U14348 (N_14348,N_9106,N_9623);
nor U14349 (N_14349,N_11733,N_10153);
or U14350 (N_14350,N_11408,N_11122);
or U14351 (N_14351,N_9326,N_9652);
xnor U14352 (N_14352,N_10353,N_10783);
nor U14353 (N_14353,N_11075,N_11498);
or U14354 (N_14354,N_9748,N_9197);
and U14355 (N_14355,N_9905,N_10706);
nor U14356 (N_14356,N_10433,N_9779);
nand U14357 (N_14357,N_10399,N_10224);
nor U14358 (N_14358,N_9686,N_9718);
nor U14359 (N_14359,N_9217,N_9804);
or U14360 (N_14360,N_11730,N_10428);
nor U14361 (N_14361,N_10677,N_9518);
xnor U14362 (N_14362,N_9292,N_10564);
nor U14363 (N_14363,N_10411,N_11428);
and U14364 (N_14364,N_10704,N_11444);
nand U14365 (N_14365,N_10910,N_11209);
nand U14366 (N_14366,N_10752,N_10060);
nand U14367 (N_14367,N_10710,N_11352);
nand U14368 (N_14368,N_10879,N_11069);
nand U14369 (N_14369,N_11690,N_10685);
or U14370 (N_14370,N_11608,N_11791);
or U14371 (N_14371,N_10805,N_11360);
xor U14372 (N_14372,N_11772,N_11572);
xor U14373 (N_14373,N_10852,N_11774);
xnor U14374 (N_14374,N_10951,N_9448);
or U14375 (N_14375,N_10376,N_9655);
nor U14376 (N_14376,N_11689,N_9438);
nand U14377 (N_14377,N_11172,N_11254);
and U14378 (N_14378,N_10379,N_9539);
nor U14379 (N_14379,N_11951,N_11080);
nor U14380 (N_14380,N_11615,N_11695);
and U14381 (N_14381,N_10317,N_9212);
or U14382 (N_14382,N_11221,N_11485);
nand U14383 (N_14383,N_10247,N_11006);
nand U14384 (N_14384,N_11891,N_10677);
nand U14385 (N_14385,N_11221,N_9790);
nand U14386 (N_14386,N_9182,N_9022);
and U14387 (N_14387,N_10569,N_11113);
nand U14388 (N_14388,N_10684,N_9887);
nand U14389 (N_14389,N_9918,N_11333);
nor U14390 (N_14390,N_11102,N_10557);
or U14391 (N_14391,N_11924,N_10189);
or U14392 (N_14392,N_11690,N_11145);
and U14393 (N_14393,N_10643,N_11569);
nand U14394 (N_14394,N_9612,N_11440);
nor U14395 (N_14395,N_9169,N_10861);
or U14396 (N_14396,N_9283,N_9161);
nand U14397 (N_14397,N_10227,N_9544);
nand U14398 (N_14398,N_9464,N_10813);
xnor U14399 (N_14399,N_9560,N_9867);
xnor U14400 (N_14400,N_9765,N_11521);
or U14401 (N_14401,N_11681,N_9126);
or U14402 (N_14402,N_10225,N_11664);
nand U14403 (N_14403,N_10646,N_11197);
or U14404 (N_14404,N_10090,N_9459);
and U14405 (N_14405,N_11886,N_9391);
or U14406 (N_14406,N_10385,N_10758);
nand U14407 (N_14407,N_11583,N_10921);
nor U14408 (N_14408,N_9803,N_10122);
nor U14409 (N_14409,N_10120,N_11088);
and U14410 (N_14410,N_10904,N_9936);
nand U14411 (N_14411,N_10436,N_11394);
and U14412 (N_14412,N_9949,N_10888);
or U14413 (N_14413,N_9274,N_9809);
or U14414 (N_14414,N_10373,N_10429);
nor U14415 (N_14415,N_11569,N_9938);
xnor U14416 (N_14416,N_9082,N_11197);
nand U14417 (N_14417,N_11489,N_9683);
or U14418 (N_14418,N_9614,N_10276);
nor U14419 (N_14419,N_10252,N_9855);
xor U14420 (N_14420,N_11421,N_10493);
nand U14421 (N_14421,N_9392,N_10796);
or U14422 (N_14422,N_9367,N_9315);
and U14423 (N_14423,N_9839,N_9188);
xnor U14424 (N_14424,N_9507,N_9332);
nand U14425 (N_14425,N_9005,N_10021);
or U14426 (N_14426,N_11950,N_10642);
or U14427 (N_14427,N_9766,N_10364);
and U14428 (N_14428,N_11087,N_9129);
nor U14429 (N_14429,N_9754,N_10946);
and U14430 (N_14430,N_11292,N_9295);
nand U14431 (N_14431,N_10287,N_9598);
nand U14432 (N_14432,N_11612,N_9718);
xnor U14433 (N_14433,N_10884,N_9207);
xor U14434 (N_14434,N_11833,N_11202);
xnor U14435 (N_14435,N_10606,N_9208);
and U14436 (N_14436,N_10570,N_10928);
nor U14437 (N_14437,N_10788,N_11952);
or U14438 (N_14438,N_11405,N_10313);
nand U14439 (N_14439,N_9516,N_11221);
nand U14440 (N_14440,N_9325,N_9348);
and U14441 (N_14441,N_9348,N_10179);
xor U14442 (N_14442,N_11156,N_9352);
xnor U14443 (N_14443,N_9381,N_10848);
nor U14444 (N_14444,N_9809,N_11774);
nor U14445 (N_14445,N_9641,N_9999);
nor U14446 (N_14446,N_10720,N_11357);
and U14447 (N_14447,N_9296,N_10969);
or U14448 (N_14448,N_9074,N_11412);
nor U14449 (N_14449,N_11189,N_10718);
nor U14450 (N_14450,N_11843,N_9808);
or U14451 (N_14451,N_9065,N_9337);
or U14452 (N_14452,N_10517,N_10468);
or U14453 (N_14453,N_11357,N_10634);
or U14454 (N_14454,N_9037,N_10390);
xnor U14455 (N_14455,N_9628,N_9061);
nand U14456 (N_14456,N_9021,N_9214);
nor U14457 (N_14457,N_11236,N_10631);
nand U14458 (N_14458,N_9361,N_10995);
or U14459 (N_14459,N_10191,N_11230);
nor U14460 (N_14460,N_11310,N_9709);
or U14461 (N_14461,N_11467,N_10683);
nor U14462 (N_14462,N_9239,N_11856);
and U14463 (N_14463,N_10397,N_11194);
nor U14464 (N_14464,N_11805,N_10039);
nor U14465 (N_14465,N_11297,N_9906);
nand U14466 (N_14466,N_10240,N_11444);
nand U14467 (N_14467,N_11881,N_10527);
and U14468 (N_14468,N_10164,N_9200);
nor U14469 (N_14469,N_9330,N_10823);
or U14470 (N_14470,N_11478,N_9521);
nor U14471 (N_14471,N_11713,N_10287);
nand U14472 (N_14472,N_11031,N_11093);
nor U14473 (N_14473,N_10882,N_9428);
nand U14474 (N_14474,N_11205,N_9736);
nor U14475 (N_14475,N_11553,N_9494);
and U14476 (N_14476,N_11015,N_9648);
nand U14477 (N_14477,N_9148,N_11442);
nor U14478 (N_14478,N_10792,N_9592);
nand U14479 (N_14479,N_11766,N_11396);
and U14480 (N_14480,N_11393,N_10557);
nor U14481 (N_14481,N_9696,N_11630);
and U14482 (N_14482,N_9937,N_9683);
and U14483 (N_14483,N_9148,N_9200);
nor U14484 (N_14484,N_10246,N_9081);
xnor U14485 (N_14485,N_9217,N_9167);
and U14486 (N_14486,N_9894,N_9801);
nand U14487 (N_14487,N_10356,N_10518);
and U14488 (N_14488,N_11456,N_11491);
or U14489 (N_14489,N_11027,N_10102);
nand U14490 (N_14490,N_9920,N_11627);
nor U14491 (N_14491,N_11922,N_11700);
nand U14492 (N_14492,N_11061,N_11287);
nand U14493 (N_14493,N_9073,N_9646);
or U14494 (N_14494,N_10849,N_9475);
nand U14495 (N_14495,N_11471,N_11166);
nor U14496 (N_14496,N_11100,N_9972);
xnor U14497 (N_14497,N_11188,N_10166);
xnor U14498 (N_14498,N_10960,N_10565);
or U14499 (N_14499,N_11742,N_9381);
nor U14500 (N_14500,N_10358,N_10979);
nand U14501 (N_14501,N_9129,N_9662);
or U14502 (N_14502,N_9449,N_11182);
nor U14503 (N_14503,N_11115,N_10400);
or U14504 (N_14504,N_9974,N_10180);
nand U14505 (N_14505,N_10341,N_11757);
and U14506 (N_14506,N_10710,N_10396);
or U14507 (N_14507,N_9201,N_10365);
nand U14508 (N_14508,N_9670,N_9540);
and U14509 (N_14509,N_11051,N_9424);
xnor U14510 (N_14510,N_9953,N_10874);
xor U14511 (N_14511,N_9721,N_9780);
xor U14512 (N_14512,N_10149,N_10107);
and U14513 (N_14513,N_9982,N_10436);
nand U14514 (N_14514,N_11063,N_11970);
nand U14515 (N_14515,N_10584,N_9241);
nor U14516 (N_14516,N_9523,N_10330);
nand U14517 (N_14517,N_9626,N_10227);
and U14518 (N_14518,N_11584,N_9839);
nor U14519 (N_14519,N_10715,N_9446);
or U14520 (N_14520,N_11481,N_11862);
xnor U14521 (N_14521,N_11080,N_10512);
and U14522 (N_14522,N_11597,N_11424);
or U14523 (N_14523,N_10302,N_11628);
xnor U14524 (N_14524,N_11634,N_11483);
nand U14525 (N_14525,N_9443,N_9637);
xnor U14526 (N_14526,N_10492,N_11218);
and U14527 (N_14527,N_9649,N_10549);
or U14528 (N_14528,N_10050,N_11907);
nand U14529 (N_14529,N_9774,N_9701);
nand U14530 (N_14530,N_11309,N_10462);
nor U14531 (N_14531,N_10641,N_11572);
nor U14532 (N_14532,N_9204,N_11004);
or U14533 (N_14533,N_10313,N_11838);
and U14534 (N_14534,N_11828,N_9828);
nor U14535 (N_14535,N_9103,N_11787);
nor U14536 (N_14536,N_9222,N_10545);
nand U14537 (N_14537,N_9618,N_11190);
xnor U14538 (N_14538,N_11917,N_10675);
xor U14539 (N_14539,N_11129,N_9152);
or U14540 (N_14540,N_10300,N_9244);
nor U14541 (N_14541,N_10699,N_9465);
or U14542 (N_14542,N_11002,N_10300);
and U14543 (N_14543,N_10850,N_10257);
nand U14544 (N_14544,N_10772,N_9435);
nor U14545 (N_14545,N_10865,N_9581);
nand U14546 (N_14546,N_11844,N_11813);
or U14547 (N_14547,N_10058,N_10025);
xnor U14548 (N_14548,N_9399,N_10474);
and U14549 (N_14549,N_10414,N_11580);
or U14550 (N_14550,N_11907,N_10852);
nand U14551 (N_14551,N_11386,N_10575);
or U14552 (N_14552,N_9716,N_9203);
and U14553 (N_14553,N_11243,N_9943);
nor U14554 (N_14554,N_9511,N_11309);
xor U14555 (N_14555,N_10965,N_10873);
and U14556 (N_14556,N_11660,N_11493);
nand U14557 (N_14557,N_11247,N_10060);
nor U14558 (N_14558,N_9633,N_10499);
nor U14559 (N_14559,N_9608,N_10611);
and U14560 (N_14560,N_11904,N_10694);
nand U14561 (N_14561,N_9154,N_9909);
nand U14562 (N_14562,N_9838,N_9606);
and U14563 (N_14563,N_11677,N_10533);
nand U14564 (N_14564,N_9796,N_11982);
nand U14565 (N_14565,N_11834,N_9028);
nand U14566 (N_14566,N_9323,N_9495);
nor U14567 (N_14567,N_11581,N_11428);
nand U14568 (N_14568,N_10705,N_10809);
nand U14569 (N_14569,N_9221,N_11064);
nand U14570 (N_14570,N_10227,N_10861);
and U14571 (N_14571,N_9181,N_9211);
and U14572 (N_14572,N_10431,N_9717);
or U14573 (N_14573,N_9359,N_10151);
nand U14574 (N_14574,N_11227,N_9836);
and U14575 (N_14575,N_11023,N_10559);
or U14576 (N_14576,N_11357,N_9126);
and U14577 (N_14577,N_9924,N_10067);
nor U14578 (N_14578,N_10519,N_9762);
or U14579 (N_14579,N_9516,N_11257);
or U14580 (N_14580,N_9508,N_11675);
xor U14581 (N_14581,N_9740,N_10196);
nand U14582 (N_14582,N_9732,N_9779);
or U14583 (N_14583,N_11444,N_10289);
nand U14584 (N_14584,N_10448,N_9675);
xnor U14585 (N_14585,N_9991,N_11392);
nand U14586 (N_14586,N_11604,N_10116);
or U14587 (N_14587,N_11900,N_9844);
and U14588 (N_14588,N_9090,N_11130);
nor U14589 (N_14589,N_9953,N_11843);
nor U14590 (N_14590,N_11557,N_9016);
and U14591 (N_14591,N_9347,N_11235);
or U14592 (N_14592,N_10555,N_9240);
and U14593 (N_14593,N_10094,N_9832);
and U14594 (N_14594,N_11852,N_11221);
or U14595 (N_14595,N_10775,N_10509);
nor U14596 (N_14596,N_9390,N_10548);
nand U14597 (N_14597,N_11855,N_10228);
and U14598 (N_14598,N_10206,N_11807);
and U14599 (N_14599,N_11013,N_10257);
or U14600 (N_14600,N_9297,N_9839);
and U14601 (N_14601,N_9129,N_11105);
or U14602 (N_14602,N_11014,N_11127);
nor U14603 (N_14603,N_11834,N_11484);
nor U14604 (N_14604,N_9107,N_10208);
nand U14605 (N_14605,N_9367,N_9203);
and U14606 (N_14606,N_9873,N_11786);
nand U14607 (N_14607,N_11322,N_11301);
nor U14608 (N_14608,N_11139,N_11912);
or U14609 (N_14609,N_9444,N_10074);
or U14610 (N_14610,N_10944,N_11866);
xnor U14611 (N_14611,N_9157,N_10671);
and U14612 (N_14612,N_11583,N_9286);
or U14613 (N_14613,N_11330,N_9168);
or U14614 (N_14614,N_11188,N_11472);
nor U14615 (N_14615,N_10273,N_11021);
nand U14616 (N_14616,N_11799,N_9485);
or U14617 (N_14617,N_9771,N_11012);
or U14618 (N_14618,N_9303,N_11741);
or U14619 (N_14619,N_11829,N_10228);
or U14620 (N_14620,N_11070,N_9785);
nand U14621 (N_14621,N_9875,N_10945);
nor U14622 (N_14622,N_10011,N_9315);
xor U14623 (N_14623,N_9762,N_9434);
or U14624 (N_14624,N_11916,N_9300);
nor U14625 (N_14625,N_11967,N_9251);
and U14626 (N_14626,N_9404,N_11952);
and U14627 (N_14627,N_11187,N_10282);
or U14628 (N_14628,N_9087,N_10350);
or U14629 (N_14629,N_9434,N_10651);
nor U14630 (N_14630,N_11340,N_9995);
nand U14631 (N_14631,N_11299,N_11579);
or U14632 (N_14632,N_9516,N_11737);
and U14633 (N_14633,N_11567,N_10988);
nor U14634 (N_14634,N_11710,N_10060);
nand U14635 (N_14635,N_10703,N_10828);
and U14636 (N_14636,N_9997,N_11415);
nor U14637 (N_14637,N_11951,N_9575);
and U14638 (N_14638,N_9381,N_9066);
nand U14639 (N_14639,N_10214,N_10766);
or U14640 (N_14640,N_9098,N_9676);
nor U14641 (N_14641,N_9320,N_10223);
xnor U14642 (N_14642,N_9364,N_10353);
nand U14643 (N_14643,N_11908,N_9910);
nor U14644 (N_14644,N_10093,N_9628);
nor U14645 (N_14645,N_11604,N_10447);
and U14646 (N_14646,N_10789,N_11115);
and U14647 (N_14647,N_9700,N_10802);
or U14648 (N_14648,N_9379,N_10585);
and U14649 (N_14649,N_11399,N_11544);
and U14650 (N_14650,N_10941,N_10218);
xor U14651 (N_14651,N_9540,N_11672);
nor U14652 (N_14652,N_10408,N_10178);
nor U14653 (N_14653,N_10903,N_9296);
xor U14654 (N_14654,N_10079,N_11187);
or U14655 (N_14655,N_9381,N_9629);
xor U14656 (N_14656,N_10896,N_9647);
and U14657 (N_14657,N_9481,N_9394);
and U14658 (N_14658,N_11400,N_11186);
nand U14659 (N_14659,N_9692,N_11033);
and U14660 (N_14660,N_11071,N_10301);
nand U14661 (N_14661,N_10336,N_11702);
and U14662 (N_14662,N_10372,N_10199);
and U14663 (N_14663,N_9322,N_10725);
or U14664 (N_14664,N_10159,N_11218);
nor U14665 (N_14665,N_11890,N_10359);
nand U14666 (N_14666,N_11616,N_11191);
xnor U14667 (N_14667,N_10860,N_11156);
or U14668 (N_14668,N_9754,N_11593);
nor U14669 (N_14669,N_9995,N_11097);
or U14670 (N_14670,N_10648,N_9621);
or U14671 (N_14671,N_10206,N_11406);
or U14672 (N_14672,N_11444,N_11411);
or U14673 (N_14673,N_10180,N_9085);
xnor U14674 (N_14674,N_11253,N_9967);
and U14675 (N_14675,N_9165,N_9009);
nor U14676 (N_14676,N_11671,N_11508);
nand U14677 (N_14677,N_9621,N_9810);
nor U14678 (N_14678,N_11408,N_9336);
or U14679 (N_14679,N_10578,N_11086);
and U14680 (N_14680,N_9076,N_10260);
xnor U14681 (N_14681,N_11377,N_9200);
nor U14682 (N_14682,N_10786,N_11686);
nor U14683 (N_14683,N_10523,N_11878);
or U14684 (N_14684,N_9237,N_9880);
or U14685 (N_14685,N_10496,N_10857);
and U14686 (N_14686,N_10385,N_10339);
or U14687 (N_14687,N_10165,N_11731);
xor U14688 (N_14688,N_10853,N_9134);
or U14689 (N_14689,N_9373,N_9000);
or U14690 (N_14690,N_10747,N_10669);
nor U14691 (N_14691,N_11816,N_10023);
nand U14692 (N_14692,N_11441,N_11098);
and U14693 (N_14693,N_11188,N_11647);
nor U14694 (N_14694,N_10597,N_9441);
nand U14695 (N_14695,N_10417,N_10491);
or U14696 (N_14696,N_10574,N_9533);
or U14697 (N_14697,N_11130,N_11205);
or U14698 (N_14698,N_11347,N_10468);
and U14699 (N_14699,N_11784,N_11809);
nand U14700 (N_14700,N_9033,N_9554);
xor U14701 (N_14701,N_11425,N_9396);
xor U14702 (N_14702,N_10640,N_9628);
and U14703 (N_14703,N_9962,N_9294);
nand U14704 (N_14704,N_10947,N_10409);
nor U14705 (N_14705,N_11519,N_9685);
and U14706 (N_14706,N_10089,N_11379);
and U14707 (N_14707,N_11585,N_10681);
and U14708 (N_14708,N_10769,N_11079);
or U14709 (N_14709,N_10297,N_10349);
nor U14710 (N_14710,N_11260,N_9191);
nor U14711 (N_14711,N_10676,N_9265);
nand U14712 (N_14712,N_9337,N_11907);
and U14713 (N_14713,N_9136,N_10963);
or U14714 (N_14714,N_11495,N_11665);
or U14715 (N_14715,N_10390,N_10526);
nand U14716 (N_14716,N_10147,N_10132);
nand U14717 (N_14717,N_10574,N_11940);
and U14718 (N_14718,N_11442,N_11736);
and U14719 (N_14719,N_9036,N_9220);
and U14720 (N_14720,N_10090,N_9134);
nor U14721 (N_14721,N_11290,N_10780);
nand U14722 (N_14722,N_10462,N_9184);
xnor U14723 (N_14723,N_10629,N_11498);
and U14724 (N_14724,N_11077,N_11031);
and U14725 (N_14725,N_9738,N_10337);
nand U14726 (N_14726,N_10305,N_9554);
or U14727 (N_14727,N_11359,N_11290);
and U14728 (N_14728,N_9551,N_11934);
nand U14729 (N_14729,N_9539,N_10529);
nand U14730 (N_14730,N_10514,N_9110);
or U14731 (N_14731,N_9033,N_11442);
nand U14732 (N_14732,N_9732,N_9229);
or U14733 (N_14733,N_9153,N_9022);
nor U14734 (N_14734,N_10400,N_10675);
or U14735 (N_14735,N_11941,N_11810);
and U14736 (N_14736,N_11624,N_10385);
or U14737 (N_14737,N_11758,N_9742);
or U14738 (N_14738,N_9450,N_11383);
nand U14739 (N_14739,N_10588,N_10070);
or U14740 (N_14740,N_9322,N_10404);
nor U14741 (N_14741,N_10697,N_11083);
nor U14742 (N_14742,N_9448,N_10286);
or U14743 (N_14743,N_9279,N_11814);
or U14744 (N_14744,N_10564,N_10645);
xor U14745 (N_14745,N_10541,N_10724);
or U14746 (N_14746,N_10436,N_11593);
nor U14747 (N_14747,N_11479,N_9247);
or U14748 (N_14748,N_9983,N_10784);
or U14749 (N_14749,N_10468,N_9467);
nor U14750 (N_14750,N_10481,N_9712);
or U14751 (N_14751,N_9168,N_11141);
xnor U14752 (N_14752,N_9767,N_10594);
nand U14753 (N_14753,N_10801,N_10855);
nor U14754 (N_14754,N_11064,N_11087);
or U14755 (N_14755,N_10365,N_10829);
or U14756 (N_14756,N_10919,N_9914);
and U14757 (N_14757,N_9957,N_11716);
or U14758 (N_14758,N_9630,N_9021);
or U14759 (N_14759,N_9919,N_10547);
and U14760 (N_14760,N_11833,N_9569);
or U14761 (N_14761,N_11936,N_10488);
and U14762 (N_14762,N_11150,N_10226);
nor U14763 (N_14763,N_11186,N_11440);
nand U14764 (N_14764,N_9088,N_11590);
nand U14765 (N_14765,N_11929,N_10618);
nand U14766 (N_14766,N_10991,N_10755);
or U14767 (N_14767,N_11516,N_9418);
or U14768 (N_14768,N_9612,N_9510);
nor U14769 (N_14769,N_11543,N_9883);
nor U14770 (N_14770,N_9461,N_11340);
and U14771 (N_14771,N_11534,N_10499);
xor U14772 (N_14772,N_9117,N_10971);
and U14773 (N_14773,N_9087,N_10961);
and U14774 (N_14774,N_11268,N_10940);
xor U14775 (N_14775,N_11535,N_10475);
nor U14776 (N_14776,N_9848,N_10177);
nor U14777 (N_14777,N_10706,N_11745);
or U14778 (N_14778,N_10211,N_11852);
nand U14779 (N_14779,N_10842,N_11670);
and U14780 (N_14780,N_9810,N_10469);
nand U14781 (N_14781,N_11851,N_10142);
nor U14782 (N_14782,N_11321,N_9091);
nand U14783 (N_14783,N_10542,N_10495);
or U14784 (N_14784,N_10468,N_9624);
nand U14785 (N_14785,N_9445,N_9115);
nand U14786 (N_14786,N_9152,N_11503);
nand U14787 (N_14787,N_10295,N_10488);
nand U14788 (N_14788,N_9918,N_9384);
and U14789 (N_14789,N_11302,N_10430);
nor U14790 (N_14790,N_9843,N_10066);
nand U14791 (N_14791,N_10771,N_10973);
nand U14792 (N_14792,N_9693,N_11164);
xor U14793 (N_14793,N_9553,N_9794);
and U14794 (N_14794,N_10523,N_11085);
nor U14795 (N_14795,N_11109,N_10579);
nand U14796 (N_14796,N_9080,N_9961);
nor U14797 (N_14797,N_11743,N_10903);
or U14798 (N_14798,N_9611,N_11391);
nand U14799 (N_14799,N_9121,N_11465);
or U14800 (N_14800,N_9508,N_10638);
and U14801 (N_14801,N_9855,N_11181);
nor U14802 (N_14802,N_11598,N_11271);
or U14803 (N_14803,N_11876,N_9870);
nand U14804 (N_14804,N_11764,N_11730);
nand U14805 (N_14805,N_11337,N_10355);
and U14806 (N_14806,N_9063,N_9967);
nand U14807 (N_14807,N_11229,N_9012);
or U14808 (N_14808,N_10203,N_9715);
xor U14809 (N_14809,N_10897,N_10510);
and U14810 (N_14810,N_11701,N_11966);
nor U14811 (N_14811,N_9122,N_11616);
nor U14812 (N_14812,N_11497,N_9971);
nor U14813 (N_14813,N_11053,N_11938);
nand U14814 (N_14814,N_9382,N_9301);
nand U14815 (N_14815,N_11791,N_9602);
and U14816 (N_14816,N_9486,N_9093);
and U14817 (N_14817,N_9491,N_9299);
and U14818 (N_14818,N_9769,N_11200);
and U14819 (N_14819,N_11086,N_9259);
nand U14820 (N_14820,N_10628,N_9033);
nand U14821 (N_14821,N_9055,N_9453);
and U14822 (N_14822,N_9177,N_11973);
and U14823 (N_14823,N_9617,N_11634);
and U14824 (N_14824,N_11564,N_10350);
nor U14825 (N_14825,N_9726,N_9532);
nor U14826 (N_14826,N_11903,N_10859);
xnor U14827 (N_14827,N_10278,N_9151);
nand U14828 (N_14828,N_11511,N_11926);
nor U14829 (N_14829,N_11705,N_9703);
or U14830 (N_14830,N_11785,N_10881);
or U14831 (N_14831,N_11926,N_11577);
and U14832 (N_14832,N_10116,N_10541);
nor U14833 (N_14833,N_10292,N_11829);
or U14834 (N_14834,N_9945,N_10963);
xnor U14835 (N_14835,N_10683,N_11430);
nand U14836 (N_14836,N_10770,N_10551);
nand U14837 (N_14837,N_11348,N_11794);
nor U14838 (N_14838,N_9128,N_9329);
and U14839 (N_14839,N_9616,N_11656);
nor U14840 (N_14840,N_11043,N_9017);
or U14841 (N_14841,N_9286,N_9685);
and U14842 (N_14842,N_11787,N_9806);
nor U14843 (N_14843,N_9607,N_9777);
nor U14844 (N_14844,N_10603,N_9542);
nand U14845 (N_14845,N_11708,N_9844);
nor U14846 (N_14846,N_11795,N_9659);
nor U14847 (N_14847,N_10754,N_9930);
or U14848 (N_14848,N_10781,N_10394);
xor U14849 (N_14849,N_10146,N_11425);
and U14850 (N_14850,N_10459,N_9275);
and U14851 (N_14851,N_10277,N_9397);
or U14852 (N_14852,N_11297,N_9444);
and U14853 (N_14853,N_10763,N_9180);
or U14854 (N_14854,N_9641,N_9077);
or U14855 (N_14855,N_9786,N_9537);
nand U14856 (N_14856,N_11702,N_11694);
nor U14857 (N_14857,N_9757,N_11387);
xnor U14858 (N_14858,N_10374,N_11939);
and U14859 (N_14859,N_9618,N_9949);
or U14860 (N_14860,N_11182,N_11639);
nor U14861 (N_14861,N_11342,N_11910);
nor U14862 (N_14862,N_10658,N_9497);
and U14863 (N_14863,N_10889,N_10394);
nand U14864 (N_14864,N_9709,N_10824);
nand U14865 (N_14865,N_10709,N_11661);
nor U14866 (N_14866,N_11088,N_11467);
nand U14867 (N_14867,N_11024,N_11732);
nand U14868 (N_14868,N_9623,N_9782);
nand U14869 (N_14869,N_11245,N_11058);
or U14870 (N_14870,N_9813,N_10948);
xnor U14871 (N_14871,N_11931,N_10115);
or U14872 (N_14872,N_10177,N_9249);
and U14873 (N_14873,N_11707,N_10930);
and U14874 (N_14874,N_11877,N_11600);
or U14875 (N_14875,N_10847,N_10906);
and U14876 (N_14876,N_9711,N_9228);
or U14877 (N_14877,N_10710,N_11300);
nor U14878 (N_14878,N_9708,N_11948);
and U14879 (N_14879,N_10990,N_10570);
nand U14880 (N_14880,N_11857,N_9320);
and U14881 (N_14881,N_9050,N_11949);
nand U14882 (N_14882,N_9220,N_9370);
or U14883 (N_14883,N_9913,N_10741);
and U14884 (N_14884,N_10125,N_10392);
nor U14885 (N_14885,N_9405,N_9464);
or U14886 (N_14886,N_10994,N_10224);
nand U14887 (N_14887,N_9368,N_10941);
or U14888 (N_14888,N_9890,N_10066);
nand U14889 (N_14889,N_10462,N_9133);
nand U14890 (N_14890,N_10541,N_9383);
nor U14891 (N_14891,N_9942,N_9211);
and U14892 (N_14892,N_10598,N_9173);
or U14893 (N_14893,N_9938,N_10051);
nor U14894 (N_14894,N_11026,N_10745);
nor U14895 (N_14895,N_9049,N_10888);
and U14896 (N_14896,N_9766,N_10880);
and U14897 (N_14897,N_9669,N_9478);
or U14898 (N_14898,N_11270,N_9543);
nor U14899 (N_14899,N_11484,N_9197);
nor U14900 (N_14900,N_9008,N_9164);
nor U14901 (N_14901,N_10513,N_10940);
and U14902 (N_14902,N_11419,N_10861);
nor U14903 (N_14903,N_10430,N_10084);
nand U14904 (N_14904,N_9309,N_10816);
and U14905 (N_14905,N_10456,N_11905);
and U14906 (N_14906,N_10829,N_9487);
nand U14907 (N_14907,N_9940,N_11205);
nor U14908 (N_14908,N_11893,N_9692);
xnor U14909 (N_14909,N_9721,N_9475);
and U14910 (N_14910,N_10726,N_9620);
nor U14911 (N_14911,N_9231,N_11585);
and U14912 (N_14912,N_11092,N_11446);
and U14913 (N_14913,N_11233,N_10954);
and U14914 (N_14914,N_9818,N_11965);
or U14915 (N_14915,N_9097,N_10972);
and U14916 (N_14916,N_9295,N_11188);
nand U14917 (N_14917,N_11861,N_10641);
nor U14918 (N_14918,N_9910,N_11608);
and U14919 (N_14919,N_9908,N_11396);
and U14920 (N_14920,N_11489,N_10120);
nor U14921 (N_14921,N_9441,N_11202);
nand U14922 (N_14922,N_9064,N_11208);
xor U14923 (N_14923,N_9633,N_9567);
xnor U14924 (N_14924,N_10521,N_10861);
and U14925 (N_14925,N_9170,N_11190);
nor U14926 (N_14926,N_10809,N_11399);
nor U14927 (N_14927,N_11237,N_9112);
and U14928 (N_14928,N_10708,N_11503);
nand U14929 (N_14929,N_11480,N_10670);
xor U14930 (N_14930,N_9688,N_9768);
nand U14931 (N_14931,N_9428,N_9986);
or U14932 (N_14932,N_11602,N_9839);
or U14933 (N_14933,N_10434,N_10260);
or U14934 (N_14934,N_10206,N_9021);
xnor U14935 (N_14935,N_11790,N_10779);
nand U14936 (N_14936,N_10478,N_9029);
nand U14937 (N_14937,N_10677,N_9239);
or U14938 (N_14938,N_10292,N_11684);
or U14939 (N_14939,N_10372,N_9549);
xnor U14940 (N_14940,N_9567,N_11169);
xor U14941 (N_14941,N_10323,N_9215);
nor U14942 (N_14942,N_9045,N_11552);
nand U14943 (N_14943,N_11937,N_11922);
xor U14944 (N_14944,N_11082,N_11250);
nand U14945 (N_14945,N_9254,N_9154);
nand U14946 (N_14946,N_10466,N_10184);
nor U14947 (N_14947,N_10220,N_10755);
nand U14948 (N_14948,N_9823,N_10506);
or U14949 (N_14949,N_10915,N_9205);
or U14950 (N_14950,N_11468,N_11164);
and U14951 (N_14951,N_10278,N_10280);
or U14952 (N_14952,N_9354,N_10130);
or U14953 (N_14953,N_11048,N_10242);
xor U14954 (N_14954,N_11480,N_11582);
and U14955 (N_14955,N_9198,N_11865);
nand U14956 (N_14956,N_9482,N_10811);
nand U14957 (N_14957,N_11973,N_11376);
or U14958 (N_14958,N_10350,N_9120);
or U14959 (N_14959,N_11008,N_11733);
nand U14960 (N_14960,N_9071,N_9656);
or U14961 (N_14961,N_9270,N_9182);
nand U14962 (N_14962,N_10122,N_9696);
nand U14963 (N_14963,N_10583,N_9505);
or U14964 (N_14964,N_9248,N_11945);
xor U14965 (N_14965,N_9600,N_11452);
xor U14966 (N_14966,N_10529,N_9587);
nand U14967 (N_14967,N_11638,N_11309);
nor U14968 (N_14968,N_10711,N_10461);
and U14969 (N_14969,N_9398,N_11310);
nand U14970 (N_14970,N_10316,N_11308);
or U14971 (N_14971,N_10828,N_11831);
nor U14972 (N_14972,N_9734,N_9154);
nand U14973 (N_14973,N_9192,N_9866);
and U14974 (N_14974,N_11650,N_11854);
nand U14975 (N_14975,N_11602,N_9345);
or U14976 (N_14976,N_10604,N_11886);
nor U14977 (N_14977,N_10681,N_9354);
and U14978 (N_14978,N_11857,N_11101);
and U14979 (N_14979,N_9029,N_11314);
nor U14980 (N_14980,N_9018,N_10507);
and U14981 (N_14981,N_10707,N_10516);
and U14982 (N_14982,N_11224,N_11357);
or U14983 (N_14983,N_10750,N_10167);
nand U14984 (N_14984,N_9788,N_9237);
and U14985 (N_14985,N_11493,N_9162);
or U14986 (N_14986,N_10362,N_10318);
nand U14987 (N_14987,N_11193,N_9573);
nor U14988 (N_14988,N_11149,N_9990);
nor U14989 (N_14989,N_10450,N_10512);
or U14990 (N_14990,N_11445,N_9595);
nor U14991 (N_14991,N_10941,N_9490);
and U14992 (N_14992,N_10972,N_10200);
or U14993 (N_14993,N_9213,N_10807);
and U14994 (N_14994,N_9585,N_9554);
nand U14995 (N_14995,N_9647,N_10207);
nor U14996 (N_14996,N_11666,N_10951);
and U14997 (N_14997,N_9559,N_11627);
nand U14998 (N_14998,N_10515,N_10393);
nor U14999 (N_14999,N_9495,N_10314);
or UO_0 (O_0,N_14560,N_14398);
nand UO_1 (O_1,N_14392,N_12815);
and UO_2 (O_2,N_13783,N_14854);
or UO_3 (O_3,N_13117,N_12560);
xnor UO_4 (O_4,N_12618,N_12296);
or UO_5 (O_5,N_13934,N_13089);
or UO_6 (O_6,N_14628,N_12727);
nor UO_7 (O_7,N_13914,N_13004);
or UO_8 (O_8,N_12260,N_14584);
or UO_9 (O_9,N_14126,N_13388);
nor UO_10 (O_10,N_12381,N_14894);
or UO_11 (O_11,N_13426,N_12382);
nor UO_12 (O_12,N_13471,N_12740);
or UO_13 (O_13,N_13191,N_12191);
or UO_14 (O_14,N_12128,N_12287);
or UO_15 (O_15,N_13266,N_12119);
nand UO_16 (O_16,N_13320,N_14355);
nand UO_17 (O_17,N_13217,N_13535);
xor UO_18 (O_18,N_13122,N_14594);
xnor UO_19 (O_19,N_13165,N_13574);
xnor UO_20 (O_20,N_13243,N_14540);
or UO_21 (O_21,N_14508,N_12485);
nand UO_22 (O_22,N_14779,N_14877);
or UO_23 (O_23,N_13995,N_14983);
and UO_24 (O_24,N_14357,N_13239);
nor UO_25 (O_25,N_14268,N_13469);
and UO_26 (O_26,N_14865,N_12734);
and UO_27 (O_27,N_13031,N_13313);
and UO_28 (O_28,N_13854,N_12476);
nor UO_29 (O_29,N_12845,N_14556);
xnor UO_30 (O_30,N_12344,N_14710);
and UO_31 (O_31,N_12141,N_13837);
and UO_32 (O_32,N_14525,N_13990);
nor UO_33 (O_33,N_13422,N_14656);
nand UO_34 (O_34,N_12208,N_13424);
nor UO_35 (O_35,N_14399,N_13068);
nand UO_36 (O_36,N_13865,N_12171);
nand UO_37 (O_37,N_14408,N_13030);
nand UO_38 (O_38,N_12543,N_14611);
nor UO_39 (O_39,N_14053,N_14499);
and UO_40 (O_40,N_14397,N_14861);
and UO_41 (O_41,N_14231,N_14310);
nand UO_42 (O_42,N_14490,N_12105);
nand UO_43 (O_43,N_14372,N_12003);
nand UO_44 (O_44,N_12684,N_12182);
nand UO_45 (O_45,N_12940,N_14706);
and UO_46 (O_46,N_14244,N_13558);
or UO_47 (O_47,N_14713,N_13070);
nand UO_48 (O_48,N_13417,N_12700);
nand UO_49 (O_49,N_13581,N_13458);
xnor UO_50 (O_50,N_13941,N_13674);
nand UO_51 (O_51,N_13472,N_13959);
nand UO_52 (O_52,N_14339,N_13354);
nand UO_53 (O_53,N_13193,N_13776);
nand UO_54 (O_54,N_12544,N_12489);
and UO_55 (O_55,N_12177,N_13221);
nor UO_56 (O_56,N_13009,N_13702);
xnor UO_57 (O_57,N_13715,N_14204);
and UO_58 (O_58,N_13843,N_13828);
and UO_59 (O_59,N_13307,N_12458);
and UO_60 (O_60,N_12307,N_13363);
nand UO_61 (O_61,N_13541,N_13306);
nand UO_62 (O_62,N_14364,N_12990);
nand UO_63 (O_63,N_13932,N_14287);
xor UO_64 (O_64,N_14825,N_13544);
nor UO_65 (O_65,N_14862,N_12947);
or UO_66 (O_66,N_12033,N_14608);
and UO_67 (O_67,N_14793,N_14463);
and UO_68 (O_68,N_13722,N_12863);
or UO_69 (O_69,N_13698,N_14187);
and UO_70 (O_70,N_12833,N_14311);
nor UO_71 (O_71,N_12397,N_14484);
nand UO_72 (O_72,N_14785,N_12504);
nor UO_73 (O_73,N_13057,N_13000);
nand UO_74 (O_74,N_13749,N_13042);
and UO_75 (O_75,N_14852,N_13358);
nor UO_76 (O_76,N_13149,N_12303);
or UO_77 (O_77,N_12665,N_14654);
nand UO_78 (O_78,N_13938,N_12991);
or UO_79 (O_79,N_14152,N_12830);
and UO_80 (O_80,N_14860,N_13509);
or UO_81 (O_81,N_13287,N_12406);
xnor UO_82 (O_82,N_13220,N_12651);
nor UO_83 (O_83,N_13410,N_13584);
or UO_84 (O_84,N_14191,N_14886);
nand UO_85 (O_85,N_12459,N_14272);
xnor UO_86 (O_86,N_13861,N_14305);
or UO_87 (O_87,N_13918,N_14294);
nand UO_88 (O_88,N_13970,N_12950);
nand UO_89 (O_89,N_13435,N_13814);
xor UO_90 (O_90,N_12978,N_13978);
nor UO_91 (O_91,N_14910,N_12660);
nor UO_92 (O_92,N_12948,N_14087);
nor UO_93 (O_93,N_14390,N_14149);
nor UO_94 (O_94,N_12573,N_14688);
nor UO_95 (O_95,N_13651,N_13807);
or UO_96 (O_96,N_13571,N_14547);
nand UO_97 (O_97,N_14143,N_12689);
or UO_98 (O_98,N_12448,N_14419);
nand UO_99 (O_99,N_12971,N_13910);
or UO_100 (O_100,N_14182,N_13947);
and UO_101 (O_101,N_12244,N_13455);
nor UO_102 (O_102,N_14210,N_13039);
or UO_103 (O_103,N_14802,N_12184);
nand UO_104 (O_104,N_14258,N_12638);
and UO_105 (O_105,N_13025,N_14570);
nand UO_106 (O_106,N_14539,N_13008);
or UO_107 (O_107,N_14964,N_13711);
and UO_108 (O_108,N_13409,N_13290);
or UO_109 (O_109,N_13633,N_13378);
and UO_110 (O_110,N_12807,N_13695);
xor UO_111 (O_111,N_12945,N_14920);
nor UO_112 (O_112,N_14068,N_14958);
nor UO_113 (O_113,N_14801,N_12616);
and UO_114 (O_114,N_14435,N_12685);
or UO_115 (O_115,N_13800,N_13953);
and UO_116 (O_116,N_12509,N_14723);
nand UO_117 (O_117,N_12376,N_14675);
nand UO_118 (O_118,N_13593,N_13218);
and UO_119 (O_119,N_13325,N_12470);
or UO_120 (O_120,N_13047,N_13163);
and UO_121 (O_121,N_12855,N_13262);
and UO_122 (O_122,N_14061,N_13931);
or UO_123 (O_123,N_14598,N_12819);
or UO_124 (O_124,N_12677,N_13791);
and UO_125 (O_125,N_12233,N_14601);
nor UO_126 (O_126,N_12876,N_14256);
nand UO_127 (O_127,N_12355,N_14571);
and UO_128 (O_128,N_13747,N_13244);
nand UO_129 (O_129,N_14366,N_14481);
or UO_130 (O_130,N_12954,N_13703);
and UO_131 (O_131,N_12768,N_13598);
xor UO_132 (O_132,N_14173,N_14795);
nand UO_133 (O_133,N_14631,N_12899);
nand UO_134 (O_134,N_12043,N_13812);
or UO_135 (O_135,N_14194,N_12275);
nand UO_136 (O_136,N_13456,N_12178);
nor UO_137 (O_137,N_14702,N_14383);
nor UO_138 (O_138,N_13059,N_14161);
and UO_139 (O_139,N_14069,N_13635);
nor UO_140 (O_140,N_12435,N_13351);
or UO_141 (O_141,N_14504,N_13147);
nand UO_142 (O_142,N_13170,N_13348);
and UO_143 (O_143,N_14190,N_13434);
xnor UO_144 (O_144,N_12230,N_14343);
nor UO_145 (O_145,N_12722,N_13957);
nand UO_146 (O_146,N_14127,N_13387);
or UO_147 (O_147,N_12391,N_13961);
nand UO_148 (O_148,N_13053,N_12084);
nor UO_149 (O_149,N_12529,N_13403);
xor UO_150 (O_150,N_13802,N_13625);
or UO_151 (O_151,N_14848,N_14563);
nor UO_152 (O_152,N_13005,N_12534);
nand UO_153 (O_153,N_13880,N_13737);
nor UO_154 (O_154,N_13329,N_14241);
nand UO_155 (O_155,N_12254,N_12196);
or UO_156 (O_156,N_14744,N_14048);
or UO_157 (O_157,N_12456,N_14909);
nand UO_158 (O_158,N_13532,N_13319);
and UO_159 (O_159,N_14774,N_14465);
nor UO_160 (O_160,N_12601,N_14216);
nand UO_161 (O_161,N_12377,N_12517);
nor UO_162 (O_162,N_14957,N_14316);
nor UO_163 (O_163,N_14113,N_14359);
or UO_164 (O_164,N_14705,N_14747);
xor UO_165 (O_165,N_14591,N_13349);
nor UO_166 (O_166,N_13413,N_14991);
or UO_167 (O_167,N_12294,N_14660);
or UO_168 (O_168,N_14427,N_12440);
xnor UO_169 (O_169,N_12108,N_14809);
nand UO_170 (O_170,N_13467,N_12310);
nand UO_171 (O_171,N_13665,N_12736);
nor UO_172 (O_172,N_12969,N_13583);
and UO_173 (O_173,N_13058,N_14773);
and UO_174 (O_174,N_13400,N_13767);
or UO_175 (O_175,N_14476,N_13666);
nand UO_176 (O_176,N_12520,N_13485);
xor UO_177 (O_177,N_12569,N_13311);
and UO_178 (O_178,N_12932,N_12896);
nor UO_179 (O_179,N_13251,N_14167);
nand UO_180 (O_180,N_13357,N_12076);
or UO_181 (O_181,N_12542,N_12921);
nand UO_182 (O_182,N_12600,N_12786);
xnor UO_183 (O_183,N_14695,N_12521);
and UO_184 (O_184,N_14042,N_12626);
nor UO_185 (O_185,N_12674,N_12372);
nand UO_186 (O_186,N_14714,N_12603);
xnor UO_187 (O_187,N_12519,N_12441);
or UO_188 (O_188,N_13759,N_12706);
and UO_189 (O_189,N_14012,N_14803);
or UO_190 (O_190,N_12443,N_12071);
nor UO_191 (O_191,N_13618,N_12868);
xnor UO_192 (O_192,N_13850,N_14922);
nor UO_193 (O_193,N_13461,N_13065);
nand UO_194 (O_194,N_13623,N_13496);
or UO_195 (O_195,N_12332,N_12758);
nor UO_196 (O_196,N_12500,N_13612);
nor UO_197 (O_197,N_12426,N_12265);
nor UO_198 (O_198,N_13282,N_13097);
or UO_199 (O_199,N_12986,N_13172);
or UO_200 (O_200,N_12578,N_12323);
xnor UO_201 (O_201,N_13564,N_13418);
and UO_202 (O_202,N_14483,N_14325);
and UO_203 (O_203,N_13798,N_12818);
nand UO_204 (O_204,N_12047,N_13464);
or UO_205 (O_205,N_14493,N_13223);
or UO_206 (O_206,N_13969,N_12078);
xnor UO_207 (O_207,N_12305,N_14373);
or UO_208 (O_208,N_12690,N_13801);
or UO_209 (O_209,N_14911,N_14545);
or UO_210 (O_210,N_13713,N_13112);
or UO_211 (O_211,N_12869,N_14426);
and UO_212 (O_212,N_14520,N_12759);
xnor UO_213 (O_213,N_14249,N_12001);
nor UO_214 (O_214,N_14291,N_14505);
xnor UO_215 (O_215,N_12789,N_12895);
xnor UO_216 (O_216,N_12125,N_12649);
nor UO_217 (O_217,N_12006,N_12809);
nand UO_218 (O_218,N_14100,N_13425);
and UO_219 (O_219,N_13062,N_12908);
nor UO_220 (O_220,N_12495,N_14623);
and UO_221 (O_221,N_12236,N_14669);
and UO_222 (O_222,N_12466,N_14332);
and UO_223 (O_223,N_14778,N_13719);
nor UO_224 (O_224,N_12175,N_14369);
nand UO_225 (O_225,N_12820,N_14972);
nand UO_226 (O_226,N_12136,N_14136);
and UO_227 (O_227,N_13599,N_14568);
xnor UO_228 (O_228,N_14170,N_13094);
nand UO_229 (O_229,N_12988,N_12050);
or UO_230 (O_230,N_12082,N_14864);
or UO_231 (O_231,N_12452,N_12639);
nor UO_232 (O_232,N_12352,N_13190);
and UO_233 (O_233,N_12715,N_12117);
or UO_234 (O_234,N_12222,N_13201);
and UO_235 (O_235,N_13528,N_13657);
and UO_236 (O_236,N_13328,N_14863);
nand UO_237 (O_237,N_13408,N_14847);
or UO_238 (O_238,N_12488,N_13984);
and UO_239 (O_239,N_14455,N_14973);
or UO_240 (O_240,N_14099,N_14333);
nor UO_241 (O_241,N_12981,N_14368);
or UO_242 (O_242,N_14122,N_14370);
xor UO_243 (O_243,N_13478,N_12747);
or UO_244 (O_244,N_14264,N_12145);
or UO_245 (O_245,N_13444,N_14507);
xnor UO_246 (O_246,N_14941,N_13310);
and UO_247 (O_247,N_12183,N_13108);
or UO_248 (O_248,N_12270,N_12198);
or UO_249 (O_249,N_13813,N_13250);
nor UO_250 (O_250,N_13705,N_12916);
xnor UO_251 (O_251,N_12015,N_14005);
or UO_252 (O_252,N_12327,N_12679);
nor UO_253 (O_253,N_14549,N_12562);
or UO_254 (O_254,N_12100,N_13613);
and UO_255 (O_255,N_13090,N_14936);
nand UO_256 (O_256,N_12064,N_13687);
nor UO_257 (O_257,N_14907,N_13234);
or UO_258 (O_258,N_12427,N_12429);
nor UO_259 (O_259,N_13894,N_14566);
nand UO_260 (O_260,N_14897,N_12831);
or UO_261 (O_261,N_13012,N_13002);
nor UO_262 (O_262,N_12235,N_12374);
xor UO_263 (O_263,N_13240,N_14689);
nand UO_264 (O_264,N_13474,N_12735);
nor UO_265 (O_265,N_13826,N_13091);
nor UO_266 (O_266,N_14386,N_14641);
and UO_267 (O_267,N_14971,N_13260);
or UO_268 (O_268,N_14596,N_14624);
or UO_269 (O_269,N_14769,N_14078);
or UO_270 (O_270,N_12246,N_12846);
and UO_271 (O_271,N_12858,N_14887);
and UO_272 (O_272,N_14914,N_13994);
and UO_273 (O_273,N_13362,N_12477);
xor UO_274 (O_274,N_14196,N_14199);
nor UO_275 (O_275,N_14954,N_14102);
nor UO_276 (O_276,N_12189,N_12319);
xor UO_277 (O_277,N_12567,N_13169);
or UO_278 (O_278,N_13536,N_14396);
nand UO_279 (O_279,N_14443,N_13207);
and UO_280 (O_280,N_14697,N_13773);
xnor UO_281 (O_281,N_13906,N_14564);
or UO_282 (O_282,N_12850,N_14625);
and UO_283 (O_283,N_12166,N_14385);
nand UO_284 (O_284,N_14721,N_14462);
nor UO_285 (O_285,N_12062,N_14965);
and UO_286 (O_286,N_13061,N_13985);
or UO_287 (O_287,N_14717,N_12396);
or UO_288 (O_288,N_12907,N_14619);
nand UO_289 (O_289,N_13324,N_14929);
nand UO_290 (O_290,N_12862,N_13189);
nand UO_291 (O_291,N_13560,N_13858);
nand UO_292 (O_292,N_13521,N_12207);
xor UO_293 (O_293,N_12240,N_14323);
nor UO_294 (O_294,N_12901,N_12425);
nor UO_295 (O_295,N_12402,N_13028);
and UO_296 (O_296,N_14447,N_14424);
and UO_297 (O_297,N_12285,N_14021);
nor UO_298 (O_298,N_12561,N_14787);
or UO_299 (O_299,N_12741,N_14019);
nand UO_300 (O_300,N_14634,N_12289);
and UO_301 (O_301,N_13762,N_12577);
nand UO_302 (O_302,N_13293,N_14094);
or UO_303 (O_303,N_13437,N_14354);
xnor UO_304 (O_304,N_13644,N_12540);
or UO_305 (O_305,N_13075,N_12770);
nand UO_306 (O_306,N_14213,N_13734);
nor UO_307 (O_307,N_14902,N_12924);
nor UO_308 (O_308,N_12952,N_14677);
xnor UO_309 (O_309,N_13219,N_14184);
nor UO_310 (O_310,N_13676,N_13871);
xnor UO_311 (O_311,N_14480,N_14763);
nand UO_312 (O_312,N_14265,N_14489);
or UO_313 (O_313,N_14812,N_13427);
nor UO_314 (O_314,N_13982,N_14144);
or UO_315 (O_315,N_14952,N_14111);
nand UO_316 (O_316,N_14351,N_13950);
nor UO_317 (O_317,N_12069,N_13284);
nor UO_318 (O_318,N_13459,N_12152);
nand UO_319 (O_319,N_14303,N_12266);
nand UO_320 (O_320,N_13852,N_12010);
xnor UO_321 (O_321,N_13176,N_13764);
or UO_322 (O_322,N_13963,N_13504);
nor UO_323 (O_323,N_12163,N_14289);
and UO_324 (O_324,N_14225,N_14903);
or UO_325 (O_325,N_12545,N_14251);
and UO_326 (O_326,N_14758,N_13516);
or UO_327 (O_327,N_12493,N_14898);
nor UO_328 (O_328,N_12056,N_13054);
or UO_329 (O_329,N_12875,N_13992);
and UO_330 (O_330,N_13026,N_12321);
and UO_331 (O_331,N_14701,N_13229);
or UO_332 (O_332,N_14526,N_14374);
xnor UO_333 (O_333,N_13182,N_13898);
or UO_334 (O_334,N_14703,N_13168);
or UO_335 (O_335,N_14263,N_12264);
xnor UO_336 (O_336,N_13882,N_14457);
and UO_337 (O_337,N_12705,N_12020);
nand UO_338 (O_338,N_14927,N_13827);
xor UO_339 (O_339,N_14070,N_14015);
and UO_340 (O_340,N_14267,N_13517);
nor UO_341 (O_341,N_14846,N_13872);
or UO_342 (O_342,N_13786,N_14642);
nand UO_343 (O_343,N_14209,N_13046);
xnor UO_344 (O_344,N_12143,N_12810);
nor UO_345 (O_345,N_14756,N_14056);
or UO_346 (O_346,N_12693,N_14776);
and UO_347 (O_347,N_12953,N_12421);
nand UO_348 (O_348,N_13505,N_14635);
xor UO_349 (O_349,N_13345,N_12547);
or UO_350 (O_350,N_14553,N_14007);
nand UO_351 (O_351,N_14032,N_14814);
and UO_352 (O_352,N_12536,N_14135);
nor UO_353 (O_353,N_14273,N_12919);
xor UO_354 (O_354,N_14996,N_13326);
nand UO_355 (O_355,N_12070,N_12090);
or UO_356 (O_356,N_14686,N_13268);
nand UO_357 (O_357,N_12822,N_13245);
nand UO_358 (O_358,N_12200,N_14630);
nor UO_359 (O_359,N_12737,N_13079);
nor UO_360 (O_360,N_12118,N_12259);
and UO_361 (O_361,N_13368,N_12676);
nor UO_362 (O_362,N_14453,N_14074);
or UO_363 (O_363,N_14737,N_13333);
or UO_364 (O_364,N_14533,N_12093);
nor UO_365 (O_365,N_12510,N_14046);
nand UO_366 (O_366,N_13033,N_12272);
nor UO_367 (O_367,N_12847,N_13991);
and UO_368 (O_368,N_14766,N_12113);
nor UO_369 (O_369,N_14708,N_13752);
or UO_370 (O_370,N_14430,N_14274);
nand UO_371 (O_371,N_13073,N_14868);
or UO_372 (O_372,N_14859,N_13267);
and UO_373 (O_373,N_14439,N_12672);
or UO_374 (O_374,N_14529,N_13529);
or UO_375 (O_375,N_14692,N_12994);
nor UO_376 (O_376,N_14201,N_13565);
nor UO_377 (O_377,N_12696,N_14726);
and UO_378 (O_378,N_14337,N_14732);
nand UO_379 (O_379,N_14017,N_13470);
or UO_380 (O_380,N_12879,N_13771);
xnor UO_381 (O_381,N_13162,N_13748);
or UO_382 (O_382,N_14978,N_12606);
nor UO_383 (O_383,N_14304,N_12774);
nand UO_384 (O_384,N_13939,N_13398);
nor UO_385 (O_385,N_13192,N_14114);
nor UO_386 (O_386,N_12106,N_14335);
nand UO_387 (O_387,N_12571,N_13161);
nor UO_388 (O_388,N_14284,N_12142);
nor UO_389 (O_389,N_14813,N_13394);
xnor UO_390 (O_390,N_14442,N_13757);
nor UO_391 (O_391,N_13256,N_14458);
or UO_392 (O_392,N_14531,N_13556);
and UO_393 (O_393,N_12837,N_12409);
nor UO_394 (O_394,N_13366,N_13851);
nand UO_395 (O_395,N_13379,N_13029);
and UO_396 (O_396,N_13453,N_14347);
nor UO_397 (O_397,N_12619,N_14674);
nand UO_398 (O_398,N_14752,N_13664);
and UO_399 (O_399,N_12457,N_13060);
nor UO_400 (O_400,N_12138,N_13297);
nor UO_401 (O_401,N_12229,N_12691);
nor UO_402 (O_402,N_12533,N_14252);
and UO_403 (O_403,N_12564,N_12782);
or UO_404 (O_404,N_14711,N_14467);
or UO_405 (O_405,N_14935,N_14821);
nand UO_406 (O_406,N_12021,N_13376);
or UO_407 (O_407,N_12135,N_12422);
or UO_408 (O_408,N_13224,N_12337);
nand UO_409 (O_409,N_14472,N_12881);
nand UO_410 (O_410,N_13672,N_13327);
or UO_411 (O_411,N_14228,N_13180);
or UO_412 (O_412,N_13130,N_14607);
and UO_413 (O_413,N_13248,N_14326);
and UO_414 (O_414,N_12357,N_13194);
or UO_415 (O_415,N_12194,N_14626);
and UO_416 (O_416,N_12394,N_14822);
and UO_417 (O_417,N_12417,N_13361);
or UO_418 (O_418,N_14924,N_12215);
and UO_419 (O_419,N_12773,N_13399);
nor UO_420 (O_420,N_13380,N_12346);
nor UO_421 (O_421,N_14120,N_12019);
or UO_422 (O_422,N_13006,N_12527);
and UO_423 (O_423,N_12008,N_14157);
nand UO_424 (O_424,N_14400,N_13578);
xor UO_425 (O_425,N_14479,N_14245);
nand UO_426 (O_426,N_13895,N_12886);
and UO_427 (O_427,N_13213,N_13304);
or UO_428 (O_428,N_12089,N_12449);
nor UO_429 (O_429,N_12300,N_12641);
or UO_430 (O_430,N_13228,N_12729);
nor UO_431 (O_431,N_13620,N_14098);
and UO_432 (O_432,N_14254,N_14150);
nand UO_433 (O_433,N_13829,N_12359);
nand UO_434 (O_434,N_12878,N_13406);
nand UO_435 (O_435,N_14579,N_12037);
nand UO_436 (O_436,N_14067,N_12046);
and UO_437 (O_437,N_14799,N_14334);
or UO_438 (O_438,N_14461,N_14110);
nor UO_439 (O_439,N_12499,N_12146);
or UO_440 (O_440,N_14878,N_12585);
or UO_441 (O_441,N_13291,N_14387);
nor UO_442 (O_442,N_13071,N_12042);
nand UO_443 (O_443,N_14299,N_14949);
and UO_444 (O_444,N_14151,N_12088);
nand UO_445 (O_445,N_13518,N_12646);
nor UO_446 (O_446,N_12877,N_12308);
xor UO_447 (O_447,N_12249,N_14140);
and UO_448 (O_448,N_14746,N_12731);
nor UO_449 (O_449,N_14904,N_12306);
and UO_450 (O_450,N_13832,N_12077);
xor UO_451 (O_451,N_12699,N_12832);
nor UO_452 (O_452,N_13525,N_12854);
or UO_453 (O_453,N_13508,N_12392);
or UO_454 (O_454,N_12928,N_13806);
nand UO_455 (O_455,N_13457,N_13374);
and UO_456 (O_456,N_14389,N_14552);
nand UO_457 (O_457,N_14593,N_12325);
or UO_458 (O_458,N_13511,N_12111);
nand UO_459 (O_459,N_14874,N_14469);
and UO_460 (O_460,N_14257,N_14066);
and UO_461 (O_461,N_14108,N_13736);
nor UO_462 (O_462,N_14976,N_14054);
nor UO_463 (O_463,N_12976,N_13247);
nand UO_464 (O_464,N_14095,N_14853);
and UO_465 (O_465,N_14464,N_12804);
nor UO_466 (O_466,N_12351,N_12378);
xor UO_467 (O_467,N_14754,N_14423);
and UO_468 (O_468,N_14057,N_13402);
nor UO_469 (O_469,N_13879,N_12282);
or UO_470 (O_470,N_14837,N_13550);
or UO_471 (O_471,N_13935,N_14008);
nand UO_472 (O_472,N_14205,N_13548);
nor UO_473 (O_473,N_13477,N_12170);
nand UO_474 (O_474,N_14819,N_14830);
xor UO_475 (O_475,N_14834,N_14168);
nand UO_476 (O_476,N_14637,N_13569);
nand UO_477 (O_477,N_12959,N_14329);
or UO_478 (O_478,N_13111,N_12623);
and UO_479 (O_479,N_12867,N_14006);
and UO_480 (O_480,N_14506,N_14503);
nand UO_481 (O_481,N_14206,N_14156);
or UO_482 (O_482,N_13308,N_14939);
and UO_483 (O_483,N_14930,N_13171);
or UO_484 (O_484,N_14432,N_12903);
nor UO_485 (O_485,N_12673,N_12256);
nand UO_486 (O_486,N_12239,N_12036);
nand UO_487 (O_487,N_14650,N_13049);
nor UO_488 (O_488,N_12217,N_12320);
or UO_489 (O_489,N_12389,N_13756);
and UO_490 (O_490,N_14722,N_12386);
nor UO_491 (O_491,N_12843,N_14159);
and UO_492 (O_492,N_13946,N_12581);
nand UO_493 (O_493,N_13448,N_13078);
and UO_494 (O_494,N_13639,N_14215);
and UO_495 (O_495,N_14912,N_14817);
nor UO_496 (O_496,N_14362,N_12432);
xor UO_497 (O_497,N_14730,N_13346);
nor UO_498 (O_498,N_13303,N_13519);
nor UO_499 (O_499,N_12293,N_12927);
or UO_500 (O_500,N_14232,N_12045);
or UO_501 (O_501,N_14306,N_14189);
nand UO_502 (O_502,N_13114,N_14818);
nor UO_503 (O_503,N_12383,N_13707);
and UO_504 (O_504,N_12995,N_14371);
or UO_505 (O_505,N_13367,N_14154);
nand UO_506 (O_506,N_14283,N_12029);
nor UO_507 (O_507,N_13021,N_13498);
nor UO_508 (O_508,N_14893,N_13634);
or UO_509 (O_509,N_14524,N_14118);
and UO_510 (O_510,N_14183,N_12962);
and UO_511 (O_511,N_14966,N_12479);
xor UO_512 (O_512,N_13967,N_14578);
nand UO_513 (O_513,N_13746,N_14792);
xor UO_514 (O_514,N_14026,N_14644);
nor UO_515 (O_515,N_14699,N_14292);
nand UO_516 (O_516,N_12686,N_13204);
nand UO_517 (O_517,N_14614,N_12551);
or UO_518 (O_518,N_13476,N_14923);
and UO_519 (O_519,N_14671,N_14459);
nor UO_520 (O_520,N_14440,N_13663);
and UO_521 (O_521,N_14690,N_14743);
nor UO_522 (O_522,N_13706,N_13123);
and UO_523 (O_523,N_14885,N_14338);
nand UO_524 (O_524,N_14694,N_12472);
nand UO_525 (O_525,N_12902,N_14079);
xor UO_526 (O_526,N_13119,N_12340);
or UO_527 (O_527,N_12148,N_12073);
or UO_528 (O_528,N_13986,N_14975);
nor UO_529 (O_529,N_12025,N_13735);
nand UO_530 (O_530,N_13236,N_12920);
nand UO_531 (O_531,N_13590,N_14024);
or UO_532 (O_532,N_13604,N_13653);
nand UO_533 (O_533,N_12284,N_12350);
nor UO_534 (O_534,N_14065,N_12756);
or UO_535 (O_535,N_13103,N_13693);
or UO_536 (O_536,N_12127,N_14655);
nor UO_537 (O_537,N_13727,N_14125);
nor UO_538 (O_538,N_13729,N_13976);
or UO_539 (O_539,N_13494,N_13622);
nand UO_540 (O_540,N_14039,N_12168);
and UO_541 (O_541,N_13808,N_12816);
nor UO_542 (O_542,N_14123,N_13159);
nor UO_543 (O_543,N_14828,N_13661);
nand UO_544 (O_544,N_13100,N_12761);
nand UO_545 (O_545,N_13125,N_13557);
and UO_546 (O_546,N_12384,N_13793);
nor UO_547 (O_547,N_12765,N_14765);
or UO_548 (O_548,N_14169,N_14038);
nand UO_549 (O_549,N_14687,N_14595);
and UO_550 (O_550,N_13272,N_12347);
or UO_551 (O_551,N_14988,N_14097);
or UO_552 (O_552,N_14133,N_14090);
and UO_553 (O_553,N_13372,N_14137);
nand UO_554 (O_554,N_13299,N_12369);
xor UO_555 (O_555,N_13777,N_14415);
or UO_556 (O_556,N_13924,N_13377);
nor UO_557 (O_557,N_13211,N_14772);
nand UO_558 (O_558,N_14380,N_13198);
nor UO_559 (O_559,N_13350,N_12982);
nor UO_560 (O_560,N_14384,N_13086);
or UO_561 (O_561,N_14648,N_14739);
and UO_562 (O_562,N_13109,N_12034);
nand UO_563 (O_563,N_14062,N_14485);
and UO_564 (O_564,N_13809,N_12890);
or UO_565 (O_565,N_12748,N_12802);
nor UO_566 (O_566,N_13241,N_13627);
nand UO_567 (O_567,N_12496,N_12212);
nand UO_568 (O_568,N_12531,N_13393);
xnor UO_569 (O_569,N_14145,N_14035);
nor UO_570 (O_570,N_13157,N_13088);
or UO_571 (O_571,N_14622,N_14022);
or UO_572 (O_572,N_13421,N_14984);
and UO_573 (O_573,N_12420,N_13700);
or UO_574 (O_574,N_12678,N_13181);
or UO_575 (O_575,N_13933,N_12027);
or UO_576 (O_576,N_14002,N_12505);
and UO_577 (O_577,N_12016,N_14959);
nand UO_578 (O_578,N_12634,N_14647);
nand UO_579 (O_579,N_13460,N_13905);
nand UO_580 (O_580,N_12147,N_14155);
or UO_581 (O_581,N_14059,N_13051);
nand UO_582 (O_582,N_12609,N_12938);
or UO_583 (O_583,N_14148,N_14314);
nand UO_584 (O_584,N_13405,N_13295);
nand UO_585 (O_585,N_14696,N_13975);
nand UO_586 (O_586,N_14796,N_14719);
xnor UO_587 (O_587,N_12398,N_12035);
nor UO_588 (O_588,N_12637,N_12710);
nor UO_589 (O_589,N_13135,N_12214);
or UO_590 (O_590,N_12436,N_13811);
or UO_591 (O_591,N_13233,N_14011);
xor UO_592 (O_592,N_14282,N_13810);
nand UO_593 (O_593,N_12974,N_13269);
nor UO_594 (O_594,N_13120,N_13129);
nor UO_595 (O_595,N_12410,N_13908);
and UO_596 (O_596,N_13154,N_14033);
and UO_597 (O_597,N_12640,N_13214);
and UO_598 (O_598,N_12838,N_14588);
xnor UO_599 (O_599,N_12155,N_12889);
xor UO_600 (O_600,N_12133,N_13506);
nand UO_601 (O_601,N_12627,N_13781);
nor UO_602 (O_602,N_13289,N_14129);
or UO_603 (O_603,N_13831,N_14301);
or UO_604 (O_604,N_14780,N_14610);
xnor UO_605 (O_605,N_14116,N_14044);
and UO_606 (O_606,N_14270,N_12644);
nand UO_607 (O_607,N_14891,N_13617);
or UO_608 (O_608,N_13024,N_12102);
or UO_609 (O_609,N_13745,N_12299);
nand UO_610 (O_610,N_14296,N_14589);
nand UO_611 (O_611,N_12271,N_13765);
and UO_612 (O_612,N_13589,N_14548);
nor UO_613 (O_613,N_14557,N_12780);
or UO_614 (O_614,N_12257,N_14475);
nand UO_615 (O_615,N_14040,N_12475);
or UO_616 (O_616,N_14816,N_14842);
or UO_617 (O_617,N_13429,N_14709);
xor UO_618 (O_618,N_14246,N_14926);
or UO_619 (O_619,N_14760,N_14544);
nand UO_620 (O_620,N_12482,N_14919);
and UO_621 (O_621,N_13956,N_13164);
or UO_622 (O_622,N_12909,N_14147);
and UO_623 (O_623,N_13277,N_13552);
nor UO_624 (O_624,N_14171,N_14071);
and UO_625 (O_625,N_12891,N_14712);
or UO_626 (O_626,N_14356,N_13188);
nor UO_627 (O_627,N_14883,N_13203);
or UO_628 (O_628,N_13775,N_14495);
and UO_629 (O_629,N_13034,N_13035);
xor UO_630 (O_630,N_13412,N_14239);
nand UO_631 (O_631,N_14016,N_13270);
nor UO_632 (O_632,N_13352,N_13597);
and UO_633 (O_633,N_12453,N_12629);
nor UO_634 (O_634,N_13927,N_12094);
nand UO_635 (O_635,N_13347,N_14676);
nand UO_636 (O_636,N_13473,N_12361);
nand UO_637 (O_637,N_14318,N_13916);
or UO_638 (O_638,N_13415,N_13731);
or UO_639 (O_639,N_13714,N_13365);
xnor UO_640 (O_640,N_12524,N_13728);
and UO_641 (O_641,N_12512,N_14288);
nor UO_642 (O_642,N_12395,N_12931);
nand UO_643 (O_643,N_14278,N_13041);
nor UO_644 (O_644,N_13726,N_12835);
or UO_645 (O_645,N_14510,N_14290);
or UO_646 (O_646,N_14679,N_12568);
nor UO_647 (O_647,N_14740,N_14163);
or UO_648 (O_648,N_12408,N_12702);
nand UO_649 (O_649,N_14961,N_12785);
nand UO_650 (O_650,N_14811,N_12615);
nand UO_651 (O_651,N_13484,N_12946);
and UO_652 (O_652,N_14025,N_13083);
or UO_653 (O_653,N_12277,N_13840);
or UO_654 (O_654,N_14072,N_13804);
xor UO_655 (O_655,N_13067,N_12742);
and UO_656 (O_656,N_13656,N_13364);
nand UO_657 (O_657,N_13834,N_12588);
or UO_658 (O_658,N_14915,N_12338);
and UO_659 (O_659,N_12525,N_14208);
nand UO_660 (O_660,N_12281,N_14195);
nand UO_661 (O_661,N_13964,N_12852);
nor UO_662 (O_662,N_14018,N_12373);
nand UO_663 (O_663,N_12176,N_12522);
xnor UO_664 (O_664,N_12213,N_14867);
and UO_665 (O_665,N_13940,N_13370);
nand UO_666 (O_666,N_14317,N_12984);
nand UO_667 (O_667,N_12328,N_12628);
and UO_668 (O_668,N_13610,N_12762);
and UO_669 (O_669,N_12468,N_14761);
xor UO_670 (O_670,N_12631,N_14050);
nor UO_671 (O_671,N_14670,N_14227);
and UO_672 (O_672,N_14166,N_12790);
nand UO_673 (O_673,N_13980,N_14720);
nor UO_674 (O_674,N_14609,N_12024);
and UO_675 (O_675,N_13397,N_14890);
xor UO_676 (O_676,N_12797,N_12059);
xnor UO_677 (O_677,N_13632,N_13842);
and UO_678 (O_678,N_14536,N_12393);
or UO_679 (O_679,N_13692,N_12013);
xor UO_680 (O_680,N_12085,N_14350);
nor UO_681 (O_681,N_13534,N_13186);
nor UO_682 (O_682,N_12546,N_14951);
or UO_683 (O_683,N_14994,N_13948);
xor UO_684 (O_684,N_12871,N_13743);
and UO_685 (O_685,N_12549,N_12801);
nand UO_686 (O_686,N_13889,N_14188);
or UO_687 (O_687,N_12095,N_12776);
nor UO_688 (O_688,N_13452,N_13690);
nand UO_689 (O_689,N_14748,N_13332);
nand UO_690 (O_690,N_14081,N_12853);
xnor UO_691 (O_691,N_14107,N_13337);
or UO_692 (O_692,N_12007,N_12554);
or UO_693 (O_693,N_13680,N_13626);
xor UO_694 (O_694,N_13580,N_13725);
or UO_695 (O_695,N_13962,N_13134);
or UO_696 (O_696,N_13921,N_13227);
and UO_697 (O_697,N_12914,N_12906);
and UO_698 (O_698,N_13118,N_14960);
or UO_699 (O_699,N_13253,N_13140);
nor UO_700 (O_700,N_13540,N_13805);
or UO_701 (O_701,N_14367,N_13003);
xnor UO_702 (O_702,N_13279,N_14341);
or UO_703 (O_703,N_13899,N_14238);
nand UO_704 (O_704,N_14698,N_12851);
nand UO_705 (O_705,N_14327,N_12080);
nand UO_706 (O_706,N_13020,N_12764);
nor UO_707 (O_707,N_12197,N_12949);
xnor UO_708 (O_708,N_13156,N_14298);
nor UO_709 (O_709,N_14049,N_12783);
nor UO_710 (O_710,N_12508,N_14352);
and UO_711 (O_711,N_12366,N_13789);
nand UO_712 (O_712,N_13179,N_14945);
or UO_713 (O_713,N_14782,N_13524);
or UO_714 (O_714,N_13208,N_14639);
and UO_715 (O_715,N_12656,N_14734);
nand UO_716 (O_716,N_12716,N_12866);
nor UO_717 (O_717,N_13616,N_14790);
or UO_718 (O_718,N_12375,N_13682);
and UO_719 (O_719,N_13642,N_12442);
nor UO_720 (O_720,N_13951,N_14434);
nor UO_721 (O_721,N_13419,N_12526);
and UO_722 (O_722,N_13433,N_14750);
nand UO_723 (O_723,N_12484,N_12597);
or UO_724 (O_724,N_14838,N_13862);
or UO_725 (O_725,N_14900,N_14603);
nor UO_726 (O_726,N_12150,N_14281);
and UO_727 (O_727,N_14103,N_12806);
xor UO_728 (O_728,N_13462,N_14857);
and UO_729 (O_729,N_13685,N_14535);
xnor UO_730 (O_730,N_14800,N_13263);
or UO_731 (O_731,N_12199,N_13280);
nor UO_732 (O_732,N_13391,N_14691);
nand UO_733 (O_733,N_14681,N_14500);
and UO_734 (O_734,N_12642,N_12424);
xnor UO_735 (O_735,N_12462,N_14083);
or UO_736 (O_736,N_14804,N_12412);
and UO_737 (O_737,N_13040,N_14775);
nand UO_738 (O_738,N_12297,N_13334);
nand UO_739 (O_739,N_12274,N_14037);
nor UO_740 (O_740,N_14003,N_13331);
and UO_741 (O_741,N_13152,N_12942);
or UO_742 (O_742,N_13960,N_13575);
or UO_743 (O_743,N_12324,N_12000);
or UO_744 (O_744,N_14770,N_13925);
nor UO_745 (O_745,N_13439,N_14134);
and UO_746 (O_746,N_13301,N_14404);
or UO_747 (O_747,N_14985,N_12552);
nand UO_748 (O_748,N_12811,N_13596);
nor UO_749 (O_749,N_14947,N_14418);
and UO_750 (O_750,N_12354,N_13937);
and UO_751 (O_751,N_13999,N_13037);
and UO_752 (O_752,N_12965,N_12912);
or UO_753 (O_753,N_13893,N_13546);
nor UO_754 (O_754,N_12329,N_12494);
nor UO_755 (O_755,N_14731,N_14096);
nand UO_756 (O_756,N_14585,N_13709);
nand UO_757 (O_757,N_13490,N_13716);
nand UO_758 (O_758,N_14365,N_14521);
xnor UO_759 (O_759,N_12356,N_14092);
nand UO_760 (O_760,N_13582,N_14875);
nand UO_761 (O_761,N_12593,N_14943);
nor UO_762 (O_762,N_13081,N_14586);
nand UO_763 (O_763,N_14582,N_14328);
or UO_764 (O_764,N_13369,N_14478);
nor UO_765 (O_765,N_13278,N_12224);
nand UO_766 (O_766,N_12662,N_13146);
or UO_767 (O_767,N_13573,N_13763);
xnor UO_768 (O_768,N_13143,N_12192);
and UO_769 (O_769,N_14575,N_14446);
or UO_770 (O_770,N_14573,N_14995);
nor UO_771 (O_771,N_12733,N_12112);
nor UO_772 (O_772,N_13958,N_13857);
nand UO_773 (O_773,N_14836,N_14313);
or UO_774 (O_774,N_12486,N_13482);
nor UO_775 (O_775,N_12712,N_14666);
and UO_776 (O_776,N_12718,N_12491);
and UO_777 (O_777,N_12583,N_14363);
or UO_778 (O_778,N_12091,N_14831);
nand UO_779 (O_779,N_14302,N_14810);
nor UO_780 (O_780,N_12513,N_14768);
or UO_781 (O_781,N_14181,N_12925);
nand UO_782 (O_782,N_14207,N_13652);
or UO_783 (O_783,N_12675,N_13202);
nand UO_784 (O_784,N_14222,N_14353);
nand UO_785 (O_785,N_13815,N_14534);
nand UO_786 (O_786,N_14621,N_14477);
nor UO_787 (O_787,N_12605,N_12709);
xnor UO_788 (O_788,N_12523,N_14844);
or UO_789 (O_789,N_13601,N_12387);
nor UO_790 (O_790,N_12796,N_14080);
nor UO_791 (O_791,N_14235,N_14659);
nand UO_792 (O_792,N_14030,N_13608);
nor UO_793 (O_793,N_13423,N_12124);
nor UO_794 (O_794,N_13848,N_12251);
nand UO_795 (O_795,N_13150,N_13835);
or UO_796 (O_796,N_14913,N_13655);
xnor UO_797 (O_797,N_14089,N_14063);
nand UO_798 (O_798,N_12798,N_13064);
nand UO_799 (O_799,N_14394,N_14987);
nand UO_800 (O_800,N_13285,N_13174);
or UO_801 (O_801,N_13515,N_12258);
nor UO_802 (O_802,N_12471,N_14488);
nor UO_803 (O_803,N_14445,N_12130);
xor UO_804 (O_804,N_13684,N_12732);
nand UO_805 (O_805,N_13151,N_13538);
and UO_806 (O_806,N_12829,N_12744);
nor UO_807 (O_807,N_14755,N_13283);
nor UO_808 (O_808,N_14277,N_13675);
xor UO_809 (O_809,N_12680,N_14513);
and UO_810 (O_810,N_13730,N_12086);
xor UO_811 (O_811,N_13316,N_12057);
nor UO_812 (O_812,N_12087,N_13670);
xor UO_813 (O_813,N_13662,N_13878);
nand UO_814 (O_814,N_14683,N_13416);
and UO_815 (O_815,N_13196,N_12447);
or UO_816 (O_816,N_14889,N_12219);
or UO_817 (O_817,N_14360,N_13259);
nand UO_818 (O_818,N_12671,N_12570);
and UO_819 (O_819,N_13440,N_13510);
xnor UO_820 (O_820,N_14522,N_12334);
nand UO_821 (O_821,N_12645,N_12014);
xor UO_822 (O_822,N_12565,N_13138);
and UO_823 (O_823,N_12295,N_14223);
or UO_824 (O_824,N_13335,N_14682);
and UO_825 (O_825,N_12985,N_13115);
nand UO_826 (O_826,N_14132,N_13979);
nor UO_827 (O_827,N_13489,N_14916);
and UO_828 (O_828,N_13401,N_14981);
nor UO_829 (O_829,N_13555,N_14617);
and UO_830 (O_830,N_13226,N_12655);
nand UO_831 (O_831,N_14105,N_12607);
and UO_832 (O_832,N_12726,N_14937);
and UO_833 (O_833,N_12772,N_12668);
nand UO_834 (O_834,N_14086,N_14892);
nand UO_835 (O_835,N_12126,N_12654);
nor UO_836 (O_836,N_14115,N_13153);
nor UO_837 (O_837,N_14829,N_13720);
and UO_838 (O_838,N_12880,N_14794);
nor UO_839 (O_839,N_13844,N_14494);
and UO_840 (O_840,N_13859,N_14855);
nand UO_841 (O_841,N_14058,N_13131);
nor UO_842 (O_842,N_13302,N_14498);
and UO_843 (O_843,N_12857,N_13336);
and UO_844 (O_844,N_12399,N_14075);
and UO_845 (O_845,N_14527,N_13847);
xnor UO_846 (O_846,N_14989,N_13928);
or UO_847 (O_847,N_12757,N_12380);
xnor UO_848 (O_848,N_14031,N_12620);
nor UO_849 (O_849,N_13760,N_13592);
nand UO_850 (O_850,N_12967,N_13124);
nor UO_851 (O_851,N_12157,N_13242);
nand UO_852 (O_852,N_14992,N_13074);
and UO_853 (O_853,N_13868,N_13874);
nor UO_854 (O_854,N_12563,N_12624);
nand UO_855 (O_855,N_13903,N_14388);
or UO_856 (O_856,N_13619,N_12390);
and UO_857 (O_857,N_14895,N_13526);
nand UO_858 (O_858,N_13993,N_13649);
and UO_859 (O_859,N_14745,N_12298);
or UO_860 (O_860,N_13629,N_12225);
nand UO_861 (O_861,N_12518,N_12683);
and UO_862 (O_862,N_12267,N_12904);
nor UO_863 (O_863,N_12633,N_14646);
or UO_864 (O_864,N_13235,N_13197);
nor UO_865 (O_865,N_12506,N_13359);
nand UO_866 (O_866,N_12548,N_13697);
nand UO_867 (O_867,N_12253,N_12874);
nor UO_868 (O_868,N_12929,N_13683);
nand UO_869 (O_869,N_13691,N_12172);
and UO_870 (O_870,N_14574,N_14806);
xnor UO_871 (O_871,N_12966,N_12193);
or UO_872 (O_872,N_13952,N_12413);
or UO_873 (O_873,N_14433,N_12511);
and UO_874 (O_874,N_14977,N_14850);
nand UO_875 (O_875,N_14602,N_14308);
or UO_876 (O_876,N_13265,N_14165);
nand UO_877 (O_877,N_13420,N_12535);
or UO_878 (O_878,N_14841,N_14091);
and UO_879 (O_879,N_14872,N_12515);
nand UO_880 (O_880,N_12079,N_14615);
and UO_881 (O_881,N_12186,N_14407);
nand UO_882 (O_882,N_13501,N_12803);
nand UO_883 (O_883,N_12316,N_12317);
xor UO_884 (O_884,N_12030,N_14509);
xnor UO_885 (O_885,N_14590,N_13258);
and UO_886 (O_886,N_13018,N_14441);
or UO_887 (O_887,N_13107,N_14876);
nand UO_888 (O_888,N_14236,N_12788);
and UO_889 (O_889,N_13917,N_12934);
or UO_890 (O_890,N_13650,N_13896);
nand UO_891 (O_891,N_13855,N_12115);
nor UO_892 (O_892,N_14516,N_12237);
and UO_893 (O_893,N_13866,N_12280);
nor UO_894 (O_894,N_14403,N_14940);
nand UO_895 (O_895,N_13249,N_13441);
nand UO_896 (O_896,N_14082,N_14474);
nand UO_897 (O_897,N_12861,N_14986);
or UO_898 (O_898,N_12314,N_13739);
and UO_899 (O_899,N_12368,N_13144);
or UO_900 (O_900,N_12800,N_13022);
nor UO_901 (O_901,N_13216,N_12576);
and UO_902 (O_902,N_13867,N_14409);
nand UO_903 (O_903,N_12066,N_12652);
or UO_904 (O_904,N_12401,N_13104);
nor UO_905 (O_905,N_14014,N_14851);
xnor UO_906 (O_906,N_14402,N_13891);
nor UO_907 (O_907,N_12828,N_12528);
nor UO_908 (O_908,N_13486,N_14175);
and UO_909 (O_909,N_14738,N_13479);
or UO_910 (O_910,N_14348,N_12977);
or UO_911 (O_911,N_12180,N_14771);
nor UO_912 (O_912,N_12701,N_13343);
nand UO_913 (O_913,N_13833,N_14473);
xor UO_914 (O_914,N_13977,N_12053);
or UO_915 (O_915,N_12582,N_14192);
nand UO_916 (O_916,N_12713,N_12721);
and UO_917 (O_917,N_12584,N_14395);
nand UO_918 (O_918,N_14456,N_12687);
nor UO_919 (O_919,N_14193,N_12698);
xor UO_920 (O_920,N_13671,N_13183);
or UO_921 (O_921,N_14088,N_13093);
and UO_922 (O_922,N_14820,N_14993);
nor UO_923 (O_923,N_14253,N_12205);
nor UO_924 (O_924,N_14587,N_14414);
or UO_925 (O_925,N_13704,N_13901);
and UO_926 (O_926,N_14320,N_14259);
nand UO_927 (O_927,N_12291,N_13092);
and UO_928 (O_928,N_14198,N_14153);
and UO_929 (O_929,N_12121,N_13606);
and UO_930 (O_930,N_12559,N_14164);
nand UO_931 (O_931,N_13015,N_13014);
xnor UO_932 (O_932,N_12075,N_12989);
xor UO_933 (O_933,N_13527,N_13797);
or UO_934 (O_934,N_12717,N_14753);
xor UO_935 (O_935,N_14979,N_14512);
and UO_936 (O_936,N_13570,N_12103);
or UO_937 (O_937,N_14345,N_12658);
nand UO_938 (O_938,N_14718,N_14186);
nor UO_939 (O_939,N_12211,N_13481);
nor UO_940 (O_940,N_12238,N_13539);
and UO_941 (O_941,N_12231,N_12541);
nand UO_942 (O_942,N_12532,N_13586);
nand UO_943 (O_943,N_12159,N_12463);
xnor UO_944 (O_944,N_13116,N_13178);
nand UO_945 (O_945,N_14962,N_13696);
nand UO_946 (O_946,N_14729,N_12017);
nand UO_947 (O_947,N_14849,N_13750);
nand UO_948 (O_948,N_12779,N_14121);
and UO_949 (O_949,N_14084,N_12161);
nor UO_950 (O_950,N_12330,N_13721);
xnor UO_951 (O_951,N_13276,N_12107);
nand UO_952 (O_952,N_12487,N_13904);
or UO_953 (O_953,N_14808,N_13373);
and UO_954 (O_954,N_13121,N_12255);
or UO_955 (O_955,N_13795,N_12026);
nor UO_956 (O_956,N_13177,N_12348);
or UO_957 (O_957,N_14869,N_13205);
and UO_958 (O_958,N_12358,N_14468);
nand UO_959 (O_959,N_14667,N_14757);
nand UO_960 (O_960,N_12589,N_12278);
or UO_961 (O_961,N_14727,N_14375);
nand UO_962 (O_962,N_14515,N_13542);
nor UO_963 (O_963,N_12414,N_14275);
or UO_964 (O_964,N_13106,N_12516);
nand UO_965 (O_965,N_13044,N_12099);
xnor UO_966 (O_966,N_14142,N_14933);
nand UO_967 (O_967,N_12501,N_12022);
or UO_968 (O_968,N_14815,N_12681);
xor UO_969 (O_969,N_13187,N_13922);
nand UO_970 (O_970,N_12575,N_14009);
and UO_971 (O_971,N_12067,N_12028);
xnor UO_972 (O_972,N_14633,N_13839);
nand UO_973 (O_973,N_12944,N_13158);
xnor UO_974 (O_974,N_12647,N_13594);
nand UO_975 (O_975,N_12725,N_14482);
or UO_976 (O_976,N_14377,N_12864);
nand UO_977 (O_977,N_13339,N_14412);
or UO_978 (O_978,N_14028,N_14824);
nand UO_979 (O_979,N_12005,N_13286);
nor UO_980 (O_980,N_14653,N_13609);
nand UO_981 (O_981,N_13988,N_13717);
and UO_982 (O_982,N_13816,N_13751);
nand UO_983 (O_983,N_13288,N_13167);
nor UO_984 (O_984,N_14085,N_13443);
nor UO_985 (O_985,N_13264,N_13860);
xnor UO_986 (O_986,N_13732,N_12311);
nor UO_987 (O_987,N_12648,N_14141);
or UO_988 (O_988,N_14751,N_14128);
nor UO_989 (O_989,N_14300,N_13493);
or UO_990 (O_990,N_12539,N_12894);
nand UO_991 (O_991,N_14523,N_12766);
and UO_992 (O_992,N_14896,N_13740);
nor UO_993 (O_993,N_12360,N_12187);
or UO_994 (O_994,N_12179,N_14177);
or UO_995 (O_995,N_14436,N_12349);
or UO_996 (O_996,N_12165,N_13392);
nand UO_997 (O_997,N_12068,N_12963);
or UO_998 (O_998,N_14429,N_12592);
nor UO_999 (O_999,N_14970,N_13066);
nor UO_1000 (O_1000,N_12714,N_14331);
and UO_1001 (O_1001,N_12302,N_12497);
nor UO_1002 (O_1002,N_13890,N_14221);
and UO_1003 (O_1003,N_13499,N_13562);
nor UO_1004 (O_1004,N_13576,N_14665);
and UO_1005 (O_1005,N_12964,N_14899);
xnor UO_1006 (O_1006,N_13257,N_14378);
and UO_1007 (O_1007,N_12220,N_12836);
or UO_1008 (O_1008,N_14358,N_13113);
and UO_1009 (O_1009,N_12923,N_12023);
and UO_1010 (O_1010,N_12490,N_12483);
nand UO_1011 (O_1011,N_12011,N_14330);
nor UO_1012 (O_1012,N_12411,N_13911);
nand UO_1013 (O_1013,N_12613,N_12893);
nor UO_1014 (O_1014,N_13631,N_14051);
nand UO_1015 (O_1015,N_14565,N_13825);
nand UO_1016 (O_1016,N_12746,N_14823);
nand UO_1017 (O_1017,N_13389,N_13579);
nand UO_1018 (O_1018,N_13699,N_13785);
nor UO_1019 (O_1019,N_13087,N_13636);
xnor UO_1020 (O_1020,N_14856,N_12362);
nor UO_1021 (O_1021,N_14997,N_14807);
nor UO_1022 (O_1022,N_13099,N_12973);
nand UO_1023 (O_1023,N_13645,N_13414);
and UO_1024 (O_1024,N_12419,N_12805);
nand UO_1025 (O_1025,N_13383,N_13381);
nand UO_1026 (O_1026,N_12247,N_13254);
nand UO_1027 (O_1027,N_14612,N_13445);
nor UO_1028 (O_1028,N_13132,N_14680);
nand UO_1029 (O_1029,N_13849,N_12750);
nor UO_1030 (O_1030,N_14733,N_14678);
and UO_1031 (O_1031,N_13710,N_12144);
nand UO_1032 (O_1032,N_12840,N_13577);
nand UO_1033 (O_1033,N_12438,N_14704);
nand UO_1034 (O_1034,N_12598,N_14783);
nor UO_1035 (O_1035,N_13870,N_13032);
or UO_1036 (O_1036,N_12911,N_13796);
xnor UO_1037 (O_1037,N_14276,N_14077);
nand UO_1038 (O_1038,N_14293,N_14884);
nor UO_1039 (O_1039,N_14045,N_12241);
or UO_1040 (O_1040,N_13794,N_12999);
xor UO_1041 (O_1041,N_13998,N_12120);
or UO_1042 (O_1042,N_12201,N_14466);
nand UO_1043 (O_1043,N_12860,N_12775);
nor UO_1044 (O_1044,N_13981,N_13587);
xnor UO_1045 (O_1045,N_13318,N_14942);
xnor UO_1046 (O_1046,N_14663,N_13819);
or UO_1047 (O_1047,N_14605,N_12926);
and UO_1048 (O_1048,N_12537,N_12009);
nand UO_1049 (O_1049,N_12481,N_14202);
and UO_1050 (O_1050,N_13900,N_12167);
and UO_1051 (O_1051,N_13063,N_14393);
nand UO_1052 (O_1052,N_12704,N_14762);
nor UO_1053 (O_1053,N_14759,N_12434);
and UO_1054 (O_1054,N_12158,N_12885);
nor UO_1055 (O_1055,N_12814,N_12454);
and UO_1056 (O_1056,N_12460,N_12322);
nor UO_1057 (O_1057,N_14376,N_13983);
nand UO_1058 (O_1058,N_13155,N_12269);
nor UO_1059 (O_1059,N_14833,N_14180);
and UO_1060 (O_1060,N_14632,N_12418);
and UO_1061 (O_1061,N_12137,N_14518);
nand UO_1062 (O_1062,N_13742,N_12273);
nor UO_1063 (O_1063,N_12983,N_14901);
or UO_1064 (O_1064,N_13317,N_13654);
nand UO_1065 (O_1065,N_13944,N_14179);
and UO_1066 (O_1066,N_14131,N_12755);
nor UO_1067 (O_1067,N_13281,N_12132);
and UO_1068 (O_1068,N_14558,N_13340);
or UO_1069 (O_1069,N_14421,N_14146);
xor UO_1070 (O_1070,N_13876,N_13133);
and UO_1071 (O_1071,N_12587,N_14955);
and UO_1072 (O_1072,N_13955,N_12371);
nor UO_1073 (O_1073,N_14448,N_12720);
nand UO_1074 (O_1074,N_13838,N_13846);
and UO_1075 (O_1075,N_13817,N_14124);
nand UO_1076 (O_1076,N_13821,N_13658);
and UO_1077 (O_1077,N_14130,N_13072);
and UO_1078 (O_1078,N_13907,N_13531);
or UO_1079 (O_1079,N_12052,N_13782);
and UO_1080 (O_1080,N_13386,N_12979);
or UO_1081 (O_1081,N_14138,N_14104);
nor UO_1082 (O_1082,N_13929,N_14487);
nand UO_1083 (O_1083,N_13585,N_14543);
or UO_1084 (O_1084,N_12290,N_12288);
or UO_1085 (O_1085,N_14528,N_12793);
and UO_1086 (O_1086,N_12002,N_14781);
or UO_1087 (O_1087,N_12813,N_14629);
nor UO_1088 (O_1088,N_13942,N_14880);
nor UO_1089 (O_1089,N_12039,N_13679);
nor UO_1090 (O_1090,N_14618,N_14237);
nor UO_1091 (O_1091,N_13522,N_12865);
xor UO_1092 (O_1092,N_14845,N_14741);
nand UO_1093 (O_1093,N_12055,N_14491);
nor UO_1094 (O_1094,N_13887,N_13897);
and UO_1095 (O_1095,N_14968,N_13628);
and UO_1096 (O_1096,N_13076,N_13342);
nor UO_1097 (O_1097,N_13514,N_14260);
and UO_1098 (O_1098,N_13430,N_13638);
nand UO_1099 (O_1099,N_12823,N_13668);
nand UO_1100 (O_1100,N_12980,N_12787);
or UO_1101 (O_1101,N_12507,N_14262);
nor UO_1102 (O_1102,N_13503,N_14411);
or UO_1103 (O_1103,N_12968,N_12958);
nor UO_1104 (O_1104,N_12131,N_14452);
and UO_1105 (O_1105,N_13502,N_12114);
nor UO_1106 (O_1106,N_13232,N_12431);
or UO_1107 (O_1107,N_13755,N_13344);
and UO_1108 (O_1108,N_12195,N_13568);
nor UO_1109 (O_1109,N_12061,N_13001);
nand UO_1110 (O_1110,N_13966,N_14174);
nor UO_1111 (O_1111,N_13972,N_13718);
and UO_1112 (O_1112,N_13744,N_13095);
nor UO_1113 (O_1113,N_13572,N_12245);
and UO_1114 (O_1114,N_14492,N_13559);
and UO_1115 (O_1115,N_14219,N_13551);
xor UO_1116 (O_1116,N_13520,N_13271);
or UO_1117 (O_1117,N_12032,N_12538);
nand UO_1118 (O_1118,N_14541,N_12096);
and UO_1119 (O_1119,N_14613,N_14597);
or UO_1120 (O_1120,N_12451,N_12415);
nor UO_1121 (O_1121,N_12313,N_14788);
and UO_1122 (O_1122,N_12664,N_13465);
nor UO_1123 (O_1123,N_12939,N_14444);
xnor UO_1124 (O_1124,N_13446,N_12385);
nand UO_1125 (O_1125,N_12849,N_14551);
and UO_1126 (O_1126,N_13255,N_12898);
and UO_1127 (O_1127,N_13330,N_14530);
and UO_1128 (O_1128,N_14176,N_12961);
nor UO_1129 (O_1129,N_13537,N_12226);
nand UO_1130 (O_1130,N_14158,N_13595);
and UO_1131 (O_1131,N_12031,N_13902);
or UO_1132 (O_1132,N_12753,N_13886);
or UO_1133 (O_1133,N_13292,N_12900);
nand UO_1134 (O_1134,N_14569,N_13199);
nand UO_1135 (O_1135,N_14664,N_12370);
nor UO_1136 (O_1136,N_14470,N_14616);
and UO_1137 (O_1137,N_14211,N_13141);
nand UO_1138 (O_1138,N_13818,N_12404);
and UO_1139 (O_1139,N_12610,N_13384);
or UO_1140 (O_1140,N_13353,N_12216);
nand UO_1141 (O_1141,N_12697,N_12834);
nand UO_1142 (O_1142,N_12763,N_13082);
nand UO_1143 (O_1143,N_12098,N_14269);
nor UO_1144 (O_1144,N_13500,N_12808);
and UO_1145 (O_1145,N_12859,N_14636);
or UO_1146 (O_1146,N_14576,N_13126);
or UO_1147 (O_1147,N_14217,N_13753);
nor UO_1148 (O_1148,N_14449,N_12692);
or UO_1149 (O_1149,N_12169,N_12723);
xnor UO_1150 (O_1150,N_14212,N_14700);
or UO_1151 (O_1151,N_14511,N_14428);
nand UO_1152 (O_1152,N_14638,N_13772);
nand UO_1153 (O_1153,N_12286,N_13974);
and UO_1154 (O_1154,N_14242,N_13523);
or UO_1155 (O_1155,N_13688,N_14542);
nor UO_1156 (O_1156,N_14220,N_13085);
xnor UO_1157 (O_1157,N_14073,N_13877);
nor UO_1158 (O_1158,N_12975,N_13778);
or UO_1159 (O_1159,N_12469,N_13145);
or UO_1160 (O_1160,N_14029,N_13210);
xor UO_1161 (O_1161,N_14160,N_12913);
nand UO_1162 (O_1162,N_13454,N_14767);
nand UO_1163 (O_1163,N_12428,N_12318);
or UO_1164 (O_1164,N_13600,N_12724);
and UO_1165 (O_1165,N_12998,N_13621);
nor UO_1166 (O_1166,N_14791,N_12937);
nor UO_1167 (O_1167,N_12888,N_14047);
nor UO_1168 (O_1168,N_14519,N_12164);
and UO_1169 (O_1169,N_13543,N_14229);
and UO_1170 (O_1170,N_13475,N_14567);
and UO_1171 (O_1171,N_12279,N_13530);
or UO_1172 (O_1172,N_12887,N_14023);
or UO_1173 (O_1173,N_14950,N_12134);
or UO_1174 (O_1174,N_14532,N_14391);
xor UO_1175 (O_1175,N_14538,N_12794);
and UO_1176 (O_1176,N_13741,N_13758);
nand UO_1177 (O_1177,N_14295,N_14580);
and UO_1178 (O_1178,N_12688,N_12997);
nor UO_1179 (O_1179,N_14266,N_12202);
and UO_1180 (O_1180,N_14420,N_13607);
nand UO_1181 (O_1181,N_12261,N_12711);
nand UO_1182 (O_1182,N_13681,N_14797);
or UO_1183 (O_1183,N_14956,N_12707);
and UO_1184 (O_1184,N_12218,N_14724);
nand UO_1185 (O_1185,N_13779,N_12405);
or UO_1186 (O_1186,N_14651,N_13451);
or UO_1187 (O_1187,N_13602,N_12708);
and UO_1188 (O_1188,N_13643,N_13404);
nor UO_1189 (O_1189,N_12918,N_12065);
nor UO_1190 (O_1190,N_12248,N_12365);
and UO_1191 (O_1191,N_14832,N_14963);
nand UO_1192 (O_1192,N_14866,N_12663);
xor UO_1193 (O_1193,N_13920,N_12635);
or UO_1194 (O_1194,N_13305,N_13382);
xnor UO_1195 (O_1195,N_13007,N_13660);
nor UO_1196 (O_1196,N_13055,N_12897);
or UO_1197 (O_1197,N_13913,N_12594);
or UO_1198 (O_1198,N_12960,N_14413);
nor UO_1199 (O_1199,N_13098,N_12204);
and UO_1200 (O_1200,N_14871,N_14685);
and UO_1201 (O_1201,N_12439,N_12503);
xnor UO_1202 (O_1202,N_12160,N_13056);
nand UO_1203 (O_1203,N_13497,N_13912);
nand UO_1204 (O_1204,N_13487,N_14707);
nor UO_1205 (O_1205,N_13640,N_12430);
nand UO_1206 (O_1206,N_12262,N_12461);
and UO_1207 (O_1207,N_12341,N_12530);
or UO_1208 (O_1208,N_14882,N_12363);
and UO_1209 (O_1209,N_13483,N_14250);
xor UO_1210 (O_1210,N_12661,N_12883);
or UO_1211 (O_1211,N_14925,N_12956);
and UO_1212 (O_1212,N_12445,N_12063);
or UO_1213 (O_1213,N_12339,N_13987);
nand UO_1214 (O_1214,N_13824,N_13468);
and UO_1215 (O_1215,N_12364,N_13296);
and UO_1216 (O_1216,N_12555,N_12596);
nand UO_1217 (O_1217,N_14905,N_14344);
nand UO_1218 (O_1218,N_14827,N_13766);
nand UO_1219 (O_1219,N_13919,N_12188);
nor UO_1220 (O_1220,N_14917,N_14309);
nand UO_1221 (O_1221,N_14101,N_12331);
and UO_1222 (O_1222,N_13774,N_12778);
and UO_1223 (O_1223,N_12149,N_14581);
or UO_1224 (O_1224,N_14798,N_13869);
nand UO_1225 (O_1225,N_12993,N_12821);
nand UO_1226 (O_1226,N_13212,N_14786);
nand UO_1227 (O_1227,N_14076,N_13780);
and UO_1228 (O_1228,N_12437,N_13356);
and UO_1229 (O_1229,N_14599,N_13677);
or UO_1230 (O_1230,N_13561,N_12074);
nand UO_1231 (O_1231,N_14554,N_14693);
and UO_1232 (O_1232,N_12038,N_13997);
xor UO_1233 (O_1233,N_14652,N_12342);
nand UO_1234 (O_1234,N_12051,N_14918);
and UO_1235 (O_1235,N_13488,N_12553);
or UO_1236 (O_1236,N_12416,N_14934);
or UO_1237 (O_1237,N_12933,N_13733);
nand UO_1238 (O_1238,N_12622,N_13637);
xor UO_1239 (O_1239,N_14931,N_13043);
or UO_1240 (O_1240,N_13611,N_14451);
or UO_1241 (O_1241,N_13648,N_13371);
or UO_1242 (O_1242,N_13396,N_14240);
and UO_1243 (O_1243,N_13139,N_12276);
nand UO_1244 (O_1244,N_13545,N_13096);
xor UO_1245 (O_1245,N_14230,N_12566);
and UO_1246 (O_1246,N_12745,N_12049);
nor UO_1247 (O_1247,N_14405,N_14982);
or UO_1248 (O_1248,N_14661,N_12617);
nand UO_1249 (O_1249,N_12630,N_13206);
nor UO_1250 (O_1250,N_14410,N_12784);
nand UO_1251 (O_1251,N_14517,N_13996);
or UO_1252 (O_1252,N_14312,N_12502);
or UO_1253 (O_1253,N_13761,N_14938);
and UO_1254 (O_1254,N_13973,N_13799);
and UO_1255 (O_1255,N_14662,N_13605);
nand UO_1256 (O_1256,N_13724,N_12930);
and UO_1257 (O_1257,N_12608,N_14742);
nor UO_1258 (O_1258,N_13315,N_14805);
nand UO_1259 (O_1259,N_12336,N_14789);
or UO_1260 (O_1260,N_12590,N_12185);
or UO_1261 (O_1261,N_12643,N_13246);
or UO_1262 (O_1262,N_12110,N_12922);
xor UO_1263 (O_1263,N_12771,N_12242);
and UO_1264 (O_1264,N_12915,N_14093);
nand UO_1265 (O_1265,N_12210,N_14501);
nor UO_1266 (O_1266,N_14234,N_12221);
and UO_1267 (O_1267,N_13312,N_13466);
and UO_1268 (O_1268,N_14200,N_13237);
and UO_1269 (O_1269,N_12333,N_12109);
and UO_1270 (O_1270,N_13968,N_14055);
or UO_1271 (O_1271,N_13110,N_13863);
and UO_1272 (O_1272,N_14381,N_14248);
nor UO_1273 (O_1273,N_12621,N_13261);
nor UO_1274 (O_1274,N_12791,N_12151);
nand UO_1275 (O_1275,N_13930,N_14946);
nor UO_1276 (O_1276,N_12799,N_13792);
nand UO_1277 (O_1277,N_14577,N_12659);
or UO_1278 (O_1278,N_14346,N_12250);
nand UO_1279 (O_1279,N_14106,N_14728);
or UO_1280 (O_1280,N_13175,N_13673);
nand UO_1281 (O_1281,N_14606,N_13230);
and UO_1282 (O_1282,N_14583,N_14921);
or UO_1283 (O_1283,N_12156,N_13385);
nand UO_1284 (O_1284,N_14401,N_13209);
or UO_1285 (O_1285,N_14261,N_12558);
and UO_1286 (O_1286,N_14572,N_12941);
nor UO_1287 (O_1287,N_14233,N_14672);
or UO_1288 (O_1288,N_12101,N_12234);
nor UO_1289 (O_1289,N_12580,N_12104);
or UO_1290 (O_1290,N_12083,N_14835);
nor UO_1291 (O_1291,N_12825,N_13915);
nand UO_1292 (O_1292,N_14340,N_12882);
and UO_1293 (O_1293,N_13105,N_13407);
or UO_1294 (O_1294,N_14948,N_12123);
or UO_1295 (O_1295,N_13954,N_13431);
and UO_1296 (O_1296,N_13708,N_12312);
nand UO_1297 (O_1297,N_12315,N_14716);
or UO_1298 (O_1298,N_12612,N_14908);
or UO_1299 (O_1299,N_13322,N_12760);
or UO_1300 (O_1300,N_12738,N_14243);
nand UO_1301 (O_1301,N_14777,N_14013);
or UO_1302 (O_1302,N_13659,N_14247);
or UO_1303 (O_1303,N_13338,N_13010);
and UO_1304 (O_1304,N_13038,N_13480);
xnor UO_1305 (O_1305,N_13856,N_12072);
or UO_1306 (O_1306,N_14112,N_12304);
or UO_1307 (O_1307,N_12367,N_12190);
and UO_1308 (O_1308,N_13507,N_13127);
or UO_1309 (O_1309,N_14271,N_12972);
xor UO_1310 (O_1310,N_14379,N_13787);
nand UO_1311 (O_1311,N_13989,N_14879);
nand UO_1312 (O_1312,N_13694,N_14321);
or UO_1313 (O_1313,N_14784,N_12228);
xnor UO_1314 (O_1314,N_12769,N_14980);
nor UO_1315 (O_1315,N_12048,N_12872);
and UO_1316 (O_1316,N_13184,N_13027);
nand UO_1317 (O_1317,N_12743,N_14843);
nand UO_1318 (O_1318,N_12996,N_12695);
or UO_1319 (O_1319,N_12767,N_12870);
or UO_1320 (O_1320,N_12595,N_13630);
and UO_1321 (O_1321,N_12379,N_14604);
or UO_1322 (O_1322,N_14497,N_12433);
nor UO_1323 (O_1323,N_13820,N_13173);
or UO_1324 (O_1324,N_13136,N_13712);
nand UO_1325 (O_1325,N_12943,N_14561);
nor UO_1326 (O_1326,N_12154,N_13275);
nand UO_1327 (O_1327,N_14658,N_13492);
nand UO_1328 (O_1328,N_12602,N_12666);
or UO_1329 (O_1329,N_14450,N_12842);
or UO_1330 (O_1330,N_13231,N_12227);
nor UO_1331 (O_1331,N_13142,N_14004);
or UO_1332 (O_1332,N_13294,N_13360);
nand UO_1333 (O_1333,N_14036,N_12206);
nand UO_1334 (O_1334,N_14214,N_14826);
and UO_1335 (O_1335,N_13395,N_12987);
nor UO_1336 (O_1336,N_12139,N_12636);
or UO_1337 (O_1337,N_12844,N_12129);
nand UO_1338 (O_1338,N_13436,N_12041);
and UO_1339 (O_1339,N_13603,N_14034);
or UO_1340 (O_1340,N_12586,N_14715);
and UO_1341 (O_1341,N_13883,N_13375);
and UO_1342 (O_1342,N_13701,N_14060);
and UO_1343 (O_1343,N_13943,N_12892);
xor UO_1344 (O_1344,N_14944,N_12335);
nand UO_1345 (O_1345,N_12116,N_14555);
nor UO_1346 (O_1346,N_12478,N_13689);
nor UO_1347 (O_1347,N_12599,N_13873);
xor UO_1348 (O_1348,N_14870,N_13888);
nor UO_1349 (O_1349,N_13841,N_12326);
or UO_1350 (O_1350,N_12464,N_14906);
nand UO_1351 (O_1351,N_13450,N_13923);
or UO_1352 (O_1352,N_12556,N_13080);
and UO_1353 (O_1353,N_13624,N_13166);
xnor UO_1354 (O_1354,N_14764,N_14990);
nand UO_1355 (O_1355,N_14406,N_12097);
nor UO_1356 (O_1356,N_14640,N_12054);
nand UO_1357 (O_1357,N_14279,N_12632);
xor UO_1358 (O_1358,N_13069,N_12754);
nand UO_1359 (O_1359,N_12574,N_14361);
nor UO_1360 (O_1360,N_12625,N_14888);
nand UO_1361 (O_1361,N_12473,N_12917);
nor UO_1362 (O_1362,N_13011,N_14562);
nor UO_1363 (O_1363,N_12181,N_12669);
nand UO_1364 (O_1364,N_13300,N_14999);
nand UO_1365 (O_1365,N_13554,N_12792);
nor UO_1366 (O_1366,N_12498,N_14342);
nor UO_1367 (O_1367,N_12650,N_14416);
or UO_1368 (O_1368,N_14203,N_13314);
xor UO_1369 (O_1369,N_14139,N_13754);
nor UO_1370 (O_1370,N_12446,N_12232);
and UO_1371 (O_1371,N_14172,N_13321);
nor UO_1372 (O_1372,N_13615,N_12730);
nor UO_1373 (O_1373,N_12884,N_13738);
or UO_1374 (O_1374,N_12781,N_12682);
or UO_1375 (O_1375,N_13438,N_14218);
nand UO_1376 (O_1376,N_12670,N_12400);
nor UO_1377 (O_1377,N_14041,N_13547);
or UO_1378 (O_1378,N_13723,N_14537);
or UO_1379 (O_1379,N_14514,N_14502);
nor UO_1380 (O_1380,N_13222,N_13971);
nand UO_1381 (O_1381,N_12252,N_14324);
nand UO_1382 (O_1382,N_13769,N_13512);
nor UO_1383 (O_1383,N_12827,N_12936);
or UO_1384 (O_1384,N_14226,N_14315);
nand UO_1385 (O_1385,N_14438,N_14162);
nor UO_1386 (O_1386,N_13200,N_13447);
nand UO_1387 (O_1387,N_12579,N_14307);
and UO_1388 (O_1388,N_14645,N_13892);
or UO_1389 (O_1389,N_14620,N_12572);
nand UO_1390 (O_1390,N_14725,N_13128);
nand UO_1391 (O_1391,N_13442,N_12812);
or UO_1392 (O_1392,N_12935,N_12841);
and UO_1393 (O_1393,N_13137,N_12203);
xnor UO_1394 (O_1394,N_14454,N_12824);
nand UO_1395 (O_1395,N_12122,N_13549);
xnor UO_1396 (O_1396,N_12703,N_14224);
nor UO_1397 (O_1397,N_13853,N_12012);
xnor UO_1398 (O_1398,N_12309,N_12423);
or UO_1399 (O_1399,N_13023,N_12719);
and UO_1400 (O_1400,N_12407,N_14000);
nand UO_1401 (O_1401,N_14431,N_13926);
nor UO_1402 (O_1402,N_14437,N_13667);
and UO_1403 (O_1403,N_12153,N_13647);
nand UO_1404 (O_1404,N_12301,N_12826);
nor UO_1405 (O_1405,N_12653,N_14974);
nand UO_1406 (O_1406,N_14336,N_13017);
and UO_1407 (O_1407,N_12444,N_13016);
or UO_1408 (O_1408,N_14873,N_13048);
nand UO_1409 (O_1409,N_13491,N_14953);
or UO_1410 (O_1410,N_13845,N_13185);
nor UO_1411 (O_1411,N_12450,N_14684);
and UO_1412 (O_1412,N_13428,N_13567);
and UO_1413 (O_1413,N_13784,N_13591);
and UO_1414 (O_1414,N_13449,N_13836);
or UO_1415 (O_1415,N_13052,N_12955);
and UO_1416 (O_1416,N_14471,N_14117);
nand UO_1417 (O_1417,N_12795,N_13252);
nand UO_1418 (O_1418,N_12343,N_12910);
and UO_1419 (O_1419,N_14027,N_12604);
or UO_1420 (O_1420,N_12403,N_14319);
nor UO_1421 (O_1421,N_14668,N_13614);
and UO_1422 (O_1422,N_14425,N_14460);
xnor UO_1423 (O_1423,N_12817,N_14840);
or UO_1424 (O_1424,N_12040,N_14255);
xnor UO_1425 (O_1425,N_12667,N_13965);
and UO_1426 (O_1426,N_14496,N_14881);
and UO_1427 (O_1427,N_14998,N_14109);
nand UO_1428 (O_1428,N_14928,N_13803);
and UO_1429 (O_1429,N_12905,N_13463);
nand UO_1430 (O_1430,N_14064,N_13884);
and UO_1431 (O_1431,N_13553,N_12174);
nor UO_1432 (O_1432,N_14600,N_13945);
nand UO_1433 (O_1433,N_13768,N_13885);
or UO_1434 (O_1434,N_13036,N_13274);
nor UO_1435 (O_1435,N_13566,N_12388);
or UO_1436 (O_1436,N_12749,N_13678);
or UO_1437 (O_1437,N_14967,N_12223);
and UO_1438 (O_1438,N_12992,N_12839);
nor UO_1439 (O_1439,N_12728,N_12856);
nor UO_1440 (O_1440,N_13533,N_13823);
nand UO_1441 (O_1441,N_14627,N_13019);
nand UO_1442 (O_1442,N_13881,N_14969);
nor UO_1443 (O_1443,N_12970,N_12353);
nor UO_1444 (O_1444,N_14052,N_12465);
or UO_1445 (O_1445,N_13646,N_13563);
and UO_1446 (O_1446,N_12283,N_14559);
and UO_1447 (O_1447,N_13875,N_12951);
or UO_1448 (O_1448,N_14932,N_12058);
and UO_1449 (O_1449,N_12957,N_14736);
and UO_1450 (O_1450,N_14858,N_13323);
or UO_1451 (O_1451,N_13588,N_13770);
nor UO_1452 (O_1452,N_14197,N_14280);
nand UO_1453 (O_1453,N_12092,N_14349);
xor UO_1454 (O_1454,N_12751,N_12848);
and UO_1455 (O_1455,N_14178,N_13495);
and UO_1456 (O_1456,N_13148,N_12018);
nor UO_1457 (O_1457,N_14422,N_12873);
and UO_1458 (O_1458,N_12060,N_12162);
xnor UO_1459 (O_1459,N_13309,N_13686);
or UO_1460 (O_1460,N_13641,N_12292);
or UO_1461 (O_1461,N_14043,N_14643);
nor UO_1462 (O_1462,N_12044,N_13432);
nor UO_1463 (O_1463,N_12268,N_12263);
nor UO_1464 (O_1464,N_13238,N_12492);
nand UO_1465 (O_1465,N_13390,N_13790);
nand UO_1466 (O_1466,N_13045,N_13215);
or UO_1467 (O_1467,N_14001,N_14322);
or UO_1468 (O_1468,N_14486,N_12591);
and UO_1469 (O_1469,N_12694,N_14735);
and UO_1470 (O_1470,N_12739,N_12345);
nor UO_1471 (O_1471,N_13195,N_14657);
nand UO_1472 (O_1472,N_14550,N_12140);
nand UO_1473 (O_1473,N_12550,N_12614);
and UO_1474 (O_1474,N_12173,N_14010);
and UO_1475 (O_1475,N_13355,N_13101);
or UO_1476 (O_1476,N_12752,N_12557);
and UO_1477 (O_1477,N_14546,N_14592);
xnor UO_1478 (O_1478,N_13160,N_12611);
or UO_1479 (O_1479,N_13225,N_12467);
and UO_1480 (O_1480,N_12657,N_13822);
nor UO_1481 (O_1481,N_12474,N_13513);
or UO_1482 (O_1482,N_12209,N_13936);
nor UO_1483 (O_1483,N_13830,N_12081);
nor UO_1484 (O_1484,N_14119,N_12480);
nand UO_1485 (O_1485,N_13273,N_14382);
nor UO_1486 (O_1486,N_12514,N_13084);
and UO_1487 (O_1487,N_14185,N_14417);
nand UO_1488 (O_1488,N_13949,N_13077);
or UO_1489 (O_1489,N_13909,N_13102);
nand UO_1490 (O_1490,N_13788,N_14839);
nor UO_1491 (O_1491,N_14285,N_14673);
and UO_1492 (O_1492,N_14286,N_13341);
xor UO_1493 (O_1493,N_12243,N_14020);
nand UO_1494 (O_1494,N_13669,N_12777);
nand UO_1495 (O_1495,N_13298,N_14749);
and UO_1496 (O_1496,N_12004,N_13411);
or UO_1497 (O_1497,N_12455,N_13050);
or UO_1498 (O_1498,N_14297,N_13864);
nand UO_1499 (O_1499,N_14649,N_13013);
xnor UO_1500 (O_1500,N_14397,N_12420);
and UO_1501 (O_1501,N_14972,N_13541);
nor UO_1502 (O_1502,N_13957,N_14010);
or UO_1503 (O_1503,N_13733,N_12954);
or UO_1504 (O_1504,N_13282,N_13653);
nand UO_1505 (O_1505,N_12161,N_14146);
nor UO_1506 (O_1506,N_12037,N_14995);
nand UO_1507 (O_1507,N_13186,N_12058);
nor UO_1508 (O_1508,N_13816,N_12158);
nand UO_1509 (O_1509,N_13719,N_12415);
nand UO_1510 (O_1510,N_12891,N_12089);
nand UO_1511 (O_1511,N_12705,N_14635);
and UO_1512 (O_1512,N_12396,N_14555);
nor UO_1513 (O_1513,N_14896,N_12492);
xnor UO_1514 (O_1514,N_12607,N_14692);
and UO_1515 (O_1515,N_12957,N_13984);
nand UO_1516 (O_1516,N_13465,N_14987);
and UO_1517 (O_1517,N_12323,N_12451);
nor UO_1518 (O_1518,N_14659,N_14600);
xor UO_1519 (O_1519,N_12675,N_12561);
or UO_1520 (O_1520,N_14403,N_14329);
and UO_1521 (O_1521,N_14370,N_14238);
nor UO_1522 (O_1522,N_13022,N_14940);
or UO_1523 (O_1523,N_14614,N_12890);
nor UO_1524 (O_1524,N_13130,N_12135);
nor UO_1525 (O_1525,N_13274,N_14698);
and UO_1526 (O_1526,N_12137,N_12186);
and UO_1527 (O_1527,N_12965,N_12341);
and UO_1528 (O_1528,N_13340,N_12806);
xnor UO_1529 (O_1529,N_12559,N_14068);
nand UO_1530 (O_1530,N_12358,N_12278);
or UO_1531 (O_1531,N_13030,N_12116);
nor UO_1532 (O_1532,N_12124,N_13332);
and UO_1533 (O_1533,N_12817,N_14727);
and UO_1534 (O_1534,N_13081,N_13864);
nand UO_1535 (O_1535,N_12543,N_12192);
nand UO_1536 (O_1536,N_12741,N_14277);
nand UO_1537 (O_1537,N_14839,N_13147);
or UO_1538 (O_1538,N_14333,N_14890);
nand UO_1539 (O_1539,N_13762,N_12780);
nand UO_1540 (O_1540,N_13283,N_13389);
or UO_1541 (O_1541,N_14803,N_13086);
or UO_1542 (O_1542,N_14067,N_14112);
nand UO_1543 (O_1543,N_12957,N_14719);
nor UO_1544 (O_1544,N_13612,N_14485);
xor UO_1545 (O_1545,N_12112,N_14253);
and UO_1546 (O_1546,N_14987,N_12339);
or UO_1547 (O_1547,N_14039,N_13644);
nand UO_1548 (O_1548,N_14400,N_13483);
and UO_1549 (O_1549,N_14738,N_12490);
nor UO_1550 (O_1550,N_13164,N_14927);
nor UO_1551 (O_1551,N_12246,N_12199);
and UO_1552 (O_1552,N_13629,N_12988);
nand UO_1553 (O_1553,N_14418,N_13515);
and UO_1554 (O_1554,N_14445,N_14754);
and UO_1555 (O_1555,N_13438,N_13505);
xnor UO_1556 (O_1556,N_14207,N_14820);
xnor UO_1557 (O_1557,N_13868,N_13941);
and UO_1558 (O_1558,N_14983,N_12329);
nand UO_1559 (O_1559,N_14653,N_13680);
xnor UO_1560 (O_1560,N_13213,N_13063);
nor UO_1561 (O_1561,N_13315,N_13626);
nor UO_1562 (O_1562,N_13448,N_12517);
and UO_1563 (O_1563,N_12083,N_14675);
xor UO_1564 (O_1564,N_12248,N_14747);
xnor UO_1565 (O_1565,N_14241,N_12782);
nand UO_1566 (O_1566,N_14130,N_14564);
nor UO_1567 (O_1567,N_14243,N_12422);
nor UO_1568 (O_1568,N_14988,N_12333);
and UO_1569 (O_1569,N_13984,N_14744);
or UO_1570 (O_1570,N_13889,N_14174);
xnor UO_1571 (O_1571,N_13359,N_12879);
nor UO_1572 (O_1572,N_12313,N_13268);
nand UO_1573 (O_1573,N_12309,N_13443);
nor UO_1574 (O_1574,N_14324,N_12606);
nor UO_1575 (O_1575,N_14901,N_13141);
nand UO_1576 (O_1576,N_14692,N_14155);
or UO_1577 (O_1577,N_13191,N_14108);
nand UO_1578 (O_1578,N_13186,N_12137);
nor UO_1579 (O_1579,N_13215,N_12636);
or UO_1580 (O_1580,N_14833,N_13080);
nand UO_1581 (O_1581,N_13105,N_13575);
and UO_1582 (O_1582,N_13623,N_14804);
or UO_1583 (O_1583,N_13149,N_12091);
nand UO_1584 (O_1584,N_13484,N_14339);
or UO_1585 (O_1585,N_12121,N_14240);
or UO_1586 (O_1586,N_13229,N_12710);
nor UO_1587 (O_1587,N_13654,N_13599);
and UO_1588 (O_1588,N_13740,N_14400);
or UO_1589 (O_1589,N_12931,N_12066);
nand UO_1590 (O_1590,N_12277,N_13615);
nand UO_1591 (O_1591,N_12601,N_13502);
nand UO_1592 (O_1592,N_12277,N_14269);
nand UO_1593 (O_1593,N_14329,N_12907);
or UO_1594 (O_1594,N_14969,N_14165);
and UO_1595 (O_1595,N_12709,N_14303);
nand UO_1596 (O_1596,N_14088,N_14153);
nand UO_1597 (O_1597,N_12257,N_13398);
xor UO_1598 (O_1598,N_12101,N_14869);
or UO_1599 (O_1599,N_13102,N_14586);
nor UO_1600 (O_1600,N_12276,N_12511);
nand UO_1601 (O_1601,N_13792,N_14428);
nand UO_1602 (O_1602,N_14448,N_14131);
xnor UO_1603 (O_1603,N_14970,N_12014);
nor UO_1604 (O_1604,N_13061,N_13281);
xnor UO_1605 (O_1605,N_12050,N_12745);
and UO_1606 (O_1606,N_14386,N_12785);
or UO_1607 (O_1607,N_14553,N_14128);
nor UO_1608 (O_1608,N_13880,N_12807);
and UO_1609 (O_1609,N_12603,N_13961);
and UO_1610 (O_1610,N_14998,N_13448);
xnor UO_1611 (O_1611,N_14012,N_13700);
nor UO_1612 (O_1612,N_14510,N_13011);
nor UO_1613 (O_1613,N_13641,N_12721);
or UO_1614 (O_1614,N_13223,N_13770);
or UO_1615 (O_1615,N_13206,N_14342);
xor UO_1616 (O_1616,N_12998,N_12677);
and UO_1617 (O_1617,N_13581,N_12209);
or UO_1618 (O_1618,N_13028,N_12573);
nand UO_1619 (O_1619,N_14278,N_12279);
nor UO_1620 (O_1620,N_12691,N_14300);
nand UO_1621 (O_1621,N_14334,N_12805);
or UO_1622 (O_1622,N_12832,N_13117);
nor UO_1623 (O_1623,N_13712,N_14594);
or UO_1624 (O_1624,N_13951,N_14906);
nand UO_1625 (O_1625,N_12295,N_14379);
nand UO_1626 (O_1626,N_14607,N_14352);
nor UO_1627 (O_1627,N_13279,N_12082);
nor UO_1628 (O_1628,N_14907,N_14350);
or UO_1629 (O_1629,N_14615,N_14609);
nor UO_1630 (O_1630,N_14312,N_12629);
and UO_1631 (O_1631,N_13716,N_13941);
or UO_1632 (O_1632,N_14797,N_13694);
or UO_1633 (O_1633,N_12114,N_12519);
and UO_1634 (O_1634,N_13637,N_14242);
nand UO_1635 (O_1635,N_12829,N_14300);
or UO_1636 (O_1636,N_13661,N_12133);
or UO_1637 (O_1637,N_13641,N_12559);
or UO_1638 (O_1638,N_12720,N_13416);
and UO_1639 (O_1639,N_12482,N_12544);
nor UO_1640 (O_1640,N_14873,N_14827);
and UO_1641 (O_1641,N_14895,N_12569);
and UO_1642 (O_1642,N_13651,N_14360);
or UO_1643 (O_1643,N_13232,N_14112);
nand UO_1644 (O_1644,N_12250,N_12995);
or UO_1645 (O_1645,N_13257,N_13308);
or UO_1646 (O_1646,N_13133,N_12099);
or UO_1647 (O_1647,N_12381,N_12053);
nand UO_1648 (O_1648,N_12521,N_12593);
nor UO_1649 (O_1649,N_14571,N_14782);
nor UO_1650 (O_1650,N_13531,N_12978);
nor UO_1651 (O_1651,N_13688,N_12256);
and UO_1652 (O_1652,N_14423,N_12396);
nor UO_1653 (O_1653,N_14871,N_12160);
nor UO_1654 (O_1654,N_12927,N_12509);
and UO_1655 (O_1655,N_13184,N_14247);
nand UO_1656 (O_1656,N_12823,N_13495);
and UO_1657 (O_1657,N_12453,N_14224);
and UO_1658 (O_1658,N_12331,N_14452);
or UO_1659 (O_1659,N_12299,N_14361);
nand UO_1660 (O_1660,N_14054,N_12313);
nor UO_1661 (O_1661,N_13947,N_14795);
nor UO_1662 (O_1662,N_12642,N_12553);
and UO_1663 (O_1663,N_13121,N_12072);
or UO_1664 (O_1664,N_13078,N_14090);
nor UO_1665 (O_1665,N_14292,N_13594);
or UO_1666 (O_1666,N_13674,N_12809);
or UO_1667 (O_1667,N_13877,N_12454);
nand UO_1668 (O_1668,N_13888,N_14745);
and UO_1669 (O_1669,N_12644,N_13359);
and UO_1670 (O_1670,N_12421,N_13508);
nand UO_1671 (O_1671,N_12291,N_13966);
and UO_1672 (O_1672,N_14428,N_12016);
nand UO_1673 (O_1673,N_12201,N_12555);
and UO_1674 (O_1674,N_12992,N_12329);
or UO_1675 (O_1675,N_13554,N_13736);
nor UO_1676 (O_1676,N_13849,N_12733);
nor UO_1677 (O_1677,N_14833,N_13040);
nor UO_1678 (O_1678,N_14753,N_12663);
and UO_1679 (O_1679,N_13053,N_13680);
nor UO_1680 (O_1680,N_12124,N_13977);
xnor UO_1681 (O_1681,N_13837,N_13880);
nand UO_1682 (O_1682,N_12839,N_14659);
and UO_1683 (O_1683,N_14127,N_13643);
nor UO_1684 (O_1684,N_13371,N_13243);
xor UO_1685 (O_1685,N_14563,N_13455);
nand UO_1686 (O_1686,N_13307,N_14319);
and UO_1687 (O_1687,N_13652,N_14864);
nor UO_1688 (O_1688,N_12456,N_12305);
or UO_1689 (O_1689,N_13814,N_12378);
nor UO_1690 (O_1690,N_13947,N_12585);
nand UO_1691 (O_1691,N_12924,N_12783);
nor UO_1692 (O_1692,N_14430,N_13967);
xor UO_1693 (O_1693,N_13044,N_14456);
xnor UO_1694 (O_1694,N_14449,N_14377);
nor UO_1695 (O_1695,N_12265,N_13411);
nor UO_1696 (O_1696,N_14013,N_12362);
nor UO_1697 (O_1697,N_12386,N_12200);
or UO_1698 (O_1698,N_12365,N_13052);
or UO_1699 (O_1699,N_13983,N_14063);
xnor UO_1700 (O_1700,N_14427,N_14331);
nor UO_1701 (O_1701,N_14625,N_12705);
and UO_1702 (O_1702,N_12814,N_13847);
nand UO_1703 (O_1703,N_14241,N_13949);
nor UO_1704 (O_1704,N_13938,N_14376);
nor UO_1705 (O_1705,N_13945,N_13298);
or UO_1706 (O_1706,N_14858,N_14161);
nor UO_1707 (O_1707,N_13443,N_12142);
and UO_1708 (O_1708,N_14090,N_14665);
nor UO_1709 (O_1709,N_13642,N_14777);
or UO_1710 (O_1710,N_14055,N_13628);
nand UO_1711 (O_1711,N_12170,N_14161);
and UO_1712 (O_1712,N_14595,N_14145);
nor UO_1713 (O_1713,N_12313,N_12211);
or UO_1714 (O_1714,N_13020,N_14247);
and UO_1715 (O_1715,N_12841,N_14472);
nand UO_1716 (O_1716,N_12958,N_13248);
nand UO_1717 (O_1717,N_14614,N_12220);
nand UO_1718 (O_1718,N_12725,N_14800);
nand UO_1719 (O_1719,N_14474,N_13075);
nor UO_1720 (O_1720,N_12855,N_14073);
nand UO_1721 (O_1721,N_14853,N_14638);
nand UO_1722 (O_1722,N_13149,N_12039);
xor UO_1723 (O_1723,N_12935,N_13369);
and UO_1724 (O_1724,N_13819,N_12967);
or UO_1725 (O_1725,N_12776,N_13005);
nor UO_1726 (O_1726,N_13742,N_13015);
nor UO_1727 (O_1727,N_12650,N_13325);
nor UO_1728 (O_1728,N_13875,N_13041);
and UO_1729 (O_1729,N_13743,N_13769);
and UO_1730 (O_1730,N_12294,N_13996);
xor UO_1731 (O_1731,N_12937,N_13932);
or UO_1732 (O_1732,N_14347,N_12309);
nor UO_1733 (O_1733,N_13473,N_13510);
and UO_1734 (O_1734,N_13834,N_14906);
and UO_1735 (O_1735,N_12568,N_12250);
nand UO_1736 (O_1736,N_14909,N_13342);
nand UO_1737 (O_1737,N_14243,N_12615);
nor UO_1738 (O_1738,N_14107,N_13340);
xnor UO_1739 (O_1739,N_12579,N_14739);
nor UO_1740 (O_1740,N_12526,N_12215);
nor UO_1741 (O_1741,N_14886,N_13218);
nand UO_1742 (O_1742,N_12816,N_14205);
nor UO_1743 (O_1743,N_14313,N_13675);
nand UO_1744 (O_1744,N_14003,N_12633);
and UO_1745 (O_1745,N_12310,N_13549);
nand UO_1746 (O_1746,N_13652,N_12707);
nand UO_1747 (O_1747,N_14380,N_14751);
and UO_1748 (O_1748,N_13425,N_12464);
or UO_1749 (O_1749,N_12826,N_14795);
nand UO_1750 (O_1750,N_12211,N_13403);
nand UO_1751 (O_1751,N_14460,N_12368);
nand UO_1752 (O_1752,N_13201,N_13308);
nand UO_1753 (O_1753,N_14433,N_13388);
nand UO_1754 (O_1754,N_12667,N_14476);
or UO_1755 (O_1755,N_14431,N_13457);
and UO_1756 (O_1756,N_12301,N_13064);
nand UO_1757 (O_1757,N_14277,N_14449);
xor UO_1758 (O_1758,N_14680,N_13136);
xor UO_1759 (O_1759,N_14030,N_13544);
nand UO_1760 (O_1760,N_13833,N_12973);
or UO_1761 (O_1761,N_12052,N_13649);
and UO_1762 (O_1762,N_12598,N_13528);
or UO_1763 (O_1763,N_12992,N_13036);
xnor UO_1764 (O_1764,N_14437,N_14042);
nand UO_1765 (O_1765,N_14873,N_12398);
or UO_1766 (O_1766,N_14249,N_12949);
or UO_1767 (O_1767,N_12408,N_14697);
nor UO_1768 (O_1768,N_14606,N_14508);
or UO_1769 (O_1769,N_14352,N_13857);
nand UO_1770 (O_1770,N_14598,N_14664);
nor UO_1771 (O_1771,N_12643,N_13251);
or UO_1772 (O_1772,N_14456,N_13101);
nand UO_1773 (O_1773,N_12279,N_14363);
nand UO_1774 (O_1774,N_14782,N_14346);
or UO_1775 (O_1775,N_12043,N_12457);
xor UO_1776 (O_1776,N_12398,N_14616);
nand UO_1777 (O_1777,N_13971,N_13797);
or UO_1778 (O_1778,N_13958,N_12349);
nor UO_1779 (O_1779,N_12624,N_13035);
or UO_1780 (O_1780,N_13915,N_13254);
xnor UO_1781 (O_1781,N_13912,N_14558);
or UO_1782 (O_1782,N_14899,N_12006);
nand UO_1783 (O_1783,N_14303,N_14667);
and UO_1784 (O_1784,N_13933,N_12320);
nand UO_1785 (O_1785,N_13891,N_12913);
nand UO_1786 (O_1786,N_13615,N_14610);
or UO_1787 (O_1787,N_13311,N_12213);
nand UO_1788 (O_1788,N_13993,N_12065);
or UO_1789 (O_1789,N_13887,N_12059);
nand UO_1790 (O_1790,N_13394,N_14229);
and UO_1791 (O_1791,N_14300,N_14546);
and UO_1792 (O_1792,N_13823,N_12161);
and UO_1793 (O_1793,N_13529,N_14508);
nor UO_1794 (O_1794,N_13375,N_13190);
nor UO_1795 (O_1795,N_12019,N_14173);
nor UO_1796 (O_1796,N_13160,N_13898);
xor UO_1797 (O_1797,N_12467,N_12431);
and UO_1798 (O_1798,N_14170,N_13441);
nand UO_1799 (O_1799,N_14914,N_13005);
xnor UO_1800 (O_1800,N_14069,N_14045);
and UO_1801 (O_1801,N_13733,N_12755);
xor UO_1802 (O_1802,N_13644,N_14009);
and UO_1803 (O_1803,N_13563,N_13377);
or UO_1804 (O_1804,N_12765,N_13234);
nand UO_1805 (O_1805,N_13911,N_13679);
nor UO_1806 (O_1806,N_14312,N_13767);
nor UO_1807 (O_1807,N_14686,N_14723);
and UO_1808 (O_1808,N_12753,N_14319);
and UO_1809 (O_1809,N_14807,N_13005);
nor UO_1810 (O_1810,N_13832,N_14926);
nand UO_1811 (O_1811,N_14845,N_14986);
xnor UO_1812 (O_1812,N_14826,N_13643);
xor UO_1813 (O_1813,N_12689,N_13389);
and UO_1814 (O_1814,N_13834,N_14219);
or UO_1815 (O_1815,N_13840,N_14830);
or UO_1816 (O_1816,N_14159,N_12256);
nor UO_1817 (O_1817,N_13480,N_13746);
or UO_1818 (O_1818,N_12716,N_13235);
nor UO_1819 (O_1819,N_13740,N_13339);
and UO_1820 (O_1820,N_13166,N_12634);
and UO_1821 (O_1821,N_14602,N_12050);
or UO_1822 (O_1822,N_13511,N_13712);
nand UO_1823 (O_1823,N_12701,N_14506);
and UO_1824 (O_1824,N_13321,N_12405);
nand UO_1825 (O_1825,N_14875,N_13089);
and UO_1826 (O_1826,N_14422,N_14767);
or UO_1827 (O_1827,N_14183,N_14539);
nor UO_1828 (O_1828,N_13561,N_12807);
nor UO_1829 (O_1829,N_14815,N_13599);
nor UO_1830 (O_1830,N_14439,N_12505);
and UO_1831 (O_1831,N_13264,N_14177);
or UO_1832 (O_1832,N_13098,N_13861);
nand UO_1833 (O_1833,N_12261,N_12348);
xnor UO_1834 (O_1834,N_14076,N_12250);
nand UO_1835 (O_1835,N_13808,N_13274);
and UO_1836 (O_1836,N_12417,N_12092);
and UO_1837 (O_1837,N_14954,N_12950);
nor UO_1838 (O_1838,N_14203,N_14983);
nand UO_1839 (O_1839,N_14252,N_13383);
nor UO_1840 (O_1840,N_13212,N_14940);
or UO_1841 (O_1841,N_14403,N_12828);
nor UO_1842 (O_1842,N_13632,N_13245);
or UO_1843 (O_1843,N_14150,N_13106);
nor UO_1844 (O_1844,N_12106,N_12282);
nor UO_1845 (O_1845,N_14606,N_13315);
nor UO_1846 (O_1846,N_14982,N_14020);
and UO_1847 (O_1847,N_13210,N_13758);
xor UO_1848 (O_1848,N_13410,N_13382);
or UO_1849 (O_1849,N_12155,N_12003);
xnor UO_1850 (O_1850,N_13435,N_14447);
nand UO_1851 (O_1851,N_13001,N_14751);
xor UO_1852 (O_1852,N_12352,N_13159);
nand UO_1853 (O_1853,N_14829,N_12869);
nor UO_1854 (O_1854,N_14319,N_13883);
nand UO_1855 (O_1855,N_14964,N_13207);
and UO_1856 (O_1856,N_13531,N_13862);
and UO_1857 (O_1857,N_12660,N_14609);
and UO_1858 (O_1858,N_13249,N_14488);
or UO_1859 (O_1859,N_13972,N_12443);
or UO_1860 (O_1860,N_13275,N_13672);
or UO_1861 (O_1861,N_12276,N_13529);
and UO_1862 (O_1862,N_14138,N_13499);
nand UO_1863 (O_1863,N_14474,N_13159);
nand UO_1864 (O_1864,N_14633,N_14128);
nand UO_1865 (O_1865,N_12192,N_12960);
and UO_1866 (O_1866,N_12978,N_13400);
or UO_1867 (O_1867,N_13604,N_13711);
nor UO_1868 (O_1868,N_13589,N_13724);
and UO_1869 (O_1869,N_12557,N_13806);
nor UO_1870 (O_1870,N_14192,N_12999);
nor UO_1871 (O_1871,N_13529,N_14827);
nand UO_1872 (O_1872,N_13404,N_12330);
or UO_1873 (O_1873,N_12313,N_14377);
or UO_1874 (O_1874,N_14531,N_14534);
and UO_1875 (O_1875,N_14848,N_12054);
nor UO_1876 (O_1876,N_14318,N_12120);
and UO_1877 (O_1877,N_12709,N_13902);
or UO_1878 (O_1878,N_13232,N_12631);
nand UO_1879 (O_1879,N_12948,N_13199);
nand UO_1880 (O_1880,N_13173,N_13791);
and UO_1881 (O_1881,N_13354,N_12834);
xor UO_1882 (O_1882,N_12281,N_12857);
nand UO_1883 (O_1883,N_13909,N_13160);
nand UO_1884 (O_1884,N_12509,N_14335);
or UO_1885 (O_1885,N_13716,N_12479);
nand UO_1886 (O_1886,N_14961,N_13242);
nand UO_1887 (O_1887,N_14078,N_14743);
or UO_1888 (O_1888,N_12892,N_14414);
xor UO_1889 (O_1889,N_13831,N_14224);
and UO_1890 (O_1890,N_13472,N_12145);
and UO_1891 (O_1891,N_14411,N_12424);
or UO_1892 (O_1892,N_12716,N_12783);
nor UO_1893 (O_1893,N_13902,N_13256);
nor UO_1894 (O_1894,N_12037,N_12549);
or UO_1895 (O_1895,N_14797,N_14495);
nor UO_1896 (O_1896,N_13035,N_14198);
or UO_1897 (O_1897,N_14845,N_13204);
and UO_1898 (O_1898,N_14063,N_12504);
or UO_1899 (O_1899,N_14370,N_12558);
nand UO_1900 (O_1900,N_12074,N_14070);
or UO_1901 (O_1901,N_14254,N_13738);
and UO_1902 (O_1902,N_12412,N_13051);
or UO_1903 (O_1903,N_12892,N_13439);
nor UO_1904 (O_1904,N_13250,N_12711);
nor UO_1905 (O_1905,N_13268,N_13221);
and UO_1906 (O_1906,N_13211,N_14829);
and UO_1907 (O_1907,N_13879,N_12467);
or UO_1908 (O_1908,N_13024,N_13479);
nor UO_1909 (O_1909,N_13246,N_12651);
xnor UO_1910 (O_1910,N_12087,N_12702);
nor UO_1911 (O_1911,N_14725,N_14221);
or UO_1912 (O_1912,N_13800,N_12918);
nand UO_1913 (O_1913,N_12951,N_14464);
nor UO_1914 (O_1914,N_14517,N_13641);
nand UO_1915 (O_1915,N_13537,N_13064);
or UO_1916 (O_1916,N_13054,N_14765);
or UO_1917 (O_1917,N_13511,N_13430);
nand UO_1918 (O_1918,N_13739,N_13636);
or UO_1919 (O_1919,N_14573,N_13141);
nand UO_1920 (O_1920,N_13343,N_12222);
nand UO_1921 (O_1921,N_14946,N_13722);
xnor UO_1922 (O_1922,N_14582,N_13790);
or UO_1923 (O_1923,N_13156,N_12857);
or UO_1924 (O_1924,N_12803,N_13097);
and UO_1925 (O_1925,N_14722,N_14422);
or UO_1926 (O_1926,N_14443,N_14698);
xor UO_1927 (O_1927,N_12638,N_12702);
nor UO_1928 (O_1928,N_13548,N_12075);
nor UO_1929 (O_1929,N_14195,N_12678);
or UO_1930 (O_1930,N_12132,N_12256);
and UO_1931 (O_1931,N_13669,N_14262);
nor UO_1932 (O_1932,N_14164,N_13415);
and UO_1933 (O_1933,N_12723,N_12102);
nand UO_1934 (O_1934,N_12265,N_12878);
or UO_1935 (O_1935,N_13443,N_12927);
and UO_1936 (O_1936,N_14255,N_14086);
nand UO_1937 (O_1937,N_13661,N_13079);
nor UO_1938 (O_1938,N_14089,N_14295);
nand UO_1939 (O_1939,N_13395,N_12274);
nor UO_1940 (O_1940,N_14580,N_14630);
nand UO_1941 (O_1941,N_14617,N_14291);
and UO_1942 (O_1942,N_12610,N_12682);
xnor UO_1943 (O_1943,N_12983,N_13793);
nand UO_1944 (O_1944,N_12650,N_14774);
or UO_1945 (O_1945,N_13163,N_12368);
or UO_1946 (O_1946,N_12631,N_12063);
nor UO_1947 (O_1947,N_13941,N_14432);
or UO_1948 (O_1948,N_13609,N_13906);
nor UO_1949 (O_1949,N_13255,N_13190);
or UO_1950 (O_1950,N_13674,N_12122);
or UO_1951 (O_1951,N_12726,N_13806);
or UO_1952 (O_1952,N_12339,N_13699);
or UO_1953 (O_1953,N_13402,N_12559);
xnor UO_1954 (O_1954,N_14009,N_12370);
nor UO_1955 (O_1955,N_12128,N_13646);
or UO_1956 (O_1956,N_13540,N_12145);
nor UO_1957 (O_1957,N_14725,N_12632);
or UO_1958 (O_1958,N_12842,N_14194);
xor UO_1959 (O_1959,N_13139,N_13997);
and UO_1960 (O_1960,N_13359,N_12369);
and UO_1961 (O_1961,N_14158,N_14179);
and UO_1962 (O_1962,N_14244,N_12411);
or UO_1963 (O_1963,N_12325,N_14192);
or UO_1964 (O_1964,N_14248,N_12092);
or UO_1965 (O_1965,N_14032,N_14997);
nand UO_1966 (O_1966,N_14513,N_14696);
nor UO_1967 (O_1967,N_14138,N_13527);
nor UO_1968 (O_1968,N_12063,N_13574);
nand UO_1969 (O_1969,N_14190,N_13551);
nand UO_1970 (O_1970,N_13985,N_14288);
nor UO_1971 (O_1971,N_12796,N_14724);
nand UO_1972 (O_1972,N_12105,N_12064);
or UO_1973 (O_1973,N_12820,N_14886);
xnor UO_1974 (O_1974,N_12122,N_13241);
nand UO_1975 (O_1975,N_14102,N_14680);
nor UO_1976 (O_1976,N_13379,N_12880);
nor UO_1977 (O_1977,N_13580,N_14571);
nand UO_1978 (O_1978,N_14661,N_14206);
nand UO_1979 (O_1979,N_14154,N_14648);
or UO_1980 (O_1980,N_13002,N_14920);
and UO_1981 (O_1981,N_12136,N_13762);
or UO_1982 (O_1982,N_13851,N_12020);
and UO_1983 (O_1983,N_14723,N_13768);
nor UO_1984 (O_1984,N_12322,N_12936);
or UO_1985 (O_1985,N_14122,N_14565);
and UO_1986 (O_1986,N_13520,N_14403);
xor UO_1987 (O_1987,N_12360,N_12399);
nand UO_1988 (O_1988,N_14661,N_12940);
xor UO_1989 (O_1989,N_14766,N_12730);
or UO_1990 (O_1990,N_14889,N_14674);
nand UO_1991 (O_1991,N_13409,N_13574);
nor UO_1992 (O_1992,N_12784,N_12026);
xnor UO_1993 (O_1993,N_13400,N_12110);
xnor UO_1994 (O_1994,N_13498,N_14001);
or UO_1995 (O_1995,N_13408,N_13906);
or UO_1996 (O_1996,N_12688,N_12147);
or UO_1997 (O_1997,N_13616,N_14019);
and UO_1998 (O_1998,N_14001,N_12021);
or UO_1999 (O_1999,N_14211,N_12892);
endmodule