module basic_750_5000_1000_10_levels_2xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nor U0 (N_0,In_425,In_336);
and U1 (N_1,In_329,In_614);
nor U2 (N_2,In_471,In_311);
or U3 (N_3,In_536,In_461);
xor U4 (N_4,In_291,In_555);
or U5 (N_5,In_300,In_695);
or U6 (N_6,In_573,In_496);
nor U7 (N_7,In_185,In_120);
or U8 (N_8,In_156,In_126);
and U9 (N_9,In_713,In_286);
nand U10 (N_10,In_320,In_4);
nand U11 (N_11,In_165,In_127);
or U12 (N_12,In_71,In_8);
nand U13 (N_13,In_369,In_107);
or U14 (N_14,In_662,In_648);
and U15 (N_15,In_433,In_638);
or U16 (N_16,In_572,In_77);
nand U17 (N_17,In_361,In_687);
and U18 (N_18,In_253,In_525);
and U19 (N_19,In_101,In_205);
or U20 (N_20,In_142,In_500);
nor U21 (N_21,In_473,In_743);
nor U22 (N_22,In_24,In_534);
nand U23 (N_23,In_181,In_492);
or U24 (N_24,In_128,In_489);
or U25 (N_25,In_299,In_593);
and U26 (N_26,In_678,In_449);
nor U27 (N_27,In_537,In_520);
or U28 (N_28,In_189,In_658);
nor U29 (N_29,In_691,In_303);
and U30 (N_30,In_356,In_481);
nor U31 (N_31,In_502,In_541);
nand U32 (N_32,In_201,In_592);
nor U33 (N_33,In_480,In_419);
nor U34 (N_34,In_531,In_222);
nand U35 (N_35,In_55,In_668);
nand U36 (N_36,In_187,In_385);
and U37 (N_37,In_600,In_718);
nor U38 (N_38,In_52,In_475);
nand U39 (N_39,In_85,In_508);
nor U40 (N_40,In_694,In_318);
or U41 (N_41,In_382,In_0);
nor U42 (N_42,In_643,In_190);
nand U43 (N_43,In_392,In_104);
or U44 (N_44,In_518,In_159);
and U45 (N_45,In_374,In_276);
and U46 (N_46,In_437,In_474);
and U47 (N_47,In_349,In_59);
and U48 (N_48,In_180,In_63);
and U49 (N_49,In_66,In_410);
and U50 (N_50,In_33,In_626);
or U51 (N_51,In_629,In_252);
nand U52 (N_52,In_554,In_417);
or U53 (N_53,In_582,In_35);
or U54 (N_54,In_423,In_549);
nor U55 (N_55,In_64,In_28);
or U56 (N_56,In_657,In_136);
or U57 (N_57,In_710,In_310);
nand U58 (N_58,In_34,In_367);
or U59 (N_59,In_606,In_133);
and U60 (N_60,In_642,In_383);
or U61 (N_61,In_357,In_169);
and U62 (N_62,In_209,In_441);
or U63 (N_63,In_655,In_337);
nand U64 (N_64,In_405,In_193);
or U65 (N_65,In_259,In_429);
nand U66 (N_66,In_664,In_47);
nand U67 (N_67,In_225,In_548);
or U68 (N_68,In_721,In_660);
or U69 (N_69,In_91,In_31);
and U70 (N_70,In_175,In_304);
nor U71 (N_71,In_350,In_238);
or U72 (N_72,In_154,In_1);
and U73 (N_73,In_714,In_191);
nand U74 (N_74,In_2,In_340);
or U75 (N_75,In_560,In_565);
nand U76 (N_76,In_211,In_711);
and U77 (N_77,In_239,In_375);
nor U78 (N_78,In_442,In_616);
nor U79 (N_79,In_21,In_503);
xor U80 (N_80,In_499,In_517);
nand U81 (N_81,In_632,In_308);
nand U82 (N_82,In_571,In_412);
nand U83 (N_83,In_79,In_727);
or U84 (N_84,In_649,In_272);
and U85 (N_85,In_654,In_697);
and U86 (N_86,In_624,In_81);
and U87 (N_87,In_168,In_333);
nand U88 (N_88,In_111,In_706);
nand U89 (N_89,In_359,In_279);
or U90 (N_90,In_670,In_148);
nor U91 (N_91,In_327,In_322);
nand U92 (N_92,In_583,In_149);
and U93 (N_93,In_484,In_637);
and U94 (N_94,In_745,In_703);
or U95 (N_95,In_73,In_87);
or U96 (N_96,In_741,In_155);
or U97 (N_97,In_716,In_603);
xnor U98 (N_98,In_158,In_666);
or U99 (N_99,In_604,In_354);
nor U100 (N_100,In_119,In_307);
nand U101 (N_101,In_455,In_365);
or U102 (N_102,In_432,In_720);
nor U103 (N_103,In_23,In_353);
nor U104 (N_104,In_132,In_709);
and U105 (N_105,In_546,In_14);
nor U106 (N_106,In_343,In_305);
or U107 (N_107,In_178,In_700);
nor U108 (N_108,In_690,In_110);
nor U109 (N_109,In_446,In_395);
or U110 (N_110,In_67,In_420);
or U111 (N_111,In_103,In_516);
nor U112 (N_112,In_617,In_182);
or U113 (N_113,In_647,In_575);
or U114 (N_114,In_522,In_498);
nor U115 (N_115,In_60,In_701);
nor U116 (N_116,In_139,In_324);
or U117 (N_117,In_94,In_366);
nand U118 (N_118,In_12,In_195);
or U119 (N_119,In_389,In_627);
nand U120 (N_120,In_287,In_373);
nor U121 (N_121,In_280,In_316);
and U122 (N_122,In_407,In_463);
nand U123 (N_123,In_39,In_730);
and U124 (N_124,In_218,In_335);
nand U125 (N_125,In_742,In_519);
nand U126 (N_126,In_220,In_271);
nor U127 (N_127,In_685,In_396);
nand U128 (N_128,In_105,In_114);
nand U129 (N_129,In_118,In_241);
nor U130 (N_130,In_598,In_384);
nor U131 (N_131,In_289,In_663);
nor U132 (N_132,In_50,In_746);
or U133 (N_133,In_436,In_521);
nand U134 (N_134,In_29,In_595);
nor U135 (N_135,In_633,In_341);
nand U136 (N_136,In_625,In_65);
and U137 (N_137,In_258,In_440);
nand U138 (N_138,In_151,In_409);
and U139 (N_139,In_696,In_58);
or U140 (N_140,In_411,In_292);
nand U141 (N_141,In_725,In_472);
or U142 (N_142,In_143,In_585);
nand U143 (N_143,In_295,In_479);
nand U144 (N_144,In_509,In_615);
and U145 (N_145,In_199,In_297);
and U146 (N_146,In_203,In_242);
or U147 (N_147,In_641,In_493);
and U148 (N_148,In_140,In_173);
nor U149 (N_149,In_27,In_360);
nor U150 (N_150,In_403,In_83);
or U151 (N_151,In_372,In_134);
nand U152 (N_152,In_49,In_216);
or U153 (N_153,In_11,In_511);
nand U154 (N_154,In_597,In_277);
nand U155 (N_155,In_646,In_547);
xnor U156 (N_156,In_402,In_273);
or U157 (N_157,In_179,In_530);
and U158 (N_158,In_732,In_426);
nand U159 (N_159,In_88,In_729);
or U160 (N_160,In_579,In_639);
nor U161 (N_161,In_48,In_213);
nor U162 (N_162,In_613,In_491);
nand U163 (N_163,In_458,In_683);
nand U164 (N_164,In_456,In_590);
or U165 (N_165,In_166,In_477);
nand U166 (N_166,In_397,In_676);
nand U167 (N_167,In_599,In_470);
nor U168 (N_168,In_284,In_505);
and U169 (N_169,In_527,In_197);
nand U170 (N_170,In_416,In_54);
or U171 (N_171,In_62,In_584);
and U172 (N_172,In_90,In_739);
or U173 (N_173,In_296,In_202);
or U174 (N_174,In_462,In_544);
nand U175 (N_175,In_468,In_724);
nor U176 (N_176,In_722,In_247);
nor U177 (N_177,In_636,In_97);
and U178 (N_178,In_338,In_635);
and U179 (N_179,In_37,In_30);
and U180 (N_180,In_427,In_109);
and U181 (N_181,In_726,In_144);
nor U182 (N_182,In_623,In_358);
or U183 (N_183,In_44,In_380);
nand U184 (N_184,In_323,In_351);
nor U185 (N_185,In_231,In_735);
and U186 (N_186,In_445,In_450);
nor U187 (N_187,In_659,In_749);
nor U188 (N_188,In_22,In_550);
nor U189 (N_189,In_589,In_306);
nor U190 (N_190,In_717,In_223);
or U191 (N_191,In_217,In_319);
nand U192 (N_192,In_390,In_192);
nor U193 (N_193,In_504,In_92);
and U194 (N_194,In_138,In_257);
nor U195 (N_195,In_609,In_112);
or U196 (N_196,In_265,In_733);
or U197 (N_197,In_125,In_290);
nand U198 (N_198,In_3,In_672);
nand U199 (N_199,In_102,In_236);
nor U200 (N_200,In_221,In_86);
nor U201 (N_201,In_495,In_130);
or U202 (N_202,In_736,In_347);
nand U203 (N_203,In_224,In_535);
nand U204 (N_204,In_577,In_457);
nor U205 (N_205,In_363,In_269);
and U206 (N_206,In_234,In_594);
nor U207 (N_207,In_237,In_131);
or U208 (N_208,In_38,In_692);
and U209 (N_209,In_653,In_334);
or U210 (N_210,In_553,In_557);
or U211 (N_211,In_215,In_418);
or U212 (N_212,In_688,In_170);
nand U213 (N_213,In_268,In_135);
or U214 (N_214,In_15,In_464);
nor U215 (N_215,In_43,In_248);
or U216 (N_216,In_20,In_123);
nand U217 (N_217,In_76,In_227);
nor U218 (N_218,In_438,In_70);
nor U219 (N_219,In_13,In_147);
nand U220 (N_220,In_294,In_152);
or U221 (N_221,In_129,In_387);
nor U222 (N_222,In_122,In_430);
or U223 (N_223,In_526,In_229);
and U224 (N_224,In_704,In_482);
or U225 (N_225,In_435,In_352);
and U226 (N_226,In_452,In_19);
nor U227 (N_227,In_567,In_57);
or U228 (N_228,In_302,In_528);
xnor U229 (N_229,In_561,In_748);
and U230 (N_230,In_232,In_26);
or U231 (N_231,In_460,In_620);
and U232 (N_232,In_42,In_78);
and U233 (N_233,In_486,In_283);
and U234 (N_234,In_431,In_562);
nand U235 (N_235,In_137,In_240);
nor U236 (N_236,In_578,In_249);
and U237 (N_237,In_740,In_93);
and U238 (N_238,In_574,In_428);
nand U239 (N_239,In_523,In_82);
nand U240 (N_240,In_424,In_538);
nand U241 (N_241,In_707,In_80);
nand U242 (N_242,In_719,In_686);
nand U243 (N_243,In_644,In_315);
nor U244 (N_244,In_98,In_210);
or U245 (N_245,In_84,In_391);
nand U246 (N_246,In_483,In_153);
or U247 (N_247,In_188,In_421);
or U248 (N_248,In_634,In_309);
nand U249 (N_249,In_621,In_747);
nor U250 (N_250,In_96,In_282);
and U251 (N_251,In_576,In_371);
nor U252 (N_252,In_293,In_61);
nor U253 (N_253,In_552,In_448);
nand U254 (N_254,In_36,In_443);
and U255 (N_255,In_494,In_618);
or U256 (N_256,In_558,In_563);
and U257 (N_257,In_399,In_117);
and U258 (N_258,In_453,In_75);
nor U259 (N_259,In_379,In_628);
nor U260 (N_260,In_362,In_246);
nand U261 (N_261,In_533,In_581);
or U262 (N_262,In_656,In_601);
or U263 (N_263,In_673,In_368);
and U264 (N_264,In_6,In_99);
xor U265 (N_265,In_512,In_51);
nand U266 (N_266,In_652,In_56);
and U267 (N_267,In_650,In_45);
nand U268 (N_268,In_9,In_524);
and U269 (N_269,In_731,In_674);
nor U270 (N_270,In_95,In_588);
or U271 (N_271,In_157,In_260);
or U272 (N_272,In_723,In_332);
or U273 (N_273,In_467,In_317);
nand U274 (N_274,In_364,In_566);
xnor U275 (N_275,In_214,In_602);
or U276 (N_276,In_619,In_532);
and U277 (N_277,In_233,In_551);
and U278 (N_278,In_121,In_556);
nor U279 (N_279,In_622,In_514);
nand U280 (N_280,In_146,In_439);
xnor U281 (N_281,In_400,In_198);
or U282 (N_282,In_734,In_465);
nor U283 (N_283,In_68,In_270);
or U284 (N_284,In_325,In_640);
and U285 (N_285,In_434,In_680);
nand U286 (N_286,In_377,In_469);
and U287 (N_287,In_422,In_207);
xor U288 (N_288,In_328,In_570);
nor U289 (N_289,In_346,In_244);
nor U290 (N_290,In_406,In_415);
xnor U291 (N_291,In_478,In_661);
nand U292 (N_292,In_261,In_728);
nor U293 (N_293,In_264,In_243);
or U294 (N_294,In_444,In_183);
nand U295 (N_295,In_580,In_7);
nand U296 (N_296,In_645,In_230);
xnor U297 (N_297,In_738,In_150);
nand U298 (N_298,In_200,In_219);
nor U299 (N_299,In_285,In_669);
nor U300 (N_300,In_507,In_681);
or U301 (N_301,In_605,In_689);
nor U302 (N_302,In_16,In_172);
nor U303 (N_303,In_342,In_607);
and U304 (N_304,In_540,In_206);
nor U305 (N_305,In_596,In_693);
or U306 (N_306,In_41,In_171);
nor U307 (N_307,In_235,In_196);
nor U308 (N_308,In_32,In_698);
or U309 (N_309,In_459,In_314);
nor U310 (N_310,In_106,In_263);
nand U311 (N_311,In_744,In_611);
nor U312 (N_312,In_141,In_559);
nor U313 (N_313,In_255,In_591);
nor U314 (N_314,In_490,In_100);
nand U315 (N_315,In_677,In_348);
or U316 (N_316,In_281,In_715);
and U317 (N_317,In_89,In_208);
nand U318 (N_318,In_665,In_254);
and U319 (N_319,In_278,In_275);
or U320 (N_320,In_321,In_331);
nand U321 (N_321,In_401,In_312);
or U322 (N_322,In_5,In_288);
or U323 (N_323,In_204,In_25);
and U324 (N_324,In_46,In_162);
and U325 (N_325,In_160,In_53);
and U326 (N_326,In_326,In_408);
and U327 (N_327,In_705,In_167);
or U328 (N_328,In_177,In_413);
nor U329 (N_329,In_69,In_339);
nor U330 (N_330,In_586,In_398);
and U331 (N_331,In_386,In_163);
nand U332 (N_332,In_497,In_447);
nand U333 (N_333,In_378,In_569);
and U334 (N_334,In_381,In_161);
and U335 (N_335,In_250,In_679);
nor U336 (N_336,In_737,In_568);
and U337 (N_337,In_513,In_488);
and U338 (N_338,In_176,In_274);
nor U339 (N_339,In_515,In_684);
nor U340 (N_340,In_18,In_245);
nand U341 (N_341,In_145,In_414);
or U342 (N_342,In_266,In_344);
nor U343 (N_343,In_506,In_330);
nand U344 (N_344,In_630,In_612);
or U345 (N_345,In_485,In_394);
nor U346 (N_346,In_115,In_501);
and U347 (N_347,In_124,In_699);
or U348 (N_348,In_376,In_451);
and U349 (N_349,In_298,In_487);
nand U350 (N_350,In_476,In_226);
nor U351 (N_351,In_671,In_587);
nor U352 (N_352,In_682,In_564);
or U353 (N_353,In_228,In_345);
nor U354 (N_354,In_186,In_164);
or U355 (N_355,In_608,In_631);
xor U356 (N_356,In_10,In_194);
nor U357 (N_357,In_355,In_212);
nand U358 (N_358,In_702,In_40);
nand U359 (N_359,In_174,In_712);
or U360 (N_360,In_667,In_256);
or U361 (N_361,In_74,In_108);
and U362 (N_362,In_388,In_675);
or U363 (N_363,In_529,In_313);
nor U364 (N_364,In_510,In_251);
and U365 (N_365,In_17,In_267);
xnor U366 (N_366,In_708,In_651);
and U367 (N_367,In_610,In_301);
nor U368 (N_368,In_393,In_116);
nand U369 (N_369,In_262,In_184);
nor U370 (N_370,In_466,In_542);
and U371 (N_371,In_543,In_404);
nand U372 (N_372,In_113,In_72);
and U373 (N_373,In_370,In_545);
or U374 (N_374,In_454,In_539);
or U375 (N_375,In_558,In_225);
and U376 (N_376,In_383,In_655);
nor U377 (N_377,In_461,In_186);
xor U378 (N_378,In_197,In_668);
nand U379 (N_379,In_549,In_664);
nand U380 (N_380,In_317,In_573);
or U381 (N_381,In_516,In_196);
nor U382 (N_382,In_29,In_467);
nor U383 (N_383,In_490,In_734);
and U384 (N_384,In_78,In_319);
xnor U385 (N_385,In_294,In_333);
nand U386 (N_386,In_164,In_94);
nand U387 (N_387,In_406,In_584);
and U388 (N_388,In_54,In_272);
and U389 (N_389,In_612,In_264);
nand U390 (N_390,In_486,In_364);
or U391 (N_391,In_444,In_205);
or U392 (N_392,In_13,In_527);
or U393 (N_393,In_437,In_79);
nand U394 (N_394,In_69,In_47);
and U395 (N_395,In_523,In_265);
and U396 (N_396,In_435,In_355);
and U397 (N_397,In_482,In_712);
nand U398 (N_398,In_330,In_549);
nand U399 (N_399,In_54,In_519);
and U400 (N_400,In_526,In_328);
or U401 (N_401,In_540,In_528);
nor U402 (N_402,In_632,In_644);
xor U403 (N_403,In_531,In_330);
xnor U404 (N_404,In_505,In_528);
nor U405 (N_405,In_576,In_162);
nor U406 (N_406,In_180,In_107);
nor U407 (N_407,In_264,In_16);
nor U408 (N_408,In_674,In_534);
nand U409 (N_409,In_734,In_516);
or U410 (N_410,In_625,In_614);
nor U411 (N_411,In_310,In_721);
and U412 (N_412,In_334,In_577);
nor U413 (N_413,In_645,In_152);
nand U414 (N_414,In_242,In_587);
or U415 (N_415,In_589,In_120);
nand U416 (N_416,In_182,In_94);
nor U417 (N_417,In_10,In_674);
nand U418 (N_418,In_114,In_633);
and U419 (N_419,In_198,In_266);
nand U420 (N_420,In_172,In_433);
nand U421 (N_421,In_592,In_54);
and U422 (N_422,In_231,In_745);
and U423 (N_423,In_113,In_263);
or U424 (N_424,In_205,In_358);
nor U425 (N_425,In_699,In_647);
nor U426 (N_426,In_663,In_407);
or U427 (N_427,In_93,In_341);
nand U428 (N_428,In_696,In_110);
nor U429 (N_429,In_671,In_83);
and U430 (N_430,In_648,In_221);
nand U431 (N_431,In_472,In_114);
and U432 (N_432,In_484,In_677);
nor U433 (N_433,In_120,In_318);
nor U434 (N_434,In_618,In_701);
nand U435 (N_435,In_28,In_492);
or U436 (N_436,In_292,In_611);
or U437 (N_437,In_200,In_465);
or U438 (N_438,In_370,In_430);
or U439 (N_439,In_58,In_371);
nor U440 (N_440,In_62,In_746);
nor U441 (N_441,In_208,In_589);
and U442 (N_442,In_614,In_393);
nor U443 (N_443,In_73,In_271);
xnor U444 (N_444,In_166,In_385);
or U445 (N_445,In_589,In_318);
and U446 (N_446,In_371,In_98);
nor U447 (N_447,In_583,In_592);
nand U448 (N_448,In_56,In_635);
nor U449 (N_449,In_629,In_704);
or U450 (N_450,In_681,In_642);
nor U451 (N_451,In_253,In_261);
nor U452 (N_452,In_413,In_343);
nand U453 (N_453,In_110,In_185);
or U454 (N_454,In_376,In_327);
xor U455 (N_455,In_717,In_124);
and U456 (N_456,In_686,In_683);
and U457 (N_457,In_427,In_657);
nor U458 (N_458,In_119,In_391);
nor U459 (N_459,In_53,In_79);
nand U460 (N_460,In_486,In_281);
nor U461 (N_461,In_61,In_630);
nor U462 (N_462,In_97,In_457);
nor U463 (N_463,In_648,In_140);
nor U464 (N_464,In_377,In_635);
nand U465 (N_465,In_744,In_259);
and U466 (N_466,In_67,In_532);
nand U467 (N_467,In_395,In_642);
or U468 (N_468,In_721,In_699);
nand U469 (N_469,In_712,In_436);
nand U470 (N_470,In_291,In_454);
nand U471 (N_471,In_29,In_378);
nand U472 (N_472,In_200,In_228);
or U473 (N_473,In_104,In_296);
nand U474 (N_474,In_267,In_426);
nand U475 (N_475,In_414,In_598);
or U476 (N_476,In_542,In_436);
or U477 (N_477,In_51,In_549);
or U478 (N_478,In_747,In_662);
and U479 (N_479,In_3,In_455);
or U480 (N_480,In_385,In_501);
nor U481 (N_481,In_285,In_465);
or U482 (N_482,In_359,In_3);
or U483 (N_483,In_123,In_558);
nand U484 (N_484,In_661,In_649);
nand U485 (N_485,In_408,In_394);
nor U486 (N_486,In_690,In_741);
nor U487 (N_487,In_30,In_207);
and U488 (N_488,In_134,In_386);
nand U489 (N_489,In_145,In_447);
and U490 (N_490,In_514,In_301);
nand U491 (N_491,In_372,In_726);
nand U492 (N_492,In_596,In_103);
nor U493 (N_493,In_26,In_385);
or U494 (N_494,In_374,In_249);
nand U495 (N_495,In_604,In_689);
and U496 (N_496,In_7,In_338);
nor U497 (N_497,In_36,In_372);
nor U498 (N_498,In_86,In_369);
and U499 (N_499,In_584,In_589);
or U500 (N_500,N_304,N_188);
nand U501 (N_501,N_299,N_444);
and U502 (N_502,N_193,N_442);
and U503 (N_503,N_359,N_405);
nand U504 (N_504,N_31,N_344);
nand U505 (N_505,N_92,N_77);
nor U506 (N_506,N_136,N_61);
and U507 (N_507,N_411,N_457);
and U508 (N_508,N_216,N_30);
nor U509 (N_509,N_182,N_176);
nor U510 (N_510,N_341,N_131);
or U511 (N_511,N_488,N_200);
or U512 (N_512,N_249,N_301);
nand U513 (N_513,N_361,N_74);
or U514 (N_514,N_379,N_451);
or U515 (N_515,N_478,N_288);
and U516 (N_516,N_35,N_48);
or U517 (N_517,N_422,N_171);
nor U518 (N_518,N_73,N_177);
nor U519 (N_519,N_192,N_204);
or U520 (N_520,N_102,N_272);
and U521 (N_521,N_378,N_179);
or U522 (N_522,N_205,N_42);
and U523 (N_523,N_101,N_401);
and U524 (N_524,N_116,N_195);
nor U525 (N_525,N_350,N_248);
and U526 (N_526,N_163,N_139);
or U527 (N_527,N_36,N_165);
and U528 (N_528,N_452,N_144);
and U529 (N_529,N_419,N_57);
and U530 (N_530,N_168,N_142);
nor U531 (N_531,N_231,N_292);
nor U532 (N_532,N_58,N_324);
nor U533 (N_533,N_426,N_275);
and U534 (N_534,N_151,N_16);
nor U535 (N_535,N_346,N_156);
or U536 (N_536,N_184,N_146);
nand U537 (N_537,N_269,N_384);
nor U538 (N_538,N_154,N_67);
nand U539 (N_539,N_187,N_4);
nand U540 (N_540,N_82,N_203);
nand U541 (N_541,N_477,N_239);
nand U542 (N_542,N_495,N_84);
nand U543 (N_543,N_313,N_402);
and U544 (N_544,N_268,N_392);
nor U545 (N_545,N_208,N_63);
nor U546 (N_546,N_110,N_99);
nand U547 (N_547,N_37,N_206);
and U548 (N_548,N_207,N_437);
nor U549 (N_549,N_271,N_215);
nand U550 (N_550,N_167,N_202);
and U551 (N_551,N_294,N_395);
and U552 (N_552,N_72,N_287);
nor U553 (N_553,N_62,N_240);
xor U554 (N_554,N_283,N_388);
or U555 (N_555,N_459,N_476);
and U556 (N_556,N_354,N_260);
and U557 (N_557,N_309,N_429);
nor U558 (N_558,N_50,N_302);
or U559 (N_559,N_129,N_172);
and U560 (N_560,N_219,N_396);
or U561 (N_561,N_64,N_486);
nand U562 (N_562,N_214,N_197);
nor U563 (N_563,N_482,N_98);
and U564 (N_564,N_170,N_270);
and U565 (N_565,N_161,N_81);
nor U566 (N_566,N_427,N_103);
nor U567 (N_567,N_499,N_27);
and U568 (N_568,N_487,N_367);
nand U569 (N_569,N_113,N_194);
or U570 (N_570,N_198,N_1);
nor U571 (N_571,N_261,N_316);
nand U572 (N_572,N_190,N_453);
nand U573 (N_573,N_162,N_211);
nand U574 (N_574,N_464,N_320);
or U575 (N_575,N_445,N_29);
nand U576 (N_576,N_138,N_147);
and U577 (N_577,N_463,N_212);
nor U578 (N_578,N_96,N_85);
and U579 (N_579,N_345,N_310);
or U580 (N_580,N_246,N_471);
nor U581 (N_581,N_185,N_125);
and U582 (N_582,N_278,N_493);
and U583 (N_583,N_276,N_404);
and U584 (N_584,N_80,N_347);
and U585 (N_585,N_264,N_335);
nor U586 (N_586,N_331,N_432);
or U587 (N_587,N_370,N_221);
nor U588 (N_588,N_155,N_173);
and U589 (N_589,N_191,N_230);
and U590 (N_590,N_224,N_52);
or U591 (N_591,N_130,N_91);
or U592 (N_592,N_222,N_468);
or U593 (N_593,N_252,N_2);
nor U594 (N_594,N_45,N_5);
or U595 (N_595,N_434,N_473);
nand U596 (N_596,N_90,N_472);
xor U597 (N_597,N_201,N_409);
and U598 (N_598,N_480,N_358);
nor U599 (N_599,N_238,N_68);
nand U600 (N_600,N_44,N_7);
nand U601 (N_601,N_466,N_108);
and U602 (N_602,N_104,N_189);
and U603 (N_603,N_412,N_49);
nor U604 (N_604,N_385,N_41);
nor U605 (N_605,N_181,N_314);
or U606 (N_606,N_100,N_234);
nand U607 (N_607,N_254,N_286);
or U608 (N_608,N_492,N_10);
nor U609 (N_609,N_306,N_343);
nor U610 (N_610,N_55,N_122);
nor U611 (N_611,N_220,N_484);
or U612 (N_612,N_20,N_134);
or U613 (N_613,N_218,N_400);
and U614 (N_614,N_428,N_75);
nor U615 (N_615,N_259,N_305);
nand U616 (N_616,N_496,N_417);
nand U617 (N_617,N_342,N_333);
nor U618 (N_618,N_114,N_469);
and U619 (N_619,N_387,N_263);
and U620 (N_620,N_8,N_356);
nand U621 (N_621,N_251,N_449);
xor U622 (N_622,N_430,N_9);
and U623 (N_623,N_365,N_3);
and U624 (N_624,N_17,N_180);
and U625 (N_625,N_112,N_307);
nor U626 (N_626,N_389,N_483);
nand U627 (N_627,N_415,N_284);
or U628 (N_628,N_298,N_321);
nor U629 (N_629,N_289,N_475);
or U630 (N_630,N_460,N_285);
and U631 (N_631,N_391,N_152);
nand U632 (N_632,N_235,N_351);
and U633 (N_633,N_330,N_209);
nor U634 (N_634,N_157,N_433);
nand U635 (N_635,N_258,N_76);
nand U636 (N_636,N_423,N_106);
or U637 (N_637,N_322,N_416);
and U638 (N_638,N_158,N_18);
and U639 (N_639,N_19,N_323);
or U640 (N_640,N_79,N_89);
or U641 (N_641,N_311,N_174);
nor U642 (N_642,N_140,N_153);
and U643 (N_643,N_373,N_266);
nand U644 (N_644,N_15,N_223);
nor U645 (N_645,N_282,N_353);
nand U646 (N_646,N_420,N_34);
xor U647 (N_647,N_414,N_47);
nand U648 (N_648,N_312,N_148);
nor U649 (N_649,N_94,N_436);
nor U650 (N_650,N_424,N_86);
nor U651 (N_651,N_107,N_454);
nand U652 (N_652,N_315,N_127);
or U653 (N_653,N_348,N_355);
and U654 (N_654,N_93,N_325);
and U655 (N_655,N_295,N_447);
or U656 (N_656,N_25,N_88);
nand U657 (N_657,N_393,N_357);
nor U658 (N_658,N_54,N_175);
or U659 (N_659,N_78,N_124);
nand U660 (N_660,N_32,N_0);
and U661 (N_661,N_274,N_398);
nor U662 (N_662,N_450,N_183);
and U663 (N_663,N_83,N_440);
and U664 (N_664,N_303,N_253);
nand U665 (N_665,N_439,N_326);
or U666 (N_666,N_40,N_228);
or U667 (N_667,N_470,N_149);
and U668 (N_668,N_115,N_105);
and U669 (N_669,N_229,N_267);
or U670 (N_670,N_280,N_245);
and U671 (N_671,N_236,N_403);
and U672 (N_672,N_293,N_51);
or U673 (N_673,N_12,N_374);
nor U674 (N_674,N_242,N_407);
or U675 (N_675,N_372,N_145);
and U676 (N_676,N_133,N_128);
and U677 (N_677,N_26,N_87);
nor U678 (N_678,N_24,N_338);
nand U679 (N_679,N_352,N_399);
or U680 (N_680,N_362,N_441);
nand U681 (N_681,N_132,N_435);
and U682 (N_682,N_377,N_277);
nand U683 (N_683,N_413,N_196);
and U684 (N_684,N_425,N_366);
or U685 (N_685,N_497,N_244);
or U686 (N_686,N_364,N_141);
or U687 (N_687,N_166,N_467);
nand U688 (N_688,N_498,N_247);
or U689 (N_689,N_406,N_21);
nand U690 (N_690,N_296,N_390);
nor U691 (N_691,N_226,N_494);
nand U692 (N_692,N_22,N_59);
and U693 (N_693,N_70,N_458);
or U694 (N_694,N_199,N_250);
nor U695 (N_695,N_371,N_318);
nand U696 (N_696,N_186,N_438);
xor U697 (N_697,N_349,N_394);
or U698 (N_698,N_290,N_479);
or U699 (N_699,N_448,N_137);
and U700 (N_700,N_317,N_337);
nor U701 (N_701,N_273,N_39);
and U702 (N_702,N_164,N_485);
or U703 (N_703,N_6,N_474);
nand U704 (N_704,N_397,N_23);
and U705 (N_705,N_363,N_360);
nand U706 (N_706,N_66,N_56);
nand U707 (N_707,N_160,N_443);
xnor U708 (N_708,N_227,N_256);
or U709 (N_709,N_334,N_233);
or U710 (N_710,N_386,N_13);
and U711 (N_711,N_237,N_418);
and U712 (N_712,N_69,N_169);
xor U713 (N_713,N_465,N_232);
nand U714 (N_714,N_241,N_421);
nand U715 (N_715,N_210,N_46);
or U716 (N_716,N_382,N_119);
nand U717 (N_717,N_143,N_28);
nand U718 (N_718,N_53,N_265);
nor U719 (N_719,N_375,N_38);
nand U720 (N_720,N_490,N_213);
and U721 (N_721,N_262,N_217);
and U722 (N_722,N_95,N_178);
or U723 (N_723,N_328,N_257);
or U724 (N_724,N_369,N_117);
nor U725 (N_725,N_135,N_491);
and U726 (N_726,N_118,N_123);
nor U727 (N_727,N_60,N_43);
or U728 (N_728,N_71,N_381);
nand U729 (N_729,N_339,N_383);
nand U730 (N_730,N_481,N_446);
or U731 (N_731,N_109,N_14);
nand U732 (N_732,N_225,N_243);
nor U733 (N_733,N_33,N_120);
or U734 (N_734,N_336,N_111);
nor U735 (N_735,N_456,N_461);
nor U736 (N_736,N_327,N_368);
nand U737 (N_737,N_11,N_300);
and U738 (N_738,N_462,N_281);
and U739 (N_739,N_255,N_126);
nor U740 (N_740,N_297,N_332);
nand U741 (N_741,N_150,N_455);
or U742 (N_742,N_489,N_408);
and U743 (N_743,N_97,N_410);
and U744 (N_744,N_65,N_376);
nor U745 (N_745,N_291,N_329);
nor U746 (N_746,N_319,N_121);
and U747 (N_747,N_279,N_380);
and U748 (N_748,N_308,N_159);
nor U749 (N_749,N_431,N_340);
or U750 (N_750,N_300,N_141);
and U751 (N_751,N_263,N_352);
and U752 (N_752,N_20,N_435);
and U753 (N_753,N_56,N_127);
xor U754 (N_754,N_423,N_203);
or U755 (N_755,N_283,N_343);
nand U756 (N_756,N_19,N_376);
and U757 (N_757,N_314,N_397);
and U758 (N_758,N_483,N_223);
and U759 (N_759,N_238,N_53);
and U760 (N_760,N_183,N_151);
nand U761 (N_761,N_343,N_86);
nand U762 (N_762,N_199,N_277);
nor U763 (N_763,N_22,N_345);
nand U764 (N_764,N_469,N_449);
and U765 (N_765,N_269,N_445);
and U766 (N_766,N_112,N_148);
nand U767 (N_767,N_284,N_14);
or U768 (N_768,N_151,N_489);
and U769 (N_769,N_62,N_252);
nand U770 (N_770,N_424,N_94);
or U771 (N_771,N_466,N_411);
nand U772 (N_772,N_403,N_286);
nor U773 (N_773,N_147,N_92);
xor U774 (N_774,N_369,N_486);
and U775 (N_775,N_185,N_15);
nand U776 (N_776,N_150,N_125);
and U777 (N_777,N_197,N_336);
nand U778 (N_778,N_289,N_50);
or U779 (N_779,N_117,N_144);
or U780 (N_780,N_255,N_25);
nor U781 (N_781,N_329,N_499);
and U782 (N_782,N_487,N_303);
nand U783 (N_783,N_34,N_8);
and U784 (N_784,N_226,N_472);
nand U785 (N_785,N_168,N_188);
or U786 (N_786,N_258,N_152);
and U787 (N_787,N_420,N_73);
nand U788 (N_788,N_494,N_61);
nor U789 (N_789,N_420,N_447);
and U790 (N_790,N_171,N_426);
nand U791 (N_791,N_256,N_401);
nand U792 (N_792,N_222,N_52);
nand U793 (N_793,N_225,N_419);
nor U794 (N_794,N_135,N_329);
nand U795 (N_795,N_80,N_277);
nand U796 (N_796,N_339,N_153);
nor U797 (N_797,N_8,N_257);
nand U798 (N_798,N_6,N_448);
nand U799 (N_799,N_238,N_355);
or U800 (N_800,N_372,N_116);
nor U801 (N_801,N_7,N_323);
nand U802 (N_802,N_143,N_310);
or U803 (N_803,N_191,N_81);
nand U804 (N_804,N_242,N_174);
or U805 (N_805,N_128,N_368);
nor U806 (N_806,N_217,N_200);
or U807 (N_807,N_70,N_202);
nor U808 (N_808,N_386,N_11);
and U809 (N_809,N_337,N_251);
nand U810 (N_810,N_187,N_171);
nor U811 (N_811,N_498,N_171);
and U812 (N_812,N_63,N_481);
nor U813 (N_813,N_331,N_116);
and U814 (N_814,N_44,N_471);
and U815 (N_815,N_479,N_424);
or U816 (N_816,N_350,N_200);
or U817 (N_817,N_99,N_363);
or U818 (N_818,N_94,N_119);
and U819 (N_819,N_45,N_217);
nand U820 (N_820,N_264,N_436);
nand U821 (N_821,N_256,N_235);
nand U822 (N_822,N_328,N_409);
nand U823 (N_823,N_101,N_496);
nor U824 (N_824,N_59,N_90);
nor U825 (N_825,N_68,N_346);
nand U826 (N_826,N_342,N_372);
nand U827 (N_827,N_98,N_317);
nor U828 (N_828,N_265,N_366);
and U829 (N_829,N_76,N_461);
nand U830 (N_830,N_487,N_431);
and U831 (N_831,N_331,N_400);
and U832 (N_832,N_423,N_174);
xor U833 (N_833,N_205,N_211);
nand U834 (N_834,N_188,N_181);
nor U835 (N_835,N_56,N_132);
nor U836 (N_836,N_315,N_215);
nand U837 (N_837,N_335,N_384);
and U838 (N_838,N_241,N_418);
and U839 (N_839,N_93,N_187);
nor U840 (N_840,N_262,N_174);
nand U841 (N_841,N_436,N_377);
nand U842 (N_842,N_426,N_314);
or U843 (N_843,N_180,N_429);
or U844 (N_844,N_169,N_184);
and U845 (N_845,N_33,N_243);
nand U846 (N_846,N_449,N_80);
nand U847 (N_847,N_39,N_306);
nand U848 (N_848,N_387,N_388);
and U849 (N_849,N_333,N_154);
and U850 (N_850,N_224,N_22);
nor U851 (N_851,N_353,N_448);
nor U852 (N_852,N_125,N_53);
xor U853 (N_853,N_447,N_59);
and U854 (N_854,N_264,N_38);
nor U855 (N_855,N_208,N_428);
and U856 (N_856,N_391,N_21);
or U857 (N_857,N_422,N_131);
and U858 (N_858,N_395,N_56);
nand U859 (N_859,N_434,N_367);
nand U860 (N_860,N_400,N_129);
and U861 (N_861,N_352,N_185);
xnor U862 (N_862,N_182,N_256);
or U863 (N_863,N_485,N_288);
nand U864 (N_864,N_326,N_155);
nor U865 (N_865,N_460,N_240);
nand U866 (N_866,N_273,N_452);
nand U867 (N_867,N_212,N_168);
or U868 (N_868,N_366,N_485);
and U869 (N_869,N_495,N_187);
xnor U870 (N_870,N_106,N_377);
nand U871 (N_871,N_442,N_369);
and U872 (N_872,N_222,N_293);
nor U873 (N_873,N_410,N_443);
or U874 (N_874,N_131,N_254);
nand U875 (N_875,N_278,N_237);
nor U876 (N_876,N_193,N_321);
or U877 (N_877,N_291,N_469);
nand U878 (N_878,N_288,N_305);
or U879 (N_879,N_103,N_82);
and U880 (N_880,N_2,N_168);
or U881 (N_881,N_106,N_256);
nand U882 (N_882,N_198,N_323);
and U883 (N_883,N_9,N_384);
nor U884 (N_884,N_317,N_479);
nor U885 (N_885,N_228,N_191);
nor U886 (N_886,N_263,N_441);
and U887 (N_887,N_267,N_130);
or U888 (N_888,N_12,N_124);
and U889 (N_889,N_21,N_402);
nand U890 (N_890,N_387,N_187);
nor U891 (N_891,N_484,N_351);
nor U892 (N_892,N_352,N_102);
nand U893 (N_893,N_67,N_105);
nand U894 (N_894,N_467,N_142);
and U895 (N_895,N_195,N_86);
or U896 (N_896,N_427,N_312);
and U897 (N_897,N_99,N_128);
nor U898 (N_898,N_474,N_379);
or U899 (N_899,N_98,N_438);
and U900 (N_900,N_171,N_179);
nor U901 (N_901,N_14,N_116);
and U902 (N_902,N_113,N_354);
or U903 (N_903,N_346,N_143);
nand U904 (N_904,N_211,N_493);
nand U905 (N_905,N_271,N_350);
nand U906 (N_906,N_399,N_462);
or U907 (N_907,N_446,N_194);
or U908 (N_908,N_449,N_87);
nor U909 (N_909,N_258,N_274);
nand U910 (N_910,N_475,N_224);
nor U911 (N_911,N_167,N_7);
nor U912 (N_912,N_279,N_396);
and U913 (N_913,N_326,N_309);
or U914 (N_914,N_403,N_30);
nand U915 (N_915,N_268,N_420);
or U916 (N_916,N_289,N_37);
or U917 (N_917,N_143,N_314);
and U918 (N_918,N_330,N_342);
or U919 (N_919,N_309,N_260);
nand U920 (N_920,N_228,N_462);
nor U921 (N_921,N_263,N_87);
or U922 (N_922,N_15,N_193);
and U923 (N_923,N_87,N_12);
and U924 (N_924,N_97,N_4);
nor U925 (N_925,N_36,N_124);
xnor U926 (N_926,N_478,N_499);
and U927 (N_927,N_118,N_284);
and U928 (N_928,N_119,N_409);
and U929 (N_929,N_476,N_397);
nor U930 (N_930,N_118,N_454);
and U931 (N_931,N_317,N_482);
nand U932 (N_932,N_375,N_427);
or U933 (N_933,N_185,N_228);
xor U934 (N_934,N_410,N_221);
nand U935 (N_935,N_263,N_54);
and U936 (N_936,N_51,N_336);
nor U937 (N_937,N_97,N_443);
nand U938 (N_938,N_339,N_361);
nor U939 (N_939,N_256,N_402);
or U940 (N_940,N_269,N_12);
nand U941 (N_941,N_410,N_319);
and U942 (N_942,N_429,N_265);
and U943 (N_943,N_115,N_289);
nor U944 (N_944,N_177,N_454);
or U945 (N_945,N_24,N_442);
or U946 (N_946,N_454,N_415);
nand U947 (N_947,N_352,N_36);
xnor U948 (N_948,N_210,N_373);
nor U949 (N_949,N_277,N_252);
nor U950 (N_950,N_168,N_194);
nor U951 (N_951,N_495,N_62);
nor U952 (N_952,N_28,N_37);
nand U953 (N_953,N_354,N_40);
and U954 (N_954,N_443,N_291);
or U955 (N_955,N_145,N_59);
or U956 (N_956,N_41,N_152);
or U957 (N_957,N_254,N_363);
and U958 (N_958,N_20,N_229);
or U959 (N_959,N_168,N_40);
or U960 (N_960,N_4,N_365);
and U961 (N_961,N_397,N_468);
or U962 (N_962,N_299,N_481);
nor U963 (N_963,N_255,N_372);
or U964 (N_964,N_477,N_62);
or U965 (N_965,N_301,N_153);
or U966 (N_966,N_189,N_50);
or U967 (N_967,N_71,N_99);
or U968 (N_968,N_211,N_70);
nand U969 (N_969,N_434,N_465);
or U970 (N_970,N_432,N_56);
or U971 (N_971,N_69,N_415);
and U972 (N_972,N_177,N_169);
nand U973 (N_973,N_442,N_434);
or U974 (N_974,N_369,N_226);
or U975 (N_975,N_9,N_227);
nand U976 (N_976,N_34,N_55);
or U977 (N_977,N_315,N_447);
or U978 (N_978,N_364,N_306);
nand U979 (N_979,N_416,N_392);
nand U980 (N_980,N_122,N_323);
nor U981 (N_981,N_282,N_271);
or U982 (N_982,N_34,N_58);
or U983 (N_983,N_138,N_283);
or U984 (N_984,N_211,N_389);
nand U985 (N_985,N_175,N_405);
nor U986 (N_986,N_290,N_90);
or U987 (N_987,N_104,N_402);
or U988 (N_988,N_110,N_336);
and U989 (N_989,N_96,N_143);
nor U990 (N_990,N_51,N_467);
and U991 (N_991,N_151,N_359);
nand U992 (N_992,N_198,N_438);
or U993 (N_993,N_301,N_137);
or U994 (N_994,N_476,N_183);
or U995 (N_995,N_226,N_323);
or U996 (N_996,N_209,N_377);
or U997 (N_997,N_63,N_422);
or U998 (N_998,N_455,N_477);
nand U999 (N_999,N_109,N_201);
nor U1000 (N_1000,N_826,N_651);
or U1001 (N_1001,N_657,N_891);
nand U1002 (N_1002,N_670,N_612);
nor U1003 (N_1003,N_985,N_962);
and U1004 (N_1004,N_923,N_789);
and U1005 (N_1005,N_580,N_759);
nand U1006 (N_1006,N_783,N_882);
nor U1007 (N_1007,N_859,N_796);
and U1008 (N_1008,N_705,N_729);
and U1009 (N_1009,N_945,N_976);
nand U1010 (N_1010,N_963,N_685);
and U1011 (N_1011,N_860,N_678);
or U1012 (N_1012,N_558,N_509);
and U1013 (N_1013,N_866,N_653);
nor U1014 (N_1014,N_706,N_782);
and U1015 (N_1015,N_843,N_936);
or U1016 (N_1016,N_967,N_553);
or U1017 (N_1017,N_850,N_511);
nor U1018 (N_1018,N_590,N_507);
and U1019 (N_1019,N_792,N_926);
xor U1020 (N_1020,N_500,N_531);
or U1021 (N_1021,N_520,N_535);
nand U1022 (N_1022,N_727,N_745);
nor U1023 (N_1023,N_547,N_775);
or U1024 (N_1024,N_510,N_751);
nor U1025 (N_1025,N_668,N_719);
or U1026 (N_1026,N_947,N_608);
and U1027 (N_1027,N_695,N_694);
nor U1028 (N_1028,N_752,N_624);
and U1029 (N_1029,N_944,N_832);
and U1030 (N_1030,N_573,N_674);
nor U1031 (N_1031,N_616,N_819);
nor U1032 (N_1032,N_880,N_790);
nor U1033 (N_1033,N_574,N_878);
nand U1034 (N_1034,N_677,N_918);
or U1035 (N_1035,N_822,N_630);
and U1036 (N_1036,N_721,N_606);
nand U1037 (N_1037,N_786,N_925);
or U1038 (N_1038,N_849,N_995);
and U1039 (N_1039,N_941,N_801);
nand U1040 (N_1040,N_662,N_516);
and U1041 (N_1041,N_858,N_997);
and U1042 (N_1042,N_907,N_597);
or U1043 (N_1043,N_897,N_660);
or U1044 (N_1044,N_802,N_661);
or U1045 (N_1045,N_732,N_702);
nand U1046 (N_1046,N_692,N_975);
xor U1047 (N_1047,N_886,N_579);
nor U1048 (N_1048,N_901,N_834);
or U1049 (N_1049,N_546,N_628);
and U1050 (N_1050,N_996,N_737);
or U1051 (N_1051,N_675,N_765);
nor U1052 (N_1052,N_581,N_687);
and U1053 (N_1053,N_747,N_723);
nand U1054 (N_1054,N_830,N_935);
nand U1055 (N_1055,N_753,N_603);
nand U1056 (N_1056,N_504,N_621);
and U1057 (N_1057,N_631,N_939);
and U1058 (N_1058,N_641,N_735);
nor U1059 (N_1059,N_593,N_549);
and U1060 (N_1060,N_742,N_953);
nand U1061 (N_1061,N_811,N_512);
nor U1062 (N_1062,N_650,N_998);
or U1063 (N_1063,N_681,N_848);
nor U1064 (N_1064,N_679,N_844);
nor U1065 (N_1065,N_760,N_680);
or U1066 (N_1066,N_835,N_594);
nand U1067 (N_1067,N_562,N_942);
nor U1068 (N_1068,N_929,N_572);
xor U1069 (N_1069,N_666,N_781);
nor U1070 (N_1070,N_837,N_618);
or U1071 (N_1071,N_887,N_709);
nand U1072 (N_1072,N_770,N_733);
nor U1073 (N_1073,N_526,N_851);
nand U1074 (N_1074,N_649,N_924);
or U1075 (N_1075,N_906,N_689);
nor U1076 (N_1076,N_656,N_805);
or U1077 (N_1077,N_505,N_896);
and U1078 (N_1078,N_913,N_537);
or U1079 (N_1079,N_544,N_845);
nor U1080 (N_1080,N_600,N_575);
nor U1081 (N_1081,N_922,N_712);
and U1082 (N_1082,N_734,N_632);
nand U1083 (N_1083,N_988,N_809);
or U1084 (N_1084,N_556,N_599);
or U1085 (N_1085,N_639,N_838);
and U1086 (N_1086,N_688,N_927);
and U1087 (N_1087,N_989,N_784);
and U1088 (N_1088,N_700,N_964);
or U1089 (N_1089,N_979,N_652);
nor U1090 (N_1090,N_748,N_771);
or U1091 (N_1091,N_539,N_659);
nor U1092 (N_1092,N_949,N_855);
or U1093 (N_1093,N_852,N_841);
xor U1094 (N_1094,N_726,N_758);
and U1095 (N_1095,N_648,N_570);
and U1096 (N_1096,N_808,N_810);
nor U1097 (N_1097,N_686,N_730);
nand U1098 (N_1098,N_676,N_794);
nor U1099 (N_1099,N_961,N_803);
and U1100 (N_1100,N_816,N_591);
xor U1101 (N_1101,N_763,N_501);
nand U1102 (N_1102,N_738,N_853);
nand U1103 (N_1103,N_946,N_746);
and U1104 (N_1104,N_879,N_950);
nand U1105 (N_1105,N_971,N_807);
nand U1106 (N_1106,N_561,N_821);
or U1107 (N_1107,N_958,N_595);
nand U1108 (N_1108,N_981,N_533);
nand U1109 (N_1109,N_955,N_614);
xnor U1110 (N_1110,N_525,N_536);
and U1111 (N_1111,N_892,N_540);
and U1112 (N_1112,N_559,N_937);
or U1113 (N_1113,N_987,N_508);
and U1114 (N_1114,N_750,N_761);
nor U1115 (N_1115,N_517,N_744);
nor U1116 (N_1116,N_611,N_881);
nand U1117 (N_1117,N_890,N_833);
nand U1118 (N_1118,N_633,N_635);
or U1119 (N_1119,N_827,N_625);
nand U1120 (N_1120,N_952,N_671);
nor U1121 (N_1121,N_626,N_663);
nand U1122 (N_1122,N_613,N_779);
or U1123 (N_1123,N_969,N_883);
nand U1124 (N_1124,N_978,N_968);
nor U1125 (N_1125,N_982,N_514);
nor U1126 (N_1126,N_715,N_755);
nor U1127 (N_1127,N_785,N_867);
nor U1128 (N_1128,N_993,N_584);
and U1129 (N_1129,N_788,N_557);
and U1130 (N_1130,N_956,N_567);
nor U1131 (N_1131,N_903,N_583);
nor U1132 (N_1132,N_701,N_601);
nor U1133 (N_1133,N_542,N_908);
nor U1134 (N_1134,N_823,N_768);
or U1135 (N_1135,N_502,N_566);
nor U1136 (N_1136,N_899,N_787);
nor U1137 (N_1137,N_762,N_813);
or U1138 (N_1138,N_840,N_871);
nor U1139 (N_1139,N_872,N_919);
or U1140 (N_1140,N_538,N_828);
and U1141 (N_1141,N_806,N_916);
and U1142 (N_1142,N_839,N_900);
nand U1143 (N_1143,N_615,N_889);
nand U1144 (N_1144,N_707,N_864);
nand U1145 (N_1145,N_912,N_731);
nand U1146 (N_1146,N_904,N_587);
nand U1147 (N_1147,N_696,N_829);
or U1148 (N_1148,N_902,N_644);
nand U1149 (N_1149,N_836,N_767);
and U1150 (N_1150,N_994,N_856);
nand U1151 (N_1151,N_921,N_714);
or U1152 (N_1152,N_999,N_716);
nor U1153 (N_1153,N_960,N_820);
and U1154 (N_1154,N_527,N_711);
nor U1155 (N_1155,N_645,N_812);
or U1156 (N_1156,N_776,N_847);
and U1157 (N_1157,N_754,N_636);
nand U1158 (N_1158,N_992,N_757);
or U1159 (N_1159,N_778,N_610);
and U1160 (N_1160,N_647,N_973);
nand U1161 (N_1161,N_582,N_586);
nor U1162 (N_1162,N_724,N_965);
nor U1163 (N_1163,N_629,N_563);
nand U1164 (N_1164,N_914,N_915);
xor U1165 (N_1165,N_898,N_515);
nand U1166 (N_1166,N_532,N_725);
nand U1167 (N_1167,N_602,N_984);
nor U1168 (N_1168,N_605,N_798);
or U1169 (N_1169,N_565,N_831);
or U1170 (N_1170,N_777,N_620);
or U1171 (N_1171,N_703,N_736);
or U1172 (N_1172,N_654,N_699);
nand U1173 (N_1173,N_627,N_682);
nor U1174 (N_1174,N_773,N_983);
nor U1175 (N_1175,N_576,N_970);
and U1176 (N_1176,N_642,N_909);
nand U1177 (N_1177,N_932,N_691);
or U1178 (N_1178,N_846,N_869);
or U1179 (N_1179,N_954,N_643);
nor U1180 (N_1180,N_664,N_519);
nand U1181 (N_1181,N_861,N_571);
nand U1182 (N_1182,N_569,N_815);
nand U1183 (N_1183,N_588,N_905);
or U1184 (N_1184,N_717,N_780);
nand U1185 (N_1185,N_877,N_894);
and U1186 (N_1186,N_534,N_528);
nor U1187 (N_1187,N_740,N_797);
nor U1188 (N_1188,N_545,N_552);
nand U1189 (N_1189,N_658,N_818);
and U1190 (N_1190,N_885,N_518);
or U1191 (N_1191,N_638,N_917);
or U1192 (N_1192,N_772,N_795);
nor U1193 (N_1193,N_870,N_920);
nand U1194 (N_1194,N_617,N_910);
nor U1195 (N_1195,N_577,N_764);
nand U1196 (N_1196,N_598,N_766);
or U1197 (N_1197,N_911,N_959);
nand U1198 (N_1198,N_875,N_986);
nor U1199 (N_1199,N_708,N_690);
or U1200 (N_1200,N_693,N_943);
and U1201 (N_1201,N_554,N_607);
or U1202 (N_1202,N_928,N_938);
or U1203 (N_1203,N_739,N_550);
xnor U1204 (N_1204,N_673,N_895);
and U1205 (N_1205,N_854,N_933);
nor U1206 (N_1206,N_756,N_560);
or U1207 (N_1207,N_966,N_722);
nand U1208 (N_1208,N_930,N_622);
nand U1209 (N_1209,N_634,N_957);
nand U1210 (N_1210,N_974,N_804);
nand U1211 (N_1211,N_698,N_585);
and U1212 (N_1212,N_876,N_684);
and U1213 (N_1213,N_541,N_506);
nor U1214 (N_1214,N_713,N_683);
or U1215 (N_1215,N_874,N_948);
nand U1216 (N_1216,N_825,N_743);
nand U1217 (N_1217,N_503,N_749);
or U1218 (N_1218,N_548,N_513);
nand U1219 (N_1219,N_523,N_972);
nor U1220 (N_1220,N_791,N_991);
nand U1221 (N_1221,N_980,N_863);
or U1222 (N_1222,N_718,N_604);
xnor U1223 (N_1223,N_868,N_619);
nor U1224 (N_1224,N_589,N_951);
nand U1225 (N_1225,N_741,N_873);
nand U1226 (N_1226,N_551,N_522);
and U1227 (N_1227,N_530,N_710);
nor U1228 (N_1228,N_637,N_842);
or U1229 (N_1229,N_728,N_555);
and U1230 (N_1230,N_521,N_931);
or U1231 (N_1231,N_529,N_568);
and U1232 (N_1232,N_814,N_609);
nor U1233 (N_1233,N_799,N_667);
nor U1234 (N_1234,N_884,N_793);
nor U1235 (N_1235,N_893,N_940);
nor U1236 (N_1236,N_857,N_774);
nand U1237 (N_1237,N_817,N_977);
nor U1238 (N_1238,N_640,N_800);
nor U1239 (N_1239,N_543,N_824);
nor U1240 (N_1240,N_655,N_934);
nand U1241 (N_1241,N_669,N_564);
nand U1242 (N_1242,N_862,N_697);
nand U1243 (N_1243,N_665,N_990);
and U1244 (N_1244,N_592,N_865);
and U1245 (N_1245,N_672,N_720);
nor U1246 (N_1246,N_769,N_524);
nor U1247 (N_1247,N_596,N_704);
nor U1248 (N_1248,N_646,N_623);
nor U1249 (N_1249,N_578,N_888);
nand U1250 (N_1250,N_750,N_757);
and U1251 (N_1251,N_781,N_566);
nor U1252 (N_1252,N_623,N_769);
or U1253 (N_1253,N_996,N_925);
nand U1254 (N_1254,N_951,N_932);
or U1255 (N_1255,N_932,N_767);
or U1256 (N_1256,N_806,N_899);
nor U1257 (N_1257,N_877,N_721);
nand U1258 (N_1258,N_685,N_631);
nor U1259 (N_1259,N_927,N_795);
or U1260 (N_1260,N_966,N_757);
or U1261 (N_1261,N_931,N_873);
or U1262 (N_1262,N_519,N_775);
nand U1263 (N_1263,N_591,N_802);
nor U1264 (N_1264,N_630,N_632);
and U1265 (N_1265,N_953,N_902);
nand U1266 (N_1266,N_941,N_992);
xor U1267 (N_1267,N_808,N_777);
nor U1268 (N_1268,N_681,N_867);
or U1269 (N_1269,N_578,N_873);
or U1270 (N_1270,N_598,N_788);
or U1271 (N_1271,N_654,N_951);
or U1272 (N_1272,N_594,N_677);
or U1273 (N_1273,N_638,N_568);
and U1274 (N_1274,N_822,N_643);
or U1275 (N_1275,N_672,N_784);
xor U1276 (N_1276,N_727,N_673);
nor U1277 (N_1277,N_817,N_710);
nor U1278 (N_1278,N_576,N_677);
or U1279 (N_1279,N_741,N_911);
nor U1280 (N_1280,N_682,N_500);
and U1281 (N_1281,N_929,N_779);
and U1282 (N_1282,N_936,N_855);
and U1283 (N_1283,N_864,N_769);
and U1284 (N_1284,N_892,N_614);
or U1285 (N_1285,N_955,N_755);
and U1286 (N_1286,N_657,N_964);
or U1287 (N_1287,N_848,N_742);
or U1288 (N_1288,N_783,N_719);
and U1289 (N_1289,N_584,N_916);
nor U1290 (N_1290,N_604,N_829);
or U1291 (N_1291,N_919,N_907);
and U1292 (N_1292,N_796,N_928);
nor U1293 (N_1293,N_709,N_865);
or U1294 (N_1294,N_720,N_588);
nor U1295 (N_1295,N_687,N_882);
and U1296 (N_1296,N_755,N_825);
nand U1297 (N_1297,N_569,N_650);
nand U1298 (N_1298,N_681,N_630);
nand U1299 (N_1299,N_841,N_843);
nor U1300 (N_1300,N_515,N_760);
and U1301 (N_1301,N_791,N_863);
and U1302 (N_1302,N_671,N_752);
or U1303 (N_1303,N_714,N_553);
nand U1304 (N_1304,N_939,N_574);
nor U1305 (N_1305,N_946,N_989);
or U1306 (N_1306,N_973,N_732);
nand U1307 (N_1307,N_618,N_563);
nand U1308 (N_1308,N_925,N_824);
and U1309 (N_1309,N_575,N_890);
and U1310 (N_1310,N_863,N_575);
xnor U1311 (N_1311,N_570,N_701);
nand U1312 (N_1312,N_731,N_899);
nor U1313 (N_1313,N_820,N_800);
nand U1314 (N_1314,N_685,N_944);
nor U1315 (N_1315,N_614,N_645);
and U1316 (N_1316,N_983,N_695);
and U1317 (N_1317,N_942,N_521);
or U1318 (N_1318,N_613,N_572);
nor U1319 (N_1319,N_824,N_821);
nand U1320 (N_1320,N_776,N_552);
nor U1321 (N_1321,N_975,N_684);
or U1322 (N_1322,N_662,N_609);
nor U1323 (N_1323,N_962,N_731);
nand U1324 (N_1324,N_689,N_519);
nor U1325 (N_1325,N_606,N_697);
and U1326 (N_1326,N_704,N_907);
and U1327 (N_1327,N_571,N_767);
nand U1328 (N_1328,N_540,N_847);
nor U1329 (N_1329,N_675,N_900);
nand U1330 (N_1330,N_673,N_594);
nand U1331 (N_1331,N_620,N_632);
and U1332 (N_1332,N_942,N_934);
xnor U1333 (N_1333,N_605,N_995);
or U1334 (N_1334,N_637,N_642);
nor U1335 (N_1335,N_605,N_553);
nor U1336 (N_1336,N_530,N_960);
nand U1337 (N_1337,N_638,N_652);
xor U1338 (N_1338,N_856,N_753);
or U1339 (N_1339,N_713,N_751);
and U1340 (N_1340,N_909,N_939);
nand U1341 (N_1341,N_960,N_941);
or U1342 (N_1342,N_787,N_687);
and U1343 (N_1343,N_508,N_575);
nor U1344 (N_1344,N_777,N_598);
nor U1345 (N_1345,N_788,N_549);
nor U1346 (N_1346,N_693,N_592);
or U1347 (N_1347,N_731,N_911);
nor U1348 (N_1348,N_587,N_751);
xnor U1349 (N_1349,N_930,N_866);
nor U1350 (N_1350,N_902,N_985);
or U1351 (N_1351,N_863,N_625);
nand U1352 (N_1352,N_972,N_865);
nor U1353 (N_1353,N_622,N_922);
and U1354 (N_1354,N_995,N_696);
and U1355 (N_1355,N_925,N_738);
xor U1356 (N_1356,N_973,N_695);
or U1357 (N_1357,N_520,N_928);
nor U1358 (N_1358,N_635,N_659);
and U1359 (N_1359,N_728,N_732);
or U1360 (N_1360,N_663,N_957);
nor U1361 (N_1361,N_923,N_884);
nand U1362 (N_1362,N_817,N_750);
nand U1363 (N_1363,N_503,N_523);
and U1364 (N_1364,N_779,N_928);
nor U1365 (N_1365,N_855,N_787);
nand U1366 (N_1366,N_667,N_790);
and U1367 (N_1367,N_852,N_525);
and U1368 (N_1368,N_838,N_621);
and U1369 (N_1369,N_601,N_593);
or U1370 (N_1370,N_601,N_999);
and U1371 (N_1371,N_522,N_796);
nor U1372 (N_1372,N_504,N_878);
nor U1373 (N_1373,N_903,N_853);
and U1374 (N_1374,N_801,N_761);
and U1375 (N_1375,N_645,N_977);
or U1376 (N_1376,N_955,N_771);
or U1377 (N_1377,N_640,N_543);
or U1378 (N_1378,N_690,N_817);
or U1379 (N_1379,N_836,N_881);
nor U1380 (N_1380,N_861,N_747);
or U1381 (N_1381,N_537,N_977);
and U1382 (N_1382,N_604,N_557);
nand U1383 (N_1383,N_663,N_940);
xnor U1384 (N_1384,N_612,N_626);
and U1385 (N_1385,N_992,N_835);
and U1386 (N_1386,N_873,N_812);
nand U1387 (N_1387,N_591,N_967);
nor U1388 (N_1388,N_963,N_700);
nor U1389 (N_1389,N_766,N_770);
nor U1390 (N_1390,N_893,N_717);
or U1391 (N_1391,N_883,N_787);
nor U1392 (N_1392,N_533,N_871);
and U1393 (N_1393,N_510,N_846);
nand U1394 (N_1394,N_930,N_745);
nor U1395 (N_1395,N_679,N_551);
nand U1396 (N_1396,N_885,N_691);
nand U1397 (N_1397,N_948,N_818);
nand U1398 (N_1398,N_793,N_504);
and U1399 (N_1399,N_889,N_613);
nor U1400 (N_1400,N_638,N_988);
and U1401 (N_1401,N_732,N_778);
nand U1402 (N_1402,N_763,N_587);
nor U1403 (N_1403,N_873,N_511);
nor U1404 (N_1404,N_509,N_560);
nand U1405 (N_1405,N_678,N_655);
or U1406 (N_1406,N_741,N_955);
or U1407 (N_1407,N_782,N_855);
and U1408 (N_1408,N_632,N_565);
nor U1409 (N_1409,N_921,N_631);
or U1410 (N_1410,N_782,N_808);
and U1411 (N_1411,N_757,N_784);
nand U1412 (N_1412,N_559,N_718);
nand U1413 (N_1413,N_724,N_780);
or U1414 (N_1414,N_812,N_532);
nand U1415 (N_1415,N_643,N_657);
nor U1416 (N_1416,N_919,N_657);
or U1417 (N_1417,N_897,N_624);
and U1418 (N_1418,N_767,N_712);
nor U1419 (N_1419,N_842,N_572);
nand U1420 (N_1420,N_624,N_661);
nand U1421 (N_1421,N_518,N_968);
or U1422 (N_1422,N_553,N_656);
or U1423 (N_1423,N_768,N_910);
and U1424 (N_1424,N_562,N_895);
nor U1425 (N_1425,N_906,N_921);
or U1426 (N_1426,N_842,N_996);
nor U1427 (N_1427,N_862,N_534);
xor U1428 (N_1428,N_617,N_779);
nor U1429 (N_1429,N_730,N_584);
or U1430 (N_1430,N_624,N_765);
and U1431 (N_1431,N_801,N_740);
or U1432 (N_1432,N_840,N_802);
nand U1433 (N_1433,N_546,N_607);
or U1434 (N_1434,N_608,N_729);
and U1435 (N_1435,N_781,N_886);
xnor U1436 (N_1436,N_971,N_771);
and U1437 (N_1437,N_755,N_860);
and U1438 (N_1438,N_649,N_638);
nand U1439 (N_1439,N_662,N_545);
nor U1440 (N_1440,N_549,N_775);
nor U1441 (N_1441,N_760,N_678);
nor U1442 (N_1442,N_742,N_602);
nor U1443 (N_1443,N_951,N_684);
or U1444 (N_1444,N_878,N_645);
xnor U1445 (N_1445,N_960,N_933);
nand U1446 (N_1446,N_791,N_684);
and U1447 (N_1447,N_577,N_795);
and U1448 (N_1448,N_691,N_653);
and U1449 (N_1449,N_857,N_733);
nor U1450 (N_1450,N_515,N_519);
xor U1451 (N_1451,N_583,N_975);
and U1452 (N_1452,N_813,N_954);
and U1453 (N_1453,N_842,N_888);
or U1454 (N_1454,N_839,N_873);
nor U1455 (N_1455,N_768,N_816);
and U1456 (N_1456,N_521,N_845);
or U1457 (N_1457,N_560,N_866);
and U1458 (N_1458,N_506,N_878);
nor U1459 (N_1459,N_735,N_510);
nand U1460 (N_1460,N_823,N_731);
or U1461 (N_1461,N_541,N_698);
and U1462 (N_1462,N_542,N_614);
or U1463 (N_1463,N_529,N_673);
nor U1464 (N_1464,N_903,N_513);
nand U1465 (N_1465,N_557,N_967);
or U1466 (N_1466,N_993,N_755);
nor U1467 (N_1467,N_769,N_927);
or U1468 (N_1468,N_603,N_952);
or U1469 (N_1469,N_769,N_873);
xor U1470 (N_1470,N_500,N_549);
or U1471 (N_1471,N_609,N_542);
xnor U1472 (N_1472,N_900,N_897);
nand U1473 (N_1473,N_670,N_822);
and U1474 (N_1474,N_582,N_572);
and U1475 (N_1475,N_883,N_860);
nand U1476 (N_1476,N_705,N_811);
xor U1477 (N_1477,N_839,N_518);
or U1478 (N_1478,N_705,N_849);
and U1479 (N_1479,N_824,N_635);
or U1480 (N_1480,N_740,N_718);
nor U1481 (N_1481,N_802,N_777);
nand U1482 (N_1482,N_740,N_705);
nor U1483 (N_1483,N_881,N_951);
nor U1484 (N_1484,N_685,N_896);
and U1485 (N_1485,N_551,N_742);
nand U1486 (N_1486,N_940,N_890);
nand U1487 (N_1487,N_836,N_729);
or U1488 (N_1488,N_848,N_808);
xor U1489 (N_1489,N_818,N_528);
or U1490 (N_1490,N_953,N_621);
and U1491 (N_1491,N_707,N_579);
and U1492 (N_1492,N_558,N_534);
or U1493 (N_1493,N_919,N_624);
and U1494 (N_1494,N_654,N_547);
or U1495 (N_1495,N_637,N_584);
or U1496 (N_1496,N_726,N_523);
nor U1497 (N_1497,N_746,N_664);
or U1498 (N_1498,N_726,N_849);
and U1499 (N_1499,N_658,N_625);
nand U1500 (N_1500,N_1165,N_1097);
or U1501 (N_1501,N_1273,N_1434);
or U1502 (N_1502,N_1267,N_1085);
nor U1503 (N_1503,N_1463,N_1124);
or U1504 (N_1504,N_1010,N_1299);
nand U1505 (N_1505,N_1318,N_1018);
nor U1506 (N_1506,N_1412,N_1208);
nand U1507 (N_1507,N_1421,N_1429);
nor U1508 (N_1508,N_1139,N_1013);
or U1509 (N_1509,N_1037,N_1190);
and U1510 (N_1510,N_1136,N_1140);
nand U1511 (N_1511,N_1402,N_1220);
nor U1512 (N_1512,N_1333,N_1035);
xor U1513 (N_1513,N_1368,N_1340);
or U1514 (N_1514,N_1493,N_1057);
nand U1515 (N_1515,N_1450,N_1388);
or U1516 (N_1516,N_1383,N_1455);
nor U1517 (N_1517,N_1117,N_1189);
nor U1518 (N_1518,N_1486,N_1128);
nor U1519 (N_1519,N_1174,N_1436);
nor U1520 (N_1520,N_1034,N_1329);
nand U1521 (N_1521,N_1243,N_1497);
nor U1522 (N_1522,N_1049,N_1047);
and U1523 (N_1523,N_1354,N_1355);
and U1524 (N_1524,N_1498,N_1431);
and U1525 (N_1525,N_1361,N_1363);
nand U1526 (N_1526,N_1286,N_1473);
or U1527 (N_1527,N_1437,N_1116);
or U1528 (N_1528,N_1425,N_1283);
nand U1529 (N_1529,N_1384,N_1126);
nor U1530 (N_1530,N_1108,N_1099);
or U1531 (N_1531,N_1216,N_1335);
nand U1532 (N_1532,N_1079,N_1033);
and U1533 (N_1533,N_1039,N_1083);
or U1534 (N_1534,N_1274,N_1161);
nor U1535 (N_1535,N_1198,N_1449);
nand U1536 (N_1536,N_1432,N_1023);
nand U1537 (N_1537,N_1435,N_1214);
nand U1538 (N_1538,N_1258,N_1186);
or U1539 (N_1539,N_1297,N_1137);
nor U1540 (N_1540,N_1387,N_1166);
and U1541 (N_1541,N_1400,N_1492);
or U1542 (N_1542,N_1251,N_1257);
and U1543 (N_1543,N_1032,N_1211);
and U1544 (N_1544,N_1285,N_1364);
and U1545 (N_1545,N_1055,N_1375);
or U1546 (N_1546,N_1464,N_1417);
nand U1547 (N_1547,N_1081,N_1224);
nor U1548 (N_1548,N_1115,N_1433);
or U1549 (N_1549,N_1247,N_1427);
nor U1550 (N_1550,N_1048,N_1359);
and U1551 (N_1551,N_1022,N_1228);
and U1552 (N_1552,N_1045,N_1327);
nor U1553 (N_1553,N_1011,N_1462);
and U1554 (N_1554,N_1014,N_1145);
and U1555 (N_1555,N_1328,N_1192);
nor U1556 (N_1556,N_1279,N_1056);
nand U1557 (N_1557,N_1106,N_1210);
nor U1558 (N_1558,N_1181,N_1317);
or U1559 (N_1559,N_1233,N_1159);
nand U1560 (N_1560,N_1397,N_1331);
and U1561 (N_1561,N_1238,N_1446);
nand U1562 (N_1562,N_1236,N_1094);
and U1563 (N_1563,N_1336,N_1206);
and U1564 (N_1564,N_1133,N_1483);
nor U1565 (N_1565,N_1420,N_1272);
nor U1566 (N_1566,N_1202,N_1180);
and U1567 (N_1567,N_1444,N_1118);
or U1568 (N_1568,N_1360,N_1231);
nand U1569 (N_1569,N_1242,N_1125);
and U1570 (N_1570,N_1287,N_1104);
nand U1571 (N_1571,N_1095,N_1170);
nor U1572 (N_1572,N_1271,N_1030);
or U1573 (N_1573,N_1374,N_1203);
nand U1574 (N_1574,N_1069,N_1093);
and U1575 (N_1575,N_1051,N_1027);
nand U1576 (N_1576,N_1149,N_1239);
nor U1577 (N_1577,N_1164,N_1175);
nor U1578 (N_1578,N_1160,N_1385);
and U1579 (N_1579,N_1487,N_1135);
nand U1580 (N_1580,N_1284,N_1304);
or U1581 (N_1581,N_1101,N_1007);
or U1582 (N_1582,N_1038,N_1046);
nand U1583 (N_1583,N_1332,N_1292);
or U1584 (N_1584,N_1087,N_1422);
nor U1585 (N_1585,N_1182,N_1004);
nor U1586 (N_1586,N_1062,N_1112);
nand U1587 (N_1587,N_1440,N_1103);
nand U1588 (N_1588,N_1218,N_1254);
nor U1589 (N_1589,N_1148,N_1219);
or U1590 (N_1590,N_1445,N_1499);
nor U1591 (N_1591,N_1119,N_1142);
and U1592 (N_1592,N_1157,N_1343);
nand U1593 (N_1593,N_1396,N_1373);
or U1594 (N_1594,N_1303,N_1330);
or U1595 (N_1595,N_1456,N_1401);
nand U1596 (N_1596,N_1480,N_1054);
and U1597 (N_1597,N_1114,N_1342);
xor U1598 (N_1598,N_1019,N_1471);
or U1599 (N_1599,N_1052,N_1447);
or U1600 (N_1600,N_1347,N_1266);
nor U1601 (N_1601,N_1452,N_1470);
nor U1602 (N_1602,N_1212,N_1351);
nand U1603 (N_1603,N_1026,N_1172);
xor U1604 (N_1604,N_1003,N_1248);
and U1605 (N_1605,N_1201,N_1454);
or U1606 (N_1606,N_1300,N_1409);
nand U1607 (N_1607,N_1098,N_1352);
and U1608 (N_1608,N_1415,N_1076);
xnor U1609 (N_1609,N_1393,N_1169);
nand U1610 (N_1610,N_1153,N_1015);
nor U1611 (N_1611,N_1316,N_1215);
nand U1612 (N_1612,N_1080,N_1065);
nand U1613 (N_1613,N_1372,N_1308);
and U1614 (N_1614,N_1105,N_1000);
nand U1615 (N_1615,N_1282,N_1245);
nor U1616 (N_1616,N_1102,N_1323);
xor U1617 (N_1617,N_1200,N_1301);
and U1618 (N_1618,N_1107,N_1269);
and U1619 (N_1619,N_1339,N_1423);
or U1620 (N_1620,N_1078,N_1349);
nand U1621 (N_1621,N_1240,N_1158);
or U1622 (N_1622,N_1197,N_1036);
nor U1623 (N_1623,N_1042,N_1461);
nor U1624 (N_1624,N_1146,N_1143);
and U1625 (N_1625,N_1195,N_1221);
nand U1626 (N_1626,N_1187,N_1082);
nor U1627 (N_1627,N_1307,N_1185);
or U1628 (N_1628,N_1399,N_1468);
nor U1629 (N_1629,N_1264,N_1009);
nor U1630 (N_1630,N_1322,N_1070);
and U1631 (N_1631,N_1320,N_1068);
and U1632 (N_1632,N_1475,N_1398);
or U1633 (N_1633,N_1426,N_1008);
or U1634 (N_1634,N_1371,N_1110);
nor U1635 (N_1635,N_1382,N_1150);
nand U1636 (N_1636,N_1326,N_1167);
nor U1637 (N_1637,N_1067,N_1088);
and U1638 (N_1638,N_1138,N_1465);
and U1639 (N_1639,N_1021,N_1122);
nor U1640 (N_1640,N_1319,N_1179);
nor U1641 (N_1641,N_1089,N_1386);
nor U1642 (N_1642,N_1071,N_1050);
nor U1643 (N_1643,N_1494,N_1005);
or U1644 (N_1644,N_1025,N_1295);
nand U1645 (N_1645,N_1152,N_1263);
and U1646 (N_1646,N_1176,N_1418);
or U1647 (N_1647,N_1155,N_1411);
or U1648 (N_1648,N_1002,N_1369);
nor U1649 (N_1649,N_1281,N_1129);
nor U1650 (N_1650,N_1296,N_1439);
nand U1651 (N_1651,N_1260,N_1496);
nand U1652 (N_1652,N_1353,N_1249);
nor U1653 (N_1653,N_1194,N_1168);
nor U1654 (N_1654,N_1490,N_1223);
nand U1655 (N_1655,N_1325,N_1261);
nand U1656 (N_1656,N_1276,N_1130);
nand U1657 (N_1657,N_1262,N_1315);
nor U1658 (N_1658,N_1121,N_1134);
nor U1659 (N_1659,N_1424,N_1495);
nor U1660 (N_1660,N_1204,N_1268);
and U1661 (N_1661,N_1059,N_1313);
nand U1662 (N_1662,N_1466,N_1484);
and U1663 (N_1663,N_1229,N_1100);
and U1664 (N_1664,N_1491,N_1278);
and U1665 (N_1665,N_1184,N_1040);
nor U1666 (N_1666,N_1171,N_1291);
nor U1667 (N_1667,N_1380,N_1123);
nand U1668 (N_1668,N_1096,N_1162);
nand U1669 (N_1669,N_1311,N_1041);
and U1670 (N_1670,N_1147,N_1132);
or U1671 (N_1671,N_1232,N_1213);
and U1672 (N_1672,N_1028,N_1092);
nand U1673 (N_1673,N_1044,N_1154);
or U1674 (N_1674,N_1031,N_1404);
nand U1675 (N_1675,N_1459,N_1151);
nor U1676 (N_1676,N_1277,N_1256);
nor U1677 (N_1677,N_1430,N_1362);
and U1678 (N_1678,N_1334,N_1479);
nor U1679 (N_1679,N_1217,N_1091);
or U1680 (N_1680,N_1414,N_1227);
or U1681 (N_1681,N_1252,N_1001);
and U1682 (N_1682,N_1016,N_1416);
nand U1683 (N_1683,N_1390,N_1207);
xnor U1684 (N_1684,N_1405,N_1310);
nor U1685 (N_1685,N_1265,N_1127);
or U1686 (N_1686,N_1073,N_1294);
nand U1687 (N_1687,N_1156,N_1410);
and U1688 (N_1688,N_1120,N_1131);
or U1689 (N_1689,N_1199,N_1477);
nand U1690 (N_1690,N_1395,N_1205);
nor U1691 (N_1691,N_1246,N_1275);
and U1692 (N_1692,N_1141,N_1244);
nor U1693 (N_1693,N_1442,N_1357);
nor U1694 (N_1694,N_1458,N_1163);
nand U1695 (N_1695,N_1481,N_1259);
and U1696 (N_1696,N_1064,N_1012);
or U1697 (N_1697,N_1366,N_1066);
or U1698 (N_1698,N_1478,N_1255);
nor U1699 (N_1699,N_1109,N_1392);
nand U1700 (N_1700,N_1072,N_1306);
and U1701 (N_1701,N_1293,N_1467);
or U1702 (N_1702,N_1309,N_1241);
and U1703 (N_1703,N_1428,N_1314);
nand U1704 (N_1704,N_1337,N_1253);
nor U1705 (N_1705,N_1234,N_1365);
nor U1706 (N_1706,N_1173,N_1188);
nand U1707 (N_1707,N_1485,N_1408);
nor U1708 (N_1708,N_1489,N_1376);
and U1709 (N_1709,N_1348,N_1075);
and U1710 (N_1710,N_1413,N_1457);
or U1711 (N_1711,N_1177,N_1191);
nand U1712 (N_1712,N_1469,N_1472);
and U1713 (N_1713,N_1448,N_1389);
and U1714 (N_1714,N_1391,N_1438);
nor U1715 (N_1715,N_1288,N_1084);
and U1716 (N_1716,N_1043,N_1367);
or U1717 (N_1717,N_1358,N_1406);
or U1718 (N_1718,N_1074,N_1237);
nand U1719 (N_1719,N_1222,N_1235);
nor U1720 (N_1720,N_1270,N_1476);
nor U1721 (N_1721,N_1058,N_1419);
and U1722 (N_1722,N_1289,N_1061);
nor U1723 (N_1723,N_1113,N_1443);
or U1724 (N_1724,N_1345,N_1090);
or U1725 (N_1725,N_1356,N_1209);
or U1726 (N_1726,N_1379,N_1341);
nor U1727 (N_1727,N_1063,N_1302);
nand U1728 (N_1728,N_1290,N_1381);
nand U1729 (N_1729,N_1346,N_1451);
nand U1730 (N_1730,N_1298,N_1488);
nand U1731 (N_1731,N_1029,N_1350);
or U1732 (N_1732,N_1111,N_1453);
and U1733 (N_1733,N_1441,N_1193);
nand U1734 (N_1734,N_1053,N_1378);
nor U1735 (N_1735,N_1060,N_1460);
and U1736 (N_1736,N_1344,N_1225);
or U1737 (N_1737,N_1338,N_1312);
nor U1738 (N_1738,N_1324,N_1086);
and U1739 (N_1739,N_1377,N_1250);
nor U1740 (N_1740,N_1474,N_1280);
nand U1741 (N_1741,N_1394,N_1020);
nand U1742 (N_1742,N_1305,N_1144);
nor U1743 (N_1743,N_1017,N_1403);
nor U1744 (N_1744,N_1226,N_1407);
nand U1745 (N_1745,N_1196,N_1183);
nand U1746 (N_1746,N_1178,N_1321);
and U1747 (N_1747,N_1230,N_1077);
or U1748 (N_1748,N_1482,N_1370);
nor U1749 (N_1749,N_1024,N_1006);
nand U1750 (N_1750,N_1070,N_1050);
or U1751 (N_1751,N_1264,N_1439);
nand U1752 (N_1752,N_1428,N_1384);
nand U1753 (N_1753,N_1341,N_1351);
or U1754 (N_1754,N_1190,N_1035);
and U1755 (N_1755,N_1045,N_1498);
nand U1756 (N_1756,N_1241,N_1448);
nor U1757 (N_1757,N_1079,N_1212);
nand U1758 (N_1758,N_1089,N_1082);
and U1759 (N_1759,N_1291,N_1147);
and U1760 (N_1760,N_1317,N_1047);
or U1761 (N_1761,N_1377,N_1150);
nand U1762 (N_1762,N_1365,N_1364);
or U1763 (N_1763,N_1291,N_1285);
xnor U1764 (N_1764,N_1028,N_1295);
nand U1765 (N_1765,N_1179,N_1180);
nor U1766 (N_1766,N_1002,N_1477);
nand U1767 (N_1767,N_1096,N_1178);
nor U1768 (N_1768,N_1202,N_1048);
and U1769 (N_1769,N_1174,N_1035);
nand U1770 (N_1770,N_1420,N_1245);
or U1771 (N_1771,N_1299,N_1078);
nor U1772 (N_1772,N_1098,N_1388);
or U1773 (N_1773,N_1267,N_1010);
or U1774 (N_1774,N_1328,N_1375);
nand U1775 (N_1775,N_1141,N_1499);
nand U1776 (N_1776,N_1197,N_1051);
and U1777 (N_1777,N_1118,N_1220);
nand U1778 (N_1778,N_1065,N_1376);
or U1779 (N_1779,N_1125,N_1109);
and U1780 (N_1780,N_1458,N_1229);
nand U1781 (N_1781,N_1133,N_1060);
or U1782 (N_1782,N_1397,N_1222);
and U1783 (N_1783,N_1107,N_1472);
nand U1784 (N_1784,N_1118,N_1097);
or U1785 (N_1785,N_1011,N_1171);
nand U1786 (N_1786,N_1089,N_1219);
and U1787 (N_1787,N_1483,N_1041);
and U1788 (N_1788,N_1159,N_1310);
nand U1789 (N_1789,N_1069,N_1237);
nor U1790 (N_1790,N_1252,N_1394);
or U1791 (N_1791,N_1120,N_1191);
or U1792 (N_1792,N_1204,N_1461);
nor U1793 (N_1793,N_1055,N_1098);
or U1794 (N_1794,N_1011,N_1166);
nand U1795 (N_1795,N_1155,N_1102);
and U1796 (N_1796,N_1267,N_1452);
nand U1797 (N_1797,N_1266,N_1019);
and U1798 (N_1798,N_1258,N_1078);
nand U1799 (N_1799,N_1121,N_1102);
nand U1800 (N_1800,N_1447,N_1261);
or U1801 (N_1801,N_1363,N_1164);
or U1802 (N_1802,N_1195,N_1136);
nand U1803 (N_1803,N_1157,N_1158);
nor U1804 (N_1804,N_1135,N_1209);
or U1805 (N_1805,N_1219,N_1154);
nand U1806 (N_1806,N_1019,N_1151);
and U1807 (N_1807,N_1474,N_1464);
nor U1808 (N_1808,N_1247,N_1056);
xnor U1809 (N_1809,N_1468,N_1137);
nor U1810 (N_1810,N_1001,N_1213);
nand U1811 (N_1811,N_1130,N_1039);
nor U1812 (N_1812,N_1053,N_1401);
or U1813 (N_1813,N_1373,N_1494);
and U1814 (N_1814,N_1474,N_1194);
and U1815 (N_1815,N_1294,N_1110);
nand U1816 (N_1816,N_1332,N_1165);
and U1817 (N_1817,N_1372,N_1316);
nor U1818 (N_1818,N_1450,N_1036);
and U1819 (N_1819,N_1456,N_1486);
and U1820 (N_1820,N_1330,N_1152);
xnor U1821 (N_1821,N_1236,N_1285);
and U1822 (N_1822,N_1001,N_1130);
and U1823 (N_1823,N_1276,N_1469);
and U1824 (N_1824,N_1483,N_1247);
nor U1825 (N_1825,N_1347,N_1144);
or U1826 (N_1826,N_1147,N_1373);
nand U1827 (N_1827,N_1296,N_1056);
and U1828 (N_1828,N_1289,N_1087);
or U1829 (N_1829,N_1466,N_1057);
nand U1830 (N_1830,N_1152,N_1359);
and U1831 (N_1831,N_1328,N_1080);
nor U1832 (N_1832,N_1335,N_1179);
xor U1833 (N_1833,N_1012,N_1297);
or U1834 (N_1834,N_1350,N_1267);
and U1835 (N_1835,N_1415,N_1413);
nor U1836 (N_1836,N_1167,N_1308);
nand U1837 (N_1837,N_1218,N_1459);
and U1838 (N_1838,N_1398,N_1026);
nand U1839 (N_1839,N_1474,N_1420);
and U1840 (N_1840,N_1400,N_1070);
and U1841 (N_1841,N_1174,N_1319);
nor U1842 (N_1842,N_1040,N_1474);
nor U1843 (N_1843,N_1154,N_1307);
or U1844 (N_1844,N_1364,N_1315);
xor U1845 (N_1845,N_1286,N_1495);
nand U1846 (N_1846,N_1107,N_1135);
nor U1847 (N_1847,N_1447,N_1053);
nor U1848 (N_1848,N_1033,N_1403);
or U1849 (N_1849,N_1174,N_1229);
nand U1850 (N_1850,N_1345,N_1343);
and U1851 (N_1851,N_1233,N_1093);
and U1852 (N_1852,N_1242,N_1494);
or U1853 (N_1853,N_1177,N_1065);
nor U1854 (N_1854,N_1306,N_1255);
nor U1855 (N_1855,N_1350,N_1409);
or U1856 (N_1856,N_1242,N_1410);
nor U1857 (N_1857,N_1239,N_1173);
nand U1858 (N_1858,N_1189,N_1324);
and U1859 (N_1859,N_1324,N_1282);
and U1860 (N_1860,N_1396,N_1269);
or U1861 (N_1861,N_1213,N_1465);
and U1862 (N_1862,N_1006,N_1384);
and U1863 (N_1863,N_1045,N_1013);
or U1864 (N_1864,N_1337,N_1144);
or U1865 (N_1865,N_1344,N_1424);
and U1866 (N_1866,N_1117,N_1084);
and U1867 (N_1867,N_1367,N_1362);
or U1868 (N_1868,N_1157,N_1474);
or U1869 (N_1869,N_1030,N_1100);
or U1870 (N_1870,N_1262,N_1309);
or U1871 (N_1871,N_1189,N_1020);
and U1872 (N_1872,N_1134,N_1451);
and U1873 (N_1873,N_1479,N_1167);
nand U1874 (N_1874,N_1255,N_1424);
nand U1875 (N_1875,N_1081,N_1478);
nand U1876 (N_1876,N_1034,N_1361);
nand U1877 (N_1877,N_1239,N_1339);
or U1878 (N_1878,N_1046,N_1366);
nor U1879 (N_1879,N_1377,N_1078);
or U1880 (N_1880,N_1375,N_1160);
and U1881 (N_1881,N_1035,N_1384);
nor U1882 (N_1882,N_1205,N_1372);
and U1883 (N_1883,N_1322,N_1392);
nand U1884 (N_1884,N_1071,N_1262);
or U1885 (N_1885,N_1375,N_1489);
or U1886 (N_1886,N_1027,N_1468);
nand U1887 (N_1887,N_1192,N_1211);
or U1888 (N_1888,N_1239,N_1288);
and U1889 (N_1889,N_1340,N_1170);
nor U1890 (N_1890,N_1387,N_1274);
nor U1891 (N_1891,N_1411,N_1312);
nand U1892 (N_1892,N_1256,N_1009);
nand U1893 (N_1893,N_1111,N_1038);
and U1894 (N_1894,N_1136,N_1062);
nor U1895 (N_1895,N_1128,N_1412);
and U1896 (N_1896,N_1006,N_1417);
nand U1897 (N_1897,N_1071,N_1077);
and U1898 (N_1898,N_1337,N_1400);
nand U1899 (N_1899,N_1025,N_1163);
nand U1900 (N_1900,N_1411,N_1224);
nand U1901 (N_1901,N_1143,N_1098);
and U1902 (N_1902,N_1141,N_1327);
and U1903 (N_1903,N_1462,N_1461);
nor U1904 (N_1904,N_1497,N_1019);
or U1905 (N_1905,N_1202,N_1263);
nor U1906 (N_1906,N_1402,N_1295);
nor U1907 (N_1907,N_1325,N_1246);
nor U1908 (N_1908,N_1058,N_1350);
and U1909 (N_1909,N_1028,N_1043);
or U1910 (N_1910,N_1304,N_1036);
nand U1911 (N_1911,N_1328,N_1041);
or U1912 (N_1912,N_1427,N_1325);
nand U1913 (N_1913,N_1017,N_1055);
or U1914 (N_1914,N_1172,N_1465);
or U1915 (N_1915,N_1032,N_1238);
nor U1916 (N_1916,N_1155,N_1097);
and U1917 (N_1917,N_1270,N_1117);
and U1918 (N_1918,N_1380,N_1235);
and U1919 (N_1919,N_1321,N_1423);
nor U1920 (N_1920,N_1155,N_1152);
nand U1921 (N_1921,N_1385,N_1401);
or U1922 (N_1922,N_1161,N_1054);
nor U1923 (N_1923,N_1441,N_1407);
and U1924 (N_1924,N_1023,N_1338);
and U1925 (N_1925,N_1034,N_1374);
nand U1926 (N_1926,N_1370,N_1219);
xnor U1927 (N_1927,N_1253,N_1043);
or U1928 (N_1928,N_1050,N_1369);
nand U1929 (N_1929,N_1324,N_1481);
nand U1930 (N_1930,N_1438,N_1383);
or U1931 (N_1931,N_1435,N_1260);
or U1932 (N_1932,N_1323,N_1307);
and U1933 (N_1933,N_1426,N_1136);
and U1934 (N_1934,N_1360,N_1274);
and U1935 (N_1935,N_1056,N_1438);
or U1936 (N_1936,N_1324,N_1152);
or U1937 (N_1937,N_1152,N_1223);
and U1938 (N_1938,N_1454,N_1262);
nand U1939 (N_1939,N_1307,N_1096);
and U1940 (N_1940,N_1247,N_1331);
and U1941 (N_1941,N_1072,N_1136);
nand U1942 (N_1942,N_1242,N_1019);
nor U1943 (N_1943,N_1370,N_1127);
nand U1944 (N_1944,N_1421,N_1183);
nor U1945 (N_1945,N_1051,N_1347);
nor U1946 (N_1946,N_1479,N_1352);
or U1947 (N_1947,N_1197,N_1174);
nor U1948 (N_1948,N_1137,N_1042);
nand U1949 (N_1949,N_1026,N_1210);
nor U1950 (N_1950,N_1114,N_1462);
nand U1951 (N_1951,N_1148,N_1013);
nand U1952 (N_1952,N_1449,N_1068);
nor U1953 (N_1953,N_1342,N_1277);
nand U1954 (N_1954,N_1158,N_1085);
nand U1955 (N_1955,N_1254,N_1183);
nand U1956 (N_1956,N_1281,N_1055);
or U1957 (N_1957,N_1013,N_1150);
nand U1958 (N_1958,N_1464,N_1357);
and U1959 (N_1959,N_1221,N_1337);
and U1960 (N_1960,N_1279,N_1369);
and U1961 (N_1961,N_1388,N_1474);
xnor U1962 (N_1962,N_1102,N_1488);
nand U1963 (N_1963,N_1214,N_1103);
nand U1964 (N_1964,N_1055,N_1407);
nand U1965 (N_1965,N_1377,N_1164);
nand U1966 (N_1966,N_1229,N_1258);
nand U1967 (N_1967,N_1304,N_1452);
and U1968 (N_1968,N_1463,N_1076);
or U1969 (N_1969,N_1133,N_1091);
nor U1970 (N_1970,N_1115,N_1020);
xnor U1971 (N_1971,N_1455,N_1208);
or U1972 (N_1972,N_1364,N_1064);
nor U1973 (N_1973,N_1419,N_1286);
nor U1974 (N_1974,N_1333,N_1401);
nor U1975 (N_1975,N_1000,N_1002);
and U1976 (N_1976,N_1027,N_1457);
nand U1977 (N_1977,N_1187,N_1110);
and U1978 (N_1978,N_1184,N_1402);
nand U1979 (N_1979,N_1385,N_1122);
and U1980 (N_1980,N_1207,N_1029);
or U1981 (N_1981,N_1015,N_1118);
nand U1982 (N_1982,N_1324,N_1355);
and U1983 (N_1983,N_1169,N_1154);
and U1984 (N_1984,N_1104,N_1478);
or U1985 (N_1985,N_1257,N_1252);
and U1986 (N_1986,N_1445,N_1039);
and U1987 (N_1987,N_1055,N_1332);
xor U1988 (N_1988,N_1135,N_1321);
and U1989 (N_1989,N_1107,N_1369);
nor U1990 (N_1990,N_1439,N_1210);
nand U1991 (N_1991,N_1354,N_1333);
or U1992 (N_1992,N_1483,N_1287);
or U1993 (N_1993,N_1323,N_1328);
nor U1994 (N_1994,N_1216,N_1051);
or U1995 (N_1995,N_1298,N_1036);
xnor U1996 (N_1996,N_1144,N_1042);
nor U1997 (N_1997,N_1410,N_1347);
nor U1998 (N_1998,N_1102,N_1340);
and U1999 (N_1999,N_1169,N_1262);
and U2000 (N_2000,N_1781,N_1942);
and U2001 (N_2001,N_1804,N_1827);
or U2002 (N_2002,N_1956,N_1696);
or U2003 (N_2003,N_1562,N_1673);
and U2004 (N_2004,N_1779,N_1637);
and U2005 (N_2005,N_1874,N_1866);
nand U2006 (N_2006,N_1701,N_1587);
nand U2007 (N_2007,N_1631,N_1854);
nor U2008 (N_2008,N_1726,N_1968);
or U2009 (N_2009,N_1853,N_1563);
nand U2010 (N_2010,N_1824,N_1740);
nand U2011 (N_2011,N_1775,N_1873);
nand U2012 (N_2012,N_1909,N_1992);
and U2013 (N_2013,N_1807,N_1962);
nor U2014 (N_2014,N_1518,N_1682);
nand U2015 (N_2015,N_1864,N_1925);
or U2016 (N_2016,N_1893,N_1744);
or U2017 (N_2017,N_1504,N_1555);
and U2018 (N_2018,N_1583,N_1738);
nand U2019 (N_2019,N_1887,N_1971);
and U2020 (N_2020,N_1612,N_1845);
and U2021 (N_2021,N_1839,N_1693);
nand U2022 (N_2022,N_1690,N_1922);
nor U2023 (N_2023,N_1525,N_1940);
nor U2024 (N_2024,N_1894,N_1783);
and U2025 (N_2025,N_1561,N_1559);
and U2026 (N_2026,N_1786,N_1952);
nor U2027 (N_2027,N_1819,N_1581);
or U2028 (N_2028,N_1769,N_1535);
xor U2029 (N_2029,N_1987,N_1538);
and U2030 (N_2030,N_1821,N_1611);
or U2031 (N_2031,N_1645,N_1772);
or U2032 (N_2032,N_1954,N_1735);
nand U2033 (N_2033,N_1536,N_1755);
or U2034 (N_2034,N_1569,N_1834);
and U2035 (N_2035,N_1960,N_1567);
and U2036 (N_2036,N_1731,N_1966);
or U2037 (N_2037,N_1680,N_1876);
nand U2038 (N_2038,N_1614,N_1549);
and U2039 (N_2039,N_1918,N_1815);
and U2040 (N_2040,N_1833,N_1941);
or U2041 (N_2041,N_1898,N_1544);
and U2042 (N_2042,N_1672,N_1566);
nor U2043 (N_2043,N_1698,N_1787);
nor U2044 (N_2044,N_1799,N_1702);
or U2045 (N_2045,N_1647,N_1610);
or U2046 (N_2046,N_1801,N_1832);
nor U2047 (N_2047,N_1802,N_1969);
nor U2048 (N_2048,N_1676,N_1595);
and U2049 (N_2049,N_1784,N_1655);
nand U2050 (N_2050,N_1985,N_1902);
nor U2051 (N_2051,N_1764,N_1939);
and U2052 (N_2052,N_1770,N_1812);
or U2053 (N_2053,N_1957,N_1677);
nand U2054 (N_2054,N_1529,N_1979);
nand U2055 (N_2055,N_1849,N_1511);
and U2056 (N_2056,N_1572,N_1554);
nor U2057 (N_2057,N_1712,N_1792);
and U2058 (N_2058,N_1661,N_1808);
nand U2059 (N_2059,N_1923,N_1919);
nand U2060 (N_2060,N_1917,N_1633);
and U2061 (N_2061,N_1644,N_1859);
nand U2062 (N_2062,N_1774,N_1888);
and U2063 (N_2063,N_1835,N_1601);
nor U2064 (N_2064,N_1656,N_1621);
and U2065 (N_2065,N_1692,N_1908);
or U2066 (N_2066,N_1506,N_1666);
nor U2067 (N_2067,N_1789,N_1658);
nor U2068 (N_2068,N_1705,N_1790);
or U2069 (N_2069,N_1773,N_1776);
nand U2070 (N_2070,N_1623,N_1648);
and U2071 (N_2071,N_1593,N_1616);
nor U2072 (N_2072,N_1896,N_1803);
or U2073 (N_2073,N_1700,N_1830);
xor U2074 (N_2074,N_1752,N_1542);
or U2075 (N_2075,N_1681,N_1951);
nand U2076 (N_2076,N_1540,N_1946);
and U2077 (N_2077,N_1732,N_1892);
and U2078 (N_2078,N_1885,N_1809);
nor U2079 (N_2079,N_1685,N_1704);
nor U2080 (N_2080,N_1708,N_1509);
and U2081 (N_2081,N_1910,N_1578);
nor U2082 (N_2082,N_1613,N_1534);
nand U2083 (N_2083,N_1972,N_1948);
or U2084 (N_2084,N_1615,N_1758);
or U2085 (N_2085,N_1724,N_1573);
nor U2086 (N_2086,N_1788,N_1862);
nand U2087 (N_2087,N_1643,N_1530);
and U2088 (N_2088,N_1521,N_1659);
and U2089 (N_2089,N_1930,N_1867);
nand U2090 (N_2090,N_1520,N_1608);
or U2091 (N_2091,N_1625,N_1991);
nand U2092 (N_2092,N_1999,N_1878);
nor U2093 (N_2093,N_1826,N_1868);
or U2094 (N_2094,N_1903,N_1975);
nand U2095 (N_2095,N_1565,N_1683);
and U2096 (N_2096,N_1844,N_1929);
and U2097 (N_2097,N_1905,N_1884);
or U2098 (N_2098,N_1765,N_1523);
nand U2099 (N_2099,N_1571,N_1590);
or U2100 (N_2100,N_1945,N_1539);
nor U2101 (N_2101,N_1852,N_1748);
nor U2102 (N_2102,N_1901,N_1718);
nand U2103 (N_2103,N_1543,N_1889);
and U2104 (N_2104,N_1635,N_1955);
and U2105 (N_2105,N_1932,N_1512);
nand U2106 (N_2106,N_1654,N_1639);
xor U2107 (N_2107,N_1517,N_1983);
nor U2108 (N_2108,N_1937,N_1707);
and U2109 (N_2109,N_1668,N_1660);
or U2110 (N_2110,N_1899,N_1519);
or U2111 (N_2111,N_1603,N_1545);
nand U2112 (N_2112,N_1716,N_1817);
nand U2113 (N_2113,N_1730,N_1736);
nor U2114 (N_2114,N_1747,N_1689);
nor U2115 (N_2115,N_1753,N_1657);
or U2116 (N_2116,N_1996,N_1665);
or U2117 (N_2117,N_1522,N_1618);
nand U2118 (N_2118,N_1632,N_1831);
or U2119 (N_2119,N_1914,N_1713);
nor U2120 (N_2120,N_1994,N_1630);
or U2121 (N_2121,N_1816,N_1594);
or U2122 (N_2122,N_1856,N_1880);
and U2123 (N_2123,N_1627,N_1727);
and U2124 (N_2124,N_1785,N_1754);
nand U2125 (N_2125,N_1751,N_1500);
and U2126 (N_2126,N_1588,N_1895);
or U2127 (N_2127,N_1911,N_1697);
and U2128 (N_2128,N_1508,N_1586);
or U2129 (N_2129,N_1861,N_1793);
nor U2130 (N_2130,N_1671,N_1725);
and U2131 (N_2131,N_1974,N_1592);
nand U2132 (N_2132,N_1503,N_1597);
nand U2133 (N_2133,N_1596,N_1794);
or U2134 (N_2134,N_1875,N_1715);
nor U2135 (N_2135,N_1970,N_1650);
nand U2136 (N_2136,N_1546,N_1737);
nor U2137 (N_2137,N_1527,N_1978);
and U2138 (N_2138,N_1977,N_1628);
nor U2139 (N_2139,N_1963,N_1965);
nor U2140 (N_2140,N_1646,N_1629);
nand U2141 (N_2141,N_1865,N_1729);
and U2142 (N_2142,N_1580,N_1904);
or U2143 (N_2143,N_1771,N_1938);
and U2144 (N_2144,N_1843,N_1762);
xor U2145 (N_2145,N_1912,N_1686);
and U2146 (N_2146,N_1515,N_1501);
nor U2147 (N_2147,N_1582,N_1589);
or U2148 (N_2148,N_1695,N_1591);
or U2149 (N_2149,N_1720,N_1797);
or U2150 (N_2150,N_1768,N_1624);
nor U2151 (N_2151,N_1675,N_1528);
xor U2152 (N_2152,N_1881,N_1921);
nor U2153 (N_2153,N_1883,N_1600);
and U2154 (N_2154,N_1850,N_1570);
nor U2155 (N_2155,N_1617,N_1800);
nor U2156 (N_2156,N_1741,N_1507);
and U2157 (N_2157,N_1961,N_1745);
nor U2158 (N_2158,N_1669,N_1778);
nand U2159 (N_2159,N_1688,N_1798);
and U2160 (N_2160,N_1717,N_1619);
xnor U2161 (N_2161,N_1560,N_1620);
nand U2162 (N_2162,N_1879,N_1605);
nor U2163 (N_2163,N_1626,N_1848);
nand U2164 (N_2164,N_1513,N_1759);
nor U2165 (N_2165,N_1743,N_1777);
nand U2166 (N_2166,N_1915,N_1557);
and U2167 (N_2167,N_1548,N_1579);
and U2168 (N_2168,N_1851,N_1944);
nor U2169 (N_2169,N_1761,N_1552);
nand U2170 (N_2170,N_1926,N_1913);
and U2171 (N_2171,N_1767,N_1606);
or U2172 (N_2172,N_1652,N_1607);
nor U2173 (N_2173,N_1739,N_1906);
nor U2174 (N_2174,N_1953,N_1634);
nor U2175 (N_2175,N_1728,N_1553);
or U2176 (N_2176,N_1870,N_1664);
or U2177 (N_2177,N_1653,N_1841);
and U2178 (N_2178,N_1810,N_1679);
and U2179 (N_2179,N_1995,N_1531);
or U2180 (N_2180,N_1746,N_1721);
or U2181 (N_2181,N_1733,N_1699);
and U2182 (N_2182,N_1763,N_1986);
xor U2183 (N_2183,N_1836,N_1818);
and U2184 (N_2184,N_1907,N_1860);
nand U2185 (N_2185,N_1928,N_1526);
nor U2186 (N_2186,N_1541,N_1976);
or U2187 (N_2187,N_1936,N_1766);
nand U2188 (N_2188,N_1709,N_1890);
xor U2189 (N_2189,N_1882,N_1998);
and U2190 (N_2190,N_1749,N_1760);
and U2191 (N_2191,N_1814,N_1828);
nor U2192 (N_2192,N_1927,N_1916);
nor U2193 (N_2193,N_1838,N_1574);
nand U2194 (N_2194,N_1959,N_1719);
nand U2195 (N_2195,N_1967,N_1703);
and U2196 (N_2196,N_1934,N_1950);
or U2197 (N_2197,N_1877,N_1842);
and U2198 (N_2198,N_1577,N_1750);
nand U2199 (N_2199,N_1510,N_1829);
or U2200 (N_2200,N_1641,N_1537);
nand U2201 (N_2201,N_1687,N_1663);
nand U2202 (N_2202,N_1640,N_1547);
and U2203 (N_2203,N_1694,N_1638);
or U2204 (N_2204,N_1516,N_1990);
and U2205 (N_2205,N_1949,N_1780);
or U2206 (N_2206,N_1920,N_1723);
nor U2207 (N_2207,N_1811,N_1872);
nand U2208 (N_2208,N_1795,N_1609);
nand U2209 (N_2209,N_1678,N_1599);
nor U2210 (N_2210,N_1989,N_1791);
or U2211 (N_2211,N_1900,N_1622);
nor U2212 (N_2212,N_1891,N_1980);
nand U2213 (N_2213,N_1931,N_1869);
nand U2214 (N_2214,N_1598,N_1973);
or U2215 (N_2215,N_1584,N_1550);
and U2216 (N_2216,N_1822,N_1651);
and U2217 (N_2217,N_1636,N_1855);
or U2218 (N_2218,N_1710,N_1984);
nand U2219 (N_2219,N_1568,N_1806);
or U2220 (N_2220,N_1602,N_1782);
and U2221 (N_2221,N_1670,N_1886);
nand U2222 (N_2222,N_1947,N_1757);
or U2223 (N_2223,N_1714,N_1564);
or U2224 (N_2224,N_1711,N_1823);
nand U2225 (N_2225,N_1691,N_1649);
nor U2226 (N_2226,N_1840,N_1863);
nand U2227 (N_2227,N_1988,N_1667);
nand U2228 (N_2228,N_1604,N_1533);
nand U2229 (N_2229,N_1684,N_1820);
or U2230 (N_2230,N_1993,N_1742);
or U2231 (N_2231,N_1924,N_1997);
and U2232 (N_2232,N_1813,N_1662);
nor U2233 (N_2233,N_1576,N_1825);
and U2234 (N_2234,N_1805,N_1964);
nor U2235 (N_2235,N_1756,N_1642);
or U2236 (N_2236,N_1722,N_1846);
nand U2237 (N_2237,N_1858,N_1674);
or U2238 (N_2238,N_1982,N_1585);
nor U2239 (N_2239,N_1556,N_1706);
nor U2240 (N_2240,N_1734,N_1935);
and U2241 (N_2241,N_1558,N_1857);
nor U2242 (N_2242,N_1505,N_1532);
nor U2243 (N_2243,N_1958,N_1933);
nand U2244 (N_2244,N_1575,N_1943);
and U2245 (N_2245,N_1871,N_1796);
nand U2246 (N_2246,N_1897,N_1502);
or U2247 (N_2247,N_1981,N_1551);
or U2248 (N_2248,N_1524,N_1837);
or U2249 (N_2249,N_1847,N_1514);
nand U2250 (N_2250,N_1981,N_1999);
nand U2251 (N_2251,N_1905,N_1780);
nor U2252 (N_2252,N_1688,N_1910);
and U2253 (N_2253,N_1640,N_1656);
nand U2254 (N_2254,N_1782,N_1524);
and U2255 (N_2255,N_1645,N_1946);
nand U2256 (N_2256,N_1874,N_1525);
nand U2257 (N_2257,N_1934,N_1886);
nand U2258 (N_2258,N_1920,N_1793);
and U2259 (N_2259,N_1905,N_1544);
nand U2260 (N_2260,N_1705,N_1769);
and U2261 (N_2261,N_1516,N_1972);
or U2262 (N_2262,N_1530,N_1668);
nand U2263 (N_2263,N_1809,N_1790);
or U2264 (N_2264,N_1999,N_1948);
nand U2265 (N_2265,N_1873,N_1500);
or U2266 (N_2266,N_1871,N_1968);
or U2267 (N_2267,N_1578,N_1630);
and U2268 (N_2268,N_1748,N_1978);
or U2269 (N_2269,N_1797,N_1746);
and U2270 (N_2270,N_1817,N_1741);
nor U2271 (N_2271,N_1985,N_1570);
nor U2272 (N_2272,N_1621,N_1663);
and U2273 (N_2273,N_1726,N_1639);
and U2274 (N_2274,N_1692,N_1956);
or U2275 (N_2275,N_1849,N_1666);
or U2276 (N_2276,N_1649,N_1534);
and U2277 (N_2277,N_1669,N_1986);
or U2278 (N_2278,N_1761,N_1896);
nand U2279 (N_2279,N_1567,N_1652);
nor U2280 (N_2280,N_1602,N_1965);
nand U2281 (N_2281,N_1843,N_1917);
nand U2282 (N_2282,N_1736,N_1792);
nand U2283 (N_2283,N_1800,N_1747);
nand U2284 (N_2284,N_1836,N_1932);
and U2285 (N_2285,N_1662,N_1909);
and U2286 (N_2286,N_1817,N_1810);
and U2287 (N_2287,N_1717,N_1553);
nand U2288 (N_2288,N_1783,N_1609);
or U2289 (N_2289,N_1757,N_1755);
and U2290 (N_2290,N_1731,N_1557);
or U2291 (N_2291,N_1834,N_1689);
nor U2292 (N_2292,N_1980,N_1890);
or U2293 (N_2293,N_1691,N_1855);
and U2294 (N_2294,N_1727,N_1721);
nor U2295 (N_2295,N_1701,N_1820);
and U2296 (N_2296,N_1623,N_1600);
nand U2297 (N_2297,N_1875,N_1603);
or U2298 (N_2298,N_1563,N_1703);
or U2299 (N_2299,N_1660,N_1559);
xnor U2300 (N_2300,N_1915,N_1725);
nor U2301 (N_2301,N_1977,N_1917);
or U2302 (N_2302,N_1979,N_1830);
and U2303 (N_2303,N_1592,N_1537);
nand U2304 (N_2304,N_1720,N_1781);
or U2305 (N_2305,N_1684,N_1779);
nor U2306 (N_2306,N_1682,N_1531);
or U2307 (N_2307,N_1752,N_1675);
or U2308 (N_2308,N_1899,N_1875);
nor U2309 (N_2309,N_1846,N_1761);
or U2310 (N_2310,N_1709,N_1817);
and U2311 (N_2311,N_1851,N_1832);
nand U2312 (N_2312,N_1993,N_1677);
nand U2313 (N_2313,N_1522,N_1584);
nand U2314 (N_2314,N_1761,N_1627);
nand U2315 (N_2315,N_1659,N_1525);
and U2316 (N_2316,N_1943,N_1573);
nor U2317 (N_2317,N_1734,N_1530);
nor U2318 (N_2318,N_1743,N_1697);
nor U2319 (N_2319,N_1965,N_1828);
nand U2320 (N_2320,N_1615,N_1652);
and U2321 (N_2321,N_1963,N_1854);
nand U2322 (N_2322,N_1537,N_1768);
and U2323 (N_2323,N_1900,N_1781);
nand U2324 (N_2324,N_1586,N_1947);
or U2325 (N_2325,N_1565,N_1984);
or U2326 (N_2326,N_1716,N_1567);
nor U2327 (N_2327,N_1545,N_1629);
and U2328 (N_2328,N_1520,N_1976);
nor U2329 (N_2329,N_1774,N_1566);
nand U2330 (N_2330,N_1598,N_1655);
and U2331 (N_2331,N_1701,N_1598);
or U2332 (N_2332,N_1701,N_1599);
or U2333 (N_2333,N_1907,N_1964);
or U2334 (N_2334,N_1924,N_1933);
or U2335 (N_2335,N_1797,N_1743);
nand U2336 (N_2336,N_1932,N_1638);
nor U2337 (N_2337,N_1578,N_1694);
nand U2338 (N_2338,N_1583,N_1676);
nor U2339 (N_2339,N_1928,N_1620);
or U2340 (N_2340,N_1837,N_1828);
or U2341 (N_2341,N_1736,N_1644);
nand U2342 (N_2342,N_1556,N_1860);
and U2343 (N_2343,N_1622,N_1898);
and U2344 (N_2344,N_1536,N_1957);
nand U2345 (N_2345,N_1809,N_1867);
nand U2346 (N_2346,N_1811,N_1581);
nor U2347 (N_2347,N_1971,N_1763);
or U2348 (N_2348,N_1770,N_1600);
and U2349 (N_2349,N_1964,N_1960);
nand U2350 (N_2350,N_1691,N_1677);
or U2351 (N_2351,N_1502,N_1620);
and U2352 (N_2352,N_1543,N_1770);
and U2353 (N_2353,N_1545,N_1932);
nor U2354 (N_2354,N_1715,N_1935);
and U2355 (N_2355,N_1790,N_1912);
nand U2356 (N_2356,N_1845,N_1500);
and U2357 (N_2357,N_1883,N_1531);
nor U2358 (N_2358,N_1735,N_1653);
nand U2359 (N_2359,N_1560,N_1698);
and U2360 (N_2360,N_1757,N_1695);
or U2361 (N_2361,N_1539,N_1799);
and U2362 (N_2362,N_1759,N_1753);
and U2363 (N_2363,N_1708,N_1948);
nor U2364 (N_2364,N_1681,N_1964);
or U2365 (N_2365,N_1685,N_1610);
nand U2366 (N_2366,N_1928,N_1762);
and U2367 (N_2367,N_1528,N_1713);
and U2368 (N_2368,N_1579,N_1952);
xor U2369 (N_2369,N_1850,N_1703);
nor U2370 (N_2370,N_1930,N_1545);
nor U2371 (N_2371,N_1716,N_1538);
and U2372 (N_2372,N_1562,N_1759);
nand U2373 (N_2373,N_1753,N_1909);
nor U2374 (N_2374,N_1759,N_1848);
and U2375 (N_2375,N_1808,N_1847);
nor U2376 (N_2376,N_1733,N_1842);
or U2377 (N_2377,N_1786,N_1837);
nand U2378 (N_2378,N_1515,N_1505);
nor U2379 (N_2379,N_1618,N_1728);
or U2380 (N_2380,N_1734,N_1801);
and U2381 (N_2381,N_1707,N_1505);
xnor U2382 (N_2382,N_1940,N_1589);
and U2383 (N_2383,N_1976,N_1754);
or U2384 (N_2384,N_1533,N_1845);
nand U2385 (N_2385,N_1512,N_1882);
nor U2386 (N_2386,N_1746,N_1928);
or U2387 (N_2387,N_1608,N_1704);
or U2388 (N_2388,N_1575,N_1656);
and U2389 (N_2389,N_1925,N_1916);
xnor U2390 (N_2390,N_1651,N_1963);
nor U2391 (N_2391,N_1831,N_1838);
nand U2392 (N_2392,N_1716,N_1642);
nor U2393 (N_2393,N_1639,N_1674);
or U2394 (N_2394,N_1530,N_1505);
nand U2395 (N_2395,N_1772,N_1545);
nor U2396 (N_2396,N_1956,N_1899);
and U2397 (N_2397,N_1690,N_1728);
nor U2398 (N_2398,N_1843,N_1635);
nand U2399 (N_2399,N_1536,N_1687);
or U2400 (N_2400,N_1652,N_1594);
nor U2401 (N_2401,N_1623,N_1722);
nor U2402 (N_2402,N_1979,N_1602);
nand U2403 (N_2403,N_1808,N_1752);
and U2404 (N_2404,N_1919,N_1756);
nor U2405 (N_2405,N_1703,N_1970);
nor U2406 (N_2406,N_1795,N_1615);
nand U2407 (N_2407,N_1867,N_1878);
nand U2408 (N_2408,N_1759,N_1683);
or U2409 (N_2409,N_1818,N_1749);
nor U2410 (N_2410,N_1885,N_1905);
nor U2411 (N_2411,N_1785,N_1905);
nand U2412 (N_2412,N_1657,N_1548);
nand U2413 (N_2413,N_1840,N_1579);
or U2414 (N_2414,N_1835,N_1660);
or U2415 (N_2415,N_1939,N_1536);
and U2416 (N_2416,N_1746,N_1518);
nor U2417 (N_2417,N_1967,N_1537);
nand U2418 (N_2418,N_1864,N_1886);
or U2419 (N_2419,N_1862,N_1951);
nor U2420 (N_2420,N_1581,N_1681);
nor U2421 (N_2421,N_1669,N_1688);
and U2422 (N_2422,N_1979,N_1588);
and U2423 (N_2423,N_1846,N_1823);
nand U2424 (N_2424,N_1934,N_1804);
nand U2425 (N_2425,N_1535,N_1694);
and U2426 (N_2426,N_1899,N_1866);
nand U2427 (N_2427,N_1889,N_1519);
or U2428 (N_2428,N_1615,N_1805);
and U2429 (N_2429,N_1800,N_1896);
nor U2430 (N_2430,N_1688,N_1595);
nand U2431 (N_2431,N_1657,N_1582);
nand U2432 (N_2432,N_1824,N_1970);
and U2433 (N_2433,N_1936,N_1753);
and U2434 (N_2434,N_1936,N_1885);
nor U2435 (N_2435,N_1838,N_1989);
or U2436 (N_2436,N_1539,N_1553);
nor U2437 (N_2437,N_1704,N_1517);
and U2438 (N_2438,N_1875,N_1837);
and U2439 (N_2439,N_1738,N_1715);
or U2440 (N_2440,N_1801,N_1781);
or U2441 (N_2441,N_1872,N_1728);
nor U2442 (N_2442,N_1625,N_1785);
or U2443 (N_2443,N_1776,N_1558);
nor U2444 (N_2444,N_1709,N_1613);
or U2445 (N_2445,N_1544,N_1836);
or U2446 (N_2446,N_1978,N_1771);
and U2447 (N_2447,N_1739,N_1697);
and U2448 (N_2448,N_1867,N_1851);
nand U2449 (N_2449,N_1627,N_1723);
or U2450 (N_2450,N_1818,N_1744);
or U2451 (N_2451,N_1553,N_1831);
nand U2452 (N_2452,N_1972,N_1943);
or U2453 (N_2453,N_1771,N_1824);
or U2454 (N_2454,N_1628,N_1563);
nor U2455 (N_2455,N_1655,N_1853);
nand U2456 (N_2456,N_1507,N_1792);
and U2457 (N_2457,N_1930,N_1660);
nand U2458 (N_2458,N_1730,N_1868);
xor U2459 (N_2459,N_1813,N_1606);
and U2460 (N_2460,N_1675,N_1875);
or U2461 (N_2461,N_1698,N_1999);
or U2462 (N_2462,N_1751,N_1830);
nand U2463 (N_2463,N_1854,N_1995);
or U2464 (N_2464,N_1507,N_1866);
and U2465 (N_2465,N_1809,N_1630);
or U2466 (N_2466,N_1647,N_1855);
nor U2467 (N_2467,N_1541,N_1943);
and U2468 (N_2468,N_1725,N_1955);
and U2469 (N_2469,N_1959,N_1694);
and U2470 (N_2470,N_1720,N_1842);
nand U2471 (N_2471,N_1748,N_1842);
and U2472 (N_2472,N_1534,N_1931);
nor U2473 (N_2473,N_1737,N_1893);
or U2474 (N_2474,N_1953,N_1511);
or U2475 (N_2475,N_1628,N_1754);
nor U2476 (N_2476,N_1796,N_1762);
nand U2477 (N_2477,N_1697,N_1805);
and U2478 (N_2478,N_1725,N_1555);
or U2479 (N_2479,N_1886,N_1717);
and U2480 (N_2480,N_1759,N_1971);
or U2481 (N_2481,N_1802,N_1717);
nand U2482 (N_2482,N_1888,N_1989);
and U2483 (N_2483,N_1561,N_1612);
or U2484 (N_2484,N_1962,N_1514);
and U2485 (N_2485,N_1686,N_1814);
or U2486 (N_2486,N_1626,N_1895);
or U2487 (N_2487,N_1584,N_1798);
and U2488 (N_2488,N_1637,N_1796);
nand U2489 (N_2489,N_1840,N_1505);
nor U2490 (N_2490,N_1769,N_1648);
and U2491 (N_2491,N_1919,N_1943);
or U2492 (N_2492,N_1653,N_1559);
and U2493 (N_2493,N_1766,N_1750);
nor U2494 (N_2494,N_1738,N_1766);
or U2495 (N_2495,N_1808,N_1713);
or U2496 (N_2496,N_1583,N_1500);
nand U2497 (N_2497,N_1726,N_1721);
and U2498 (N_2498,N_1588,N_1661);
or U2499 (N_2499,N_1857,N_1532);
nand U2500 (N_2500,N_2157,N_2162);
or U2501 (N_2501,N_2088,N_2321);
or U2502 (N_2502,N_2420,N_2163);
or U2503 (N_2503,N_2059,N_2236);
or U2504 (N_2504,N_2017,N_2091);
and U2505 (N_2505,N_2192,N_2378);
nand U2506 (N_2506,N_2415,N_2367);
and U2507 (N_2507,N_2285,N_2290);
and U2508 (N_2508,N_2366,N_2279);
and U2509 (N_2509,N_2408,N_2156);
nand U2510 (N_2510,N_2451,N_2147);
nor U2511 (N_2511,N_2254,N_2388);
nand U2512 (N_2512,N_2233,N_2095);
and U2513 (N_2513,N_2151,N_2448);
nand U2514 (N_2514,N_2122,N_2427);
nand U2515 (N_2515,N_2120,N_2019);
nor U2516 (N_2516,N_2127,N_2387);
nand U2517 (N_2517,N_2014,N_2208);
and U2518 (N_2518,N_2328,N_2010);
nand U2519 (N_2519,N_2214,N_2093);
and U2520 (N_2520,N_2228,N_2286);
nand U2521 (N_2521,N_2131,N_2354);
or U2522 (N_2522,N_2237,N_2128);
nand U2523 (N_2523,N_2124,N_2073);
nor U2524 (N_2524,N_2260,N_2270);
xor U2525 (N_2525,N_2339,N_2158);
and U2526 (N_2526,N_2170,N_2206);
and U2527 (N_2527,N_2240,N_2198);
or U2528 (N_2528,N_2202,N_2497);
or U2529 (N_2529,N_2089,N_2035);
nor U2530 (N_2530,N_2051,N_2160);
and U2531 (N_2531,N_2074,N_2449);
or U2532 (N_2532,N_2075,N_2345);
nand U2533 (N_2533,N_2047,N_2469);
nor U2534 (N_2534,N_2334,N_2435);
and U2535 (N_2535,N_2018,N_2331);
and U2536 (N_2536,N_2273,N_2213);
or U2537 (N_2537,N_2101,N_2249);
and U2538 (N_2538,N_2087,N_2210);
nor U2539 (N_2539,N_2402,N_2178);
nand U2540 (N_2540,N_2168,N_2302);
nor U2541 (N_2541,N_2486,N_2048);
nor U2542 (N_2542,N_2252,N_2153);
or U2543 (N_2543,N_2409,N_2284);
nor U2544 (N_2544,N_2262,N_2108);
and U2545 (N_2545,N_2460,N_2023);
xnor U2546 (N_2546,N_2197,N_2139);
or U2547 (N_2547,N_2426,N_2396);
or U2548 (N_2548,N_2340,N_2322);
nand U2549 (N_2549,N_2096,N_2114);
nor U2550 (N_2550,N_2304,N_2195);
nand U2551 (N_2551,N_2294,N_2133);
or U2552 (N_2552,N_2393,N_2244);
or U2553 (N_2553,N_2433,N_2394);
or U2554 (N_2554,N_2134,N_2490);
nand U2555 (N_2555,N_2314,N_2392);
nand U2556 (N_2556,N_2453,N_2476);
and U2557 (N_2557,N_2105,N_2325);
and U2558 (N_2558,N_2312,N_2385);
nand U2559 (N_2559,N_2376,N_2319);
nor U2560 (N_2560,N_2186,N_2231);
and U2561 (N_2561,N_2026,N_2188);
or U2562 (N_2562,N_2422,N_2012);
or U2563 (N_2563,N_2103,N_2100);
and U2564 (N_2564,N_2138,N_2078);
and U2565 (N_2565,N_2474,N_2099);
nor U2566 (N_2566,N_2002,N_2226);
nand U2567 (N_2567,N_2011,N_2470);
or U2568 (N_2568,N_2232,N_2291);
or U2569 (N_2569,N_2377,N_2152);
xnor U2570 (N_2570,N_2230,N_2225);
or U2571 (N_2571,N_2116,N_2301);
nand U2572 (N_2572,N_2203,N_2084);
or U2573 (N_2573,N_2318,N_2067);
nor U2574 (N_2574,N_2382,N_2375);
and U2575 (N_2575,N_2117,N_2481);
nor U2576 (N_2576,N_2159,N_2185);
nand U2577 (N_2577,N_2347,N_2038);
and U2578 (N_2578,N_2052,N_2429);
nand U2579 (N_2579,N_2313,N_2349);
or U2580 (N_2580,N_2438,N_2261);
nand U2581 (N_2581,N_2494,N_2234);
nor U2582 (N_2582,N_2498,N_2459);
or U2583 (N_2583,N_2403,N_2115);
or U2584 (N_2584,N_2140,N_2293);
or U2585 (N_2585,N_2055,N_2323);
or U2586 (N_2586,N_2330,N_2274);
or U2587 (N_2587,N_2471,N_2348);
and U2588 (N_2588,N_2063,N_2370);
nor U2589 (N_2589,N_2399,N_2257);
nand U2590 (N_2590,N_2480,N_2253);
nand U2591 (N_2591,N_2043,N_2307);
xnor U2592 (N_2592,N_2295,N_2412);
nand U2593 (N_2593,N_2364,N_2373);
nor U2594 (N_2594,N_2411,N_2276);
or U2595 (N_2595,N_2424,N_2333);
nand U2596 (N_2596,N_2033,N_2166);
nand U2597 (N_2597,N_2468,N_2109);
nor U2598 (N_2598,N_2269,N_2071);
or U2599 (N_2599,N_2280,N_2265);
and U2600 (N_2600,N_2037,N_2288);
and U2601 (N_2601,N_2219,N_2430);
nor U2602 (N_2602,N_2007,N_2371);
or U2603 (N_2603,N_2241,N_2341);
or U2604 (N_2604,N_2344,N_2191);
nand U2605 (N_2605,N_2224,N_2369);
or U2606 (N_2606,N_2303,N_2275);
nor U2607 (N_2607,N_2094,N_2024);
nor U2608 (N_2608,N_2085,N_2003);
nor U2609 (N_2609,N_2172,N_2077);
and U2610 (N_2610,N_2229,N_2287);
and U2611 (N_2611,N_2247,N_2455);
nand U2612 (N_2612,N_2358,N_2218);
nor U2613 (N_2613,N_2194,N_2404);
and U2614 (N_2614,N_2296,N_2183);
and U2615 (N_2615,N_2031,N_2278);
nand U2616 (N_2616,N_2040,N_2221);
and U2617 (N_2617,N_2246,N_2362);
or U2618 (N_2618,N_2454,N_2013);
nor U2619 (N_2619,N_2395,N_2467);
nand U2620 (N_2620,N_2222,N_2060);
nor U2621 (N_2621,N_2053,N_2189);
nand U2622 (N_2622,N_2000,N_2207);
and U2623 (N_2623,N_2169,N_2416);
nand U2624 (N_2624,N_2125,N_2315);
nand U2625 (N_2625,N_2058,N_2390);
or U2626 (N_2626,N_2311,N_2054);
and U2627 (N_2627,N_2363,N_2006);
nor U2628 (N_2628,N_2201,N_2450);
nand U2629 (N_2629,N_2266,N_2118);
or U2630 (N_2630,N_2021,N_2272);
and U2631 (N_2631,N_2346,N_2149);
and U2632 (N_2632,N_2457,N_2258);
xor U2633 (N_2633,N_2475,N_2329);
or U2634 (N_2634,N_2143,N_2335);
or U2635 (N_2635,N_2056,N_2381);
and U2636 (N_2636,N_2405,N_2015);
or U2637 (N_2637,N_2097,N_2352);
and U2638 (N_2638,N_2282,N_2167);
and U2639 (N_2639,N_2034,N_2179);
nand U2640 (N_2640,N_2441,N_2235);
or U2641 (N_2641,N_2401,N_2025);
xor U2642 (N_2642,N_2081,N_2400);
or U2643 (N_2643,N_2123,N_2478);
or U2644 (N_2644,N_2466,N_2144);
nor U2645 (N_2645,N_2150,N_2141);
nor U2646 (N_2646,N_2112,N_2428);
and U2647 (N_2647,N_2447,N_2041);
or U2648 (N_2648,N_2050,N_2181);
nand U2649 (N_2649,N_2022,N_2004);
and U2650 (N_2650,N_2142,N_2297);
nor U2651 (N_2651,N_2353,N_2332);
nand U2652 (N_2652,N_2001,N_2223);
or U2653 (N_2653,N_2417,N_2174);
and U2654 (N_2654,N_2456,N_2431);
nand U2655 (N_2655,N_2492,N_2308);
and U2656 (N_2656,N_2436,N_2082);
and U2657 (N_2657,N_2320,N_2028);
nor U2658 (N_2658,N_2488,N_2386);
or U2659 (N_2659,N_2104,N_2343);
or U2660 (N_2660,N_2046,N_2391);
nor U2661 (N_2661,N_2227,N_2365);
and U2662 (N_2662,N_2016,N_2216);
nand U2663 (N_2663,N_2200,N_2472);
and U2664 (N_2664,N_2215,N_2355);
nand U2665 (N_2665,N_2477,N_2379);
or U2666 (N_2666,N_2171,N_2076);
nand U2667 (N_2667,N_2398,N_2102);
nand U2668 (N_2668,N_2305,N_2439);
nor U2669 (N_2669,N_2268,N_2072);
xnor U2670 (N_2670,N_2337,N_2482);
or U2671 (N_2671,N_2238,N_2175);
nor U2672 (N_2672,N_2090,N_2298);
or U2673 (N_2673,N_2130,N_2137);
and U2674 (N_2674,N_2299,N_2092);
nand U2675 (N_2675,N_2211,N_2489);
nand U2676 (N_2676,N_2368,N_2487);
nor U2677 (N_2677,N_2380,N_2042);
or U2678 (N_2678,N_2154,N_2190);
and U2679 (N_2679,N_2389,N_2484);
nor U2680 (N_2680,N_2316,N_2248);
or U2681 (N_2681,N_2180,N_2289);
nor U2682 (N_2682,N_2145,N_2239);
nand U2683 (N_2683,N_2267,N_2086);
nor U2684 (N_2684,N_2446,N_2057);
nand U2685 (N_2685,N_2132,N_2217);
nor U2686 (N_2686,N_2107,N_2350);
nor U2687 (N_2687,N_2164,N_2464);
or U2688 (N_2688,N_2111,N_2044);
or U2689 (N_2689,N_2277,N_2309);
and U2690 (N_2690,N_2220,N_2106);
nand U2691 (N_2691,N_2342,N_2418);
and U2692 (N_2692,N_2136,N_2423);
or U2693 (N_2693,N_2281,N_2338);
or U2694 (N_2694,N_2271,N_2126);
and U2695 (N_2695,N_2483,N_2110);
and U2696 (N_2696,N_2351,N_2146);
and U2697 (N_2697,N_2184,N_2205);
nor U2698 (N_2698,N_2425,N_2256);
nand U2699 (N_2699,N_2324,N_2173);
nand U2700 (N_2700,N_2264,N_2327);
nand U2701 (N_2701,N_2283,N_2204);
and U2702 (N_2702,N_2461,N_2070);
and U2703 (N_2703,N_2442,N_2473);
and U2704 (N_2704,N_2199,N_2493);
nor U2705 (N_2705,N_2036,N_2255);
and U2706 (N_2706,N_2361,N_2119);
nand U2707 (N_2707,N_2458,N_2129);
or U2708 (N_2708,N_2030,N_2432);
or U2709 (N_2709,N_2182,N_2005);
nand U2710 (N_2710,N_2359,N_2064);
and U2711 (N_2711,N_2406,N_2374);
nand U2712 (N_2712,N_2300,N_2434);
nor U2713 (N_2713,N_2029,N_2360);
nand U2714 (N_2714,N_2080,N_2135);
xnor U2715 (N_2715,N_2496,N_2336);
or U2716 (N_2716,N_2421,N_2068);
or U2717 (N_2717,N_2397,N_2292);
xnor U2718 (N_2718,N_2049,N_2485);
nand U2719 (N_2719,N_2009,N_2414);
nand U2720 (N_2720,N_2243,N_2209);
nor U2721 (N_2721,N_2020,N_2263);
nor U2722 (N_2722,N_2465,N_2027);
and U2723 (N_2723,N_2039,N_2245);
and U2724 (N_2724,N_2413,N_2079);
or U2725 (N_2725,N_2445,N_2407);
and U2726 (N_2726,N_2383,N_2251);
or U2727 (N_2727,N_2032,N_2410);
and U2728 (N_2728,N_2065,N_2193);
or U2729 (N_2729,N_2499,N_2187);
or U2730 (N_2730,N_2155,N_2443);
and U2731 (N_2731,N_2419,N_2495);
or U2732 (N_2732,N_2452,N_2463);
and U2733 (N_2733,N_2491,N_2098);
and U2734 (N_2734,N_2444,N_2310);
nor U2735 (N_2735,N_2306,N_2196);
and U2736 (N_2736,N_2357,N_2069);
nor U2737 (N_2737,N_2121,N_2045);
nor U2738 (N_2738,N_2326,N_2440);
and U2739 (N_2739,N_2250,N_2177);
nand U2740 (N_2740,N_2462,N_2165);
nor U2741 (N_2741,N_2437,N_2317);
nand U2742 (N_2742,N_2061,N_2356);
nand U2743 (N_2743,N_2066,N_2148);
nor U2744 (N_2744,N_2008,N_2161);
and U2745 (N_2745,N_2176,N_2212);
and U2746 (N_2746,N_2083,N_2242);
and U2747 (N_2747,N_2372,N_2384);
nor U2748 (N_2748,N_2479,N_2259);
nor U2749 (N_2749,N_2062,N_2113);
and U2750 (N_2750,N_2401,N_2044);
and U2751 (N_2751,N_2121,N_2040);
or U2752 (N_2752,N_2408,N_2357);
or U2753 (N_2753,N_2355,N_2477);
nand U2754 (N_2754,N_2322,N_2039);
and U2755 (N_2755,N_2351,N_2045);
nand U2756 (N_2756,N_2087,N_2348);
xnor U2757 (N_2757,N_2091,N_2246);
nand U2758 (N_2758,N_2285,N_2261);
nand U2759 (N_2759,N_2499,N_2143);
nand U2760 (N_2760,N_2142,N_2070);
and U2761 (N_2761,N_2367,N_2368);
nor U2762 (N_2762,N_2442,N_2216);
and U2763 (N_2763,N_2465,N_2217);
and U2764 (N_2764,N_2088,N_2296);
and U2765 (N_2765,N_2494,N_2291);
and U2766 (N_2766,N_2306,N_2406);
nor U2767 (N_2767,N_2119,N_2348);
or U2768 (N_2768,N_2420,N_2192);
nand U2769 (N_2769,N_2120,N_2497);
and U2770 (N_2770,N_2041,N_2223);
or U2771 (N_2771,N_2140,N_2443);
nor U2772 (N_2772,N_2109,N_2450);
nor U2773 (N_2773,N_2370,N_2410);
nand U2774 (N_2774,N_2430,N_2264);
and U2775 (N_2775,N_2203,N_2019);
nor U2776 (N_2776,N_2411,N_2331);
and U2777 (N_2777,N_2168,N_2332);
xnor U2778 (N_2778,N_2009,N_2167);
and U2779 (N_2779,N_2492,N_2309);
nor U2780 (N_2780,N_2457,N_2331);
and U2781 (N_2781,N_2313,N_2410);
nor U2782 (N_2782,N_2254,N_2054);
nand U2783 (N_2783,N_2208,N_2394);
nor U2784 (N_2784,N_2380,N_2384);
nand U2785 (N_2785,N_2418,N_2201);
nor U2786 (N_2786,N_2214,N_2005);
nor U2787 (N_2787,N_2096,N_2389);
nor U2788 (N_2788,N_2310,N_2076);
and U2789 (N_2789,N_2095,N_2108);
and U2790 (N_2790,N_2177,N_2118);
and U2791 (N_2791,N_2463,N_2462);
nand U2792 (N_2792,N_2320,N_2402);
nor U2793 (N_2793,N_2417,N_2469);
and U2794 (N_2794,N_2321,N_2427);
nand U2795 (N_2795,N_2319,N_2275);
or U2796 (N_2796,N_2083,N_2425);
or U2797 (N_2797,N_2139,N_2391);
and U2798 (N_2798,N_2425,N_2141);
nand U2799 (N_2799,N_2222,N_2429);
or U2800 (N_2800,N_2429,N_2416);
nand U2801 (N_2801,N_2304,N_2208);
nor U2802 (N_2802,N_2433,N_2290);
and U2803 (N_2803,N_2074,N_2424);
nor U2804 (N_2804,N_2172,N_2295);
nand U2805 (N_2805,N_2462,N_2000);
nor U2806 (N_2806,N_2069,N_2264);
and U2807 (N_2807,N_2460,N_2190);
nor U2808 (N_2808,N_2258,N_2093);
nor U2809 (N_2809,N_2183,N_2098);
and U2810 (N_2810,N_2496,N_2451);
and U2811 (N_2811,N_2417,N_2429);
and U2812 (N_2812,N_2494,N_2183);
nor U2813 (N_2813,N_2326,N_2470);
nor U2814 (N_2814,N_2279,N_2234);
nor U2815 (N_2815,N_2420,N_2161);
and U2816 (N_2816,N_2238,N_2282);
nand U2817 (N_2817,N_2085,N_2488);
nand U2818 (N_2818,N_2095,N_2440);
or U2819 (N_2819,N_2250,N_2016);
or U2820 (N_2820,N_2276,N_2157);
nor U2821 (N_2821,N_2225,N_2190);
xnor U2822 (N_2822,N_2119,N_2320);
nand U2823 (N_2823,N_2382,N_2332);
or U2824 (N_2824,N_2170,N_2319);
or U2825 (N_2825,N_2420,N_2250);
nand U2826 (N_2826,N_2078,N_2043);
and U2827 (N_2827,N_2340,N_2258);
nor U2828 (N_2828,N_2286,N_2116);
and U2829 (N_2829,N_2004,N_2024);
nor U2830 (N_2830,N_2368,N_2252);
and U2831 (N_2831,N_2387,N_2466);
nand U2832 (N_2832,N_2275,N_2350);
nand U2833 (N_2833,N_2305,N_2095);
and U2834 (N_2834,N_2347,N_2080);
xor U2835 (N_2835,N_2476,N_2123);
nand U2836 (N_2836,N_2453,N_2468);
nand U2837 (N_2837,N_2168,N_2370);
or U2838 (N_2838,N_2370,N_2258);
and U2839 (N_2839,N_2000,N_2224);
nor U2840 (N_2840,N_2392,N_2066);
and U2841 (N_2841,N_2135,N_2294);
nand U2842 (N_2842,N_2280,N_2215);
xnor U2843 (N_2843,N_2400,N_2467);
xor U2844 (N_2844,N_2269,N_2281);
nor U2845 (N_2845,N_2309,N_2230);
nand U2846 (N_2846,N_2477,N_2178);
nor U2847 (N_2847,N_2466,N_2425);
nor U2848 (N_2848,N_2441,N_2432);
nor U2849 (N_2849,N_2057,N_2100);
nor U2850 (N_2850,N_2321,N_2131);
nand U2851 (N_2851,N_2029,N_2275);
and U2852 (N_2852,N_2326,N_2206);
nor U2853 (N_2853,N_2491,N_2285);
and U2854 (N_2854,N_2292,N_2479);
nor U2855 (N_2855,N_2385,N_2278);
or U2856 (N_2856,N_2028,N_2355);
nor U2857 (N_2857,N_2026,N_2135);
and U2858 (N_2858,N_2404,N_2166);
nand U2859 (N_2859,N_2288,N_2378);
nand U2860 (N_2860,N_2152,N_2409);
or U2861 (N_2861,N_2033,N_2394);
and U2862 (N_2862,N_2188,N_2466);
nand U2863 (N_2863,N_2463,N_2419);
or U2864 (N_2864,N_2021,N_2461);
xnor U2865 (N_2865,N_2293,N_2055);
xnor U2866 (N_2866,N_2005,N_2442);
or U2867 (N_2867,N_2089,N_2086);
nand U2868 (N_2868,N_2194,N_2137);
or U2869 (N_2869,N_2297,N_2229);
or U2870 (N_2870,N_2496,N_2195);
nand U2871 (N_2871,N_2425,N_2115);
nand U2872 (N_2872,N_2072,N_2449);
or U2873 (N_2873,N_2101,N_2109);
and U2874 (N_2874,N_2158,N_2084);
nor U2875 (N_2875,N_2050,N_2227);
and U2876 (N_2876,N_2405,N_2158);
nand U2877 (N_2877,N_2050,N_2283);
nor U2878 (N_2878,N_2124,N_2299);
and U2879 (N_2879,N_2445,N_2153);
nand U2880 (N_2880,N_2084,N_2016);
and U2881 (N_2881,N_2359,N_2369);
or U2882 (N_2882,N_2276,N_2453);
nand U2883 (N_2883,N_2244,N_2012);
and U2884 (N_2884,N_2494,N_2499);
or U2885 (N_2885,N_2392,N_2481);
xnor U2886 (N_2886,N_2415,N_2118);
and U2887 (N_2887,N_2391,N_2168);
nor U2888 (N_2888,N_2368,N_2361);
nor U2889 (N_2889,N_2481,N_2166);
nor U2890 (N_2890,N_2458,N_2071);
or U2891 (N_2891,N_2371,N_2412);
nand U2892 (N_2892,N_2212,N_2138);
nand U2893 (N_2893,N_2001,N_2083);
nand U2894 (N_2894,N_2067,N_2404);
nand U2895 (N_2895,N_2213,N_2184);
or U2896 (N_2896,N_2477,N_2015);
nand U2897 (N_2897,N_2101,N_2296);
nor U2898 (N_2898,N_2492,N_2365);
and U2899 (N_2899,N_2218,N_2350);
nor U2900 (N_2900,N_2329,N_2278);
nor U2901 (N_2901,N_2050,N_2039);
or U2902 (N_2902,N_2119,N_2116);
and U2903 (N_2903,N_2328,N_2011);
nand U2904 (N_2904,N_2095,N_2105);
nor U2905 (N_2905,N_2053,N_2177);
and U2906 (N_2906,N_2477,N_2485);
and U2907 (N_2907,N_2438,N_2015);
nor U2908 (N_2908,N_2167,N_2164);
nor U2909 (N_2909,N_2181,N_2008);
and U2910 (N_2910,N_2434,N_2139);
nor U2911 (N_2911,N_2033,N_2064);
and U2912 (N_2912,N_2023,N_2195);
or U2913 (N_2913,N_2037,N_2116);
or U2914 (N_2914,N_2018,N_2402);
nor U2915 (N_2915,N_2311,N_2401);
nor U2916 (N_2916,N_2451,N_2069);
and U2917 (N_2917,N_2036,N_2317);
or U2918 (N_2918,N_2204,N_2371);
or U2919 (N_2919,N_2302,N_2011);
nor U2920 (N_2920,N_2114,N_2100);
and U2921 (N_2921,N_2122,N_2015);
xnor U2922 (N_2922,N_2266,N_2394);
nor U2923 (N_2923,N_2404,N_2157);
nand U2924 (N_2924,N_2455,N_2197);
nand U2925 (N_2925,N_2179,N_2396);
or U2926 (N_2926,N_2387,N_2006);
nor U2927 (N_2927,N_2262,N_2210);
and U2928 (N_2928,N_2031,N_2438);
or U2929 (N_2929,N_2395,N_2328);
nand U2930 (N_2930,N_2325,N_2410);
nand U2931 (N_2931,N_2497,N_2072);
and U2932 (N_2932,N_2042,N_2221);
nand U2933 (N_2933,N_2034,N_2441);
nand U2934 (N_2934,N_2349,N_2095);
nand U2935 (N_2935,N_2186,N_2289);
or U2936 (N_2936,N_2340,N_2371);
nand U2937 (N_2937,N_2415,N_2470);
or U2938 (N_2938,N_2495,N_2094);
or U2939 (N_2939,N_2096,N_2299);
nand U2940 (N_2940,N_2200,N_2491);
nor U2941 (N_2941,N_2264,N_2433);
nor U2942 (N_2942,N_2148,N_2155);
nor U2943 (N_2943,N_2417,N_2416);
or U2944 (N_2944,N_2176,N_2354);
or U2945 (N_2945,N_2097,N_2398);
nor U2946 (N_2946,N_2239,N_2341);
or U2947 (N_2947,N_2348,N_2166);
or U2948 (N_2948,N_2019,N_2218);
and U2949 (N_2949,N_2117,N_2118);
nand U2950 (N_2950,N_2076,N_2446);
nor U2951 (N_2951,N_2325,N_2095);
nand U2952 (N_2952,N_2137,N_2207);
nor U2953 (N_2953,N_2157,N_2328);
or U2954 (N_2954,N_2043,N_2488);
or U2955 (N_2955,N_2037,N_2370);
and U2956 (N_2956,N_2254,N_2185);
or U2957 (N_2957,N_2342,N_2019);
and U2958 (N_2958,N_2100,N_2276);
nor U2959 (N_2959,N_2098,N_2114);
nor U2960 (N_2960,N_2130,N_2435);
nor U2961 (N_2961,N_2008,N_2035);
and U2962 (N_2962,N_2261,N_2367);
and U2963 (N_2963,N_2226,N_2026);
and U2964 (N_2964,N_2394,N_2203);
nor U2965 (N_2965,N_2372,N_2367);
nor U2966 (N_2966,N_2375,N_2303);
nand U2967 (N_2967,N_2062,N_2033);
nand U2968 (N_2968,N_2039,N_2314);
or U2969 (N_2969,N_2114,N_2264);
nand U2970 (N_2970,N_2381,N_2497);
nor U2971 (N_2971,N_2075,N_2104);
or U2972 (N_2972,N_2053,N_2067);
nor U2973 (N_2973,N_2299,N_2339);
and U2974 (N_2974,N_2035,N_2138);
nand U2975 (N_2975,N_2462,N_2458);
nor U2976 (N_2976,N_2031,N_2315);
and U2977 (N_2977,N_2005,N_2193);
or U2978 (N_2978,N_2149,N_2182);
nor U2979 (N_2979,N_2027,N_2377);
nand U2980 (N_2980,N_2058,N_2370);
and U2981 (N_2981,N_2364,N_2214);
or U2982 (N_2982,N_2173,N_2272);
and U2983 (N_2983,N_2265,N_2273);
and U2984 (N_2984,N_2150,N_2248);
or U2985 (N_2985,N_2455,N_2442);
nand U2986 (N_2986,N_2499,N_2212);
nand U2987 (N_2987,N_2411,N_2113);
nand U2988 (N_2988,N_2360,N_2377);
nand U2989 (N_2989,N_2096,N_2439);
and U2990 (N_2990,N_2110,N_2164);
or U2991 (N_2991,N_2124,N_2395);
nand U2992 (N_2992,N_2356,N_2379);
nor U2993 (N_2993,N_2235,N_2095);
or U2994 (N_2994,N_2121,N_2102);
and U2995 (N_2995,N_2227,N_2299);
nand U2996 (N_2996,N_2011,N_2129);
and U2997 (N_2997,N_2027,N_2061);
and U2998 (N_2998,N_2132,N_2200);
nor U2999 (N_2999,N_2175,N_2386);
or U3000 (N_3000,N_2583,N_2530);
and U3001 (N_3001,N_2769,N_2717);
nor U3002 (N_3002,N_2925,N_2928);
nand U3003 (N_3003,N_2724,N_2625);
nor U3004 (N_3004,N_2945,N_2779);
nand U3005 (N_3005,N_2525,N_2721);
nand U3006 (N_3006,N_2771,N_2567);
or U3007 (N_3007,N_2834,N_2923);
or U3008 (N_3008,N_2636,N_2993);
nor U3009 (N_3009,N_2689,N_2927);
nand U3010 (N_3010,N_2648,N_2504);
nand U3011 (N_3011,N_2615,N_2803);
nor U3012 (N_3012,N_2888,N_2586);
nand U3013 (N_3013,N_2835,N_2992);
or U3014 (N_3014,N_2705,N_2505);
nor U3015 (N_3015,N_2612,N_2661);
nor U3016 (N_3016,N_2841,N_2884);
nand U3017 (N_3017,N_2672,N_2654);
nor U3018 (N_3018,N_2783,N_2799);
nand U3019 (N_3019,N_2570,N_2849);
xnor U3020 (N_3020,N_2641,N_2669);
nand U3021 (N_3021,N_2957,N_2659);
or U3022 (N_3022,N_2629,N_2919);
and U3023 (N_3023,N_2962,N_2643);
and U3024 (N_3024,N_2785,N_2857);
and U3025 (N_3025,N_2934,N_2743);
and U3026 (N_3026,N_2577,N_2819);
nand U3027 (N_3027,N_2832,N_2891);
and U3028 (N_3028,N_2594,N_2810);
and U3029 (N_3029,N_2549,N_2958);
nor U3030 (N_3030,N_2870,N_2618);
and U3031 (N_3031,N_2538,N_2844);
xnor U3032 (N_3032,N_2572,N_2741);
nor U3033 (N_3033,N_2806,N_2939);
nand U3034 (N_3034,N_2775,N_2529);
nand U3035 (N_3035,N_2909,N_2889);
or U3036 (N_3036,N_2528,N_2926);
nand U3037 (N_3037,N_2540,N_2951);
nand U3038 (N_3038,N_2593,N_2534);
or U3039 (N_3039,N_2850,N_2952);
or U3040 (N_3040,N_2881,N_2754);
and U3041 (N_3041,N_2997,N_2644);
nor U3042 (N_3042,N_2559,N_2837);
and U3043 (N_3043,N_2851,N_2535);
and U3044 (N_3044,N_2773,N_2899);
nor U3045 (N_3045,N_2581,N_2893);
or U3046 (N_3046,N_2956,N_2500);
and U3047 (N_3047,N_2790,N_2770);
xor U3048 (N_3048,N_2918,N_2886);
nand U3049 (N_3049,N_2902,N_2807);
nor U3050 (N_3050,N_2970,N_2591);
xor U3051 (N_3051,N_2633,N_2587);
nand U3052 (N_3052,N_2766,N_2917);
nor U3053 (N_3053,N_2627,N_2679);
or U3054 (N_3054,N_2816,N_2793);
or U3055 (N_3055,N_2710,N_2647);
and U3056 (N_3056,N_2592,N_2969);
or U3057 (N_3057,N_2777,N_2712);
or U3058 (N_3058,N_2818,N_2650);
nor U3059 (N_3059,N_2795,N_2550);
nand U3060 (N_3060,N_2551,N_2616);
nor U3061 (N_3061,N_2565,N_2573);
and U3062 (N_3062,N_2621,N_2745);
or U3063 (N_3063,N_2516,N_2905);
nor U3064 (N_3064,N_2598,N_2554);
and U3065 (N_3065,N_2742,N_2960);
nand U3066 (N_3066,N_2630,N_2825);
or U3067 (N_3067,N_2739,N_2836);
xnor U3068 (N_3068,N_2533,N_2804);
nand U3069 (N_3069,N_2977,N_2781);
or U3070 (N_3070,N_2617,N_2578);
or U3071 (N_3071,N_2558,N_2678);
nand U3072 (N_3072,N_2757,N_2976);
nand U3073 (N_3073,N_2996,N_2874);
nor U3074 (N_3074,N_2674,N_2588);
nand U3075 (N_3075,N_2882,N_2937);
or U3076 (N_3076,N_2685,N_2511);
nand U3077 (N_3077,N_2994,N_2989);
nand U3078 (N_3078,N_2557,N_2652);
nor U3079 (N_3079,N_2916,N_2722);
nor U3080 (N_3080,N_2896,N_2580);
nand U3081 (N_3081,N_2846,N_2920);
nand U3082 (N_3082,N_2703,N_2760);
nor U3083 (N_3083,N_2887,N_2751);
nor U3084 (N_3084,N_2828,N_2520);
nand U3085 (N_3085,N_2871,N_2866);
or U3086 (N_3086,N_2892,N_2966);
and U3087 (N_3087,N_2744,N_2830);
nand U3088 (N_3088,N_2833,N_2515);
nor U3089 (N_3089,N_2726,N_2898);
nand U3090 (N_3090,N_2660,N_2856);
nand U3091 (N_3091,N_2566,N_2562);
nor U3092 (N_3092,N_2853,N_2708);
nor U3093 (N_3093,N_2702,N_2801);
and U3094 (N_3094,N_2933,N_2658);
or U3095 (N_3095,N_2676,N_2692);
nor U3096 (N_3096,N_2522,N_2548);
nand U3097 (N_3097,N_2867,N_2811);
and U3098 (N_3098,N_2847,N_2576);
and U3099 (N_3099,N_2915,N_2512);
or U3100 (N_3100,N_2827,N_2817);
or U3101 (N_3101,N_2805,N_2697);
nor U3102 (N_3102,N_2946,N_2510);
or U3103 (N_3103,N_2711,N_2634);
or U3104 (N_3104,N_2675,N_2842);
nand U3105 (N_3105,N_2603,N_2747);
nor U3106 (N_3106,N_2531,N_2610);
nor U3107 (N_3107,N_2963,N_2690);
and U3108 (N_3108,N_2686,N_2571);
nor U3109 (N_3109,N_2719,N_2608);
and U3110 (N_3110,N_2714,N_2619);
and U3111 (N_3111,N_2526,N_2517);
nor U3112 (N_3112,N_2713,N_2738);
or U3113 (N_3113,N_2954,N_2749);
nor U3114 (N_3114,N_2746,N_2862);
and U3115 (N_3115,N_2631,N_2778);
nand U3116 (N_3116,N_2519,N_2536);
nand U3117 (N_3117,N_2651,N_2601);
nor U3118 (N_3118,N_2735,N_2514);
nor U3119 (N_3119,N_2907,N_2840);
and U3120 (N_3120,N_2824,N_2663);
nand U3121 (N_3121,N_2639,N_2829);
nand U3122 (N_3122,N_2877,N_2575);
or U3123 (N_3123,N_2750,N_2967);
or U3124 (N_3124,N_2931,N_2688);
nand U3125 (N_3125,N_2869,N_2502);
or U3126 (N_3126,N_2947,N_2622);
nor U3127 (N_3127,N_2890,N_2667);
nand U3128 (N_3128,N_2873,N_2681);
or U3129 (N_3129,N_2910,N_2929);
nand U3130 (N_3130,N_2823,N_2600);
nor U3131 (N_3131,N_2673,N_2604);
nor U3132 (N_3132,N_2642,N_2791);
or U3133 (N_3133,N_2728,N_2949);
xnor U3134 (N_3134,N_2879,N_2765);
nor U3135 (N_3135,N_2950,N_2809);
or U3136 (N_3136,N_2808,N_2941);
or U3137 (N_3137,N_2607,N_2852);
nor U3138 (N_3138,N_2547,N_2718);
nor U3139 (N_3139,N_2943,N_2944);
nand U3140 (N_3140,N_2518,N_2684);
nor U3141 (N_3141,N_2831,N_2839);
and U3142 (N_3142,N_2734,N_2503);
and U3143 (N_3143,N_2513,N_2971);
and U3144 (N_3144,N_2843,N_2983);
nand U3145 (N_3145,N_2693,N_2677);
nor U3146 (N_3146,N_2999,N_2552);
or U3147 (N_3147,N_2820,N_2863);
nand U3148 (N_3148,N_2758,N_2964);
nand U3149 (N_3149,N_2691,N_2628);
and U3150 (N_3150,N_2921,N_2982);
or U3151 (N_3151,N_2759,N_2680);
or U3152 (N_3152,N_2620,N_2955);
and U3153 (N_3153,N_2640,N_2782);
or U3154 (N_3154,N_2815,N_2730);
nor U3155 (N_3155,N_2995,N_2582);
or U3156 (N_3156,N_2541,N_2872);
and U3157 (N_3157,N_2894,N_2657);
nor U3158 (N_3158,N_2737,N_2848);
nand U3159 (N_3159,N_2696,N_2605);
or U3160 (N_3160,N_2859,N_2990);
and U3161 (N_3161,N_2796,N_2595);
and U3162 (N_3162,N_2865,N_2885);
or U3163 (N_3163,N_2638,N_2720);
and U3164 (N_3164,N_2984,N_2752);
nor U3165 (N_3165,N_2875,N_2932);
nor U3166 (N_3166,N_2699,N_2539);
xnor U3167 (N_3167,N_2509,N_2922);
and U3168 (N_3168,N_2597,N_2501);
nor U3169 (N_3169,N_2901,N_2784);
nand U3170 (N_3170,N_2537,N_2764);
xnor U3171 (N_3171,N_2774,N_2991);
and U3172 (N_3172,N_2731,N_2948);
nand U3173 (N_3173,N_2798,N_2561);
nand U3174 (N_3174,N_2864,N_2786);
or U3175 (N_3175,N_2821,N_2506);
and U3176 (N_3176,N_2579,N_2861);
nand U3177 (N_3177,N_2568,N_2792);
nand U3178 (N_3178,N_2961,N_2645);
or U3179 (N_3179,N_2683,N_2632);
nor U3180 (N_3180,N_2706,N_2911);
nand U3181 (N_3181,N_2736,N_2942);
nor U3182 (N_3182,N_2613,N_2838);
or U3183 (N_3183,N_2544,N_2802);
nand U3184 (N_3184,N_2606,N_2975);
nand U3185 (N_3185,N_2546,N_2761);
nand U3186 (N_3186,N_2780,N_2704);
and U3187 (N_3187,N_2959,N_2596);
nand U3188 (N_3188,N_2987,N_2671);
nand U3189 (N_3189,N_2972,N_2687);
nor U3190 (N_3190,N_2564,N_2930);
or U3191 (N_3191,N_2740,N_2878);
nand U3192 (N_3192,N_2755,N_2988);
nor U3193 (N_3193,N_2936,N_2725);
or U3194 (N_3194,N_2543,N_2813);
nand U3195 (N_3195,N_2858,N_2553);
and U3196 (N_3196,N_2729,N_2906);
or U3197 (N_3197,N_2748,N_2590);
nand U3198 (N_3198,N_2584,N_2854);
and U3199 (N_3199,N_2602,N_2521);
and U3200 (N_3200,N_2763,N_2695);
nand U3201 (N_3201,N_2637,N_2787);
and U3202 (N_3202,N_2822,N_2940);
nand U3203 (N_3203,N_2698,N_2973);
nor U3204 (N_3204,N_2979,N_2707);
or U3205 (N_3205,N_2814,N_2666);
nor U3206 (N_3206,N_2694,N_2980);
nand U3207 (N_3207,N_2904,N_2938);
and U3208 (N_3208,N_2880,N_2794);
and U3209 (N_3209,N_2649,N_2998);
nor U3210 (N_3210,N_2756,N_2589);
or U3211 (N_3211,N_2935,N_2924);
and U3212 (N_3212,N_2981,N_2527);
or U3213 (N_3213,N_2732,N_2709);
or U3214 (N_3214,N_2913,N_2665);
nand U3215 (N_3215,N_2767,N_2635);
or U3216 (N_3216,N_2701,N_2903);
nand U3217 (N_3217,N_2855,N_2845);
nand U3218 (N_3218,N_2953,N_2646);
nand U3219 (N_3219,N_2614,N_2965);
nand U3220 (N_3220,N_2883,N_2670);
nand U3221 (N_3221,N_2555,N_2868);
nand U3222 (N_3222,N_2560,N_2978);
and U3223 (N_3223,N_2900,N_2507);
nand U3224 (N_3224,N_2623,N_2800);
xor U3225 (N_3225,N_2532,N_2524);
nor U3226 (N_3226,N_2716,N_2753);
nand U3227 (N_3227,N_2542,N_2599);
or U3228 (N_3228,N_2723,N_2609);
or U3229 (N_3229,N_2876,N_2789);
nor U3230 (N_3230,N_2776,N_2569);
nand U3231 (N_3231,N_2897,N_2733);
or U3232 (N_3232,N_2655,N_2768);
and U3233 (N_3233,N_2611,N_2556);
and U3234 (N_3234,N_2700,N_2986);
and U3235 (N_3235,N_2788,N_2727);
nor U3236 (N_3236,N_2860,N_2653);
nand U3237 (N_3237,N_2715,N_2662);
nor U3238 (N_3238,N_2912,N_2826);
nor U3239 (N_3239,N_2656,N_2772);
and U3240 (N_3240,N_2682,N_2664);
nand U3241 (N_3241,N_2668,N_2985);
xor U3242 (N_3242,N_2968,N_2895);
nor U3243 (N_3243,N_2574,N_2626);
and U3244 (N_3244,N_2585,N_2812);
or U3245 (N_3245,N_2762,N_2624);
nor U3246 (N_3246,N_2914,N_2797);
nor U3247 (N_3247,N_2563,N_2908);
nor U3248 (N_3248,N_2974,N_2523);
xor U3249 (N_3249,N_2508,N_2545);
or U3250 (N_3250,N_2927,N_2973);
nand U3251 (N_3251,N_2501,N_2910);
nand U3252 (N_3252,N_2788,N_2502);
nand U3253 (N_3253,N_2664,N_2540);
and U3254 (N_3254,N_2675,N_2960);
and U3255 (N_3255,N_2589,N_2546);
nand U3256 (N_3256,N_2753,N_2659);
xnor U3257 (N_3257,N_2698,N_2964);
and U3258 (N_3258,N_2862,N_2995);
nand U3259 (N_3259,N_2961,N_2538);
and U3260 (N_3260,N_2871,N_2625);
and U3261 (N_3261,N_2675,N_2572);
nor U3262 (N_3262,N_2811,N_2693);
nand U3263 (N_3263,N_2703,N_2846);
or U3264 (N_3264,N_2844,N_2765);
and U3265 (N_3265,N_2612,N_2547);
or U3266 (N_3266,N_2767,N_2513);
nor U3267 (N_3267,N_2690,N_2915);
and U3268 (N_3268,N_2837,N_2674);
and U3269 (N_3269,N_2635,N_2579);
nand U3270 (N_3270,N_2710,N_2633);
or U3271 (N_3271,N_2681,N_2559);
nor U3272 (N_3272,N_2930,N_2745);
nor U3273 (N_3273,N_2918,N_2875);
nor U3274 (N_3274,N_2965,N_2973);
nor U3275 (N_3275,N_2581,N_2904);
or U3276 (N_3276,N_2934,N_2609);
or U3277 (N_3277,N_2855,N_2716);
nor U3278 (N_3278,N_2936,N_2649);
xor U3279 (N_3279,N_2715,N_2951);
nor U3280 (N_3280,N_2507,N_2707);
and U3281 (N_3281,N_2852,N_2727);
nand U3282 (N_3282,N_2945,N_2669);
or U3283 (N_3283,N_2752,N_2683);
or U3284 (N_3284,N_2650,N_2642);
and U3285 (N_3285,N_2852,N_2647);
nor U3286 (N_3286,N_2705,N_2633);
or U3287 (N_3287,N_2597,N_2817);
xnor U3288 (N_3288,N_2948,N_2597);
and U3289 (N_3289,N_2668,N_2986);
or U3290 (N_3290,N_2827,N_2738);
nand U3291 (N_3291,N_2893,N_2641);
or U3292 (N_3292,N_2878,N_2800);
nand U3293 (N_3293,N_2828,N_2545);
xnor U3294 (N_3294,N_2869,N_2794);
and U3295 (N_3295,N_2856,N_2527);
nor U3296 (N_3296,N_2647,N_2625);
and U3297 (N_3297,N_2805,N_2632);
or U3298 (N_3298,N_2964,N_2511);
nor U3299 (N_3299,N_2921,N_2722);
or U3300 (N_3300,N_2525,N_2941);
nor U3301 (N_3301,N_2557,N_2897);
nor U3302 (N_3302,N_2539,N_2977);
nand U3303 (N_3303,N_2838,N_2676);
and U3304 (N_3304,N_2851,N_2556);
or U3305 (N_3305,N_2990,N_2508);
nand U3306 (N_3306,N_2856,N_2553);
nor U3307 (N_3307,N_2769,N_2559);
and U3308 (N_3308,N_2939,N_2729);
nand U3309 (N_3309,N_2985,N_2663);
nor U3310 (N_3310,N_2502,N_2946);
nor U3311 (N_3311,N_2620,N_2807);
and U3312 (N_3312,N_2698,N_2803);
nand U3313 (N_3313,N_2810,N_2566);
or U3314 (N_3314,N_2783,N_2526);
nor U3315 (N_3315,N_2754,N_2512);
or U3316 (N_3316,N_2742,N_2895);
and U3317 (N_3317,N_2997,N_2868);
and U3318 (N_3318,N_2946,N_2971);
or U3319 (N_3319,N_2531,N_2938);
nor U3320 (N_3320,N_2722,N_2956);
nand U3321 (N_3321,N_2528,N_2566);
nor U3322 (N_3322,N_2564,N_2928);
or U3323 (N_3323,N_2913,N_2849);
nor U3324 (N_3324,N_2721,N_2562);
and U3325 (N_3325,N_2511,N_2819);
or U3326 (N_3326,N_2527,N_2624);
nand U3327 (N_3327,N_2697,N_2782);
or U3328 (N_3328,N_2883,N_2825);
nand U3329 (N_3329,N_2880,N_2741);
and U3330 (N_3330,N_2888,N_2889);
xor U3331 (N_3331,N_2994,N_2757);
nor U3332 (N_3332,N_2582,N_2574);
and U3333 (N_3333,N_2763,N_2608);
nor U3334 (N_3334,N_2903,N_2890);
and U3335 (N_3335,N_2793,N_2991);
nor U3336 (N_3336,N_2918,N_2806);
nand U3337 (N_3337,N_2985,N_2984);
nand U3338 (N_3338,N_2645,N_2526);
nor U3339 (N_3339,N_2657,N_2654);
nand U3340 (N_3340,N_2652,N_2848);
nor U3341 (N_3341,N_2519,N_2679);
and U3342 (N_3342,N_2871,N_2854);
and U3343 (N_3343,N_2626,N_2991);
or U3344 (N_3344,N_2529,N_2926);
or U3345 (N_3345,N_2897,N_2551);
or U3346 (N_3346,N_2693,N_2882);
nand U3347 (N_3347,N_2980,N_2789);
xnor U3348 (N_3348,N_2899,N_2949);
xnor U3349 (N_3349,N_2866,N_2654);
nand U3350 (N_3350,N_2912,N_2679);
or U3351 (N_3351,N_2911,N_2500);
nor U3352 (N_3352,N_2647,N_2991);
or U3353 (N_3353,N_2709,N_2935);
xnor U3354 (N_3354,N_2778,N_2651);
and U3355 (N_3355,N_2790,N_2723);
and U3356 (N_3356,N_2755,N_2734);
nand U3357 (N_3357,N_2940,N_2582);
nand U3358 (N_3358,N_2532,N_2519);
nand U3359 (N_3359,N_2542,N_2651);
nor U3360 (N_3360,N_2500,N_2964);
nand U3361 (N_3361,N_2969,N_2707);
nand U3362 (N_3362,N_2784,N_2612);
nand U3363 (N_3363,N_2523,N_2658);
nand U3364 (N_3364,N_2854,N_2754);
nand U3365 (N_3365,N_2991,N_2660);
or U3366 (N_3366,N_2739,N_2889);
or U3367 (N_3367,N_2621,N_2586);
and U3368 (N_3368,N_2645,N_2707);
nand U3369 (N_3369,N_2778,N_2856);
nand U3370 (N_3370,N_2853,N_2527);
and U3371 (N_3371,N_2585,N_2737);
or U3372 (N_3372,N_2765,N_2825);
and U3373 (N_3373,N_2610,N_2855);
or U3374 (N_3374,N_2840,N_2943);
and U3375 (N_3375,N_2768,N_2632);
nor U3376 (N_3376,N_2687,N_2558);
or U3377 (N_3377,N_2629,N_2532);
nand U3378 (N_3378,N_2524,N_2570);
or U3379 (N_3379,N_2736,N_2743);
or U3380 (N_3380,N_2921,N_2814);
and U3381 (N_3381,N_2550,N_2502);
nor U3382 (N_3382,N_2972,N_2668);
or U3383 (N_3383,N_2952,N_2659);
or U3384 (N_3384,N_2888,N_2976);
nand U3385 (N_3385,N_2720,N_2851);
nor U3386 (N_3386,N_2692,N_2787);
or U3387 (N_3387,N_2674,N_2629);
or U3388 (N_3388,N_2540,N_2546);
xor U3389 (N_3389,N_2799,N_2579);
or U3390 (N_3390,N_2996,N_2830);
and U3391 (N_3391,N_2793,N_2933);
and U3392 (N_3392,N_2882,N_2540);
or U3393 (N_3393,N_2543,N_2965);
nor U3394 (N_3394,N_2627,N_2566);
nor U3395 (N_3395,N_2602,N_2781);
nor U3396 (N_3396,N_2678,N_2857);
or U3397 (N_3397,N_2669,N_2685);
nor U3398 (N_3398,N_2791,N_2735);
nor U3399 (N_3399,N_2890,N_2928);
nand U3400 (N_3400,N_2503,N_2845);
nand U3401 (N_3401,N_2907,N_2991);
or U3402 (N_3402,N_2728,N_2621);
or U3403 (N_3403,N_2948,N_2755);
nor U3404 (N_3404,N_2707,N_2883);
and U3405 (N_3405,N_2911,N_2984);
or U3406 (N_3406,N_2755,N_2774);
nand U3407 (N_3407,N_2800,N_2996);
and U3408 (N_3408,N_2632,N_2985);
nand U3409 (N_3409,N_2864,N_2895);
nand U3410 (N_3410,N_2539,N_2545);
or U3411 (N_3411,N_2761,N_2833);
nor U3412 (N_3412,N_2886,N_2773);
or U3413 (N_3413,N_2828,N_2965);
nand U3414 (N_3414,N_2868,N_2882);
or U3415 (N_3415,N_2935,N_2515);
or U3416 (N_3416,N_2714,N_2834);
and U3417 (N_3417,N_2658,N_2960);
and U3418 (N_3418,N_2770,N_2564);
nand U3419 (N_3419,N_2975,N_2779);
or U3420 (N_3420,N_2874,N_2532);
or U3421 (N_3421,N_2853,N_2773);
or U3422 (N_3422,N_2714,N_2640);
nand U3423 (N_3423,N_2529,N_2647);
and U3424 (N_3424,N_2529,N_2934);
or U3425 (N_3425,N_2598,N_2926);
nand U3426 (N_3426,N_2588,N_2836);
nor U3427 (N_3427,N_2919,N_2549);
nand U3428 (N_3428,N_2743,N_2950);
or U3429 (N_3429,N_2840,N_2556);
or U3430 (N_3430,N_2504,N_2521);
nand U3431 (N_3431,N_2825,N_2774);
nand U3432 (N_3432,N_2941,N_2800);
nor U3433 (N_3433,N_2811,N_2662);
nand U3434 (N_3434,N_2947,N_2979);
nand U3435 (N_3435,N_2729,N_2739);
or U3436 (N_3436,N_2896,N_2512);
nand U3437 (N_3437,N_2547,N_2735);
nor U3438 (N_3438,N_2647,N_2865);
nor U3439 (N_3439,N_2878,N_2884);
nand U3440 (N_3440,N_2507,N_2988);
nor U3441 (N_3441,N_2941,N_2908);
xor U3442 (N_3442,N_2725,N_2557);
or U3443 (N_3443,N_2603,N_2723);
or U3444 (N_3444,N_2524,N_2779);
nor U3445 (N_3445,N_2939,N_2526);
and U3446 (N_3446,N_2523,N_2582);
and U3447 (N_3447,N_2826,N_2781);
nand U3448 (N_3448,N_2952,N_2801);
or U3449 (N_3449,N_2684,N_2829);
or U3450 (N_3450,N_2730,N_2570);
nand U3451 (N_3451,N_2639,N_2526);
nor U3452 (N_3452,N_2722,N_2946);
or U3453 (N_3453,N_2680,N_2744);
nor U3454 (N_3454,N_2917,N_2899);
and U3455 (N_3455,N_2505,N_2990);
and U3456 (N_3456,N_2642,N_2760);
nand U3457 (N_3457,N_2866,N_2886);
nand U3458 (N_3458,N_2909,N_2617);
nand U3459 (N_3459,N_2766,N_2524);
nand U3460 (N_3460,N_2787,N_2779);
nor U3461 (N_3461,N_2620,N_2729);
nand U3462 (N_3462,N_2788,N_2537);
or U3463 (N_3463,N_2578,N_2644);
and U3464 (N_3464,N_2595,N_2635);
nor U3465 (N_3465,N_2728,N_2798);
nor U3466 (N_3466,N_2731,N_2689);
and U3467 (N_3467,N_2605,N_2822);
and U3468 (N_3468,N_2672,N_2767);
nor U3469 (N_3469,N_2579,N_2973);
nand U3470 (N_3470,N_2997,N_2773);
and U3471 (N_3471,N_2819,N_2918);
and U3472 (N_3472,N_2817,N_2821);
nor U3473 (N_3473,N_2982,N_2711);
or U3474 (N_3474,N_2531,N_2930);
nor U3475 (N_3475,N_2815,N_2922);
or U3476 (N_3476,N_2653,N_2990);
nor U3477 (N_3477,N_2825,N_2588);
nand U3478 (N_3478,N_2558,N_2930);
or U3479 (N_3479,N_2775,N_2924);
nand U3480 (N_3480,N_2874,N_2903);
xor U3481 (N_3481,N_2805,N_2765);
nor U3482 (N_3482,N_2836,N_2674);
or U3483 (N_3483,N_2968,N_2763);
or U3484 (N_3484,N_2904,N_2582);
nor U3485 (N_3485,N_2732,N_2669);
or U3486 (N_3486,N_2687,N_2866);
nand U3487 (N_3487,N_2898,N_2561);
nor U3488 (N_3488,N_2885,N_2803);
nand U3489 (N_3489,N_2823,N_2929);
and U3490 (N_3490,N_2593,N_2764);
nand U3491 (N_3491,N_2570,N_2568);
or U3492 (N_3492,N_2873,N_2656);
nand U3493 (N_3493,N_2901,N_2688);
or U3494 (N_3494,N_2828,N_2623);
nand U3495 (N_3495,N_2685,N_2703);
or U3496 (N_3496,N_2506,N_2553);
xor U3497 (N_3497,N_2607,N_2544);
nor U3498 (N_3498,N_2607,N_2706);
or U3499 (N_3499,N_2694,N_2623);
or U3500 (N_3500,N_3357,N_3170);
nor U3501 (N_3501,N_3255,N_3020);
nand U3502 (N_3502,N_3189,N_3308);
nand U3503 (N_3503,N_3193,N_3346);
and U3504 (N_3504,N_3251,N_3479);
or U3505 (N_3505,N_3028,N_3235);
nand U3506 (N_3506,N_3403,N_3187);
and U3507 (N_3507,N_3067,N_3476);
nor U3508 (N_3508,N_3086,N_3448);
and U3509 (N_3509,N_3492,N_3405);
nand U3510 (N_3510,N_3000,N_3042);
nor U3511 (N_3511,N_3152,N_3425);
xor U3512 (N_3512,N_3485,N_3160);
and U3513 (N_3513,N_3444,N_3490);
and U3514 (N_3514,N_3175,N_3285);
or U3515 (N_3515,N_3385,N_3266);
nor U3516 (N_3516,N_3353,N_3267);
or U3517 (N_3517,N_3331,N_3096);
nand U3518 (N_3518,N_3103,N_3375);
or U3519 (N_3519,N_3198,N_3117);
nor U3520 (N_3520,N_3234,N_3363);
nand U3521 (N_3521,N_3345,N_3048);
or U3522 (N_3522,N_3219,N_3292);
nor U3523 (N_3523,N_3093,N_3128);
or U3524 (N_3524,N_3078,N_3462);
or U3525 (N_3525,N_3121,N_3194);
nand U3526 (N_3526,N_3108,N_3314);
nor U3527 (N_3527,N_3423,N_3428);
nor U3528 (N_3528,N_3356,N_3342);
xor U3529 (N_3529,N_3228,N_3414);
or U3530 (N_3530,N_3461,N_3062);
nand U3531 (N_3531,N_3070,N_3066);
or U3532 (N_3532,N_3333,N_3144);
or U3533 (N_3533,N_3147,N_3489);
nor U3534 (N_3534,N_3404,N_3418);
nor U3535 (N_3535,N_3413,N_3008);
nor U3536 (N_3536,N_3453,N_3268);
and U3537 (N_3537,N_3374,N_3452);
nand U3538 (N_3538,N_3010,N_3214);
nor U3539 (N_3539,N_3229,N_3386);
nand U3540 (N_3540,N_3191,N_3242);
or U3541 (N_3541,N_3208,N_3347);
nor U3542 (N_3542,N_3141,N_3301);
or U3543 (N_3543,N_3222,N_3341);
or U3544 (N_3544,N_3315,N_3409);
nand U3545 (N_3545,N_3188,N_3303);
nand U3546 (N_3546,N_3282,N_3220);
or U3547 (N_3547,N_3233,N_3468);
nand U3548 (N_3548,N_3149,N_3159);
or U3549 (N_3549,N_3259,N_3287);
nor U3550 (N_3550,N_3125,N_3090);
or U3551 (N_3551,N_3081,N_3394);
nand U3552 (N_3552,N_3202,N_3161);
or U3553 (N_3553,N_3158,N_3100);
nor U3554 (N_3554,N_3408,N_3289);
xnor U3555 (N_3555,N_3249,N_3092);
or U3556 (N_3556,N_3169,N_3022);
nand U3557 (N_3557,N_3465,N_3098);
nor U3558 (N_3558,N_3024,N_3046);
nand U3559 (N_3559,N_3358,N_3480);
nand U3560 (N_3560,N_3009,N_3215);
nand U3561 (N_3561,N_3364,N_3398);
nor U3562 (N_3562,N_3354,N_3377);
and U3563 (N_3563,N_3304,N_3473);
xnor U3564 (N_3564,N_3486,N_3260);
and U3565 (N_3565,N_3148,N_3069);
nand U3566 (N_3566,N_3439,N_3097);
nand U3567 (N_3567,N_3043,N_3326);
or U3568 (N_3568,N_3184,N_3372);
nor U3569 (N_3569,N_3004,N_3278);
nand U3570 (N_3570,N_3178,N_3309);
nor U3571 (N_3571,N_3477,N_3102);
nor U3572 (N_3572,N_3002,N_3467);
xor U3573 (N_3573,N_3493,N_3094);
and U3574 (N_3574,N_3054,N_3416);
or U3575 (N_3575,N_3114,N_3167);
nor U3576 (N_3576,N_3052,N_3401);
or U3577 (N_3577,N_3018,N_3129);
and U3578 (N_3578,N_3196,N_3120);
and U3579 (N_3579,N_3231,N_3343);
and U3580 (N_3580,N_3006,N_3300);
or U3581 (N_3581,N_3154,N_3387);
nand U3582 (N_3582,N_3362,N_3424);
nor U3583 (N_3583,N_3080,N_3012);
or U3584 (N_3584,N_3302,N_3321);
nor U3585 (N_3585,N_3361,N_3082);
nand U3586 (N_3586,N_3256,N_3051);
nor U3587 (N_3587,N_3047,N_3407);
or U3588 (N_3588,N_3174,N_3327);
nand U3589 (N_3589,N_3436,N_3366);
nand U3590 (N_3590,N_3291,N_3232);
nand U3591 (N_3591,N_3437,N_3324);
and U3592 (N_3592,N_3258,N_3293);
xnor U3593 (N_3593,N_3201,N_3388);
nor U3594 (N_3594,N_3262,N_3107);
or U3595 (N_3595,N_3145,N_3296);
and U3596 (N_3596,N_3335,N_3030);
or U3597 (N_3597,N_3495,N_3143);
or U3598 (N_3598,N_3338,N_3063);
or U3599 (N_3599,N_3137,N_3118);
and U3600 (N_3600,N_3195,N_3084);
nand U3601 (N_3601,N_3391,N_3435);
or U3602 (N_3602,N_3433,N_3494);
nand U3603 (N_3603,N_3491,N_3384);
nand U3604 (N_3604,N_3019,N_3325);
nor U3605 (N_3605,N_3471,N_3180);
or U3606 (N_3606,N_3487,N_3127);
nor U3607 (N_3607,N_3101,N_3211);
nor U3608 (N_3608,N_3199,N_3206);
nand U3609 (N_3609,N_3172,N_3420);
or U3610 (N_3610,N_3334,N_3163);
and U3611 (N_3611,N_3038,N_3183);
and U3612 (N_3612,N_3350,N_3085);
nor U3613 (N_3613,N_3115,N_3273);
nor U3614 (N_3614,N_3369,N_3298);
or U3615 (N_3615,N_3091,N_3438);
nand U3616 (N_3616,N_3079,N_3365);
and U3617 (N_3617,N_3498,N_3056);
nor U3618 (N_3618,N_3213,N_3087);
nand U3619 (N_3619,N_3227,N_3105);
or U3620 (N_3620,N_3089,N_3319);
or U3621 (N_3621,N_3045,N_3252);
nand U3622 (N_3622,N_3032,N_3253);
nor U3623 (N_3623,N_3224,N_3328);
nand U3624 (N_3624,N_3445,N_3257);
or U3625 (N_3625,N_3277,N_3254);
and U3626 (N_3626,N_3075,N_3162);
nand U3627 (N_3627,N_3349,N_3431);
nor U3628 (N_3628,N_3049,N_3432);
nor U3629 (N_3629,N_3496,N_3223);
nand U3630 (N_3630,N_3015,N_3441);
xor U3631 (N_3631,N_3068,N_3122);
or U3632 (N_3632,N_3400,N_3332);
or U3633 (N_3633,N_3368,N_3171);
or U3634 (N_3634,N_3322,N_3352);
nor U3635 (N_3635,N_3135,N_3442);
nand U3636 (N_3636,N_3157,N_3204);
and U3637 (N_3637,N_3458,N_3339);
xnor U3638 (N_3638,N_3410,N_3397);
or U3639 (N_3639,N_3455,N_3497);
nand U3640 (N_3640,N_3113,N_3310);
and U3641 (N_3641,N_3168,N_3123);
or U3642 (N_3642,N_3451,N_3212);
nand U3643 (N_3643,N_3316,N_3399);
or U3644 (N_3644,N_3481,N_3271);
nor U3645 (N_3645,N_3381,N_3041);
or U3646 (N_3646,N_3280,N_3336);
or U3647 (N_3647,N_3389,N_3126);
or U3648 (N_3648,N_3313,N_3340);
nand U3649 (N_3649,N_3053,N_3348);
nor U3650 (N_3650,N_3272,N_3274);
and U3651 (N_3651,N_3449,N_3402);
nor U3652 (N_3652,N_3360,N_3155);
nand U3653 (N_3653,N_3236,N_3151);
or U3654 (N_3654,N_3474,N_3482);
and U3655 (N_3655,N_3412,N_3221);
or U3656 (N_3656,N_3165,N_3294);
and U3657 (N_3657,N_3112,N_3083);
or U3658 (N_3658,N_3380,N_3475);
nand U3659 (N_3659,N_3025,N_3031);
nor U3660 (N_3660,N_3237,N_3001);
or U3661 (N_3661,N_3469,N_3246);
or U3662 (N_3662,N_3430,N_3422);
nor U3663 (N_3663,N_3176,N_3472);
and U3664 (N_3664,N_3337,N_3139);
nor U3665 (N_3665,N_3446,N_3150);
or U3666 (N_3666,N_3460,N_3059);
nor U3667 (N_3667,N_3205,N_3450);
and U3668 (N_3668,N_3440,N_3421);
xor U3669 (N_3669,N_3110,N_3265);
and U3670 (N_3670,N_3013,N_3396);
or U3671 (N_3671,N_3393,N_3478);
nor U3672 (N_3672,N_3383,N_3415);
or U3673 (N_3673,N_3134,N_3027);
or U3674 (N_3674,N_3014,N_3177);
nand U3675 (N_3675,N_3029,N_3136);
nor U3676 (N_3676,N_3036,N_3317);
or U3677 (N_3677,N_3099,N_3207);
nand U3678 (N_3678,N_3104,N_3005);
nand U3679 (N_3679,N_3179,N_3153);
or U3680 (N_3680,N_3464,N_3146);
or U3681 (N_3681,N_3359,N_3297);
or U3682 (N_3682,N_3210,N_3240);
or U3683 (N_3683,N_3016,N_3131);
and U3684 (N_3684,N_3484,N_3351);
nand U3685 (N_3685,N_3065,N_3017);
nor U3686 (N_3686,N_3261,N_3499);
nand U3687 (N_3687,N_3044,N_3088);
nor U3688 (N_3688,N_3230,N_3058);
nor U3689 (N_3689,N_3248,N_3281);
and U3690 (N_3690,N_3329,N_3186);
or U3691 (N_3691,N_3488,N_3138);
nor U3692 (N_3692,N_3344,N_3071);
nand U3693 (N_3693,N_3459,N_3197);
nand U3694 (N_3694,N_3367,N_3320);
or U3695 (N_3695,N_3132,N_3390);
or U3696 (N_3696,N_3106,N_3284);
nand U3697 (N_3697,N_3037,N_3454);
nor U3698 (N_3698,N_3306,N_3241);
nor U3699 (N_3699,N_3318,N_3406);
nor U3700 (N_3700,N_3033,N_3263);
or U3701 (N_3701,N_3243,N_3039);
and U3702 (N_3702,N_3130,N_3264);
nand U3703 (N_3703,N_3111,N_3239);
nor U3704 (N_3704,N_3003,N_3164);
nand U3705 (N_3705,N_3192,N_3182);
nor U3706 (N_3706,N_3483,N_3463);
and U3707 (N_3707,N_3076,N_3305);
or U3708 (N_3708,N_3269,N_3200);
or U3709 (N_3709,N_3295,N_3392);
or U3710 (N_3710,N_3209,N_3077);
xnor U3711 (N_3711,N_3156,N_3119);
or U3712 (N_3712,N_3311,N_3288);
and U3713 (N_3713,N_3074,N_3286);
nor U3714 (N_3714,N_3244,N_3116);
and U3715 (N_3715,N_3378,N_3216);
nand U3716 (N_3716,N_3011,N_3140);
nand U3717 (N_3717,N_3419,N_3190);
nand U3718 (N_3718,N_3142,N_3427);
and U3719 (N_3719,N_3443,N_3040);
nor U3720 (N_3720,N_3095,N_3064);
nand U3721 (N_3721,N_3370,N_3371);
nor U3722 (N_3722,N_3376,N_3447);
nand U3723 (N_3723,N_3417,N_3456);
nor U3724 (N_3724,N_3270,N_3250);
nor U3725 (N_3725,N_3133,N_3073);
nor U3726 (N_3726,N_3035,N_3023);
or U3727 (N_3727,N_3021,N_3060);
xor U3728 (N_3728,N_3457,N_3247);
nor U3729 (N_3729,N_3061,N_3217);
xor U3730 (N_3730,N_3290,N_3185);
and U3731 (N_3731,N_3109,N_3166);
or U3732 (N_3732,N_3373,N_3072);
and U3733 (N_3733,N_3429,N_3203);
and U3734 (N_3734,N_3379,N_3279);
or U3735 (N_3735,N_3330,N_3218);
and U3736 (N_3736,N_3238,N_3466);
and U3737 (N_3737,N_3323,N_3055);
or U3738 (N_3738,N_3276,N_3057);
nor U3739 (N_3739,N_3173,N_3050);
nand U3740 (N_3740,N_3275,N_3226);
nor U3741 (N_3741,N_3007,N_3312);
nor U3742 (N_3742,N_3181,N_3395);
or U3743 (N_3743,N_3434,N_3124);
or U3744 (N_3744,N_3283,N_3034);
nor U3745 (N_3745,N_3245,N_3225);
xor U3746 (N_3746,N_3026,N_3426);
nor U3747 (N_3747,N_3470,N_3382);
nand U3748 (N_3748,N_3355,N_3307);
or U3749 (N_3749,N_3411,N_3299);
nand U3750 (N_3750,N_3109,N_3139);
nand U3751 (N_3751,N_3340,N_3117);
nor U3752 (N_3752,N_3352,N_3365);
and U3753 (N_3753,N_3387,N_3356);
or U3754 (N_3754,N_3452,N_3486);
nor U3755 (N_3755,N_3005,N_3361);
nor U3756 (N_3756,N_3224,N_3062);
nand U3757 (N_3757,N_3306,N_3152);
or U3758 (N_3758,N_3011,N_3473);
and U3759 (N_3759,N_3429,N_3149);
or U3760 (N_3760,N_3004,N_3141);
and U3761 (N_3761,N_3396,N_3129);
or U3762 (N_3762,N_3190,N_3427);
or U3763 (N_3763,N_3206,N_3400);
and U3764 (N_3764,N_3465,N_3270);
nand U3765 (N_3765,N_3400,N_3016);
nor U3766 (N_3766,N_3138,N_3255);
or U3767 (N_3767,N_3394,N_3369);
nand U3768 (N_3768,N_3464,N_3411);
and U3769 (N_3769,N_3235,N_3452);
or U3770 (N_3770,N_3144,N_3350);
nand U3771 (N_3771,N_3335,N_3140);
or U3772 (N_3772,N_3311,N_3313);
nor U3773 (N_3773,N_3239,N_3292);
nor U3774 (N_3774,N_3038,N_3075);
and U3775 (N_3775,N_3216,N_3388);
nand U3776 (N_3776,N_3351,N_3237);
and U3777 (N_3777,N_3403,N_3428);
nor U3778 (N_3778,N_3135,N_3068);
nand U3779 (N_3779,N_3397,N_3482);
nand U3780 (N_3780,N_3263,N_3206);
nand U3781 (N_3781,N_3060,N_3467);
or U3782 (N_3782,N_3339,N_3259);
and U3783 (N_3783,N_3371,N_3018);
nand U3784 (N_3784,N_3071,N_3222);
nor U3785 (N_3785,N_3095,N_3061);
nand U3786 (N_3786,N_3003,N_3419);
nor U3787 (N_3787,N_3215,N_3318);
nor U3788 (N_3788,N_3419,N_3273);
nor U3789 (N_3789,N_3140,N_3002);
or U3790 (N_3790,N_3021,N_3002);
nand U3791 (N_3791,N_3110,N_3257);
or U3792 (N_3792,N_3048,N_3410);
nand U3793 (N_3793,N_3033,N_3253);
and U3794 (N_3794,N_3081,N_3123);
or U3795 (N_3795,N_3218,N_3257);
and U3796 (N_3796,N_3292,N_3486);
and U3797 (N_3797,N_3465,N_3427);
nand U3798 (N_3798,N_3384,N_3123);
nor U3799 (N_3799,N_3456,N_3309);
and U3800 (N_3800,N_3286,N_3136);
nand U3801 (N_3801,N_3049,N_3214);
nor U3802 (N_3802,N_3126,N_3299);
nor U3803 (N_3803,N_3489,N_3224);
nand U3804 (N_3804,N_3429,N_3137);
and U3805 (N_3805,N_3418,N_3300);
and U3806 (N_3806,N_3447,N_3275);
nand U3807 (N_3807,N_3017,N_3422);
nand U3808 (N_3808,N_3371,N_3350);
or U3809 (N_3809,N_3122,N_3268);
or U3810 (N_3810,N_3104,N_3313);
nor U3811 (N_3811,N_3115,N_3493);
nand U3812 (N_3812,N_3107,N_3130);
nand U3813 (N_3813,N_3441,N_3147);
and U3814 (N_3814,N_3430,N_3416);
nor U3815 (N_3815,N_3282,N_3406);
nor U3816 (N_3816,N_3054,N_3477);
nand U3817 (N_3817,N_3340,N_3301);
nand U3818 (N_3818,N_3223,N_3209);
or U3819 (N_3819,N_3460,N_3448);
nand U3820 (N_3820,N_3053,N_3280);
xor U3821 (N_3821,N_3330,N_3364);
and U3822 (N_3822,N_3401,N_3090);
nor U3823 (N_3823,N_3096,N_3456);
and U3824 (N_3824,N_3210,N_3186);
and U3825 (N_3825,N_3208,N_3265);
nor U3826 (N_3826,N_3090,N_3240);
nand U3827 (N_3827,N_3454,N_3387);
and U3828 (N_3828,N_3406,N_3175);
nand U3829 (N_3829,N_3095,N_3126);
or U3830 (N_3830,N_3443,N_3103);
nor U3831 (N_3831,N_3349,N_3015);
nor U3832 (N_3832,N_3294,N_3490);
nor U3833 (N_3833,N_3396,N_3429);
nor U3834 (N_3834,N_3106,N_3214);
and U3835 (N_3835,N_3448,N_3300);
and U3836 (N_3836,N_3361,N_3184);
or U3837 (N_3837,N_3109,N_3185);
or U3838 (N_3838,N_3056,N_3476);
nor U3839 (N_3839,N_3201,N_3005);
nor U3840 (N_3840,N_3436,N_3194);
or U3841 (N_3841,N_3132,N_3011);
and U3842 (N_3842,N_3087,N_3341);
or U3843 (N_3843,N_3307,N_3101);
and U3844 (N_3844,N_3099,N_3033);
xnor U3845 (N_3845,N_3435,N_3021);
nor U3846 (N_3846,N_3186,N_3314);
nor U3847 (N_3847,N_3216,N_3026);
nand U3848 (N_3848,N_3432,N_3442);
and U3849 (N_3849,N_3108,N_3420);
nand U3850 (N_3850,N_3037,N_3443);
nor U3851 (N_3851,N_3064,N_3013);
xnor U3852 (N_3852,N_3208,N_3337);
nand U3853 (N_3853,N_3220,N_3440);
or U3854 (N_3854,N_3479,N_3191);
and U3855 (N_3855,N_3305,N_3318);
nor U3856 (N_3856,N_3279,N_3237);
and U3857 (N_3857,N_3142,N_3308);
nor U3858 (N_3858,N_3067,N_3023);
nor U3859 (N_3859,N_3400,N_3277);
or U3860 (N_3860,N_3169,N_3080);
or U3861 (N_3861,N_3213,N_3334);
nand U3862 (N_3862,N_3057,N_3412);
xor U3863 (N_3863,N_3086,N_3461);
and U3864 (N_3864,N_3333,N_3014);
and U3865 (N_3865,N_3481,N_3131);
nand U3866 (N_3866,N_3410,N_3377);
and U3867 (N_3867,N_3275,N_3311);
and U3868 (N_3868,N_3396,N_3376);
and U3869 (N_3869,N_3485,N_3116);
or U3870 (N_3870,N_3112,N_3290);
or U3871 (N_3871,N_3366,N_3274);
or U3872 (N_3872,N_3475,N_3353);
or U3873 (N_3873,N_3437,N_3179);
nand U3874 (N_3874,N_3276,N_3060);
xnor U3875 (N_3875,N_3086,N_3480);
nand U3876 (N_3876,N_3219,N_3427);
and U3877 (N_3877,N_3341,N_3057);
and U3878 (N_3878,N_3017,N_3048);
nor U3879 (N_3879,N_3300,N_3394);
nor U3880 (N_3880,N_3087,N_3115);
and U3881 (N_3881,N_3052,N_3031);
nor U3882 (N_3882,N_3119,N_3234);
nand U3883 (N_3883,N_3396,N_3062);
and U3884 (N_3884,N_3437,N_3425);
or U3885 (N_3885,N_3313,N_3417);
and U3886 (N_3886,N_3443,N_3057);
and U3887 (N_3887,N_3021,N_3388);
and U3888 (N_3888,N_3481,N_3374);
nor U3889 (N_3889,N_3038,N_3005);
nand U3890 (N_3890,N_3149,N_3009);
or U3891 (N_3891,N_3029,N_3293);
nand U3892 (N_3892,N_3328,N_3341);
nor U3893 (N_3893,N_3098,N_3118);
xor U3894 (N_3894,N_3197,N_3021);
nand U3895 (N_3895,N_3399,N_3059);
nor U3896 (N_3896,N_3125,N_3044);
and U3897 (N_3897,N_3407,N_3410);
nor U3898 (N_3898,N_3074,N_3072);
or U3899 (N_3899,N_3169,N_3037);
or U3900 (N_3900,N_3085,N_3300);
and U3901 (N_3901,N_3262,N_3159);
nor U3902 (N_3902,N_3323,N_3202);
and U3903 (N_3903,N_3463,N_3180);
nand U3904 (N_3904,N_3072,N_3289);
or U3905 (N_3905,N_3225,N_3439);
and U3906 (N_3906,N_3120,N_3117);
nand U3907 (N_3907,N_3260,N_3448);
and U3908 (N_3908,N_3150,N_3363);
and U3909 (N_3909,N_3361,N_3344);
or U3910 (N_3910,N_3143,N_3225);
or U3911 (N_3911,N_3404,N_3334);
nor U3912 (N_3912,N_3157,N_3063);
nand U3913 (N_3913,N_3425,N_3179);
nor U3914 (N_3914,N_3080,N_3282);
nand U3915 (N_3915,N_3073,N_3013);
and U3916 (N_3916,N_3344,N_3260);
nor U3917 (N_3917,N_3151,N_3398);
nand U3918 (N_3918,N_3175,N_3090);
and U3919 (N_3919,N_3446,N_3314);
and U3920 (N_3920,N_3190,N_3377);
or U3921 (N_3921,N_3174,N_3160);
and U3922 (N_3922,N_3202,N_3263);
nor U3923 (N_3923,N_3286,N_3176);
nand U3924 (N_3924,N_3099,N_3172);
and U3925 (N_3925,N_3189,N_3096);
and U3926 (N_3926,N_3498,N_3442);
and U3927 (N_3927,N_3326,N_3170);
nor U3928 (N_3928,N_3471,N_3171);
nand U3929 (N_3929,N_3422,N_3074);
xor U3930 (N_3930,N_3013,N_3279);
and U3931 (N_3931,N_3182,N_3482);
nand U3932 (N_3932,N_3151,N_3187);
and U3933 (N_3933,N_3287,N_3106);
and U3934 (N_3934,N_3232,N_3190);
and U3935 (N_3935,N_3236,N_3429);
nor U3936 (N_3936,N_3314,N_3209);
and U3937 (N_3937,N_3128,N_3064);
nor U3938 (N_3938,N_3252,N_3161);
nor U3939 (N_3939,N_3090,N_3305);
and U3940 (N_3940,N_3169,N_3067);
nand U3941 (N_3941,N_3001,N_3373);
or U3942 (N_3942,N_3282,N_3217);
or U3943 (N_3943,N_3049,N_3320);
nand U3944 (N_3944,N_3144,N_3222);
nor U3945 (N_3945,N_3184,N_3054);
or U3946 (N_3946,N_3085,N_3488);
nor U3947 (N_3947,N_3273,N_3127);
and U3948 (N_3948,N_3314,N_3432);
and U3949 (N_3949,N_3179,N_3329);
or U3950 (N_3950,N_3319,N_3463);
nor U3951 (N_3951,N_3309,N_3175);
or U3952 (N_3952,N_3040,N_3129);
nand U3953 (N_3953,N_3468,N_3302);
nor U3954 (N_3954,N_3069,N_3039);
or U3955 (N_3955,N_3002,N_3213);
nor U3956 (N_3956,N_3400,N_3185);
and U3957 (N_3957,N_3131,N_3249);
nand U3958 (N_3958,N_3269,N_3084);
and U3959 (N_3959,N_3219,N_3061);
and U3960 (N_3960,N_3078,N_3438);
and U3961 (N_3961,N_3291,N_3410);
nor U3962 (N_3962,N_3314,N_3220);
or U3963 (N_3963,N_3183,N_3410);
and U3964 (N_3964,N_3153,N_3357);
xnor U3965 (N_3965,N_3265,N_3045);
nor U3966 (N_3966,N_3371,N_3424);
or U3967 (N_3967,N_3046,N_3402);
nor U3968 (N_3968,N_3011,N_3100);
and U3969 (N_3969,N_3476,N_3022);
or U3970 (N_3970,N_3341,N_3299);
nand U3971 (N_3971,N_3104,N_3122);
or U3972 (N_3972,N_3384,N_3416);
nor U3973 (N_3973,N_3267,N_3496);
nor U3974 (N_3974,N_3189,N_3405);
nand U3975 (N_3975,N_3000,N_3204);
nor U3976 (N_3976,N_3453,N_3415);
or U3977 (N_3977,N_3255,N_3150);
or U3978 (N_3978,N_3206,N_3100);
or U3979 (N_3979,N_3181,N_3001);
nor U3980 (N_3980,N_3002,N_3248);
or U3981 (N_3981,N_3135,N_3186);
nand U3982 (N_3982,N_3294,N_3138);
and U3983 (N_3983,N_3078,N_3205);
xnor U3984 (N_3984,N_3021,N_3097);
and U3985 (N_3985,N_3128,N_3120);
and U3986 (N_3986,N_3141,N_3045);
and U3987 (N_3987,N_3439,N_3155);
and U3988 (N_3988,N_3132,N_3091);
or U3989 (N_3989,N_3408,N_3077);
nand U3990 (N_3990,N_3022,N_3378);
nand U3991 (N_3991,N_3091,N_3106);
nand U3992 (N_3992,N_3254,N_3175);
nand U3993 (N_3993,N_3141,N_3247);
nor U3994 (N_3994,N_3271,N_3069);
and U3995 (N_3995,N_3077,N_3230);
or U3996 (N_3996,N_3459,N_3335);
and U3997 (N_3997,N_3491,N_3073);
or U3998 (N_3998,N_3120,N_3123);
or U3999 (N_3999,N_3411,N_3338);
nor U4000 (N_4000,N_3668,N_3508);
nor U4001 (N_4001,N_3927,N_3566);
nor U4002 (N_4002,N_3999,N_3857);
or U4003 (N_4003,N_3829,N_3963);
or U4004 (N_4004,N_3997,N_3686);
or U4005 (N_4005,N_3856,N_3659);
nor U4006 (N_4006,N_3626,N_3915);
xnor U4007 (N_4007,N_3894,N_3802);
nor U4008 (N_4008,N_3582,N_3913);
nand U4009 (N_4009,N_3684,N_3959);
or U4010 (N_4010,N_3890,N_3561);
and U4011 (N_4011,N_3767,N_3682);
nand U4012 (N_4012,N_3575,N_3747);
and U4013 (N_4013,N_3733,N_3522);
nand U4014 (N_4014,N_3955,N_3661);
nor U4015 (N_4015,N_3641,N_3712);
and U4016 (N_4016,N_3681,N_3614);
nor U4017 (N_4017,N_3655,N_3899);
or U4018 (N_4018,N_3618,N_3987);
or U4019 (N_4019,N_3644,N_3720);
or U4020 (N_4020,N_3816,N_3678);
nand U4021 (N_4021,N_3893,N_3706);
and U4022 (N_4022,N_3810,N_3625);
nor U4023 (N_4023,N_3578,N_3705);
and U4024 (N_4024,N_3576,N_3945);
nor U4025 (N_4025,N_3635,N_3548);
nand U4026 (N_4026,N_3710,N_3600);
nor U4027 (N_4027,N_3836,N_3536);
nand U4028 (N_4028,N_3962,N_3629);
nand U4029 (N_4029,N_3845,N_3778);
nor U4030 (N_4030,N_3921,N_3691);
nand U4031 (N_4031,N_3617,N_3695);
or U4032 (N_4032,N_3862,N_3953);
or U4033 (N_4033,N_3771,N_3672);
and U4034 (N_4034,N_3872,N_3773);
or U4035 (N_4035,N_3852,N_3537);
nor U4036 (N_4036,N_3571,N_3774);
nand U4037 (N_4037,N_3886,N_3685);
nor U4038 (N_4038,N_3850,N_3606);
and U4039 (N_4039,N_3723,N_3966);
or U4040 (N_4040,N_3881,N_3725);
or U4041 (N_4041,N_3879,N_3669);
nand U4042 (N_4042,N_3823,N_3734);
nor U4043 (N_4043,N_3524,N_3516);
and U4044 (N_4044,N_3506,N_3671);
nand U4045 (N_4045,N_3935,N_3752);
or U4046 (N_4046,N_3923,N_3533);
nand U4047 (N_4047,N_3636,N_3517);
and U4048 (N_4048,N_3621,N_3787);
or U4049 (N_4049,N_3589,N_3758);
nor U4050 (N_4050,N_3924,N_3643);
or U4051 (N_4051,N_3690,N_3878);
and U4052 (N_4052,N_3901,N_3854);
and U4053 (N_4053,N_3900,N_3860);
nand U4054 (N_4054,N_3974,N_3992);
nor U4055 (N_4055,N_3883,N_3592);
nor U4056 (N_4056,N_3744,N_3870);
or U4057 (N_4057,N_3528,N_3590);
nor U4058 (N_4058,N_3531,N_3847);
nor U4059 (N_4059,N_3970,N_3545);
and U4060 (N_4060,N_3735,N_3568);
nor U4061 (N_4061,N_3912,N_3563);
nor U4062 (N_4062,N_3888,N_3613);
nand U4063 (N_4063,N_3967,N_3965);
nand U4064 (N_4064,N_3941,N_3689);
nor U4065 (N_4065,N_3952,N_3549);
nor U4066 (N_4066,N_3944,N_3801);
and U4067 (N_4067,N_3832,N_3835);
nand U4068 (N_4068,N_3708,N_3718);
nand U4069 (N_4069,N_3687,N_3793);
and U4070 (N_4070,N_3866,N_3756);
xor U4071 (N_4071,N_3510,N_3607);
and U4072 (N_4072,N_3822,N_3925);
and U4073 (N_4073,N_3650,N_3514);
nand U4074 (N_4074,N_3849,N_3831);
nor U4075 (N_4075,N_3784,N_3954);
and U4076 (N_4076,N_3791,N_3730);
nor U4077 (N_4077,N_3694,N_3633);
nor U4078 (N_4078,N_3620,N_3931);
and U4079 (N_4079,N_3885,N_3754);
and U4080 (N_4080,N_3585,N_3868);
nor U4081 (N_4081,N_3760,N_3581);
or U4082 (N_4082,N_3875,N_3554);
nand U4083 (N_4083,N_3765,N_3601);
and U4084 (N_4084,N_3977,N_3948);
and U4085 (N_4085,N_3707,N_3658);
and U4086 (N_4086,N_3530,N_3846);
and U4087 (N_4087,N_3559,N_3859);
and U4088 (N_4088,N_3930,N_3666);
and U4089 (N_4089,N_3587,N_3887);
nand U4090 (N_4090,N_3824,N_3975);
nor U4091 (N_4091,N_3942,N_3813);
nor U4092 (N_4092,N_3664,N_3610);
nor U4093 (N_4093,N_3830,N_3500);
or U4094 (N_4094,N_3919,N_3764);
nor U4095 (N_4095,N_3855,N_3892);
nor U4096 (N_4096,N_3978,N_3591);
nand U4097 (N_4097,N_3586,N_3947);
and U4098 (N_4098,N_3603,N_3909);
nor U4099 (N_4099,N_3827,N_3688);
nor U4100 (N_4100,N_3848,N_3969);
nor U4101 (N_4101,N_3539,N_3740);
nor U4102 (N_4102,N_3692,N_3837);
and U4103 (N_4103,N_3529,N_3809);
nand U4104 (N_4104,N_3958,N_3526);
and U4105 (N_4105,N_3918,N_3577);
or U4106 (N_4106,N_3991,N_3745);
nand U4107 (N_4107,N_3680,N_3535);
nor U4108 (N_4108,N_3786,N_3615);
nand U4109 (N_4109,N_3709,N_3818);
or U4110 (N_4110,N_3632,N_3768);
and U4111 (N_4111,N_3906,N_3917);
nor U4112 (N_4112,N_3739,N_3979);
nor U4113 (N_4113,N_3724,N_3657);
nor U4114 (N_4114,N_3637,N_3843);
nand U4115 (N_4115,N_3731,N_3891);
and U4116 (N_4116,N_3544,N_3904);
xor U4117 (N_4117,N_3513,N_3776);
and U4118 (N_4118,N_3540,N_3598);
nand U4119 (N_4119,N_3588,N_3616);
nor U4120 (N_4120,N_3871,N_3792);
xnor U4121 (N_4121,N_3634,N_3895);
and U4122 (N_4122,N_3583,N_3567);
or U4123 (N_4123,N_3701,N_3580);
nor U4124 (N_4124,N_3509,N_3574);
nor U4125 (N_4125,N_3700,N_3926);
nor U4126 (N_4126,N_3933,N_3702);
and U4127 (N_4127,N_3646,N_3570);
and U4128 (N_4128,N_3749,N_3806);
or U4129 (N_4129,N_3884,N_3649);
nor U4130 (N_4130,N_3775,N_3897);
nor U4131 (N_4131,N_3814,N_3565);
nor U4132 (N_4132,N_3647,N_3815);
or U4133 (N_4133,N_3799,N_3914);
or U4134 (N_4134,N_3717,N_3555);
or U4135 (N_4135,N_3782,N_3766);
and U4136 (N_4136,N_3622,N_3770);
nor U4137 (N_4137,N_3783,N_3863);
and U4138 (N_4138,N_3777,N_3715);
nand U4139 (N_4139,N_3907,N_3826);
nand U4140 (N_4140,N_3676,N_3785);
or U4141 (N_4141,N_3796,N_3867);
and U4142 (N_4142,N_3989,N_3800);
and U4143 (N_4143,N_3572,N_3932);
or U4144 (N_4144,N_3543,N_3980);
nor U4145 (N_4145,N_3627,N_3609);
nand U4146 (N_4146,N_3780,N_3808);
nand U4147 (N_4147,N_3515,N_3504);
or U4148 (N_4148,N_3821,N_3518);
nor U4149 (N_4149,N_3556,N_3828);
or U4150 (N_4150,N_3812,N_3679);
and U4151 (N_4151,N_3584,N_3746);
nor U4152 (N_4152,N_3753,N_3865);
or U4153 (N_4153,N_3699,N_3726);
xor U4154 (N_4154,N_3790,N_3788);
nor U4155 (N_4155,N_3558,N_3950);
nor U4156 (N_4156,N_3769,N_3599);
xor U4157 (N_4157,N_3505,N_3928);
nor U4158 (N_4158,N_3520,N_3990);
nand U4159 (N_4159,N_3527,N_3663);
and U4160 (N_4160,N_3961,N_3779);
nor U4161 (N_4161,N_3825,N_3569);
and U4162 (N_4162,N_3939,N_3631);
or U4163 (N_4163,N_3971,N_3525);
nand U4164 (N_4164,N_3596,N_3721);
and U4165 (N_4165,N_3946,N_3757);
nand U4166 (N_4166,N_3630,N_3929);
and U4167 (N_4167,N_3562,N_3956);
or U4168 (N_4168,N_3738,N_3957);
nor U4169 (N_4169,N_3984,N_3640);
or U4170 (N_4170,N_3960,N_3993);
xnor U4171 (N_4171,N_3716,N_3869);
and U4172 (N_4172,N_3507,N_3998);
nor U4173 (N_4173,N_3604,N_3882);
and U4174 (N_4174,N_3936,N_3789);
and U4175 (N_4175,N_3541,N_3665);
nor U4176 (N_4176,N_3732,N_3523);
nand U4177 (N_4177,N_3645,N_3713);
and U4178 (N_4178,N_3841,N_3602);
nor U4179 (N_4179,N_3711,N_3943);
nor U4180 (N_4180,N_3593,N_3803);
nor U4181 (N_4181,N_3542,N_3864);
nor U4182 (N_4182,N_3898,N_3910);
nand U4183 (N_4183,N_3838,N_3795);
nor U4184 (N_4184,N_3794,N_3755);
or U4185 (N_4185,N_3889,N_3759);
nand U4186 (N_4186,N_3639,N_3719);
xnor U4187 (N_4187,N_3751,N_3858);
nor U4188 (N_4188,N_3512,N_3762);
nor U4189 (N_4189,N_3612,N_3781);
or U4190 (N_4190,N_3982,N_3628);
and U4191 (N_4191,N_3638,N_3673);
nand U4192 (N_4192,N_3534,N_3696);
and U4193 (N_4193,N_3920,N_3693);
nor U4194 (N_4194,N_3853,N_3597);
nand U4195 (N_4195,N_3938,N_3877);
and U4196 (N_4196,N_3934,N_3972);
or U4197 (N_4197,N_3903,N_3807);
nor U4198 (N_4198,N_3922,N_3557);
and U4199 (N_4199,N_3896,N_3729);
nand U4200 (N_4200,N_3874,N_3996);
or U4201 (N_4201,N_3611,N_3538);
or U4202 (N_4202,N_3994,N_3595);
nor U4203 (N_4203,N_3703,N_3624);
nor U4204 (N_4204,N_3653,N_3727);
nand U4205 (N_4205,N_3761,N_3547);
and U4206 (N_4206,N_3840,N_3763);
and U4207 (N_4207,N_3573,N_3820);
nand U4208 (N_4208,N_3937,N_3750);
or U4209 (N_4209,N_3605,N_3623);
nor U4210 (N_4210,N_3742,N_3503);
nor U4211 (N_4211,N_3797,N_3861);
nand U4212 (N_4212,N_3819,N_3667);
or U4213 (N_4213,N_3741,N_3670);
or U4214 (N_4214,N_3880,N_3648);
and U4215 (N_4215,N_3553,N_3683);
or U4216 (N_4216,N_3839,N_3842);
xor U4217 (N_4217,N_3654,N_3642);
and U4218 (N_4218,N_3652,N_3697);
and U4219 (N_4219,N_3662,N_3737);
or U4220 (N_4220,N_3981,N_3594);
or U4221 (N_4221,N_3968,N_3675);
and U4222 (N_4222,N_3834,N_3736);
or U4223 (N_4223,N_3940,N_3552);
nor U4224 (N_4224,N_3714,N_3546);
nor U4225 (N_4225,N_3772,N_3988);
xor U4226 (N_4226,N_3651,N_3911);
nor U4227 (N_4227,N_3985,N_3951);
and U4228 (N_4228,N_3817,N_3674);
nand U4229 (N_4229,N_3983,N_3916);
nor U4230 (N_4230,N_3564,N_3619);
nand U4231 (N_4231,N_3722,N_3851);
and U4232 (N_4232,N_3551,N_3833);
nor U4233 (N_4233,N_3743,N_3728);
nand U4234 (N_4234,N_3511,N_3908);
nand U4235 (N_4235,N_3805,N_3502);
nor U4236 (N_4236,N_3811,N_3579);
or U4237 (N_4237,N_3550,N_3521);
nor U4238 (N_4238,N_3804,N_3973);
and U4239 (N_4239,N_3532,N_3560);
xor U4240 (N_4240,N_3844,N_3986);
nand U4241 (N_4241,N_3501,N_3748);
and U4242 (N_4242,N_3608,N_3698);
or U4243 (N_4243,N_3873,N_3976);
and U4244 (N_4244,N_3902,N_3656);
nor U4245 (N_4245,N_3949,N_3876);
or U4246 (N_4246,N_3519,N_3660);
and U4247 (N_4247,N_3905,N_3677);
nor U4248 (N_4248,N_3704,N_3995);
nor U4249 (N_4249,N_3798,N_3964);
nand U4250 (N_4250,N_3509,N_3583);
and U4251 (N_4251,N_3974,N_3905);
nor U4252 (N_4252,N_3871,N_3667);
nor U4253 (N_4253,N_3741,N_3666);
and U4254 (N_4254,N_3902,N_3566);
and U4255 (N_4255,N_3778,N_3704);
or U4256 (N_4256,N_3921,N_3965);
and U4257 (N_4257,N_3815,N_3544);
and U4258 (N_4258,N_3592,N_3947);
or U4259 (N_4259,N_3774,N_3664);
and U4260 (N_4260,N_3677,N_3872);
xor U4261 (N_4261,N_3786,N_3565);
or U4262 (N_4262,N_3987,N_3984);
and U4263 (N_4263,N_3635,N_3944);
nand U4264 (N_4264,N_3875,N_3924);
or U4265 (N_4265,N_3504,N_3773);
and U4266 (N_4266,N_3946,N_3805);
or U4267 (N_4267,N_3840,N_3934);
xnor U4268 (N_4268,N_3956,N_3844);
nand U4269 (N_4269,N_3597,N_3634);
nand U4270 (N_4270,N_3617,N_3680);
nor U4271 (N_4271,N_3934,N_3529);
or U4272 (N_4272,N_3792,N_3961);
nor U4273 (N_4273,N_3597,N_3846);
nand U4274 (N_4274,N_3981,N_3774);
and U4275 (N_4275,N_3849,N_3730);
nand U4276 (N_4276,N_3737,N_3773);
nand U4277 (N_4277,N_3656,N_3881);
or U4278 (N_4278,N_3854,N_3674);
nand U4279 (N_4279,N_3806,N_3559);
nor U4280 (N_4280,N_3896,N_3509);
or U4281 (N_4281,N_3649,N_3668);
and U4282 (N_4282,N_3980,N_3598);
and U4283 (N_4283,N_3792,N_3925);
or U4284 (N_4284,N_3653,N_3919);
or U4285 (N_4285,N_3560,N_3503);
nand U4286 (N_4286,N_3601,N_3941);
or U4287 (N_4287,N_3569,N_3519);
nor U4288 (N_4288,N_3980,N_3523);
xor U4289 (N_4289,N_3773,N_3786);
nor U4290 (N_4290,N_3520,N_3933);
and U4291 (N_4291,N_3759,N_3907);
nor U4292 (N_4292,N_3942,N_3768);
nor U4293 (N_4293,N_3725,N_3752);
nand U4294 (N_4294,N_3518,N_3773);
nand U4295 (N_4295,N_3546,N_3756);
and U4296 (N_4296,N_3758,N_3985);
nor U4297 (N_4297,N_3921,N_3637);
and U4298 (N_4298,N_3964,N_3605);
and U4299 (N_4299,N_3808,N_3907);
nor U4300 (N_4300,N_3674,N_3571);
nand U4301 (N_4301,N_3564,N_3957);
and U4302 (N_4302,N_3852,N_3525);
nor U4303 (N_4303,N_3897,N_3969);
nand U4304 (N_4304,N_3606,N_3804);
or U4305 (N_4305,N_3805,N_3537);
or U4306 (N_4306,N_3541,N_3962);
nand U4307 (N_4307,N_3632,N_3532);
nor U4308 (N_4308,N_3652,N_3919);
nand U4309 (N_4309,N_3741,N_3838);
or U4310 (N_4310,N_3628,N_3821);
nand U4311 (N_4311,N_3789,N_3630);
nand U4312 (N_4312,N_3677,N_3867);
or U4313 (N_4313,N_3511,N_3504);
and U4314 (N_4314,N_3907,N_3795);
xor U4315 (N_4315,N_3545,N_3676);
and U4316 (N_4316,N_3758,N_3587);
or U4317 (N_4317,N_3745,N_3907);
nand U4318 (N_4318,N_3513,N_3904);
or U4319 (N_4319,N_3968,N_3534);
nand U4320 (N_4320,N_3715,N_3684);
nor U4321 (N_4321,N_3713,N_3586);
nor U4322 (N_4322,N_3554,N_3668);
or U4323 (N_4323,N_3970,N_3596);
and U4324 (N_4324,N_3905,N_3706);
nor U4325 (N_4325,N_3536,N_3572);
nand U4326 (N_4326,N_3993,N_3566);
or U4327 (N_4327,N_3946,N_3642);
and U4328 (N_4328,N_3519,N_3656);
nor U4329 (N_4329,N_3710,N_3555);
nor U4330 (N_4330,N_3624,N_3693);
and U4331 (N_4331,N_3705,N_3940);
nand U4332 (N_4332,N_3587,N_3763);
nor U4333 (N_4333,N_3577,N_3964);
nor U4334 (N_4334,N_3947,N_3662);
or U4335 (N_4335,N_3769,N_3513);
or U4336 (N_4336,N_3617,N_3917);
nand U4337 (N_4337,N_3963,N_3773);
nor U4338 (N_4338,N_3908,N_3860);
nor U4339 (N_4339,N_3536,N_3804);
nand U4340 (N_4340,N_3872,N_3632);
nand U4341 (N_4341,N_3528,N_3922);
nor U4342 (N_4342,N_3730,N_3959);
nand U4343 (N_4343,N_3846,N_3723);
nand U4344 (N_4344,N_3579,N_3525);
nand U4345 (N_4345,N_3545,N_3830);
nor U4346 (N_4346,N_3926,N_3616);
nand U4347 (N_4347,N_3896,N_3836);
and U4348 (N_4348,N_3886,N_3854);
and U4349 (N_4349,N_3589,N_3518);
and U4350 (N_4350,N_3763,N_3793);
or U4351 (N_4351,N_3937,N_3970);
nor U4352 (N_4352,N_3839,N_3702);
nor U4353 (N_4353,N_3533,N_3914);
and U4354 (N_4354,N_3767,N_3713);
nor U4355 (N_4355,N_3817,N_3597);
nand U4356 (N_4356,N_3975,N_3937);
nor U4357 (N_4357,N_3677,N_3574);
nor U4358 (N_4358,N_3526,N_3667);
or U4359 (N_4359,N_3552,N_3796);
and U4360 (N_4360,N_3973,N_3770);
nor U4361 (N_4361,N_3983,N_3617);
or U4362 (N_4362,N_3787,N_3805);
and U4363 (N_4363,N_3946,N_3814);
and U4364 (N_4364,N_3529,N_3776);
nand U4365 (N_4365,N_3836,N_3842);
nand U4366 (N_4366,N_3858,N_3551);
nor U4367 (N_4367,N_3947,N_3911);
nor U4368 (N_4368,N_3852,N_3676);
nor U4369 (N_4369,N_3670,N_3552);
and U4370 (N_4370,N_3561,N_3842);
nor U4371 (N_4371,N_3690,N_3939);
or U4372 (N_4372,N_3720,N_3558);
nor U4373 (N_4373,N_3878,N_3602);
and U4374 (N_4374,N_3735,N_3790);
nor U4375 (N_4375,N_3608,N_3553);
and U4376 (N_4376,N_3693,N_3761);
nor U4377 (N_4377,N_3682,N_3684);
or U4378 (N_4378,N_3534,N_3564);
and U4379 (N_4379,N_3781,N_3892);
or U4380 (N_4380,N_3697,N_3542);
nor U4381 (N_4381,N_3554,N_3909);
or U4382 (N_4382,N_3819,N_3563);
nor U4383 (N_4383,N_3869,N_3829);
nand U4384 (N_4384,N_3812,N_3774);
or U4385 (N_4385,N_3670,N_3526);
or U4386 (N_4386,N_3668,N_3841);
nand U4387 (N_4387,N_3547,N_3870);
nor U4388 (N_4388,N_3553,N_3769);
nand U4389 (N_4389,N_3741,N_3722);
or U4390 (N_4390,N_3752,N_3697);
and U4391 (N_4391,N_3607,N_3702);
nand U4392 (N_4392,N_3832,N_3834);
or U4393 (N_4393,N_3718,N_3682);
and U4394 (N_4394,N_3513,N_3859);
nand U4395 (N_4395,N_3838,N_3821);
and U4396 (N_4396,N_3773,N_3946);
or U4397 (N_4397,N_3983,N_3954);
nand U4398 (N_4398,N_3808,N_3858);
nor U4399 (N_4399,N_3651,N_3646);
nand U4400 (N_4400,N_3836,N_3957);
or U4401 (N_4401,N_3883,N_3506);
and U4402 (N_4402,N_3864,N_3784);
and U4403 (N_4403,N_3961,N_3981);
nor U4404 (N_4404,N_3553,N_3896);
nor U4405 (N_4405,N_3776,N_3937);
nor U4406 (N_4406,N_3517,N_3949);
nor U4407 (N_4407,N_3704,N_3963);
nor U4408 (N_4408,N_3863,N_3800);
nand U4409 (N_4409,N_3908,N_3628);
nor U4410 (N_4410,N_3580,N_3803);
nand U4411 (N_4411,N_3693,N_3989);
or U4412 (N_4412,N_3647,N_3947);
and U4413 (N_4413,N_3563,N_3933);
nand U4414 (N_4414,N_3578,N_3699);
xor U4415 (N_4415,N_3726,N_3766);
and U4416 (N_4416,N_3874,N_3998);
or U4417 (N_4417,N_3747,N_3931);
nor U4418 (N_4418,N_3521,N_3513);
and U4419 (N_4419,N_3966,N_3870);
nor U4420 (N_4420,N_3695,N_3975);
nor U4421 (N_4421,N_3775,N_3674);
or U4422 (N_4422,N_3756,N_3878);
or U4423 (N_4423,N_3507,N_3598);
nor U4424 (N_4424,N_3692,N_3999);
or U4425 (N_4425,N_3970,N_3756);
or U4426 (N_4426,N_3666,N_3503);
nand U4427 (N_4427,N_3696,N_3582);
and U4428 (N_4428,N_3546,N_3836);
nor U4429 (N_4429,N_3649,N_3756);
or U4430 (N_4430,N_3563,N_3923);
nand U4431 (N_4431,N_3663,N_3705);
and U4432 (N_4432,N_3557,N_3937);
or U4433 (N_4433,N_3767,N_3620);
and U4434 (N_4434,N_3510,N_3911);
xor U4435 (N_4435,N_3666,N_3711);
nand U4436 (N_4436,N_3507,N_3937);
and U4437 (N_4437,N_3552,N_3571);
and U4438 (N_4438,N_3680,N_3631);
nand U4439 (N_4439,N_3522,N_3611);
or U4440 (N_4440,N_3573,N_3824);
and U4441 (N_4441,N_3627,N_3505);
and U4442 (N_4442,N_3572,N_3587);
nor U4443 (N_4443,N_3574,N_3535);
or U4444 (N_4444,N_3597,N_3744);
or U4445 (N_4445,N_3884,N_3951);
nand U4446 (N_4446,N_3529,N_3741);
nand U4447 (N_4447,N_3505,N_3722);
or U4448 (N_4448,N_3738,N_3728);
or U4449 (N_4449,N_3732,N_3592);
nor U4450 (N_4450,N_3580,N_3847);
or U4451 (N_4451,N_3779,N_3589);
and U4452 (N_4452,N_3825,N_3954);
nand U4453 (N_4453,N_3856,N_3627);
xor U4454 (N_4454,N_3968,N_3773);
and U4455 (N_4455,N_3572,N_3686);
nor U4456 (N_4456,N_3517,N_3723);
nor U4457 (N_4457,N_3887,N_3744);
nor U4458 (N_4458,N_3592,N_3664);
xnor U4459 (N_4459,N_3798,N_3850);
and U4460 (N_4460,N_3501,N_3667);
or U4461 (N_4461,N_3971,N_3598);
nor U4462 (N_4462,N_3659,N_3505);
nand U4463 (N_4463,N_3794,N_3539);
or U4464 (N_4464,N_3780,N_3548);
nor U4465 (N_4465,N_3604,N_3593);
and U4466 (N_4466,N_3517,N_3615);
nor U4467 (N_4467,N_3801,N_3590);
and U4468 (N_4468,N_3721,N_3816);
or U4469 (N_4469,N_3863,N_3923);
and U4470 (N_4470,N_3587,N_3967);
nor U4471 (N_4471,N_3830,N_3989);
and U4472 (N_4472,N_3700,N_3738);
and U4473 (N_4473,N_3892,N_3739);
and U4474 (N_4474,N_3876,N_3737);
nand U4475 (N_4475,N_3997,N_3555);
nor U4476 (N_4476,N_3616,N_3916);
nor U4477 (N_4477,N_3512,N_3866);
and U4478 (N_4478,N_3567,N_3652);
and U4479 (N_4479,N_3931,N_3880);
nor U4480 (N_4480,N_3881,N_3864);
nor U4481 (N_4481,N_3875,N_3952);
and U4482 (N_4482,N_3994,N_3652);
or U4483 (N_4483,N_3713,N_3788);
nor U4484 (N_4484,N_3659,N_3653);
nor U4485 (N_4485,N_3676,N_3960);
nor U4486 (N_4486,N_3650,N_3915);
or U4487 (N_4487,N_3555,N_3587);
nand U4488 (N_4488,N_3596,N_3987);
or U4489 (N_4489,N_3945,N_3834);
or U4490 (N_4490,N_3809,N_3736);
nand U4491 (N_4491,N_3781,N_3716);
nand U4492 (N_4492,N_3629,N_3559);
nor U4493 (N_4493,N_3943,N_3604);
nor U4494 (N_4494,N_3748,N_3670);
or U4495 (N_4495,N_3930,N_3501);
nand U4496 (N_4496,N_3654,N_3774);
nand U4497 (N_4497,N_3612,N_3912);
and U4498 (N_4498,N_3864,N_3675);
nand U4499 (N_4499,N_3628,N_3696);
nand U4500 (N_4500,N_4325,N_4459);
or U4501 (N_4501,N_4029,N_4027);
nand U4502 (N_4502,N_4187,N_4490);
nor U4503 (N_4503,N_4494,N_4139);
nor U4504 (N_4504,N_4387,N_4236);
nand U4505 (N_4505,N_4167,N_4271);
nand U4506 (N_4506,N_4243,N_4478);
nand U4507 (N_4507,N_4200,N_4178);
and U4508 (N_4508,N_4204,N_4405);
nand U4509 (N_4509,N_4451,N_4359);
nand U4510 (N_4510,N_4026,N_4152);
nor U4511 (N_4511,N_4061,N_4153);
nor U4512 (N_4512,N_4313,N_4009);
nand U4513 (N_4513,N_4277,N_4496);
or U4514 (N_4514,N_4253,N_4293);
or U4515 (N_4515,N_4446,N_4372);
nor U4516 (N_4516,N_4196,N_4177);
nor U4517 (N_4517,N_4437,N_4242);
nor U4518 (N_4518,N_4415,N_4240);
and U4519 (N_4519,N_4488,N_4302);
nor U4520 (N_4520,N_4104,N_4191);
nand U4521 (N_4521,N_4054,N_4355);
nor U4522 (N_4522,N_4378,N_4186);
xor U4523 (N_4523,N_4474,N_4057);
and U4524 (N_4524,N_4477,N_4422);
or U4525 (N_4525,N_4332,N_4462);
and U4526 (N_4526,N_4099,N_4020);
nor U4527 (N_4527,N_4141,N_4450);
nand U4528 (N_4528,N_4369,N_4364);
and U4529 (N_4529,N_4129,N_4388);
xor U4530 (N_4530,N_4258,N_4376);
nand U4531 (N_4531,N_4118,N_4173);
xor U4532 (N_4532,N_4226,N_4321);
nand U4533 (N_4533,N_4328,N_4263);
nand U4534 (N_4534,N_4100,N_4439);
nor U4535 (N_4535,N_4008,N_4247);
or U4536 (N_4536,N_4434,N_4012);
xor U4537 (N_4537,N_4154,N_4259);
and U4538 (N_4538,N_4047,N_4498);
and U4539 (N_4539,N_4333,N_4163);
and U4540 (N_4540,N_4071,N_4194);
nand U4541 (N_4541,N_4175,N_4386);
nor U4542 (N_4542,N_4018,N_4048);
nor U4543 (N_4543,N_4400,N_4398);
or U4544 (N_4544,N_4032,N_4377);
or U4545 (N_4545,N_4119,N_4114);
and U4546 (N_4546,N_4475,N_4250);
nor U4547 (N_4547,N_4438,N_4116);
and U4548 (N_4548,N_4463,N_4429);
and U4549 (N_4549,N_4076,N_4025);
nor U4550 (N_4550,N_4455,N_4158);
and U4551 (N_4551,N_4288,N_4481);
nand U4552 (N_4552,N_4416,N_4456);
and U4553 (N_4553,N_4228,N_4397);
and U4554 (N_4554,N_4296,N_4207);
or U4555 (N_4555,N_4329,N_4334);
nand U4556 (N_4556,N_4130,N_4350);
nor U4557 (N_4557,N_4442,N_4410);
nor U4558 (N_4558,N_4469,N_4436);
or U4559 (N_4559,N_4335,N_4148);
nor U4560 (N_4560,N_4093,N_4495);
nand U4561 (N_4561,N_4004,N_4034);
or U4562 (N_4562,N_4491,N_4384);
nand U4563 (N_4563,N_4183,N_4294);
or U4564 (N_4564,N_4246,N_4021);
nor U4565 (N_4565,N_4430,N_4274);
nand U4566 (N_4566,N_4460,N_4322);
nand U4567 (N_4567,N_4337,N_4185);
nand U4568 (N_4568,N_4443,N_4316);
and U4569 (N_4569,N_4353,N_4087);
or U4570 (N_4570,N_4064,N_4107);
or U4571 (N_4571,N_4180,N_4171);
nand U4572 (N_4572,N_4361,N_4188);
nand U4573 (N_4573,N_4075,N_4233);
and U4574 (N_4574,N_4159,N_4134);
or U4575 (N_4575,N_4345,N_4254);
nor U4576 (N_4576,N_4380,N_4111);
nor U4577 (N_4577,N_4275,N_4371);
nor U4578 (N_4578,N_4120,N_4062);
and U4579 (N_4579,N_4352,N_4417);
and U4580 (N_4580,N_4035,N_4287);
and U4581 (N_4581,N_4065,N_4454);
or U4582 (N_4582,N_4298,N_4000);
and U4583 (N_4583,N_4007,N_4015);
nor U4584 (N_4584,N_4037,N_4382);
nor U4585 (N_4585,N_4425,N_4343);
and U4586 (N_4586,N_4472,N_4217);
and U4587 (N_4587,N_4470,N_4391);
nand U4588 (N_4588,N_4096,N_4081);
or U4589 (N_4589,N_4110,N_4338);
nor U4590 (N_4590,N_4305,N_4255);
and U4591 (N_4591,N_4390,N_4401);
and U4592 (N_4592,N_4273,N_4205);
nor U4593 (N_4593,N_4402,N_4306);
and U4594 (N_4594,N_4272,N_4069);
and U4595 (N_4595,N_4349,N_4143);
or U4596 (N_4596,N_4435,N_4010);
nor U4597 (N_4597,N_4101,N_4304);
and U4598 (N_4598,N_4458,N_4105);
or U4599 (N_4599,N_4484,N_4112);
and U4600 (N_4600,N_4059,N_4176);
nor U4601 (N_4601,N_4285,N_4145);
xor U4602 (N_4602,N_4042,N_4465);
and U4603 (N_4603,N_4385,N_4219);
and U4604 (N_4604,N_4136,N_4082);
nand U4605 (N_4605,N_4419,N_4327);
and U4606 (N_4606,N_4016,N_4482);
nand U4607 (N_4607,N_4256,N_4072);
and U4608 (N_4608,N_4138,N_4168);
or U4609 (N_4609,N_4408,N_4150);
or U4610 (N_4610,N_4108,N_4146);
and U4611 (N_4611,N_4166,N_4039);
nand U4612 (N_4612,N_4080,N_4097);
and U4613 (N_4613,N_4070,N_4311);
or U4614 (N_4614,N_4467,N_4210);
or U4615 (N_4615,N_4428,N_4133);
or U4616 (N_4616,N_4006,N_4374);
nor U4617 (N_4617,N_4055,N_4307);
and U4618 (N_4618,N_4461,N_4457);
nand U4619 (N_4619,N_4289,N_4440);
and U4620 (N_4620,N_4238,N_4297);
and U4621 (N_4621,N_4487,N_4199);
nor U4622 (N_4622,N_4208,N_4041);
nor U4623 (N_4623,N_4278,N_4261);
nor U4624 (N_4624,N_4124,N_4348);
or U4625 (N_4625,N_4181,N_4286);
nor U4626 (N_4626,N_4389,N_4373);
nand U4627 (N_4627,N_4149,N_4002);
and U4628 (N_4628,N_4418,N_4339);
or U4629 (N_4629,N_4170,N_4357);
or U4630 (N_4630,N_4427,N_4431);
and U4631 (N_4631,N_4028,N_4203);
or U4632 (N_4632,N_4342,N_4227);
nor U4633 (N_4633,N_4392,N_4091);
nand U4634 (N_4634,N_4038,N_4403);
or U4635 (N_4635,N_4314,N_4040);
nand U4636 (N_4636,N_4106,N_4090);
nor U4637 (N_4637,N_4235,N_4368);
xnor U4638 (N_4638,N_4165,N_4320);
or U4639 (N_4639,N_4365,N_4407);
nand U4640 (N_4640,N_4102,N_4162);
or U4641 (N_4641,N_4326,N_4137);
nand U4642 (N_4642,N_4354,N_4395);
or U4643 (N_4643,N_4471,N_4366);
or U4644 (N_4644,N_4157,N_4115);
nor U4645 (N_4645,N_4346,N_4221);
and U4646 (N_4646,N_4237,N_4156);
or U4647 (N_4647,N_4098,N_4411);
nand U4648 (N_4648,N_4375,N_4014);
nand U4649 (N_4649,N_4089,N_4497);
and U4650 (N_4650,N_4270,N_4249);
and U4651 (N_4651,N_4290,N_4225);
nand U4652 (N_4652,N_4161,N_4300);
nor U4653 (N_4653,N_4051,N_4449);
or U4654 (N_4654,N_4215,N_4022);
or U4655 (N_4655,N_4444,N_4312);
or U4656 (N_4656,N_4267,N_4045);
xor U4657 (N_4657,N_4229,N_4309);
and U4658 (N_4658,N_4182,N_4257);
nor U4659 (N_4659,N_4117,N_4193);
nor U4660 (N_4660,N_4414,N_4299);
nor U4661 (N_4661,N_4142,N_4190);
nand U4662 (N_4662,N_4383,N_4426);
nor U4663 (N_4663,N_4283,N_4077);
and U4664 (N_4664,N_4030,N_4031);
nand U4665 (N_4665,N_4011,N_4239);
or U4666 (N_4666,N_4245,N_4362);
or U4667 (N_4667,N_4052,N_4131);
nand U4668 (N_4668,N_4127,N_4195);
nor U4669 (N_4669,N_4284,N_4485);
xor U4670 (N_4670,N_4399,N_4085);
and U4671 (N_4671,N_4269,N_4220);
nand U4672 (N_4672,N_4432,N_4151);
or U4673 (N_4673,N_4086,N_4232);
or U4674 (N_4674,N_4192,N_4358);
or U4675 (N_4675,N_4295,N_4292);
nor U4676 (N_4676,N_4073,N_4447);
nand U4677 (N_4677,N_4356,N_4466);
nor U4678 (N_4678,N_4340,N_4452);
nand U4679 (N_4679,N_4056,N_4172);
nor U4680 (N_4680,N_4063,N_4140);
and U4681 (N_4681,N_4291,N_4370);
nand U4682 (N_4682,N_4214,N_4360);
and U4683 (N_4683,N_4406,N_4480);
and U4684 (N_4684,N_4084,N_4351);
nor U4685 (N_4685,N_4019,N_4202);
or U4686 (N_4686,N_4336,N_4103);
nor U4687 (N_4687,N_4174,N_4024);
nand U4688 (N_4688,N_4394,N_4265);
or U4689 (N_4689,N_4079,N_4260);
nand U4690 (N_4690,N_4088,N_4067);
nor U4691 (N_4691,N_4135,N_4033);
or U4692 (N_4692,N_4218,N_4280);
nor U4693 (N_4693,N_4412,N_4264);
and U4694 (N_4694,N_4147,N_4424);
nor U4695 (N_4695,N_4363,N_4367);
nor U4696 (N_4696,N_4169,N_4144);
nand U4697 (N_4697,N_4441,N_4486);
and U4698 (N_4698,N_4068,N_4310);
and U4699 (N_4699,N_4160,N_4303);
or U4700 (N_4700,N_4381,N_4060);
xnor U4701 (N_4701,N_4268,N_4379);
or U4702 (N_4702,N_4341,N_4074);
and U4703 (N_4703,N_4433,N_4128);
or U4704 (N_4704,N_4483,N_4109);
or U4705 (N_4705,N_4420,N_4211);
nor U4706 (N_4706,N_4083,N_4184);
nor U4707 (N_4707,N_4492,N_4445);
nand U4708 (N_4708,N_4213,N_4094);
nand U4709 (N_4709,N_4262,N_4164);
xor U4710 (N_4710,N_4315,N_4050);
nand U4711 (N_4711,N_4058,N_4234);
nand U4712 (N_4712,N_4036,N_4252);
and U4713 (N_4713,N_4248,N_4005);
nor U4714 (N_4714,N_4493,N_4013);
and U4715 (N_4715,N_4003,N_4223);
and U4716 (N_4716,N_4319,N_4421);
nand U4717 (N_4717,N_4023,N_4053);
xnor U4718 (N_4718,N_4476,N_4231);
nor U4719 (N_4719,N_4046,N_4241);
or U4720 (N_4720,N_4281,N_4330);
and U4721 (N_4721,N_4279,N_4409);
nor U4722 (N_4722,N_4201,N_4230);
nand U4723 (N_4723,N_4301,N_4122);
and U4724 (N_4724,N_4323,N_4423);
nor U4725 (N_4725,N_4224,N_4282);
nor U4726 (N_4726,N_4043,N_4078);
nand U4727 (N_4727,N_4212,N_4113);
or U4728 (N_4728,N_4198,N_4473);
and U4729 (N_4729,N_4197,N_4448);
xnor U4730 (N_4730,N_4206,N_4393);
and U4731 (N_4731,N_4266,N_4404);
nor U4732 (N_4732,N_4464,N_4479);
or U4733 (N_4733,N_4044,N_4347);
and U4734 (N_4734,N_4155,N_4189);
nand U4735 (N_4735,N_4017,N_4413);
nand U4736 (N_4736,N_4216,N_4179);
nor U4737 (N_4737,N_4396,N_4251);
and U4738 (N_4738,N_4276,N_4317);
nand U4739 (N_4739,N_4132,N_4344);
or U4740 (N_4740,N_4121,N_4244);
nand U4741 (N_4741,N_4489,N_4066);
nor U4742 (N_4742,N_4125,N_4092);
and U4743 (N_4743,N_4324,N_4308);
xor U4744 (N_4744,N_4499,N_4095);
or U4745 (N_4745,N_4209,N_4468);
and U4746 (N_4746,N_4222,N_4049);
nor U4747 (N_4747,N_4453,N_4123);
nand U4748 (N_4748,N_4126,N_4001);
xor U4749 (N_4749,N_4318,N_4331);
or U4750 (N_4750,N_4475,N_4213);
or U4751 (N_4751,N_4202,N_4407);
nand U4752 (N_4752,N_4453,N_4243);
nor U4753 (N_4753,N_4321,N_4083);
or U4754 (N_4754,N_4242,N_4303);
nand U4755 (N_4755,N_4437,N_4036);
or U4756 (N_4756,N_4439,N_4466);
or U4757 (N_4757,N_4044,N_4394);
or U4758 (N_4758,N_4208,N_4122);
and U4759 (N_4759,N_4022,N_4331);
or U4760 (N_4760,N_4186,N_4361);
and U4761 (N_4761,N_4444,N_4417);
and U4762 (N_4762,N_4032,N_4394);
nor U4763 (N_4763,N_4192,N_4114);
and U4764 (N_4764,N_4234,N_4424);
nand U4765 (N_4765,N_4181,N_4028);
and U4766 (N_4766,N_4394,N_4136);
or U4767 (N_4767,N_4045,N_4110);
nor U4768 (N_4768,N_4179,N_4088);
nor U4769 (N_4769,N_4106,N_4000);
nand U4770 (N_4770,N_4138,N_4430);
and U4771 (N_4771,N_4240,N_4436);
and U4772 (N_4772,N_4294,N_4264);
nor U4773 (N_4773,N_4040,N_4247);
nor U4774 (N_4774,N_4218,N_4363);
nor U4775 (N_4775,N_4067,N_4335);
nor U4776 (N_4776,N_4458,N_4251);
nand U4777 (N_4777,N_4121,N_4374);
or U4778 (N_4778,N_4242,N_4461);
nand U4779 (N_4779,N_4439,N_4163);
xor U4780 (N_4780,N_4278,N_4262);
and U4781 (N_4781,N_4234,N_4343);
or U4782 (N_4782,N_4117,N_4433);
nand U4783 (N_4783,N_4069,N_4395);
nand U4784 (N_4784,N_4373,N_4105);
nor U4785 (N_4785,N_4010,N_4407);
nor U4786 (N_4786,N_4117,N_4327);
and U4787 (N_4787,N_4454,N_4278);
or U4788 (N_4788,N_4063,N_4294);
nand U4789 (N_4789,N_4407,N_4275);
nand U4790 (N_4790,N_4396,N_4350);
or U4791 (N_4791,N_4367,N_4078);
nand U4792 (N_4792,N_4187,N_4076);
nor U4793 (N_4793,N_4484,N_4122);
or U4794 (N_4794,N_4108,N_4480);
and U4795 (N_4795,N_4308,N_4191);
or U4796 (N_4796,N_4263,N_4427);
and U4797 (N_4797,N_4152,N_4122);
or U4798 (N_4798,N_4410,N_4068);
nor U4799 (N_4799,N_4233,N_4498);
and U4800 (N_4800,N_4428,N_4282);
and U4801 (N_4801,N_4203,N_4363);
or U4802 (N_4802,N_4175,N_4370);
xnor U4803 (N_4803,N_4456,N_4423);
nor U4804 (N_4804,N_4020,N_4492);
nand U4805 (N_4805,N_4203,N_4191);
nand U4806 (N_4806,N_4248,N_4193);
or U4807 (N_4807,N_4351,N_4142);
nand U4808 (N_4808,N_4096,N_4263);
nand U4809 (N_4809,N_4102,N_4237);
nor U4810 (N_4810,N_4478,N_4102);
nor U4811 (N_4811,N_4297,N_4149);
nand U4812 (N_4812,N_4012,N_4317);
nand U4813 (N_4813,N_4230,N_4113);
or U4814 (N_4814,N_4112,N_4103);
and U4815 (N_4815,N_4374,N_4158);
and U4816 (N_4816,N_4032,N_4096);
nand U4817 (N_4817,N_4327,N_4136);
and U4818 (N_4818,N_4317,N_4100);
nor U4819 (N_4819,N_4401,N_4385);
nand U4820 (N_4820,N_4410,N_4076);
and U4821 (N_4821,N_4176,N_4251);
nor U4822 (N_4822,N_4118,N_4094);
and U4823 (N_4823,N_4326,N_4108);
nand U4824 (N_4824,N_4175,N_4372);
and U4825 (N_4825,N_4156,N_4307);
and U4826 (N_4826,N_4101,N_4452);
or U4827 (N_4827,N_4495,N_4019);
nor U4828 (N_4828,N_4188,N_4337);
or U4829 (N_4829,N_4238,N_4423);
nor U4830 (N_4830,N_4398,N_4177);
or U4831 (N_4831,N_4492,N_4402);
and U4832 (N_4832,N_4442,N_4269);
and U4833 (N_4833,N_4238,N_4270);
and U4834 (N_4834,N_4214,N_4053);
and U4835 (N_4835,N_4174,N_4148);
nand U4836 (N_4836,N_4181,N_4144);
xor U4837 (N_4837,N_4269,N_4257);
nand U4838 (N_4838,N_4059,N_4038);
nor U4839 (N_4839,N_4087,N_4336);
and U4840 (N_4840,N_4065,N_4422);
nor U4841 (N_4841,N_4013,N_4416);
and U4842 (N_4842,N_4413,N_4483);
nand U4843 (N_4843,N_4377,N_4224);
nor U4844 (N_4844,N_4224,N_4136);
or U4845 (N_4845,N_4180,N_4291);
nor U4846 (N_4846,N_4047,N_4049);
and U4847 (N_4847,N_4097,N_4104);
or U4848 (N_4848,N_4311,N_4379);
and U4849 (N_4849,N_4483,N_4419);
or U4850 (N_4850,N_4157,N_4444);
nor U4851 (N_4851,N_4295,N_4037);
nor U4852 (N_4852,N_4116,N_4257);
nand U4853 (N_4853,N_4263,N_4327);
and U4854 (N_4854,N_4005,N_4488);
nor U4855 (N_4855,N_4276,N_4026);
and U4856 (N_4856,N_4204,N_4075);
nand U4857 (N_4857,N_4397,N_4402);
or U4858 (N_4858,N_4385,N_4382);
nand U4859 (N_4859,N_4160,N_4496);
nand U4860 (N_4860,N_4237,N_4338);
nand U4861 (N_4861,N_4069,N_4485);
xnor U4862 (N_4862,N_4190,N_4030);
nor U4863 (N_4863,N_4278,N_4225);
nor U4864 (N_4864,N_4218,N_4084);
nor U4865 (N_4865,N_4211,N_4421);
nor U4866 (N_4866,N_4326,N_4343);
nand U4867 (N_4867,N_4180,N_4218);
nor U4868 (N_4868,N_4140,N_4217);
nand U4869 (N_4869,N_4393,N_4051);
or U4870 (N_4870,N_4359,N_4395);
and U4871 (N_4871,N_4013,N_4232);
and U4872 (N_4872,N_4154,N_4416);
nand U4873 (N_4873,N_4470,N_4025);
or U4874 (N_4874,N_4041,N_4414);
nor U4875 (N_4875,N_4201,N_4287);
nand U4876 (N_4876,N_4132,N_4011);
or U4877 (N_4877,N_4420,N_4062);
or U4878 (N_4878,N_4016,N_4423);
nand U4879 (N_4879,N_4229,N_4362);
and U4880 (N_4880,N_4462,N_4221);
nor U4881 (N_4881,N_4381,N_4469);
or U4882 (N_4882,N_4251,N_4410);
and U4883 (N_4883,N_4169,N_4365);
nand U4884 (N_4884,N_4063,N_4251);
nor U4885 (N_4885,N_4463,N_4498);
xnor U4886 (N_4886,N_4186,N_4483);
and U4887 (N_4887,N_4152,N_4282);
and U4888 (N_4888,N_4372,N_4399);
xor U4889 (N_4889,N_4228,N_4026);
and U4890 (N_4890,N_4485,N_4271);
nor U4891 (N_4891,N_4205,N_4191);
and U4892 (N_4892,N_4308,N_4340);
nand U4893 (N_4893,N_4312,N_4136);
nor U4894 (N_4894,N_4478,N_4281);
or U4895 (N_4895,N_4413,N_4251);
and U4896 (N_4896,N_4428,N_4279);
and U4897 (N_4897,N_4113,N_4438);
and U4898 (N_4898,N_4158,N_4160);
nor U4899 (N_4899,N_4283,N_4009);
nor U4900 (N_4900,N_4098,N_4437);
or U4901 (N_4901,N_4227,N_4311);
nor U4902 (N_4902,N_4248,N_4273);
nor U4903 (N_4903,N_4463,N_4237);
nor U4904 (N_4904,N_4259,N_4162);
and U4905 (N_4905,N_4036,N_4418);
or U4906 (N_4906,N_4418,N_4153);
nand U4907 (N_4907,N_4482,N_4437);
and U4908 (N_4908,N_4448,N_4081);
nor U4909 (N_4909,N_4155,N_4049);
nand U4910 (N_4910,N_4038,N_4367);
or U4911 (N_4911,N_4396,N_4153);
nand U4912 (N_4912,N_4038,N_4127);
or U4913 (N_4913,N_4142,N_4171);
and U4914 (N_4914,N_4128,N_4167);
nor U4915 (N_4915,N_4047,N_4309);
nand U4916 (N_4916,N_4367,N_4343);
or U4917 (N_4917,N_4419,N_4016);
nor U4918 (N_4918,N_4081,N_4134);
or U4919 (N_4919,N_4113,N_4117);
and U4920 (N_4920,N_4268,N_4114);
or U4921 (N_4921,N_4493,N_4329);
nor U4922 (N_4922,N_4061,N_4299);
nor U4923 (N_4923,N_4495,N_4127);
nor U4924 (N_4924,N_4187,N_4142);
nand U4925 (N_4925,N_4300,N_4359);
and U4926 (N_4926,N_4369,N_4217);
or U4927 (N_4927,N_4250,N_4451);
nand U4928 (N_4928,N_4071,N_4374);
and U4929 (N_4929,N_4448,N_4470);
nor U4930 (N_4930,N_4040,N_4412);
and U4931 (N_4931,N_4160,N_4401);
nor U4932 (N_4932,N_4438,N_4008);
and U4933 (N_4933,N_4101,N_4124);
nand U4934 (N_4934,N_4126,N_4178);
or U4935 (N_4935,N_4465,N_4298);
and U4936 (N_4936,N_4442,N_4002);
or U4937 (N_4937,N_4183,N_4105);
or U4938 (N_4938,N_4477,N_4175);
nor U4939 (N_4939,N_4096,N_4476);
nand U4940 (N_4940,N_4209,N_4293);
or U4941 (N_4941,N_4057,N_4293);
nand U4942 (N_4942,N_4047,N_4396);
nor U4943 (N_4943,N_4259,N_4257);
nand U4944 (N_4944,N_4306,N_4006);
nand U4945 (N_4945,N_4168,N_4072);
and U4946 (N_4946,N_4152,N_4079);
or U4947 (N_4947,N_4314,N_4193);
and U4948 (N_4948,N_4023,N_4436);
nor U4949 (N_4949,N_4197,N_4393);
nand U4950 (N_4950,N_4246,N_4301);
and U4951 (N_4951,N_4242,N_4314);
nand U4952 (N_4952,N_4132,N_4039);
nor U4953 (N_4953,N_4347,N_4489);
and U4954 (N_4954,N_4463,N_4297);
or U4955 (N_4955,N_4009,N_4134);
nand U4956 (N_4956,N_4327,N_4166);
nand U4957 (N_4957,N_4282,N_4160);
nor U4958 (N_4958,N_4357,N_4030);
nor U4959 (N_4959,N_4390,N_4468);
or U4960 (N_4960,N_4173,N_4087);
and U4961 (N_4961,N_4409,N_4244);
nor U4962 (N_4962,N_4063,N_4249);
and U4963 (N_4963,N_4009,N_4462);
nand U4964 (N_4964,N_4249,N_4314);
nand U4965 (N_4965,N_4457,N_4008);
nand U4966 (N_4966,N_4066,N_4223);
nand U4967 (N_4967,N_4374,N_4425);
or U4968 (N_4968,N_4385,N_4201);
and U4969 (N_4969,N_4226,N_4056);
nand U4970 (N_4970,N_4156,N_4242);
nor U4971 (N_4971,N_4287,N_4215);
and U4972 (N_4972,N_4130,N_4462);
or U4973 (N_4973,N_4074,N_4089);
or U4974 (N_4974,N_4087,N_4102);
nand U4975 (N_4975,N_4290,N_4413);
or U4976 (N_4976,N_4035,N_4332);
nand U4977 (N_4977,N_4058,N_4169);
or U4978 (N_4978,N_4360,N_4305);
nor U4979 (N_4979,N_4319,N_4000);
nor U4980 (N_4980,N_4229,N_4121);
nor U4981 (N_4981,N_4348,N_4419);
or U4982 (N_4982,N_4152,N_4112);
or U4983 (N_4983,N_4248,N_4132);
or U4984 (N_4984,N_4167,N_4402);
or U4985 (N_4985,N_4212,N_4384);
or U4986 (N_4986,N_4070,N_4095);
nor U4987 (N_4987,N_4087,N_4023);
or U4988 (N_4988,N_4346,N_4152);
nor U4989 (N_4989,N_4039,N_4113);
nand U4990 (N_4990,N_4016,N_4153);
and U4991 (N_4991,N_4438,N_4149);
nand U4992 (N_4992,N_4493,N_4148);
nand U4993 (N_4993,N_4251,N_4435);
or U4994 (N_4994,N_4451,N_4407);
nand U4995 (N_4995,N_4052,N_4214);
and U4996 (N_4996,N_4093,N_4385);
or U4997 (N_4997,N_4270,N_4005);
and U4998 (N_4998,N_4057,N_4312);
or U4999 (N_4999,N_4413,N_4382);
and UO_0 (O_0,N_4967,N_4599);
xnor UO_1 (O_1,N_4532,N_4804);
and UO_2 (O_2,N_4616,N_4627);
nor UO_3 (O_3,N_4564,N_4988);
nor UO_4 (O_4,N_4632,N_4869);
or UO_5 (O_5,N_4536,N_4764);
nor UO_6 (O_6,N_4876,N_4574);
nand UO_7 (O_7,N_4663,N_4946);
or UO_8 (O_8,N_4662,N_4711);
or UO_9 (O_9,N_4707,N_4612);
and UO_10 (O_10,N_4505,N_4693);
nor UO_11 (O_11,N_4813,N_4636);
nand UO_12 (O_12,N_4940,N_4509);
xor UO_13 (O_13,N_4676,N_4561);
nor UO_14 (O_14,N_4805,N_4782);
nand UO_15 (O_15,N_4892,N_4987);
nand UO_16 (O_16,N_4559,N_4969);
and UO_17 (O_17,N_4793,N_4728);
or UO_18 (O_18,N_4611,N_4710);
and UO_19 (O_19,N_4571,N_4588);
nand UO_20 (O_20,N_4580,N_4642);
and UO_21 (O_21,N_4698,N_4515);
or UO_22 (O_22,N_4885,N_4689);
or UO_23 (O_23,N_4590,N_4744);
nand UO_24 (O_24,N_4553,N_4774);
nor UO_25 (O_25,N_4942,N_4667);
nor UO_26 (O_26,N_4949,N_4752);
and UO_27 (O_27,N_4842,N_4549);
nor UO_28 (O_28,N_4816,N_4558);
or UO_29 (O_29,N_4657,N_4702);
nor UO_30 (O_30,N_4933,N_4716);
nor UO_31 (O_31,N_4851,N_4589);
nor UO_32 (O_32,N_4618,N_4672);
nand UO_33 (O_33,N_4637,N_4759);
nand UO_34 (O_34,N_4850,N_4978);
or UO_35 (O_35,N_4706,N_4932);
or UO_36 (O_36,N_4777,N_4890);
or UO_37 (O_37,N_4545,N_4837);
and UO_38 (O_38,N_4897,N_4770);
nand UO_39 (O_39,N_4838,N_4535);
or UO_40 (O_40,N_4790,N_4779);
and UO_41 (O_41,N_4605,N_4660);
and UO_42 (O_42,N_4846,N_4715);
nand UO_43 (O_43,N_4854,N_4938);
and UO_44 (O_44,N_4852,N_4824);
and UO_45 (O_45,N_4704,N_4740);
nand UO_46 (O_46,N_4576,N_4925);
or UO_47 (O_47,N_4802,N_4986);
or UO_48 (O_48,N_4705,N_4750);
nor UO_49 (O_49,N_4908,N_4621);
and UO_50 (O_50,N_4921,N_4628);
nor UO_51 (O_51,N_4748,N_4501);
nor UO_52 (O_52,N_4718,N_4794);
nor UO_53 (O_53,N_4993,N_4861);
or UO_54 (O_54,N_4935,N_4954);
or UO_55 (O_55,N_4769,N_4555);
and UO_56 (O_56,N_4845,N_4812);
or UO_57 (O_57,N_4626,N_4709);
nand UO_58 (O_58,N_4739,N_4664);
nand UO_59 (O_59,N_4904,N_4862);
nor UO_60 (O_60,N_4955,N_4582);
or UO_61 (O_61,N_4650,N_4806);
nor UO_62 (O_62,N_4609,N_4974);
and UO_63 (O_63,N_4570,N_4738);
nor UO_64 (O_64,N_4755,N_4581);
nor UO_65 (O_65,N_4893,N_4595);
and UO_66 (O_66,N_4931,N_4714);
and UO_67 (O_67,N_4525,N_4602);
and UO_68 (O_68,N_4977,N_4508);
nor UO_69 (O_69,N_4849,N_4763);
xor UO_70 (O_70,N_4873,N_4953);
or UO_71 (O_71,N_4780,N_4810);
nand UO_72 (O_72,N_4903,N_4701);
and UO_73 (O_73,N_4533,N_4573);
and UO_74 (O_74,N_4947,N_4819);
or UO_75 (O_75,N_4775,N_4733);
xnor UO_76 (O_76,N_4756,N_4964);
or UO_77 (O_77,N_4762,N_4922);
nor UO_78 (O_78,N_4907,N_4784);
and UO_79 (O_79,N_4649,N_4853);
nand UO_80 (O_80,N_4587,N_4843);
or UO_81 (O_81,N_4923,N_4644);
xnor UO_82 (O_82,N_4634,N_4631);
or UO_83 (O_83,N_4550,N_4537);
nand UO_84 (O_84,N_4567,N_4717);
or UO_85 (O_85,N_4735,N_4982);
nor UO_86 (O_86,N_4924,N_4792);
nor UO_87 (O_87,N_4523,N_4615);
xnor UO_88 (O_88,N_4963,N_4504);
and UO_89 (O_89,N_4512,N_4554);
and UO_90 (O_90,N_4655,N_4510);
nand UO_91 (O_91,N_4699,N_4857);
nor UO_92 (O_92,N_4965,N_4884);
nand UO_93 (O_93,N_4678,N_4679);
nor UO_94 (O_94,N_4668,N_4630);
or UO_95 (O_95,N_4591,N_4917);
and UO_96 (O_96,N_4848,N_4839);
nor UO_97 (O_97,N_4785,N_4973);
or UO_98 (O_98,N_4633,N_4765);
nor UO_99 (O_99,N_4592,N_4860);
or UO_100 (O_100,N_4522,N_4865);
nor UO_101 (O_101,N_4970,N_4541);
or UO_102 (O_102,N_4640,N_4795);
xor UO_103 (O_103,N_4999,N_4788);
nor UO_104 (O_104,N_4868,N_4825);
nor UO_105 (O_105,N_4513,N_4514);
nand UO_106 (O_106,N_4786,N_4635);
or UO_107 (O_107,N_4856,N_4529);
or UO_108 (O_108,N_4871,N_4641);
nor UO_109 (O_109,N_4872,N_4734);
nor UO_110 (O_110,N_4929,N_4697);
nor UO_111 (O_111,N_4844,N_4817);
or UO_112 (O_112,N_4915,N_4959);
nor UO_113 (O_113,N_4858,N_4766);
or UO_114 (O_114,N_4749,N_4874);
nor UO_115 (O_115,N_4530,N_4606);
nand UO_116 (O_116,N_4593,N_4563);
nor UO_117 (O_117,N_4654,N_4565);
nand UO_118 (O_118,N_4518,N_4724);
and UO_119 (O_119,N_4544,N_4562);
nand UO_120 (O_120,N_4551,N_4556);
or UO_121 (O_121,N_4507,N_4761);
nor UO_122 (O_122,N_4661,N_4961);
or UO_123 (O_123,N_4934,N_4998);
nand UO_124 (O_124,N_4913,N_4952);
and UO_125 (O_125,N_4771,N_4539);
or UO_126 (O_126,N_4997,N_4741);
nor UO_127 (O_127,N_4936,N_4624);
nand UO_128 (O_128,N_4737,N_4579);
nand UO_129 (O_129,N_4877,N_4975);
or UO_130 (O_130,N_4822,N_4976);
nand UO_131 (O_131,N_4727,N_4866);
nand UO_132 (O_132,N_4500,N_4673);
nor UO_133 (O_133,N_4909,N_4905);
or UO_134 (O_134,N_4878,N_4894);
nand UO_135 (O_135,N_4680,N_4972);
and UO_136 (O_136,N_4674,N_4677);
or UO_137 (O_137,N_4503,N_4538);
and UO_138 (O_138,N_4597,N_4653);
nand UO_139 (O_139,N_4826,N_4557);
nor UO_140 (O_140,N_4891,N_4989);
xor UO_141 (O_141,N_4623,N_4746);
nand UO_142 (O_142,N_4617,N_4614);
or UO_143 (O_143,N_4902,N_4984);
or UO_144 (O_144,N_4966,N_4683);
and UO_145 (O_145,N_4800,N_4596);
xnor UO_146 (O_146,N_4773,N_4552);
or UO_147 (O_147,N_4656,N_4991);
nand UO_148 (O_148,N_4979,N_4586);
and UO_149 (O_149,N_4747,N_4910);
nor UO_150 (O_150,N_4753,N_4781);
or UO_151 (O_151,N_4524,N_4815);
nand UO_152 (O_152,N_4543,N_4708);
nor UO_153 (O_153,N_4814,N_4540);
or UO_154 (O_154,N_4758,N_4566);
nand UO_155 (O_155,N_4939,N_4951);
nand UO_156 (O_156,N_4686,N_4888);
and UO_157 (O_157,N_4918,N_4990);
nand UO_158 (O_158,N_4883,N_4681);
or UO_159 (O_159,N_4807,N_4569);
or UO_160 (O_160,N_4945,N_4783);
nor UO_161 (O_161,N_4911,N_4767);
or UO_162 (O_162,N_4721,N_4809);
nand UO_163 (O_163,N_4604,N_4643);
nand UO_164 (O_164,N_4958,N_4742);
and UO_165 (O_165,N_4687,N_4896);
or UO_166 (O_166,N_4542,N_4887);
and UO_167 (O_167,N_4517,N_4534);
nor UO_168 (O_168,N_4886,N_4808);
and UO_169 (O_169,N_4731,N_4516);
nor UO_170 (O_170,N_4692,N_4801);
xnor UO_171 (O_171,N_4684,N_4906);
or UO_172 (O_172,N_4700,N_4743);
or UO_173 (O_173,N_4578,N_4688);
nor UO_174 (O_174,N_4960,N_4528);
and UO_175 (O_175,N_4875,N_4797);
nor UO_176 (O_176,N_4919,N_4996);
nand UO_177 (O_177,N_4796,N_4620);
nor UO_178 (O_178,N_4899,N_4726);
nor UO_179 (O_179,N_4927,N_4703);
or UO_180 (O_180,N_4778,N_4527);
nor UO_181 (O_181,N_4603,N_4895);
and UO_182 (O_182,N_4732,N_4898);
nand UO_183 (O_183,N_4520,N_4572);
nor UO_184 (O_184,N_4880,N_4713);
nand UO_185 (O_185,N_4560,N_4675);
nor UO_186 (O_186,N_4859,N_4694);
xor UO_187 (O_187,N_4828,N_4625);
nor UO_188 (O_188,N_4629,N_4995);
nand UO_189 (O_189,N_4519,N_4983);
nor UO_190 (O_190,N_4803,N_4696);
or UO_191 (O_191,N_4811,N_4568);
nor UO_192 (O_192,N_4751,N_4834);
nor UO_193 (O_193,N_4730,N_4831);
and UO_194 (O_194,N_4651,N_4864);
nand UO_195 (O_195,N_4992,N_4584);
or UO_196 (O_196,N_4745,N_4548);
and UO_197 (O_197,N_4912,N_4546);
or UO_198 (O_198,N_4882,N_4670);
or UO_199 (O_199,N_4900,N_4720);
and UO_200 (O_200,N_4506,N_4956);
nand UO_201 (O_201,N_4855,N_4941);
nor UO_202 (O_202,N_4926,N_4729);
or UO_203 (O_203,N_4712,N_4647);
nor UO_204 (O_204,N_4685,N_4928);
nand UO_205 (O_205,N_4980,N_4547);
nand UO_206 (O_206,N_4521,N_4968);
and UO_207 (O_207,N_4682,N_4648);
nor UO_208 (O_208,N_4818,N_4948);
and UO_209 (O_209,N_4971,N_4832);
and UO_210 (O_210,N_4690,N_4607);
or UO_211 (O_211,N_4619,N_4601);
and UO_212 (O_212,N_4823,N_4881);
nor UO_213 (O_213,N_4669,N_4836);
and UO_214 (O_214,N_4608,N_4526);
nor UO_215 (O_215,N_4914,N_4666);
nand UO_216 (O_216,N_4994,N_4798);
nor UO_217 (O_217,N_4930,N_4821);
or UO_218 (O_218,N_4920,N_4827);
and UO_219 (O_219,N_4867,N_4610);
and UO_220 (O_220,N_4622,N_4870);
and UO_221 (O_221,N_4950,N_4943);
nand UO_222 (O_222,N_4985,N_4916);
nor UO_223 (O_223,N_4695,N_4768);
and UO_224 (O_224,N_4772,N_4829);
nand UO_225 (O_225,N_4665,N_4671);
nand UO_226 (O_226,N_4840,N_4613);
nor UO_227 (O_227,N_4598,N_4638);
and UO_228 (O_228,N_4719,N_4639);
nand UO_229 (O_229,N_4577,N_4502);
nor UO_230 (O_230,N_4799,N_4658);
or UO_231 (O_231,N_4723,N_4937);
and UO_232 (O_232,N_4889,N_4981);
and UO_233 (O_233,N_4594,N_4944);
or UO_234 (O_234,N_4847,N_4645);
nor UO_235 (O_235,N_4820,N_4791);
or UO_236 (O_236,N_4835,N_4511);
nand UO_237 (O_237,N_4600,N_4841);
nor UO_238 (O_238,N_4725,N_4879);
nand UO_239 (O_239,N_4776,N_4901);
or UO_240 (O_240,N_4830,N_4957);
and UO_241 (O_241,N_4583,N_4833);
and UO_242 (O_242,N_4760,N_4585);
or UO_243 (O_243,N_4787,N_4646);
nor UO_244 (O_244,N_4575,N_4652);
and UO_245 (O_245,N_4736,N_4757);
nand UO_246 (O_246,N_4962,N_4531);
or UO_247 (O_247,N_4722,N_4659);
nor UO_248 (O_248,N_4754,N_4789);
or UO_249 (O_249,N_4691,N_4863);
nand UO_250 (O_250,N_4560,N_4945);
nand UO_251 (O_251,N_4952,N_4729);
nand UO_252 (O_252,N_4624,N_4639);
and UO_253 (O_253,N_4783,N_4756);
nand UO_254 (O_254,N_4562,N_4644);
or UO_255 (O_255,N_4856,N_4769);
or UO_256 (O_256,N_4872,N_4912);
nand UO_257 (O_257,N_4623,N_4564);
nand UO_258 (O_258,N_4749,N_4595);
nand UO_259 (O_259,N_4659,N_4956);
nor UO_260 (O_260,N_4608,N_4545);
and UO_261 (O_261,N_4853,N_4877);
nor UO_262 (O_262,N_4957,N_4658);
or UO_263 (O_263,N_4976,N_4891);
nor UO_264 (O_264,N_4779,N_4999);
or UO_265 (O_265,N_4927,N_4974);
nor UO_266 (O_266,N_4999,N_4547);
and UO_267 (O_267,N_4670,N_4702);
and UO_268 (O_268,N_4752,N_4853);
nor UO_269 (O_269,N_4560,N_4690);
nor UO_270 (O_270,N_4837,N_4656);
nor UO_271 (O_271,N_4979,N_4631);
or UO_272 (O_272,N_4964,N_4581);
and UO_273 (O_273,N_4963,N_4960);
nand UO_274 (O_274,N_4721,N_4556);
and UO_275 (O_275,N_4635,N_4951);
and UO_276 (O_276,N_4849,N_4664);
nor UO_277 (O_277,N_4928,N_4627);
or UO_278 (O_278,N_4830,N_4719);
xnor UO_279 (O_279,N_4525,N_4746);
and UO_280 (O_280,N_4595,N_4950);
or UO_281 (O_281,N_4539,N_4554);
nor UO_282 (O_282,N_4880,N_4825);
nand UO_283 (O_283,N_4556,N_4698);
nor UO_284 (O_284,N_4859,N_4606);
nor UO_285 (O_285,N_4564,N_4647);
nand UO_286 (O_286,N_4916,N_4594);
or UO_287 (O_287,N_4554,N_4867);
and UO_288 (O_288,N_4510,N_4954);
nand UO_289 (O_289,N_4988,N_4643);
and UO_290 (O_290,N_4989,N_4554);
and UO_291 (O_291,N_4840,N_4837);
nor UO_292 (O_292,N_4583,N_4937);
or UO_293 (O_293,N_4919,N_4631);
nand UO_294 (O_294,N_4661,N_4845);
nand UO_295 (O_295,N_4727,N_4746);
nand UO_296 (O_296,N_4561,N_4960);
nor UO_297 (O_297,N_4958,N_4833);
nand UO_298 (O_298,N_4812,N_4682);
or UO_299 (O_299,N_4985,N_4542);
nor UO_300 (O_300,N_4651,N_4980);
and UO_301 (O_301,N_4544,N_4903);
or UO_302 (O_302,N_4939,N_4597);
nand UO_303 (O_303,N_4634,N_4717);
nor UO_304 (O_304,N_4779,N_4687);
or UO_305 (O_305,N_4753,N_4963);
nor UO_306 (O_306,N_4536,N_4761);
or UO_307 (O_307,N_4682,N_4594);
nor UO_308 (O_308,N_4975,N_4954);
nand UO_309 (O_309,N_4881,N_4641);
nor UO_310 (O_310,N_4785,N_4776);
and UO_311 (O_311,N_4620,N_4854);
nand UO_312 (O_312,N_4865,N_4827);
nand UO_313 (O_313,N_4666,N_4902);
nand UO_314 (O_314,N_4683,N_4599);
and UO_315 (O_315,N_4921,N_4677);
nor UO_316 (O_316,N_4513,N_4848);
nor UO_317 (O_317,N_4860,N_4578);
nand UO_318 (O_318,N_4622,N_4907);
nand UO_319 (O_319,N_4652,N_4833);
nand UO_320 (O_320,N_4602,N_4579);
nand UO_321 (O_321,N_4515,N_4542);
or UO_322 (O_322,N_4718,N_4744);
nor UO_323 (O_323,N_4720,N_4825);
and UO_324 (O_324,N_4597,N_4980);
nand UO_325 (O_325,N_4771,N_4803);
or UO_326 (O_326,N_4917,N_4689);
or UO_327 (O_327,N_4702,N_4799);
and UO_328 (O_328,N_4883,N_4536);
nor UO_329 (O_329,N_4941,N_4977);
nor UO_330 (O_330,N_4537,N_4866);
and UO_331 (O_331,N_4861,N_4789);
nand UO_332 (O_332,N_4749,N_4691);
or UO_333 (O_333,N_4793,N_4729);
xnor UO_334 (O_334,N_4638,N_4832);
and UO_335 (O_335,N_4839,N_4747);
nor UO_336 (O_336,N_4518,N_4995);
and UO_337 (O_337,N_4638,N_4803);
nand UO_338 (O_338,N_4716,N_4664);
and UO_339 (O_339,N_4845,N_4583);
and UO_340 (O_340,N_4703,N_4998);
nor UO_341 (O_341,N_4708,N_4647);
nor UO_342 (O_342,N_4850,N_4801);
nand UO_343 (O_343,N_4621,N_4501);
or UO_344 (O_344,N_4694,N_4858);
or UO_345 (O_345,N_4664,N_4757);
or UO_346 (O_346,N_4858,N_4893);
nor UO_347 (O_347,N_4752,N_4920);
nor UO_348 (O_348,N_4545,N_4740);
nor UO_349 (O_349,N_4930,N_4912);
and UO_350 (O_350,N_4959,N_4700);
nand UO_351 (O_351,N_4708,N_4680);
nor UO_352 (O_352,N_4729,N_4995);
nor UO_353 (O_353,N_4542,N_4732);
and UO_354 (O_354,N_4861,N_4658);
and UO_355 (O_355,N_4581,N_4590);
or UO_356 (O_356,N_4712,N_4919);
or UO_357 (O_357,N_4653,N_4772);
and UO_358 (O_358,N_4989,N_4671);
or UO_359 (O_359,N_4792,N_4845);
and UO_360 (O_360,N_4515,N_4623);
nand UO_361 (O_361,N_4503,N_4959);
nand UO_362 (O_362,N_4679,N_4854);
nand UO_363 (O_363,N_4621,N_4856);
nand UO_364 (O_364,N_4991,N_4921);
xnor UO_365 (O_365,N_4683,N_4525);
and UO_366 (O_366,N_4825,N_4867);
or UO_367 (O_367,N_4911,N_4867);
and UO_368 (O_368,N_4654,N_4981);
and UO_369 (O_369,N_4654,N_4608);
and UO_370 (O_370,N_4657,N_4915);
nor UO_371 (O_371,N_4698,N_4863);
nor UO_372 (O_372,N_4682,N_4913);
nand UO_373 (O_373,N_4953,N_4613);
nand UO_374 (O_374,N_4828,N_4967);
and UO_375 (O_375,N_4929,N_4591);
nand UO_376 (O_376,N_4586,N_4624);
and UO_377 (O_377,N_4802,N_4866);
and UO_378 (O_378,N_4976,N_4832);
nand UO_379 (O_379,N_4722,N_4829);
or UO_380 (O_380,N_4603,N_4528);
nor UO_381 (O_381,N_4560,N_4996);
or UO_382 (O_382,N_4882,N_4836);
nor UO_383 (O_383,N_4733,N_4564);
nor UO_384 (O_384,N_4931,N_4686);
nor UO_385 (O_385,N_4512,N_4809);
or UO_386 (O_386,N_4682,N_4521);
nor UO_387 (O_387,N_4843,N_4940);
or UO_388 (O_388,N_4716,N_4872);
and UO_389 (O_389,N_4511,N_4501);
xor UO_390 (O_390,N_4748,N_4710);
nor UO_391 (O_391,N_4592,N_4914);
or UO_392 (O_392,N_4953,N_4745);
nor UO_393 (O_393,N_4942,N_4786);
and UO_394 (O_394,N_4515,N_4664);
nand UO_395 (O_395,N_4572,N_4595);
nand UO_396 (O_396,N_4531,N_4789);
or UO_397 (O_397,N_4961,N_4685);
or UO_398 (O_398,N_4848,N_4917);
and UO_399 (O_399,N_4620,N_4821);
or UO_400 (O_400,N_4630,N_4609);
and UO_401 (O_401,N_4825,N_4860);
and UO_402 (O_402,N_4964,N_4595);
and UO_403 (O_403,N_4981,N_4799);
nor UO_404 (O_404,N_4714,N_4871);
nor UO_405 (O_405,N_4742,N_4999);
nand UO_406 (O_406,N_4926,N_4777);
nand UO_407 (O_407,N_4962,N_4916);
nor UO_408 (O_408,N_4856,N_4661);
or UO_409 (O_409,N_4568,N_4979);
and UO_410 (O_410,N_4642,N_4893);
nand UO_411 (O_411,N_4835,N_4567);
and UO_412 (O_412,N_4537,N_4738);
or UO_413 (O_413,N_4842,N_4657);
and UO_414 (O_414,N_4533,N_4959);
nor UO_415 (O_415,N_4836,N_4506);
or UO_416 (O_416,N_4701,N_4904);
or UO_417 (O_417,N_4982,N_4845);
xnor UO_418 (O_418,N_4957,N_4511);
or UO_419 (O_419,N_4792,N_4713);
or UO_420 (O_420,N_4555,N_4603);
and UO_421 (O_421,N_4940,N_4515);
and UO_422 (O_422,N_4590,N_4529);
nor UO_423 (O_423,N_4852,N_4883);
and UO_424 (O_424,N_4786,N_4718);
and UO_425 (O_425,N_4580,N_4701);
or UO_426 (O_426,N_4700,N_4982);
nor UO_427 (O_427,N_4670,N_4644);
nor UO_428 (O_428,N_4550,N_4954);
nand UO_429 (O_429,N_4868,N_4685);
nand UO_430 (O_430,N_4620,N_4536);
nand UO_431 (O_431,N_4992,N_4700);
nor UO_432 (O_432,N_4858,N_4556);
or UO_433 (O_433,N_4981,N_4503);
nor UO_434 (O_434,N_4644,N_4580);
or UO_435 (O_435,N_4938,N_4678);
or UO_436 (O_436,N_4772,N_4934);
nor UO_437 (O_437,N_4644,N_4588);
nor UO_438 (O_438,N_4996,N_4947);
or UO_439 (O_439,N_4861,N_4958);
nand UO_440 (O_440,N_4685,N_4752);
or UO_441 (O_441,N_4779,N_4676);
nand UO_442 (O_442,N_4938,N_4939);
nor UO_443 (O_443,N_4804,N_4976);
nand UO_444 (O_444,N_4797,N_4877);
nor UO_445 (O_445,N_4721,N_4550);
and UO_446 (O_446,N_4919,N_4647);
nand UO_447 (O_447,N_4978,N_4564);
nand UO_448 (O_448,N_4643,N_4535);
nand UO_449 (O_449,N_4876,N_4593);
or UO_450 (O_450,N_4569,N_4672);
and UO_451 (O_451,N_4797,N_4847);
nor UO_452 (O_452,N_4729,N_4976);
nand UO_453 (O_453,N_4724,N_4627);
nor UO_454 (O_454,N_4663,N_4507);
or UO_455 (O_455,N_4832,N_4550);
nand UO_456 (O_456,N_4781,N_4759);
and UO_457 (O_457,N_4918,N_4745);
and UO_458 (O_458,N_4525,N_4788);
and UO_459 (O_459,N_4989,N_4633);
or UO_460 (O_460,N_4586,N_4836);
and UO_461 (O_461,N_4682,N_4746);
nor UO_462 (O_462,N_4827,N_4662);
nor UO_463 (O_463,N_4708,N_4640);
or UO_464 (O_464,N_4981,N_4644);
and UO_465 (O_465,N_4618,N_4635);
xnor UO_466 (O_466,N_4850,N_4859);
nand UO_467 (O_467,N_4982,N_4751);
and UO_468 (O_468,N_4639,N_4621);
nand UO_469 (O_469,N_4914,N_4915);
or UO_470 (O_470,N_4871,N_4874);
nand UO_471 (O_471,N_4799,N_4554);
nand UO_472 (O_472,N_4996,N_4610);
nand UO_473 (O_473,N_4869,N_4556);
nor UO_474 (O_474,N_4678,N_4889);
and UO_475 (O_475,N_4822,N_4929);
nor UO_476 (O_476,N_4960,N_4582);
and UO_477 (O_477,N_4990,N_4662);
nand UO_478 (O_478,N_4713,N_4689);
and UO_479 (O_479,N_4910,N_4694);
or UO_480 (O_480,N_4993,N_4923);
or UO_481 (O_481,N_4756,N_4546);
or UO_482 (O_482,N_4639,N_4783);
nor UO_483 (O_483,N_4637,N_4854);
nand UO_484 (O_484,N_4735,N_4971);
and UO_485 (O_485,N_4989,N_4640);
nand UO_486 (O_486,N_4738,N_4544);
nor UO_487 (O_487,N_4576,N_4641);
nand UO_488 (O_488,N_4562,N_4732);
nor UO_489 (O_489,N_4897,N_4536);
and UO_490 (O_490,N_4763,N_4725);
nand UO_491 (O_491,N_4601,N_4774);
and UO_492 (O_492,N_4654,N_4548);
and UO_493 (O_493,N_4790,N_4787);
nand UO_494 (O_494,N_4635,N_4525);
and UO_495 (O_495,N_4787,N_4502);
or UO_496 (O_496,N_4895,N_4759);
nand UO_497 (O_497,N_4527,N_4629);
and UO_498 (O_498,N_4669,N_4939);
nand UO_499 (O_499,N_4507,N_4757);
or UO_500 (O_500,N_4707,N_4563);
and UO_501 (O_501,N_4780,N_4876);
nor UO_502 (O_502,N_4715,N_4891);
nor UO_503 (O_503,N_4816,N_4713);
or UO_504 (O_504,N_4672,N_4969);
and UO_505 (O_505,N_4777,N_4606);
xor UO_506 (O_506,N_4855,N_4598);
nand UO_507 (O_507,N_4637,N_4950);
nor UO_508 (O_508,N_4785,N_4919);
or UO_509 (O_509,N_4834,N_4889);
or UO_510 (O_510,N_4640,N_4523);
nor UO_511 (O_511,N_4906,N_4522);
nor UO_512 (O_512,N_4806,N_4884);
or UO_513 (O_513,N_4607,N_4705);
and UO_514 (O_514,N_4777,N_4960);
and UO_515 (O_515,N_4867,N_4738);
nand UO_516 (O_516,N_4807,N_4776);
nor UO_517 (O_517,N_4510,N_4513);
and UO_518 (O_518,N_4531,N_4671);
or UO_519 (O_519,N_4903,N_4512);
nor UO_520 (O_520,N_4606,N_4602);
nand UO_521 (O_521,N_4505,N_4785);
or UO_522 (O_522,N_4590,N_4530);
nand UO_523 (O_523,N_4863,N_4532);
nor UO_524 (O_524,N_4817,N_4969);
nand UO_525 (O_525,N_4668,N_4707);
and UO_526 (O_526,N_4572,N_4707);
and UO_527 (O_527,N_4568,N_4729);
nand UO_528 (O_528,N_4537,N_4970);
nand UO_529 (O_529,N_4736,N_4536);
and UO_530 (O_530,N_4751,N_4804);
nor UO_531 (O_531,N_4857,N_4602);
or UO_532 (O_532,N_4849,N_4807);
nor UO_533 (O_533,N_4609,N_4626);
and UO_534 (O_534,N_4678,N_4891);
nor UO_535 (O_535,N_4834,N_4878);
and UO_536 (O_536,N_4969,N_4976);
and UO_537 (O_537,N_4763,N_4778);
nor UO_538 (O_538,N_4836,N_4952);
or UO_539 (O_539,N_4921,N_4912);
xor UO_540 (O_540,N_4702,N_4811);
nor UO_541 (O_541,N_4849,N_4648);
or UO_542 (O_542,N_4767,N_4988);
or UO_543 (O_543,N_4822,N_4813);
nor UO_544 (O_544,N_4665,N_4641);
nor UO_545 (O_545,N_4953,N_4814);
and UO_546 (O_546,N_4893,N_4775);
or UO_547 (O_547,N_4507,N_4613);
or UO_548 (O_548,N_4510,N_4759);
or UO_549 (O_549,N_4995,N_4685);
and UO_550 (O_550,N_4673,N_4755);
or UO_551 (O_551,N_4614,N_4592);
and UO_552 (O_552,N_4522,N_4795);
and UO_553 (O_553,N_4524,N_4519);
and UO_554 (O_554,N_4745,N_4655);
nor UO_555 (O_555,N_4786,N_4536);
nand UO_556 (O_556,N_4651,N_4737);
nand UO_557 (O_557,N_4756,N_4568);
nand UO_558 (O_558,N_4688,N_4736);
nand UO_559 (O_559,N_4827,N_4639);
or UO_560 (O_560,N_4670,N_4729);
and UO_561 (O_561,N_4967,N_4693);
and UO_562 (O_562,N_4944,N_4537);
and UO_563 (O_563,N_4574,N_4518);
and UO_564 (O_564,N_4569,N_4836);
and UO_565 (O_565,N_4502,N_4742);
nand UO_566 (O_566,N_4923,N_4515);
or UO_567 (O_567,N_4683,N_4953);
or UO_568 (O_568,N_4819,N_4716);
or UO_569 (O_569,N_4598,N_4537);
xor UO_570 (O_570,N_4610,N_4539);
nor UO_571 (O_571,N_4796,N_4937);
or UO_572 (O_572,N_4910,N_4544);
and UO_573 (O_573,N_4855,N_4521);
or UO_574 (O_574,N_4995,N_4846);
nand UO_575 (O_575,N_4641,N_4733);
or UO_576 (O_576,N_4751,N_4767);
and UO_577 (O_577,N_4739,N_4702);
nor UO_578 (O_578,N_4761,N_4838);
nor UO_579 (O_579,N_4564,N_4793);
and UO_580 (O_580,N_4869,N_4785);
nor UO_581 (O_581,N_4586,N_4998);
nand UO_582 (O_582,N_4654,N_4927);
or UO_583 (O_583,N_4509,N_4831);
and UO_584 (O_584,N_4858,N_4537);
or UO_585 (O_585,N_4526,N_4538);
nor UO_586 (O_586,N_4703,N_4981);
and UO_587 (O_587,N_4868,N_4886);
and UO_588 (O_588,N_4896,N_4613);
nor UO_589 (O_589,N_4679,N_4638);
nor UO_590 (O_590,N_4722,N_4696);
nand UO_591 (O_591,N_4803,N_4779);
nand UO_592 (O_592,N_4687,N_4904);
nand UO_593 (O_593,N_4988,N_4620);
nor UO_594 (O_594,N_4987,N_4604);
nor UO_595 (O_595,N_4896,N_4504);
and UO_596 (O_596,N_4839,N_4645);
or UO_597 (O_597,N_4588,N_4707);
and UO_598 (O_598,N_4603,N_4553);
nand UO_599 (O_599,N_4997,N_4758);
or UO_600 (O_600,N_4574,N_4898);
nand UO_601 (O_601,N_4622,N_4943);
nor UO_602 (O_602,N_4657,N_4512);
or UO_603 (O_603,N_4805,N_4809);
nand UO_604 (O_604,N_4963,N_4613);
or UO_605 (O_605,N_4809,N_4573);
nor UO_606 (O_606,N_4875,N_4779);
nand UO_607 (O_607,N_4824,N_4792);
nand UO_608 (O_608,N_4972,N_4861);
nand UO_609 (O_609,N_4601,N_4902);
or UO_610 (O_610,N_4623,N_4779);
or UO_611 (O_611,N_4782,N_4669);
nand UO_612 (O_612,N_4840,N_4928);
nand UO_613 (O_613,N_4941,N_4932);
nor UO_614 (O_614,N_4932,N_4683);
nor UO_615 (O_615,N_4934,N_4952);
nor UO_616 (O_616,N_4833,N_4657);
nor UO_617 (O_617,N_4696,N_4530);
nor UO_618 (O_618,N_4952,N_4863);
or UO_619 (O_619,N_4697,N_4614);
nand UO_620 (O_620,N_4820,N_4921);
nand UO_621 (O_621,N_4680,N_4518);
xor UO_622 (O_622,N_4974,N_4830);
nand UO_623 (O_623,N_4657,N_4554);
nand UO_624 (O_624,N_4764,N_4773);
and UO_625 (O_625,N_4746,N_4879);
nor UO_626 (O_626,N_4963,N_4527);
and UO_627 (O_627,N_4989,N_4659);
nand UO_628 (O_628,N_4642,N_4894);
and UO_629 (O_629,N_4784,N_4823);
nand UO_630 (O_630,N_4702,N_4614);
nand UO_631 (O_631,N_4967,N_4648);
or UO_632 (O_632,N_4946,N_4774);
nand UO_633 (O_633,N_4762,N_4752);
or UO_634 (O_634,N_4819,N_4857);
xor UO_635 (O_635,N_4692,N_4985);
nor UO_636 (O_636,N_4974,N_4627);
or UO_637 (O_637,N_4981,N_4767);
xor UO_638 (O_638,N_4643,N_4508);
nand UO_639 (O_639,N_4838,N_4587);
nor UO_640 (O_640,N_4969,N_4914);
and UO_641 (O_641,N_4772,N_4563);
or UO_642 (O_642,N_4701,N_4810);
or UO_643 (O_643,N_4807,N_4767);
or UO_644 (O_644,N_4867,N_4676);
xnor UO_645 (O_645,N_4965,N_4533);
xnor UO_646 (O_646,N_4813,N_4732);
or UO_647 (O_647,N_4975,N_4998);
and UO_648 (O_648,N_4929,N_4992);
and UO_649 (O_649,N_4925,N_4751);
nor UO_650 (O_650,N_4758,N_4588);
nand UO_651 (O_651,N_4993,N_4860);
and UO_652 (O_652,N_4715,N_4912);
nor UO_653 (O_653,N_4736,N_4907);
or UO_654 (O_654,N_4765,N_4753);
or UO_655 (O_655,N_4812,N_4827);
nand UO_656 (O_656,N_4830,N_4747);
or UO_657 (O_657,N_4599,N_4781);
nor UO_658 (O_658,N_4997,N_4561);
and UO_659 (O_659,N_4759,N_4593);
or UO_660 (O_660,N_4938,N_4888);
or UO_661 (O_661,N_4614,N_4803);
nor UO_662 (O_662,N_4674,N_4851);
nor UO_663 (O_663,N_4921,N_4581);
nor UO_664 (O_664,N_4745,N_4607);
xnor UO_665 (O_665,N_4666,N_4899);
nor UO_666 (O_666,N_4596,N_4968);
nand UO_667 (O_667,N_4619,N_4551);
nor UO_668 (O_668,N_4549,N_4568);
xor UO_669 (O_669,N_4836,N_4875);
or UO_670 (O_670,N_4632,N_4551);
and UO_671 (O_671,N_4608,N_4880);
nor UO_672 (O_672,N_4507,N_4981);
or UO_673 (O_673,N_4794,N_4542);
nand UO_674 (O_674,N_4510,N_4972);
and UO_675 (O_675,N_4706,N_4952);
or UO_676 (O_676,N_4900,N_4990);
nor UO_677 (O_677,N_4682,N_4672);
nand UO_678 (O_678,N_4867,N_4669);
nand UO_679 (O_679,N_4941,N_4646);
xnor UO_680 (O_680,N_4760,N_4874);
nor UO_681 (O_681,N_4573,N_4553);
nand UO_682 (O_682,N_4859,N_4965);
nor UO_683 (O_683,N_4707,N_4710);
nand UO_684 (O_684,N_4613,N_4978);
or UO_685 (O_685,N_4577,N_4737);
nand UO_686 (O_686,N_4806,N_4557);
or UO_687 (O_687,N_4664,N_4685);
nand UO_688 (O_688,N_4593,N_4542);
nand UO_689 (O_689,N_4560,N_4707);
nor UO_690 (O_690,N_4544,N_4775);
or UO_691 (O_691,N_4935,N_4771);
and UO_692 (O_692,N_4681,N_4662);
xor UO_693 (O_693,N_4588,N_4869);
nor UO_694 (O_694,N_4812,N_4548);
or UO_695 (O_695,N_4930,N_4684);
and UO_696 (O_696,N_4742,N_4641);
and UO_697 (O_697,N_4837,N_4666);
nand UO_698 (O_698,N_4645,N_4572);
nand UO_699 (O_699,N_4680,N_4715);
or UO_700 (O_700,N_4766,N_4630);
and UO_701 (O_701,N_4703,N_4582);
or UO_702 (O_702,N_4514,N_4559);
nand UO_703 (O_703,N_4764,N_4587);
nand UO_704 (O_704,N_4662,N_4838);
and UO_705 (O_705,N_4856,N_4933);
or UO_706 (O_706,N_4724,N_4921);
xor UO_707 (O_707,N_4725,N_4559);
and UO_708 (O_708,N_4822,N_4512);
and UO_709 (O_709,N_4891,N_4792);
nand UO_710 (O_710,N_4750,N_4505);
and UO_711 (O_711,N_4650,N_4711);
nand UO_712 (O_712,N_4848,N_4534);
and UO_713 (O_713,N_4861,N_4920);
nor UO_714 (O_714,N_4666,N_4501);
and UO_715 (O_715,N_4636,N_4573);
nor UO_716 (O_716,N_4915,N_4908);
nand UO_717 (O_717,N_4601,N_4718);
or UO_718 (O_718,N_4659,N_4526);
nor UO_719 (O_719,N_4551,N_4980);
and UO_720 (O_720,N_4668,N_4511);
nand UO_721 (O_721,N_4929,N_4631);
and UO_722 (O_722,N_4668,N_4805);
or UO_723 (O_723,N_4638,N_4978);
and UO_724 (O_724,N_4675,N_4719);
and UO_725 (O_725,N_4585,N_4845);
nor UO_726 (O_726,N_4580,N_4611);
or UO_727 (O_727,N_4750,N_4749);
nand UO_728 (O_728,N_4631,N_4516);
nor UO_729 (O_729,N_4913,N_4713);
or UO_730 (O_730,N_4973,N_4570);
nor UO_731 (O_731,N_4673,N_4845);
and UO_732 (O_732,N_4699,N_4891);
or UO_733 (O_733,N_4904,N_4969);
nor UO_734 (O_734,N_4654,N_4944);
nor UO_735 (O_735,N_4567,N_4862);
and UO_736 (O_736,N_4835,N_4766);
nor UO_737 (O_737,N_4704,N_4701);
nor UO_738 (O_738,N_4508,N_4677);
or UO_739 (O_739,N_4700,N_4774);
and UO_740 (O_740,N_4898,N_4782);
nand UO_741 (O_741,N_4690,N_4614);
nor UO_742 (O_742,N_4915,N_4899);
nand UO_743 (O_743,N_4789,N_4939);
nor UO_744 (O_744,N_4683,N_4846);
or UO_745 (O_745,N_4516,N_4605);
nor UO_746 (O_746,N_4921,N_4854);
or UO_747 (O_747,N_4845,N_4681);
and UO_748 (O_748,N_4892,N_4567);
nor UO_749 (O_749,N_4733,N_4872);
and UO_750 (O_750,N_4638,N_4608);
nand UO_751 (O_751,N_4967,N_4709);
or UO_752 (O_752,N_4727,N_4784);
and UO_753 (O_753,N_4847,N_4542);
nor UO_754 (O_754,N_4908,N_4921);
nand UO_755 (O_755,N_4587,N_4872);
or UO_756 (O_756,N_4693,N_4549);
and UO_757 (O_757,N_4759,N_4631);
or UO_758 (O_758,N_4816,N_4594);
and UO_759 (O_759,N_4913,N_4724);
xor UO_760 (O_760,N_4748,N_4554);
or UO_761 (O_761,N_4689,N_4696);
and UO_762 (O_762,N_4517,N_4943);
and UO_763 (O_763,N_4754,N_4776);
nand UO_764 (O_764,N_4990,N_4542);
nor UO_765 (O_765,N_4731,N_4810);
and UO_766 (O_766,N_4527,N_4648);
nand UO_767 (O_767,N_4748,N_4770);
nand UO_768 (O_768,N_4884,N_4519);
or UO_769 (O_769,N_4634,N_4743);
nand UO_770 (O_770,N_4681,N_4595);
and UO_771 (O_771,N_4797,N_4627);
or UO_772 (O_772,N_4512,N_4990);
nand UO_773 (O_773,N_4522,N_4743);
and UO_774 (O_774,N_4586,N_4578);
nor UO_775 (O_775,N_4803,N_4539);
or UO_776 (O_776,N_4898,N_4588);
nor UO_777 (O_777,N_4978,N_4870);
xnor UO_778 (O_778,N_4896,N_4826);
or UO_779 (O_779,N_4832,N_4762);
and UO_780 (O_780,N_4889,N_4677);
or UO_781 (O_781,N_4659,N_4742);
nor UO_782 (O_782,N_4980,N_4809);
or UO_783 (O_783,N_4946,N_4823);
or UO_784 (O_784,N_4989,N_4756);
and UO_785 (O_785,N_4671,N_4851);
nand UO_786 (O_786,N_4523,N_4778);
or UO_787 (O_787,N_4742,N_4598);
and UO_788 (O_788,N_4503,N_4542);
or UO_789 (O_789,N_4962,N_4511);
and UO_790 (O_790,N_4797,N_4604);
or UO_791 (O_791,N_4791,N_4587);
nand UO_792 (O_792,N_4740,N_4757);
and UO_793 (O_793,N_4520,N_4778);
and UO_794 (O_794,N_4984,N_4648);
nand UO_795 (O_795,N_4827,N_4702);
or UO_796 (O_796,N_4697,N_4547);
and UO_797 (O_797,N_4568,N_4551);
or UO_798 (O_798,N_4967,N_4583);
nor UO_799 (O_799,N_4579,N_4545);
nor UO_800 (O_800,N_4822,N_4515);
or UO_801 (O_801,N_4988,N_4715);
or UO_802 (O_802,N_4921,N_4748);
and UO_803 (O_803,N_4845,N_4623);
and UO_804 (O_804,N_4733,N_4998);
nor UO_805 (O_805,N_4607,N_4875);
or UO_806 (O_806,N_4587,N_4858);
nand UO_807 (O_807,N_4708,N_4984);
nor UO_808 (O_808,N_4918,N_4926);
nor UO_809 (O_809,N_4601,N_4763);
or UO_810 (O_810,N_4517,N_4592);
nand UO_811 (O_811,N_4935,N_4956);
nand UO_812 (O_812,N_4561,N_4900);
nor UO_813 (O_813,N_4932,N_4608);
or UO_814 (O_814,N_4722,N_4665);
or UO_815 (O_815,N_4774,N_4880);
nor UO_816 (O_816,N_4775,N_4989);
nor UO_817 (O_817,N_4997,N_4579);
or UO_818 (O_818,N_4786,N_4602);
nor UO_819 (O_819,N_4532,N_4836);
nor UO_820 (O_820,N_4513,N_4949);
or UO_821 (O_821,N_4854,N_4720);
and UO_822 (O_822,N_4568,N_4623);
or UO_823 (O_823,N_4736,N_4602);
or UO_824 (O_824,N_4531,N_4607);
xor UO_825 (O_825,N_4632,N_4879);
and UO_826 (O_826,N_4824,N_4850);
nor UO_827 (O_827,N_4753,N_4998);
nand UO_828 (O_828,N_4532,N_4577);
or UO_829 (O_829,N_4657,N_4782);
nor UO_830 (O_830,N_4669,N_4881);
nor UO_831 (O_831,N_4915,N_4668);
xor UO_832 (O_832,N_4997,N_4708);
or UO_833 (O_833,N_4813,N_4976);
or UO_834 (O_834,N_4655,N_4652);
or UO_835 (O_835,N_4590,N_4803);
or UO_836 (O_836,N_4745,N_4860);
xnor UO_837 (O_837,N_4541,N_4531);
nor UO_838 (O_838,N_4781,N_4694);
nor UO_839 (O_839,N_4746,N_4763);
nand UO_840 (O_840,N_4612,N_4588);
nand UO_841 (O_841,N_4992,N_4798);
or UO_842 (O_842,N_4906,N_4927);
or UO_843 (O_843,N_4960,N_4834);
nor UO_844 (O_844,N_4750,N_4502);
nand UO_845 (O_845,N_4950,N_4737);
nor UO_846 (O_846,N_4609,N_4577);
or UO_847 (O_847,N_4624,N_4655);
nor UO_848 (O_848,N_4649,N_4505);
nand UO_849 (O_849,N_4812,N_4940);
or UO_850 (O_850,N_4774,N_4792);
nor UO_851 (O_851,N_4718,N_4570);
nor UO_852 (O_852,N_4717,N_4797);
nand UO_853 (O_853,N_4974,N_4681);
or UO_854 (O_854,N_4927,N_4668);
or UO_855 (O_855,N_4588,N_4682);
xor UO_856 (O_856,N_4688,N_4760);
and UO_857 (O_857,N_4595,N_4765);
nor UO_858 (O_858,N_4546,N_4599);
nor UO_859 (O_859,N_4899,N_4896);
or UO_860 (O_860,N_4782,N_4541);
nand UO_861 (O_861,N_4818,N_4612);
and UO_862 (O_862,N_4940,N_4780);
and UO_863 (O_863,N_4525,N_4557);
nor UO_864 (O_864,N_4536,N_4776);
nor UO_865 (O_865,N_4635,N_4882);
xnor UO_866 (O_866,N_4800,N_4926);
nand UO_867 (O_867,N_4941,N_4544);
nand UO_868 (O_868,N_4810,N_4840);
or UO_869 (O_869,N_4963,N_4820);
nor UO_870 (O_870,N_4870,N_4535);
or UO_871 (O_871,N_4678,N_4706);
and UO_872 (O_872,N_4730,N_4945);
or UO_873 (O_873,N_4623,N_4833);
or UO_874 (O_874,N_4998,N_4524);
and UO_875 (O_875,N_4594,N_4538);
and UO_876 (O_876,N_4648,N_4555);
nand UO_877 (O_877,N_4570,N_4931);
nor UO_878 (O_878,N_4701,N_4859);
or UO_879 (O_879,N_4695,N_4575);
nor UO_880 (O_880,N_4614,N_4975);
or UO_881 (O_881,N_4793,N_4890);
nand UO_882 (O_882,N_4993,N_4951);
nand UO_883 (O_883,N_4876,N_4897);
or UO_884 (O_884,N_4744,N_4824);
and UO_885 (O_885,N_4972,N_4974);
and UO_886 (O_886,N_4740,N_4655);
nor UO_887 (O_887,N_4649,N_4798);
and UO_888 (O_888,N_4758,N_4770);
and UO_889 (O_889,N_4644,N_4802);
nor UO_890 (O_890,N_4564,N_4804);
or UO_891 (O_891,N_4516,N_4896);
xor UO_892 (O_892,N_4705,N_4577);
or UO_893 (O_893,N_4582,N_4559);
or UO_894 (O_894,N_4908,N_4747);
nand UO_895 (O_895,N_4556,N_4826);
or UO_896 (O_896,N_4582,N_4915);
nand UO_897 (O_897,N_4632,N_4846);
nand UO_898 (O_898,N_4512,N_4908);
or UO_899 (O_899,N_4979,N_4542);
nor UO_900 (O_900,N_4569,N_4943);
or UO_901 (O_901,N_4859,N_4910);
nand UO_902 (O_902,N_4985,N_4849);
and UO_903 (O_903,N_4547,N_4559);
or UO_904 (O_904,N_4597,N_4864);
nor UO_905 (O_905,N_4584,N_4746);
nand UO_906 (O_906,N_4583,N_4777);
or UO_907 (O_907,N_4798,N_4579);
nand UO_908 (O_908,N_4963,N_4935);
or UO_909 (O_909,N_4834,N_4535);
or UO_910 (O_910,N_4675,N_4723);
nand UO_911 (O_911,N_4570,N_4819);
or UO_912 (O_912,N_4973,N_4631);
nor UO_913 (O_913,N_4863,N_4554);
nand UO_914 (O_914,N_4878,N_4818);
nand UO_915 (O_915,N_4584,N_4991);
nor UO_916 (O_916,N_4675,N_4987);
nand UO_917 (O_917,N_4965,N_4563);
and UO_918 (O_918,N_4874,N_4511);
nor UO_919 (O_919,N_4598,N_4688);
nand UO_920 (O_920,N_4710,N_4708);
nand UO_921 (O_921,N_4862,N_4831);
nand UO_922 (O_922,N_4789,N_4866);
and UO_923 (O_923,N_4975,N_4596);
and UO_924 (O_924,N_4689,N_4639);
nor UO_925 (O_925,N_4984,N_4527);
or UO_926 (O_926,N_4732,N_4986);
and UO_927 (O_927,N_4582,N_4999);
or UO_928 (O_928,N_4532,N_4870);
and UO_929 (O_929,N_4503,N_4833);
nor UO_930 (O_930,N_4998,N_4873);
and UO_931 (O_931,N_4571,N_4666);
and UO_932 (O_932,N_4850,N_4718);
nor UO_933 (O_933,N_4948,N_4902);
nor UO_934 (O_934,N_4543,N_4792);
nor UO_935 (O_935,N_4862,N_4532);
nand UO_936 (O_936,N_4501,N_4702);
and UO_937 (O_937,N_4994,N_4512);
and UO_938 (O_938,N_4572,N_4552);
or UO_939 (O_939,N_4964,N_4858);
or UO_940 (O_940,N_4583,N_4553);
nor UO_941 (O_941,N_4941,N_4838);
nor UO_942 (O_942,N_4792,N_4795);
nand UO_943 (O_943,N_4778,N_4695);
nor UO_944 (O_944,N_4628,N_4505);
nor UO_945 (O_945,N_4979,N_4960);
nand UO_946 (O_946,N_4574,N_4792);
or UO_947 (O_947,N_4970,N_4665);
or UO_948 (O_948,N_4921,N_4602);
nor UO_949 (O_949,N_4745,N_4729);
nor UO_950 (O_950,N_4709,N_4556);
xnor UO_951 (O_951,N_4837,N_4883);
nand UO_952 (O_952,N_4535,N_4678);
and UO_953 (O_953,N_4768,N_4509);
or UO_954 (O_954,N_4959,N_4991);
and UO_955 (O_955,N_4918,N_4912);
or UO_956 (O_956,N_4864,N_4673);
nand UO_957 (O_957,N_4644,N_4617);
nor UO_958 (O_958,N_4942,N_4879);
nor UO_959 (O_959,N_4660,N_4535);
nand UO_960 (O_960,N_4560,N_4994);
or UO_961 (O_961,N_4630,N_4516);
nand UO_962 (O_962,N_4670,N_4536);
nor UO_963 (O_963,N_4736,N_4571);
or UO_964 (O_964,N_4547,N_4700);
and UO_965 (O_965,N_4986,N_4729);
and UO_966 (O_966,N_4825,N_4946);
xor UO_967 (O_967,N_4612,N_4648);
and UO_968 (O_968,N_4993,N_4746);
nor UO_969 (O_969,N_4813,N_4957);
and UO_970 (O_970,N_4596,N_4858);
or UO_971 (O_971,N_4693,N_4844);
or UO_972 (O_972,N_4808,N_4917);
or UO_973 (O_973,N_4578,N_4837);
and UO_974 (O_974,N_4614,N_4863);
or UO_975 (O_975,N_4636,N_4578);
nor UO_976 (O_976,N_4773,N_4976);
nor UO_977 (O_977,N_4756,N_4875);
and UO_978 (O_978,N_4871,N_4823);
nand UO_979 (O_979,N_4676,N_4501);
nor UO_980 (O_980,N_4655,N_4893);
and UO_981 (O_981,N_4868,N_4708);
or UO_982 (O_982,N_4608,N_4670);
xor UO_983 (O_983,N_4937,N_4831);
or UO_984 (O_984,N_4923,N_4770);
nand UO_985 (O_985,N_4968,N_4547);
nor UO_986 (O_986,N_4748,N_4520);
or UO_987 (O_987,N_4955,N_4978);
nor UO_988 (O_988,N_4552,N_4779);
nand UO_989 (O_989,N_4768,N_4952);
and UO_990 (O_990,N_4882,N_4915);
and UO_991 (O_991,N_4552,N_4803);
and UO_992 (O_992,N_4680,N_4853);
or UO_993 (O_993,N_4630,N_4746);
nor UO_994 (O_994,N_4804,N_4928);
or UO_995 (O_995,N_4778,N_4760);
nor UO_996 (O_996,N_4577,N_4834);
and UO_997 (O_997,N_4834,N_4573);
and UO_998 (O_998,N_4933,N_4684);
nor UO_999 (O_999,N_4820,N_4833);
endmodule