module basic_1000_10000_1500_2_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5003,N_5005,N_5007,N_5008,N_5009,N_5010,N_5012,N_5016,N_5019,N_5020,N_5021,N_5024,N_5025,N_5026,N_5027,N_5029,N_5030,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5040,N_5043,N_5044,N_5045,N_5046,N_5048,N_5050,N_5051,N_5052,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5061,N_5062,N_5064,N_5065,N_5068,N_5072,N_5073,N_5074,N_5076,N_5077,N_5078,N_5079,N_5080,N_5082,N_5084,N_5085,N_5086,N_5087,N_5089,N_5091,N_5092,N_5093,N_5095,N_5097,N_5100,N_5101,N_5102,N_5103,N_5104,N_5108,N_5109,N_5110,N_5111,N_5114,N_5115,N_5118,N_5120,N_5121,N_5122,N_5126,N_5128,N_5130,N_5131,N_5134,N_5135,N_5136,N_5138,N_5139,N_5140,N_5142,N_5144,N_5145,N_5147,N_5148,N_5150,N_5151,N_5152,N_5153,N_5155,N_5157,N_5159,N_5161,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5172,N_5174,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5184,N_5185,N_5186,N_5188,N_5191,N_5193,N_5195,N_5197,N_5198,N_5201,N_5204,N_5206,N_5212,N_5213,N_5214,N_5215,N_5216,N_5218,N_5219,N_5220,N_5221,N_5222,N_5224,N_5225,N_5226,N_5231,N_5232,N_5233,N_5235,N_5236,N_5237,N_5238,N_5240,N_5243,N_5245,N_5249,N_5250,N_5255,N_5256,N_5257,N_5259,N_5260,N_5261,N_5263,N_5264,N_5266,N_5267,N_5270,N_5271,N_5273,N_5274,N_5275,N_5276,N_5278,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5292,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5305,N_5306,N_5309,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5320,N_5322,N_5324,N_5326,N_5327,N_5328,N_5330,N_5332,N_5333,N_5335,N_5336,N_5337,N_5338,N_5341,N_5342,N_5346,N_5349,N_5350,N_5352,N_5354,N_5355,N_5357,N_5358,N_5359,N_5361,N_5362,N_5363,N_5364,N_5365,N_5368,N_5369,N_5370,N_5371,N_5374,N_5375,N_5376,N_5379,N_5381,N_5382,N_5383,N_5384,N_5385,N_5387,N_5389,N_5390,N_5392,N_5393,N_5394,N_5397,N_5399,N_5401,N_5402,N_5403,N_5404,N_5405,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5420,N_5422,N_5423,N_5424,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5436,N_5437,N_5441,N_5442,N_5443,N_5448,N_5449,N_5450,N_5453,N_5459,N_5460,N_5461,N_5463,N_5468,N_5469,N_5470,N_5471,N_5473,N_5476,N_5478,N_5479,N_5480,N_5482,N_5485,N_5486,N_5487,N_5489,N_5492,N_5493,N_5494,N_5495,N_5496,N_5498,N_5499,N_5500,N_5502,N_5503,N_5504,N_5505,N_5506,N_5508,N_5509,N_5511,N_5512,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5523,N_5527,N_5529,N_5531,N_5533,N_5537,N_5539,N_5540,N_5541,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5553,N_5554,N_5558,N_5560,N_5561,N_5563,N_5565,N_5570,N_5571,N_5572,N_5573,N_5575,N_5576,N_5577,N_5578,N_5579,N_5583,N_5584,N_5586,N_5588,N_5589,N_5590,N_5592,N_5594,N_5597,N_5601,N_5602,N_5603,N_5606,N_5607,N_5609,N_5610,N_5611,N_5612,N_5613,N_5616,N_5621,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5634,N_5635,N_5636,N_5637,N_5641,N_5644,N_5646,N_5648,N_5650,N_5651,N_5653,N_5654,N_5655,N_5658,N_5662,N_5664,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5677,N_5678,N_5679,N_5687,N_5688,N_5690,N_5692,N_5701,N_5702,N_5704,N_5705,N_5706,N_5707,N_5712,N_5715,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5724,N_5727,N_5729,N_5730,N_5731,N_5733,N_5734,N_5735,N_5737,N_5739,N_5741,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5752,N_5753,N_5754,N_5755,N_5757,N_5758,N_5760,N_5761,N_5762,N_5764,N_5765,N_5767,N_5771,N_5773,N_5774,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5797,N_5802,N_5804,N_5807,N_5809,N_5810,N_5811,N_5814,N_5815,N_5817,N_5820,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5829,N_5831,N_5832,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5844,N_5845,N_5848,N_5849,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5868,N_5873,N_5875,N_5876,N_5877,N_5879,N_5880,N_5882,N_5883,N_5885,N_5886,N_5887,N_5888,N_5890,N_5892,N_5893,N_5894,N_5895,N_5896,N_5898,N_5899,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5908,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5918,N_5919,N_5921,N_5925,N_5927,N_5928,N_5929,N_5933,N_5936,N_5937,N_5938,N_5939,N_5941,N_5943,N_5944,N_5946,N_5948,N_5949,N_5951,N_5952,N_5953,N_5954,N_5955,N_5957,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5966,N_5967,N_5968,N_5970,N_5974,N_5975,N_5977,N_5978,N_5979,N_5980,N_5982,N_5985,N_5986,N_5988,N_5989,N_5994,N_5995,N_5996,N_5999,N_6000,N_6001,N_6002,N_6003,N_6005,N_6006,N_6008,N_6010,N_6013,N_6015,N_6016,N_6017,N_6019,N_6020,N_6023,N_6025,N_6026,N_6027,N_6030,N_6031,N_6035,N_6036,N_6039,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6052,N_6053,N_6054,N_6055,N_6057,N_6058,N_6059,N_6061,N_6062,N_6066,N_6068,N_6069,N_6070,N_6072,N_6074,N_6075,N_6077,N_6078,N_6079,N_6080,N_6081,N_6084,N_6089,N_6090,N_6091,N_6093,N_6094,N_6096,N_6097,N_6098,N_6099,N_6100,N_6104,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6113,N_6114,N_6116,N_6117,N_6120,N_6122,N_6124,N_6125,N_6126,N_6127,N_6129,N_6130,N_6131,N_6134,N_6135,N_6136,N_6138,N_6139,N_6140,N_6142,N_6144,N_6146,N_6148,N_6149,N_6150,N_6152,N_6155,N_6157,N_6159,N_6160,N_6161,N_6162,N_6164,N_6165,N_6166,N_6167,N_6169,N_6170,N_6171,N_6175,N_6176,N_6178,N_6181,N_6182,N_6183,N_6185,N_6186,N_6188,N_6189,N_6191,N_6192,N_6195,N_6198,N_6199,N_6203,N_6204,N_6205,N_6206,N_6207,N_6210,N_6211,N_6213,N_6216,N_6217,N_6218,N_6219,N_6222,N_6224,N_6226,N_6229,N_6230,N_6232,N_6234,N_6236,N_6237,N_6239,N_6240,N_6241,N_6243,N_6244,N_6245,N_6246,N_6248,N_6249,N_6251,N_6252,N_6254,N_6255,N_6256,N_6258,N_6259,N_6260,N_6262,N_6263,N_6264,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6277,N_6278,N_6279,N_6280,N_6282,N_6283,N_6284,N_6285,N_6286,N_6289,N_6290,N_6291,N_6292,N_6294,N_6295,N_6296,N_6297,N_6299,N_6300,N_6301,N_6302,N_6304,N_6306,N_6307,N_6308,N_6312,N_6313,N_6314,N_6318,N_6319,N_6322,N_6323,N_6325,N_6328,N_6329,N_6331,N_6337,N_6339,N_6342,N_6343,N_6345,N_6346,N_6348,N_6349,N_6351,N_6353,N_6354,N_6355,N_6356,N_6358,N_6359,N_6360,N_6361,N_6364,N_6366,N_6367,N_6369,N_6372,N_6373,N_6374,N_6377,N_6378,N_6382,N_6383,N_6385,N_6386,N_6387,N_6388,N_6391,N_6392,N_6395,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6407,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6416,N_6417,N_6418,N_6420,N_6422,N_6423,N_6424,N_6425,N_6427,N_6430,N_6433,N_6434,N_6435,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6448,N_6449,N_6451,N_6453,N_6454,N_6455,N_6457,N_6458,N_6460,N_6461,N_6463,N_6467,N_6469,N_6470,N_6475,N_6476,N_6479,N_6481,N_6484,N_6485,N_6486,N_6487,N_6489,N_6490,N_6492,N_6493,N_6496,N_6497,N_6499,N_6500,N_6504,N_6505,N_6506,N_6507,N_6510,N_6513,N_6515,N_6518,N_6520,N_6522,N_6524,N_6528,N_6529,N_6531,N_6532,N_6533,N_6535,N_6536,N_6537,N_6539,N_6540,N_6541,N_6543,N_6544,N_6545,N_6546,N_6549,N_6550,N_6551,N_6552,N_6554,N_6556,N_6557,N_6558,N_6561,N_6562,N_6563,N_6564,N_6567,N_6569,N_6570,N_6571,N_6575,N_6576,N_6577,N_6578,N_6579,N_6581,N_6584,N_6585,N_6587,N_6589,N_6590,N_6591,N_6592,N_6594,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6606,N_6607,N_6611,N_6612,N_6614,N_6615,N_6617,N_6620,N_6624,N_6627,N_6630,N_6631,N_6633,N_6634,N_6636,N_6640,N_6641,N_6642,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6651,N_6652,N_6654,N_6655,N_6658,N_6659,N_6660,N_6661,N_6663,N_6664,N_6665,N_6666,N_6668,N_6669,N_6671,N_6672,N_6673,N_6674,N_6676,N_6677,N_6678,N_6679,N_6680,N_6682,N_6683,N_6684,N_6685,N_6686,N_6691,N_6696,N_6699,N_6700,N_6704,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6717,N_6718,N_6719,N_6720,N_6726,N_6728,N_6729,N_6731,N_6732,N_6734,N_6735,N_6737,N_6738,N_6739,N_6740,N_6743,N_6744,N_6745,N_6746,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6755,N_6756,N_6757,N_6758,N_6759,N_6761,N_6764,N_6765,N_6767,N_6768,N_6772,N_6773,N_6775,N_6778,N_6780,N_6781,N_6784,N_6786,N_6788,N_6790,N_6793,N_6795,N_6798,N_6800,N_6802,N_6803,N_6805,N_6806,N_6807,N_6808,N_6812,N_6813,N_6814,N_6817,N_6818,N_6819,N_6822,N_6827,N_6828,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6838,N_6840,N_6841,N_6844,N_6846,N_6848,N_6849,N_6850,N_6852,N_6854,N_6856,N_6858,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6867,N_6868,N_6871,N_6872,N_6874,N_6875,N_6876,N_6877,N_6879,N_6880,N_6882,N_6884,N_6887,N_6888,N_6889,N_6890,N_6891,N_6893,N_6894,N_6896,N_6897,N_6899,N_6900,N_6901,N_6902,N_6907,N_6909,N_6910,N_6912,N_6916,N_6917,N_6919,N_6920,N_6921,N_6923,N_6924,N_6925,N_6927,N_6928,N_6929,N_6930,N_6932,N_6933,N_6934,N_6935,N_6937,N_6938,N_6940,N_6942,N_6943,N_6944,N_6945,N_6948,N_6949,N_6951,N_6956,N_6958,N_6961,N_6963,N_6966,N_6967,N_6968,N_6969,N_6970,N_6973,N_6974,N_6975,N_6976,N_6977,N_6979,N_6980,N_6983,N_6984,N_6986,N_6987,N_6989,N_6990,N_6992,N_6993,N_6995,N_6997,N_7000,N_7001,N_7003,N_7004,N_7005,N_7006,N_7010,N_7017,N_7018,N_7019,N_7023,N_7025,N_7026,N_7030,N_7033,N_7034,N_7036,N_7040,N_7041,N_7044,N_7047,N_7048,N_7049,N_7050,N_7052,N_7055,N_7056,N_7057,N_7058,N_7062,N_7063,N_7064,N_7065,N_7067,N_7069,N_7071,N_7076,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7090,N_7091,N_7092,N_7094,N_7095,N_7096,N_7098,N_7100,N_7103,N_7104,N_7107,N_7109,N_7110,N_7112,N_7115,N_7116,N_7117,N_7118,N_7121,N_7125,N_7129,N_7130,N_7131,N_7135,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7150,N_7151,N_7152,N_7153,N_7156,N_7160,N_7161,N_7163,N_7164,N_7165,N_7166,N_7167,N_7169,N_7170,N_7172,N_7173,N_7174,N_7176,N_7179,N_7180,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7189,N_7190,N_7192,N_7193,N_7194,N_7195,N_7198,N_7199,N_7202,N_7204,N_7206,N_7209,N_7210,N_7212,N_7213,N_7214,N_7215,N_7216,N_7221,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7231,N_7233,N_7237,N_7238,N_7240,N_7242,N_7245,N_7250,N_7252,N_7253,N_7254,N_7256,N_7257,N_7258,N_7260,N_7261,N_7262,N_7267,N_7268,N_7269,N_7270,N_7272,N_7278,N_7279,N_7282,N_7283,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7293,N_7294,N_7296,N_7297,N_7298,N_7299,N_7301,N_7302,N_7303,N_7305,N_7309,N_7310,N_7311,N_7313,N_7316,N_7319,N_7320,N_7321,N_7326,N_7328,N_7329,N_7330,N_7331,N_7332,N_7334,N_7336,N_7337,N_7339,N_7340,N_7341,N_7346,N_7347,N_7349,N_7352,N_7353,N_7358,N_7359,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7369,N_7370,N_7371,N_7373,N_7374,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7384,N_7387,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7396,N_7398,N_7399,N_7400,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7411,N_7412,N_7415,N_7417,N_7418,N_7419,N_7420,N_7424,N_7425,N_7426,N_7427,N_7430,N_7431,N_7432,N_7433,N_7436,N_7437,N_7439,N_7440,N_7441,N_7446,N_7447,N_7449,N_7451,N_7452,N_7453,N_7455,N_7457,N_7459,N_7460,N_7461,N_7462,N_7463,N_7468,N_7471,N_7473,N_7475,N_7479,N_7480,N_7481,N_7483,N_7484,N_7486,N_7490,N_7492,N_7493,N_7497,N_7498,N_7499,N_7501,N_7503,N_7504,N_7507,N_7509,N_7511,N_7512,N_7514,N_7515,N_7516,N_7518,N_7519,N_7522,N_7523,N_7526,N_7528,N_7529,N_7531,N_7533,N_7535,N_7537,N_7538,N_7542,N_7545,N_7546,N_7547,N_7548,N_7549,N_7552,N_7553,N_7556,N_7557,N_7558,N_7559,N_7561,N_7562,N_7566,N_7567,N_7568,N_7570,N_7572,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7584,N_7586,N_7588,N_7590,N_7591,N_7594,N_7595,N_7597,N_7599,N_7600,N_7605,N_7606,N_7607,N_7608,N_7611,N_7614,N_7618,N_7620,N_7622,N_7624,N_7625,N_7628,N_7629,N_7630,N_7631,N_7634,N_7635,N_7638,N_7639,N_7640,N_7643,N_7644,N_7645,N_7646,N_7648,N_7650,N_7651,N_7652,N_7653,N_7655,N_7656,N_7657,N_7658,N_7659,N_7661,N_7664,N_7665,N_7666,N_7667,N_7672,N_7673,N_7676,N_7677,N_7678,N_7680,N_7681,N_7685,N_7686,N_7688,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7699,N_7700,N_7701,N_7702,N_7704,N_7705,N_7706,N_7708,N_7709,N_7710,N_7715,N_7717,N_7721,N_7722,N_7723,N_7724,N_7725,N_7727,N_7728,N_7729,N_7731,N_7734,N_7736,N_7737,N_7738,N_7741,N_7742,N_7743,N_7744,N_7745,N_7747,N_7750,N_7752,N_7753,N_7754,N_7756,N_7757,N_7758,N_7761,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7771,N_7772,N_7773,N_7774,N_7775,N_7777,N_7779,N_7780,N_7781,N_7783,N_7784,N_7785,N_7786,N_7790,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7799,N_7800,N_7804,N_7805,N_7807,N_7808,N_7809,N_7811,N_7812,N_7813,N_7814,N_7815,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7824,N_7826,N_7829,N_7830,N_7831,N_7832,N_7834,N_7836,N_7837,N_7838,N_7841,N_7842,N_7843,N_7844,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7859,N_7861,N_7862,N_7864,N_7866,N_7869,N_7870,N_7872,N_7874,N_7875,N_7880,N_7881,N_7883,N_7884,N_7886,N_7887,N_7888,N_7890,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7903,N_7904,N_7905,N_7906,N_7908,N_7910,N_7911,N_7914,N_7915,N_7916,N_7917,N_7920,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7931,N_7932,N_7936,N_7937,N_7938,N_7939,N_7941,N_7943,N_7944,N_7945,N_7947,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7957,N_7958,N_7960,N_7961,N_7963,N_7964,N_7965,N_7967,N_7968,N_7970,N_7971,N_7973,N_7974,N_7975,N_7976,N_7980,N_7983,N_7984,N_7985,N_7988,N_7990,N_7992,N_7993,N_7995,N_7996,N_7997,N_7998,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8009,N_8012,N_8013,N_8014,N_8015,N_8016,N_8019,N_8020,N_8023,N_8025,N_8026,N_8028,N_8029,N_8031,N_8033,N_8035,N_8037,N_8042,N_8044,N_8045,N_8048,N_8050,N_8051,N_8052,N_8053,N_8055,N_8056,N_8059,N_8061,N_8063,N_8065,N_8066,N_8070,N_8073,N_8075,N_8076,N_8078,N_8081,N_8082,N_8083,N_8086,N_8088,N_8089,N_8090,N_8093,N_8095,N_8096,N_8097,N_8098,N_8100,N_8101,N_8102,N_8106,N_8107,N_8109,N_8110,N_8111,N_8112,N_8113,N_8115,N_8117,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8136,N_8137,N_8139,N_8140,N_8146,N_8148,N_8149,N_8151,N_8152,N_8157,N_8159,N_8161,N_8162,N_8163,N_8166,N_8169,N_8170,N_8171,N_8173,N_8174,N_8175,N_8176,N_8178,N_8179,N_8180,N_8182,N_8184,N_8186,N_8188,N_8189,N_8193,N_8194,N_8198,N_8199,N_8200,N_8202,N_8204,N_8205,N_8207,N_8209,N_8213,N_8214,N_8217,N_8218,N_8220,N_8221,N_8222,N_8225,N_8226,N_8227,N_8228,N_8230,N_8231,N_8233,N_8234,N_8235,N_8237,N_8238,N_8239,N_8244,N_8245,N_8246,N_8248,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8266,N_8267,N_8268,N_8275,N_8279,N_8282,N_8284,N_8285,N_8286,N_8287,N_8288,N_8290,N_8291,N_8292,N_8296,N_8302,N_8305,N_8307,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8319,N_8320,N_8321,N_8322,N_8324,N_8325,N_8326,N_8327,N_8329,N_8330,N_8336,N_8338,N_8339,N_8340,N_8341,N_8342,N_8344,N_8345,N_8348,N_8349,N_8350,N_8351,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8366,N_8369,N_8371,N_8372,N_8375,N_8376,N_8377,N_8380,N_8381,N_8382,N_8384,N_8385,N_8386,N_8387,N_8389,N_8390,N_8391,N_8392,N_8395,N_8396,N_8397,N_8398,N_8400,N_8402,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8414,N_8415,N_8417,N_8419,N_8420,N_8421,N_8422,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8431,N_8432,N_8434,N_8435,N_8436,N_8437,N_8441,N_8442,N_8443,N_8446,N_8447,N_8448,N_8451,N_8452,N_8455,N_8456,N_8457,N_8460,N_8463,N_8464,N_8466,N_8467,N_8468,N_8470,N_8471,N_8472,N_8474,N_8476,N_8477,N_8479,N_8480,N_8481,N_8483,N_8484,N_8485,N_8490,N_8492,N_8494,N_8495,N_8499,N_8501,N_8503,N_8504,N_8505,N_8510,N_8511,N_8512,N_8513,N_8514,N_8516,N_8517,N_8518,N_8527,N_8528,N_8530,N_8531,N_8535,N_8538,N_8540,N_8543,N_8544,N_8547,N_8549,N_8550,N_8552,N_8553,N_8561,N_8563,N_8564,N_8566,N_8568,N_8572,N_8580,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8594,N_8596,N_8597,N_8598,N_8600,N_8602,N_8603,N_8604,N_8608,N_8609,N_8610,N_8611,N_8614,N_8616,N_8618,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8630,N_8633,N_8635,N_8636,N_8637,N_8639,N_8640,N_8643,N_8647,N_8648,N_8649,N_8653,N_8655,N_8657,N_8658,N_8662,N_8663,N_8664,N_8667,N_8669,N_8670,N_8673,N_8676,N_8677,N_8680,N_8681,N_8684,N_8686,N_8687,N_8690,N_8691,N_8692,N_8695,N_8696,N_8697,N_8699,N_8700,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8714,N_8715,N_8720,N_8721,N_8722,N_8724,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8741,N_8743,N_8744,N_8745,N_8748,N_8750,N_8754,N_8755,N_8757,N_8759,N_8761,N_8762,N_8763,N_8764,N_8767,N_8768,N_8769,N_8771,N_8773,N_8774,N_8776,N_8778,N_8779,N_8780,N_8782,N_8783,N_8784,N_8787,N_8788,N_8789,N_8791,N_8792,N_8794,N_8795,N_8799,N_8801,N_8802,N_8803,N_8804,N_8805,N_8808,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8818,N_8819,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8831,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8843,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8860,N_8861,N_8862,N_8863,N_8864,N_8866,N_8867,N_8868,N_8869,N_8870,N_8872,N_8873,N_8874,N_8877,N_8878,N_8879,N_8881,N_8883,N_8884,N_8886,N_8888,N_8890,N_8891,N_8892,N_8893,N_8896,N_8897,N_8900,N_8902,N_8906,N_8907,N_8909,N_8910,N_8911,N_8913,N_8914,N_8915,N_8916,N_8919,N_8920,N_8921,N_8922,N_8923,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8934,N_8935,N_8936,N_8937,N_8938,N_8942,N_8943,N_8945,N_8946,N_8947,N_8949,N_8950,N_8951,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8966,N_8968,N_8970,N_8971,N_8972,N_8973,N_8975,N_8979,N_8981,N_8982,N_8987,N_8990,N_8992,N_8995,N_8996,N_8997,N_8998,N_9000,N_9002,N_9003,N_9007,N_9010,N_9012,N_9013,N_9014,N_9015,N_9020,N_9022,N_9023,N_9024,N_9026,N_9028,N_9029,N_9031,N_9033,N_9034,N_9036,N_9037,N_9038,N_9039,N_9041,N_9042,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9052,N_9053,N_9056,N_9059,N_9066,N_9067,N_9068,N_9071,N_9075,N_9076,N_9078,N_9080,N_9083,N_9086,N_9087,N_9088,N_9092,N_9093,N_9094,N_9096,N_9098,N_9102,N_9103,N_9104,N_9105,N_9107,N_9108,N_9110,N_9111,N_9112,N_9114,N_9116,N_9117,N_9118,N_9119,N_9120,N_9122,N_9124,N_9125,N_9126,N_9127,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9137,N_9138,N_9139,N_9140,N_9142,N_9143,N_9145,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9155,N_9156,N_9157,N_9159,N_9160,N_9161,N_9162,N_9165,N_9166,N_9169,N_9171,N_9172,N_9173,N_9174,N_9177,N_9179,N_9180,N_9184,N_9185,N_9186,N_9187,N_9189,N_9192,N_9193,N_9194,N_9195,N_9197,N_9202,N_9203,N_9204,N_9207,N_9209,N_9211,N_9214,N_9216,N_9217,N_9218,N_9219,N_9220,N_9225,N_9229,N_9231,N_9237,N_9238,N_9239,N_9241,N_9245,N_9247,N_9248,N_9249,N_9251,N_9257,N_9261,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9278,N_9280,N_9281,N_9282,N_9285,N_9288,N_9289,N_9292,N_9294,N_9295,N_9296,N_9298,N_9300,N_9301,N_9303,N_9305,N_9306,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9328,N_9329,N_9331,N_9332,N_9333,N_9334,N_9336,N_9338,N_9339,N_9342,N_9343,N_9346,N_9348,N_9352,N_9354,N_9355,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9368,N_9369,N_9371,N_9372,N_9373,N_9374,N_9376,N_9379,N_9380,N_9381,N_9382,N_9383,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9397,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9406,N_9409,N_9410,N_9412,N_9414,N_9416,N_9419,N_9422,N_9425,N_9426,N_9427,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9437,N_9439,N_9440,N_9441,N_9442,N_9444,N_9446,N_9447,N_9449,N_9450,N_9451,N_9452,N_9454,N_9455,N_9458,N_9459,N_9460,N_9461,N_9464,N_9465,N_9467,N_9469,N_9470,N_9471,N_9473,N_9475,N_9476,N_9478,N_9480,N_9482,N_9483,N_9485,N_9486,N_9488,N_9494,N_9495,N_9496,N_9500,N_9502,N_9503,N_9506,N_9507,N_9509,N_9510,N_9513,N_9514,N_9515,N_9516,N_9517,N_9519,N_9520,N_9521,N_9523,N_9525,N_9526,N_9530,N_9531,N_9532,N_9533,N_9534,N_9536,N_9537,N_9538,N_9539,N_9540,N_9542,N_9543,N_9544,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9555,N_9556,N_9557,N_9558,N_9559,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9581,N_9582,N_9583,N_9586,N_9587,N_9588,N_9589,N_9594,N_9595,N_9597,N_9598,N_9600,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9621,N_9622,N_9624,N_9625,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9634,N_9635,N_9637,N_9638,N_9639,N_9640,N_9641,N_9645,N_9647,N_9648,N_9649,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9661,N_9664,N_9665,N_9668,N_9670,N_9671,N_9672,N_9677,N_9681,N_9685,N_9686,N_9689,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9701,N_9702,N_9704,N_9705,N_9706,N_9708,N_9709,N_9713,N_9715,N_9716,N_9717,N_9719,N_9722,N_9723,N_9724,N_9727,N_9728,N_9729,N_9735,N_9736,N_9738,N_9741,N_9742,N_9746,N_9747,N_9749,N_9750,N_9752,N_9754,N_9755,N_9759,N_9760,N_9763,N_9764,N_9765,N_9767,N_9768,N_9771,N_9772,N_9774,N_9775,N_9777,N_9779,N_9780,N_9782,N_9783,N_9784,N_9785,N_9786,N_9791,N_9794,N_9795,N_9797,N_9798,N_9799,N_9800,N_9803,N_9804,N_9808,N_9809,N_9810,N_9811,N_9812,N_9814,N_9815,N_9816,N_9817,N_9820,N_9825,N_9826,N_9827,N_9828,N_9829,N_9831,N_9834,N_9836,N_9838,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9851,N_9852,N_9853,N_9854,N_9856,N_9857,N_9859,N_9861,N_9864,N_9865,N_9866,N_9869,N_9870,N_9873,N_9874,N_9877,N_9879,N_9880,N_9881,N_9882,N_9883,N_9885,N_9887,N_9888,N_9889,N_9893,N_9894,N_9895,N_9898,N_9900,N_9901,N_9903,N_9904,N_9906,N_9907,N_9908,N_9910,N_9912,N_9913,N_9915,N_9917,N_9919,N_9920,N_9921,N_9922,N_9923,N_9926,N_9929,N_9931,N_9932,N_9934,N_9935,N_9938,N_9939,N_9940,N_9942,N_9943,N_9944,N_9945,N_9946,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9960,N_9961,N_9966,N_9969,N_9970,N_9972,N_9974,N_9975,N_9976,N_9977,N_9981,N_9983,N_9984,N_9985,N_9986,N_9987,N_9991,N_9992,N_9993,N_9994,N_9996,N_9998,N_9999;
xnor U0 (N_0,In_547,In_112);
or U1 (N_1,In_167,In_451);
or U2 (N_2,In_751,In_1);
nor U3 (N_3,In_797,In_526);
nor U4 (N_4,In_268,In_453);
or U5 (N_5,In_370,In_975);
nand U6 (N_6,In_884,In_59);
nand U7 (N_7,In_179,In_645);
or U8 (N_8,In_554,In_696);
xor U9 (N_9,In_474,In_796);
nand U10 (N_10,In_262,In_338);
xor U11 (N_11,In_378,In_33);
and U12 (N_12,In_950,In_923);
nor U13 (N_13,In_424,In_106);
or U14 (N_14,In_72,In_701);
nand U15 (N_15,In_94,In_45);
nand U16 (N_16,In_164,In_443);
nor U17 (N_17,In_551,In_707);
nand U18 (N_18,In_345,In_865);
xnor U19 (N_19,In_694,In_208);
or U20 (N_20,In_716,In_736);
nand U21 (N_21,In_902,In_987);
and U22 (N_22,In_661,In_662);
and U23 (N_23,In_286,In_559);
xor U24 (N_24,In_663,In_320);
xor U25 (N_25,In_592,In_122);
nand U26 (N_26,In_698,In_416);
nor U27 (N_27,In_355,In_74);
nor U28 (N_28,In_798,In_450);
and U29 (N_29,In_905,In_613);
and U30 (N_30,In_56,In_580);
or U31 (N_31,In_408,In_172);
or U32 (N_32,In_974,In_487);
nor U33 (N_33,In_389,In_478);
nor U34 (N_34,In_337,In_692);
nor U35 (N_35,In_608,In_568);
and U36 (N_36,In_757,In_388);
or U37 (N_37,In_273,In_103);
xnor U38 (N_38,In_814,In_271);
or U39 (N_39,In_555,In_577);
and U40 (N_40,In_753,In_600);
nand U41 (N_41,In_894,In_236);
or U42 (N_42,In_898,In_848);
xnor U43 (N_43,In_965,In_540);
nand U44 (N_44,In_823,In_418);
and U45 (N_45,In_657,In_879);
or U46 (N_46,In_145,In_911);
and U47 (N_47,In_35,In_223);
nor U48 (N_48,In_260,In_705);
xor U49 (N_49,In_219,In_447);
nand U50 (N_50,In_149,In_459);
and U51 (N_51,In_855,In_252);
xnor U52 (N_52,In_25,In_926);
or U53 (N_53,In_952,In_326);
nor U54 (N_54,In_254,In_788);
or U55 (N_55,In_825,In_70);
nor U56 (N_56,In_27,In_805);
or U57 (N_57,In_88,In_976);
or U58 (N_58,In_482,In_431);
nor U59 (N_59,In_383,In_50);
nor U60 (N_60,In_312,In_517);
and U61 (N_61,In_503,In_209);
xor U62 (N_62,In_293,In_55);
and U63 (N_63,In_935,In_634);
or U64 (N_64,In_651,In_615);
nor U65 (N_65,In_372,In_405);
or U66 (N_66,In_476,In_31);
nand U67 (N_67,In_17,In_168);
or U68 (N_68,In_496,In_841);
nand U69 (N_69,In_708,In_192);
and U70 (N_70,In_81,In_834);
nor U71 (N_71,In_135,In_231);
or U72 (N_72,In_959,In_259);
nor U73 (N_73,In_175,In_358);
nand U74 (N_74,In_494,In_614);
nand U75 (N_75,In_560,In_748);
xnor U76 (N_76,In_785,In_737);
nor U77 (N_77,In_656,In_346);
xor U78 (N_78,In_318,In_774);
and U79 (N_79,In_703,In_221);
xnor U80 (N_80,In_996,In_137);
xnor U81 (N_81,In_261,In_756);
or U82 (N_82,In_816,In_321);
nand U83 (N_83,In_573,In_795);
nor U84 (N_84,In_764,In_782);
xnor U85 (N_85,In_104,In_632);
or U86 (N_86,In_586,In_4);
and U87 (N_87,In_549,In_15);
and U88 (N_88,In_497,In_384);
nand U89 (N_89,In_859,In_518);
nand U90 (N_90,In_124,In_21);
xor U91 (N_91,In_724,In_763);
or U92 (N_92,In_28,In_619);
nor U93 (N_93,In_30,In_413);
or U94 (N_94,In_427,In_151);
nor U95 (N_95,In_118,In_896);
or U96 (N_96,In_771,In_519);
xnor U97 (N_97,In_341,In_620);
and U98 (N_98,In_304,In_361);
xor U99 (N_99,In_604,In_465);
nand U100 (N_100,In_462,In_150);
nand U101 (N_101,In_759,In_166);
or U102 (N_102,In_277,In_366);
or U103 (N_103,In_817,In_516);
or U104 (N_104,In_979,In_210);
and U105 (N_105,In_811,In_942);
or U106 (N_106,In_909,In_311);
nor U107 (N_107,In_69,In_793);
nand U108 (N_108,In_181,In_198);
or U109 (N_109,In_704,In_919);
and U110 (N_110,In_875,In_300);
xor U111 (N_111,In_351,In_733);
xnor U112 (N_112,In_644,In_787);
nor U113 (N_113,In_892,In_120);
nand U114 (N_114,In_729,In_943);
nand U115 (N_115,In_316,In_769);
nand U116 (N_116,In_882,In_635);
nand U117 (N_117,In_544,In_618);
nor U118 (N_118,In_853,In_993);
nand U119 (N_119,In_468,In_3);
or U120 (N_120,In_477,In_813);
nor U121 (N_121,In_62,In_415);
xor U122 (N_122,In_359,In_65);
xnor U123 (N_123,In_131,In_486);
xnor U124 (N_124,In_889,In_189);
and U125 (N_125,In_750,In_713);
or U126 (N_126,In_801,In_781);
and U127 (N_127,In_414,In_435);
nand U128 (N_128,In_490,In_812);
and U129 (N_129,In_669,In_360);
nand U130 (N_130,In_58,In_583);
xor U131 (N_131,In_404,In_836);
or U132 (N_132,In_23,In_986);
nor U133 (N_133,In_948,In_152);
xnor U134 (N_134,In_49,In_350);
xnor U135 (N_135,In_863,In_80);
xnor U136 (N_136,In_754,In_977);
or U137 (N_137,In_832,In_876);
nand U138 (N_138,In_457,In_978);
nand U139 (N_139,In_401,In_740);
nand U140 (N_140,In_125,In_340);
nand U141 (N_141,In_44,In_274);
or U142 (N_142,In_946,In_711);
and U143 (N_143,In_446,In_157);
xnor U144 (N_144,In_130,In_772);
and U145 (N_145,In_76,In_229);
and U146 (N_146,In_406,In_913);
xnor U147 (N_147,In_387,In_883);
nor U148 (N_148,In_988,In_745);
nor U149 (N_149,In_190,In_934);
and U150 (N_150,In_289,In_224);
nand U151 (N_151,In_660,In_222);
nor U152 (N_152,In_114,In_994);
and U153 (N_153,In_347,In_242);
and U154 (N_154,In_333,In_217);
nor U155 (N_155,In_502,In_362);
xor U156 (N_156,In_365,In_225);
nand U157 (N_157,In_957,In_835);
and U158 (N_158,In_538,In_593);
xor U159 (N_159,In_524,In_680);
or U160 (N_160,In_63,In_531);
xnor U161 (N_161,In_279,In_721);
nor U162 (N_162,In_510,In_777);
nor U163 (N_163,In_275,In_546);
or U164 (N_164,In_99,In_655);
and U165 (N_165,In_310,In_438);
and U166 (N_166,In_639,In_958);
xor U167 (N_167,In_200,In_390);
and U168 (N_168,In_379,In_43);
or U169 (N_169,In_471,In_970);
nor U170 (N_170,In_68,In_990);
nand U171 (N_171,In_671,In_565);
nand U172 (N_172,In_407,In_216);
xor U173 (N_173,In_392,In_897);
xor U174 (N_174,In_205,In_283);
xnor U175 (N_175,In_837,In_397);
or U176 (N_176,In_563,In_709);
nand U177 (N_177,In_344,In_850);
and U178 (N_178,In_215,In_421);
xnor U179 (N_179,In_877,In_686);
nor U180 (N_180,In_849,In_95);
xor U181 (N_181,In_203,In_770);
and U182 (N_182,In_910,In_691);
nor U183 (N_183,In_47,In_238);
nor U184 (N_184,In_758,In_423);
or U185 (N_185,In_108,In_985);
and U186 (N_186,In_339,In_206);
and U187 (N_187,In_308,In_628);
nor U188 (N_188,In_891,In_927);
and U189 (N_189,In_609,In_322);
nand U190 (N_190,In_687,In_410);
xnor U191 (N_191,In_434,In_802);
nand U192 (N_192,In_980,In_40);
or U193 (N_193,In_429,In_41);
nand U194 (N_194,In_539,In_412);
or U195 (N_195,In_285,In_963);
nor U196 (N_196,In_741,In_845);
or U197 (N_197,In_685,In_621);
and U198 (N_198,In_810,In_141);
or U199 (N_199,In_684,In_469);
nand U200 (N_200,In_806,In_601);
nor U201 (N_201,In_827,In_643);
or U202 (N_202,In_140,In_689);
and U203 (N_203,In_162,In_36);
or U204 (N_204,In_336,In_473);
and U205 (N_205,In_679,In_101);
or U206 (N_206,In_562,In_386);
nor U207 (N_207,In_314,In_96);
xnor U208 (N_208,In_278,In_235);
xor U209 (N_209,In_641,In_523);
or U210 (N_210,In_944,In_234);
nor U211 (N_211,In_245,In_638);
nor U212 (N_212,In_218,In_204);
or U213 (N_213,In_485,In_54);
and U214 (N_214,In_38,In_323);
nor U215 (N_215,In_342,In_940);
and U216 (N_216,In_301,In_881);
xor U217 (N_217,In_255,In_739);
xor U218 (N_218,In_852,In_16);
and U219 (N_219,In_989,In_822);
and U220 (N_220,In_553,In_437);
nand U221 (N_221,In_887,In_624);
and U222 (N_222,In_981,In_281);
xor U223 (N_223,In_195,In_177);
and U224 (N_224,In_594,In_633);
nor U225 (N_225,In_706,In_269);
or U226 (N_226,In_481,In_442);
nand U227 (N_227,In_2,In_374);
nor U228 (N_228,In_385,In_265);
nor U229 (N_229,In_847,In_839);
nand U230 (N_230,In_995,In_129);
nand U231 (N_231,In_143,In_931);
and U232 (N_232,In_182,In_629);
nand U233 (N_233,In_287,In_393);
xor U234 (N_234,In_332,In_677);
and U235 (N_235,In_147,In_452);
and U236 (N_236,In_417,In_295);
nand U237 (N_237,In_697,In_664);
nor U238 (N_238,In_612,In_299);
and U239 (N_239,In_918,In_34);
nand U240 (N_240,In_610,In_906);
and U241 (N_241,In_296,In_991);
nor U242 (N_242,In_676,In_302);
or U243 (N_243,In_566,In_78);
or U244 (N_244,In_420,In_776);
nor U245 (N_245,In_317,In_541);
xor U246 (N_246,In_57,In_860);
nand U247 (N_247,In_922,In_77);
or U248 (N_248,In_5,In_331);
nand U249 (N_249,In_693,In_640);
or U250 (N_250,In_213,In_305);
nand U251 (N_251,In_82,In_495);
or U252 (N_252,In_232,In_515);
nand U253 (N_253,In_498,In_91);
or U254 (N_254,In_804,In_6);
or U255 (N_255,In_702,In_840);
or U256 (N_256,In_212,In_960);
and U257 (N_257,In_0,In_504);
nor U258 (N_258,In_144,In_844);
and U259 (N_259,In_792,In_874);
nand U260 (N_260,In_900,In_667);
or U261 (N_261,In_303,In_492);
or U262 (N_262,In_20,In_880);
nor U263 (N_263,In_869,In_688);
xor U264 (N_264,In_542,In_507);
and U265 (N_265,In_917,In_857);
or U266 (N_266,In_622,In_732);
nor U267 (N_267,In_324,In_760);
nor U268 (N_268,In_357,In_7);
xor U269 (N_269,In_163,In_712);
or U270 (N_270,In_982,In_132);
and U271 (N_271,In_574,In_521);
or U272 (N_272,In_11,In_98);
nor U273 (N_273,In_747,In_42);
and U274 (N_274,In_230,In_647);
or U275 (N_275,In_949,In_363);
nand U276 (N_276,In_867,In_66);
xor U277 (N_277,In_587,In_250);
and U278 (N_278,In_327,In_211);
nor U279 (N_279,In_961,In_779);
xor U280 (N_280,In_846,In_522);
nor U281 (N_281,In_461,In_530);
nor U282 (N_282,In_199,In_155);
nor U283 (N_283,In_470,In_878);
nand U284 (N_284,In_625,In_557);
nor U285 (N_285,In_734,In_354);
nor U286 (N_286,In_176,In_695);
nor U287 (N_287,In_642,In_945);
nand U288 (N_288,In_121,In_315);
and U289 (N_289,In_650,In_403);
xor U290 (N_290,In_10,In_356);
and U291 (N_291,In_353,In_956);
nor U292 (N_292,In_514,In_89);
or U293 (N_293,In_821,In_570);
and U294 (N_294,In_173,In_824);
nor U295 (N_295,In_46,In_202);
xnor U296 (N_296,In_738,In_616);
nand U297 (N_297,In_529,In_93);
and U298 (N_298,In_105,In_445);
and U299 (N_299,In_9,In_267);
nor U300 (N_300,In_18,In_425);
nand U301 (N_301,In_8,In_999);
and U302 (N_302,In_138,In_449);
and U303 (N_303,In_29,In_433);
nand U304 (N_304,In_228,In_527);
xor U305 (N_305,In_842,In_765);
and U306 (N_306,In_491,In_607);
nand U307 (N_307,In_588,In_307);
nand U308 (N_308,In_895,In_75);
or U309 (N_309,In_84,In_107);
or U310 (N_310,In_264,In_746);
xor U311 (N_311,In_675,In_964);
or U312 (N_312,In_24,In_272);
nand U313 (N_313,In_391,In_537);
xor U314 (N_314,In_501,In_325);
xnor U315 (N_315,In_297,In_456);
xnor U316 (N_316,In_672,In_731);
nor U317 (N_317,In_159,In_561);
and U318 (N_318,In_398,In_444);
and U319 (N_319,In_833,In_901);
or U320 (N_320,In_862,In_794);
and U321 (N_321,In_637,In_253);
nand U322 (N_322,In_51,In_558);
or U323 (N_323,In_489,In_146);
and U324 (N_324,In_903,In_484);
and U325 (N_325,In_668,In_371);
nor U326 (N_326,In_678,In_448);
or U327 (N_327,In_119,In_730);
or U328 (N_328,In_64,In_111);
xnor U329 (N_329,In_419,In_670);
and U330 (N_330,In_767,In_455);
xnor U331 (N_331,In_270,In_611);
nor U332 (N_332,In_207,In_480);
nor U333 (N_333,In_174,In_467);
nor U334 (N_334,In_117,In_727);
or U335 (N_335,In_893,In_382);
nor U336 (N_336,In_441,In_997);
xnor U337 (N_337,In_178,In_907);
and U338 (N_338,In_890,In_761);
nor U339 (N_339,In_921,In_630);
or U340 (N_340,In_830,In_520);
nor U341 (N_341,In_735,In_888);
or U342 (N_342,In_631,In_483);
nor U343 (N_343,In_400,In_838);
nand U344 (N_344,In_717,In_169);
nor U345 (N_345,In_930,In_590);
xnor U346 (N_346,In_116,In_87);
and U347 (N_347,In_13,In_636);
xnor U348 (N_348,In_807,In_962);
and U349 (N_349,In_505,In_886);
or U350 (N_350,In_723,In_605);
and U351 (N_351,In_575,In_872);
nor U352 (N_352,In_201,In_532);
and U353 (N_353,In_376,In_153);
nor U354 (N_354,In_422,In_67);
or U355 (N_355,In_591,In_368);
and U356 (N_356,In_440,In_599);
and U357 (N_357,In_369,In_248);
nand U358 (N_358,In_596,In_428);
nand U359 (N_359,In_185,In_773);
nand U360 (N_360,In_955,In_920);
nor U361 (N_361,In_809,In_623);
or U362 (N_362,In_556,In_196);
nor U363 (N_363,In_819,In_464);
or U364 (N_364,In_381,In_873);
nand U365 (N_365,In_720,In_330);
and U366 (N_366,In_743,In_983);
or U367 (N_367,In_184,In_61);
nor U368 (N_368,In_969,In_187);
and U369 (N_369,In_183,In_744);
xor U370 (N_370,In_899,In_939);
nand U371 (N_371,In_992,In_439);
nor U372 (N_372,In_60,In_953);
nor U373 (N_373,In_924,In_193);
or U374 (N_374,In_180,In_512);
or U375 (N_375,In_597,In_722);
or U376 (N_376,In_430,In_399);
or U377 (N_377,In_161,In_752);
xor U378 (N_378,In_276,In_598);
and U379 (N_379,In_170,In_571);
nor U380 (N_380,In_53,In_227);
xnor U381 (N_381,In_142,In_375);
or U382 (N_382,In_954,In_197);
nor U383 (N_383,In_941,In_778);
and U384 (N_384,In_719,In_742);
nor U385 (N_385,In_683,In_126);
xnor U386 (N_386,In_348,In_460);
xor U387 (N_387,In_97,In_584);
or U388 (N_388,In_432,In_247);
or U389 (N_389,In_866,In_528);
xor U390 (N_390,In_102,In_938);
nand U391 (N_391,In_606,In_912);
nor U392 (N_392,In_352,In_755);
and U393 (N_393,In_851,In_682);
xnor U394 (N_394,In_39,In_659);
or U395 (N_395,In_789,In_309);
nand U396 (N_396,In_513,In_52);
nor U397 (N_397,In_90,In_715);
nand U398 (N_398,In_240,In_475);
xnor U399 (N_399,In_578,In_158);
or U400 (N_400,In_665,In_349);
nor U401 (N_401,In_256,In_402);
or U402 (N_402,In_454,In_826);
nor U403 (N_403,In_288,In_820);
xnor U404 (N_404,In_506,In_576);
xor U405 (N_405,In_831,In_829);
and U406 (N_406,In_466,In_329);
and U407 (N_407,In_127,In_725);
and U408 (N_408,In_110,In_582);
nand U409 (N_409,In_914,In_726);
xor U410 (N_410,In_666,In_552);
xor U411 (N_411,In_649,In_548);
xor U412 (N_412,In_535,In_967);
nand U413 (N_413,In_718,In_92);
nand U414 (N_414,In_728,In_856);
and U415 (N_415,In_626,In_12);
or U416 (N_416,In_762,In_808);
xnor U417 (N_417,In_569,In_479);
nand U418 (N_418,In_783,In_377);
nand U419 (N_419,In_343,In_589);
nand U420 (N_420,In_904,In_239);
nor U421 (N_421,In_710,In_280);
and U422 (N_422,In_291,In_328);
nor U423 (N_423,In_803,In_188);
and U424 (N_424,In_937,In_115);
and U425 (N_425,In_160,In_436);
or U426 (N_426,In_648,In_395);
nand U427 (N_427,In_700,In_257);
and U428 (N_428,In_998,In_973);
xnor U429 (N_429,In_171,In_928);
xnor U430 (N_430,In_37,In_673);
xor U431 (N_431,In_32,In_861);
and U432 (N_432,In_916,In_463);
nor U433 (N_433,In_780,In_885);
and U434 (N_434,In_864,In_251);
and U435 (N_435,In_100,In_191);
and U436 (N_436,In_133,In_972);
xor U437 (N_437,In_19,In_306);
and U438 (N_438,In_85,In_654);
xor U439 (N_439,In_749,In_83);
or U440 (N_440,In_699,In_411);
nand U441 (N_441,In_595,In_367);
nand U442 (N_442,In_653,In_714);
nor U443 (N_443,In_843,In_237);
nor U444 (N_444,In_543,In_136);
nor U445 (N_445,In_123,In_334);
nor U446 (N_446,In_984,In_373);
xor U447 (N_447,In_22,In_244);
nor U448 (N_448,In_165,In_775);
and U449 (N_449,In_766,In_791);
and U450 (N_450,In_627,In_603);
nand U451 (N_451,In_364,In_525);
xor U452 (N_452,In_585,In_500);
nor U453 (N_453,In_932,In_858);
nor U454 (N_454,In_14,In_263);
nand U455 (N_455,In_292,In_550);
xnor U456 (N_456,In_249,In_214);
and U457 (N_457,In_380,In_396);
or U458 (N_458,In_233,In_488);
nor U459 (N_459,In_545,In_567);
nor U460 (N_460,In_186,In_971);
xnor U461 (N_461,In_915,In_674);
nor U462 (N_462,In_109,In_226);
nor U463 (N_463,In_966,In_243);
and U464 (N_464,In_784,In_394);
nand U465 (N_465,In_426,In_790);
and U466 (N_466,In_48,In_951);
nor U467 (N_467,In_246,In_908);
and U468 (N_468,In_786,In_868);
and U469 (N_469,In_282,In_508);
nor U470 (N_470,In_290,In_536);
and U471 (N_471,In_26,In_579);
and U472 (N_472,In_968,In_113);
xor U473 (N_473,In_148,In_870);
xnor U474 (N_474,In_134,In_499);
or U475 (N_475,In_800,In_313);
and U476 (N_476,In_818,In_258);
nand U477 (N_477,In_71,In_564);
or U478 (N_478,In_319,In_572);
nand U479 (N_479,In_294,In_690);
or U480 (N_480,In_828,In_936);
or U481 (N_481,In_86,In_509);
nor U482 (N_482,In_581,In_241);
xnor U483 (N_483,In_511,In_658);
or U484 (N_484,In_947,In_156);
or U485 (N_485,In_933,In_194);
or U486 (N_486,In_458,In_128);
or U487 (N_487,In_602,In_493);
xor U488 (N_488,In_854,In_154);
nand U489 (N_489,In_652,In_73);
or U490 (N_490,In_284,In_79);
or U491 (N_491,In_220,In_139);
or U492 (N_492,In_929,In_298);
nor U493 (N_493,In_617,In_409);
xnor U494 (N_494,In_335,In_472);
nand U495 (N_495,In_646,In_681);
or U496 (N_496,In_815,In_799);
nand U497 (N_497,In_533,In_768);
or U498 (N_498,In_925,In_266);
nand U499 (N_499,In_871,In_534);
or U500 (N_500,In_123,In_172);
nand U501 (N_501,In_968,In_139);
nor U502 (N_502,In_309,In_569);
nor U503 (N_503,In_908,In_258);
xnor U504 (N_504,In_437,In_663);
or U505 (N_505,In_272,In_664);
or U506 (N_506,In_156,In_470);
nor U507 (N_507,In_688,In_63);
nor U508 (N_508,In_59,In_872);
or U509 (N_509,In_579,In_712);
and U510 (N_510,In_750,In_719);
nand U511 (N_511,In_849,In_493);
nor U512 (N_512,In_833,In_968);
or U513 (N_513,In_569,In_440);
or U514 (N_514,In_445,In_381);
nor U515 (N_515,In_825,In_415);
nor U516 (N_516,In_699,In_111);
and U517 (N_517,In_943,In_87);
or U518 (N_518,In_902,In_562);
nor U519 (N_519,In_423,In_855);
nor U520 (N_520,In_129,In_866);
xnor U521 (N_521,In_465,In_194);
nand U522 (N_522,In_718,In_301);
xnor U523 (N_523,In_920,In_310);
nand U524 (N_524,In_56,In_680);
and U525 (N_525,In_144,In_958);
nor U526 (N_526,In_41,In_674);
nand U527 (N_527,In_72,In_792);
nand U528 (N_528,In_436,In_628);
or U529 (N_529,In_68,In_50);
and U530 (N_530,In_703,In_651);
xnor U531 (N_531,In_529,In_83);
nand U532 (N_532,In_222,In_34);
nand U533 (N_533,In_706,In_264);
nand U534 (N_534,In_938,In_215);
nor U535 (N_535,In_133,In_648);
nor U536 (N_536,In_720,In_498);
nand U537 (N_537,In_503,In_514);
nand U538 (N_538,In_481,In_395);
nor U539 (N_539,In_678,In_129);
nor U540 (N_540,In_378,In_225);
and U541 (N_541,In_740,In_222);
or U542 (N_542,In_232,In_968);
nor U543 (N_543,In_739,In_479);
and U544 (N_544,In_310,In_315);
xor U545 (N_545,In_613,In_190);
and U546 (N_546,In_964,In_860);
nor U547 (N_547,In_900,In_717);
xnor U548 (N_548,In_999,In_145);
xnor U549 (N_549,In_698,In_351);
xnor U550 (N_550,In_495,In_680);
xor U551 (N_551,In_651,In_351);
nor U552 (N_552,In_362,In_963);
nor U553 (N_553,In_58,In_355);
or U554 (N_554,In_46,In_760);
nor U555 (N_555,In_355,In_534);
or U556 (N_556,In_613,In_400);
xnor U557 (N_557,In_135,In_38);
nor U558 (N_558,In_830,In_996);
or U559 (N_559,In_350,In_256);
xor U560 (N_560,In_351,In_631);
nand U561 (N_561,In_497,In_871);
xnor U562 (N_562,In_711,In_667);
xnor U563 (N_563,In_559,In_661);
nor U564 (N_564,In_820,In_691);
nand U565 (N_565,In_339,In_990);
xnor U566 (N_566,In_984,In_970);
xor U567 (N_567,In_305,In_827);
nand U568 (N_568,In_284,In_886);
or U569 (N_569,In_978,In_887);
and U570 (N_570,In_448,In_196);
nand U571 (N_571,In_803,In_81);
xor U572 (N_572,In_238,In_723);
nor U573 (N_573,In_235,In_128);
or U574 (N_574,In_48,In_570);
nor U575 (N_575,In_397,In_764);
nor U576 (N_576,In_318,In_974);
and U577 (N_577,In_561,In_42);
nor U578 (N_578,In_619,In_398);
or U579 (N_579,In_41,In_212);
or U580 (N_580,In_255,In_887);
nand U581 (N_581,In_466,In_219);
and U582 (N_582,In_925,In_333);
and U583 (N_583,In_368,In_283);
xnor U584 (N_584,In_717,In_155);
and U585 (N_585,In_648,In_95);
and U586 (N_586,In_556,In_33);
nor U587 (N_587,In_107,In_263);
xor U588 (N_588,In_961,In_673);
nand U589 (N_589,In_421,In_386);
nand U590 (N_590,In_77,In_253);
or U591 (N_591,In_558,In_19);
nand U592 (N_592,In_904,In_905);
or U593 (N_593,In_737,In_382);
or U594 (N_594,In_375,In_835);
nor U595 (N_595,In_661,In_506);
nor U596 (N_596,In_536,In_451);
nand U597 (N_597,In_66,In_633);
nor U598 (N_598,In_887,In_357);
and U599 (N_599,In_598,In_830);
nor U600 (N_600,In_922,In_289);
or U601 (N_601,In_492,In_207);
or U602 (N_602,In_165,In_890);
or U603 (N_603,In_691,In_985);
xor U604 (N_604,In_389,In_196);
nand U605 (N_605,In_709,In_168);
nand U606 (N_606,In_740,In_839);
nor U607 (N_607,In_289,In_971);
and U608 (N_608,In_827,In_149);
and U609 (N_609,In_642,In_14);
nand U610 (N_610,In_846,In_204);
nand U611 (N_611,In_542,In_772);
or U612 (N_612,In_879,In_549);
and U613 (N_613,In_800,In_527);
and U614 (N_614,In_619,In_278);
and U615 (N_615,In_18,In_831);
or U616 (N_616,In_985,In_959);
nand U617 (N_617,In_254,In_228);
or U618 (N_618,In_358,In_584);
nor U619 (N_619,In_788,In_268);
or U620 (N_620,In_977,In_713);
xnor U621 (N_621,In_526,In_738);
or U622 (N_622,In_158,In_410);
nor U623 (N_623,In_148,In_701);
or U624 (N_624,In_560,In_724);
nand U625 (N_625,In_629,In_924);
nor U626 (N_626,In_928,In_846);
xnor U627 (N_627,In_698,In_126);
or U628 (N_628,In_977,In_4);
xnor U629 (N_629,In_617,In_849);
nor U630 (N_630,In_498,In_185);
or U631 (N_631,In_452,In_536);
nand U632 (N_632,In_363,In_701);
or U633 (N_633,In_341,In_235);
xnor U634 (N_634,In_160,In_943);
xor U635 (N_635,In_881,In_233);
xnor U636 (N_636,In_405,In_618);
nand U637 (N_637,In_234,In_780);
nand U638 (N_638,In_877,In_44);
and U639 (N_639,In_198,In_189);
and U640 (N_640,In_14,In_527);
or U641 (N_641,In_16,In_915);
or U642 (N_642,In_464,In_512);
nor U643 (N_643,In_370,In_447);
and U644 (N_644,In_56,In_214);
nor U645 (N_645,In_9,In_633);
nor U646 (N_646,In_774,In_646);
xor U647 (N_647,In_163,In_197);
and U648 (N_648,In_861,In_411);
xnor U649 (N_649,In_430,In_388);
nor U650 (N_650,In_70,In_664);
and U651 (N_651,In_729,In_318);
nor U652 (N_652,In_195,In_810);
nand U653 (N_653,In_513,In_538);
or U654 (N_654,In_188,In_216);
xor U655 (N_655,In_708,In_793);
and U656 (N_656,In_142,In_755);
or U657 (N_657,In_193,In_279);
or U658 (N_658,In_259,In_924);
xnor U659 (N_659,In_256,In_223);
nand U660 (N_660,In_737,In_283);
nand U661 (N_661,In_218,In_235);
nand U662 (N_662,In_386,In_516);
and U663 (N_663,In_59,In_339);
and U664 (N_664,In_750,In_15);
xnor U665 (N_665,In_246,In_227);
nand U666 (N_666,In_184,In_452);
nand U667 (N_667,In_607,In_721);
nand U668 (N_668,In_465,In_522);
nor U669 (N_669,In_595,In_132);
or U670 (N_670,In_749,In_509);
or U671 (N_671,In_295,In_556);
nand U672 (N_672,In_442,In_101);
xor U673 (N_673,In_705,In_958);
and U674 (N_674,In_865,In_600);
xor U675 (N_675,In_298,In_353);
nor U676 (N_676,In_671,In_801);
nor U677 (N_677,In_20,In_250);
nand U678 (N_678,In_374,In_281);
nand U679 (N_679,In_403,In_800);
nor U680 (N_680,In_39,In_972);
and U681 (N_681,In_661,In_80);
or U682 (N_682,In_735,In_436);
nand U683 (N_683,In_45,In_249);
and U684 (N_684,In_291,In_90);
and U685 (N_685,In_448,In_80);
and U686 (N_686,In_339,In_928);
or U687 (N_687,In_337,In_474);
xnor U688 (N_688,In_28,In_511);
or U689 (N_689,In_48,In_290);
or U690 (N_690,In_366,In_292);
nor U691 (N_691,In_201,In_874);
and U692 (N_692,In_168,In_724);
or U693 (N_693,In_895,In_804);
xor U694 (N_694,In_485,In_119);
xor U695 (N_695,In_380,In_100);
and U696 (N_696,In_562,In_306);
and U697 (N_697,In_490,In_135);
xor U698 (N_698,In_241,In_211);
nor U699 (N_699,In_374,In_316);
xor U700 (N_700,In_859,In_41);
and U701 (N_701,In_857,In_451);
nor U702 (N_702,In_865,In_240);
nor U703 (N_703,In_95,In_397);
nand U704 (N_704,In_90,In_428);
nor U705 (N_705,In_275,In_62);
and U706 (N_706,In_242,In_612);
or U707 (N_707,In_522,In_371);
or U708 (N_708,In_167,In_368);
nand U709 (N_709,In_870,In_537);
nand U710 (N_710,In_395,In_701);
nand U711 (N_711,In_961,In_487);
and U712 (N_712,In_589,In_59);
nor U713 (N_713,In_712,In_529);
and U714 (N_714,In_600,In_611);
nor U715 (N_715,In_970,In_846);
nand U716 (N_716,In_0,In_592);
nand U717 (N_717,In_883,In_47);
xor U718 (N_718,In_129,In_632);
nor U719 (N_719,In_314,In_650);
or U720 (N_720,In_146,In_926);
or U721 (N_721,In_73,In_326);
nor U722 (N_722,In_644,In_816);
xor U723 (N_723,In_682,In_366);
and U724 (N_724,In_126,In_598);
xnor U725 (N_725,In_512,In_212);
or U726 (N_726,In_195,In_706);
or U727 (N_727,In_374,In_131);
and U728 (N_728,In_325,In_644);
nand U729 (N_729,In_54,In_888);
xnor U730 (N_730,In_250,In_202);
xnor U731 (N_731,In_152,In_176);
nor U732 (N_732,In_301,In_159);
nand U733 (N_733,In_476,In_676);
or U734 (N_734,In_662,In_876);
xnor U735 (N_735,In_311,In_177);
nand U736 (N_736,In_458,In_165);
nand U737 (N_737,In_172,In_542);
and U738 (N_738,In_679,In_986);
nor U739 (N_739,In_15,In_670);
and U740 (N_740,In_208,In_388);
or U741 (N_741,In_891,In_428);
nor U742 (N_742,In_895,In_145);
nand U743 (N_743,In_207,In_795);
nor U744 (N_744,In_519,In_858);
and U745 (N_745,In_819,In_301);
and U746 (N_746,In_77,In_985);
and U747 (N_747,In_907,In_236);
nor U748 (N_748,In_825,In_244);
nand U749 (N_749,In_906,In_79);
and U750 (N_750,In_616,In_389);
nor U751 (N_751,In_91,In_624);
or U752 (N_752,In_837,In_5);
or U753 (N_753,In_710,In_698);
xor U754 (N_754,In_571,In_981);
and U755 (N_755,In_857,In_23);
xnor U756 (N_756,In_176,In_343);
xor U757 (N_757,In_609,In_923);
xor U758 (N_758,In_577,In_621);
or U759 (N_759,In_427,In_584);
and U760 (N_760,In_877,In_510);
and U761 (N_761,In_944,In_626);
nand U762 (N_762,In_495,In_523);
and U763 (N_763,In_100,In_446);
nor U764 (N_764,In_900,In_151);
xor U765 (N_765,In_541,In_370);
and U766 (N_766,In_156,In_481);
nand U767 (N_767,In_382,In_500);
and U768 (N_768,In_29,In_494);
nand U769 (N_769,In_35,In_287);
xor U770 (N_770,In_329,In_42);
nor U771 (N_771,In_966,In_134);
and U772 (N_772,In_509,In_260);
or U773 (N_773,In_259,In_991);
or U774 (N_774,In_528,In_936);
nand U775 (N_775,In_684,In_644);
xnor U776 (N_776,In_614,In_30);
xnor U777 (N_777,In_967,In_21);
nand U778 (N_778,In_613,In_43);
or U779 (N_779,In_122,In_861);
or U780 (N_780,In_106,In_84);
or U781 (N_781,In_451,In_684);
nor U782 (N_782,In_711,In_575);
nand U783 (N_783,In_760,In_260);
or U784 (N_784,In_979,In_681);
xnor U785 (N_785,In_383,In_365);
nand U786 (N_786,In_20,In_297);
xor U787 (N_787,In_284,In_719);
nor U788 (N_788,In_266,In_893);
and U789 (N_789,In_469,In_706);
and U790 (N_790,In_207,In_639);
or U791 (N_791,In_491,In_373);
xnor U792 (N_792,In_642,In_463);
and U793 (N_793,In_250,In_249);
and U794 (N_794,In_904,In_695);
or U795 (N_795,In_892,In_200);
xnor U796 (N_796,In_552,In_499);
nand U797 (N_797,In_28,In_17);
or U798 (N_798,In_441,In_847);
nor U799 (N_799,In_632,In_332);
nand U800 (N_800,In_805,In_598);
nor U801 (N_801,In_567,In_577);
nand U802 (N_802,In_313,In_59);
nand U803 (N_803,In_614,In_340);
nand U804 (N_804,In_641,In_912);
xor U805 (N_805,In_280,In_411);
xnor U806 (N_806,In_548,In_38);
nand U807 (N_807,In_454,In_718);
nand U808 (N_808,In_755,In_665);
nand U809 (N_809,In_463,In_886);
or U810 (N_810,In_894,In_664);
nor U811 (N_811,In_440,In_268);
xor U812 (N_812,In_487,In_779);
or U813 (N_813,In_778,In_36);
nand U814 (N_814,In_246,In_894);
and U815 (N_815,In_671,In_433);
nand U816 (N_816,In_961,In_688);
and U817 (N_817,In_422,In_947);
or U818 (N_818,In_246,In_740);
xor U819 (N_819,In_437,In_984);
and U820 (N_820,In_168,In_390);
nand U821 (N_821,In_112,In_537);
nor U822 (N_822,In_488,In_974);
and U823 (N_823,In_683,In_213);
and U824 (N_824,In_668,In_616);
xor U825 (N_825,In_56,In_952);
xnor U826 (N_826,In_348,In_64);
and U827 (N_827,In_702,In_10);
xnor U828 (N_828,In_77,In_355);
xnor U829 (N_829,In_41,In_563);
and U830 (N_830,In_87,In_762);
or U831 (N_831,In_202,In_740);
nand U832 (N_832,In_408,In_852);
and U833 (N_833,In_949,In_375);
and U834 (N_834,In_241,In_334);
or U835 (N_835,In_744,In_480);
nand U836 (N_836,In_106,In_440);
nor U837 (N_837,In_982,In_978);
or U838 (N_838,In_296,In_552);
and U839 (N_839,In_445,In_60);
nor U840 (N_840,In_466,In_943);
nor U841 (N_841,In_158,In_433);
nand U842 (N_842,In_171,In_61);
or U843 (N_843,In_253,In_818);
xnor U844 (N_844,In_433,In_81);
nand U845 (N_845,In_770,In_882);
nand U846 (N_846,In_26,In_358);
or U847 (N_847,In_970,In_279);
nand U848 (N_848,In_807,In_402);
xor U849 (N_849,In_311,In_42);
nor U850 (N_850,In_677,In_550);
xnor U851 (N_851,In_316,In_690);
xnor U852 (N_852,In_872,In_723);
nor U853 (N_853,In_941,In_649);
or U854 (N_854,In_827,In_347);
or U855 (N_855,In_733,In_988);
nand U856 (N_856,In_300,In_155);
nand U857 (N_857,In_909,In_748);
or U858 (N_858,In_874,In_942);
or U859 (N_859,In_667,In_705);
xnor U860 (N_860,In_9,In_173);
nand U861 (N_861,In_218,In_684);
and U862 (N_862,In_131,In_648);
nor U863 (N_863,In_435,In_979);
nor U864 (N_864,In_955,In_428);
nand U865 (N_865,In_570,In_276);
nor U866 (N_866,In_261,In_260);
nand U867 (N_867,In_436,In_273);
nor U868 (N_868,In_376,In_388);
xor U869 (N_869,In_648,In_399);
nor U870 (N_870,In_739,In_709);
xnor U871 (N_871,In_357,In_84);
and U872 (N_872,In_348,In_19);
and U873 (N_873,In_326,In_774);
xnor U874 (N_874,In_106,In_645);
nand U875 (N_875,In_638,In_178);
and U876 (N_876,In_205,In_774);
or U877 (N_877,In_420,In_932);
or U878 (N_878,In_755,In_424);
nor U879 (N_879,In_352,In_31);
and U880 (N_880,In_102,In_991);
nor U881 (N_881,In_474,In_641);
and U882 (N_882,In_324,In_798);
or U883 (N_883,In_531,In_535);
xor U884 (N_884,In_281,In_476);
nand U885 (N_885,In_799,In_788);
nor U886 (N_886,In_654,In_249);
and U887 (N_887,In_858,In_428);
and U888 (N_888,In_19,In_640);
or U889 (N_889,In_267,In_952);
nand U890 (N_890,In_156,In_345);
or U891 (N_891,In_812,In_363);
and U892 (N_892,In_633,In_513);
and U893 (N_893,In_748,In_808);
xor U894 (N_894,In_30,In_139);
or U895 (N_895,In_168,In_559);
and U896 (N_896,In_465,In_82);
nand U897 (N_897,In_389,In_152);
nand U898 (N_898,In_518,In_677);
and U899 (N_899,In_169,In_959);
nor U900 (N_900,In_808,In_536);
or U901 (N_901,In_23,In_297);
nor U902 (N_902,In_472,In_707);
or U903 (N_903,In_85,In_445);
and U904 (N_904,In_940,In_464);
nand U905 (N_905,In_579,In_379);
nor U906 (N_906,In_706,In_674);
or U907 (N_907,In_244,In_956);
nand U908 (N_908,In_57,In_50);
xnor U909 (N_909,In_96,In_283);
xnor U910 (N_910,In_66,In_697);
xor U911 (N_911,In_706,In_510);
nand U912 (N_912,In_20,In_772);
nand U913 (N_913,In_283,In_441);
nand U914 (N_914,In_771,In_115);
nand U915 (N_915,In_778,In_770);
and U916 (N_916,In_856,In_242);
and U917 (N_917,In_557,In_678);
nand U918 (N_918,In_321,In_156);
nor U919 (N_919,In_685,In_449);
and U920 (N_920,In_825,In_450);
or U921 (N_921,In_132,In_668);
xor U922 (N_922,In_741,In_250);
and U923 (N_923,In_483,In_226);
nor U924 (N_924,In_371,In_729);
nand U925 (N_925,In_378,In_754);
nand U926 (N_926,In_139,In_313);
xor U927 (N_927,In_427,In_809);
or U928 (N_928,In_508,In_618);
or U929 (N_929,In_995,In_113);
nand U930 (N_930,In_554,In_90);
or U931 (N_931,In_38,In_142);
or U932 (N_932,In_245,In_425);
or U933 (N_933,In_233,In_133);
xor U934 (N_934,In_447,In_478);
nor U935 (N_935,In_534,In_723);
and U936 (N_936,In_851,In_53);
nand U937 (N_937,In_170,In_165);
and U938 (N_938,In_875,In_532);
and U939 (N_939,In_514,In_909);
nor U940 (N_940,In_177,In_724);
nor U941 (N_941,In_165,In_285);
and U942 (N_942,In_912,In_538);
or U943 (N_943,In_413,In_348);
nand U944 (N_944,In_497,In_558);
nand U945 (N_945,In_167,In_193);
nand U946 (N_946,In_74,In_874);
xor U947 (N_947,In_855,In_653);
or U948 (N_948,In_657,In_750);
and U949 (N_949,In_261,In_672);
nand U950 (N_950,In_687,In_287);
and U951 (N_951,In_118,In_19);
xor U952 (N_952,In_365,In_143);
nor U953 (N_953,In_872,In_949);
xnor U954 (N_954,In_783,In_947);
nand U955 (N_955,In_729,In_21);
and U956 (N_956,In_891,In_279);
and U957 (N_957,In_603,In_217);
nand U958 (N_958,In_823,In_200);
nor U959 (N_959,In_170,In_16);
nor U960 (N_960,In_269,In_159);
and U961 (N_961,In_473,In_600);
nor U962 (N_962,In_248,In_426);
or U963 (N_963,In_10,In_986);
xnor U964 (N_964,In_19,In_971);
or U965 (N_965,In_721,In_605);
and U966 (N_966,In_912,In_210);
or U967 (N_967,In_395,In_285);
xnor U968 (N_968,In_142,In_405);
nor U969 (N_969,In_323,In_767);
nand U970 (N_970,In_820,In_975);
nand U971 (N_971,In_66,In_520);
xnor U972 (N_972,In_122,In_491);
and U973 (N_973,In_985,In_522);
nor U974 (N_974,In_179,In_440);
nand U975 (N_975,In_352,In_730);
or U976 (N_976,In_202,In_817);
xnor U977 (N_977,In_194,In_887);
xnor U978 (N_978,In_133,In_514);
nor U979 (N_979,In_701,In_774);
and U980 (N_980,In_444,In_300);
xor U981 (N_981,In_483,In_770);
and U982 (N_982,In_688,In_433);
nand U983 (N_983,In_298,In_488);
nor U984 (N_984,In_698,In_179);
xor U985 (N_985,In_268,In_909);
or U986 (N_986,In_108,In_14);
and U987 (N_987,In_491,In_245);
nor U988 (N_988,In_179,In_105);
nor U989 (N_989,In_218,In_374);
and U990 (N_990,In_43,In_656);
nand U991 (N_991,In_403,In_951);
or U992 (N_992,In_974,In_603);
xnor U993 (N_993,In_664,In_394);
nand U994 (N_994,In_131,In_655);
and U995 (N_995,In_874,In_293);
xor U996 (N_996,In_10,In_909);
nor U997 (N_997,In_361,In_211);
nand U998 (N_998,In_762,In_508);
and U999 (N_999,In_877,In_7);
xor U1000 (N_1000,In_694,In_248);
nand U1001 (N_1001,In_277,In_444);
and U1002 (N_1002,In_164,In_479);
or U1003 (N_1003,In_305,In_45);
nor U1004 (N_1004,In_854,In_114);
nor U1005 (N_1005,In_45,In_523);
or U1006 (N_1006,In_796,In_495);
nand U1007 (N_1007,In_186,In_312);
and U1008 (N_1008,In_152,In_4);
nand U1009 (N_1009,In_757,In_627);
xnor U1010 (N_1010,In_449,In_311);
xor U1011 (N_1011,In_362,In_619);
and U1012 (N_1012,In_255,In_290);
xor U1013 (N_1013,In_8,In_179);
and U1014 (N_1014,In_139,In_808);
and U1015 (N_1015,In_345,In_454);
or U1016 (N_1016,In_597,In_582);
nand U1017 (N_1017,In_321,In_163);
and U1018 (N_1018,In_323,In_30);
and U1019 (N_1019,In_309,In_51);
xor U1020 (N_1020,In_524,In_273);
or U1021 (N_1021,In_683,In_993);
xnor U1022 (N_1022,In_229,In_679);
nor U1023 (N_1023,In_825,In_683);
nor U1024 (N_1024,In_790,In_776);
nand U1025 (N_1025,In_235,In_427);
nand U1026 (N_1026,In_277,In_506);
or U1027 (N_1027,In_439,In_789);
nand U1028 (N_1028,In_968,In_858);
and U1029 (N_1029,In_733,In_953);
xnor U1030 (N_1030,In_531,In_753);
nand U1031 (N_1031,In_416,In_864);
nand U1032 (N_1032,In_365,In_391);
and U1033 (N_1033,In_528,In_872);
or U1034 (N_1034,In_193,In_115);
xor U1035 (N_1035,In_502,In_634);
and U1036 (N_1036,In_581,In_916);
and U1037 (N_1037,In_463,In_113);
nor U1038 (N_1038,In_400,In_836);
nor U1039 (N_1039,In_796,In_850);
or U1040 (N_1040,In_796,In_448);
xor U1041 (N_1041,In_706,In_495);
nand U1042 (N_1042,In_368,In_923);
and U1043 (N_1043,In_482,In_767);
or U1044 (N_1044,In_811,In_729);
or U1045 (N_1045,In_742,In_519);
nand U1046 (N_1046,In_528,In_804);
xnor U1047 (N_1047,In_850,In_894);
nand U1048 (N_1048,In_983,In_774);
or U1049 (N_1049,In_509,In_297);
xnor U1050 (N_1050,In_74,In_564);
or U1051 (N_1051,In_988,In_903);
nor U1052 (N_1052,In_597,In_87);
xnor U1053 (N_1053,In_475,In_864);
nor U1054 (N_1054,In_320,In_818);
xnor U1055 (N_1055,In_893,In_924);
or U1056 (N_1056,In_850,In_564);
and U1057 (N_1057,In_497,In_710);
nor U1058 (N_1058,In_685,In_797);
or U1059 (N_1059,In_179,In_120);
or U1060 (N_1060,In_35,In_203);
or U1061 (N_1061,In_58,In_281);
nor U1062 (N_1062,In_124,In_407);
nor U1063 (N_1063,In_749,In_88);
and U1064 (N_1064,In_975,In_458);
xor U1065 (N_1065,In_303,In_453);
xor U1066 (N_1066,In_818,In_914);
or U1067 (N_1067,In_792,In_343);
xor U1068 (N_1068,In_441,In_201);
nand U1069 (N_1069,In_58,In_232);
xor U1070 (N_1070,In_49,In_302);
or U1071 (N_1071,In_260,In_273);
and U1072 (N_1072,In_783,In_181);
nor U1073 (N_1073,In_331,In_961);
and U1074 (N_1074,In_164,In_440);
nor U1075 (N_1075,In_339,In_617);
and U1076 (N_1076,In_648,In_201);
or U1077 (N_1077,In_607,In_623);
xor U1078 (N_1078,In_755,In_906);
and U1079 (N_1079,In_587,In_235);
nor U1080 (N_1080,In_486,In_229);
nor U1081 (N_1081,In_394,In_241);
nor U1082 (N_1082,In_632,In_215);
or U1083 (N_1083,In_642,In_532);
nand U1084 (N_1084,In_140,In_851);
and U1085 (N_1085,In_667,In_588);
nor U1086 (N_1086,In_576,In_661);
xor U1087 (N_1087,In_608,In_381);
or U1088 (N_1088,In_342,In_212);
xor U1089 (N_1089,In_744,In_216);
nor U1090 (N_1090,In_559,In_635);
nand U1091 (N_1091,In_904,In_484);
or U1092 (N_1092,In_144,In_45);
and U1093 (N_1093,In_79,In_925);
xor U1094 (N_1094,In_343,In_200);
nor U1095 (N_1095,In_200,In_99);
nand U1096 (N_1096,In_702,In_911);
nand U1097 (N_1097,In_627,In_969);
nor U1098 (N_1098,In_345,In_875);
and U1099 (N_1099,In_722,In_875);
xnor U1100 (N_1100,In_32,In_924);
nand U1101 (N_1101,In_222,In_542);
nor U1102 (N_1102,In_439,In_171);
or U1103 (N_1103,In_93,In_473);
or U1104 (N_1104,In_433,In_340);
xnor U1105 (N_1105,In_495,In_318);
or U1106 (N_1106,In_450,In_316);
xnor U1107 (N_1107,In_836,In_388);
nor U1108 (N_1108,In_346,In_271);
nor U1109 (N_1109,In_256,In_899);
nand U1110 (N_1110,In_172,In_880);
and U1111 (N_1111,In_395,In_242);
nor U1112 (N_1112,In_439,In_653);
nor U1113 (N_1113,In_834,In_110);
or U1114 (N_1114,In_325,In_389);
and U1115 (N_1115,In_537,In_353);
nand U1116 (N_1116,In_45,In_540);
or U1117 (N_1117,In_42,In_959);
and U1118 (N_1118,In_763,In_587);
or U1119 (N_1119,In_467,In_120);
nand U1120 (N_1120,In_945,In_950);
or U1121 (N_1121,In_943,In_155);
nand U1122 (N_1122,In_975,In_205);
nor U1123 (N_1123,In_827,In_55);
or U1124 (N_1124,In_861,In_545);
or U1125 (N_1125,In_202,In_482);
nand U1126 (N_1126,In_991,In_273);
and U1127 (N_1127,In_965,In_467);
xnor U1128 (N_1128,In_410,In_13);
xor U1129 (N_1129,In_802,In_445);
or U1130 (N_1130,In_27,In_991);
xor U1131 (N_1131,In_652,In_871);
nor U1132 (N_1132,In_258,In_361);
xnor U1133 (N_1133,In_167,In_585);
and U1134 (N_1134,In_820,In_13);
nand U1135 (N_1135,In_292,In_229);
nand U1136 (N_1136,In_566,In_489);
or U1137 (N_1137,In_246,In_648);
nor U1138 (N_1138,In_158,In_856);
and U1139 (N_1139,In_110,In_37);
xor U1140 (N_1140,In_348,In_983);
nand U1141 (N_1141,In_260,In_171);
or U1142 (N_1142,In_946,In_628);
nand U1143 (N_1143,In_990,In_968);
or U1144 (N_1144,In_530,In_682);
nand U1145 (N_1145,In_847,In_239);
nor U1146 (N_1146,In_493,In_534);
and U1147 (N_1147,In_681,In_41);
nand U1148 (N_1148,In_411,In_750);
or U1149 (N_1149,In_187,In_62);
xnor U1150 (N_1150,In_743,In_974);
nand U1151 (N_1151,In_344,In_719);
nand U1152 (N_1152,In_712,In_623);
or U1153 (N_1153,In_669,In_374);
nor U1154 (N_1154,In_653,In_661);
and U1155 (N_1155,In_744,In_605);
nor U1156 (N_1156,In_54,In_588);
and U1157 (N_1157,In_24,In_769);
and U1158 (N_1158,In_941,In_202);
and U1159 (N_1159,In_826,In_343);
nor U1160 (N_1160,In_711,In_390);
xor U1161 (N_1161,In_940,In_302);
nor U1162 (N_1162,In_368,In_459);
nand U1163 (N_1163,In_109,In_627);
nand U1164 (N_1164,In_222,In_702);
xnor U1165 (N_1165,In_15,In_559);
nor U1166 (N_1166,In_427,In_281);
and U1167 (N_1167,In_666,In_603);
and U1168 (N_1168,In_307,In_822);
nand U1169 (N_1169,In_804,In_287);
and U1170 (N_1170,In_722,In_657);
xnor U1171 (N_1171,In_606,In_329);
and U1172 (N_1172,In_982,In_901);
xor U1173 (N_1173,In_606,In_268);
xnor U1174 (N_1174,In_146,In_288);
xnor U1175 (N_1175,In_288,In_149);
nand U1176 (N_1176,In_861,In_628);
or U1177 (N_1177,In_619,In_687);
nor U1178 (N_1178,In_827,In_868);
nand U1179 (N_1179,In_903,In_580);
xor U1180 (N_1180,In_850,In_157);
and U1181 (N_1181,In_479,In_499);
nor U1182 (N_1182,In_587,In_392);
nand U1183 (N_1183,In_749,In_563);
nand U1184 (N_1184,In_52,In_280);
xor U1185 (N_1185,In_870,In_987);
xor U1186 (N_1186,In_49,In_785);
or U1187 (N_1187,In_591,In_29);
xor U1188 (N_1188,In_11,In_612);
or U1189 (N_1189,In_730,In_212);
and U1190 (N_1190,In_919,In_3);
or U1191 (N_1191,In_579,In_349);
and U1192 (N_1192,In_433,In_617);
xnor U1193 (N_1193,In_574,In_578);
nand U1194 (N_1194,In_191,In_635);
and U1195 (N_1195,In_230,In_996);
xor U1196 (N_1196,In_732,In_858);
nor U1197 (N_1197,In_737,In_562);
nor U1198 (N_1198,In_778,In_872);
xnor U1199 (N_1199,In_695,In_583);
or U1200 (N_1200,In_842,In_962);
or U1201 (N_1201,In_174,In_797);
nand U1202 (N_1202,In_254,In_210);
xnor U1203 (N_1203,In_840,In_849);
nand U1204 (N_1204,In_816,In_542);
nor U1205 (N_1205,In_952,In_146);
and U1206 (N_1206,In_222,In_340);
xor U1207 (N_1207,In_599,In_334);
nand U1208 (N_1208,In_960,In_280);
or U1209 (N_1209,In_236,In_784);
nor U1210 (N_1210,In_955,In_944);
or U1211 (N_1211,In_882,In_815);
nor U1212 (N_1212,In_459,In_235);
and U1213 (N_1213,In_913,In_318);
or U1214 (N_1214,In_125,In_687);
xnor U1215 (N_1215,In_935,In_588);
nor U1216 (N_1216,In_366,In_161);
nand U1217 (N_1217,In_398,In_301);
or U1218 (N_1218,In_307,In_898);
and U1219 (N_1219,In_182,In_256);
or U1220 (N_1220,In_259,In_793);
nor U1221 (N_1221,In_649,In_991);
xnor U1222 (N_1222,In_531,In_80);
xor U1223 (N_1223,In_222,In_203);
nor U1224 (N_1224,In_245,In_89);
and U1225 (N_1225,In_965,In_265);
and U1226 (N_1226,In_503,In_252);
nor U1227 (N_1227,In_108,In_263);
and U1228 (N_1228,In_852,In_548);
nand U1229 (N_1229,In_141,In_467);
or U1230 (N_1230,In_319,In_819);
and U1231 (N_1231,In_363,In_953);
and U1232 (N_1232,In_839,In_506);
nand U1233 (N_1233,In_190,In_743);
xnor U1234 (N_1234,In_848,In_88);
or U1235 (N_1235,In_574,In_362);
nand U1236 (N_1236,In_737,In_835);
and U1237 (N_1237,In_496,In_671);
nand U1238 (N_1238,In_560,In_267);
or U1239 (N_1239,In_695,In_115);
nand U1240 (N_1240,In_760,In_667);
nand U1241 (N_1241,In_854,In_909);
nor U1242 (N_1242,In_804,In_921);
nor U1243 (N_1243,In_763,In_726);
xnor U1244 (N_1244,In_979,In_857);
and U1245 (N_1245,In_215,In_595);
or U1246 (N_1246,In_973,In_433);
or U1247 (N_1247,In_991,In_842);
nand U1248 (N_1248,In_486,In_69);
nor U1249 (N_1249,In_16,In_782);
or U1250 (N_1250,In_814,In_626);
and U1251 (N_1251,In_850,In_332);
or U1252 (N_1252,In_460,In_169);
and U1253 (N_1253,In_908,In_340);
nor U1254 (N_1254,In_39,In_445);
nand U1255 (N_1255,In_722,In_309);
or U1256 (N_1256,In_189,In_151);
nor U1257 (N_1257,In_79,In_354);
and U1258 (N_1258,In_74,In_89);
and U1259 (N_1259,In_621,In_971);
nand U1260 (N_1260,In_737,In_621);
nor U1261 (N_1261,In_941,In_529);
nand U1262 (N_1262,In_341,In_848);
xnor U1263 (N_1263,In_62,In_436);
or U1264 (N_1264,In_906,In_330);
nor U1265 (N_1265,In_797,In_661);
xor U1266 (N_1266,In_323,In_124);
xnor U1267 (N_1267,In_1,In_112);
and U1268 (N_1268,In_616,In_906);
nor U1269 (N_1269,In_93,In_648);
nand U1270 (N_1270,In_655,In_170);
and U1271 (N_1271,In_251,In_48);
xnor U1272 (N_1272,In_412,In_484);
xor U1273 (N_1273,In_497,In_693);
and U1274 (N_1274,In_922,In_208);
nand U1275 (N_1275,In_272,In_219);
nor U1276 (N_1276,In_122,In_401);
nor U1277 (N_1277,In_263,In_644);
and U1278 (N_1278,In_601,In_96);
nor U1279 (N_1279,In_515,In_546);
nor U1280 (N_1280,In_447,In_306);
nor U1281 (N_1281,In_604,In_552);
xor U1282 (N_1282,In_776,In_475);
and U1283 (N_1283,In_506,In_88);
nor U1284 (N_1284,In_543,In_498);
nor U1285 (N_1285,In_963,In_15);
nand U1286 (N_1286,In_727,In_427);
nand U1287 (N_1287,In_9,In_266);
and U1288 (N_1288,In_436,In_207);
or U1289 (N_1289,In_268,In_661);
or U1290 (N_1290,In_757,In_812);
nand U1291 (N_1291,In_33,In_531);
xor U1292 (N_1292,In_561,In_681);
nand U1293 (N_1293,In_467,In_578);
nand U1294 (N_1294,In_985,In_371);
or U1295 (N_1295,In_89,In_229);
nand U1296 (N_1296,In_770,In_891);
nor U1297 (N_1297,In_687,In_370);
nor U1298 (N_1298,In_485,In_844);
or U1299 (N_1299,In_131,In_154);
nor U1300 (N_1300,In_41,In_855);
nand U1301 (N_1301,In_408,In_810);
nor U1302 (N_1302,In_497,In_72);
nand U1303 (N_1303,In_596,In_812);
nand U1304 (N_1304,In_928,In_652);
and U1305 (N_1305,In_973,In_876);
and U1306 (N_1306,In_372,In_111);
nor U1307 (N_1307,In_948,In_596);
and U1308 (N_1308,In_472,In_624);
xor U1309 (N_1309,In_620,In_635);
or U1310 (N_1310,In_843,In_621);
xnor U1311 (N_1311,In_507,In_302);
nor U1312 (N_1312,In_65,In_522);
and U1313 (N_1313,In_594,In_838);
xnor U1314 (N_1314,In_253,In_6);
nor U1315 (N_1315,In_345,In_831);
nand U1316 (N_1316,In_49,In_790);
and U1317 (N_1317,In_714,In_316);
and U1318 (N_1318,In_297,In_890);
or U1319 (N_1319,In_788,In_472);
nor U1320 (N_1320,In_627,In_93);
and U1321 (N_1321,In_35,In_952);
xnor U1322 (N_1322,In_97,In_978);
nand U1323 (N_1323,In_186,In_301);
xnor U1324 (N_1324,In_345,In_934);
nand U1325 (N_1325,In_710,In_596);
or U1326 (N_1326,In_11,In_315);
and U1327 (N_1327,In_787,In_426);
nand U1328 (N_1328,In_614,In_113);
nor U1329 (N_1329,In_125,In_239);
nand U1330 (N_1330,In_785,In_252);
or U1331 (N_1331,In_48,In_936);
xnor U1332 (N_1332,In_33,In_106);
xnor U1333 (N_1333,In_244,In_12);
nand U1334 (N_1334,In_197,In_348);
nor U1335 (N_1335,In_629,In_590);
and U1336 (N_1336,In_484,In_697);
or U1337 (N_1337,In_557,In_996);
nor U1338 (N_1338,In_94,In_537);
and U1339 (N_1339,In_795,In_323);
xor U1340 (N_1340,In_445,In_256);
xor U1341 (N_1341,In_749,In_250);
and U1342 (N_1342,In_561,In_823);
xor U1343 (N_1343,In_308,In_439);
xor U1344 (N_1344,In_223,In_490);
or U1345 (N_1345,In_553,In_970);
or U1346 (N_1346,In_338,In_824);
and U1347 (N_1347,In_824,In_948);
or U1348 (N_1348,In_792,In_54);
and U1349 (N_1349,In_445,In_109);
xor U1350 (N_1350,In_878,In_631);
nor U1351 (N_1351,In_369,In_326);
xor U1352 (N_1352,In_631,In_563);
xor U1353 (N_1353,In_430,In_789);
and U1354 (N_1354,In_927,In_937);
and U1355 (N_1355,In_798,In_958);
nand U1356 (N_1356,In_588,In_912);
or U1357 (N_1357,In_833,In_313);
or U1358 (N_1358,In_752,In_358);
nand U1359 (N_1359,In_950,In_728);
or U1360 (N_1360,In_418,In_236);
and U1361 (N_1361,In_14,In_333);
or U1362 (N_1362,In_69,In_281);
nor U1363 (N_1363,In_346,In_546);
and U1364 (N_1364,In_318,In_451);
or U1365 (N_1365,In_551,In_74);
or U1366 (N_1366,In_849,In_66);
and U1367 (N_1367,In_710,In_91);
and U1368 (N_1368,In_270,In_691);
or U1369 (N_1369,In_71,In_219);
nor U1370 (N_1370,In_50,In_278);
xnor U1371 (N_1371,In_760,In_552);
nand U1372 (N_1372,In_124,In_750);
and U1373 (N_1373,In_517,In_117);
nor U1374 (N_1374,In_437,In_752);
or U1375 (N_1375,In_517,In_333);
or U1376 (N_1376,In_394,In_805);
nand U1377 (N_1377,In_590,In_355);
or U1378 (N_1378,In_5,In_375);
xor U1379 (N_1379,In_143,In_231);
or U1380 (N_1380,In_461,In_427);
nand U1381 (N_1381,In_306,In_489);
nor U1382 (N_1382,In_806,In_653);
nor U1383 (N_1383,In_54,In_733);
and U1384 (N_1384,In_381,In_960);
nor U1385 (N_1385,In_27,In_401);
nor U1386 (N_1386,In_892,In_927);
nand U1387 (N_1387,In_37,In_872);
or U1388 (N_1388,In_410,In_830);
xor U1389 (N_1389,In_460,In_777);
nand U1390 (N_1390,In_244,In_53);
and U1391 (N_1391,In_73,In_681);
xnor U1392 (N_1392,In_181,In_85);
and U1393 (N_1393,In_736,In_94);
nand U1394 (N_1394,In_317,In_919);
nand U1395 (N_1395,In_67,In_492);
or U1396 (N_1396,In_293,In_109);
and U1397 (N_1397,In_579,In_648);
xor U1398 (N_1398,In_175,In_692);
nor U1399 (N_1399,In_833,In_83);
and U1400 (N_1400,In_584,In_339);
or U1401 (N_1401,In_140,In_995);
or U1402 (N_1402,In_822,In_889);
xnor U1403 (N_1403,In_334,In_30);
and U1404 (N_1404,In_300,In_595);
and U1405 (N_1405,In_166,In_658);
or U1406 (N_1406,In_808,In_407);
and U1407 (N_1407,In_55,In_67);
nor U1408 (N_1408,In_594,In_755);
nand U1409 (N_1409,In_38,In_378);
nand U1410 (N_1410,In_103,In_123);
or U1411 (N_1411,In_617,In_323);
or U1412 (N_1412,In_801,In_961);
nand U1413 (N_1413,In_889,In_279);
and U1414 (N_1414,In_214,In_328);
xor U1415 (N_1415,In_752,In_205);
nand U1416 (N_1416,In_749,In_387);
nor U1417 (N_1417,In_346,In_695);
and U1418 (N_1418,In_40,In_681);
nor U1419 (N_1419,In_356,In_2);
nand U1420 (N_1420,In_935,In_88);
nor U1421 (N_1421,In_488,In_212);
xnor U1422 (N_1422,In_435,In_285);
and U1423 (N_1423,In_567,In_654);
and U1424 (N_1424,In_209,In_808);
and U1425 (N_1425,In_642,In_991);
or U1426 (N_1426,In_881,In_816);
xor U1427 (N_1427,In_374,In_223);
nand U1428 (N_1428,In_231,In_14);
and U1429 (N_1429,In_136,In_848);
or U1430 (N_1430,In_494,In_584);
xnor U1431 (N_1431,In_877,In_523);
or U1432 (N_1432,In_917,In_105);
nor U1433 (N_1433,In_959,In_637);
and U1434 (N_1434,In_627,In_565);
nor U1435 (N_1435,In_832,In_794);
or U1436 (N_1436,In_896,In_48);
nor U1437 (N_1437,In_182,In_467);
xor U1438 (N_1438,In_234,In_400);
or U1439 (N_1439,In_280,In_638);
xor U1440 (N_1440,In_622,In_620);
or U1441 (N_1441,In_664,In_587);
nor U1442 (N_1442,In_504,In_657);
xnor U1443 (N_1443,In_304,In_533);
xor U1444 (N_1444,In_550,In_374);
and U1445 (N_1445,In_405,In_549);
xnor U1446 (N_1446,In_745,In_161);
and U1447 (N_1447,In_533,In_468);
or U1448 (N_1448,In_498,In_532);
and U1449 (N_1449,In_845,In_265);
nand U1450 (N_1450,In_48,In_649);
and U1451 (N_1451,In_322,In_438);
nand U1452 (N_1452,In_777,In_543);
nor U1453 (N_1453,In_442,In_290);
nand U1454 (N_1454,In_252,In_780);
or U1455 (N_1455,In_302,In_15);
and U1456 (N_1456,In_604,In_143);
xnor U1457 (N_1457,In_936,In_51);
nor U1458 (N_1458,In_831,In_286);
and U1459 (N_1459,In_706,In_421);
nor U1460 (N_1460,In_234,In_966);
xnor U1461 (N_1461,In_366,In_113);
nand U1462 (N_1462,In_482,In_230);
or U1463 (N_1463,In_176,In_266);
or U1464 (N_1464,In_971,In_677);
or U1465 (N_1465,In_976,In_275);
and U1466 (N_1466,In_623,In_102);
xor U1467 (N_1467,In_342,In_382);
and U1468 (N_1468,In_158,In_470);
xnor U1469 (N_1469,In_97,In_252);
nor U1470 (N_1470,In_209,In_622);
and U1471 (N_1471,In_317,In_341);
or U1472 (N_1472,In_792,In_614);
and U1473 (N_1473,In_626,In_857);
xor U1474 (N_1474,In_187,In_626);
or U1475 (N_1475,In_788,In_340);
nor U1476 (N_1476,In_675,In_354);
nand U1477 (N_1477,In_969,In_922);
and U1478 (N_1478,In_896,In_822);
and U1479 (N_1479,In_115,In_96);
or U1480 (N_1480,In_126,In_839);
nor U1481 (N_1481,In_819,In_310);
nor U1482 (N_1482,In_854,In_347);
nand U1483 (N_1483,In_418,In_865);
nor U1484 (N_1484,In_142,In_882);
and U1485 (N_1485,In_428,In_850);
nand U1486 (N_1486,In_66,In_738);
or U1487 (N_1487,In_733,In_162);
nand U1488 (N_1488,In_897,In_120);
or U1489 (N_1489,In_809,In_209);
or U1490 (N_1490,In_518,In_50);
or U1491 (N_1491,In_949,In_945);
nand U1492 (N_1492,In_13,In_840);
and U1493 (N_1493,In_184,In_55);
nand U1494 (N_1494,In_109,In_251);
or U1495 (N_1495,In_411,In_928);
xnor U1496 (N_1496,In_264,In_512);
and U1497 (N_1497,In_263,In_882);
nor U1498 (N_1498,In_215,In_634);
or U1499 (N_1499,In_239,In_340);
xnor U1500 (N_1500,In_933,In_237);
nand U1501 (N_1501,In_838,In_267);
nor U1502 (N_1502,In_716,In_422);
nor U1503 (N_1503,In_314,In_360);
or U1504 (N_1504,In_84,In_872);
or U1505 (N_1505,In_460,In_304);
xor U1506 (N_1506,In_843,In_458);
nor U1507 (N_1507,In_373,In_161);
and U1508 (N_1508,In_174,In_349);
xor U1509 (N_1509,In_943,In_617);
and U1510 (N_1510,In_397,In_820);
nor U1511 (N_1511,In_283,In_333);
xor U1512 (N_1512,In_587,In_916);
and U1513 (N_1513,In_979,In_781);
and U1514 (N_1514,In_481,In_403);
xnor U1515 (N_1515,In_875,In_113);
or U1516 (N_1516,In_295,In_525);
xor U1517 (N_1517,In_59,In_809);
and U1518 (N_1518,In_536,In_675);
or U1519 (N_1519,In_716,In_724);
nand U1520 (N_1520,In_367,In_351);
nand U1521 (N_1521,In_699,In_576);
nor U1522 (N_1522,In_588,In_323);
and U1523 (N_1523,In_4,In_561);
and U1524 (N_1524,In_558,In_693);
or U1525 (N_1525,In_739,In_270);
xor U1526 (N_1526,In_698,In_55);
nand U1527 (N_1527,In_528,In_64);
or U1528 (N_1528,In_633,In_74);
nand U1529 (N_1529,In_172,In_866);
nor U1530 (N_1530,In_640,In_284);
or U1531 (N_1531,In_617,In_914);
and U1532 (N_1532,In_838,In_522);
or U1533 (N_1533,In_501,In_19);
and U1534 (N_1534,In_580,In_880);
xnor U1535 (N_1535,In_54,In_516);
and U1536 (N_1536,In_26,In_413);
nand U1537 (N_1537,In_901,In_897);
xor U1538 (N_1538,In_138,In_262);
xor U1539 (N_1539,In_875,In_515);
xnor U1540 (N_1540,In_9,In_278);
and U1541 (N_1541,In_66,In_141);
nor U1542 (N_1542,In_504,In_420);
or U1543 (N_1543,In_760,In_792);
nand U1544 (N_1544,In_765,In_303);
xor U1545 (N_1545,In_110,In_52);
nor U1546 (N_1546,In_168,In_190);
xor U1547 (N_1547,In_978,In_604);
nand U1548 (N_1548,In_359,In_520);
and U1549 (N_1549,In_900,In_659);
and U1550 (N_1550,In_524,In_585);
or U1551 (N_1551,In_175,In_385);
xor U1552 (N_1552,In_427,In_165);
and U1553 (N_1553,In_359,In_957);
xnor U1554 (N_1554,In_783,In_787);
nand U1555 (N_1555,In_1,In_608);
xor U1556 (N_1556,In_866,In_300);
nand U1557 (N_1557,In_758,In_235);
xor U1558 (N_1558,In_395,In_810);
xor U1559 (N_1559,In_44,In_608);
and U1560 (N_1560,In_916,In_992);
nor U1561 (N_1561,In_104,In_895);
or U1562 (N_1562,In_115,In_993);
and U1563 (N_1563,In_148,In_816);
nand U1564 (N_1564,In_940,In_237);
nand U1565 (N_1565,In_740,In_590);
or U1566 (N_1566,In_807,In_410);
nor U1567 (N_1567,In_490,In_95);
nand U1568 (N_1568,In_683,In_855);
and U1569 (N_1569,In_320,In_637);
nor U1570 (N_1570,In_358,In_714);
or U1571 (N_1571,In_593,In_726);
and U1572 (N_1572,In_334,In_576);
nor U1573 (N_1573,In_982,In_959);
or U1574 (N_1574,In_455,In_126);
xnor U1575 (N_1575,In_133,In_733);
xor U1576 (N_1576,In_727,In_358);
nor U1577 (N_1577,In_746,In_36);
xor U1578 (N_1578,In_125,In_306);
nor U1579 (N_1579,In_837,In_102);
nor U1580 (N_1580,In_322,In_632);
or U1581 (N_1581,In_416,In_692);
nor U1582 (N_1582,In_657,In_87);
nor U1583 (N_1583,In_450,In_237);
xnor U1584 (N_1584,In_884,In_704);
or U1585 (N_1585,In_757,In_811);
or U1586 (N_1586,In_990,In_400);
xnor U1587 (N_1587,In_999,In_30);
nand U1588 (N_1588,In_672,In_95);
xor U1589 (N_1589,In_56,In_993);
nor U1590 (N_1590,In_735,In_515);
nand U1591 (N_1591,In_547,In_421);
nand U1592 (N_1592,In_239,In_956);
xnor U1593 (N_1593,In_171,In_518);
nor U1594 (N_1594,In_852,In_958);
nand U1595 (N_1595,In_168,In_611);
and U1596 (N_1596,In_398,In_121);
nand U1597 (N_1597,In_468,In_522);
nand U1598 (N_1598,In_783,In_194);
and U1599 (N_1599,In_274,In_724);
and U1600 (N_1600,In_285,In_712);
nand U1601 (N_1601,In_594,In_472);
xor U1602 (N_1602,In_807,In_949);
xor U1603 (N_1603,In_800,In_205);
nor U1604 (N_1604,In_274,In_49);
nor U1605 (N_1605,In_146,In_381);
or U1606 (N_1606,In_716,In_11);
or U1607 (N_1607,In_960,In_391);
xor U1608 (N_1608,In_213,In_132);
xnor U1609 (N_1609,In_805,In_907);
xnor U1610 (N_1610,In_932,In_765);
nor U1611 (N_1611,In_250,In_65);
nand U1612 (N_1612,In_116,In_443);
nor U1613 (N_1613,In_317,In_794);
and U1614 (N_1614,In_451,In_77);
nand U1615 (N_1615,In_337,In_688);
or U1616 (N_1616,In_855,In_691);
xnor U1617 (N_1617,In_991,In_775);
or U1618 (N_1618,In_592,In_740);
nor U1619 (N_1619,In_979,In_991);
nor U1620 (N_1620,In_903,In_262);
nand U1621 (N_1621,In_471,In_614);
and U1622 (N_1622,In_843,In_72);
nand U1623 (N_1623,In_177,In_572);
or U1624 (N_1624,In_173,In_769);
nand U1625 (N_1625,In_393,In_652);
nand U1626 (N_1626,In_946,In_330);
xor U1627 (N_1627,In_304,In_498);
or U1628 (N_1628,In_649,In_752);
nor U1629 (N_1629,In_263,In_635);
or U1630 (N_1630,In_332,In_555);
and U1631 (N_1631,In_893,In_340);
nor U1632 (N_1632,In_915,In_584);
or U1633 (N_1633,In_609,In_56);
or U1634 (N_1634,In_459,In_483);
and U1635 (N_1635,In_584,In_504);
xnor U1636 (N_1636,In_310,In_40);
nand U1637 (N_1637,In_937,In_87);
or U1638 (N_1638,In_862,In_897);
xnor U1639 (N_1639,In_232,In_588);
and U1640 (N_1640,In_15,In_442);
nand U1641 (N_1641,In_267,In_581);
and U1642 (N_1642,In_570,In_636);
or U1643 (N_1643,In_987,In_137);
xnor U1644 (N_1644,In_66,In_455);
xor U1645 (N_1645,In_710,In_680);
nand U1646 (N_1646,In_74,In_799);
xnor U1647 (N_1647,In_834,In_819);
xor U1648 (N_1648,In_760,In_133);
or U1649 (N_1649,In_468,In_720);
nor U1650 (N_1650,In_403,In_577);
nor U1651 (N_1651,In_589,In_928);
or U1652 (N_1652,In_249,In_411);
nor U1653 (N_1653,In_888,In_648);
nand U1654 (N_1654,In_410,In_15);
xor U1655 (N_1655,In_55,In_900);
xor U1656 (N_1656,In_666,In_514);
nand U1657 (N_1657,In_393,In_164);
or U1658 (N_1658,In_595,In_817);
or U1659 (N_1659,In_851,In_938);
and U1660 (N_1660,In_306,In_798);
nor U1661 (N_1661,In_670,In_644);
or U1662 (N_1662,In_187,In_975);
xor U1663 (N_1663,In_687,In_77);
xnor U1664 (N_1664,In_542,In_129);
xor U1665 (N_1665,In_865,In_110);
nor U1666 (N_1666,In_517,In_713);
or U1667 (N_1667,In_828,In_310);
nand U1668 (N_1668,In_169,In_43);
or U1669 (N_1669,In_415,In_109);
xor U1670 (N_1670,In_704,In_997);
nor U1671 (N_1671,In_495,In_941);
or U1672 (N_1672,In_183,In_36);
or U1673 (N_1673,In_361,In_108);
and U1674 (N_1674,In_125,In_218);
nand U1675 (N_1675,In_350,In_22);
nand U1676 (N_1676,In_558,In_67);
nand U1677 (N_1677,In_524,In_604);
or U1678 (N_1678,In_988,In_732);
nand U1679 (N_1679,In_654,In_298);
nor U1680 (N_1680,In_338,In_511);
xor U1681 (N_1681,In_270,In_729);
or U1682 (N_1682,In_188,In_58);
nor U1683 (N_1683,In_783,In_802);
nor U1684 (N_1684,In_89,In_331);
nand U1685 (N_1685,In_211,In_346);
nor U1686 (N_1686,In_414,In_378);
and U1687 (N_1687,In_999,In_996);
and U1688 (N_1688,In_678,In_120);
and U1689 (N_1689,In_244,In_986);
nand U1690 (N_1690,In_155,In_462);
and U1691 (N_1691,In_499,In_914);
nand U1692 (N_1692,In_532,In_291);
or U1693 (N_1693,In_821,In_792);
nor U1694 (N_1694,In_5,In_88);
xor U1695 (N_1695,In_175,In_193);
xor U1696 (N_1696,In_409,In_107);
nor U1697 (N_1697,In_700,In_225);
and U1698 (N_1698,In_243,In_370);
nor U1699 (N_1699,In_130,In_99);
xor U1700 (N_1700,In_132,In_803);
nand U1701 (N_1701,In_442,In_663);
or U1702 (N_1702,In_100,In_804);
and U1703 (N_1703,In_152,In_373);
or U1704 (N_1704,In_634,In_346);
and U1705 (N_1705,In_478,In_473);
or U1706 (N_1706,In_542,In_335);
or U1707 (N_1707,In_719,In_832);
and U1708 (N_1708,In_533,In_979);
nand U1709 (N_1709,In_727,In_715);
xor U1710 (N_1710,In_504,In_493);
nand U1711 (N_1711,In_113,In_277);
and U1712 (N_1712,In_406,In_823);
and U1713 (N_1713,In_815,In_645);
nand U1714 (N_1714,In_675,In_981);
nand U1715 (N_1715,In_629,In_604);
or U1716 (N_1716,In_808,In_519);
and U1717 (N_1717,In_861,In_978);
and U1718 (N_1718,In_310,In_311);
nand U1719 (N_1719,In_176,In_871);
xor U1720 (N_1720,In_826,In_568);
nor U1721 (N_1721,In_435,In_958);
xor U1722 (N_1722,In_891,In_550);
and U1723 (N_1723,In_636,In_879);
or U1724 (N_1724,In_874,In_188);
xnor U1725 (N_1725,In_244,In_417);
nand U1726 (N_1726,In_729,In_342);
nand U1727 (N_1727,In_737,In_330);
nor U1728 (N_1728,In_216,In_33);
nor U1729 (N_1729,In_918,In_639);
and U1730 (N_1730,In_596,In_766);
or U1731 (N_1731,In_365,In_153);
and U1732 (N_1732,In_359,In_977);
xnor U1733 (N_1733,In_116,In_363);
nor U1734 (N_1734,In_348,In_281);
nor U1735 (N_1735,In_583,In_36);
xnor U1736 (N_1736,In_743,In_232);
and U1737 (N_1737,In_187,In_856);
nor U1738 (N_1738,In_391,In_86);
and U1739 (N_1739,In_608,In_306);
xnor U1740 (N_1740,In_423,In_710);
and U1741 (N_1741,In_248,In_291);
xor U1742 (N_1742,In_467,In_908);
or U1743 (N_1743,In_526,In_749);
xnor U1744 (N_1744,In_351,In_270);
nor U1745 (N_1745,In_257,In_381);
nor U1746 (N_1746,In_8,In_144);
and U1747 (N_1747,In_604,In_737);
xor U1748 (N_1748,In_316,In_842);
nor U1749 (N_1749,In_384,In_91);
and U1750 (N_1750,In_348,In_870);
xor U1751 (N_1751,In_304,In_997);
nor U1752 (N_1752,In_224,In_346);
xor U1753 (N_1753,In_795,In_3);
xor U1754 (N_1754,In_864,In_970);
nor U1755 (N_1755,In_581,In_584);
nor U1756 (N_1756,In_216,In_633);
xor U1757 (N_1757,In_373,In_950);
and U1758 (N_1758,In_839,In_596);
or U1759 (N_1759,In_730,In_431);
or U1760 (N_1760,In_985,In_798);
and U1761 (N_1761,In_118,In_665);
nand U1762 (N_1762,In_457,In_181);
nand U1763 (N_1763,In_336,In_901);
xnor U1764 (N_1764,In_167,In_317);
xnor U1765 (N_1765,In_555,In_536);
nor U1766 (N_1766,In_149,In_966);
nor U1767 (N_1767,In_211,In_154);
nand U1768 (N_1768,In_582,In_901);
nor U1769 (N_1769,In_823,In_609);
xnor U1770 (N_1770,In_420,In_55);
or U1771 (N_1771,In_386,In_509);
nor U1772 (N_1772,In_497,In_236);
nor U1773 (N_1773,In_553,In_456);
nand U1774 (N_1774,In_810,In_102);
or U1775 (N_1775,In_244,In_740);
xor U1776 (N_1776,In_166,In_879);
or U1777 (N_1777,In_512,In_65);
and U1778 (N_1778,In_308,In_39);
xnor U1779 (N_1779,In_803,In_21);
nor U1780 (N_1780,In_29,In_87);
or U1781 (N_1781,In_426,In_303);
xnor U1782 (N_1782,In_457,In_857);
nand U1783 (N_1783,In_18,In_214);
or U1784 (N_1784,In_761,In_618);
xor U1785 (N_1785,In_145,In_854);
or U1786 (N_1786,In_593,In_213);
xor U1787 (N_1787,In_234,In_357);
nor U1788 (N_1788,In_442,In_391);
xnor U1789 (N_1789,In_757,In_303);
xnor U1790 (N_1790,In_24,In_168);
nand U1791 (N_1791,In_833,In_97);
nor U1792 (N_1792,In_52,In_554);
nand U1793 (N_1793,In_146,In_964);
and U1794 (N_1794,In_189,In_860);
and U1795 (N_1795,In_960,In_649);
nand U1796 (N_1796,In_880,In_766);
nor U1797 (N_1797,In_629,In_602);
nor U1798 (N_1798,In_609,In_18);
and U1799 (N_1799,In_851,In_562);
and U1800 (N_1800,In_390,In_696);
and U1801 (N_1801,In_210,In_388);
or U1802 (N_1802,In_833,In_834);
nor U1803 (N_1803,In_385,In_537);
xor U1804 (N_1804,In_529,In_807);
and U1805 (N_1805,In_849,In_966);
and U1806 (N_1806,In_505,In_511);
xnor U1807 (N_1807,In_280,In_867);
xor U1808 (N_1808,In_531,In_926);
and U1809 (N_1809,In_730,In_719);
and U1810 (N_1810,In_94,In_382);
and U1811 (N_1811,In_396,In_769);
or U1812 (N_1812,In_491,In_258);
and U1813 (N_1813,In_649,In_578);
nor U1814 (N_1814,In_866,In_584);
and U1815 (N_1815,In_980,In_854);
and U1816 (N_1816,In_192,In_89);
xnor U1817 (N_1817,In_500,In_887);
or U1818 (N_1818,In_670,In_106);
nand U1819 (N_1819,In_229,In_207);
nor U1820 (N_1820,In_758,In_439);
xor U1821 (N_1821,In_913,In_166);
nor U1822 (N_1822,In_310,In_235);
nor U1823 (N_1823,In_103,In_687);
xor U1824 (N_1824,In_409,In_318);
and U1825 (N_1825,In_518,In_510);
or U1826 (N_1826,In_781,In_991);
and U1827 (N_1827,In_52,In_302);
nand U1828 (N_1828,In_990,In_328);
nand U1829 (N_1829,In_391,In_380);
nor U1830 (N_1830,In_218,In_972);
xnor U1831 (N_1831,In_596,In_975);
and U1832 (N_1832,In_234,In_575);
nand U1833 (N_1833,In_415,In_781);
and U1834 (N_1834,In_681,In_194);
and U1835 (N_1835,In_733,In_273);
xnor U1836 (N_1836,In_586,In_553);
xor U1837 (N_1837,In_441,In_669);
xor U1838 (N_1838,In_933,In_45);
or U1839 (N_1839,In_436,In_452);
xor U1840 (N_1840,In_945,In_658);
nand U1841 (N_1841,In_838,In_207);
and U1842 (N_1842,In_387,In_237);
nor U1843 (N_1843,In_699,In_249);
or U1844 (N_1844,In_399,In_233);
xnor U1845 (N_1845,In_583,In_548);
nor U1846 (N_1846,In_620,In_610);
xnor U1847 (N_1847,In_320,In_861);
and U1848 (N_1848,In_418,In_591);
xnor U1849 (N_1849,In_813,In_52);
nor U1850 (N_1850,In_421,In_800);
xnor U1851 (N_1851,In_46,In_565);
xnor U1852 (N_1852,In_744,In_776);
or U1853 (N_1853,In_215,In_744);
xnor U1854 (N_1854,In_614,In_497);
and U1855 (N_1855,In_142,In_303);
nor U1856 (N_1856,In_672,In_815);
nor U1857 (N_1857,In_973,In_728);
nand U1858 (N_1858,In_151,In_698);
nand U1859 (N_1859,In_553,In_368);
xnor U1860 (N_1860,In_217,In_501);
and U1861 (N_1861,In_3,In_165);
xnor U1862 (N_1862,In_981,In_249);
xor U1863 (N_1863,In_90,In_886);
or U1864 (N_1864,In_972,In_181);
xnor U1865 (N_1865,In_5,In_31);
and U1866 (N_1866,In_108,In_788);
nand U1867 (N_1867,In_330,In_561);
and U1868 (N_1868,In_583,In_535);
and U1869 (N_1869,In_55,In_291);
nor U1870 (N_1870,In_970,In_709);
nand U1871 (N_1871,In_339,In_551);
xor U1872 (N_1872,In_201,In_797);
or U1873 (N_1873,In_251,In_616);
nand U1874 (N_1874,In_200,In_522);
or U1875 (N_1875,In_41,In_583);
or U1876 (N_1876,In_149,In_474);
nand U1877 (N_1877,In_638,In_98);
and U1878 (N_1878,In_321,In_72);
nor U1879 (N_1879,In_514,In_106);
and U1880 (N_1880,In_814,In_912);
nand U1881 (N_1881,In_129,In_566);
or U1882 (N_1882,In_94,In_644);
xor U1883 (N_1883,In_40,In_399);
nand U1884 (N_1884,In_534,In_194);
and U1885 (N_1885,In_338,In_990);
nor U1886 (N_1886,In_391,In_191);
xnor U1887 (N_1887,In_354,In_250);
nor U1888 (N_1888,In_45,In_761);
or U1889 (N_1889,In_711,In_580);
xnor U1890 (N_1890,In_195,In_136);
and U1891 (N_1891,In_43,In_812);
xor U1892 (N_1892,In_780,In_647);
xnor U1893 (N_1893,In_439,In_801);
nor U1894 (N_1894,In_876,In_106);
xnor U1895 (N_1895,In_461,In_650);
and U1896 (N_1896,In_625,In_199);
nor U1897 (N_1897,In_478,In_3);
nor U1898 (N_1898,In_64,In_4);
nor U1899 (N_1899,In_944,In_38);
nor U1900 (N_1900,In_611,In_22);
nor U1901 (N_1901,In_807,In_498);
nand U1902 (N_1902,In_221,In_8);
or U1903 (N_1903,In_576,In_737);
nor U1904 (N_1904,In_274,In_172);
and U1905 (N_1905,In_106,In_827);
nand U1906 (N_1906,In_346,In_73);
and U1907 (N_1907,In_183,In_824);
nor U1908 (N_1908,In_972,In_691);
xnor U1909 (N_1909,In_514,In_820);
and U1910 (N_1910,In_216,In_841);
nor U1911 (N_1911,In_659,In_668);
nand U1912 (N_1912,In_357,In_436);
xor U1913 (N_1913,In_698,In_941);
nand U1914 (N_1914,In_320,In_881);
nor U1915 (N_1915,In_150,In_26);
nor U1916 (N_1916,In_797,In_451);
or U1917 (N_1917,In_425,In_182);
and U1918 (N_1918,In_311,In_430);
or U1919 (N_1919,In_530,In_284);
nor U1920 (N_1920,In_250,In_447);
and U1921 (N_1921,In_654,In_677);
nand U1922 (N_1922,In_616,In_916);
and U1923 (N_1923,In_115,In_30);
nand U1924 (N_1924,In_994,In_687);
nand U1925 (N_1925,In_717,In_338);
or U1926 (N_1926,In_470,In_21);
xor U1927 (N_1927,In_874,In_560);
or U1928 (N_1928,In_290,In_686);
nor U1929 (N_1929,In_374,In_856);
and U1930 (N_1930,In_78,In_372);
nor U1931 (N_1931,In_839,In_180);
or U1932 (N_1932,In_487,In_178);
and U1933 (N_1933,In_358,In_520);
and U1934 (N_1934,In_956,In_961);
xor U1935 (N_1935,In_647,In_266);
xor U1936 (N_1936,In_586,In_251);
and U1937 (N_1937,In_114,In_170);
and U1938 (N_1938,In_448,In_943);
or U1939 (N_1939,In_190,In_514);
nor U1940 (N_1940,In_791,In_682);
or U1941 (N_1941,In_98,In_276);
and U1942 (N_1942,In_142,In_810);
nand U1943 (N_1943,In_22,In_949);
and U1944 (N_1944,In_976,In_787);
nor U1945 (N_1945,In_861,In_789);
or U1946 (N_1946,In_478,In_494);
or U1947 (N_1947,In_706,In_802);
nor U1948 (N_1948,In_833,In_310);
and U1949 (N_1949,In_61,In_319);
or U1950 (N_1950,In_67,In_421);
xor U1951 (N_1951,In_932,In_655);
xnor U1952 (N_1952,In_100,In_71);
xnor U1953 (N_1953,In_434,In_596);
or U1954 (N_1954,In_274,In_802);
and U1955 (N_1955,In_625,In_417);
and U1956 (N_1956,In_239,In_436);
xnor U1957 (N_1957,In_774,In_827);
and U1958 (N_1958,In_890,In_140);
nand U1959 (N_1959,In_592,In_654);
or U1960 (N_1960,In_996,In_958);
nor U1961 (N_1961,In_250,In_695);
nand U1962 (N_1962,In_921,In_910);
nand U1963 (N_1963,In_308,In_807);
nand U1964 (N_1964,In_57,In_108);
and U1965 (N_1965,In_861,In_898);
nor U1966 (N_1966,In_164,In_986);
or U1967 (N_1967,In_142,In_155);
nand U1968 (N_1968,In_180,In_10);
xor U1969 (N_1969,In_58,In_773);
nand U1970 (N_1970,In_526,In_910);
nor U1971 (N_1971,In_770,In_583);
nor U1972 (N_1972,In_973,In_591);
nand U1973 (N_1973,In_275,In_192);
xnor U1974 (N_1974,In_425,In_200);
or U1975 (N_1975,In_823,In_844);
xor U1976 (N_1976,In_75,In_960);
or U1977 (N_1977,In_64,In_324);
nor U1978 (N_1978,In_661,In_468);
nor U1979 (N_1979,In_20,In_840);
nand U1980 (N_1980,In_813,In_74);
xor U1981 (N_1981,In_534,In_288);
and U1982 (N_1982,In_888,In_650);
and U1983 (N_1983,In_217,In_312);
and U1984 (N_1984,In_210,In_480);
or U1985 (N_1985,In_149,In_8);
nand U1986 (N_1986,In_467,In_676);
and U1987 (N_1987,In_994,In_356);
nand U1988 (N_1988,In_63,In_393);
and U1989 (N_1989,In_365,In_528);
xor U1990 (N_1990,In_276,In_139);
xor U1991 (N_1991,In_147,In_447);
or U1992 (N_1992,In_607,In_965);
and U1993 (N_1993,In_652,In_135);
xor U1994 (N_1994,In_324,In_383);
and U1995 (N_1995,In_211,In_455);
nand U1996 (N_1996,In_311,In_499);
or U1997 (N_1997,In_765,In_200);
nor U1998 (N_1998,In_985,In_424);
nor U1999 (N_1999,In_163,In_37);
or U2000 (N_2000,In_784,In_612);
nand U2001 (N_2001,In_93,In_774);
nand U2002 (N_2002,In_720,In_647);
nor U2003 (N_2003,In_11,In_603);
and U2004 (N_2004,In_585,In_707);
nor U2005 (N_2005,In_427,In_181);
and U2006 (N_2006,In_688,In_372);
and U2007 (N_2007,In_391,In_757);
xnor U2008 (N_2008,In_88,In_929);
nor U2009 (N_2009,In_700,In_526);
xor U2010 (N_2010,In_980,In_906);
or U2011 (N_2011,In_688,In_620);
nand U2012 (N_2012,In_337,In_887);
xnor U2013 (N_2013,In_956,In_341);
and U2014 (N_2014,In_374,In_883);
and U2015 (N_2015,In_14,In_841);
nand U2016 (N_2016,In_205,In_35);
xnor U2017 (N_2017,In_56,In_989);
or U2018 (N_2018,In_55,In_752);
or U2019 (N_2019,In_381,In_282);
xnor U2020 (N_2020,In_238,In_711);
nand U2021 (N_2021,In_531,In_812);
xor U2022 (N_2022,In_230,In_409);
or U2023 (N_2023,In_279,In_33);
nor U2024 (N_2024,In_452,In_752);
and U2025 (N_2025,In_761,In_231);
xor U2026 (N_2026,In_738,In_618);
xor U2027 (N_2027,In_593,In_625);
nor U2028 (N_2028,In_702,In_531);
nand U2029 (N_2029,In_219,In_153);
or U2030 (N_2030,In_214,In_750);
and U2031 (N_2031,In_646,In_33);
xor U2032 (N_2032,In_12,In_773);
nor U2033 (N_2033,In_356,In_341);
nor U2034 (N_2034,In_224,In_844);
and U2035 (N_2035,In_56,In_412);
nand U2036 (N_2036,In_146,In_562);
nand U2037 (N_2037,In_445,In_130);
nand U2038 (N_2038,In_293,In_739);
or U2039 (N_2039,In_2,In_48);
or U2040 (N_2040,In_746,In_470);
xor U2041 (N_2041,In_805,In_457);
and U2042 (N_2042,In_964,In_223);
nand U2043 (N_2043,In_492,In_812);
and U2044 (N_2044,In_429,In_500);
nor U2045 (N_2045,In_34,In_167);
and U2046 (N_2046,In_670,In_579);
xnor U2047 (N_2047,In_850,In_62);
and U2048 (N_2048,In_179,In_974);
xnor U2049 (N_2049,In_838,In_754);
xor U2050 (N_2050,In_400,In_204);
and U2051 (N_2051,In_778,In_884);
xor U2052 (N_2052,In_78,In_869);
or U2053 (N_2053,In_593,In_973);
xnor U2054 (N_2054,In_284,In_256);
and U2055 (N_2055,In_484,In_76);
or U2056 (N_2056,In_82,In_719);
nor U2057 (N_2057,In_230,In_534);
nand U2058 (N_2058,In_768,In_76);
nor U2059 (N_2059,In_51,In_13);
nor U2060 (N_2060,In_619,In_45);
nor U2061 (N_2061,In_557,In_691);
xor U2062 (N_2062,In_739,In_912);
xor U2063 (N_2063,In_392,In_236);
or U2064 (N_2064,In_393,In_256);
nor U2065 (N_2065,In_426,In_82);
xnor U2066 (N_2066,In_166,In_733);
nor U2067 (N_2067,In_304,In_787);
nand U2068 (N_2068,In_864,In_429);
nor U2069 (N_2069,In_464,In_275);
nor U2070 (N_2070,In_33,In_228);
xnor U2071 (N_2071,In_409,In_882);
nor U2072 (N_2072,In_963,In_946);
nor U2073 (N_2073,In_708,In_957);
nand U2074 (N_2074,In_302,In_740);
nand U2075 (N_2075,In_857,In_380);
xor U2076 (N_2076,In_299,In_807);
or U2077 (N_2077,In_122,In_833);
xnor U2078 (N_2078,In_834,In_706);
xor U2079 (N_2079,In_204,In_380);
xor U2080 (N_2080,In_800,In_906);
nor U2081 (N_2081,In_162,In_153);
nand U2082 (N_2082,In_634,In_901);
or U2083 (N_2083,In_169,In_175);
nand U2084 (N_2084,In_795,In_359);
nand U2085 (N_2085,In_660,In_33);
nor U2086 (N_2086,In_216,In_127);
nor U2087 (N_2087,In_73,In_282);
and U2088 (N_2088,In_459,In_620);
nand U2089 (N_2089,In_93,In_84);
or U2090 (N_2090,In_54,In_274);
and U2091 (N_2091,In_555,In_642);
xor U2092 (N_2092,In_274,In_732);
and U2093 (N_2093,In_230,In_286);
xor U2094 (N_2094,In_550,In_105);
nor U2095 (N_2095,In_999,In_192);
or U2096 (N_2096,In_122,In_767);
nor U2097 (N_2097,In_201,In_871);
nand U2098 (N_2098,In_163,In_798);
and U2099 (N_2099,In_116,In_159);
xor U2100 (N_2100,In_610,In_374);
nor U2101 (N_2101,In_942,In_903);
xnor U2102 (N_2102,In_732,In_52);
nor U2103 (N_2103,In_794,In_677);
and U2104 (N_2104,In_626,In_365);
nor U2105 (N_2105,In_964,In_661);
nand U2106 (N_2106,In_148,In_842);
or U2107 (N_2107,In_154,In_814);
or U2108 (N_2108,In_283,In_188);
and U2109 (N_2109,In_225,In_403);
and U2110 (N_2110,In_786,In_301);
and U2111 (N_2111,In_97,In_946);
and U2112 (N_2112,In_424,In_927);
nor U2113 (N_2113,In_960,In_269);
and U2114 (N_2114,In_452,In_468);
nor U2115 (N_2115,In_193,In_989);
and U2116 (N_2116,In_443,In_147);
xnor U2117 (N_2117,In_438,In_185);
nand U2118 (N_2118,In_747,In_957);
and U2119 (N_2119,In_324,In_609);
xor U2120 (N_2120,In_297,In_967);
xor U2121 (N_2121,In_481,In_306);
xor U2122 (N_2122,In_306,In_372);
xnor U2123 (N_2123,In_457,In_700);
and U2124 (N_2124,In_308,In_85);
or U2125 (N_2125,In_470,In_377);
or U2126 (N_2126,In_959,In_356);
nor U2127 (N_2127,In_269,In_701);
or U2128 (N_2128,In_962,In_573);
or U2129 (N_2129,In_427,In_685);
nand U2130 (N_2130,In_874,In_796);
xnor U2131 (N_2131,In_352,In_125);
nor U2132 (N_2132,In_60,In_28);
and U2133 (N_2133,In_134,In_557);
nor U2134 (N_2134,In_860,In_387);
xnor U2135 (N_2135,In_96,In_307);
or U2136 (N_2136,In_634,In_879);
xor U2137 (N_2137,In_142,In_510);
or U2138 (N_2138,In_403,In_619);
nand U2139 (N_2139,In_69,In_226);
or U2140 (N_2140,In_15,In_149);
xnor U2141 (N_2141,In_76,In_204);
nor U2142 (N_2142,In_927,In_246);
or U2143 (N_2143,In_516,In_337);
or U2144 (N_2144,In_956,In_181);
and U2145 (N_2145,In_136,In_989);
nand U2146 (N_2146,In_510,In_153);
and U2147 (N_2147,In_296,In_300);
nand U2148 (N_2148,In_935,In_713);
nor U2149 (N_2149,In_845,In_928);
xor U2150 (N_2150,In_677,In_376);
and U2151 (N_2151,In_525,In_171);
or U2152 (N_2152,In_673,In_922);
or U2153 (N_2153,In_435,In_303);
nor U2154 (N_2154,In_244,In_528);
or U2155 (N_2155,In_310,In_706);
xnor U2156 (N_2156,In_866,In_512);
nor U2157 (N_2157,In_17,In_893);
or U2158 (N_2158,In_996,In_95);
or U2159 (N_2159,In_168,In_571);
nand U2160 (N_2160,In_681,In_81);
nor U2161 (N_2161,In_938,In_986);
xnor U2162 (N_2162,In_140,In_888);
xor U2163 (N_2163,In_73,In_362);
nand U2164 (N_2164,In_916,In_867);
or U2165 (N_2165,In_728,In_138);
or U2166 (N_2166,In_298,In_222);
nand U2167 (N_2167,In_295,In_603);
or U2168 (N_2168,In_559,In_551);
and U2169 (N_2169,In_119,In_452);
or U2170 (N_2170,In_952,In_725);
nor U2171 (N_2171,In_253,In_257);
nand U2172 (N_2172,In_365,In_75);
xnor U2173 (N_2173,In_314,In_814);
or U2174 (N_2174,In_708,In_802);
and U2175 (N_2175,In_687,In_616);
nand U2176 (N_2176,In_864,In_109);
and U2177 (N_2177,In_314,In_725);
and U2178 (N_2178,In_507,In_96);
or U2179 (N_2179,In_874,In_371);
xor U2180 (N_2180,In_465,In_903);
xnor U2181 (N_2181,In_365,In_683);
and U2182 (N_2182,In_759,In_28);
nand U2183 (N_2183,In_522,In_800);
nand U2184 (N_2184,In_384,In_449);
xnor U2185 (N_2185,In_530,In_246);
or U2186 (N_2186,In_983,In_969);
nand U2187 (N_2187,In_7,In_987);
or U2188 (N_2188,In_532,In_713);
nand U2189 (N_2189,In_57,In_324);
nand U2190 (N_2190,In_745,In_822);
nor U2191 (N_2191,In_971,In_372);
xnor U2192 (N_2192,In_831,In_443);
or U2193 (N_2193,In_817,In_467);
xor U2194 (N_2194,In_929,In_452);
nand U2195 (N_2195,In_277,In_971);
xor U2196 (N_2196,In_583,In_115);
or U2197 (N_2197,In_450,In_805);
nand U2198 (N_2198,In_863,In_853);
xnor U2199 (N_2199,In_460,In_164);
xor U2200 (N_2200,In_624,In_185);
and U2201 (N_2201,In_403,In_732);
xor U2202 (N_2202,In_172,In_305);
nand U2203 (N_2203,In_312,In_286);
xor U2204 (N_2204,In_447,In_931);
or U2205 (N_2205,In_372,In_123);
and U2206 (N_2206,In_780,In_637);
and U2207 (N_2207,In_456,In_203);
or U2208 (N_2208,In_339,In_200);
and U2209 (N_2209,In_534,In_996);
nand U2210 (N_2210,In_606,In_782);
nand U2211 (N_2211,In_612,In_810);
nand U2212 (N_2212,In_172,In_309);
xor U2213 (N_2213,In_951,In_777);
nor U2214 (N_2214,In_437,In_783);
and U2215 (N_2215,In_937,In_83);
nand U2216 (N_2216,In_523,In_909);
xnor U2217 (N_2217,In_552,In_147);
or U2218 (N_2218,In_152,In_862);
nand U2219 (N_2219,In_779,In_3);
nand U2220 (N_2220,In_641,In_980);
and U2221 (N_2221,In_592,In_25);
and U2222 (N_2222,In_107,In_933);
or U2223 (N_2223,In_542,In_623);
nor U2224 (N_2224,In_741,In_667);
nor U2225 (N_2225,In_729,In_821);
xor U2226 (N_2226,In_740,In_30);
nand U2227 (N_2227,In_280,In_749);
xnor U2228 (N_2228,In_874,In_576);
nor U2229 (N_2229,In_156,In_103);
and U2230 (N_2230,In_518,In_960);
or U2231 (N_2231,In_670,In_974);
or U2232 (N_2232,In_475,In_212);
nor U2233 (N_2233,In_921,In_544);
and U2234 (N_2234,In_803,In_208);
nand U2235 (N_2235,In_484,In_842);
nor U2236 (N_2236,In_757,In_67);
or U2237 (N_2237,In_610,In_239);
xor U2238 (N_2238,In_680,In_979);
nor U2239 (N_2239,In_958,In_163);
xnor U2240 (N_2240,In_691,In_244);
nand U2241 (N_2241,In_587,In_650);
nand U2242 (N_2242,In_525,In_574);
xnor U2243 (N_2243,In_920,In_814);
and U2244 (N_2244,In_69,In_905);
xnor U2245 (N_2245,In_667,In_110);
and U2246 (N_2246,In_819,In_9);
xor U2247 (N_2247,In_472,In_147);
nand U2248 (N_2248,In_544,In_794);
xnor U2249 (N_2249,In_375,In_861);
xor U2250 (N_2250,In_478,In_163);
nand U2251 (N_2251,In_24,In_369);
nor U2252 (N_2252,In_774,In_560);
and U2253 (N_2253,In_576,In_239);
or U2254 (N_2254,In_607,In_431);
or U2255 (N_2255,In_969,In_106);
xnor U2256 (N_2256,In_685,In_294);
and U2257 (N_2257,In_245,In_305);
nor U2258 (N_2258,In_420,In_509);
and U2259 (N_2259,In_74,In_991);
xor U2260 (N_2260,In_376,In_572);
nand U2261 (N_2261,In_186,In_777);
and U2262 (N_2262,In_97,In_587);
nor U2263 (N_2263,In_137,In_177);
nand U2264 (N_2264,In_782,In_342);
or U2265 (N_2265,In_283,In_860);
nor U2266 (N_2266,In_783,In_105);
nand U2267 (N_2267,In_131,In_431);
nor U2268 (N_2268,In_518,In_942);
or U2269 (N_2269,In_799,In_61);
or U2270 (N_2270,In_883,In_938);
or U2271 (N_2271,In_357,In_755);
xnor U2272 (N_2272,In_174,In_86);
and U2273 (N_2273,In_784,In_547);
nor U2274 (N_2274,In_591,In_842);
nand U2275 (N_2275,In_553,In_361);
nand U2276 (N_2276,In_26,In_658);
nand U2277 (N_2277,In_204,In_544);
xor U2278 (N_2278,In_314,In_243);
and U2279 (N_2279,In_308,In_723);
nor U2280 (N_2280,In_562,In_819);
nand U2281 (N_2281,In_612,In_285);
xnor U2282 (N_2282,In_234,In_9);
nand U2283 (N_2283,In_93,In_426);
or U2284 (N_2284,In_268,In_578);
and U2285 (N_2285,In_520,In_972);
or U2286 (N_2286,In_579,In_495);
xnor U2287 (N_2287,In_274,In_676);
xor U2288 (N_2288,In_188,In_814);
xor U2289 (N_2289,In_508,In_132);
nand U2290 (N_2290,In_739,In_188);
nor U2291 (N_2291,In_750,In_905);
or U2292 (N_2292,In_718,In_391);
xor U2293 (N_2293,In_855,In_114);
nor U2294 (N_2294,In_976,In_456);
nor U2295 (N_2295,In_13,In_103);
xor U2296 (N_2296,In_703,In_239);
or U2297 (N_2297,In_85,In_642);
nor U2298 (N_2298,In_801,In_218);
nand U2299 (N_2299,In_115,In_402);
nor U2300 (N_2300,In_749,In_718);
or U2301 (N_2301,In_697,In_968);
or U2302 (N_2302,In_266,In_41);
and U2303 (N_2303,In_815,In_933);
and U2304 (N_2304,In_730,In_534);
or U2305 (N_2305,In_633,In_680);
or U2306 (N_2306,In_691,In_525);
xor U2307 (N_2307,In_722,In_811);
nand U2308 (N_2308,In_735,In_354);
nor U2309 (N_2309,In_704,In_493);
xor U2310 (N_2310,In_886,In_479);
and U2311 (N_2311,In_606,In_39);
nor U2312 (N_2312,In_621,In_179);
or U2313 (N_2313,In_258,In_932);
or U2314 (N_2314,In_336,In_949);
and U2315 (N_2315,In_163,In_314);
nor U2316 (N_2316,In_384,In_846);
xor U2317 (N_2317,In_812,In_721);
xor U2318 (N_2318,In_113,In_873);
xnor U2319 (N_2319,In_76,In_991);
or U2320 (N_2320,In_883,In_792);
and U2321 (N_2321,In_983,In_590);
or U2322 (N_2322,In_157,In_849);
xor U2323 (N_2323,In_292,In_401);
or U2324 (N_2324,In_707,In_94);
nor U2325 (N_2325,In_746,In_800);
xor U2326 (N_2326,In_68,In_974);
nand U2327 (N_2327,In_541,In_903);
nor U2328 (N_2328,In_151,In_287);
xnor U2329 (N_2329,In_227,In_786);
or U2330 (N_2330,In_365,In_975);
or U2331 (N_2331,In_825,In_31);
nand U2332 (N_2332,In_242,In_273);
and U2333 (N_2333,In_589,In_398);
xor U2334 (N_2334,In_681,In_554);
nor U2335 (N_2335,In_428,In_372);
nand U2336 (N_2336,In_194,In_211);
and U2337 (N_2337,In_627,In_898);
and U2338 (N_2338,In_34,In_125);
nor U2339 (N_2339,In_83,In_790);
or U2340 (N_2340,In_275,In_895);
xor U2341 (N_2341,In_95,In_130);
and U2342 (N_2342,In_478,In_180);
xor U2343 (N_2343,In_37,In_32);
or U2344 (N_2344,In_99,In_832);
xor U2345 (N_2345,In_54,In_227);
nand U2346 (N_2346,In_983,In_888);
and U2347 (N_2347,In_864,In_443);
nor U2348 (N_2348,In_476,In_808);
xnor U2349 (N_2349,In_749,In_994);
and U2350 (N_2350,In_215,In_98);
xor U2351 (N_2351,In_129,In_720);
or U2352 (N_2352,In_233,In_611);
and U2353 (N_2353,In_945,In_712);
and U2354 (N_2354,In_560,In_542);
nor U2355 (N_2355,In_774,In_910);
nand U2356 (N_2356,In_976,In_136);
nand U2357 (N_2357,In_626,In_952);
and U2358 (N_2358,In_8,In_53);
nand U2359 (N_2359,In_358,In_894);
nor U2360 (N_2360,In_687,In_495);
nor U2361 (N_2361,In_190,In_624);
and U2362 (N_2362,In_683,In_100);
and U2363 (N_2363,In_10,In_696);
and U2364 (N_2364,In_933,In_240);
nor U2365 (N_2365,In_635,In_81);
or U2366 (N_2366,In_750,In_632);
nor U2367 (N_2367,In_944,In_946);
and U2368 (N_2368,In_103,In_664);
and U2369 (N_2369,In_259,In_477);
or U2370 (N_2370,In_939,In_138);
nand U2371 (N_2371,In_22,In_206);
or U2372 (N_2372,In_276,In_691);
nand U2373 (N_2373,In_950,In_33);
nand U2374 (N_2374,In_149,In_270);
nand U2375 (N_2375,In_893,In_139);
nand U2376 (N_2376,In_647,In_940);
nor U2377 (N_2377,In_683,In_975);
nand U2378 (N_2378,In_875,In_378);
xnor U2379 (N_2379,In_977,In_573);
or U2380 (N_2380,In_960,In_128);
nor U2381 (N_2381,In_989,In_858);
nand U2382 (N_2382,In_189,In_631);
nand U2383 (N_2383,In_324,In_959);
nor U2384 (N_2384,In_827,In_424);
nand U2385 (N_2385,In_989,In_896);
or U2386 (N_2386,In_470,In_277);
and U2387 (N_2387,In_228,In_951);
or U2388 (N_2388,In_426,In_601);
or U2389 (N_2389,In_464,In_659);
xnor U2390 (N_2390,In_547,In_903);
xor U2391 (N_2391,In_289,In_410);
or U2392 (N_2392,In_371,In_747);
nor U2393 (N_2393,In_453,In_484);
or U2394 (N_2394,In_151,In_515);
and U2395 (N_2395,In_654,In_265);
and U2396 (N_2396,In_944,In_61);
and U2397 (N_2397,In_635,In_22);
and U2398 (N_2398,In_1,In_13);
nand U2399 (N_2399,In_928,In_509);
xnor U2400 (N_2400,In_557,In_296);
xor U2401 (N_2401,In_222,In_731);
nor U2402 (N_2402,In_110,In_436);
nand U2403 (N_2403,In_856,In_555);
or U2404 (N_2404,In_511,In_287);
xnor U2405 (N_2405,In_868,In_699);
nor U2406 (N_2406,In_299,In_444);
xnor U2407 (N_2407,In_654,In_850);
and U2408 (N_2408,In_961,In_777);
or U2409 (N_2409,In_989,In_80);
xnor U2410 (N_2410,In_237,In_336);
nor U2411 (N_2411,In_343,In_290);
and U2412 (N_2412,In_3,In_416);
or U2413 (N_2413,In_935,In_190);
nor U2414 (N_2414,In_487,In_513);
and U2415 (N_2415,In_606,In_258);
nor U2416 (N_2416,In_885,In_586);
and U2417 (N_2417,In_455,In_780);
and U2418 (N_2418,In_642,In_763);
nor U2419 (N_2419,In_127,In_806);
and U2420 (N_2420,In_638,In_301);
and U2421 (N_2421,In_667,In_21);
xor U2422 (N_2422,In_436,In_174);
xnor U2423 (N_2423,In_316,In_478);
nand U2424 (N_2424,In_991,In_690);
nor U2425 (N_2425,In_928,In_848);
nor U2426 (N_2426,In_220,In_375);
and U2427 (N_2427,In_886,In_663);
xnor U2428 (N_2428,In_439,In_351);
and U2429 (N_2429,In_340,In_730);
and U2430 (N_2430,In_569,In_244);
nor U2431 (N_2431,In_962,In_381);
nand U2432 (N_2432,In_435,In_122);
or U2433 (N_2433,In_444,In_926);
or U2434 (N_2434,In_398,In_517);
nor U2435 (N_2435,In_899,In_284);
xnor U2436 (N_2436,In_744,In_704);
nand U2437 (N_2437,In_952,In_413);
xnor U2438 (N_2438,In_480,In_968);
nor U2439 (N_2439,In_868,In_725);
or U2440 (N_2440,In_971,In_299);
nand U2441 (N_2441,In_326,In_822);
nor U2442 (N_2442,In_30,In_691);
nand U2443 (N_2443,In_785,In_881);
nand U2444 (N_2444,In_653,In_492);
and U2445 (N_2445,In_598,In_548);
and U2446 (N_2446,In_703,In_982);
xor U2447 (N_2447,In_615,In_457);
or U2448 (N_2448,In_308,In_824);
and U2449 (N_2449,In_512,In_949);
nor U2450 (N_2450,In_222,In_391);
and U2451 (N_2451,In_840,In_24);
and U2452 (N_2452,In_883,In_647);
nand U2453 (N_2453,In_609,In_893);
nor U2454 (N_2454,In_747,In_443);
nand U2455 (N_2455,In_679,In_813);
nand U2456 (N_2456,In_864,In_710);
or U2457 (N_2457,In_132,In_854);
nor U2458 (N_2458,In_506,In_398);
nand U2459 (N_2459,In_595,In_70);
nand U2460 (N_2460,In_931,In_286);
and U2461 (N_2461,In_761,In_214);
or U2462 (N_2462,In_960,In_617);
nand U2463 (N_2463,In_189,In_386);
xnor U2464 (N_2464,In_645,In_223);
xor U2465 (N_2465,In_463,In_154);
xor U2466 (N_2466,In_290,In_80);
or U2467 (N_2467,In_355,In_245);
and U2468 (N_2468,In_374,In_882);
nor U2469 (N_2469,In_937,In_966);
xnor U2470 (N_2470,In_213,In_966);
or U2471 (N_2471,In_590,In_664);
nand U2472 (N_2472,In_846,In_989);
xor U2473 (N_2473,In_889,In_832);
xnor U2474 (N_2474,In_899,In_830);
nor U2475 (N_2475,In_161,In_31);
nand U2476 (N_2476,In_469,In_389);
and U2477 (N_2477,In_201,In_367);
nand U2478 (N_2478,In_778,In_702);
and U2479 (N_2479,In_654,In_264);
nor U2480 (N_2480,In_348,In_351);
nand U2481 (N_2481,In_942,In_415);
or U2482 (N_2482,In_471,In_609);
or U2483 (N_2483,In_346,In_786);
and U2484 (N_2484,In_505,In_746);
or U2485 (N_2485,In_226,In_668);
nand U2486 (N_2486,In_40,In_561);
nor U2487 (N_2487,In_217,In_476);
or U2488 (N_2488,In_163,In_290);
nand U2489 (N_2489,In_448,In_363);
and U2490 (N_2490,In_197,In_517);
xnor U2491 (N_2491,In_879,In_492);
and U2492 (N_2492,In_422,In_950);
xor U2493 (N_2493,In_523,In_831);
xnor U2494 (N_2494,In_878,In_213);
or U2495 (N_2495,In_987,In_907);
xor U2496 (N_2496,In_684,In_648);
nand U2497 (N_2497,In_998,In_828);
nand U2498 (N_2498,In_557,In_829);
xor U2499 (N_2499,In_644,In_704);
xor U2500 (N_2500,In_53,In_716);
nand U2501 (N_2501,In_216,In_437);
or U2502 (N_2502,In_347,In_306);
nand U2503 (N_2503,In_599,In_20);
nor U2504 (N_2504,In_70,In_273);
or U2505 (N_2505,In_893,In_861);
nor U2506 (N_2506,In_704,In_243);
or U2507 (N_2507,In_834,In_120);
xor U2508 (N_2508,In_27,In_624);
xnor U2509 (N_2509,In_410,In_968);
or U2510 (N_2510,In_568,In_43);
and U2511 (N_2511,In_307,In_714);
nor U2512 (N_2512,In_93,In_397);
nor U2513 (N_2513,In_217,In_393);
nand U2514 (N_2514,In_316,In_743);
or U2515 (N_2515,In_825,In_872);
nand U2516 (N_2516,In_942,In_55);
xnor U2517 (N_2517,In_256,In_268);
nor U2518 (N_2518,In_817,In_602);
or U2519 (N_2519,In_708,In_85);
nand U2520 (N_2520,In_49,In_672);
and U2521 (N_2521,In_197,In_501);
xor U2522 (N_2522,In_829,In_510);
and U2523 (N_2523,In_768,In_941);
nor U2524 (N_2524,In_671,In_483);
or U2525 (N_2525,In_554,In_621);
or U2526 (N_2526,In_57,In_831);
nor U2527 (N_2527,In_301,In_39);
and U2528 (N_2528,In_401,In_74);
nor U2529 (N_2529,In_235,In_74);
and U2530 (N_2530,In_447,In_469);
xor U2531 (N_2531,In_364,In_127);
and U2532 (N_2532,In_295,In_803);
and U2533 (N_2533,In_6,In_83);
xor U2534 (N_2534,In_613,In_100);
and U2535 (N_2535,In_441,In_656);
or U2536 (N_2536,In_373,In_483);
nor U2537 (N_2537,In_247,In_924);
nor U2538 (N_2538,In_894,In_895);
xor U2539 (N_2539,In_91,In_292);
nand U2540 (N_2540,In_601,In_450);
or U2541 (N_2541,In_167,In_752);
nor U2542 (N_2542,In_193,In_765);
xor U2543 (N_2543,In_185,In_414);
nor U2544 (N_2544,In_827,In_205);
xnor U2545 (N_2545,In_25,In_875);
xor U2546 (N_2546,In_573,In_213);
and U2547 (N_2547,In_577,In_717);
xnor U2548 (N_2548,In_784,In_967);
and U2549 (N_2549,In_522,In_509);
and U2550 (N_2550,In_220,In_778);
and U2551 (N_2551,In_590,In_997);
or U2552 (N_2552,In_794,In_359);
xnor U2553 (N_2553,In_126,In_165);
or U2554 (N_2554,In_836,In_143);
or U2555 (N_2555,In_664,In_983);
xor U2556 (N_2556,In_58,In_176);
and U2557 (N_2557,In_333,In_516);
xor U2558 (N_2558,In_79,In_26);
or U2559 (N_2559,In_496,In_165);
and U2560 (N_2560,In_737,In_649);
or U2561 (N_2561,In_346,In_154);
nor U2562 (N_2562,In_939,In_629);
nor U2563 (N_2563,In_690,In_907);
nand U2564 (N_2564,In_325,In_45);
nor U2565 (N_2565,In_870,In_62);
xor U2566 (N_2566,In_13,In_368);
and U2567 (N_2567,In_711,In_551);
nor U2568 (N_2568,In_220,In_460);
and U2569 (N_2569,In_283,In_524);
nor U2570 (N_2570,In_291,In_979);
xor U2571 (N_2571,In_887,In_418);
nand U2572 (N_2572,In_17,In_342);
and U2573 (N_2573,In_744,In_333);
xnor U2574 (N_2574,In_146,In_837);
xor U2575 (N_2575,In_489,In_856);
and U2576 (N_2576,In_941,In_246);
xnor U2577 (N_2577,In_522,In_344);
or U2578 (N_2578,In_343,In_970);
nor U2579 (N_2579,In_606,In_170);
xor U2580 (N_2580,In_615,In_745);
or U2581 (N_2581,In_671,In_811);
or U2582 (N_2582,In_659,In_388);
or U2583 (N_2583,In_484,In_607);
and U2584 (N_2584,In_825,In_115);
nor U2585 (N_2585,In_991,In_613);
nor U2586 (N_2586,In_247,In_746);
nand U2587 (N_2587,In_845,In_795);
or U2588 (N_2588,In_680,In_910);
and U2589 (N_2589,In_728,In_407);
or U2590 (N_2590,In_793,In_546);
nand U2591 (N_2591,In_809,In_2);
and U2592 (N_2592,In_497,In_355);
or U2593 (N_2593,In_958,In_465);
nor U2594 (N_2594,In_848,In_304);
nand U2595 (N_2595,In_130,In_137);
xor U2596 (N_2596,In_25,In_928);
nand U2597 (N_2597,In_100,In_451);
and U2598 (N_2598,In_437,In_384);
or U2599 (N_2599,In_647,In_375);
xor U2600 (N_2600,In_29,In_833);
nand U2601 (N_2601,In_939,In_837);
xor U2602 (N_2602,In_731,In_254);
and U2603 (N_2603,In_332,In_874);
nand U2604 (N_2604,In_731,In_207);
and U2605 (N_2605,In_764,In_312);
nor U2606 (N_2606,In_613,In_620);
or U2607 (N_2607,In_765,In_15);
and U2608 (N_2608,In_882,In_441);
and U2609 (N_2609,In_876,In_217);
and U2610 (N_2610,In_545,In_460);
and U2611 (N_2611,In_265,In_560);
nand U2612 (N_2612,In_349,In_531);
and U2613 (N_2613,In_392,In_33);
nor U2614 (N_2614,In_507,In_929);
nor U2615 (N_2615,In_590,In_982);
xnor U2616 (N_2616,In_220,In_447);
nor U2617 (N_2617,In_95,In_481);
nor U2618 (N_2618,In_490,In_775);
and U2619 (N_2619,In_367,In_119);
and U2620 (N_2620,In_110,In_333);
xnor U2621 (N_2621,In_311,In_617);
and U2622 (N_2622,In_243,In_215);
and U2623 (N_2623,In_116,In_285);
and U2624 (N_2624,In_743,In_381);
nor U2625 (N_2625,In_202,In_937);
nand U2626 (N_2626,In_411,In_16);
or U2627 (N_2627,In_518,In_530);
xnor U2628 (N_2628,In_624,In_713);
or U2629 (N_2629,In_3,In_423);
nand U2630 (N_2630,In_352,In_982);
nor U2631 (N_2631,In_385,In_757);
or U2632 (N_2632,In_267,In_325);
and U2633 (N_2633,In_829,In_959);
xor U2634 (N_2634,In_495,In_211);
nor U2635 (N_2635,In_113,In_108);
xnor U2636 (N_2636,In_848,In_781);
xor U2637 (N_2637,In_85,In_212);
nand U2638 (N_2638,In_355,In_552);
nor U2639 (N_2639,In_157,In_274);
nor U2640 (N_2640,In_299,In_579);
xnor U2641 (N_2641,In_1,In_768);
or U2642 (N_2642,In_931,In_540);
nand U2643 (N_2643,In_26,In_577);
and U2644 (N_2644,In_889,In_890);
or U2645 (N_2645,In_50,In_862);
or U2646 (N_2646,In_893,In_878);
and U2647 (N_2647,In_758,In_118);
and U2648 (N_2648,In_950,In_481);
nor U2649 (N_2649,In_50,In_415);
or U2650 (N_2650,In_239,In_786);
and U2651 (N_2651,In_842,In_860);
or U2652 (N_2652,In_121,In_552);
nor U2653 (N_2653,In_228,In_718);
nand U2654 (N_2654,In_366,In_845);
and U2655 (N_2655,In_303,In_367);
and U2656 (N_2656,In_158,In_381);
and U2657 (N_2657,In_780,In_199);
nand U2658 (N_2658,In_363,In_259);
nor U2659 (N_2659,In_9,In_128);
and U2660 (N_2660,In_379,In_622);
nand U2661 (N_2661,In_439,In_12);
xnor U2662 (N_2662,In_584,In_900);
nand U2663 (N_2663,In_164,In_531);
xnor U2664 (N_2664,In_475,In_592);
nor U2665 (N_2665,In_65,In_773);
or U2666 (N_2666,In_516,In_196);
nor U2667 (N_2667,In_525,In_429);
nor U2668 (N_2668,In_789,In_340);
and U2669 (N_2669,In_677,In_567);
or U2670 (N_2670,In_728,In_26);
and U2671 (N_2671,In_651,In_125);
and U2672 (N_2672,In_220,In_328);
nor U2673 (N_2673,In_824,In_727);
xor U2674 (N_2674,In_250,In_314);
nor U2675 (N_2675,In_590,In_311);
or U2676 (N_2676,In_469,In_767);
nor U2677 (N_2677,In_895,In_241);
nand U2678 (N_2678,In_970,In_260);
and U2679 (N_2679,In_644,In_563);
nand U2680 (N_2680,In_205,In_347);
nor U2681 (N_2681,In_19,In_474);
nand U2682 (N_2682,In_303,In_744);
xnor U2683 (N_2683,In_959,In_739);
xnor U2684 (N_2684,In_582,In_631);
or U2685 (N_2685,In_325,In_844);
or U2686 (N_2686,In_252,In_413);
nand U2687 (N_2687,In_779,In_508);
and U2688 (N_2688,In_283,In_265);
xor U2689 (N_2689,In_143,In_464);
nor U2690 (N_2690,In_687,In_988);
and U2691 (N_2691,In_805,In_568);
nor U2692 (N_2692,In_136,In_425);
or U2693 (N_2693,In_422,In_541);
xor U2694 (N_2694,In_817,In_540);
nand U2695 (N_2695,In_580,In_8);
xnor U2696 (N_2696,In_88,In_689);
xnor U2697 (N_2697,In_605,In_421);
xnor U2698 (N_2698,In_920,In_68);
and U2699 (N_2699,In_289,In_775);
or U2700 (N_2700,In_124,In_449);
and U2701 (N_2701,In_208,In_211);
nor U2702 (N_2702,In_81,In_190);
nand U2703 (N_2703,In_273,In_57);
or U2704 (N_2704,In_443,In_579);
or U2705 (N_2705,In_167,In_960);
and U2706 (N_2706,In_148,In_548);
nor U2707 (N_2707,In_825,In_684);
xor U2708 (N_2708,In_415,In_6);
and U2709 (N_2709,In_607,In_161);
nand U2710 (N_2710,In_926,In_325);
and U2711 (N_2711,In_109,In_48);
nand U2712 (N_2712,In_348,In_916);
nor U2713 (N_2713,In_895,In_590);
and U2714 (N_2714,In_615,In_3);
nand U2715 (N_2715,In_42,In_433);
and U2716 (N_2716,In_248,In_539);
and U2717 (N_2717,In_472,In_580);
xnor U2718 (N_2718,In_410,In_62);
xnor U2719 (N_2719,In_595,In_649);
nand U2720 (N_2720,In_913,In_79);
nor U2721 (N_2721,In_208,In_931);
nor U2722 (N_2722,In_894,In_341);
nand U2723 (N_2723,In_770,In_101);
nand U2724 (N_2724,In_295,In_791);
or U2725 (N_2725,In_38,In_984);
xor U2726 (N_2726,In_521,In_32);
and U2727 (N_2727,In_669,In_457);
xnor U2728 (N_2728,In_578,In_339);
nor U2729 (N_2729,In_311,In_905);
nand U2730 (N_2730,In_947,In_417);
nor U2731 (N_2731,In_963,In_996);
xnor U2732 (N_2732,In_217,In_236);
nor U2733 (N_2733,In_788,In_815);
nand U2734 (N_2734,In_311,In_303);
nor U2735 (N_2735,In_624,In_338);
nor U2736 (N_2736,In_803,In_379);
nand U2737 (N_2737,In_839,In_946);
nand U2738 (N_2738,In_782,In_607);
and U2739 (N_2739,In_672,In_303);
xor U2740 (N_2740,In_646,In_867);
xor U2741 (N_2741,In_32,In_95);
xnor U2742 (N_2742,In_483,In_168);
and U2743 (N_2743,In_912,In_731);
nand U2744 (N_2744,In_50,In_172);
or U2745 (N_2745,In_919,In_776);
nor U2746 (N_2746,In_405,In_323);
nand U2747 (N_2747,In_669,In_652);
xnor U2748 (N_2748,In_67,In_490);
nor U2749 (N_2749,In_8,In_942);
or U2750 (N_2750,In_712,In_888);
or U2751 (N_2751,In_663,In_992);
nand U2752 (N_2752,In_67,In_351);
nand U2753 (N_2753,In_234,In_645);
and U2754 (N_2754,In_972,In_711);
or U2755 (N_2755,In_216,In_210);
or U2756 (N_2756,In_379,In_939);
nor U2757 (N_2757,In_152,In_694);
nand U2758 (N_2758,In_812,In_788);
or U2759 (N_2759,In_56,In_409);
or U2760 (N_2760,In_908,In_792);
and U2761 (N_2761,In_662,In_130);
nand U2762 (N_2762,In_986,In_415);
or U2763 (N_2763,In_302,In_148);
nor U2764 (N_2764,In_951,In_366);
xor U2765 (N_2765,In_176,In_436);
nor U2766 (N_2766,In_336,In_541);
and U2767 (N_2767,In_816,In_989);
xnor U2768 (N_2768,In_838,In_2);
xor U2769 (N_2769,In_868,In_491);
or U2770 (N_2770,In_317,In_717);
and U2771 (N_2771,In_861,In_211);
and U2772 (N_2772,In_256,In_152);
nor U2773 (N_2773,In_798,In_963);
xnor U2774 (N_2774,In_138,In_486);
or U2775 (N_2775,In_913,In_642);
nor U2776 (N_2776,In_127,In_137);
xor U2777 (N_2777,In_123,In_731);
xor U2778 (N_2778,In_279,In_90);
xor U2779 (N_2779,In_294,In_237);
xor U2780 (N_2780,In_22,In_228);
nor U2781 (N_2781,In_996,In_67);
nand U2782 (N_2782,In_484,In_911);
and U2783 (N_2783,In_192,In_643);
nand U2784 (N_2784,In_891,In_299);
nor U2785 (N_2785,In_516,In_521);
xor U2786 (N_2786,In_786,In_79);
xnor U2787 (N_2787,In_704,In_748);
or U2788 (N_2788,In_881,In_10);
xor U2789 (N_2789,In_225,In_577);
and U2790 (N_2790,In_998,In_197);
xnor U2791 (N_2791,In_378,In_519);
xnor U2792 (N_2792,In_649,In_412);
and U2793 (N_2793,In_955,In_403);
nand U2794 (N_2794,In_482,In_347);
and U2795 (N_2795,In_513,In_245);
nor U2796 (N_2796,In_901,In_841);
nor U2797 (N_2797,In_227,In_372);
nor U2798 (N_2798,In_330,In_564);
xnor U2799 (N_2799,In_724,In_251);
or U2800 (N_2800,In_291,In_288);
xor U2801 (N_2801,In_759,In_37);
or U2802 (N_2802,In_80,In_952);
nand U2803 (N_2803,In_618,In_965);
nor U2804 (N_2804,In_724,In_132);
and U2805 (N_2805,In_771,In_40);
nor U2806 (N_2806,In_760,In_931);
and U2807 (N_2807,In_544,In_289);
xor U2808 (N_2808,In_685,In_366);
and U2809 (N_2809,In_439,In_363);
or U2810 (N_2810,In_800,In_392);
nor U2811 (N_2811,In_457,In_140);
xnor U2812 (N_2812,In_926,In_663);
and U2813 (N_2813,In_441,In_720);
nor U2814 (N_2814,In_680,In_95);
or U2815 (N_2815,In_418,In_419);
nand U2816 (N_2816,In_833,In_141);
or U2817 (N_2817,In_411,In_106);
nor U2818 (N_2818,In_895,In_43);
xnor U2819 (N_2819,In_215,In_531);
xnor U2820 (N_2820,In_668,In_501);
and U2821 (N_2821,In_949,In_198);
nand U2822 (N_2822,In_105,In_168);
nor U2823 (N_2823,In_452,In_684);
xor U2824 (N_2824,In_446,In_120);
or U2825 (N_2825,In_687,In_964);
nand U2826 (N_2826,In_639,In_51);
xnor U2827 (N_2827,In_261,In_585);
nor U2828 (N_2828,In_295,In_143);
xor U2829 (N_2829,In_17,In_731);
xnor U2830 (N_2830,In_966,In_237);
and U2831 (N_2831,In_192,In_732);
and U2832 (N_2832,In_911,In_305);
or U2833 (N_2833,In_855,In_639);
nand U2834 (N_2834,In_994,In_228);
xor U2835 (N_2835,In_316,In_40);
xnor U2836 (N_2836,In_299,In_51);
nor U2837 (N_2837,In_781,In_427);
and U2838 (N_2838,In_739,In_323);
xor U2839 (N_2839,In_211,In_376);
and U2840 (N_2840,In_998,In_341);
xnor U2841 (N_2841,In_453,In_729);
nor U2842 (N_2842,In_65,In_46);
xnor U2843 (N_2843,In_949,In_192);
nand U2844 (N_2844,In_82,In_790);
xnor U2845 (N_2845,In_106,In_815);
xnor U2846 (N_2846,In_699,In_603);
nor U2847 (N_2847,In_411,In_582);
or U2848 (N_2848,In_12,In_209);
and U2849 (N_2849,In_98,In_672);
and U2850 (N_2850,In_655,In_686);
xnor U2851 (N_2851,In_460,In_98);
or U2852 (N_2852,In_138,In_101);
or U2853 (N_2853,In_889,In_719);
nor U2854 (N_2854,In_405,In_189);
nor U2855 (N_2855,In_322,In_516);
xor U2856 (N_2856,In_652,In_715);
nand U2857 (N_2857,In_931,In_963);
nor U2858 (N_2858,In_869,In_389);
nand U2859 (N_2859,In_329,In_519);
xnor U2860 (N_2860,In_64,In_897);
nor U2861 (N_2861,In_916,In_898);
nand U2862 (N_2862,In_550,In_415);
nand U2863 (N_2863,In_554,In_638);
nand U2864 (N_2864,In_819,In_191);
xnor U2865 (N_2865,In_224,In_156);
nand U2866 (N_2866,In_57,In_136);
or U2867 (N_2867,In_228,In_788);
and U2868 (N_2868,In_780,In_472);
xnor U2869 (N_2869,In_325,In_435);
xnor U2870 (N_2870,In_554,In_372);
or U2871 (N_2871,In_759,In_595);
or U2872 (N_2872,In_593,In_81);
or U2873 (N_2873,In_783,In_348);
and U2874 (N_2874,In_854,In_943);
xnor U2875 (N_2875,In_777,In_601);
xor U2876 (N_2876,In_624,In_509);
nor U2877 (N_2877,In_414,In_598);
nor U2878 (N_2878,In_742,In_124);
nor U2879 (N_2879,In_61,In_284);
or U2880 (N_2880,In_485,In_768);
nor U2881 (N_2881,In_596,In_654);
nor U2882 (N_2882,In_706,In_569);
nand U2883 (N_2883,In_674,In_350);
xnor U2884 (N_2884,In_667,In_447);
nor U2885 (N_2885,In_486,In_3);
or U2886 (N_2886,In_638,In_507);
xnor U2887 (N_2887,In_662,In_860);
nor U2888 (N_2888,In_278,In_905);
or U2889 (N_2889,In_767,In_527);
nand U2890 (N_2890,In_409,In_895);
nand U2891 (N_2891,In_102,In_356);
and U2892 (N_2892,In_326,In_945);
or U2893 (N_2893,In_414,In_675);
nand U2894 (N_2894,In_33,In_872);
nor U2895 (N_2895,In_511,In_374);
nor U2896 (N_2896,In_907,In_777);
nand U2897 (N_2897,In_488,In_544);
or U2898 (N_2898,In_420,In_104);
xnor U2899 (N_2899,In_869,In_626);
and U2900 (N_2900,In_982,In_213);
nand U2901 (N_2901,In_366,In_733);
or U2902 (N_2902,In_627,In_923);
and U2903 (N_2903,In_947,In_619);
and U2904 (N_2904,In_194,In_961);
nand U2905 (N_2905,In_430,In_169);
and U2906 (N_2906,In_415,In_584);
nand U2907 (N_2907,In_459,In_382);
and U2908 (N_2908,In_401,In_899);
or U2909 (N_2909,In_16,In_646);
nand U2910 (N_2910,In_922,In_821);
nor U2911 (N_2911,In_743,In_725);
and U2912 (N_2912,In_867,In_249);
or U2913 (N_2913,In_697,In_684);
or U2914 (N_2914,In_619,In_982);
nand U2915 (N_2915,In_781,In_129);
nor U2916 (N_2916,In_472,In_910);
and U2917 (N_2917,In_572,In_126);
nor U2918 (N_2918,In_903,In_475);
xor U2919 (N_2919,In_561,In_967);
xor U2920 (N_2920,In_873,In_30);
nor U2921 (N_2921,In_6,In_800);
and U2922 (N_2922,In_948,In_586);
nor U2923 (N_2923,In_964,In_800);
nand U2924 (N_2924,In_402,In_604);
nor U2925 (N_2925,In_684,In_572);
nand U2926 (N_2926,In_430,In_503);
nor U2927 (N_2927,In_741,In_186);
or U2928 (N_2928,In_635,In_46);
xnor U2929 (N_2929,In_97,In_904);
nand U2930 (N_2930,In_332,In_229);
xnor U2931 (N_2931,In_366,In_428);
or U2932 (N_2932,In_657,In_9);
xor U2933 (N_2933,In_958,In_569);
xor U2934 (N_2934,In_926,In_239);
and U2935 (N_2935,In_751,In_135);
nand U2936 (N_2936,In_181,In_873);
or U2937 (N_2937,In_629,In_178);
or U2938 (N_2938,In_299,In_535);
xnor U2939 (N_2939,In_55,In_999);
or U2940 (N_2940,In_224,In_94);
nand U2941 (N_2941,In_797,In_327);
or U2942 (N_2942,In_677,In_195);
and U2943 (N_2943,In_426,In_48);
xnor U2944 (N_2944,In_839,In_776);
xor U2945 (N_2945,In_410,In_457);
or U2946 (N_2946,In_279,In_224);
or U2947 (N_2947,In_418,In_462);
nor U2948 (N_2948,In_47,In_654);
nand U2949 (N_2949,In_63,In_77);
nor U2950 (N_2950,In_143,In_445);
xnor U2951 (N_2951,In_263,In_473);
and U2952 (N_2952,In_683,In_257);
xor U2953 (N_2953,In_331,In_561);
nand U2954 (N_2954,In_147,In_847);
nand U2955 (N_2955,In_66,In_918);
xnor U2956 (N_2956,In_9,In_32);
nand U2957 (N_2957,In_7,In_605);
xnor U2958 (N_2958,In_710,In_771);
xor U2959 (N_2959,In_748,In_188);
xor U2960 (N_2960,In_742,In_501);
nor U2961 (N_2961,In_736,In_95);
and U2962 (N_2962,In_993,In_457);
nor U2963 (N_2963,In_394,In_897);
and U2964 (N_2964,In_670,In_870);
nor U2965 (N_2965,In_949,In_100);
xor U2966 (N_2966,In_100,In_68);
xnor U2967 (N_2967,In_145,In_888);
and U2968 (N_2968,In_205,In_607);
and U2969 (N_2969,In_202,In_383);
nor U2970 (N_2970,In_809,In_741);
nand U2971 (N_2971,In_193,In_203);
xnor U2972 (N_2972,In_891,In_707);
xnor U2973 (N_2973,In_282,In_451);
or U2974 (N_2974,In_473,In_55);
nor U2975 (N_2975,In_742,In_945);
nor U2976 (N_2976,In_299,In_249);
or U2977 (N_2977,In_907,In_386);
and U2978 (N_2978,In_951,In_63);
or U2979 (N_2979,In_172,In_978);
xnor U2980 (N_2980,In_882,In_802);
nor U2981 (N_2981,In_68,In_892);
or U2982 (N_2982,In_194,In_752);
and U2983 (N_2983,In_842,In_434);
and U2984 (N_2984,In_556,In_997);
or U2985 (N_2985,In_26,In_352);
and U2986 (N_2986,In_322,In_495);
xnor U2987 (N_2987,In_613,In_105);
and U2988 (N_2988,In_875,In_638);
xnor U2989 (N_2989,In_549,In_981);
or U2990 (N_2990,In_223,In_681);
xor U2991 (N_2991,In_922,In_977);
and U2992 (N_2992,In_442,In_853);
xor U2993 (N_2993,In_966,In_614);
nor U2994 (N_2994,In_487,In_434);
or U2995 (N_2995,In_449,In_997);
xnor U2996 (N_2996,In_855,In_772);
or U2997 (N_2997,In_320,In_688);
nor U2998 (N_2998,In_872,In_957);
xnor U2999 (N_2999,In_412,In_481);
nor U3000 (N_3000,In_802,In_186);
xor U3001 (N_3001,In_841,In_357);
and U3002 (N_3002,In_292,In_818);
nand U3003 (N_3003,In_280,In_20);
nand U3004 (N_3004,In_926,In_854);
nor U3005 (N_3005,In_228,In_618);
or U3006 (N_3006,In_691,In_586);
and U3007 (N_3007,In_21,In_632);
nand U3008 (N_3008,In_678,In_34);
nand U3009 (N_3009,In_554,In_679);
and U3010 (N_3010,In_756,In_326);
xor U3011 (N_3011,In_110,In_798);
xnor U3012 (N_3012,In_139,In_774);
and U3013 (N_3013,In_589,In_673);
nand U3014 (N_3014,In_562,In_24);
and U3015 (N_3015,In_472,In_573);
or U3016 (N_3016,In_91,In_521);
xor U3017 (N_3017,In_780,In_844);
or U3018 (N_3018,In_561,In_652);
nand U3019 (N_3019,In_569,In_961);
xor U3020 (N_3020,In_759,In_981);
nor U3021 (N_3021,In_324,In_260);
xnor U3022 (N_3022,In_235,In_292);
nor U3023 (N_3023,In_473,In_145);
nand U3024 (N_3024,In_520,In_615);
nand U3025 (N_3025,In_688,In_813);
nand U3026 (N_3026,In_807,In_771);
xnor U3027 (N_3027,In_188,In_198);
xor U3028 (N_3028,In_241,In_845);
nand U3029 (N_3029,In_994,In_341);
or U3030 (N_3030,In_965,In_534);
nor U3031 (N_3031,In_217,In_184);
nor U3032 (N_3032,In_700,In_669);
nor U3033 (N_3033,In_796,In_715);
and U3034 (N_3034,In_242,In_171);
or U3035 (N_3035,In_214,In_523);
nand U3036 (N_3036,In_229,In_466);
or U3037 (N_3037,In_142,In_226);
nand U3038 (N_3038,In_114,In_652);
nor U3039 (N_3039,In_290,In_752);
nand U3040 (N_3040,In_763,In_334);
nand U3041 (N_3041,In_950,In_142);
and U3042 (N_3042,In_362,In_408);
nor U3043 (N_3043,In_532,In_400);
nor U3044 (N_3044,In_170,In_569);
and U3045 (N_3045,In_288,In_160);
and U3046 (N_3046,In_596,In_714);
nand U3047 (N_3047,In_27,In_466);
nand U3048 (N_3048,In_173,In_774);
and U3049 (N_3049,In_186,In_323);
nor U3050 (N_3050,In_782,In_394);
or U3051 (N_3051,In_215,In_286);
nor U3052 (N_3052,In_856,In_390);
and U3053 (N_3053,In_367,In_744);
nand U3054 (N_3054,In_810,In_31);
nor U3055 (N_3055,In_565,In_309);
and U3056 (N_3056,In_942,In_975);
xor U3057 (N_3057,In_656,In_751);
xnor U3058 (N_3058,In_985,In_324);
xor U3059 (N_3059,In_493,In_323);
xor U3060 (N_3060,In_35,In_424);
or U3061 (N_3061,In_812,In_608);
xnor U3062 (N_3062,In_665,In_145);
or U3063 (N_3063,In_732,In_7);
nor U3064 (N_3064,In_760,In_721);
xor U3065 (N_3065,In_981,In_151);
nor U3066 (N_3066,In_571,In_765);
nor U3067 (N_3067,In_986,In_752);
or U3068 (N_3068,In_941,In_498);
xor U3069 (N_3069,In_151,In_15);
or U3070 (N_3070,In_174,In_711);
or U3071 (N_3071,In_488,In_872);
or U3072 (N_3072,In_591,In_940);
nand U3073 (N_3073,In_818,In_210);
nand U3074 (N_3074,In_754,In_115);
or U3075 (N_3075,In_612,In_850);
nor U3076 (N_3076,In_323,In_985);
and U3077 (N_3077,In_906,In_763);
or U3078 (N_3078,In_976,In_199);
and U3079 (N_3079,In_394,In_706);
and U3080 (N_3080,In_734,In_829);
or U3081 (N_3081,In_494,In_443);
xor U3082 (N_3082,In_901,In_81);
nor U3083 (N_3083,In_519,In_582);
and U3084 (N_3084,In_909,In_470);
and U3085 (N_3085,In_5,In_401);
xor U3086 (N_3086,In_86,In_818);
nor U3087 (N_3087,In_122,In_273);
xnor U3088 (N_3088,In_456,In_84);
nor U3089 (N_3089,In_180,In_134);
and U3090 (N_3090,In_765,In_249);
nand U3091 (N_3091,In_130,In_724);
and U3092 (N_3092,In_219,In_41);
nand U3093 (N_3093,In_573,In_916);
nand U3094 (N_3094,In_822,In_387);
and U3095 (N_3095,In_735,In_301);
and U3096 (N_3096,In_201,In_961);
and U3097 (N_3097,In_355,In_988);
nor U3098 (N_3098,In_243,In_115);
or U3099 (N_3099,In_15,In_993);
or U3100 (N_3100,In_944,In_734);
nand U3101 (N_3101,In_39,In_478);
and U3102 (N_3102,In_342,In_708);
and U3103 (N_3103,In_237,In_753);
or U3104 (N_3104,In_231,In_618);
nor U3105 (N_3105,In_535,In_353);
xnor U3106 (N_3106,In_118,In_435);
and U3107 (N_3107,In_0,In_665);
xor U3108 (N_3108,In_592,In_588);
nand U3109 (N_3109,In_504,In_211);
and U3110 (N_3110,In_555,In_892);
and U3111 (N_3111,In_16,In_400);
and U3112 (N_3112,In_149,In_430);
nor U3113 (N_3113,In_432,In_398);
and U3114 (N_3114,In_514,In_739);
nor U3115 (N_3115,In_765,In_611);
nand U3116 (N_3116,In_792,In_70);
nor U3117 (N_3117,In_920,In_508);
xor U3118 (N_3118,In_89,In_406);
and U3119 (N_3119,In_348,In_850);
and U3120 (N_3120,In_604,In_87);
and U3121 (N_3121,In_90,In_834);
nand U3122 (N_3122,In_372,In_454);
xnor U3123 (N_3123,In_452,In_60);
xnor U3124 (N_3124,In_333,In_224);
nor U3125 (N_3125,In_498,In_374);
nor U3126 (N_3126,In_79,In_139);
and U3127 (N_3127,In_811,In_76);
nand U3128 (N_3128,In_530,In_605);
nor U3129 (N_3129,In_645,In_844);
xnor U3130 (N_3130,In_511,In_633);
nand U3131 (N_3131,In_791,In_858);
xnor U3132 (N_3132,In_789,In_419);
and U3133 (N_3133,In_689,In_159);
nor U3134 (N_3134,In_418,In_930);
nor U3135 (N_3135,In_76,In_597);
or U3136 (N_3136,In_227,In_286);
or U3137 (N_3137,In_91,In_935);
nand U3138 (N_3138,In_879,In_667);
xor U3139 (N_3139,In_84,In_166);
xor U3140 (N_3140,In_363,In_28);
and U3141 (N_3141,In_884,In_368);
xor U3142 (N_3142,In_179,In_262);
or U3143 (N_3143,In_361,In_448);
and U3144 (N_3144,In_572,In_873);
nand U3145 (N_3145,In_392,In_553);
or U3146 (N_3146,In_337,In_47);
or U3147 (N_3147,In_692,In_133);
or U3148 (N_3148,In_144,In_349);
xor U3149 (N_3149,In_508,In_529);
nand U3150 (N_3150,In_548,In_461);
and U3151 (N_3151,In_401,In_429);
nor U3152 (N_3152,In_370,In_627);
xor U3153 (N_3153,In_195,In_948);
xnor U3154 (N_3154,In_34,In_629);
nor U3155 (N_3155,In_683,In_81);
nand U3156 (N_3156,In_633,In_38);
and U3157 (N_3157,In_635,In_91);
xnor U3158 (N_3158,In_662,In_515);
xor U3159 (N_3159,In_708,In_256);
nor U3160 (N_3160,In_502,In_99);
and U3161 (N_3161,In_427,In_486);
nor U3162 (N_3162,In_248,In_103);
nand U3163 (N_3163,In_699,In_349);
xnor U3164 (N_3164,In_437,In_237);
xor U3165 (N_3165,In_989,In_742);
nor U3166 (N_3166,In_890,In_843);
nor U3167 (N_3167,In_738,In_237);
xor U3168 (N_3168,In_246,In_773);
nor U3169 (N_3169,In_666,In_788);
nand U3170 (N_3170,In_155,In_503);
and U3171 (N_3171,In_501,In_384);
nor U3172 (N_3172,In_907,In_305);
and U3173 (N_3173,In_911,In_567);
nand U3174 (N_3174,In_607,In_829);
and U3175 (N_3175,In_802,In_341);
xnor U3176 (N_3176,In_527,In_140);
xor U3177 (N_3177,In_417,In_894);
or U3178 (N_3178,In_245,In_553);
and U3179 (N_3179,In_738,In_468);
or U3180 (N_3180,In_338,In_715);
and U3181 (N_3181,In_806,In_615);
and U3182 (N_3182,In_384,In_854);
and U3183 (N_3183,In_499,In_623);
nor U3184 (N_3184,In_438,In_666);
nor U3185 (N_3185,In_666,In_268);
nand U3186 (N_3186,In_722,In_828);
and U3187 (N_3187,In_799,In_55);
or U3188 (N_3188,In_738,In_483);
and U3189 (N_3189,In_164,In_168);
xor U3190 (N_3190,In_309,In_480);
and U3191 (N_3191,In_458,In_616);
nand U3192 (N_3192,In_819,In_422);
xnor U3193 (N_3193,In_300,In_537);
nor U3194 (N_3194,In_183,In_59);
xnor U3195 (N_3195,In_91,In_725);
xnor U3196 (N_3196,In_97,In_251);
xor U3197 (N_3197,In_265,In_447);
or U3198 (N_3198,In_506,In_313);
xor U3199 (N_3199,In_155,In_585);
nand U3200 (N_3200,In_690,In_117);
nor U3201 (N_3201,In_516,In_163);
xor U3202 (N_3202,In_913,In_868);
xnor U3203 (N_3203,In_351,In_323);
xnor U3204 (N_3204,In_385,In_366);
nor U3205 (N_3205,In_436,In_800);
nand U3206 (N_3206,In_415,In_754);
nand U3207 (N_3207,In_273,In_104);
xor U3208 (N_3208,In_220,In_629);
xor U3209 (N_3209,In_468,In_49);
nor U3210 (N_3210,In_799,In_776);
nor U3211 (N_3211,In_725,In_946);
nor U3212 (N_3212,In_420,In_864);
xnor U3213 (N_3213,In_137,In_628);
or U3214 (N_3214,In_407,In_317);
or U3215 (N_3215,In_84,In_727);
or U3216 (N_3216,In_839,In_854);
and U3217 (N_3217,In_953,In_417);
or U3218 (N_3218,In_103,In_661);
or U3219 (N_3219,In_614,In_177);
xnor U3220 (N_3220,In_466,In_749);
xor U3221 (N_3221,In_300,In_67);
xor U3222 (N_3222,In_401,In_324);
or U3223 (N_3223,In_983,In_157);
nor U3224 (N_3224,In_515,In_197);
or U3225 (N_3225,In_900,In_156);
and U3226 (N_3226,In_73,In_195);
xnor U3227 (N_3227,In_770,In_709);
or U3228 (N_3228,In_410,In_973);
or U3229 (N_3229,In_26,In_831);
nand U3230 (N_3230,In_469,In_463);
nand U3231 (N_3231,In_441,In_718);
xor U3232 (N_3232,In_263,In_435);
xnor U3233 (N_3233,In_426,In_22);
or U3234 (N_3234,In_636,In_888);
nor U3235 (N_3235,In_737,In_297);
or U3236 (N_3236,In_493,In_696);
nor U3237 (N_3237,In_125,In_642);
nand U3238 (N_3238,In_981,In_455);
or U3239 (N_3239,In_875,In_972);
or U3240 (N_3240,In_579,In_268);
and U3241 (N_3241,In_461,In_478);
nand U3242 (N_3242,In_658,In_369);
nand U3243 (N_3243,In_461,In_828);
or U3244 (N_3244,In_755,In_463);
xor U3245 (N_3245,In_753,In_548);
nor U3246 (N_3246,In_540,In_607);
nor U3247 (N_3247,In_745,In_100);
xor U3248 (N_3248,In_591,In_747);
nor U3249 (N_3249,In_193,In_353);
and U3250 (N_3250,In_652,In_625);
nand U3251 (N_3251,In_804,In_307);
nand U3252 (N_3252,In_437,In_796);
or U3253 (N_3253,In_809,In_9);
nand U3254 (N_3254,In_312,In_998);
and U3255 (N_3255,In_490,In_973);
xor U3256 (N_3256,In_404,In_96);
xnor U3257 (N_3257,In_25,In_632);
and U3258 (N_3258,In_183,In_945);
nor U3259 (N_3259,In_342,In_490);
nand U3260 (N_3260,In_51,In_295);
nand U3261 (N_3261,In_186,In_754);
nand U3262 (N_3262,In_883,In_534);
or U3263 (N_3263,In_525,In_425);
nand U3264 (N_3264,In_895,In_420);
and U3265 (N_3265,In_671,In_389);
xor U3266 (N_3266,In_741,In_954);
and U3267 (N_3267,In_534,In_593);
and U3268 (N_3268,In_92,In_574);
and U3269 (N_3269,In_697,In_218);
xnor U3270 (N_3270,In_453,In_347);
and U3271 (N_3271,In_223,In_553);
or U3272 (N_3272,In_921,In_855);
nand U3273 (N_3273,In_954,In_74);
or U3274 (N_3274,In_479,In_141);
or U3275 (N_3275,In_280,In_347);
nand U3276 (N_3276,In_493,In_653);
and U3277 (N_3277,In_544,In_898);
nor U3278 (N_3278,In_392,In_845);
or U3279 (N_3279,In_368,In_711);
nand U3280 (N_3280,In_254,In_873);
nor U3281 (N_3281,In_372,In_103);
and U3282 (N_3282,In_619,In_890);
xor U3283 (N_3283,In_363,In_431);
nor U3284 (N_3284,In_743,In_290);
nor U3285 (N_3285,In_521,In_932);
xor U3286 (N_3286,In_74,In_357);
nand U3287 (N_3287,In_411,In_35);
nor U3288 (N_3288,In_70,In_926);
or U3289 (N_3289,In_488,In_350);
nor U3290 (N_3290,In_416,In_165);
and U3291 (N_3291,In_49,In_477);
or U3292 (N_3292,In_254,In_872);
nand U3293 (N_3293,In_548,In_319);
or U3294 (N_3294,In_757,In_21);
xnor U3295 (N_3295,In_18,In_74);
and U3296 (N_3296,In_417,In_757);
and U3297 (N_3297,In_327,In_570);
xnor U3298 (N_3298,In_382,In_769);
and U3299 (N_3299,In_420,In_857);
or U3300 (N_3300,In_156,In_715);
and U3301 (N_3301,In_891,In_988);
and U3302 (N_3302,In_322,In_984);
and U3303 (N_3303,In_716,In_469);
nand U3304 (N_3304,In_229,In_863);
xor U3305 (N_3305,In_91,In_888);
xnor U3306 (N_3306,In_953,In_862);
and U3307 (N_3307,In_159,In_491);
xnor U3308 (N_3308,In_453,In_700);
and U3309 (N_3309,In_839,In_673);
nand U3310 (N_3310,In_144,In_450);
or U3311 (N_3311,In_55,In_427);
nor U3312 (N_3312,In_903,In_897);
and U3313 (N_3313,In_745,In_2);
or U3314 (N_3314,In_820,In_439);
nand U3315 (N_3315,In_258,In_113);
or U3316 (N_3316,In_199,In_573);
or U3317 (N_3317,In_654,In_892);
and U3318 (N_3318,In_941,In_852);
xnor U3319 (N_3319,In_589,In_803);
or U3320 (N_3320,In_474,In_168);
or U3321 (N_3321,In_422,In_730);
xor U3322 (N_3322,In_382,In_395);
and U3323 (N_3323,In_501,In_221);
and U3324 (N_3324,In_542,In_833);
xor U3325 (N_3325,In_959,In_54);
nand U3326 (N_3326,In_758,In_583);
nand U3327 (N_3327,In_964,In_176);
nand U3328 (N_3328,In_967,In_267);
xor U3329 (N_3329,In_19,In_218);
or U3330 (N_3330,In_604,In_715);
or U3331 (N_3331,In_583,In_236);
xor U3332 (N_3332,In_797,In_642);
or U3333 (N_3333,In_252,In_697);
and U3334 (N_3334,In_216,In_281);
and U3335 (N_3335,In_817,In_477);
or U3336 (N_3336,In_132,In_319);
nand U3337 (N_3337,In_305,In_835);
or U3338 (N_3338,In_536,In_409);
xnor U3339 (N_3339,In_451,In_302);
nor U3340 (N_3340,In_681,In_655);
nand U3341 (N_3341,In_849,In_418);
and U3342 (N_3342,In_12,In_617);
and U3343 (N_3343,In_13,In_546);
xnor U3344 (N_3344,In_730,In_641);
nand U3345 (N_3345,In_374,In_327);
and U3346 (N_3346,In_659,In_112);
xor U3347 (N_3347,In_628,In_778);
nand U3348 (N_3348,In_678,In_784);
nand U3349 (N_3349,In_280,In_124);
xor U3350 (N_3350,In_851,In_317);
or U3351 (N_3351,In_834,In_240);
nor U3352 (N_3352,In_202,In_847);
nor U3353 (N_3353,In_926,In_650);
nand U3354 (N_3354,In_749,In_871);
xnor U3355 (N_3355,In_350,In_927);
or U3356 (N_3356,In_581,In_465);
or U3357 (N_3357,In_777,In_625);
xor U3358 (N_3358,In_333,In_476);
nor U3359 (N_3359,In_854,In_747);
xor U3360 (N_3360,In_909,In_404);
or U3361 (N_3361,In_70,In_485);
nand U3362 (N_3362,In_781,In_576);
and U3363 (N_3363,In_106,In_672);
and U3364 (N_3364,In_238,In_214);
and U3365 (N_3365,In_144,In_543);
or U3366 (N_3366,In_423,In_893);
and U3367 (N_3367,In_676,In_188);
xnor U3368 (N_3368,In_838,In_837);
xnor U3369 (N_3369,In_246,In_967);
xor U3370 (N_3370,In_54,In_235);
or U3371 (N_3371,In_959,In_905);
nor U3372 (N_3372,In_386,In_376);
xor U3373 (N_3373,In_989,In_931);
or U3374 (N_3374,In_496,In_410);
and U3375 (N_3375,In_331,In_540);
nor U3376 (N_3376,In_948,In_295);
and U3377 (N_3377,In_949,In_596);
or U3378 (N_3378,In_882,In_125);
nand U3379 (N_3379,In_321,In_416);
nor U3380 (N_3380,In_993,In_521);
or U3381 (N_3381,In_487,In_874);
and U3382 (N_3382,In_637,In_889);
and U3383 (N_3383,In_752,In_571);
xor U3384 (N_3384,In_512,In_133);
and U3385 (N_3385,In_406,In_728);
and U3386 (N_3386,In_818,In_945);
nand U3387 (N_3387,In_962,In_2);
nand U3388 (N_3388,In_694,In_703);
and U3389 (N_3389,In_297,In_651);
and U3390 (N_3390,In_535,In_669);
nand U3391 (N_3391,In_349,In_151);
xor U3392 (N_3392,In_583,In_740);
xnor U3393 (N_3393,In_478,In_374);
nor U3394 (N_3394,In_992,In_432);
and U3395 (N_3395,In_945,In_111);
or U3396 (N_3396,In_515,In_344);
or U3397 (N_3397,In_316,In_902);
or U3398 (N_3398,In_977,In_877);
xnor U3399 (N_3399,In_375,In_427);
and U3400 (N_3400,In_578,In_924);
or U3401 (N_3401,In_888,In_991);
nand U3402 (N_3402,In_49,In_722);
nand U3403 (N_3403,In_994,In_715);
or U3404 (N_3404,In_747,In_580);
nand U3405 (N_3405,In_577,In_550);
nand U3406 (N_3406,In_22,In_775);
and U3407 (N_3407,In_925,In_106);
or U3408 (N_3408,In_663,In_706);
and U3409 (N_3409,In_523,In_398);
nor U3410 (N_3410,In_317,In_171);
xnor U3411 (N_3411,In_5,In_310);
nor U3412 (N_3412,In_232,In_134);
and U3413 (N_3413,In_717,In_989);
and U3414 (N_3414,In_330,In_529);
xnor U3415 (N_3415,In_507,In_443);
and U3416 (N_3416,In_720,In_296);
xor U3417 (N_3417,In_723,In_8);
or U3418 (N_3418,In_670,In_542);
xor U3419 (N_3419,In_859,In_851);
nand U3420 (N_3420,In_240,In_435);
nand U3421 (N_3421,In_506,In_682);
xor U3422 (N_3422,In_503,In_10);
xnor U3423 (N_3423,In_131,In_37);
nor U3424 (N_3424,In_432,In_933);
xnor U3425 (N_3425,In_309,In_543);
nand U3426 (N_3426,In_426,In_399);
or U3427 (N_3427,In_92,In_752);
nor U3428 (N_3428,In_925,In_731);
nand U3429 (N_3429,In_740,In_699);
or U3430 (N_3430,In_951,In_481);
nand U3431 (N_3431,In_212,In_457);
nor U3432 (N_3432,In_998,In_508);
xor U3433 (N_3433,In_290,In_260);
and U3434 (N_3434,In_564,In_957);
or U3435 (N_3435,In_489,In_632);
xor U3436 (N_3436,In_723,In_434);
nor U3437 (N_3437,In_517,In_535);
nor U3438 (N_3438,In_880,In_662);
xor U3439 (N_3439,In_31,In_560);
nand U3440 (N_3440,In_707,In_423);
nand U3441 (N_3441,In_608,In_712);
nand U3442 (N_3442,In_567,In_302);
xor U3443 (N_3443,In_347,In_943);
or U3444 (N_3444,In_595,In_273);
or U3445 (N_3445,In_884,In_22);
nand U3446 (N_3446,In_888,In_810);
and U3447 (N_3447,In_778,In_695);
nand U3448 (N_3448,In_399,In_693);
or U3449 (N_3449,In_237,In_896);
and U3450 (N_3450,In_781,In_683);
nor U3451 (N_3451,In_500,In_893);
xnor U3452 (N_3452,In_412,In_456);
and U3453 (N_3453,In_518,In_687);
or U3454 (N_3454,In_481,In_898);
xor U3455 (N_3455,In_822,In_97);
or U3456 (N_3456,In_425,In_250);
or U3457 (N_3457,In_285,In_511);
nor U3458 (N_3458,In_651,In_90);
or U3459 (N_3459,In_930,In_259);
and U3460 (N_3460,In_4,In_235);
and U3461 (N_3461,In_612,In_452);
nor U3462 (N_3462,In_812,In_519);
nor U3463 (N_3463,In_926,In_679);
nor U3464 (N_3464,In_824,In_361);
and U3465 (N_3465,In_100,In_964);
and U3466 (N_3466,In_673,In_576);
and U3467 (N_3467,In_668,In_950);
and U3468 (N_3468,In_740,In_731);
nor U3469 (N_3469,In_752,In_252);
or U3470 (N_3470,In_919,In_712);
and U3471 (N_3471,In_179,In_151);
nand U3472 (N_3472,In_229,In_279);
or U3473 (N_3473,In_860,In_566);
nor U3474 (N_3474,In_786,In_785);
nor U3475 (N_3475,In_543,In_928);
or U3476 (N_3476,In_696,In_45);
nor U3477 (N_3477,In_580,In_643);
nand U3478 (N_3478,In_402,In_930);
and U3479 (N_3479,In_916,In_407);
xnor U3480 (N_3480,In_861,In_988);
xnor U3481 (N_3481,In_593,In_157);
nand U3482 (N_3482,In_274,In_372);
xnor U3483 (N_3483,In_521,In_34);
and U3484 (N_3484,In_342,In_964);
nor U3485 (N_3485,In_887,In_321);
nor U3486 (N_3486,In_680,In_672);
or U3487 (N_3487,In_214,In_32);
and U3488 (N_3488,In_364,In_799);
nand U3489 (N_3489,In_698,In_768);
nand U3490 (N_3490,In_450,In_574);
or U3491 (N_3491,In_363,In_885);
and U3492 (N_3492,In_168,In_925);
nand U3493 (N_3493,In_898,In_528);
and U3494 (N_3494,In_720,In_779);
or U3495 (N_3495,In_179,In_56);
nand U3496 (N_3496,In_453,In_0);
xnor U3497 (N_3497,In_372,In_331);
or U3498 (N_3498,In_323,In_350);
xnor U3499 (N_3499,In_371,In_103);
and U3500 (N_3500,In_7,In_113);
or U3501 (N_3501,In_156,In_405);
and U3502 (N_3502,In_609,In_24);
nand U3503 (N_3503,In_961,In_653);
and U3504 (N_3504,In_478,In_595);
nand U3505 (N_3505,In_354,In_209);
and U3506 (N_3506,In_429,In_11);
and U3507 (N_3507,In_75,In_403);
nand U3508 (N_3508,In_145,In_293);
nand U3509 (N_3509,In_581,In_455);
nor U3510 (N_3510,In_956,In_930);
nand U3511 (N_3511,In_547,In_766);
xor U3512 (N_3512,In_56,In_310);
xnor U3513 (N_3513,In_631,In_108);
nor U3514 (N_3514,In_634,In_63);
nor U3515 (N_3515,In_246,In_565);
xor U3516 (N_3516,In_690,In_370);
or U3517 (N_3517,In_530,In_122);
or U3518 (N_3518,In_697,In_874);
xor U3519 (N_3519,In_245,In_177);
nand U3520 (N_3520,In_511,In_396);
nor U3521 (N_3521,In_346,In_883);
nor U3522 (N_3522,In_523,In_303);
or U3523 (N_3523,In_320,In_273);
or U3524 (N_3524,In_54,In_122);
or U3525 (N_3525,In_731,In_210);
nand U3526 (N_3526,In_746,In_482);
or U3527 (N_3527,In_616,In_592);
and U3528 (N_3528,In_973,In_438);
and U3529 (N_3529,In_43,In_923);
nand U3530 (N_3530,In_389,In_763);
or U3531 (N_3531,In_865,In_295);
and U3532 (N_3532,In_320,In_442);
and U3533 (N_3533,In_961,In_478);
nand U3534 (N_3534,In_725,In_913);
nor U3535 (N_3535,In_822,In_960);
nand U3536 (N_3536,In_267,In_868);
or U3537 (N_3537,In_953,In_272);
xnor U3538 (N_3538,In_810,In_709);
nor U3539 (N_3539,In_821,In_351);
nor U3540 (N_3540,In_675,In_696);
xnor U3541 (N_3541,In_584,In_220);
nand U3542 (N_3542,In_972,In_417);
xor U3543 (N_3543,In_432,In_648);
and U3544 (N_3544,In_596,In_162);
nand U3545 (N_3545,In_356,In_275);
nor U3546 (N_3546,In_911,In_332);
or U3547 (N_3547,In_986,In_137);
or U3548 (N_3548,In_880,In_523);
nor U3549 (N_3549,In_501,In_788);
nand U3550 (N_3550,In_677,In_501);
and U3551 (N_3551,In_495,In_413);
nand U3552 (N_3552,In_464,In_58);
nand U3553 (N_3553,In_146,In_433);
nand U3554 (N_3554,In_17,In_423);
nor U3555 (N_3555,In_294,In_569);
xnor U3556 (N_3556,In_879,In_946);
or U3557 (N_3557,In_71,In_680);
and U3558 (N_3558,In_818,In_385);
and U3559 (N_3559,In_714,In_846);
or U3560 (N_3560,In_476,In_325);
or U3561 (N_3561,In_74,In_81);
or U3562 (N_3562,In_509,In_664);
and U3563 (N_3563,In_863,In_249);
or U3564 (N_3564,In_466,In_425);
nand U3565 (N_3565,In_370,In_650);
nor U3566 (N_3566,In_663,In_712);
or U3567 (N_3567,In_792,In_221);
nand U3568 (N_3568,In_214,In_984);
nor U3569 (N_3569,In_715,In_493);
or U3570 (N_3570,In_482,In_687);
xnor U3571 (N_3571,In_807,In_542);
nand U3572 (N_3572,In_74,In_278);
or U3573 (N_3573,In_62,In_213);
and U3574 (N_3574,In_471,In_428);
xnor U3575 (N_3575,In_953,In_766);
or U3576 (N_3576,In_919,In_421);
xnor U3577 (N_3577,In_561,In_588);
xnor U3578 (N_3578,In_909,In_910);
nand U3579 (N_3579,In_144,In_767);
nand U3580 (N_3580,In_292,In_593);
xor U3581 (N_3581,In_39,In_376);
or U3582 (N_3582,In_491,In_87);
and U3583 (N_3583,In_667,In_762);
and U3584 (N_3584,In_307,In_596);
xnor U3585 (N_3585,In_93,In_771);
nand U3586 (N_3586,In_828,In_47);
nand U3587 (N_3587,In_390,In_532);
nand U3588 (N_3588,In_709,In_234);
or U3589 (N_3589,In_554,In_982);
and U3590 (N_3590,In_187,In_334);
or U3591 (N_3591,In_549,In_792);
or U3592 (N_3592,In_807,In_451);
nand U3593 (N_3593,In_709,In_641);
or U3594 (N_3594,In_281,In_895);
and U3595 (N_3595,In_871,In_632);
xnor U3596 (N_3596,In_614,In_938);
nor U3597 (N_3597,In_246,In_586);
and U3598 (N_3598,In_282,In_882);
or U3599 (N_3599,In_564,In_951);
nand U3600 (N_3600,In_978,In_441);
nor U3601 (N_3601,In_857,In_911);
nor U3602 (N_3602,In_47,In_83);
xor U3603 (N_3603,In_399,In_375);
or U3604 (N_3604,In_809,In_451);
nand U3605 (N_3605,In_877,In_139);
nand U3606 (N_3606,In_693,In_188);
xor U3607 (N_3607,In_895,In_642);
nand U3608 (N_3608,In_197,In_661);
or U3609 (N_3609,In_301,In_942);
nor U3610 (N_3610,In_710,In_888);
and U3611 (N_3611,In_939,In_319);
and U3612 (N_3612,In_898,In_631);
xnor U3613 (N_3613,In_638,In_676);
nor U3614 (N_3614,In_136,In_918);
nand U3615 (N_3615,In_648,In_523);
xnor U3616 (N_3616,In_244,In_309);
xnor U3617 (N_3617,In_358,In_985);
and U3618 (N_3618,In_393,In_389);
nand U3619 (N_3619,In_677,In_388);
or U3620 (N_3620,In_760,In_153);
nor U3621 (N_3621,In_662,In_382);
or U3622 (N_3622,In_411,In_586);
and U3623 (N_3623,In_210,In_241);
nor U3624 (N_3624,In_115,In_353);
and U3625 (N_3625,In_240,In_437);
xor U3626 (N_3626,In_475,In_360);
xor U3627 (N_3627,In_585,In_710);
xor U3628 (N_3628,In_353,In_855);
or U3629 (N_3629,In_250,In_133);
and U3630 (N_3630,In_22,In_978);
xor U3631 (N_3631,In_866,In_928);
nor U3632 (N_3632,In_132,In_200);
nor U3633 (N_3633,In_622,In_540);
or U3634 (N_3634,In_442,In_577);
or U3635 (N_3635,In_711,In_645);
or U3636 (N_3636,In_943,In_207);
nor U3637 (N_3637,In_507,In_502);
or U3638 (N_3638,In_703,In_948);
nor U3639 (N_3639,In_95,In_778);
and U3640 (N_3640,In_802,In_200);
nand U3641 (N_3641,In_432,In_812);
or U3642 (N_3642,In_36,In_97);
and U3643 (N_3643,In_899,In_890);
xnor U3644 (N_3644,In_568,In_706);
nand U3645 (N_3645,In_679,In_248);
nor U3646 (N_3646,In_999,In_708);
or U3647 (N_3647,In_622,In_340);
nand U3648 (N_3648,In_172,In_280);
nand U3649 (N_3649,In_729,In_84);
or U3650 (N_3650,In_765,In_301);
or U3651 (N_3651,In_55,In_950);
nor U3652 (N_3652,In_312,In_986);
xnor U3653 (N_3653,In_651,In_64);
nor U3654 (N_3654,In_848,In_526);
nor U3655 (N_3655,In_927,In_98);
nand U3656 (N_3656,In_151,In_944);
xnor U3657 (N_3657,In_517,In_434);
xor U3658 (N_3658,In_170,In_494);
nor U3659 (N_3659,In_499,In_680);
nand U3660 (N_3660,In_531,In_699);
xnor U3661 (N_3661,In_570,In_624);
nand U3662 (N_3662,In_23,In_320);
xor U3663 (N_3663,In_147,In_571);
xor U3664 (N_3664,In_310,In_297);
nor U3665 (N_3665,In_470,In_424);
xor U3666 (N_3666,In_582,In_841);
nand U3667 (N_3667,In_705,In_681);
and U3668 (N_3668,In_227,In_143);
nand U3669 (N_3669,In_759,In_88);
nand U3670 (N_3670,In_560,In_89);
and U3671 (N_3671,In_380,In_782);
nor U3672 (N_3672,In_982,In_649);
or U3673 (N_3673,In_153,In_941);
xnor U3674 (N_3674,In_656,In_348);
xor U3675 (N_3675,In_806,In_817);
xnor U3676 (N_3676,In_15,In_678);
nor U3677 (N_3677,In_492,In_175);
nor U3678 (N_3678,In_947,In_56);
and U3679 (N_3679,In_235,In_634);
xnor U3680 (N_3680,In_983,In_709);
nor U3681 (N_3681,In_918,In_948);
nand U3682 (N_3682,In_104,In_63);
xor U3683 (N_3683,In_740,In_544);
nor U3684 (N_3684,In_643,In_935);
xnor U3685 (N_3685,In_994,In_148);
xnor U3686 (N_3686,In_960,In_369);
nor U3687 (N_3687,In_78,In_443);
nand U3688 (N_3688,In_213,In_93);
or U3689 (N_3689,In_884,In_132);
nand U3690 (N_3690,In_885,In_790);
or U3691 (N_3691,In_522,In_629);
xnor U3692 (N_3692,In_427,In_753);
nor U3693 (N_3693,In_619,In_258);
nor U3694 (N_3694,In_411,In_246);
nand U3695 (N_3695,In_991,In_431);
or U3696 (N_3696,In_397,In_40);
and U3697 (N_3697,In_834,In_718);
or U3698 (N_3698,In_586,In_275);
nand U3699 (N_3699,In_560,In_988);
nor U3700 (N_3700,In_842,In_879);
or U3701 (N_3701,In_36,In_993);
or U3702 (N_3702,In_965,In_414);
or U3703 (N_3703,In_676,In_205);
nand U3704 (N_3704,In_514,In_500);
xor U3705 (N_3705,In_243,In_57);
and U3706 (N_3706,In_525,In_267);
nand U3707 (N_3707,In_250,In_608);
nand U3708 (N_3708,In_218,In_181);
or U3709 (N_3709,In_713,In_601);
nand U3710 (N_3710,In_643,In_517);
nand U3711 (N_3711,In_561,In_473);
nand U3712 (N_3712,In_693,In_375);
nor U3713 (N_3713,In_115,In_276);
nor U3714 (N_3714,In_603,In_424);
nor U3715 (N_3715,In_200,In_67);
xnor U3716 (N_3716,In_247,In_783);
nor U3717 (N_3717,In_992,In_272);
or U3718 (N_3718,In_254,In_406);
nor U3719 (N_3719,In_295,In_459);
or U3720 (N_3720,In_65,In_59);
or U3721 (N_3721,In_697,In_84);
nand U3722 (N_3722,In_748,In_492);
xor U3723 (N_3723,In_811,In_870);
nand U3724 (N_3724,In_599,In_293);
nand U3725 (N_3725,In_552,In_617);
xnor U3726 (N_3726,In_154,In_27);
and U3727 (N_3727,In_437,In_838);
nor U3728 (N_3728,In_206,In_449);
and U3729 (N_3729,In_609,In_238);
nor U3730 (N_3730,In_868,In_139);
or U3731 (N_3731,In_251,In_732);
xnor U3732 (N_3732,In_2,In_701);
xnor U3733 (N_3733,In_17,In_133);
nand U3734 (N_3734,In_500,In_439);
xor U3735 (N_3735,In_679,In_915);
and U3736 (N_3736,In_283,In_71);
xor U3737 (N_3737,In_416,In_127);
xnor U3738 (N_3738,In_322,In_656);
nor U3739 (N_3739,In_552,In_409);
nand U3740 (N_3740,In_575,In_961);
and U3741 (N_3741,In_296,In_851);
nand U3742 (N_3742,In_85,In_485);
or U3743 (N_3743,In_259,In_876);
xnor U3744 (N_3744,In_223,In_148);
nor U3745 (N_3745,In_686,In_320);
nor U3746 (N_3746,In_633,In_122);
nand U3747 (N_3747,In_719,In_851);
nand U3748 (N_3748,In_133,In_656);
nor U3749 (N_3749,In_256,In_951);
nor U3750 (N_3750,In_527,In_863);
and U3751 (N_3751,In_320,In_456);
and U3752 (N_3752,In_132,In_992);
nor U3753 (N_3753,In_602,In_674);
and U3754 (N_3754,In_472,In_739);
and U3755 (N_3755,In_886,In_68);
and U3756 (N_3756,In_378,In_468);
nand U3757 (N_3757,In_998,In_272);
xnor U3758 (N_3758,In_580,In_130);
nor U3759 (N_3759,In_718,In_642);
and U3760 (N_3760,In_36,In_54);
nand U3761 (N_3761,In_865,In_855);
nand U3762 (N_3762,In_936,In_645);
nand U3763 (N_3763,In_90,In_621);
nor U3764 (N_3764,In_172,In_684);
and U3765 (N_3765,In_446,In_136);
xnor U3766 (N_3766,In_878,In_481);
nor U3767 (N_3767,In_95,In_585);
xnor U3768 (N_3768,In_899,In_177);
nor U3769 (N_3769,In_562,In_256);
nand U3770 (N_3770,In_87,In_958);
xnor U3771 (N_3771,In_245,In_866);
nand U3772 (N_3772,In_13,In_796);
or U3773 (N_3773,In_506,In_23);
or U3774 (N_3774,In_880,In_27);
xor U3775 (N_3775,In_831,In_944);
or U3776 (N_3776,In_406,In_486);
nor U3777 (N_3777,In_914,In_538);
and U3778 (N_3778,In_188,In_999);
and U3779 (N_3779,In_476,In_677);
and U3780 (N_3780,In_583,In_946);
xor U3781 (N_3781,In_341,In_288);
or U3782 (N_3782,In_561,In_319);
xnor U3783 (N_3783,In_324,In_302);
nand U3784 (N_3784,In_983,In_198);
xor U3785 (N_3785,In_489,In_33);
nor U3786 (N_3786,In_704,In_590);
or U3787 (N_3787,In_697,In_266);
xor U3788 (N_3788,In_450,In_64);
or U3789 (N_3789,In_862,In_97);
and U3790 (N_3790,In_621,In_443);
or U3791 (N_3791,In_718,In_692);
nand U3792 (N_3792,In_990,In_424);
nand U3793 (N_3793,In_553,In_429);
nand U3794 (N_3794,In_322,In_416);
nor U3795 (N_3795,In_710,In_617);
and U3796 (N_3796,In_840,In_679);
nor U3797 (N_3797,In_550,In_648);
nand U3798 (N_3798,In_646,In_553);
and U3799 (N_3799,In_459,In_724);
nor U3800 (N_3800,In_251,In_764);
xnor U3801 (N_3801,In_414,In_841);
xor U3802 (N_3802,In_432,In_559);
xor U3803 (N_3803,In_936,In_434);
nand U3804 (N_3804,In_231,In_426);
and U3805 (N_3805,In_973,In_387);
or U3806 (N_3806,In_214,In_948);
xor U3807 (N_3807,In_884,In_420);
nand U3808 (N_3808,In_77,In_953);
xor U3809 (N_3809,In_28,In_815);
nand U3810 (N_3810,In_258,In_216);
nor U3811 (N_3811,In_576,In_917);
nand U3812 (N_3812,In_583,In_677);
nor U3813 (N_3813,In_354,In_954);
and U3814 (N_3814,In_577,In_427);
xor U3815 (N_3815,In_538,In_985);
xnor U3816 (N_3816,In_340,In_937);
nand U3817 (N_3817,In_314,In_255);
xor U3818 (N_3818,In_89,In_892);
nand U3819 (N_3819,In_767,In_10);
and U3820 (N_3820,In_870,In_183);
and U3821 (N_3821,In_766,In_862);
or U3822 (N_3822,In_823,In_932);
and U3823 (N_3823,In_794,In_966);
xor U3824 (N_3824,In_991,In_957);
nand U3825 (N_3825,In_704,In_946);
or U3826 (N_3826,In_296,In_510);
nand U3827 (N_3827,In_612,In_477);
xnor U3828 (N_3828,In_667,In_922);
and U3829 (N_3829,In_184,In_706);
xor U3830 (N_3830,In_752,In_333);
nand U3831 (N_3831,In_301,In_727);
or U3832 (N_3832,In_808,In_856);
nand U3833 (N_3833,In_416,In_305);
or U3834 (N_3834,In_35,In_799);
nor U3835 (N_3835,In_55,In_790);
xnor U3836 (N_3836,In_4,In_344);
and U3837 (N_3837,In_74,In_79);
and U3838 (N_3838,In_114,In_429);
nand U3839 (N_3839,In_965,In_719);
and U3840 (N_3840,In_394,In_354);
nand U3841 (N_3841,In_824,In_46);
xor U3842 (N_3842,In_615,In_136);
and U3843 (N_3843,In_812,In_146);
xor U3844 (N_3844,In_291,In_912);
nand U3845 (N_3845,In_798,In_24);
xor U3846 (N_3846,In_465,In_536);
xor U3847 (N_3847,In_722,In_486);
or U3848 (N_3848,In_666,In_127);
xnor U3849 (N_3849,In_576,In_983);
or U3850 (N_3850,In_363,In_404);
xor U3851 (N_3851,In_882,In_52);
or U3852 (N_3852,In_207,In_763);
nor U3853 (N_3853,In_137,In_546);
and U3854 (N_3854,In_492,In_915);
or U3855 (N_3855,In_513,In_747);
or U3856 (N_3856,In_634,In_316);
and U3857 (N_3857,In_565,In_242);
nor U3858 (N_3858,In_735,In_620);
nand U3859 (N_3859,In_673,In_457);
and U3860 (N_3860,In_207,In_384);
nand U3861 (N_3861,In_288,In_762);
and U3862 (N_3862,In_456,In_241);
or U3863 (N_3863,In_397,In_152);
and U3864 (N_3864,In_460,In_368);
nor U3865 (N_3865,In_85,In_674);
nor U3866 (N_3866,In_988,In_184);
nand U3867 (N_3867,In_565,In_172);
and U3868 (N_3868,In_549,In_708);
nor U3869 (N_3869,In_702,In_238);
xor U3870 (N_3870,In_43,In_847);
and U3871 (N_3871,In_413,In_550);
nor U3872 (N_3872,In_473,In_690);
xor U3873 (N_3873,In_623,In_466);
nor U3874 (N_3874,In_426,In_141);
nor U3875 (N_3875,In_531,In_484);
xor U3876 (N_3876,In_792,In_269);
xor U3877 (N_3877,In_445,In_270);
and U3878 (N_3878,In_419,In_33);
nor U3879 (N_3879,In_249,In_557);
xor U3880 (N_3880,In_460,In_660);
and U3881 (N_3881,In_59,In_124);
and U3882 (N_3882,In_588,In_522);
or U3883 (N_3883,In_260,In_617);
nand U3884 (N_3884,In_164,In_351);
or U3885 (N_3885,In_357,In_467);
and U3886 (N_3886,In_281,In_379);
or U3887 (N_3887,In_682,In_290);
nand U3888 (N_3888,In_910,In_626);
nand U3889 (N_3889,In_837,In_988);
or U3890 (N_3890,In_539,In_699);
or U3891 (N_3891,In_895,In_502);
xor U3892 (N_3892,In_886,In_821);
or U3893 (N_3893,In_834,In_65);
xnor U3894 (N_3894,In_289,In_749);
nand U3895 (N_3895,In_642,In_171);
nor U3896 (N_3896,In_647,In_677);
or U3897 (N_3897,In_700,In_872);
nor U3898 (N_3898,In_959,In_309);
xor U3899 (N_3899,In_451,In_501);
xor U3900 (N_3900,In_912,In_422);
and U3901 (N_3901,In_970,In_475);
or U3902 (N_3902,In_46,In_682);
xnor U3903 (N_3903,In_914,In_183);
xor U3904 (N_3904,In_669,In_143);
xnor U3905 (N_3905,In_91,In_652);
nand U3906 (N_3906,In_744,In_434);
or U3907 (N_3907,In_634,In_556);
and U3908 (N_3908,In_411,In_160);
or U3909 (N_3909,In_127,In_592);
nor U3910 (N_3910,In_105,In_784);
nor U3911 (N_3911,In_385,In_641);
or U3912 (N_3912,In_673,In_231);
nand U3913 (N_3913,In_605,In_975);
nor U3914 (N_3914,In_52,In_34);
nand U3915 (N_3915,In_165,In_483);
or U3916 (N_3916,In_636,In_154);
nor U3917 (N_3917,In_234,In_85);
or U3918 (N_3918,In_287,In_213);
and U3919 (N_3919,In_675,In_747);
xnor U3920 (N_3920,In_634,In_793);
xnor U3921 (N_3921,In_418,In_304);
nor U3922 (N_3922,In_873,In_365);
xnor U3923 (N_3923,In_240,In_376);
xor U3924 (N_3924,In_585,In_411);
xnor U3925 (N_3925,In_519,In_626);
nor U3926 (N_3926,In_329,In_814);
or U3927 (N_3927,In_486,In_309);
nor U3928 (N_3928,In_966,In_593);
and U3929 (N_3929,In_156,In_737);
nand U3930 (N_3930,In_944,In_143);
nor U3931 (N_3931,In_987,In_944);
or U3932 (N_3932,In_790,In_859);
or U3933 (N_3933,In_244,In_716);
or U3934 (N_3934,In_606,In_632);
xnor U3935 (N_3935,In_955,In_573);
nor U3936 (N_3936,In_13,In_261);
nand U3937 (N_3937,In_365,In_376);
or U3938 (N_3938,In_154,In_266);
nand U3939 (N_3939,In_49,In_545);
nor U3940 (N_3940,In_395,In_643);
xor U3941 (N_3941,In_797,In_438);
or U3942 (N_3942,In_806,In_48);
or U3943 (N_3943,In_924,In_624);
nand U3944 (N_3944,In_464,In_875);
xnor U3945 (N_3945,In_139,In_383);
and U3946 (N_3946,In_562,In_711);
or U3947 (N_3947,In_30,In_210);
and U3948 (N_3948,In_229,In_483);
nor U3949 (N_3949,In_879,In_883);
nor U3950 (N_3950,In_600,In_804);
or U3951 (N_3951,In_84,In_396);
nor U3952 (N_3952,In_520,In_314);
nor U3953 (N_3953,In_289,In_415);
nor U3954 (N_3954,In_660,In_296);
nor U3955 (N_3955,In_663,In_409);
nand U3956 (N_3956,In_353,In_397);
or U3957 (N_3957,In_148,In_241);
or U3958 (N_3958,In_401,In_206);
or U3959 (N_3959,In_936,In_416);
xor U3960 (N_3960,In_956,In_375);
or U3961 (N_3961,In_91,In_800);
xnor U3962 (N_3962,In_880,In_747);
nand U3963 (N_3963,In_854,In_644);
nand U3964 (N_3964,In_20,In_872);
or U3965 (N_3965,In_455,In_442);
nand U3966 (N_3966,In_431,In_230);
nand U3967 (N_3967,In_893,In_75);
or U3968 (N_3968,In_101,In_686);
nor U3969 (N_3969,In_601,In_626);
nand U3970 (N_3970,In_864,In_741);
xor U3971 (N_3971,In_154,In_3);
and U3972 (N_3972,In_569,In_363);
nor U3973 (N_3973,In_759,In_829);
or U3974 (N_3974,In_137,In_38);
xnor U3975 (N_3975,In_894,In_113);
nand U3976 (N_3976,In_563,In_626);
or U3977 (N_3977,In_360,In_657);
and U3978 (N_3978,In_970,In_559);
xnor U3979 (N_3979,In_135,In_796);
nand U3980 (N_3980,In_86,In_645);
nand U3981 (N_3981,In_184,In_497);
xor U3982 (N_3982,In_268,In_434);
nor U3983 (N_3983,In_51,In_440);
xnor U3984 (N_3984,In_498,In_938);
or U3985 (N_3985,In_641,In_243);
and U3986 (N_3986,In_175,In_999);
nor U3987 (N_3987,In_453,In_135);
or U3988 (N_3988,In_164,In_540);
nand U3989 (N_3989,In_277,In_918);
nand U3990 (N_3990,In_12,In_345);
or U3991 (N_3991,In_548,In_962);
nor U3992 (N_3992,In_454,In_833);
or U3993 (N_3993,In_109,In_290);
or U3994 (N_3994,In_381,In_657);
or U3995 (N_3995,In_20,In_632);
or U3996 (N_3996,In_772,In_775);
nand U3997 (N_3997,In_241,In_130);
nor U3998 (N_3998,In_846,In_732);
nand U3999 (N_3999,In_329,In_24);
xor U4000 (N_4000,In_538,In_614);
and U4001 (N_4001,In_356,In_224);
and U4002 (N_4002,In_39,In_579);
and U4003 (N_4003,In_877,In_572);
nand U4004 (N_4004,In_584,In_186);
xor U4005 (N_4005,In_449,In_237);
or U4006 (N_4006,In_973,In_399);
xnor U4007 (N_4007,In_324,In_303);
nor U4008 (N_4008,In_155,In_534);
nand U4009 (N_4009,In_453,In_765);
and U4010 (N_4010,In_664,In_132);
and U4011 (N_4011,In_454,In_306);
and U4012 (N_4012,In_847,In_88);
or U4013 (N_4013,In_407,In_897);
nand U4014 (N_4014,In_428,In_166);
nor U4015 (N_4015,In_802,In_603);
xor U4016 (N_4016,In_865,In_799);
nand U4017 (N_4017,In_237,In_822);
nand U4018 (N_4018,In_829,In_817);
nand U4019 (N_4019,In_699,In_322);
and U4020 (N_4020,In_31,In_339);
nand U4021 (N_4021,In_174,In_355);
xnor U4022 (N_4022,In_600,In_520);
or U4023 (N_4023,In_500,In_925);
and U4024 (N_4024,In_108,In_929);
xor U4025 (N_4025,In_13,In_492);
nor U4026 (N_4026,In_205,In_396);
and U4027 (N_4027,In_139,In_854);
xnor U4028 (N_4028,In_285,In_490);
and U4029 (N_4029,In_400,In_753);
or U4030 (N_4030,In_474,In_906);
xnor U4031 (N_4031,In_106,In_758);
or U4032 (N_4032,In_489,In_216);
nor U4033 (N_4033,In_756,In_799);
nor U4034 (N_4034,In_401,In_738);
xnor U4035 (N_4035,In_63,In_140);
xnor U4036 (N_4036,In_44,In_605);
and U4037 (N_4037,In_516,In_458);
and U4038 (N_4038,In_613,In_501);
or U4039 (N_4039,In_642,In_745);
and U4040 (N_4040,In_482,In_728);
or U4041 (N_4041,In_518,In_584);
or U4042 (N_4042,In_9,In_570);
and U4043 (N_4043,In_647,In_101);
nor U4044 (N_4044,In_280,In_176);
nand U4045 (N_4045,In_212,In_649);
and U4046 (N_4046,In_170,In_626);
nor U4047 (N_4047,In_58,In_252);
and U4048 (N_4048,In_447,In_671);
nor U4049 (N_4049,In_674,In_225);
nand U4050 (N_4050,In_145,In_425);
nor U4051 (N_4051,In_16,In_756);
xnor U4052 (N_4052,In_650,In_377);
or U4053 (N_4053,In_779,In_99);
or U4054 (N_4054,In_358,In_148);
xor U4055 (N_4055,In_257,In_922);
xor U4056 (N_4056,In_245,In_155);
xnor U4057 (N_4057,In_419,In_817);
nand U4058 (N_4058,In_383,In_818);
or U4059 (N_4059,In_464,In_787);
nor U4060 (N_4060,In_801,In_894);
xor U4061 (N_4061,In_621,In_4);
and U4062 (N_4062,In_162,In_145);
or U4063 (N_4063,In_504,In_732);
or U4064 (N_4064,In_367,In_551);
xor U4065 (N_4065,In_945,In_179);
nor U4066 (N_4066,In_796,In_134);
and U4067 (N_4067,In_934,In_412);
or U4068 (N_4068,In_301,In_671);
and U4069 (N_4069,In_454,In_431);
and U4070 (N_4070,In_766,In_674);
or U4071 (N_4071,In_456,In_819);
or U4072 (N_4072,In_170,In_914);
or U4073 (N_4073,In_19,In_890);
nand U4074 (N_4074,In_359,In_353);
nand U4075 (N_4075,In_718,In_59);
and U4076 (N_4076,In_993,In_367);
nor U4077 (N_4077,In_920,In_892);
or U4078 (N_4078,In_736,In_433);
xnor U4079 (N_4079,In_871,In_217);
and U4080 (N_4080,In_35,In_37);
nand U4081 (N_4081,In_765,In_883);
nand U4082 (N_4082,In_938,In_512);
and U4083 (N_4083,In_385,In_835);
nor U4084 (N_4084,In_254,In_834);
and U4085 (N_4085,In_252,In_148);
nand U4086 (N_4086,In_789,In_275);
and U4087 (N_4087,In_470,In_915);
and U4088 (N_4088,In_904,In_445);
nand U4089 (N_4089,In_933,In_720);
nand U4090 (N_4090,In_194,In_229);
xnor U4091 (N_4091,In_882,In_251);
or U4092 (N_4092,In_232,In_418);
xor U4093 (N_4093,In_196,In_88);
nand U4094 (N_4094,In_356,In_612);
xnor U4095 (N_4095,In_151,In_83);
and U4096 (N_4096,In_278,In_13);
xnor U4097 (N_4097,In_503,In_184);
and U4098 (N_4098,In_997,In_680);
nand U4099 (N_4099,In_793,In_587);
or U4100 (N_4100,In_193,In_26);
nor U4101 (N_4101,In_239,In_810);
nor U4102 (N_4102,In_598,In_98);
nor U4103 (N_4103,In_436,In_616);
nor U4104 (N_4104,In_81,In_943);
nand U4105 (N_4105,In_143,In_563);
nor U4106 (N_4106,In_915,In_302);
nor U4107 (N_4107,In_851,In_558);
nand U4108 (N_4108,In_201,In_540);
nor U4109 (N_4109,In_211,In_533);
nand U4110 (N_4110,In_867,In_173);
or U4111 (N_4111,In_709,In_132);
and U4112 (N_4112,In_974,In_912);
nand U4113 (N_4113,In_481,In_252);
nand U4114 (N_4114,In_965,In_642);
xnor U4115 (N_4115,In_198,In_289);
and U4116 (N_4116,In_440,In_311);
and U4117 (N_4117,In_533,In_331);
nand U4118 (N_4118,In_552,In_711);
or U4119 (N_4119,In_317,In_364);
nor U4120 (N_4120,In_930,In_295);
or U4121 (N_4121,In_202,In_8);
or U4122 (N_4122,In_29,In_529);
xor U4123 (N_4123,In_444,In_585);
nor U4124 (N_4124,In_369,In_185);
or U4125 (N_4125,In_747,In_311);
and U4126 (N_4126,In_585,In_367);
or U4127 (N_4127,In_914,In_895);
xnor U4128 (N_4128,In_916,In_545);
nand U4129 (N_4129,In_13,In_9);
xor U4130 (N_4130,In_85,In_145);
or U4131 (N_4131,In_256,In_106);
and U4132 (N_4132,In_271,In_985);
nor U4133 (N_4133,In_206,In_954);
or U4134 (N_4134,In_594,In_412);
xor U4135 (N_4135,In_826,In_821);
or U4136 (N_4136,In_537,In_985);
nor U4137 (N_4137,In_740,In_195);
and U4138 (N_4138,In_471,In_55);
nand U4139 (N_4139,In_177,In_651);
xnor U4140 (N_4140,In_446,In_842);
nand U4141 (N_4141,In_891,In_511);
nor U4142 (N_4142,In_374,In_76);
or U4143 (N_4143,In_962,In_696);
or U4144 (N_4144,In_617,In_897);
nor U4145 (N_4145,In_152,In_853);
nand U4146 (N_4146,In_18,In_242);
or U4147 (N_4147,In_79,In_203);
or U4148 (N_4148,In_435,In_966);
and U4149 (N_4149,In_6,In_605);
or U4150 (N_4150,In_788,In_951);
or U4151 (N_4151,In_705,In_82);
or U4152 (N_4152,In_680,In_459);
and U4153 (N_4153,In_623,In_108);
nor U4154 (N_4154,In_131,In_938);
nor U4155 (N_4155,In_273,In_172);
xnor U4156 (N_4156,In_15,In_158);
nand U4157 (N_4157,In_763,In_234);
or U4158 (N_4158,In_930,In_194);
nor U4159 (N_4159,In_38,In_336);
nor U4160 (N_4160,In_988,In_321);
or U4161 (N_4161,In_262,In_803);
nand U4162 (N_4162,In_944,In_317);
xor U4163 (N_4163,In_661,In_256);
nand U4164 (N_4164,In_404,In_214);
nand U4165 (N_4165,In_485,In_573);
or U4166 (N_4166,In_194,In_653);
or U4167 (N_4167,In_907,In_370);
nand U4168 (N_4168,In_485,In_420);
or U4169 (N_4169,In_440,In_675);
nand U4170 (N_4170,In_208,In_953);
nor U4171 (N_4171,In_262,In_1);
nor U4172 (N_4172,In_867,In_203);
nand U4173 (N_4173,In_542,In_884);
nand U4174 (N_4174,In_15,In_335);
or U4175 (N_4175,In_994,In_272);
xnor U4176 (N_4176,In_978,In_281);
and U4177 (N_4177,In_938,In_416);
xnor U4178 (N_4178,In_750,In_996);
nand U4179 (N_4179,In_309,In_982);
or U4180 (N_4180,In_534,In_233);
xnor U4181 (N_4181,In_680,In_223);
or U4182 (N_4182,In_116,In_909);
xnor U4183 (N_4183,In_614,In_910);
or U4184 (N_4184,In_29,In_166);
and U4185 (N_4185,In_916,In_548);
nand U4186 (N_4186,In_966,In_546);
xor U4187 (N_4187,In_781,In_230);
nand U4188 (N_4188,In_820,In_953);
or U4189 (N_4189,In_732,In_389);
and U4190 (N_4190,In_422,In_160);
xor U4191 (N_4191,In_36,In_421);
nor U4192 (N_4192,In_951,In_796);
or U4193 (N_4193,In_796,In_757);
and U4194 (N_4194,In_946,In_154);
and U4195 (N_4195,In_389,In_31);
nor U4196 (N_4196,In_137,In_267);
or U4197 (N_4197,In_47,In_655);
nand U4198 (N_4198,In_532,In_395);
nor U4199 (N_4199,In_456,In_770);
nor U4200 (N_4200,In_554,In_475);
or U4201 (N_4201,In_38,In_544);
nor U4202 (N_4202,In_32,In_872);
nor U4203 (N_4203,In_265,In_323);
nand U4204 (N_4204,In_143,In_157);
or U4205 (N_4205,In_204,In_920);
or U4206 (N_4206,In_395,In_356);
and U4207 (N_4207,In_157,In_652);
nor U4208 (N_4208,In_684,In_284);
nand U4209 (N_4209,In_464,In_113);
xnor U4210 (N_4210,In_673,In_91);
xnor U4211 (N_4211,In_905,In_44);
nand U4212 (N_4212,In_888,In_410);
and U4213 (N_4213,In_7,In_803);
xor U4214 (N_4214,In_175,In_694);
xor U4215 (N_4215,In_221,In_120);
and U4216 (N_4216,In_622,In_110);
nand U4217 (N_4217,In_664,In_416);
or U4218 (N_4218,In_736,In_737);
nor U4219 (N_4219,In_701,In_652);
nor U4220 (N_4220,In_145,In_931);
or U4221 (N_4221,In_438,In_281);
and U4222 (N_4222,In_801,In_876);
or U4223 (N_4223,In_770,In_469);
or U4224 (N_4224,In_882,In_318);
and U4225 (N_4225,In_208,In_755);
and U4226 (N_4226,In_304,In_714);
and U4227 (N_4227,In_809,In_786);
xnor U4228 (N_4228,In_874,In_409);
or U4229 (N_4229,In_606,In_655);
nor U4230 (N_4230,In_627,In_50);
nor U4231 (N_4231,In_619,In_197);
nand U4232 (N_4232,In_583,In_605);
xor U4233 (N_4233,In_485,In_272);
nand U4234 (N_4234,In_435,In_57);
or U4235 (N_4235,In_711,In_434);
nor U4236 (N_4236,In_402,In_945);
nand U4237 (N_4237,In_936,In_454);
and U4238 (N_4238,In_788,In_857);
nor U4239 (N_4239,In_697,In_973);
xnor U4240 (N_4240,In_775,In_520);
nand U4241 (N_4241,In_672,In_23);
xor U4242 (N_4242,In_417,In_618);
nor U4243 (N_4243,In_207,In_26);
nor U4244 (N_4244,In_744,In_190);
nor U4245 (N_4245,In_497,In_274);
xor U4246 (N_4246,In_853,In_217);
xor U4247 (N_4247,In_681,In_317);
nor U4248 (N_4248,In_984,In_855);
or U4249 (N_4249,In_365,In_19);
nand U4250 (N_4250,In_618,In_35);
and U4251 (N_4251,In_645,In_292);
xnor U4252 (N_4252,In_542,In_209);
or U4253 (N_4253,In_652,In_937);
or U4254 (N_4254,In_175,In_880);
and U4255 (N_4255,In_849,In_233);
or U4256 (N_4256,In_393,In_933);
nand U4257 (N_4257,In_57,In_262);
xnor U4258 (N_4258,In_996,In_288);
nand U4259 (N_4259,In_820,In_232);
nand U4260 (N_4260,In_515,In_236);
xor U4261 (N_4261,In_421,In_259);
xor U4262 (N_4262,In_869,In_383);
and U4263 (N_4263,In_141,In_32);
nor U4264 (N_4264,In_57,In_833);
and U4265 (N_4265,In_90,In_885);
and U4266 (N_4266,In_603,In_121);
nand U4267 (N_4267,In_961,In_102);
or U4268 (N_4268,In_54,In_132);
nor U4269 (N_4269,In_201,In_669);
or U4270 (N_4270,In_537,In_358);
xnor U4271 (N_4271,In_220,In_647);
xor U4272 (N_4272,In_164,In_543);
xnor U4273 (N_4273,In_427,In_208);
nor U4274 (N_4274,In_668,In_813);
and U4275 (N_4275,In_794,In_849);
nor U4276 (N_4276,In_986,In_436);
and U4277 (N_4277,In_805,In_636);
nor U4278 (N_4278,In_666,In_692);
xnor U4279 (N_4279,In_686,In_476);
or U4280 (N_4280,In_508,In_136);
or U4281 (N_4281,In_777,In_603);
nand U4282 (N_4282,In_929,In_766);
nor U4283 (N_4283,In_937,In_409);
xnor U4284 (N_4284,In_871,In_996);
xor U4285 (N_4285,In_35,In_569);
nor U4286 (N_4286,In_679,In_617);
nor U4287 (N_4287,In_201,In_526);
nand U4288 (N_4288,In_334,In_903);
xor U4289 (N_4289,In_647,In_466);
xor U4290 (N_4290,In_560,In_600);
or U4291 (N_4291,In_179,In_927);
nand U4292 (N_4292,In_580,In_322);
nor U4293 (N_4293,In_516,In_606);
xnor U4294 (N_4294,In_374,In_197);
nand U4295 (N_4295,In_603,In_934);
or U4296 (N_4296,In_777,In_396);
nor U4297 (N_4297,In_595,In_822);
and U4298 (N_4298,In_743,In_863);
and U4299 (N_4299,In_74,In_422);
and U4300 (N_4300,In_970,In_844);
or U4301 (N_4301,In_977,In_803);
nor U4302 (N_4302,In_795,In_111);
or U4303 (N_4303,In_171,In_932);
nor U4304 (N_4304,In_394,In_355);
xnor U4305 (N_4305,In_124,In_982);
nand U4306 (N_4306,In_56,In_901);
and U4307 (N_4307,In_516,In_791);
or U4308 (N_4308,In_635,In_848);
xnor U4309 (N_4309,In_65,In_902);
or U4310 (N_4310,In_928,In_309);
and U4311 (N_4311,In_816,In_973);
nand U4312 (N_4312,In_249,In_221);
or U4313 (N_4313,In_636,In_368);
and U4314 (N_4314,In_530,In_11);
nor U4315 (N_4315,In_730,In_307);
nand U4316 (N_4316,In_673,In_400);
xnor U4317 (N_4317,In_941,In_199);
xor U4318 (N_4318,In_787,In_793);
xor U4319 (N_4319,In_654,In_662);
nor U4320 (N_4320,In_155,In_236);
nor U4321 (N_4321,In_14,In_457);
or U4322 (N_4322,In_443,In_468);
xnor U4323 (N_4323,In_502,In_436);
and U4324 (N_4324,In_120,In_187);
or U4325 (N_4325,In_684,In_279);
nand U4326 (N_4326,In_470,In_456);
nand U4327 (N_4327,In_558,In_924);
nand U4328 (N_4328,In_405,In_557);
nor U4329 (N_4329,In_671,In_609);
xnor U4330 (N_4330,In_798,In_887);
nor U4331 (N_4331,In_71,In_269);
and U4332 (N_4332,In_480,In_590);
nand U4333 (N_4333,In_403,In_979);
nor U4334 (N_4334,In_75,In_667);
and U4335 (N_4335,In_161,In_59);
nor U4336 (N_4336,In_191,In_101);
or U4337 (N_4337,In_228,In_301);
nand U4338 (N_4338,In_105,In_944);
nor U4339 (N_4339,In_168,In_74);
xnor U4340 (N_4340,In_260,In_146);
or U4341 (N_4341,In_511,In_271);
nor U4342 (N_4342,In_717,In_568);
nor U4343 (N_4343,In_857,In_532);
or U4344 (N_4344,In_332,In_408);
or U4345 (N_4345,In_929,In_264);
or U4346 (N_4346,In_899,In_474);
nor U4347 (N_4347,In_610,In_724);
nand U4348 (N_4348,In_46,In_47);
nor U4349 (N_4349,In_433,In_222);
and U4350 (N_4350,In_893,In_635);
or U4351 (N_4351,In_645,In_788);
or U4352 (N_4352,In_92,In_745);
or U4353 (N_4353,In_133,In_668);
nand U4354 (N_4354,In_284,In_188);
and U4355 (N_4355,In_801,In_879);
nor U4356 (N_4356,In_895,In_865);
nand U4357 (N_4357,In_706,In_666);
xor U4358 (N_4358,In_673,In_648);
nand U4359 (N_4359,In_701,In_670);
and U4360 (N_4360,In_453,In_437);
nor U4361 (N_4361,In_978,In_371);
nand U4362 (N_4362,In_596,In_643);
or U4363 (N_4363,In_688,In_947);
or U4364 (N_4364,In_728,In_447);
and U4365 (N_4365,In_892,In_699);
nor U4366 (N_4366,In_936,In_193);
and U4367 (N_4367,In_936,In_202);
or U4368 (N_4368,In_317,In_665);
nor U4369 (N_4369,In_625,In_317);
and U4370 (N_4370,In_256,In_4);
nand U4371 (N_4371,In_125,In_980);
xor U4372 (N_4372,In_463,In_947);
xnor U4373 (N_4373,In_825,In_860);
nor U4374 (N_4374,In_193,In_531);
and U4375 (N_4375,In_892,In_886);
nor U4376 (N_4376,In_160,In_236);
nand U4377 (N_4377,In_126,In_388);
xnor U4378 (N_4378,In_901,In_760);
nor U4379 (N_4379,In_891,In_787);
or U4380 (N_4380,In_281,In_505);
nand U4381 (N_4381,In_17,In_953);
and U4382 (N_4382,In_47,In_904);
or U4383 (N_4383,In_979,In_958);
xnor U4384 (N_4384,In_804,In_377);
xor U4385 (N_4385,In_351,In_474);
xnor U4386 (N_4386,In_737,In_445);
xnor U4387 (N_4387,In_234,In_534);
and U4388 (N_4388,In_149,In_927);
nand U4389 (N_4389,In_358,In_634);
xnor U4390 (N_4390,In_378,In_905);
and U4391 (N_4391,In_665,In_886);
and U4392 (N_4392,In_821,In_378);
nor U4393 (N_4393,In_161,In_33);
nor U4394 (N_4394,In_566,In_449);
and U4395 (N_4395,In_237,In_555);
nor U4396 (N_4396,In_753,In_266);
nand U4397 (N_4397,In_840,In_88);
xnor U4398 (N_4398,In_312,In_290);
and U4399 (N_4399,In_976,In_505);
xor U4400 (N_4400,In_206,In_823);
nand U4401 (N_4401,In_899,In_589);
or U4402 (N_4402,In_202,In_685);
or U4403 (N_4403,In_61,In_241);
and U4404 (N_4404,In_597,In_784);
nor U4405 (N_4405,In_43,In_933);
nor U4406 (N_4406,In_42,In_884);
xnor U4407 (N_4407,In_62,In_566);
nand U4408 (N_4408,In_952,In_518);
or U4409 (N_4409,In_606,In_462);
nor U4410 (N_4410,In_617,In_397);
nand U4411 (N_4411,In_758,In_569);
nand U4412 (N_4412,In_948,In_710);
nand U4413 (N_4413,In_928,In_92);
and U4414 (N_4414,In_989,In_934);
nand U4415 (N_4415,In_784,In_564);
and U4416 (N_4416,In_840,In_955);
xnor U4417 (N_4417,In_95,In_930);
and U4418 (N_4418,In_370,In_636);
or U4419 (N_4419,In_444,In_879);
nor U4420 (N_4420,In_318,In_874);
or U4421 (N_4421,In_744,In_106);
xnor U4422 (N_4422,In_678,In_694);
and U4423 (N_4423,In_246,In_774);
nand U4424 (N_4424,In_91,In_778);
nor U4425 (N_4425,In_828,In_785);
and U4426 (N_4426,In_600,In_947);
and U4427 (N_4427,In_996,In_334);
and U4428 (N_4428,In_710,In_875);
and U4429 (N_4429,In_187,In_371);
and U4430 (N_4430,In_936,In_525);
nand U4431 (N_4431,In_258,In_777);
nor U4432 (N_4432,In_343,In_68);
xor U4433 (N_4433,In_864,In_270);
or U4434 (N_4434,In_865,In_544);
or U4435 (N_4435,In_314,In_434);
xor U4436 (N_4436,In_26,In_574);
and U4437 (N_4437,In_53,In_201);
xor U4438 (N_4438,In_422,In_951);
and U4439 (N_4439,In_519,In_234);
xor U4440 (N_4440,In_961,In_854);
xnor U4441 (N_4441,In_871,In_890);
and U4442 (N_4442,In_662,In_262);
or U4443 (N_4443,In_775,In_995);
or U4444 (N_4444,In_538,In_22);
xnor U4445 (N_4445,In_815,In_30);
nor U4446 (N_4446,In_680,In_943);
and U4447 (N_4447,In_591,In_613);
xnor U4448 (N_4448,In_325,In_927);
and U4449 (N_4449,In_165,In_340);
nor U4450 (N_4450,In_442,In_734);
and U4451 (N_4451,In_333,In_714);
nand U4452 (N_4452,In_645,In_77);
nor U4453 (N_4453,In_106,In_676);
nor U4454 (N_4454,In_666,In_204);
nor U4455 (N_4455,In_463,In_661);
xnor U4456 (N_4456,In_289,In_227);
xnor U4457 (N_4457,In_577,In_614);
nor U4458 (N_4458,In_915,In_893);
or U4459 (N_4459,In_34,In_16);
nor U4460 (N_4460,In_60,In_919);
nor U4461 (N_4461,In_315,In_764);
and U4462 (N_4462,In_939,In_973);
nand U4463 (N_4463,In_408,In_908);
nor U4464 (N_4464,In_432,In_869);
xor U4465 (N_4465,In_846,In_908);
and U4466 (N_4466,In_902,In_875);
nor U4467 (N_4467,In_755,In_26);
nor U4468 (N_4468,In_699,In_898);
xor U4469 (N_4469,In_852,In_867);
nand U4470 (N_4470,In_671,In_326);
xnor U4471 (N_4471,In_318,In_820);
nor U4472 (N_4472,In_823,In_990);
and U4473 (N_4473,In_154,In_368);
and U4474 (N_4474,In_724,In_845);
xor U4475 (N_4475,In_146,In_827);
nand U4476 (N_4476,In_51,In_701);
or U4477 (N_4477,In_247,In_113);
xor U4478 (N_4478,In_970,In_44);
and U4479 (N_4479,In_633,In_248);
nor U4480 (N_4480,In_245,In_800);
nand U4481 (N_4481,In_632,In_116);
nand U4482 (N_4482,In_223,In_43);
nand U4483 (N_4483,In_518,In_587);
xnor U4484 (N_4484,In_572,In_373);
nand U4485 (N_4485,In_12,In_869);
nand U4486 (N_4486,In_327,In_697);
nand U4487 (N_4487,In_269,In_822);
and U4488 (N_4488,In_859,In_643);
nand U4489 (N_4489,In_760,In_415);
or U4490 (N_4490,In_439,In_258);
and U4491 (N_4491,In_938,In_32);
xor U4492 (N_4492,In_941,In_954);
xnor U4493 (N_4493,In_910,In_144);
xnor U4494 (N_4494,In_893,In_722);
and U4495 (N_4495,In_115,In_204);
xor U4496 (N_4496,In_784,In_890);
and U4497 (N_4497,In_218,In_243);
and U4498 (N_4498,In_924,In_806);
and U4499 (N_4499,In_345,In_249);
and U4500 (N_4500,In_90,In_274);
xor U4501 (N_4501,In_902,In_353);
xnor U4502 (N_4502,In_440,In_93);
xnor U4503 (N_4503,In_699,In_700);
or U4504 (N_4504,In_476,In_941);
xor U4505 (N_4505,In_196,In_69);
or U4506 (N_4506,In_968,In_661);
nor U4507 (N_4507,In_940,In_263);
or U4508 (N_4508,In_572,In_154);
or U4509 (N_4509,In_759,In_741);
xnor U4510 (N_4510,In_206,In_292);
or U4511 (N_4511,In_41,In_522);
nand U4512 (N_4512,In_42,In_892);
and U4513 (N_4513,In_802,In_937);
nor U4514 (N_4514,In_331,In_748);
and U4515 (N_4515,In_810,In_921);
nor U4516 (N_4516,In_761,In_334);
nor U4517 (N_4517,In_466,In_816);
xnor U4518 (N_4518,In_67,In_760);
nand U4519 (N_4519,In_741,In_941);
xnor U4520 (N_4520,In_909,In_166);
nand U4521 (N_4521,In_682,In_431);
and U4522 (N_4522,In_512,In_156);
and U4523 (N_4523,In_36,In_343);
nor U4524 (N_4524,In_723,In_200);
xnor U4525 (N_4525,In_122,In_781);
nor U4526 (N_4526,In_23,In_282);
or U4527 (N_4527,In_491,In_155);
nor U4528 (N_4528,In_200,In_1);
nand U4529 (N_4529,In_528,In_163);
xnor U4530 (N_4530,In_288,In_959);
and U4531 (N_4531,In_281,In_640);
or U4532 (N_4532,In_204,In_279);
nand U4533 (N_4533,In_417,In_718);
or U4534 (N_4534,In_339,In_102);
xor U4535 (N_4535,In_268,In_366);
nor U4536 (N_4536,In_387,In_178);
or U4537 (N_4537,In_114,In_963);
or U4538 (N_4538,In_171,In_227);
nor U4539 (N_4539,In_380,In_941);
or U4540 (N_4540,In_699,In_380);
nand U4541 (N_4541,In_525,In_186);
and U4542 (N_4542,In_995,In_532);
xnor U4543 (N_4543,In_1,In_25);
nor U4544 (N_4544,In_468,In_445);
or U4545 (N_4545,In_122,In_142);
xnor U4546 (N_4546,In_48,In_479);
or U4547 (N_4547,In_90,In_268);
and U4548 (N_4548,In_737,In_507);
xor U4549 (N_4549,In_741,In_185);
or U4550 (N_4550,In_927,In_597);
nand U4551 (N_4551,In_181,In_613);
and U4552 (N_4552,In_987,In_358);
nor U4553 (N_4553,In_677,In_300);
and U4554 (N_4554,In_98,In_328);
nand U4555 (N_4555,In_991,In_132);
nand U4556 (N_4556,In_932,In_176);
or U4557 (N_4557,In_48,In_958);
or U4558 (N_4558,In_574,In_537);
or U4559 (N_4559,In_473,In_106);
nand U4560 (N_4560,In_828,In_356);
or U4561 (N_4561,In_257,In_727);
xor U4562 (N_4562,In_795,In_870);
or U4563 (N_4563,In_496,In_772);
xor U4564 (N_4564,In_869,In_436);
nor U4565 (N_4565,In_27,In_132);
nor U4566 (N_4566,In_547,In_168);
or U4567 (N_4567,In_10,In_645);
xor U4568 (N_4568,In_683,In_620);
or U4569 (N_4569,In_249,In_189);
or U4570 (N_4570,In_834,In_272);
nor U4571 (N_4571,In_204,In_513);
nor U4572 (N_4572,In_313,In_936);
and U4573 (N_4573,In_436,In_335);
nor U4574 (N_4574,In_342,In_354);
or U4575 (N_4575,In_984,In_414);
or U4576 (N_4576,In_809,In_64);
xnor U4577 (N_4577,In_525,In_597);
and U4578 (N_4578,In_729,In_861);
or U4579 (N_4579,In_589,In_332);
nor U4580 (N_4580,In_109,In_411);
and U4581 (N_4581,In_965,In_539);
and U4582 (N_4582,In_998,In_792);
and U4583 (N_4583,In_434,In_768);
and U4584 (N_4584,In_764,In_775);
nand U4585 (N_4585,In_560,In_747);
and U4586 (N_4586,In_175,In_973);
xor U4587 (N_4587,In_2,In_302);
xor U4588 (N_4588,In_305,In_379);
and U4589 (N_4589,In_190,In_517);
nor U4590 (N_4590,In_794,In_662);
nand U4591 (N_4591,In_826,In_642);
xnor U4592 (N_4592,In_986,In_843);
nand U4593 (N_4593,In_313,In_771);
xnor U4594 (N_4594,In_256,In_939);
nor U4595 (N_4595,In_658,In_896);
xor U4596 (N_4596,In_328,In_621);
xor U4597 (N_4597,In_253,In_266);
nor U4598 (N_4598,In_426,In_856);
nand U4599 (N_4599,In_55,In_865);
or U4600 (N_4600,In_810,In_343);
or U4601 (N_4601,In_905,In_273);
and U4602 (N_4602,In_355,In_957);
and U4603 (N_4603,In_940,In_228);
and U4604 (N_4604,In_650,In_788);
and U4605 (N_4605,In_764,In_992);
or U4606 (N_4606,In_72,In_418);
and U4607 (N_4607,In_77,In_300);
and U4608 (N_4608,In_658,In_575);
xor U4609 (N_4609,In_925,In_220);
or U4610 (N_4610,In_832,In_516);
or U4611 (N_4611,In_912,In_930);
and U4612 (N_4612,In_388,In_961);
or U4613 (N_4613,In_629,In_618);
nand U4614 (N_4614,In_649,In_46);
nand U4615 (N_4615,In_176,In_714);
nor U4616 (N_4616,In_941,In_321);
xor U4617 (N_4617,In_308,In_752);
nor U4618 (N_4618,In_266,In_435);
xor U4619 (N_4619,In_986,In_31);
nor U4620 (N_4620,In_33,In_103);
or U4621 (N_4621,In_846,In_961);
nand U4622 (N_4622,In_334,In_712);
and U4623 (N_4623,In_409,In_538);
or U4624 (N_4624,In_542,In_533);
nand U4625 (N_4625,In_49,In_780);
and U4626 (N_4626,In_268,In_844);
nand U4627 (N_4627,In_218,In_395);
or U4628 (N_4628,In_942,In_437);
xor U4629 (N_4629,In_851,In_776);
xnor U4630 (N_4630,In_760,In_8);
nor U4631 (N_4631,In_128,In_81);
nor U4632 (N_4632,In_975,In_652);
or U4633 (N_4633,In_548,In_630);
nand U4634 (N_4634,In_415,In_581);
xnor U4635 (N_4635,In_303,In_136);
nand U4636 (N_4636,In_37,In_268);
nand U4637 (N_4637,In_141,In_212);
or U4638 (N_4638,In_216,In_359);
nor U4639 (N_4639,In_161,In_302);
nand U4640 (N_4640,In_844,In_328);
nor U4641 (N_4641,In_510,In_132);
nor U4642 (N_4642,In_348,In_770);
xnor U4643 (N_4643,In_3,In_968);
and U4644 (N_4644,In_435,In_562);
nor U4645 (N_4645,In_471,In_56);
or U4646 (N_4646,In_513,In_913);
nor U4647 (N_4647,In_902,In_977);
xnor U4648 (N_4648,In_134,In_907);
and U4649 (N_4649,In_438,In_749);
xor U4650 (N_4650,In_66,In_244);
and U4651 (N_4651,In_542,In_592);
and U4652 (N_4652,In_217,In_222);
or U4653 (N_4653,In_778,In_499);
nor U4654 (N_4654,In_806,In_334);
nor U4655 (N_4655,In_817,In_252);
xor U4656 (N_4656,In_784,In_984);
xnor U4657 (N_4657,In_790,In_678);
xor U4658 (N_4658,In_666,In_106);
nand U4659 (N_4659,In_939,In_343);
and U4660 (N_4660,In_278,In_931);
nor U4661 (N_4661,In_536,In_540);
and U4662 (N_4662,In_348,In_691);
xnor U4663 (N_4663,In_965,In_401);
and U4664 (N_4664,In_517,In_687);
nand U4665 (N_4665,In_632,In_519);
nand U4666 (N_4666,In_801,In_851);
xor U4667 (N_4667,In_120,In_102);
or U4668 (N_4668,In_460,In_225);
and U4669 (N_4669,In_78,In_984);
or U4670 (N_4670,In_479,In_788);
xor U4671 (N_4671,In_124,In_536);
or U4672 (N_4672,In_977,In_669);
xnor U4673 (N_4673,In_970,In_396);
xor U4674 (N_4674,In_344,In_507);
or U4675 (N_4675,In_688,In_371);
or U4676 (N_4676,In_917,In_729);
or U4677 (N_4677,In_687,In_258);
nand U4678 (N_4678,In_41,In_285);
nor U4679 (N_4679,In_65,In_188);
xor U4680 (N_4680,In_702,In_746);
xor U4681 (N_4681,In_24,In_382);
nor U4682 (N_4682,In_722,In_225);
xor U4683 (N_4683,In_78,In_22);
and U4684 (N_4684,In_713,In_780);
nand U4685 (N_4685,In_110,In_589);
xor U4686 (N_4686,In_51,In_420);
and U4687 (N_4687,In_546,In_984);
xnor U4688 (N_4688,In_427,In_815);
xnor U4689 (N_4689,In_947,In_647);
xor U4690 (N_4690,In_251,In_514);
nand U4691 (N_4691,In_267,In_959);
and U4692 (N_4692,In_988,In_680);
xnor U4693 (N_4693,In_644,In_227);
nand U4694 (N_4694,In_610,In_763);
nor U4695 (N_4695,In_4,In_892);
or U4696 (N_4696,In_780,In_810);
nand U4697 (N_4697,In_898,In_355);
nand U4698 (N_4698,In_608,In_89);
nor U4699 (N_4699,In_658,In_140);
nand U4700 (N_4700,In_222,In_765);
and U4701 (N_4701,In_703,In_432);
xnor U4702 (N_4702,In_855,In_840);
nor U4703 (N_4703,In_271,In_732);
or U4704 (N_4704,In_435,In_694);
nor U4705 (N_4705,In_634,In_659);
nor U4706 (N_4706,In_30,In_226);
and U4707 (N_4707,In_641,In_119);
and U4708 (N_4708,In_718,In_357);
nand U4709 (N_4709,In_360,In_283);
and U4710 (N_4710,In_941,In_319);
nor U4711 (N_4711,In_346,In_699);
nand U4712 (N_4712,In_200,In_679);
xor U4713 (N_4713,In_353,In_753);
nor U4714 (N_4714,In_427,In_898);
or U4715 (N_4715,In_478,In_643);
nand U4716 (N_4716,In_195,In_330);
and U4717 (N_4717,In_102,In_973);
and U4718 (N_4718,In_796,In_316);
nand U4719 (N_4719,In_165,In_774);
xnor U4720 (N_4720,In_816,In_203);
nand U4721 (N_4721,In_854,In_871);
or U4722 (N_4722,In_917,In_441);
and U4723 (N_4723,In_528,In_948);
xor U4724 (N_4724,In_566,In_427);
xnor U4725 (N_4725,In_580,In_775);
and U4726 (N_4726,In_839,In_798);
nor U4727 (N_4727,In_269,In_100);
nor U4728 (N_4728,In_218,In_793);
nor U4729 (N_4729,In_583,In_302);
xnor U4730 (N_4730,In_663,In_832);
and U4731 (N_4731,In_421,In_90);
and U4732 (N_4732,In_605,In_242);
and U4733 (N_4733,In_960,In_211);
nand U4734 (N_4734,In_253,In_166);
or U4735 (N_4735,In_8,In_655);
xnor U4736 (N_4736,In_318,In_559);
nor U4737 (N_4737,In_786,In_246);
nor U4738 (N_4738,In_307,In_770);
nor U4739 (N_4739,In_663,In_490);
or U4740 (N_4740,In_321,In_965);
or U4741 (N_4741,In_880,In_249);
xor U4742 (N_4742,In_70,In_248);
nor U4743 (N_4743,In_58,In_208);
or U4744 (N_4744,In_975,In_219);
nand U4745 (N_4745,In_912,In_154);
xor U4746 (N_4746,In_406,In_78);
nand U4747 (N_4747,In_429,In_602);
xor U4748 (N_4748,In_922,In_556);
or U4749 (N_4749,In_756,In_773);
and U4750 (N_4750,In_105,In_295);
and U4751 (N_4751,In_235,In_799);
nand U4752 (N_4752,In_9,In_804);
nor U4753 (N_4753,In_108,In_460);
nor U4754 (N_4754,In_92,In_220);
nand U4755 (N_4755,In_73,In_181);
and U4756 (N_4756,In_602,In_795);
and U4757 (N_4757,In_77,In_577);
nor U4758 (N_4758,In_654,In_39);
nor U4759 (N_4759,In_403,In_599);
and U4760 (N_4760,In_346,In_719);
nand U4761 (N_4761,In_450,In_70);
nor U4762 (N_4762,In_554,In_882);
nand U4763 (N_4763,In_731,In_506);
or U4764 (N_4764,In_136,In_481);
xnor U4765 (N_4765,In_99,In_968);
or U4766 (N_4766,In_505,In_974);
and U4767 (N_4767,In_216,In_471);
xor U4768 (N_4768,In_560,In_518);
and U4769 (N_4769,In_842,In_946);
or U4770 (N_4770,In_332,In_213);
nand U4771 (N_4771,In_677,In_699);
or U4772 (N_4772,In_213,In_246);
nand U4773 (N_4773,In_861,In_51);
and U4774 (N_4774,In_859,In_152);
and U4775 (N_4775,In_709,In_400);
xnor U4776 (N_4776,In_440,In_45);
nand U4777 (N_4777,In_399,In_97);
nand U4778 (N_4778,In_654,In_822);
nand U4779 (N_4779,In_956,In_697);
or U4780 (N_4780,In_248,In_90);
xor U4781 (N_4781,In_4,In_882);
and U4782 (N_4782,In_425,In_368);
or U4783 (N_4783,In_618,In_213);
xnor U4784 (N_4784,In_193,In_865);
nor U4785 (N_4785,In_63,In_879);
nand U4786 (N_4786,In_434,In_171);
or U4787 (N_4787,In_325,In_816);
and U4788 (N_4788,In_322,In_616);
nor U4789 (N_4789,In_718,In_575);
xor U4790 (N_4790,In_57,In_719);
or U4791 (N_4791,In_350,In_266);
and U4792 (N_4792,In_617,In_458);
nand U4793 (N_4793,In_719,In_902);
xnor U4794 (N_4794,In_150,In_919);
and U4795 (N_4795,In_879,In_971);
nor U4796 (N_4796,In_388,In_19);
or U4797 (N_4797,In_130,In_361);
xnor U4798 (N_4798,In_813,In_323);
xnor U4799 (N_4799,In_614,In_9);
nand U4800 (N_4800,In_251,In_986);
or U4801 (N_4801,In_706,In_484);
nor U4802 (N_4802,In_11,In_137);
xnor U4803 (N_4803,In_463,In_897);
nor U4804 (N_4804,In_615,In_739);
or U4805 (N_4805,In_614,In_422);
and U4806 (N_4806,In_58,In_467);
xor U4807 (N_4807,In_66,In_523);
or U4808 (N_4808,In_459,In_131);
nand U4809 (N_4809,In_378,In_243);
and U4810 (N_4810,In_261,In_809);
xnor U4811 (N_4811,In_869,In_10);
xor U4812 (N_4812,In_734,In_889);
nand U4813 (N_4813,In_961,In_479);
nand U4814 (N_4814,In_120,In_81);
xnor U4815 (N_4815,In_642,In_255);
and U4816 (N_4816,In_734,In_100);
nand U4817 (N_4817,In_40,In_917);
xor U4818 (N_4818,In_395,In_783);
nor U4819 (N_4819,In_11,In_382);
and U4820 (N_4820,In_148,In_247);
and U4821 (N_4821,In_809,In_898);
xnor U4822 (N_4822,In_207,In_580);
xnor U4823 (N_4823,In_650,In_256);
nand U4824 (N_4824,In_108,In_42);
or U4825 (N_4825,In_597,In_909);
xor U4826 (N_4826,In_971,In_146);
nand U4827 (N_4827,In_985,In_557);
or U4828 (N_4828,In_76,In_215);
xor U4829 (N_4829,In_857,In_21);
and U4830 (N_4830,In_484,In_131);
or U4831 (N_4831,In_400,In_940);
nand U4832 (N_4832,In_955,In_789);
nand U4833 (N_4833,In_873,In_178);
or U4834 (N_4834,In_714,In_425);
xor U4835 (N_4835,In_540,In_115);
or U4836 (N_4836,In_7,In_892);
nor U4837 (N_4837,In_135,In_468);
nor U4838 (N_4838,In_584,In_13);
xor U4839 (N_4839,In_733,In_525);
xor U4840 (N_4840,In_615,In_80);
xor U4841 (N_4841,In_368,In_262);
xor U4842 (N_4842,In_922,In_870);
nand U4843 (N_4843,In_420,In_746);
nand U4844 (N_4844,In_191,In_904);
nor U4845 (N_4845,In_277,In_47);
and U4846 (N_4846,In_774,In_483);
nand U4847 (N_4847,In_876,In_371);
nor U4848 (N_4848,In_394,In_404);
and U4849 (N_4849,In_296,In_702);
and U4850 (N_4850,In_146,In_407);
or U4851 (N_4851,In_728,In_289);
xnor U4852 (N_4852,In_790,In_234);
and U4853 (N_4853,In_98,In_902);
and U4854 (N_4854,In_978,In_503);
or U4855 (N_4855,In_783,In_355);
nor U4856 (N_4856,In_139,In_766);
and U4857 (N_4857,In_278,In_356);
or U4858 (N_4858,In_368,In_194);
nor U4859 (N_4859,In_535,In_19);
nor U4860 (N_4860,In_953,In_826);
xnor U4861 (N_4861,In_732,In_928);
nand U4862 (N_4862,In_284,In_74);
or U4863 (N_4863,In_550,In_175);
or U4864 (N_4864,In_168,In_508);
and U4865 (N_4865,In_174,In_362);
xnor U4866 (N_4866,In_216,In_613);
xnor U4867 (N_4867,In_88,In_444);
or U4868 (N_4868,In_487,In_137);
nor U4869 (N_4869,In_733,In_572);
nor U4870 (N_4870,In_758,In_422);
and U4871 (N_4871,In_340,In_467);
nand U4872 (N_4872,In_530,In_393);
nor U4873 (N_4873,In_677,In_702);
or U4874 (N_4874,In_403,In_646);
nand U4875 (N_4875,In_592,In_630);
xnor U4876 (N_4876,In_877,In_993);
nor U4877 (N_4877,In_108,In_724);
or U4878 (N_4878,In_107,In_534);
nor U4879 (N_4879,In_811,In_45);
and U4880 (N_4880,In_149,In_584);
and U4881 (N_4881,In_443,In_560);
nand U4882 (N_4882,In_838,In_163);
nand U4883 (N_4883,In_318,In_227);
or U4884 (N_4884,In_276,In_642);
nand U4885 (N_4885,In_684,In_855);
or U4886 (N_4886,In_244,In_141);
nor U4887 (N_4887,In_427,In_498);
nand U4888 (N_4888,In_76,In_738);
xnor U4889 (N_4889,In_246,In_138);
nor U4890 (N_4890,In_325,In_97);
nand U4891 (N_4891,In_458,In_923);
nand U4892 (N_4892,In_548,In_12);
xor U4893 (N_4893,In_574,In_896);
xor U4894 (N_4894,In_341,In_477);
nor U4895 (N_4895,In_427,In_298);
xor U4896 (N_4896,In_867,In_506);
nor U4897 (N_4897,In_354,In_986);
or U4898 (N_4898,In_856,In_689);
nor U4899 (N_4899,In_428,In_993);
nor U4900 (N_4900,In_217,In_289);
nor U4901 (N_4901,In_186,In_776);
nor U4902 (N_4902,In_430,In_827);
nor U4903 (N_4903,In_474,In_66);
nand U4904 (N_4904,In_233,In_483);
nand U4905 (N_4905,In_843,In_859);
nor U4906 (N_4906,In_889,In_334);
or U4907 (N_4907,In_696,In_266);
and U4908 (N_4908,In_595,In_745);
nor U4909 (N_4909,In_317,In_125);
and U4910 (N_4910,In_771,In_69);
nor U4911 (N_4911,In_458,In_393);
and U4912 (N_4912,In_504,In_930);
nor U4913 (N_4913,In_497,In_215);
xor U4914 (N_4914,In_754,In_704);
nor U4915 (N_4915,In_571,In_640);
nor U4916 (N_4916,In_976,In_301);
or U4917 (N_4917,In_898,In_450);
or U4918 (N_4918,In_45,In_396);
xnor U4919 (N_4919,In_208,In_610);
nor U4920 (N_4920,In_857,In_488);
nor U4921 (N_4921,In_408,In_155);
nor U4922 (N_4922,In_449,In_564);
xnor U4923 (N_4923,In_202,In_336);
xnor U4924 (N_4924,In_176,In_830);
or U4925 (N_4925,In_80,In_70);
or U4926 (N_4926,In_513,In_205);
nand U4927 (N_4927,In_34,In_334);
or U4928 (N_4928,In_328,In_333);
xor U4929 (N_4929,In_807,In_196);
xor U4930 (N_4930,In_96,In_753);
nor U4931 (N_4931,In_492,In_304);
nor U4932 (N_4932,In_721,In_570);
nor U4933 (N_4933,In_252,In_69);
xnor U4934 (N_4934,In_987,In_3);
nor U4935 (N_4935,In_29,In_563);
xor U4936 (N_4936,In_124,In_981);
and U4937 (N_4937,In_323,In_77);
xor U4938 (N_4938,In_81,In_431);
or U4939 (N_4939,In_469,In_823);
or U4940 (N_4940,In_955,In_319);
nand U4941 (N_4941,In_736,In_298);
and U4942 (N_4942,In_912,In_515);
and U4943 (N_4943,In_372,In_96);
nand U4944 (N_4944,In_532,In_432);
or U4945 (N_4945,In_957,In_50);
or U4946 (N_4946,In_239,In_252);
nor U4947 (N_4947,In_694,In_999);
and U4948 (N_4948,In_246,In_237);
and U4949 (N_4949,In_429,In_636);
xnor U4950 (N_4950,In_190,In_456);
xnor U4951 (N_4951,In_221,In_605);
and U4952 (N_4952,In_634,In_460);
or U4953 (N_4953,In_225,In_364);
and U4954 (N_4954,In_112,In_554);
or U4955 (N_4955,In_974,In_481);
or U4956 (N_4956,In_26,In_123);
nand U4957 (N_4957,In_957,In_750);
xor U4958 (N_4958,In_358,In_583);
or U4959 (N_4959,In_871,In_178);
and U4960 (N_4960,In_524,In_997);
nor U4961 (N_4961,In_88,In_806);
and U4962 (N_4962,In_261,In_621);
or U4963 (N_4963,In_618,In_325);
and U4964 (N_4964,In_976,In_785);
or U4965 (N_4965,In_969,In_414);
nand U4966 (N_4966,In_23,In_248);
nor U4967 (N_4967,In_205,In_650);
xor U4968 (N_4968,In_652,In_523);
and U4969 (N_4969,In_225,In_92);
and U4970 (N_4970,In_333,In_372);
nand U4971 (N_4971,In_230,In_764);
xor U4972 (N_4972,In_365,In_289);
xnor U4973 (N_4973,In_337,In_137);
xnor U4974 (N_4974,In_441,In_819);
and U4975 (N_4975,In_936,In_689);
xnor U4976 (N_4976,In_473,In_754);
nand U4977 (N_4977,In_667,In_968);
nand U4978 (N_4978,In_394,In_191);
nor U4979 (N_4979,In_822,In_435);
xor U4980 (N_4980,In_106,In_680);
or U4981 (N_4981,In_319,In_520);
or U4982 (N_4982,In_162,In_630);
or U4983 (N_4983,In_431,In_21);
nor U4984 (N_4984,In_582,In_292);
or U4985 (N_4985,In_536,In_813);
xnor U4986 (N_4986,In_298,In_927);
and U4987 (N_4987,In_394,In_360);
xor U4988 (N_4988,In_297,In_533);
and U4989 (N_4989,In_509,In_91);
or U4990 (N_4990,In_431,In_551);
or U4991 (N_4991,In_343,In_712);
or U4992 (N_4992,In_437,In_767);
nor U4993 (N_4993,In_461,In_134);
or U4994 (N_4994,In_89,In_531);
xnor U4995 (N_4995,In_90,In_536);
nand U4996 (N_4996,In_54,In_863);
or U4997 (N_4997,In_118,In_929);
nor U4998 (N_4998,In_731,In_662);
xnor U4999 (N_4999,In_909,In_273);
nor U5000 (N_5000,N_4017,N_2709);
nor U5001 (N_5001,N_2379,N_1000);
nand U5002 (N_5002,N_3220,N_3725);
xor U5003 (N_5003,N_4040,N_681);
xor U5004 (N_5004,N_836,N_1487);
nor U5005 (N_5005,N_75,N_391);
nor U5006 (N_5006,N_528,N_4671);
and U5007 (N_5007,N_3983,N_1151);
nand U5008 (N_5008,N_273,N_1865);
or U5009 (N_5009,N_2079,N_3146);
nand U5010 (N_5010,N_1166,N_113);
nand U5011 (N_5011,N_850,N_426);
or U5012 (N_5012,N_780,N_1667);
nor U5013 (N_5013,N_3831,N_1163);
xor U5014 (N_5014,N_2319,N_3540);
or U5015 (N_5015,N_2367,N_2559);
xnor U5016 (N_5016,N_2392,N_1748);
and U5017 (N_5017,N_4542,N_4161);
nand U5018 (N_5018,N_4035,N_4014);
nand U5019 (N_5019,N_4759,N_2721);
nor U5020 (N_5020,N_408,N_4493);
nor U5021 (N_5021,N_3187,N_2703);
and U5022 (N_5022,N_4084,N_1822);
or U5023 (N_5023,N_3616,N_3171);
nand U5024 (N_5024,N_3375,N_1564);
xnor U5025 (N_5025,N_2355,N_2714);
xor U5026 (N_5026,N_643,N_131);
nand U5027 (N_5027,N_2269,N_2277);
and U5028 (N_5028,N_1732,N_4038);
and U5029 (N_5029,N_20,N_3521);
and U5030 (N_5030,N_3826,N_3297);
nor U5031 (N_5031,N_1897,N_4162);
xnor U5032 (N_5032,N_1292,N_2739);
nor U5033 (N_5033,N_3541,N_4041);
xnor U5034 (N_5034,N_649,N_4636);
nor U5035 (N_5035,N_2009,N_4332);
nor U5036 (N_5036,N_376,N_1334);
xor U5037 (N_5037,N_2543,N_578);
or U5038 (N_5038,N_3109,N_4496);
and U5039 (N_5039,N_3931,N_3096);
nand U5040 (N_5040,N_2560,N_4186);
or U5041 (N_5041,N_190,N_3288);
and U5042 (N_5042,N_1598,N_999);
xor U5043 (N_5043,N_134,N_3781);
xor U5044 (N_5044,N_4795,N_37);
xnor U5045 (N_5045,N_1825,N_1757);
or U5046 (N_5046,N_2478,N_2592);
or U5047 (N_5047,N_1423,N_1331);
and U5048 (N_5048,N_4103,N_1669);
nand U5049 (N_5049,N_2587,N_4319);
and U5050 (N_5050,N_958,N_1416);
nor U5051 (N_5051,N_4902,N_1880);
or U5052 (N_5052,N_2931,N_2608);
nor U5053 (N_5053,N_3650,N_2964);
and U5054 (N_5054,N_1996,N_2273);
nand U5055 (N_5055,N_4485,N_438);
or U5056 (N_5056,N_2554,N_2737);
or U5057 (N_5057,N_1124,N_3319);
nor U5058 (N_5058,N_1,N_1907);
xnor U5059 (N_5059,N_1447,N_1039);
nor U5060 (N_5060,N_4997,N_4942);
and U5061 (N_5061,N_1122,N_1273);
nand U5062 (N_5062,N_4466,N_825);
nand U5063 (N_5063,N_497,N_2803);
xor U5064 (N_5064,N_3088,N_3859);
or U5065 (N_5065,N_3897,N_339);
xor U5066 (N_5066,N_3480,N_3251);
and U5067 (N_5067,N_4555,N_2087);
nor U5068 (N_5068,N_259,N_4864);
nor U5069 (N_5069,N_1439,N_2762);
or U5070 (N_5070,N_4118,N_87);
xor U5071 (N_5071,N_316,N_900);
nand U5072 (N_5072,N_2730,N_3986);
and U5073 (N_5073,N_493,N_4741);
and U5074 (N_5074,N_806,N_1486);
or U5075 (N_5075,N_2380,N_1235);
nor U5076 (N_5076,N_926,N_4432);
xnor U5077 (N_5077,N_2779,N_4621);
xor U5078 (N_5078,N_4817,N_4700);
nor U5079 (N_5079,N_716,N_1692);
nand U5080 (N_5080,N_2756,N_753);
and U5081 (N_5081,N_1370,N_1280);
nor U5082 (N_5082,N_119,N_4483);
or U5083 (N_5083,N_3179,N_2781);
nand U5084 (N_5084,N_818,N_1206);
nor U5085 (N_5085,N_963,N_4701);
nor U5086 (N_5086,N_1275,N_3399);
xnor U5087 (N_5087,N_2020,N_2274);
nor U5088 (N_5088,N_30,N_3891);
nand U5089 (N_5089,N_1925,N_2580);
and U5090 (N_5090,N_82,N_2778);
nand U5091 (N_5091,N_2664,N_226);
and U5092 (N_5092,N_3531,N_4940);
nand U5093 (N_5093,N_3230,N_3783);
nor U5094 (N_5094,N_3873,N_2589);
or U5095 (N_5095,N_3849,N_821);
nand U5096 (N_5096,N_1726,N_4495);
xor U5097 (N_5097,N_3972,N_3762);
nor U5098 (N_5098,N_4052,N_2825);
or U5099 (N_5099,N_3116,N_651);
and U5100 (N_5100,N_3255,N_1195);
nand U5101 (N_5101,N_2814,N_3680);
nand U5102 (N_5102,N_1856,N_689);
nor U5103 (N_5103,N_873,N_4650);
xor U5104 (N_5104,N_4673,N_1350);
nand U5105 (N_5105,N_2080,N_1159);
and U5106 (N_5106,N_2424,N_1583);
nand U5107 (N_5107,N_4094,N_2045);
nor U5108 (N_5108,N_3684,N_3236);
and U5109 (N_5109,N_4302,N_3430);
nor U5110 (N_5110,N_1218,N_2035);
or U5111 (N_5111,N_2283,N_2887);
xnor U5112 (N_5112,N_851,N_937);
and U5113 (N_5113,N_667,N_2753);
or U5114 (N_5114,N_1332,N_1449);
nand U5115 (N_5115,N_419,N_2783);
nor U5116 (N_5116,N_3393,N_2894);
or U5117 (N_5117,N_1099,N_2883);
xor U5118 (N_5118,N_4210,N_362);
nand U5119 (N_5119,N_3510,N_919);
xor U5120 (N_5120,N_4891,N_2001);
or U5121 (N_5121,N_3271,N_1462);
xor U5122 (N_5122,N_560,N_214);
xor U5123 (N_5123,N_4488,N_3401);
and U5124 (N_5124,N_4919,N_4776);
nor U5125 (N_5125,N_3313,N_155);
nand U5126 (N_5126,N_3615,N_1635);
xor U5127 (N_5127,N_3342,N_4489);
nor U5128 (N_5128,N_787,N_2793);
xor U5129 (N_5129,N_3696,N_3981);
nand U5130 (N_5130,N_2695,N_572);
xor U5131 (N_5131,N_3561,N_601);
and U5132 (N_5132,N_774,N_4175);
nor U5133 (N_5133,N_1860,N_2491);
xnor U5134 (N_5134,N_2909,N_48);
or U5135 (N_5135,N_1857,N_3738);
or U5136 (N_5136,N_3119,N_3155);
or U5137 (N_5137,N_4365,N_3790);
or U5138 (N_5138,N_195,N_3530);
nand U5139 (N_5139,N_3926,N_2575);
nor U5140 (N_5140,N_3069,N_4346);
xor U5141 (N_5141,N_4824,N_1576);
nor U5142 (N_5142,N_538,N_2757);
xor U5143 (N_5143,N_2497,N_1894);
or U5144 (N_5144,N_3045,N_4760);
xnor U5145 (N_5145,N_137,N_1140);
nor U5146 (N_5146,N_2263,N_4949);
nor U5147 (N_5147,N_1797,N_345);
nor U5148 (N_5148,N_3570,N_211);
or U5149 (N_5149,N_2178,N_4096);
or U5150 (N_5150,N_2351,N_2854);
or U5151 (N_5151,N_1468,N_4032);
xnor U5152 (N_5152,N_4178,N_203);
xor U5153 (N_5153,N_1740,N_2493);
xor U5154 (N_5154,N_4648,N_2994);
and U5155 (N_5155,N_1200,N_3678);
nor U5156 (N_5156,N_272,N_3779);
or U5157 (N_5157,N_3161,N_2846);
or U5158 (N_5158,N_109,N_2679);
nand U5159 (N_5159,N_1213,N_3989);
or U5160 (N_5160,N_3285,N_4623);
nand U5161 (N_5161,N_2058,N_432);
and U5162 (N_5162,N_4672,N_3755);
xnor U5163 (N_5163,N_3660,N_4085);
or U5164 (N_5164,N_2605,N_2905);
and U5165 (N_5165,N_182,N_430);
nor U5166 (N_5166,N_1982,N_2595);
nor U5167 (N_5167,N_511,N_2794);
nand U5168 (N_5168,N_1814,N_3511);
xor U5169 (N_5169,N_2717,N_4606);
xnor U5170 (N_5170,N_1677,N_284);
nand U5171 (N_5171,N_2998,N_3265);
or U5172 (N_5172,N_1440,N_3574);
nand U5173 (N_5173,N_1939,N_4237);
nand U5174 (N_5174,N_2089,N_1083);
nor U5175 (N_5175,N_1062,N_4125);
nand U5176 (N_5176,N_2629,N_1067);
and U5177 (N_5177,N_3205,N_4529);
or U5178 (N_5178,N_4472,N_3785);
nor U5179 (N_5179,N_4951,N_3889);
and U5180 (N_5180,N_2397,N_111);
and U5181 (N_5181,N_3331,N_2594);
xor U5182 (N_5182,N_3083,N_3805);
nand U5183 (N_5183,N_1172,N_610);
nor U5184 (N_5184,N_2271,N_4239);
or U5185 (N_5185,N_863,N_4455);
or U5186 (N_5186,N_329,N_4867);
or U5187 (N_5187,N_292,N_3139);
nor U5188 (N_5188,N_635,N_696);
or U5189 (N_5189,N_2667,N_3031);
nand U5190 (N_5190,N_1290,N_287);
nand U5191 (N_5191,N_4163,N_3573);
and U5192 (N_5192,N_4042,N_4301);
nor U5193 (N_5193,N_2201,N_987);
xnor U5194 (N_5194,N_144,N_923);
nand U5195 (N_5195,N_650,N_428);
nor U5196 (N_5196,N_2970,N_2226);
nor U5197 (N_5197,N_3488,N_1176);
nand U5198 (N_5198,N_823,N_658);
or U5199 (N_5199,N_1919,N_3659);
nor U5200 (N_5200,N_1443,N_72);
nand U5201 (N_5201,N_3752,N_97);
nand U5202 (N_5202,N_767,N_3944);
or U5203 (N_5203,N_13,N_4519);
nand U5204 (N_5204,N_185,N_1652);
nor U5205 (N_5205,N_4725,N_2929);
or U5206 (N_5206,N_4266,N_3396);
or U5207 (N_5207,N_1126,N_3671);
nor U5208 (N_5208,N_504,N_1616);
nor U5209 (N_5209,N_1364,N_811);
nand U5210 (N_5210,N_4670,N_314);
or U5211 (N_5211,N_4727,N_2036);
xor U5212 (N_5212,N_359,N_3104);
xor U5213 (N_5213,N_1619,N_2431);
and U5214 (N_5214,N_726,N_1271);
or U5215 (N_5215,N_348,N_3851);
and U5216 (N_5216,N_2853,N_4960);
or U5217 (N_5217,N_1578,N_2078);
and U5218 (N_5218,N_2577,N_194);
xnor U5219 (N_5219,N_3166,N_1916);
and U5220 (N_5220,N_2621,N_1697);
xnor U5221 (N_5221,N_3692,N_4077);
nor U5222 (N_5222,N_573,N_2054);
nor U5223 (N_5223,N_4200,N_3913);
xor U5224 (N_5224,N_1935,N_404);
nor U5225 (N_5225,N_4990,N_2785);
or U5226 (N_5226,N_2437,N_3387);
nand U5227 (N_5227,N_3745,N_4187);
nand U5228 (N_5228,N_4950,N_602);
nor U5229 (N_5229,N_4201,N_4611);
and U5230 (N_5230,N_549,N_2933);
or U5231 (N_5231,N_2396,N_3793);
nor U5232 (N_5232,N_4977,N_1719);
or U5233 (N_5233,N_2689,N_4664);
and U5234 (N_5234,N_964,N_3699);
xor U5235 (N_5235,N_1211,N_2221);
nand U5236 (N_5236,N_3612,N_2027);
nand U5237 (N_5237,N_4157,N_1018);
nor U5238 (N_5238,N_764,N_2362);
nor U5239 (N_5239,N_1193,N_877);
and U5240 (N_5240,N_1506,N_4141);
xnor U5241 (N_5241,N_533,N_3299);
or U5242 (N_5242,N_1904,N_714);
or U5243 (N_5243,N_1735,N_4587);
nand U5244 (N_5244,N_544,N_4144);
nor U5245 (N_5245,N_4686,N_1027);
and U5246 (N_5246,N_3443,N_1401);
xor U5247 (N_5247,N_3553,N_2122);
nor U5248 (N_5248,N_2411,N_2687);
nand U5249 (N_5249,N_4427,N_1221);
or U5250 (N_5250,N_3829,N_906);
or U5251 (N_5251,N_3625,N_510);
nor U5252 (N_5252,N_1541,N_286);
and U5253 (N_5253,N_3941,N_4568);
or U5254 (N_5254,N_4932,N_2816);
nand U5255 (N_5255,N_3321,N_3405);
nor U5256 (N_5256,N_2923,N_2726);
nand U5257 (N_5257,N_606,N_4454);
nor U5258 (N_5258,N_3898,N_1479);
nor U5259 (N_5259,N_1951,N_2983);
or U5260 (N_5260,N_3766,N_1472);
nor U5261 (N_5261,N_1703,N_1941);
nand U5262 (N_5262,N_3635,N_3148);
and U5263 (N_5263,N_4441,N_4331);
or U5264 (N_5264,N_3736,N_4874);
nand U5265 (N_5265,N_1307,N_413);
or U5266 (N_5266,N_4895,N_232);
nand U5267 (N_5267,N_928,N_1674);
or U5268 (N_5268,N_1185,N_2200);
and U5269 (N_5269,N_116,N_1016);
or U5270 (N_5270,N_1261,N_4112);
xnor U5271 (N_5271,N_49,N_932);
nor U5272 (N_5272,N_2331,N_540);
xnor U5273 (N_5273,N_976,N_1045);
or U5274 (N_5274,N_3722,N_1041);
nor U5275 (N_5275,N_1670,N_4504);
nand U5276 (N_5276,N_2536,N_1641);
nor U5277 (N_5277,N_3072,N_4634);
xor U5278 (N_5278,N_29,N_4242);
nor U5279 (N_5279,N_2451,N_4000);
or U5280 (N_5280,N_1482,N_4637);
nand U5281 (N_5281,N_1249,N_584);
xnor U5282 (N_5282,N_3472,N_2272);
nor U5283 (N_5283,N_3191,N_4889);
xor U5284 (N_5284,N_735,N_4207);
or U5285 (N_5285,N_3821,N_4602);
or U5286 (N_5286,N_3994,N_4436);
xor U5287 (N_5287,N_3451,N_566);
nand U5288 (N_5288,N_1555,N_1223);
or U5289 (N_5289,N_465,N_2899);
xnor U5290 (N_5290,N_2059,N_882);
or U5291 (N_5291,N_4835,N_2350);
nor U5292 (N_5292,N_4667,N_4786);
nor U5293 (N_5293,N_632,N_4620);
and U5294 (N_5294,N_2289,N_4048);
and U5295 (N_5295,N_3720,N_3964);
and U5296 (N_5296,N_2332,N_3606);
xor U5297 (N_5297,N_126,N_400);
nor U5298 (N_5298,N_2658,N_2214);
xnor U5299 (N_5299,N_1933,N_4294);
or U5300 (N_5300,N_977,N_4596);
xnor U5301 (N_5301,N_3860,N_1442);
xnor U5302 (N_5302,N_1244,N_741);
nand U5303 (N_5303,N_3291,N_123);
and U5304 (N_5304,N_3946,N_3904);
nand U5305 (N_5305,N_2494,N_3093);
and U5306 (N_5306,N_4063,N_4995);
or U5307 (N_5307,N_2549,N_571);
or U5308 (N_5308,N_4516,N_2680);
nor U5309 (N_5309,N_2908,N_1325);
and U5310 (N_5310,N_2836,N_450);
nand U5311 (N_5311,N_1068,N_3927);
or U5312 (N_5312,N_3518,N_1278);
and U5313 (N_5313,N_379,N_3346);
xnor U5314 (N_5314,N_1397,N_1646);
nand U5315 (N_5315,N_220,N_2100);
nand U5316 (N_5316,N_910,N_4477);
xor U5317 (N_5317,N_4561,N_4378);
xor U5318 (N_5318,N_2305,N_4298);
nand U5319 (N_5319,N_3463,N_4235);
xnor U5320 (N_5320,N_542,N_14);
xor U5321 (N_5321,N_3277,N_921);
nor U5322 (N_5322,N_4751,N_3653);
xnor U5323 (N_5323,N_633,N_3234);
xnor U5324 (N_5324,N_4215,N_940);
and U5325 (N_5325,N_5,N_2316);
nand U5326 (N_5326,N_4719,N_3905);
and U5327 (N_5327,N_1942,N_1102);
nand U5328 (N_5328,N_1171,N_26);
xor U5329 (N_5329,N_1672,N_464);
xnor U5330 (N_5330,N_4087,N_570);
and U5331 (N_5331,N_1196,N_304);
nor U5332 (N_5332,N_2537,N_3359);
or U5333 (N_5333,N_1205,N_2037);
xor U5334 (N_5334,N_672,N_388);
and U5335 (N_5335,N_4961,N_3007);
or U5336 (N_5336,N_4081,N_2284);
and U5337 (N_5337,N_2903,N_2789);
nor U5338 (N_5338,N_2383,N_4846);
or U5339 (N_5339,N_4146,N_3380);
nor U5340 (N_5340,N_2950,N_179);
and U5341 (N_5341,N_2506,N_1477);
xor U5342 (N_5342,N_3169,N_2718);
or U5343 (N_5343,N_4383,N_1167);
nor U5344 (N_5344,N_4020,N_1313);
xor U5345 (N_5345,N_224,N_4548);
nand U5346 (N_5346,N_2241,N_656);
or U5347 (N_5347,N_95,N_908);
and U5348 (N_5348,N_4557,N_1187);
xor U5349 (N_5349,N_1130,N_3124);
xor U5350 (N_5350,N_1512,N_449);
or U5351 (N_5351,N_2732,N_38);
and U5352 (N_5352,N_712,N_4199);
and U5353 (N_5353,N_1484,N_2186);
nand U5354 (N_5354,N_4828,N_1323);
nor U5355 (N_5355,N_1297,N_733);
or U5356 (N_5356,N_1728,N_1216);
nand U5357 (N_5357,N_4797,N_499);
nor U5358 (N_5358,N_1329,N_3497);
or U5359 (N_5359,N_243,N_4560);
xor U5360 (N_5360,N_496,N_1805);
nand U5361 (N_5361,N_1994,N_4883);
or U5362 (N_5362,N_4204,N_1121);
nor U5363 (N_5363,N_4617,N_800);
xnor U5364 (N_5364,N_3878,N_104);
nor U5365 (N_5365,N_3508,N_1766);
and U5366 (N_5366,N_2364,N_1553);
nor U5367 (N_5367,N_1967,N_4149);
or U5368 (N_5368,N_2865,N_2008);
or U5369 (N_5369,N_358,N_3170);
nor U5370 (N_5370,N_2922,N_983);
nand U5371 (N_5371,N_4385,N_3952);
xor U5372 (N_5372,N_1687,N_1113);
xor U5373 (N_5373,N_235,N_3403);
or U5374 (N_5374,N_709,N_630);
nor U5375 (N_5375,N_2611,N_4982);
nand U5376 (N_5376,N_2070,N_53);
xnor U5377 (N_5377,N_3685,N_2467);
nand U5378 (N_5378,N_1471,N_4419);
nor U5379 (N_5379,N_138,N_161);
and U5380 (N_5380,N_4171,N_4382);
nand U5381 (N_5381,N_1414,N_4736);
nor U5382 (N_5382,N_1819,N_853);
or U5383 (N_5383,N_3440,N_2955);
nand U5384 (N_5384,N_688,N_4845);
and U5385 (N_5385,N_4822,N_2336);
and U5386 (N_5386,N_1617,N_4304);
nor U5387 (N_5387,N_4910,N_3414);
nand U5388 (N_5388,N_1095,N_1758);
nand U5389 (N_5389,N_2418,N_3156);
xor U5390 (N_5390,N_3406,N_1545);
or U5391 (N_5391,N_110,N_607);
nand U5392 (N_5392,N_1745,N_4377);
nor U5393 (N_5393,N_3791,N_4779);
nor U5394 (N_5394,N_4854,N_1508);
nor U5395 (N_5395,N_4863,N_2645);
and U5396 (N_5396,N_2823,N_4393);
and U5397 (N_5397,N_3172,N_4726);
nor U5398 (N_5398,N_4979,N_4807);
xor U5399 (N_5399,N_986,N_3818);
or U5400 (N_5400,N_3566,N_308);
or U5401 (N_5401,N_4296,N_2192);
and U5402 (N_5402,N_2498,N_4855);
xor U5403 (N_5403,N_4735,N_1702);
nor U5404 (N_5404,N_722,N_4934);
and U5405 (N_5405,N_1247,N_2999);
or U5406 (N_5406,N_608,N_2564);
xor U5407 (N_5407,N_2280,N_177);
xor U5408 (N_5408,N_180,N_1286);
nand U5409 (N_5409,N_3127,N_4254);
and U5410 (N_5410,N_2673,N_4694);
and U5411 (N_5411,N_789,N_2633);
or U5412 (N_5412,N_120,N_1843);
nor U5413 (N_5413,N_3437,N_1523);
xnor U5414 (N_5414,N_3605,N_4517);
xor U5415 (N_5415,N_2897,N_3435);
nand U5416 (N_5416,N_677,N_4320);
and U5417 (N_5417,N_3395,N_2652);
nor U5418 (N_5418,N_3002,N_364);
nand U5419 (N_5419,N_4335,N_3495);
nand U5420 (N_5420,N_4827,N_886);
nor U5421 (N_5421,N_4282,N_3385);
xnor U5422 (N_5422,N_2496,N_4033);
or U5423 (N_5423,N_1750,N_508);
nor U5424 (N_5424,N_3374,N_2407);
nand U5425 (N_5425,N_2215,N_1043);
xnor U5426 (N_5426,N_567,N_4881);
xor U5427 (N_5427,N_3028,N_3054);
and U5428 (N_5428,N_4330,N_852);
xor U5429 (N_5429,N_2770,N_4473);
xnor U5430 (N_5430,N_2625,N_363);
or U5431 (N_5431,N_1474,N_2076);
nor U5432 (N_5432,N_3492,N_3353);
nand U5433 (N_5433,N_2578,N_4306);
nor U5434 (N_5434,N_2528,N_1047);
nor U5435 (N_5435,N_4177,N_424);
nor U5436 (N_5436,N_1052,N_1312);
and U5437 (N_5437,N_257,N_2886);
xor U5438 (N_5438,N_4089,N_1006);
and U5439 (N_5439,N_4747,N_2401);
or U5440 (N_5440,N_827,N_2838);
xor U5441 (N_5441,N_7,N_1026);
or U5442 (N_5442,N_4915,N_3065);
xnor U5443 (N_5443,N_2047,N_1838);
xnor U5444 (N_5444,N_2262,N_3997);
and U5445 (N_5445,N_1567,N_4030);
nand U5446 (N_5446,N_2649,N_4921);
or U5447 (N_5447,N_4375,N_2101);
nor U5448 (N_5448,N_2552,N_283);
nand U5449 (N_5449,N_4061,N_3258);
xnor U5450 (N_5450,N_1815,N_1975);
or U5451 (N_5451,N_4692,N_3349);
or U5452 (N_5452,N_4170,N_383);
and U5453 (N_5453,N_4322,N_4948);
nand U5454 (N_5454,N_1174,N_2841);
xor U5455 (N_5455,N_4413,N_824);
nor U5456 (N_5456,N_3158,N_4798);
xnor U5457 (N_5457,N_4334,N_2585);
or U5458 (N_5458,N_3494,N_462);
and U5459 (N_5459,N_2884,N_3063);
or U5460 (N_5460,N_3876,N_4724);
or U5461 (N_5461,N_4789,N_609);
and U5462 (N_5462,N_3862,N_3647);
and U5463 (N_5463,N_1178,N_3423);
nor U5464 (N_5464,N_2084,N_2827);
nand U5465 (N_5465,N_4840,N_4222);
xor U5466 (N_5466,N_4831,N_4649);
nand U5467 (N_5467,N_4842,N_2250);
or U5468 (N_5468,N_2438,N_2421);
nor U5469 (N_5469,N_3903,N_2697);
or U5470 (N_5470,N_3122,N_3982);
nor U5471 (N_5471,N_83,N_3775);
xor U5472 (N_5472,N_4197,N_3858);
or U5473 (N_5473,N_2270,N_2470);
and U5474 (N_5474,N_2461,N_833);
and U5475 (N_5475,N_1820,N_1530);
xor U5476 (N_5476,N_377,N_2160);
and U5477 (N_5477,N_1554,N_61);
and U5478 (N_5478,N_1355,N_4261);
nor U5479 (N_5479,N_4507,N_763);
and U5480 (N_5480,N_3526,N_4646);
xor U5481 (N_5481,N_4396,N_3677);
xnor U5482 (N_5482,N_603,N_1966);
nor U5483 (N_5483,N_3144,N_2690);
nand U5484 (N_5484,N_845,N_3491);
xnor U5485 (N_5485,N_2677,N_3928);
nand U5486 (N_5486,N_4312,N_3970);
or U5487 (N_5487,N_563,N_1862);
or U5488 (N_5488,N_1182,N_1696);
and U5489 (N_5489,N_808,N_1763);
nand U5490 (N_5490,N_1876,N_4916);
nand U5491 (N_5491,N_1315,N_3565);
nor U5492 (N_5492,N_2052,N_1795);
or U5493 (N_5493,N_135,N_2602);
and U5494 (N_5494,N_1295,N_4364);
and U5495 (N_5495,N_3436,N_223);
nand U5496 (N_5496,N_3233,N_2131);
nor U5497 (N_5497,N_664,N_1230);
xnor U5498 (N_5498,N_3525,N_2228);
and U5499 (N_5499,N_918,N_1563);
or U5500 (N_5500,N_4425,N_4248);
and U5501 (N_5501,N_4043,N_4734);
and U5502 (N_5502,N_2788,N_3949);
nand U5503 (N_5503,N_4669,N_158);
and U5504 (N_5504,N_3863,N_4788);
nor U5505 (N_5505,N_3895,N_3922);
nor U5506 (N_5506,N_2685,N_472);
xor U5507 (N_5507,N_3129,N_1873);
xor U5508 (N_5508,N_835,N_2161);
nand U5509 (N_5509,N_991,N_142);
and U5510 (N_5510,N_736,N_4820);
xor U5511 (N_5511,N_1535,N_3792);
nor U5512 (N_5512,N_3594,N_3939);
and U5513 (N_5513,N_893,N_3598);
xnor U5514 (N_5514,N_3910,N_3820);
nor U5515 (N_5515,N_4398,N_2796);
and U5516 (N_5516,N_1761,N_1037);
or U5517 (N_5517,N_4344,N_1452);
xnor U5518 (N_5518,N_1606,N_434);
nor U5519 (N_5519,N_673,N_3587);
xor U5520 (N_5520,N_4013,N_545);
or U5521 (N_5521,N_1139,N_2700);
nor U5522 (N_5522,N_1888,N_268);
nand U5523 (N_5523,N_3382,N_2212);
xor U5524 (N_5524,N_3663,N_406);
or U5525 (N_5525,N_2405,N_4627);
nor U5526 (N_5526,N_2410,N_4037);
nand U5527 (N_5527,N_4525,N_1234);
nand U5528 (N_5528,N_4815,N_222);
nor U5529 (N_5529,N_2268,N_139);
nand U5530 (N_5530,N_2541,N_1499);
or U5531 (N_5531,N_3771,N_2239);
or U5532 (N_5532,N_3830,N_3059);
or U5533 (N_5533,N_2728,N_3115);
xor U5534 (N_5534,N_3824,N_1365);
nor U5535 (N_5535,N_1491,N_1800);
xnor U5536 (N_5536,N_834,N_4771);
and U5537 (N_5537,N_2957,N_2486);
nand U5538 (N_5538,N_3003,N_1009);
xnor U5539 (N_5539,N_4601,N_4464);
xor U5540 (N_5540,N_1028,N_997);
nand U5541 (N_5541,N_4238,N_1188);
or U5542 (N_5542,N_1731,N_4810);
or U5543 (N_5543,N_2701,N_690);
nor U5544 (N_5544,N_3468,N_1534);
and U5545 (N_5545,N_4702,N_1330);
nor U5546 (N_5546,N_1293,N_409);
nor U5547 (N_5547,N_4720,N_346);
and U5548 (N_5548,N_898,N_1605);
nor U5549 (N_5549,N_2156,N_4938);
nand U5550 (N_5550,N_4415,N_1893);
nor U5551 (N_5551,N_3199,N_1609);
or U5552 (N_5552,N_2207,N_648);
nand U5553 (N_5553,N_3428,N_1391);
xor U5554 (N_5554,N_11,N_1417);
or U5555 (N_5555,N_1746,N_1510);
xnor U5556 (N_5556,N_1021,N_3740);
and U5557 (N_5557,N_4984,N_4209);
xor U5558 (N_5558,N_546,N_1723);
xor U5559 (N_5559,N_2514,N_436);
or U5560 (N_5560,N_4270,N_739);
or U5561 (N_5561,N_227,N_1127);
nor U5562 (N_5562,N_270,N_697);
or U5563 (N_5563,N_757,N_183);
xor U5564 (N_5564,N_952,N_1870);
and U5565 (N_5565,N_1445,N_740);
or U5566 (N_5566,N_641,N_2213);
xnor U5567 (N_5567,N_3193,N_2871);
xnor U5568 (N_5568,N_1078,N_4317);
xor U5569 (N_5569,N_1179,N_3668);
or U5570 (N_5570,N_1648,N_4880);
xor U5571 (N_5571,N_4046,N_4812);
or U5572 (N_5572,N_4931,N_1281);
and U5573 (N_5573,N_3052,N_4808);
or U5574 (N_5574,N_1850,N_4185);
and U5575 (N_5575,N_225,N_2847);
xor U5576 (N_5576,N_2632,N_1053);
nor U5577 (N_5577,N_3424,N_3339);
or U5578 (N_5578,N_2218,N_3082);
and U5579 (N_5579,N_1082,N_2137);
or U5580 (N_5580,N_441,N_995);
xor U5581 (N_5581,N_1560,N_176);
and U5582 (N_5582,N_469,N_2414);
or U5583 (N_5583,N_3954,N_2256);
nand U5584 (N_5584,N_4687,N_2574);
or U5585 (N_5585,N_2820,N_148);
nor U5586 (N_5586,N_541,N_3106);
nor U5587 (N_5587,N_773,N_2110);
or U5588 (N_5588,N_4025,N_2551);
or U5589 (N_5589,N_2936,N_3355);
and U5590 (N_5590,N_4293,N_122);
xor U5591 (N_5591,N_3704,N_2900);
xnor U5592 (N_5592,N_4232,N_4656);
xnor U5593 (N_5593,N_2863,N_380);
or U5594 (N_5594,N_2729,N_3312);
nand U5595 (N_5595,N_4109,N_4408);
nand U5596 (N_5596,N_2453,N_3914);
nand U5597 (N_5597,N_708,N_4878);
nor U5598 (N_5598,N_35,N_0);
nand U5599 (N_5599,N_4326,N_317);
and U5600 (N_5600,N_1917,N_231);
nor U5601 (N_5601,N_598,N_3066);
nor U5602 (N_5602,N_2004,N_4183);
xor U5603 (N_5603,N_1833,N_1373);
and U5604 (N_5604,N_2126,N_3037);
nand U5605 (N_5605,N_1937,N_1135);
nor U5606 (N_5606,N_3017,N_3426);
xor U5607 (N_5607,N_915,N_4562);
and U5608 (N_5608,N_2091,N_2614);
and U5609 (N_5609,N_2310,N_4676);
nor U5610 (N_5610,N_3962,N_2859);
xnor U5611 (N_5611,N_786,N_40);
nor U5612 (N_5612,N_3978,N_2507);
nor U5613 (N_5613,N_509,N_2092);
xor U5614 (N_5614,N_1237,N_2889);
and U5615 (N_5615,N_1448,N_700);
or U5616 (N_5616,N_2304,N_2485);
nor U5617 (N_5617,N_4578,N_298);
nand U5618 (N_5618,N_4230,N_1025);
xor U5619 (N_5619,N_4541,N_3310);
nor U5620 (N_5620,N_3588,N_39);
and U5621 (N_5621,N_4906,N_1515);
or U5622 (N_5622,N_732,N_3642);
nand U5623 (N_5623,N_3673,N_2107);
and U5624 (N_5624,N_1575,N_1705);
xor U5625 (N_5625,N_1529,N_1324);
nand U5626 (N_5626,N_4543,N_1342);
nor U5627 (N_5627,N_2763,N_4384);
nor U5628 (N_5628,N_1611,N_814);
nor U5629 (N_5629,N_4368,N_1625);
and U5630 (N_5630,N_1304,N_475);
nand U5631 (N_5631,N_711,N_2518);
and U5632 (N_5632,N_4869,N_2376);
and U5633 (N_5633,N_1358,N_4939);
and U5634 (N_5634,N_378,N_1158);
and U5635 (N_5635,N_3599,N_2266);
xor U5636 (N_5636,N_3875,N_2622);
and U5637 (N_5637,N_4536,N_2267);
nor U5638 (N_5638,N_4865,N_2898);
xnor U5639 (N_5639,N_4742,N_3996);
xor U5640 (N_5640,N_4615,N_4675);
nand U5641 (N_5641,N_3885,N_3603);
nor U5642 (N_5642,N_3636,N_3500);
nor U5643 (N_5643,N_282,N_178);
and U5644 (N_5644,N_4604,N_2174);
and U5645 (N_5645,N_2879,N_1019);
nor U5646 (N_5646,N_1347,N_1110);
nor U5647 (N_5647,N_386,N_1120);
and U5648 (N_5648,N_2230,N_680);
nor U5649 (N_5649,N_473,N_3883);
nand U5650 (N_5650,N_4758,N_4862);
nand U5651 (N_5651,N_2402,N_106);
or U5652 (N_5652,N_4011,N_4336);
and U5653 (N_5653,N_3164,N_4856);
nor U5654 (N_5654,N_4651,N_3427);
nand U5655 (N_5655,N_1377,N_4754);
and U5656 (N_5656,N_3577,N_385);
xor U5657 (N_5657,N_3712,N_4376);
nor U5658 (N_5658,N_2741,N_4928);
nand U5659 (N_5659,N_210,N_1075);
or U5660 (N_5660,N_2727,N_3206);
or U5661 (N_5661,N_2590,N_4446);
xnor U5662 (N_5662,N_2686,N_3223);
nor U5663 (N_5663,N_2363,N_2663);
nand U5664 (N_5664,N_3089,N_4021);
nand U5665 (N_5665,N_3120,N_498);
and U5666 (N_5666,N_361,N_1400);
nor U5667 (N_5667,N_3078,N_1867);
and U5668 (N_5668,N_1715,N_1973);
and U5669 (N_5669,N_1177,N_2806);
nand U5670 (N_5670,N_3138,N_731);
xnor U5671 (N_5671,N_2223,N_4221);
xnor U5672 (N_5672,N_4139,N_4327);
nand U5673 (N_5673,N_191,N_4381);
or U5674 (N_5674,N_1918,N_24);
nand U5675 (N_5675,N_4164,N_4533);
or U5676 (N_5676,N_2172,N_1115);
or U5677 (N_5677,N_1503,N_644);
or U5678 (N_5678,N_3029,N_2031);
xnor U5679 (N_5679,N_1309,N_3690);
and U5680 (N_5680,N_2007,N_68);
or U5681 (N_5681,N_2761,N_55);
and U5682 (N_5682,N_4612,N_4229);
nor U5683 (N_5683,N_1734,N_3522);
and U5684 (N_5684,N_1724,N_1895);
nand U5685 (N_5685,N_4526,N_206);
and U5686 (N_5686,N_3631,N_16);
or U5687 (N_5687,N_439,N_2921);
and U5688 (N_5688,N_245,N_4947);
and U5689 (N_5689,N_2579,N_4060);
nand U5690 (N_5690,N_1054,N_4954);
xnor U5691 (N_5691,N_3036,N_1861);
xnor U5692 (N_5692,N_4803,N_569);
nor U5693 (N_5693,N_788,N_2720);
nor U5694 (N_5694,N_4964,N_3016);
nand U5695 (N_5695,N_3533,N_2066);
nand U5696 (N_5696,N_219,N_2055);
xor U5697 (N_5697,N_2260,N_2006);
or U5698 (N_5698,N_250,N_3765);
xor U5699 (N_5699,N_3343,N_4739);
nor U5700 (N_5700,N_1081,N_4274);
or U5701 (N_5701,N_147,N_1656);
or U5702 (N_5702,N_2340,N_2534);
xor U5703 (N_5703,N_1228,N_4339);
nand U5704 (N_5704,N_1266,N_3918);
or U5705 (N_5705,N_1481,N_3283);
nand U5706 (N_5706,N_1357,N_702);
nand U5707 (N_5707,N_2981,N_4360);
xnor U5708 (N_5708,N_4511,N_4674);
xnor U5709 (N_5709,N_3298,N_3703);
nor U5710 (N_5710,N_4328,N_2769);
nor U5711 (N_5711,N_216,N_1532);
nor U5712 (N_5712,N_604,N_1591);
and U5713 (N_5713,N_1760,N_3366);
or U5714 (N_5714,N_4622,N_4475);
and U5715 (N_5715,N_3788,N_4768);
nor U5716 (N_5716,N_4629,N_3950);
xor U5717 (N_5717,N_645,N_2302);
nor U5718 (N_5718,N_1055,N_81);
nor U5719 (N_5719,N_2154,N_230);
and U5720 (N_5720,N_1394,N_3912);
xor U5721 (N_5721,N_3743,N_3539);
nor U5722 (N_5722,N_207,N_278);
xor U5723 (N_5723,N_1804,N_2206);
nand U5724 (N_5724,N_1594,N_4826);
nand U5725 (N_5725,N_2802,N_3993);
and U5726 (N_5726,N_3955,N_4420);
nor U5727 (N_5727,N_4564,N_2293);
xor U5728 (N_5728,N_4787,N_1149);
and U5729 (N_5729,N_4945,N_23);
nor U5730 (N_5730,N_1792,N_3284);
xor U5731 (N_5731,N_927,N_3689);
or U5732 (N_5732,N_895,N_3611);
and U5733 (N_5733,N_2851,N_3691);
nor U5734 (N_5734,N_3308,N_12);
nor U5735 (N_5735,N_421,N_3789);
and U5736 (N_5736,N_369,N_1410);
xor U5737 (N_5737,N_4731,N_4028);
and U5738 (N_5738,N_2452,N_803);
or U5739 (N_5739,N_2106,N_1385);
xor U5740 (N_5740,N_796,N_2935);
nand U5741 (N_5741,N_638,N_3364);
or U5742 (N_5742,N_1954,N_149);
and U5743 (N_5743,N_870,N_2191);
and U5744 (N_5744,N_3006,N_1117);
nor U5745 (N_5745,N_1579,N_1964);
xor U5746 (N_5746,N_1610,N_628);
xnor U5747 (N_5747,N_1306,N_2033);
and U5748 (N_5748,N_1953,N_3850);
nand U5749 (N_5749,N_4753,N_4442);
or U5750 (N_5750,N_2666,N_1752);
nor U5751 (N_5751,N_729,N_2759);
nand U5752 (N_5752,N_3763,N_1574);
or U5753 (N_5753,N_2942,N_2837);
xnor U5754 (N_5754,N_1989,N_2301);
nand U5755 (N_5755,N_576,N_1318);
or U5756 (N_5756,N_3180,N_1832);
nand U5757 (N_5757,N_351,N_2219);
xnor U5758 (N_5758,N_4609,N_202);
nand U5759 (N_5759,N_3709,N_1806);
and U5760 (N_5760,N_4850,N_969);
nand U5761 (N_5761,N_1778,N_1602);
and U5762 (N_5762,N_4966,N_856);
nor U5763 (N_5763,N_461,N_1040);
nand U5764 (N_5764,N_10,N_4099);
and U5765 (N_5765,N_1721,N_1842);
and U5766 (N_5766,N_3019,N_3422);
and U5767 (N_5767,N_4591,N_1681);
xor U5768 (N_5768,N_2555,N_382);
or U5769 (N_5769,N_3460,N_4635);
nand U5770 (N_5770,N_1094,N_4342);
or U5771 (N_5771,N_3336,N_2620);
nor U5772 (N_5772,N_4859,N_1232);
and U5773 (N_5773,N_2255,N_4174);
nor U5774 (N_5774,N_1008,N_3051);
nor U5775 (N_5775,N_2312,N_3784);
and U5776 (N_5776,N_4528,N_2890);
nor U5777 (N_5777,N_2990,N_761);
nor U5778 (N_5778,N_1713,N_4521);
and U5779 (N_5779,N_2162,N_988);
nor U5780 (N_5780,N_4349,N_4265);
nand U5781 (N_5781,N_4655,N_2164);
and U5782 (N_5782,N_1346,N_4416);
nor U5783 (N_5783,N_1517,N_1316);
nand U5784 (N_5784,N_1759,N_2915);
or U5785 (N_5785,N_127,N_1181);
and U5786 (N_5786,N_3413,N_54);
and U5787 (N_5787,N_162,N_3173);
or U5788 (N_5788,N_4657,N_1464);
and U5789 (N_5789,N_2278,N_300);
xnor U5790 (N_5790,N_2930,N_3022);
xnor U5791 (N_5791,N_1339,N_3556);
and U5792 (N_5792,N_3356,N_2247);
nand U5793 (N_5793,N_4610,N_3142);
xor U5794 (N_5794,N_167,N_4431);
nand U5795 (N_5795,N_4486,N_917);
nand U5796 (N_5796,N_2896,N_3125);
or U5797 (N_5797,N_2446,N_420);
or U5798 (N_5798,N_1751,N_394);
or U5799 (N_5799,N_2867,N_3177);
nand U5800 (N_5800,N_4500,N_4860);
xor U5801 (N_5801,N_166,N_512);
nand U5802 (N_5802,N_51,N_96);
nor U5803 (N_5803,N_1900,N_2641);
xor U5804 (N_5804,N_2653,N_2603);
xor U5805 (N_5805,N_4031,N_1500);
nand U5806 (N_5806,N_4918,N_3959);
nand U5807 (N_5807,N_2320,N_1733);
or U5808 (N_5808,N_2702,N_2630);
xnor U5809 (N_5809,N_4417,N_4884);
nand U5810 (N_5810,N_1106,N_3749);
and U5811 (N_5811,N_864,N_2395);
or U5812 (N_5812,N_1255,N_1546);
and U5813 (N_5813,N_2022,N_1566);
and U5814 (N_5814,N_1175,N_89);
xnor U5815 (N_5815,N_169,N_4581);
nor U5816 (N_5816,N_2142,N_4218);
xor U5817 (N_5817,N_4600,N_4211);
or U5818 (N_5818,N_1321,N_2596);
xor U5819 (N_5819,N_2075,N_3698);
and U5820 (N_5820,N_1317,N_2869);
nor U5821 (N_5821,N_4315,N_4728);
or U5822 (N_5822,N_2557,N_417);
nand U5823 (N_5823,N_4074,N_170);
nand U5824 (N_5824,N_4523,N_1887);
nand U5825 (N_5825,N_4078,N_256);
and U5826 (N_5826,N_2264,N_3881);
nand U5827 (N_5827,N_3618,N_1049);
nand U5828 (N_5828,N_431,N_3293);
and U5829 (N_5829,N_4203,N_4633);
nor U5830 (N_5830,N_1497,N_2374);
xor U5831 (N_5831,N_1301,N_2443);
and U5832 (N_5832,N_776,N_2844);
and U5833 (N_5833,N_3114,N_2030);
xor U5834 (N_5834,N_1582,N_3386);
nand U5835 (N_5835,N_4316,N_3165);
or U5836 (N_5836,N_4115,N_3134);
and U5837 (N_5837,N_1402,N_890);
and U5838 (N_5838,N_3545,N_4848);
xor U5839 (N_5839,N_752,N_3055);
xnor U5840 (N_5840,N_820,N_2540);
or U5841 (N_5841,N_2891,N_189);
or U5842 (N_5842,N_1498,N_1944);
nand U5843 (N_5843,N_805,N_2561);
nor U5844 (N_5844,N_466,N_3803);
and U5845 (N_5845,N_3550,N_2098);
and U5846 (N_5846,N_659,N_2082);
xnor U5847 (N_5847,N_762,N_3536);
and U5848 (N_5848,N_4882,N_1389);
nand U5849 (N_5849,N_4257,N_1454);
nor U5850 (N_5850,N_2094,N_1461);
or U5851 (N_5851,N_849,N_1993);
xor U5852 (N_5852,N_1654,N_2032);
nand U5853 (N_5853,N_652,N_3474);
nand U5854 (N_5854,N_1565,N_3);
and U5855 (N_5855,N_289,N_979);
xor U5856 (N_5856,N_1198,N_2668);
nor U5857 (N_5857,N_1708,N_1056);
nand U5858 (N_5858,N_474,N_375);
nor U5859 (N_5859,N_1088,N_916);
xnor U5860 (N_5860,N_2097,N_42);
xor U5861 (N_5861,N_455,N_325);
xnor U5862 (N_5862,N_2225,N_4463);
xor U5863 (N_5863,N_2904,N_1505);
and U5864 (N_5864,N_3340,N_4027);
or U5865 (N_5865,N_4573,N_1785);
or U5866 (N_5866,N_76,N_1112);
nor U5867 (N_5867,N_1877,N_244);
xor U5868 (N_5868,N_4075,N_2023);
xor U5869 (N_5869,N_4216,N_1684);
or U5870 (N_5870,N_4550,N_3563);
xnor U5871 (N_5871,N_2440,N_2743);
nand U5872 (N_5872,N_4213,N_1540);
or U5873 (N_5873,N_2133,N_1243);
and U5874 (N_5874,N_3084,N_1914);
nor U5875 (N_5875,N_3044,N_3450);
or U5876 (N_5876,N_1104,N_1803);
or U5877 (N_5877,N_1507,N_1087);
nor U5878 (N_5878,N_840,N_2758);
and U5879 (N_5879,N_3924,N_2112);
nand U5880 (N_5880,N_1011,N_240);
or U5881 (N_5881,N_3257,N_3503);
xor U5882 (N_5882,N_1896,N_1097);
nor U5883 (N_5883,N_4278,N_1974);
xor U5884 (N_5884,N_4062,N_267);
xor U5885 (N_5885,N_2723,N_1716);
and U5886 (N_5886,N_1640,N_574);
xnor U5887 (N_5887,N_2403,N_4182);
and U5888 (N_5888,N_3639,N_1061);
and U5889 (N_5889,N_1816,N_3275);
or U5890 (N_5890,N_3879,N_3196);
or U5891 (N_5891,N_3936,N_3442);
nor U5892 (N_5892,N_3221,N_1133);
or U5893 (N_5893,N_2170,N_347);
and U5894 (N_5894,N_3519,N_2384);
or U5895 (N_5895,N_4625,N_993);
nor U5896 (N_5896,N_1644,N_1291);
nor U5897 (N_5897,N_3326,N_3209);
nor U5898 (N_5898,N_2670,N_3204);
nor U5899 (N_5899,N_3447,N_2361);
nand U5900 (N_5900,N_925,N_184);
xor U5901 (N_5901,N_454,N_4654);
nand U5902 (N_5902,N_2372,N_675);
xnor U5903 (N_5903,N_4794,N_4151);
and U5904 (N_5904,N_2143,N_3013);
xnor U5905 (N_5905,N_2538,N_1753);
nand U5906 (N_5906,N_305,N_2323);
xor U5907 (N_5907,N_3833,N_302);
and U5908 (N_5908,N_2817,N_3021);
or U5909 (N_5909,N_2074,N_2581);
or U5910 (N_5910,N_4233,N_1621);
nand U5911 (N_5911,N_3661,N_4530);
xor U5912 (N_5912,N_2085,N_3365);
nand U5913 (N_5913,N_2683,N_19);
xor U5914 (N_5914,N_3369,N_839);
or U5915 (N_5915,N_1841,N_1977);
xnor U5916 (N_5916,N_1164,N_4036);
or U5917 (N_5917,N_2750,N_3759);
and U5918 (N_5918,N_3415,N_3329);
xnor U5919 (N_5919,N_2997,N_838);
or U5920 (N_5920,N_4088,N_1851);
nand U5921 (N_5921,N_1992,N_1453);
and U5922 (N_5922,N_4538,N_3942);
and U5923 (N_5923,N_4994,N_3181);
nor U5924 (N_5924,N_407,N_4769);
xor U5925 (N_5925,N_74,N_4481);
or U5926 (N_5926,N_1284,N_2134);
nor U5927 (N_5927,N_4870,N_2885);
nor U5928 (N_5928,N_1990,N_4225);
and U5929 (N_5929,N_3517,N_3067);
and U5930 (N_5930,N_2533,N_887);
and U5931 (N_5931,N_1184,N_1380);
and U5932 (N_5932,N_4491,N_3734);
and U5933 (N_5933,N_654,N_4688);
nor U5934 (N_5934,N_3589,N_4300);
nand U5935 (N_5935,N_4004,N_78);
and U5936 (N_5936,N_4616,N_4572);
xnor U5937 (N_5937,N_2926,N_4965);
xor U5938 (N_5938,N_1496,N_1709);
or U5939 (N_5939,N_1148,N_517);
or U5940 (N_5940,N_3584,N_3056);
nand U5941 (N_5941,N_1710,N_2642);
or U5942 (N_5942,N_2694,N_2171);
nand U5943 (N_5943,N_3461,N_3554);
and U5944 (N_5944,N_1738,N_4404);
nor U5945 (N_5945,N_1265,N_1398);
xnor U5946 (N_5946,N_4076,N_482);
nand U5947 (N_5947,N_4016,N_3376);
nor U5948 (N_5948,N_738,N_1231);
xnor U5949 (N_5949,N_3132,N_425);
or U5950 (N_5950,N_457,N_4080);
or U5951 (N_5951,N_1959,N_4836);
nor U5952 (N_5952,N_3350,N_3813);
xnor U5953 (N_5953,N_15,N_3802);
and U5954 (N_5954,N_4876,N_1201);
nand U5955 (N_5955,N_616,N_1957);
nor U5956 (N_5956,N_2708,N_1593);
nand U5957 (N_5957,N_810,N_4885);
or U5958 (N_5958,N_301,N_1879);
nand U5959 (N_5959,N_4871,N_371);
or U5960 (N_5960,N_3068,N_1683);
or U5961 (N_5961,N_4422,N_587);
xnor U5962 (N_5962,N_2742,N_2040);
xor U5963 (N_5963,N_150,N_3770);
or U5964 (N_5964,N_543,N_4588);
or U5965 (N_5965,N_1922,N_3136);
nand U5966 (N_5966,N_912,N_1589);
xnor U5967 (N_5967,N_4923,N_2805);
or U5968 (N_5968,N_2522,N_2845);
nor U5969 (N_5969,N_3664,N_4073);
nor U5970 (N_5970,N_3371,N_4277);
or U5971 (N_5971,N_3727,N_2872);
xnor U5972 (N_5972,N_3231,N_3182);
and U5973 (N_5973,N_826,N_3609);
or U5974 (N_5974,N_448,N_4012);
xnor U5975 (N_5975,N_1456,N_2299);
and U5976 (N_5976,N_3807,N_1046);
or U5977 (N_5977,N_1180,N_2477);
nor U5978 (N_5978,N_4685,N_3062);
or U5979 (N_5979,N_4886,N_1412);
and U5980 (N_5980,N_1520,N_4539);
nor U5981 (N_5981,N_28,N_4269);
or U5982 (N_5982,N_165,N_4907);
and U5983 (N_5983,N_3634,N_3098);
or U5984 (N_5984,N_1359,N_2982);
nand U5985 (N_5985,N_3102,N_564);
or U5986 (N_5986,N_605,N_154);
and U5987 (N_5987,N_3564,N_1580);
and U5988 (N_5988,N_4323,N_3620);
or U5989 (N_5989,N_1287,N_4575);
nor U5990 (N_5990,N_4240,N_2960);
xor U5991 (N_5991,N_2953,N_3894);
or U5992 (N_5992,N_4049,N_3864);
or U5993 (N_5993,N_2011,N_523);
and U5994 (N_5994,N_199,N_2724);
or U5995 (N_5995,N_3837,N_744);
xnor U5996 (N_5996,N_2951,N_4647);
nand U5997 (N_5997,N_4212,N_1915);
nand U5998 (N_5998,N_3215,N_4105);
and U5999 (N_5999,N_1311,N_32);
nand U6000 (N_6000,N_2345,N_807);
nor U6001 (N_6001,N_3869,N_1767);
nand U6002 (N_6002,N_4468,N_4476);
nor U6003 (N_6003,N_3624,N_1882);
or U6004 (N_6004,N_1926,N_4640);
and U6005 (N_6005,N_1988,N_1361);
and U6006 (N_6006,N_312,N_4487);
and U6007 (N_6007,N_1253,N_4324);
nand U6008 (N_6008,N_2940,N_357);
xnor U6009 (N_6009,N_4399,N_4142);
nor U6010 (N_6010,N_1240,N_1675);
or U6011 (N_6011,N_3152,N_4098);
and U6012 (N_6012,N_754,N_2547);
and U6013 (N_6013,N_255,N_3842);
and U6014 (N_6014,N_2456,N_1036);
or U6015 (N_6015,N_4310,N_4433);
or U6016 (N_6016,N_18,N_676);
or U6017 (N_6017,N_4262,N_2400);
xor U6018 (N_6018,N_368,N_3706);
xor U6019 (N_6019,N_3189,N_483);
nor U6020 (N_6020,N_2593,N_1269);
nand U6021 (N_6021,N_3777,N_3613);
nand U6022 (N_6022,N_1747,N_1141);
xor U6023 (N_6023,N_3501,N_247);
nand U6024 (N_6024,N_3621,N_1855);
and U6025 (N_6025,N_3344,N_4217);
xnor U6026 (N_6026,N_463,N_4356);
and U6027 (N_6027,N_2371,N_4914);
nand U6028 (N_6028,N_2962,N_4518);
xnor U6029 (N_6029,N_1060,N_3153);
nand U6030 (N_6030,N_902,N_3466);
nor U6031 (N_6031,N_3535,N_3943);
nand U6032 (N_6032,N_2906,N_568);
or U6033 (N_6033,N_324,N_595);
and U6034 (N_6034,N_4639,N_1943);
or U6035 (N_6035,N_2979,N_580);
or U6036 (N_6036,N_859,N_3933);
xor U6037 (N_6037,N_577,N_1662);
nor U6038 (N_6038,N_4129,N_4843);
nor U6039 (N_6039,N_1790,N_1511);
or U6040 (N_6040,N_3039,N_3940);
xnor U6041 (N_6041,N_620,N_781);
or U6042 (N_6042,N_2546,N_1813);
or U6043 (N_6043,N_1488,N_3354);
nor U6044 (N_6044,N_4968,N_2989);
nand U6045 (N_6045,N_2291,N_3750);
xnor U6046 (N_6046,N_2946,N_4226);
xor U6047 (N_6047,N_1881,N_4861);
xnor U6048 (N_6048,N_2196,N_2888);
nand U6049 (N_6049,N_3578,N_4369);
and U6050 (N_6050,N_1421,N_2197);
and U6051 (N_6051,N_4227,N_486);
nor U6052 (N_6052,N_934,N_4577);
or U6053 (N_6053,N_1592,N_1132);
or U6054 (N_6054,N_2944,N_4717);
xor U6055 (N_6055,N_1676,N_1772);
xor U6056 (N_6056,N_440,N_506);
xnor U6057 (N_6057,N_4273,N_3640);
and U6058 (N_6058,N_1420,N_4508);
and U6059 (N_6059,N_4819,N_4104);
or U6060 (N_6060,N_1298,N_2113);
nand U6061 (N_6061,N_3324,N_524);
nand U6062 (N_6062,N_3103,N_913);
or U6063 (N_6063,N_2240,N_1587);
xnor U6064 (N_6064,N_1129,N_333);
or U6065 (N_6065,N_4447,N_897);
nand U6066 (N_6066,N_2468,N_3361);
and U6067 (N_6067,N_617,N_3600);
nor U6068 (N_6068,N_1277,N_4341);
nand U6069 (N_6069,N_3841,N_4959);
or U6070 (N_6070,N_4411,N_3248);
and U6071 (N_6071,N_2051,N_2773);
or U6072 (N_6072,N_1693,N_2792);
and U6073 (N_6073,N_4985,N_130);
nand U6074 (N_6074,N_4113,N_3010);
nor U6075 (N_6075,N_1072,N_2665);
nor U6076 (N_6076,N_307,N_978);
nand U6077 (N_6077,N_2125,N_2254);
and U6078 (N_6078,N_4890,N_3483);
or U6079 (N_6079,N_971,N_1035);
xnor U6080 (N_6080,N_4571,N_4246);
nand U6081 (N_6081,N_3855,N_2130);
nand U6082 (N_6082,N_1694,N_956);
and U6083 (N_6083,N_2502,N_3053);
and U6084 (N_6084,N_1351,N_56);
and U6085 (N_6085,N_1319,N_3645);
xnor U6086 (N_6086,N_791,N_3729);
nand U6087 (N_6087,N_4791,N_2612);
nand U6088 (N_6088,N_624,N_3034);
nor U6089 (N_6089,N_1076,N_4292);
and U6090 (N_6090,N_1390,N_901);
and U6091 (N_6091,N_3987,N_3195);
or U6092 (N_6092,N_4284,N_1699);
and U6093 (N_6093,N_4409,N_3726);
xor U6094 (N_6094,N_2591,N_4683);
and U6095 (N_6095,N_2086,N_728);
or U6096 (N_6096,N_3429,N_3278);
nand U6097 (N_6097,N_2881,N_4263);
and U6098 (N_6098,N_2830,N_2145);
or U6099 (N_6099,N_2674,N_71);
xor U6100 (N_6100,N_1559,N_2043);
or U6101 (N_6101,N_961,N_815);
nand U6102 (N_6102,N_500,N_4841);
nor U6103 (N_6103,N_4395,N_4547);
xor U6104 (N_6104,N_4772,N_100);
xor U6105 (N_6105,N_2500,N_3527);
xor U6106 (N_6106,N_1455,N_1714);
nor U6107 (N_6107,N_2993,N_2460);
or U6108 (N_6108,N_3967,N_1701);
xnor U6109 (N_6109,N_4490,N_4108);
nor U6110 (N_6110,N_1226,N_596);
and U6111 (N_6111,N_3741,N_200);
or U6112 (N_6112,N_4998,N_4662);
and U6113 (N_6113,N_2672,N_4554);
nor U6114 (N_6114,N_3101,N_720);
or U6115 (N_6115,N_1326,N_4132);
and U6116 (N_6116,N_2013,N_957);
xor U6117 (N_6117,N_2984,N_4018);
nor U6118 (N_6118,N_4703,N_4321);
and U6119 (N_6119,N_623,N_1502);
nor U6120 (N_6120,N_4297,N_3105);
nor U6121 (N_6121,N_1012,N_1736);
nand U6122 (N_6122,N_2617,N_4338);
and U6123 (N_6123,N_4206,N_1634);
nor U6124 (N_6124,N_2389,N_2121);
nor U6125 (N_6125,N_3087,N_1658);
xnor U6126 (N_6126,N_2607,N_303);
xor U6127 (N_6127,N_2,N_60);
nand U6128 (N_6128,N_2764,N_4952);
nor U6129 (N_6129,N_4755,N_548);
and U6130 (N_6130,N_1558,N_4872);
or U6131 (N_6131,N_4461,N_2159);
xnor U6132 (N_6132,N_2553,N_3345);
nand U6133 (N_6133,N_3814,N_3484);
xnor U6134 (N_6134,N_841,N_1123);
and U6135 (N_6135,N_3327,N_1469);
xnor U6136 (N_6136,N_4603,N_1542);
nor U6137 (N_6137,N_750,N_4469);
or U6138 (N_6138,N_989,N_3118);
nor U6139 (N_6139,N_4181,N_3623);
xor U6140 (N_6140,N_335,N_175);
and U6141 (N_6141,N_1430,N_1912);
xnor U6142 (N_6142,N_2740,N_4912);
nand U6143 (N_6143,N_3033,N_67);
nand U6144 (N_6144,N_2190,N_3097);
nor U6145 (N_6145,N_2710,N_1089);
and U6146 (N_6146,N_1531,N_4241);
nor U6147 (N_6147,N_4287,N_2615);
nand U6148 (N_6148,N_2671,N_3688);
or U6149 (N_6149,N_3617,N_3485);
nor U6150 (N_6150,N_1781,N_2378);
and U6151 (N_6151,N_112,N_1688);
nor U6152 (N_6152,N_942,N_4325);
nand U6153 (N_6153,N_1783,N_4471);
xnor U6154 (N_6154,N_1970,N_2864);
nand U6155 (N_6155,N_924,N_1930);
and U6156 (N_6156,N_114,N_3744);
and U6157 (N_6157,N_271,N_1899);
nand U6158 (N_6158,N_1866,N_4250);
or U6159 (N_6159,N_3932,N_848);
nor U6160 (N_6160,N_4773,N_1603);
nor U6161 (N_6161,N_4857,N_1613);
xnor U6162 (N_6162,N_2140,N_2425);
and U6163 (N_6163,N_3254,N_4093);
nor U6164 (N_6164,N_3225,N_4069);
xnor U6165 (N_6165,N_132,N_1690);
nand U6166 (N_6166,N_4055,N_2354);
nand U6167 (N_6167,N_790,N_1396);
and U6168 (N_6168,N_3757,N_4145);
xnor U6169 (N_6169,N_2662,N_1161);
nor U6170 (N_6170,N_1077,N_4598);
nand U6171 (N_6171,N_2977,N_1818);
nand U6172 (N_6172,N_1650,N_2141);
nor U6173 (N_6173,N_2048,N_4540);
and U6174 (N_6174,N_3551,N_2246);
or U6175 (N_6175,N_246,N_2188);
xor U6176 (N_6176,N_2834,N_3746);
xnor U6177 (N_6177,N_1848,N_1073);
nor U6178 (N_6178,N_1388,N_4830);
or U6179 (N_6179,N_3081,N_2120);
nor U6180 (N_6180,N_4534,N_4823);
or U6181 (N_6181,N_1849,N_3686);
nand U6182 (N_6182,N_2050,N_3515);
nand U6183 (N_6183,N_666,N_3368);
nand U6184 (N_6184,N_621,N_817);
and U6185 (N_6185,N_1777,N_1521);
nor U6186 (N_6186,N_1577,N_2483);
nor U6187 (N_6187,N_3333,N_2568);
xor U6188 (N_6188,N_2531,N_4056);
and U6189 (N_6189,N_349,N_1775);
xor U6190 (N_6190,N_2346,N_4097);
and U6191 (N_6191,N_1614,N_1630);
nand U6192 (N_6192,N_3938,N_3159);
nand U6193 (N_6193,N_1418,N_2765);
or U6194 (N_6194,N_2439,N_3925);
nand U6195 (N_6195,N_1769,N_3362);
nor U6196 (N_6196,N_4520,N_4574);
nand U6197 (N_6197,N_1597,N_3670);
nand U6198 (N_6198,N_1257,N_4352);
nor U6199 (N_6199,N_4192,N_4766);
xnor U6200 (N_6200,N_2866,N_3218);
and U6201 (N_6201,N_1241,N_1415);
nand U6202 (N_6202,N_2822,N_2068);
nand U6203 (N_6203,N_503,N_4567);
and U6204 (N_6204,N_266,N_1042);
xnor U6205 (N_6205,N_2153,N_395);
nor U6206 (N_6206,N_3887,N_3701);
nand U6207 (N_6207,N_1787,N_4258);
and U6208 (N_6208,N_2628,N_3868);
xor U6209 (N_6209,N_4936,N_1322);
nand U6210 (N_6210,N_1945,N_2807);
or U6211 (N_6211,N_22,N_2459);
xor U6212 (N_6212,N_1005,N_2285);
nand U6213 (N_6213,N_3030,N_1438);
nand U6214 (N_6214,N_489,N_2046);
nand U6215 (N_6215,N_4917,N_737);
or U6216 (N_6216,N_2184,N_4981);
xnor U6217 (N_6217,N_3282,N_1972);
xnor U6218 (N_6218,N_2321,N_4608);
and U6219 (N_6219,N_261,N_4645);
nor U6220 (N_6220,N_140,N_3649);
nor U6221 (N_6221,N_557,N_3141);
nor U6222 (N_6222,N_756,N_4276);
or U6223 (N_6223,N_1408,N_2501);
and U6224 (N_6224,N_1636,N_1927);
and U6225 (N_6225,N_1419,N_2187);
or U6226 (N_6226,N_25,N_3758);
nor U6227 (N_6227,N_960,N_3804);
xnor U6228 (N_6228,N_1010,N_4879);
nand U6229 (N_6229,N_4150,N_4927);
and U6230 (N_6230,N_2146,N_2503);
xor U6231 (N_6231,N_1015,N_2116);
nand U6232 (N_6232,N_1871,N_3538);
xnor U6233 (N_6233,N_2385,N_1770);
and U6234 (N_6234,N_922,N_2588);
or U6235 (N_6235,N_562,N_254);
nand U6236 (N_6236,N_3751,N_285);
nand U6237 (N_6237,N_515,N_4972);
xnor U6238 (N_6238,N_1711,N_4245);
nor U6239 (N_6239,N_2787,N_2901);
nor U6240 (N_6240,N_1823,N_2678);
nor U6241 (N_6241,N_872,N_1289);
and U6242 (N_6242,N_205,N_2474);
xnor U6243 (N_6243,N_4839,N_4291);
nand U6244 (N_6244,N_1938,N_3979);
or U6245 (N_6245,N_3871,N_2911);
or U6246 (N_6246,N_3502,N_3730);
or U6247 (N_6247,N_366,N_4390);
or U6248 (N_6248,N_2203,N_121);
nand U6249 (N_6249,N_4458,N_2209);
nand U6250 (N_6250,N_1936,N_3462);
or U6251 (N_6251,N_101,N_1519);
nor U6252 (N_6252,N_3108,N_3608);
xor U6253 (N_6253,N_414,N_2529);
nor U6254 (N_6254,N_360,N_1495);
and U6255 (N_6255,N_3004,N_3245);
or U6256 (N_6256,N_4400,N_4582);
or U6257 (N_6257,N_3795,N_4437);
nand U6258 (N_6258,N_1030,N_3041);
nor U6259 (N_6259,N_1509,N_2127);
nand U6260 (N_6260,N_4228,N_2099);
nor U6261 (N_6261,N_981,N_4946);
xor U6262 (N_6262,N_4551,N_3185);
or U6263 (N_6263,N_858,N_2712);
nor U6264 (N_6264,N_276,N_1432);
nand U6265 (N_6265,N_929,N_1490);
or U6266 (N_6266,N_487,N_3467);
xor U6267 (N_6267,N_3482,N_3575);
nor U6268 (N_6268,N_4642,N_3135);
xor U6269 (N_6269,N_322,N_2676);
nor U6270 (N_6270,N_263,N_723);
xnor U6271 (N_6271,N_4897,N_4631);
xor U6272 (N_6272,N_828,N_2489);
nor U6273 (N_6273,N_2815,N_1620);
xor U6274 (N_6274,N_1048,N_2426);
and U6275 (N_6275,N_4318,N_4499);
and U6276 (N_6276,N_3514,N_2335);
nand U6277 (N_6277,N_725,N_2311);
or U6278 (N_6278,N_1923,N_813);
and U6279 (N_6279,N_1274,N_4353);
or U6280 (N_6280,N_124,N_2123);
and U6281 (N_6281,N_1387,N_2609);
or U6282 (N_6282,N_3705,N_2812);
xor U6283 (N_6283,N_3687,N_2826);
or U6284 (N_6284,N_117,N_1704);
nor U6285 (N_6285,N_1601,N_4333);
or U6286 (N_6286,N_3397,N_519);
xor U6287 (N_6287,N_837,N_3504);
nand U6288 (N_6288,N_3838,N_354);
xor U6289 (N_6289,N_4244,N_2902);
and U6290 (N_6290,N_2369,N_3292);
nor U6291 (N_6291,N_2455,N_1405);
or U6292 (N_6292,N_1080,N_1340);
nand U6293 (N_6293,N_1649,N_291);
and U6294 (N_6294,N_1668,N_2512);
nor U6295 (N_6295,N_3214,N_3268);
nor U6296 (N_6296,N_2416,N_3899);
or U6297 (N_6297,N_2563,N_1362);
and U6298 (N_6298,N_1940,N_3079);
xor U6299 (N_6299,N_9,N_4295);
xnor U6300 (N_6300,N_3543,N_3459);
or U6301 (N_6301,N_1891,N_2584);
nand U6302 (N_6302,N_3207,N_3552);
and U6303 (N_6303,N_1628,N_905);
nand U6304 (N_6304,N_1070,N_4818);
xor U6305 (N_6305,N_547,N_3672);
or U6306 (N_6306,N_3937,N_1834);
xnor U6307 (N_6307,N_529,N_883);
nor U6308 (N_6308,N_3643,N_4790);
nand U6309 (N_6309,N_2018,N_1590);
and U6310 (N_6310,N_626,N_4503);
or U6311 (N_6311,N_3176,N_2640);
nor U6312 (N_6312,N_3075,N_4943);
nor U6313 (N_6313,N_966,N_2938);
nor U6314 (N_6314,N_1997,N_4971);
nor U6315 (N_6315,N_2650,N_3806);
and U6316 (N_6316,N_612,N_2479);
xor U6317 (N_6317,N_4793,N_1673);
nor U6318 (N_6318,N_1707,N_4064);
and U6319 (N_6319,N_3822,N_3658);
nor U6320 (N_6320,N_3493,N_416);
nor U6321 (N_6321,N_2343,N_3085);
nor U6322 (N_6322,N_1367,N_1706);
xnor U6323 (N_6323,N_3562,N_2417);
and U6324 (N_6324,N_3558,N_4357);
and U6325 (N_6325,N_3682,N_2359);
xnor U6326 (N_6326,N_3547,N_3614);
or U6327 (N_6327,N_581,N_4806);
nand U6328 (N_6328,N_197,N_62);
and U6329 (N_6329,N_1639,N_2654);
xnor U6330 (N_6330,N_2176,N_3920);
nand U6331 (N_6331,N_4774,N_4762);
and U6332 (N_6332,N_3464,N_3711);
and U6333 (N_6333,N_4264,N_1303);
nor U6334 (N_6334,N_1562,N_1128);
or U6335 (N_6335,N_3130,N_2567);
xnor U6336 (N_6336,N_4280,N_865);
and U6337 (N_6337,N_3025,N_1911);
or U6338 (N_6338,N_4372,N_1020);
nand U6339 (N_6339,N_2604,N_4993);
or U6340 (N_6340,N_4289,N_2275);
nor U6341 (N_6341,N_3095,N_3761);
xnor U6342 (N_6342,N_1971,N_1262);
xnor U6343 (N_6343,N_228,N_793);
nand U6344 (N_6344,N_3290,N_2786);
nand U6345 (N_6345,N_1968,N_2638);
nor U6346 (N_6346,N_514,N_2029);
nand U6347 (N_6347,N_2992,N_2492);
nor U6348 (N_6348,N_2713,N_1371);
xor U6349 (N_6349,N_2644,N_1831);
and U6350 (N_6350,N_2010,N_2314);
or U6351 (N_6351,N_4418,N_1150);
xor U6352 (N_6352,N_935,N_2095);
xor U6353 (N_6353,N_411,N_4307);
or U6354 (N_6354,N_2980,N_804);
or U6355 (N_6355,N_1963,N_1145);
or U6356 (N_6356,N_755,N_3301);
and U6357 (N_6357,N_2704,N_1413);
nand U6358 (N_6358,N_484,N_3874);
or U6359 (N_6359,N_2352,N_4799);
nand U6360 (N_6360,N_1627,N_962);
or U6361 (N_6361,N_2943,N_4777);
nor U6362 (N_6362,N_2860,N_4337);
nand U6363 (N_6363,N_311,N_4379);
nand U6364 (N_6364,N_842,N_442);
nand U6365 (N_6365,N_3560,N_1680);
nor U6366 (N_6366,N_3882,N_3825);
and U6367 (N_6367,N_4677,N_3190);
or U6368 (N_6368,N_2458,N_4630);
or U6369 (N_6369,N_4722,N_779);
nand U6370 (N_6370,N_2978,N_4748);
or U6371 (N_6371,N_2755,N_293);
nand U6372 (N_6372,N_1717,N_2177);
or U6373 (N_6373,N_2829,N_4193);
nand U6374 (N_6374,N_2344,N_1858);
or U6375 (N_6375,N_3227,N_717);
or U6376 (N_6376,N_1267,N_458);
nand U6377 (N_6377,N_3404,N_4925);
nor U6378 (N_6378,N_1771,N_2329);
xor U6379 (N_6379,N_4082,N_2932);
nor U6380 (N_6380,N_1985,N_3953);
and U6381 (N_6381,N_4484,N_90);
xor U6382 (N_6382,N_2071,N_1369);
or U6383 (N_6383,N_3799,N_2169);
nand U6384 (N_6384,N_2441,N_1908);
nand U6385 (N_6385,N_1547,N_4594);
xnor U6386 (N_6386,N_552,N_4015);
nor U6387 (N_6387,N_2135,N_1264);
nor U6388 (N_6388,N_2913,N_992);
nand U6389 (N_6389,N_4737,N_260);
nand U6390 (N_6390,N_4905,N_668);
and U6391 (N_6391,N_2877,N_1764);
nor U6392 (N_6392,N_2391,N_3147);
and U6393 (N_6393,N_1561,N_2996);
nand U6394 (N_6394,N_2038,N_2811);
or U6395 (N_6395,N_1754,N_4371);
nor U6396 (N_6396,N_3145,N_3985);
xor U6397 (N_6397,N_880,N_4045);
or U6398 (N_6398,N_3975,N_4663);
nand U6399 (N_6399,N_3303,N_2914);
nand U6400 (N_6400,N_4899,N_3438);
nand U6401 (N_6401,N_4767,N_1607);
or U6402 (N_6402,N_3200,N_1153);
or U6403 (N_6403,N_1642,N_3372);
xor U6404 (N_6404,N_4563,N_192);
xnor U6405 (N_6405,N_698,N_861);
xor U6406 (N_6406,N_4770,N_710);
and U6407 (N_6407,N_427,N_513);
or U6408 (N_6408,N_4370,N_2382);
nand U6409 (N_6409,N_2292,N_2988);
and U6410 (N_6410,N_614,N_972);
or U6411 (N_6411,N_3845,N_4169);
xnor U6412 (N_6412,N_2053,N_3747);
and U6413 (N_6413,N_4579,N_4457);
xor U6414 (N_6414,N_2655,N_3971);
or U6415 (N_6415,N_3796,N_4359);
and U6416 (N_6416,N_1376,N_4976);
and U6417 (N_6417,N_2800,N_3753);
nor U6418 (N_6418,N_1780,N_4279);
and U6419 (N_6419,N_4019,N_342);
nor U6420 (N_6420,N_4832,N_3123);
nand U6421 (N_6421,N_3241,N_2910);
nand U6422 (N_6422,N_4054,N_3923);
and U6423 (N_6423,N_4851,N_2360);
xnor U6424 (N_6424,N_4552,N_1215);
xor U6425 (N_6425,N_141,N_2959);
nand U6426 (N_6426,N_2349,N_2151);
or U6427 (N_6427,N_1160,N_4351);
and U6428 (N_6428,N_468,N_4482);
nor U6429 (N_6429,N_537,N_4194);
nor U6430 (N_6430,N_3419,N_3453);
nor U6431 (N_6431,N_4980,N_857);
nor U6432 (N_6432,N_3266,N_2855);
or U6433 (N_6433,N_3317,N_4309);
nand U6434 (N_6434,N_3247,N_1183);
nand U6435 (N_6435,N_3812,N_3073);
xnor U6436 (N_6436,N_3801,N_4853);
nor U6437 (N_6437,N_4763,N_3595);
or U6438 (N_6438,N_3381,N_3377);
nand U6439 (N_6439,N_1492,N_4583);
xnor U6440 (N_6440,N_3237,N_4944);
xor U6441 (N_6441,N_2224,N_181);
nor U6442 (N_6442,N_869,N_3934);
nand U6443 (N_6443,N_1155,N_4584);
xor U6444 (N_6444,N_1156,N_3012);
nor U6445 (N_6445,N_4401,N_3456);
xor U6446 (N_6446,N_1437,N_4721);
nor U6447 (N_6447,N_4699,N_2719);
or U6448 (N_6448,N_3601,N_2012);
nand U6449 (N_6449,N_4430,N_2282);
and U6450 (N_6450,N_2434,N_221);
and U6451 (N_6451,N_3133,N_3186);
nand U6452 (N_6452,N_3637,N_1906);
or U6453 (N_6453,N_3990,N_2813);
or U6454 (N_6454,N_3040,N_4071);
nand U6455 (N_6455,N_4986,N_2791);
nand U6456 (N_6456,N_2716,N_3035);
xnor U6457 (N_6457,N_2969,N_2429);
nand U6458 (N_6458,N_1395,N_365);
nor U6459 (N_6459,N_2103,N_4003);
or U6460 (N_6460,N_660,N_4196);
xnor U6461 (N_6461,N_3585,N_2034);
xor U6462 (N_6462,N_3198,N_3769);
or U6463 (N_6463,N_2448,N_446);
nand U6464 (N_6464,N_4920,N_4067);
or U6465 (N_6465,N_2472,N_3272);
xor U6466 (N_6466,N_1864,N_1202);
xor U6467 (N_6467,N_3316,N_381);
xnor U6468 (N_6468,N_2469,N_3911);
nand U6469 (N_6469,N_4101,N_1762);
nor U6470 (N_6470,N_1784,N_4120);
and U6471 (N_6471,N_4470,N_3654);
nor U6472 (N_6472,N_4983,N_3294);
and U6473 (N_6473,N_2639,N_526);
and U6474 (N_6474,N_3490,N_2017);
xnor U6475 (N_6475,N_4970,N_695);
nor U6476 (N_6476,N_3679,N_2136);
or U6477 (N_6477,N_1103,N_3626);
nand U6478 (N_6478,N_3880,N_4707);
or U6479 (N_6479,N_2158,N_4852);
or U6480 (N_6480,N_2398,N_525);
nand U6481 (N_6481,N_874,N_2208);
and U6482 (N_6482,N_4605,N_3242);
nor U6483 (N_6483,N_494,N_2318);
or U6484 (N_6484,N_4888,N_777);
and U6485 (N_6485,N_2623,N_1242);
nor U6486 (N_6486,N_108,N_782);
nor U6487 (N_6487,N_4973,N_3188);
nor U6488 (N_6488,N_4128,N_3202);
or U6489 (N_6489,N_1727,N_1466);
or U6490 (N_6490,N_4537,N_3131);
nor U6491 (N_6491,N_4044,N_3091);
or U6492 (N_6492,N_1435,N_1422);
nor U6493 (N_6493,N_480,N_1638);
nand U6494 (N_6494,N_1379,N_3828);
and U6495 (N_6495,N_994,N_1320);
or U6496 (N_6496,N_536,N_2342);
nor U6497 (N_6497,N_168,N_3998);
nor U6498 (N_6498,N_2044,N_2582);
and U6499 (N_6499,N_531,N_2804);
or U6500 (N_6500,N_2111,N_171);
nand U6501 (N_6501,N_253,N_707);
and U6502 (N_6502,N_2109,N_1208);
nor U6503 (N_6503,N_4825,N_878);
and U6504 (N_6504,N_2028,N_784);
xnor U6505 (N_6505,N_479,N_3718);
nand U6506 (N_6506,N_2784,N_2334);
or U6507 (N_6507,N_3798,N_1791);
or U6508 (N_6508,N_471,N_4272);
xor U6509 (N_6509,N_3270,N_4350);
or U6510 (N_6510,N_3390,N_4975);
nor U6511 (N_6511,N_4858,N_3347);
and U6512 (N_6512,N_2132,N_2586);
nand U6513 (N_6513,N_1288,N_1283);
nand U6514 (N_6514,N_2801,N_1485);
xor U6515 (N_6515,N_588,N_3756);
and U6516 (N_6516,N_387,N_911);
nand U6517 (N_6517,N_642,N_1032);
or U6518 (N_6518,N_4148,N_1154);
or U6519 (N_6519,N_4176,N_3507);
nor U6520 (N_6520,N_4387,N_4290);
xor U6521 (N_6521,N_1279,N_2745);
and U6522 (N_6522,N_3416,N_691);
nand U6523 (N_6523,N_453,N_3154);
nor U6524 (N_6524,N_625,N_551);
and U6525 (N_6525,N_6,N_694);
xnor U6526 (N_6526,N_3867,N_2298);
and U6527 (N_6527,N_2016,N_4231);
or U6528 (N_6528,N_3816,N_451);
and U6529 (N_6529,N_2705,N_3057);
nor U6530 (N_6530,N_2279,N_1450);
and U6531 (N_6531,N_3632,N_1929);
xor U6532 (N_6532,N_43,N_1909);
and U6533 (N_6533,N_2062,N_4709);
nand U6534 (N_6534,N_4569,N_1958);
xor U6535 (N_6535,N_3956,N_3418);
and U6536 (N_6536,N_3273,N_904);
or U6537 (N_6537,N_4665,N_157);
xor U6538 (N_6538,N_903,N_4224);
nand U6539 (N_6539,N_3457,N_1700);
nand U6540 (N_6540,N_1429,N_1136);
xnor U6541 (N_6541,N_1859,N_1483);
nand U6542 (N_6542,N_2808,N_4053);
and U6543 (N_6543,N_3398,N_4991);
nor U6544 (N_6544,N_4632,N_1570);
and U6545 (N_6545,N_582,N_555);
xor U6546 (N_6546,N_535,N_3721);
nor U6547 (N_6547,N_3479,N_1004);
nor U6548 (N_6548,N_1679,N_3175);
and U6549 (N_6549,N_2165,N_452);
and U6550 (N_6550,N_1524,N_3410);
nand U6551 (N_6551,N_1444,N_2061);
nand U6552 (N_6552,N_2965,N_2843);
and U6553 (N_6553,N_3583,N_4440);
and U6554 (N_6554,N_2775,N_1272);
and U6555 (N_6555,N_1504,N_4066);
xor U6556 (N_6556,N_4354,N_2991);
nor U6557 (N_6557,N_355,N_953);
nand U6558 (N_6558,N_1363,N_2571);
and U6559 (N_6559,N_3246,N_3921);
xor U6560 (N_6560,N_1360,N_2265);
nand U6561 (N_6561,N_646,N_2248);
nand U6562 (N_6562,N_1573,N_819);
nand U6563 (N_6563,N_3866,N_4223);
xnor U6564 (N_6564,N_4285,N_1932);
or U6565 (N_6565,N_460,N_4435);
nand U6566 (N_6566,N_193,N_640);
and U6567 (N_6567,N_3724,N_4140);
and U6568 (N_6568,N_2516,N_2419);
nor U6569 (N_6569,N_4188,N_1802);
or U6570 (N_6570,N_1720,N_2019);
and U6571 (N_6571,N_3945,N_3070);
nor U6572 (N_6572,N_4219,N_4515);
nand U6573 (N_6573,N_343,N_1840);
and U6574 (N_6574,N_3496,N_3137);
nand U6575 (N_6575,N_3058,N_3648);
and U6576 (N_6576,N_2303,N_1537);
or U6577 (N_6577,N_3217,N_2527);
xnor U6578 (N_6578,N_748,N_1064);
or U6579 (N_6579,N_2832,N_943);
xor U6580 (N_6580,N_1756,N_611);
and U6581 (N_6581,N_3287,N_4002);
nand U6582 (N_6582,N_4355,N_2892);
or U6583 (N_6583,N_1743,N_2482);
nor U6584 (N_6584,N_2963,N_478);
xnor U6585 (N_6585,N_1463,N_860);
nor U6586 (N_6586,N_1259,N_3229);
or U6587 (N_6587,N_3071,N_146);
nand U6588 (N_6588,N_2194,N_1029);
nand U6589 (N_6589,N_4746,N_1556);
or U6590 (N_6590,N_2919,N_4513);
nor U6591 (N_6591,N_2181,N_593);
and U6592 (N_6592,N_2976,N_4478);
nor U6593 (N_6593,N_4243,N_745);
xnor U6594 (N_6594,N_4136,N_4116);
nand U6595 (N_6595,N_188,N_758);
or U6596 (N_6596,N_4714,N_36);
xnor U6597 (N_6597,N_485,N_759);
and U6598 (N_6598,N_2878,N_3274);
and U6599 (N_6599,N_3592,N_3676);
nand U6600 (N_6600,N_3384,N_2873);
xor U6601 (N_6601,N_1886,N_2646);
xnor U6602 (N_6602,N_401,N_275);
nand U6603 (N_6603,N_1755,N_4260);
nor U6604 (N_6604,N_2907,N_1730);
nand U6605 (N_6605,N_2317,N_3984);
xor U6606 (N_6606,N_470,N_4065);
nor U6607 (N_6607,N_2744,N_2918);
nor U6608 (N_6608,N_4903,N_4868);
or U6609 (N_6609,N_1467,N_2858);
nand U6610 (N_6610,N_3338,N_3958);
xnor U6611 (N_6611,N_209,N_1138);
and U6612 (N_6612,N_1236,N_4556);
or U6613 (N_6613,N_3208,N_706);
xor U6614 (N_6614,N_1260,N_2952);
nor U6615 (N_6615,N_4743,N_3219);
or U6616 (N_6616,N_3980,N_1661);
nor U6617 (N_6617,N_152,N_2150);
nand U6618 (N_6618,N_701,N_3827);
xnor U6619 (N_6619,N_1878,N_1824);
or U6620 (N_6620,N_950,N_47);
nor U6621 (N_6621,N_3325,N_57);
or U6622 (N_6622,N_1473,N_2324);
nand U6623 (N_6623,N_816,N_4034);
or U6624 (N_6624,N_3253,N_85);
nor U6625 (N_6625,N_4765,N_4022);
xnor U6626 (N_6626,N_4589,N_3719);
and U6627 (N_6627,N_4834,N_3445);
and U6628 (N_6628,N_3315,N_4723);
nor U6629 (N_6629,N_3764,N_4811);
nand U6630 (N_6630,N_2373,N_2420);
nor U6631 (N_6631,N_4172,N_2227);
xnor U6632 (N_6632,N_306,N_3908);
or U6633 (N_6633,N_742,N_3884);
xor U6634 (N_6634,N_3968,N_1338);
xnor U6635 (N_6635,N_2511,N_143);
nand U6636 (N_6636,N_3259,N_2287);
nor U6637 (N_6637,N_4780,N_429);
and U6638 (N_6638,N_4875,N_3800);
and U6639 (N_6639,N_4198,N_1898);
or U6640 (N_6640,N_2357,N_4208);
nor U6641 (N_6641,N_1111,N_4716);
and U6642 (N_6642,N_33,N_3707);
and U6643 (N_6643,N_3475,N_1655);
or U6644 (N_6644,N_532,N_3295);
nand U6645 (N_6645,N_1057,N_1698);
or U6646 (N_6646,N_946,N_1476);
nand U6647 (N_6647,N_4585,N_4057);
nand U6648 (N_6648,N_561,N_2404);
and U6649 (N_6649,N_2216,N_1203);
and U6650 (N_6650,N_4429,N_3262);
nand U6651 (N_6651,N_4796,N_115);
xor U6652 (N_6652,N_704,N_2168);
and U6653 (N_6653,N_2436,N_3935);
and U6654 (N_6654,N_4070,N_990);
or U6655 (N_6655,N_3693,N_4214);
nand U6656 (N_6656,N_4999,N_338);
or U6657 (N_6657,N_4343,N_172);
or U6658 (N_6658,N_91,N_3126);
nor U6659 (N_6659,N_724,N_1101);
or U6660 (N_6660,N_2124,N_2104);
and U6661 (N_6661,N_3973,N_1071);
nor U6662 (N_6662,N_1829,N_3420);
nor U6663 (N_6663,N_2487,N_1596);
nand U6664 (N_6664,N_4814,N_3449);
or U6665 (N_6665,N_4405,N_1460);
nand U6666 (N_6666,N_3276,N_684);
or U6667 (N_6667,N_4641,N_507);
or U6668 (N_6668,N_4532,N_4374);
xor U6669 (N_6669,N_3113,N_2682);
or U6670 (N_6670,N_1984,N_2647);
nand U6671 (N_6671,N_4363,N_2139);
xor U6672 (N_6672,N_4179,N_4090);
xnor U6673 (N_6673,N_133,N_1965);
xor U6674 (N_6674,N_3005,N_98);
or U6675 (N_6675,N_2618,N_973);
or U6676 (N_6676,N_1191,N_129);
nor U6677 (N_6677,N_3400,N_1426);
and U6678 (N_6678,N_3549,N_4821);
xnor U6679 (N_6679,N_4695,N_1671);
or U6680 (N_6680,N_422,N_2971);
or U6681 (N_6681,N_4660,N_3168);
or U6682 (N_6682,N_2597,N_3559);
or U6683 (N_6683,N_1987,N_2573);
nor U6684 (N_6684,N_443,N_662);
nand U6685 (N_6685,N_52,N_2848);
nor U6686 (N_6686,N_1934,N_4974);
and U6687 (N_6687,N_352,N_3357);
nor U6688 (N_6688,N_1853,N_318);
and U6689 (N_6689,N_554,N_249);
nor U6690 (N_6690,N_1425,N_2423);
xnor U6691 (N_6691,N_705,N_4558);
xnor U6692 (N_6692,N_3094,N_1768);
and U6693 (N_6693,N_4593,N_3630);
nand U6694 (N_6694,N_45,N_1382);
or U6695 (N_6695,N_2544,N_4988);
nand U6696 (N_6696,N_4406,N_399);
nand U6697 (N_6697,N_3655,N_2242);
xor U6698 (N_6698,N_3020,N_3590);
xnor U6699 (N_6699,N_4782,N_3768);
nor U6700 (N_6700,N_871,N_669);
nand U6701 (N_6701,N_4524,N_4205);
and U6702 (N_6702,N_2149,N_415);
and U6703 (N_6703,N_1585,N_4904);
xnor U6704 (N_6704,N_3409,N_550);
and U6705 (N_6705,N_3957,N_4421);
nor U6706 (N_6706,N_213,N_3774);
xnor U6707 (N_6707,N_350,N_3710);
and U6708 (N_6708,N_1839,N_367);
and U6709 (N_6709,N_2333,N_1065);
and U6710 (N_6710,N_727,N_2175);
nor U6711 (N_6711,N_4166,N_944);
xor U6712 (N_6712,N_892,N_3015);
xor U6713 (N_6713,N_2338,N_3992);
nor U6714 (N_6714,N_1165,N_70);
nand U6715 (N_6715,N_4679,N_3572);
or U6716 (N_6716,N_565,N_947);
xnor U6717 (N_6717,N_3662,N_3014);
xor U6718 (N_6718,N_4718,N_3977);
and U6719 (N_6719,N_1090,N_2570);
xnor U6720 (N_6720,N_1884,N_4873);
xnor U6721 (N_6721,N_1263,N_3162);
nor U6722 (N_6722,N_456,N_1774);
or U6723 (N_6723,N_2189,N_1663);
xor U6724 (N_6724,N_2939,N_2691);
and U6725 (N_6725,N_2449,N_326);
and U6726 (N_6726,N_79,N_590);
xor U6727 (N_6727,N_1910,N_4236);
nor U6728 (N_6728,N_418,N_3512);
xor U6729 (N_6729,N_3714,N_955);
or U6730 (N_6730,N_2797,N_2096);
xor U6731 (N_6731,N_3330,N_518);
and U6732 (N_6732,N_1599,N_2715);
and U6733 (N_6733,N_829,N_1868);
xor U6734 (N_6734,N_2005,N_4570);
or U6735 (N_6735,N_2237,N_3969);
and U6736 (N_6736,N_4626,N_3596);
and U6737 (N_6737,N_1863,N_998);
nand U6738 (N_6738,N_539,N_847);
nor U6739 (N_6739,N_1333,N_1114);
or U6740 (N_6740,N_2810,N_1875);
xnor U6741 (N_6741,N_2294,N_3470);
nand U6742 (N_6742,N_1314,N_2505);
nor U6743 (N_6743,N_1522,N_1250);
nor U6744 (N_6744,N_2067,N_4361);
or U6745 (N_6745,N_1436,N_3455);
xnor U6746 (N_6746,N_3023,N_1854);
and U6747 (N_6747,N_1501,N_579);
and U6748 (N_6748,N_2381,N_3742);
or U6749 (N_6749,N_4838,N_3439);
nand U6750 (N_6750,N_2637,N_2707);
or U6751 (N_6751,N_2772,N_4311);
nand U6752 (N_6752,N_3481,N_760);
and U6753 (N_6753,N_4165,N_1817);
and U6754 (N_6754,N_1374,N_685);
nor U6755 (N_6755,N_3392,N_769);
and U6756 (N_6756,N_3064,N_583);
nand U6757 (N_6757,N_2824,N_4110);
or U6758 (N_6758,N_3024,N_4449);
nand U6759 (N_6759,N_2412,N_982);
nor U6760 (N_6760,N_980,N_4816);
or U6761 (N_6761,N_2108,N_1424);
nor U6762 (N_6762,N_1033,N_277);
nor U6763 (N_6763,N_2842,N_3099);
nor U6764 (N_6764,N_3309,N_3776);
nand U6765 (N_6765,N_1034,N_4804);
and U6766 (N_6766,N_1828,N_4083);
nor U6767 (N_6767,N_3633,N_1622);
nor U6768 (N_6768,N_715,N_4592);
or U6769 (N_6769,N_4628,N_801);
nand U6770 (N_6770,N_502,N_3391);
xor U6771 (N_6771,N_1168,N_2526);
nand U6772 (N_6772,N_3840,N_4450);
xnor U6773 (N_6773,N_3454,N_4465);
nor U6774 (N_6774,N_330,N_3665);
and U6775 (N_6775,N_3854,N_3568);
xor U6776 (N_6776,N_1651,N_3732);
and U6777 (N_6777,N_4092,N_3244);
nor U6778 (N_6778,N_370,N_299);
nand U6779 (N_6779,N_1192,N_402);
and U6780 (N_6780,N_2432,N_1353);
nand U6781 (N_6781,N_2093,N_1017);
nand U6782 (N_6782,N_3197,N_846);
xnor U6783 (N_6783,N_3622,N_3947);
or U6784 (N_6784,N_2308,N_3352);
nand U6785 (N_6785,N_3388,N_4281);
xnor U6786 (N_6786,N_4729,N_2358);
or U6787 (N_6787,N_3853,N_933);
xnor U6788 (N_6788,N_3834,N_4391);
xnor U6789 (N_6789,N_4479,N_2057);
or U6790 (N_6790,N_3960,N_4249);
xor U6791 (N_6791,N_4941,N_3074);
xnor U6792 (N_6792,N_2464,N_2809);
and U6793 (N_6793,N_2445,N_3961);
nand U6794 (N_6794,N_2839,N_2819);
and U6795 (N_6795,N_4467,N_1014);
or U6796 (N_6796,N_4373,N_4740);
nand U6797 (N_6797,N_4691,N_1513);
nand U6798 (N_6798,N_3008,N_1798);
or U6799 (N_6799,N_4607,N_1737);
or U6800 (N_6800,N_4522,N_3657);
or U6801 (N_6801,N_4697,N_2069);
xor U6802 (N_6802,N_3226,N_4829);
xor U6803 (N_6803,N_2833,N_3334);
nor U6804 (N_6804,N_1100,N_2849);
nor U6805 (N_6805,N_3269,N_4586);
nand U6806 (N_6806,N_792,N_713);
nor U6807 (N_6807,N_410,N_2210);
or U6808 (N_6808,N_3117,N_1525);
and U6809 (N_6809,N_3652,N_4696);
nor U6810 (N_6810,N_2183,N_1664);
nand U6811 (N_6811,N_1956,N_2347);
and U6812 (N_6812,N_4565,N_2152);
and U6813 (N_6813,N_4783,N_1031);
nand U6814 (N_6814,N_3542,N_4893);
nand U6815 (N_6815,N_334,N_4314);
nand U6816 (N_6816,N_3184,N_4792);
nand U6817 (N_6817,N_4137,N_2949);
nand U6818 (N_6818,N_3077,N_520);
xor U6819 (N_6819,N_2138,N_2163);
nor U6820 (N_6820,N_3042,N_770);
or U6821 (N_6821,N_1961,N_1296);
or U6822 (N_6822,N_1222,N_389);
nand U6823 (N_6823,N_1969,N_2558);
nand U6824 (N_6824,N_3651,N_4158);
nand U6825 (N_6825,N_1572,N_337);
and U6826 (N_6826,N_1407,N_592);
xnor U6827 (N_6827,N_2693,N_2258);
or U6828 (N_6828,N_2388,N_4580);
xnor U6829 (N_6829,N_4704,N_889);
and U6830 (N_6830,N_2114,N_3892);
and U6831 (N_6831,N_4143,N_1901);
xor U6832 (N_6832,N_65,N_3280);
xor U6833 (N_6833,N_4809,N_1384);
and U6834 (N_6834,N_2295,N_885);
nor U6835 (N_6835,N_1108,N_3893);
and U6836 (N_6836,N_1003,N_2002);
nor U6837 (N_6837,N_218,N_4531);
or U6838 (N_6838,N_2771,N_1209);
nor U6839 (N_6839,N_1403,N_3080);
nand U6840 (N_6840,N_822,N_1392);
or U6841 (N_6841,N_1354,N_1588);
nand U6842 (N_6842,N_2916,N_2243);
and U6843 (N_6843,N_1786,N_4614);
nand U6844 (N_6844,N_3644,N_1044);
or U6845 (N_6845,N_66,N_4407);
nor U6846 (N_6846,N_59,N_4251);
nor U6847 (N_6847,N_843,N_3856);
nand U6848 (N_6848,N_3394,N_1372);
nor U6849 (N_6849,N_1084,N_3465);
nand U6850 (N_6850,N_4989,N_3809);
nor U6851 (N_6851,N_4978,N_1826);
or U6852 (N_6852,N_2856,N_1143);
or U6853 (N_6853,N_4778,N_374);
xor U6854 (N_6854,N_4424,N_3311);
nand U6855 (N_6855,N_3772,N_2920);
or U6856 (N_6856,N_661,N_4505);
nor U6857 (N_6857,N_4549,N_3576);
and U6858 (N_6858,N_522,N_495);
or U6859 (N_6859,N_4618,N_4544);
nor U6860 (N_6860,N_3011,N_968);
and U6861 (N_6861,N_174,N_3794);
or U6862 (N_6862,N_1960,N_1950);
or U6863 (N_6863,N_3900,N_1059);
nor U6864 (N_6864,N_4658,N_3001);
xor U6865 (N_6865,N_3110,N_1119);
or U6866 (N_6866,N_1170,N_236);
nand U6867 (N_6867,N_2199,N_4160);
nor U6868 (N_6868,N_1796,N_4833);
nand U6869 (N_6869,N_2520,N_151);
nor U6870 (N_6870,N_2259,N_3713);
or U6871 (N_6871,N_4268,N_627);
and U6872 (N_6872,N_1789,N_248);
nand U6873 (N_6873,N_251,N_4438);
nor U6874 (N_6874,N_686,N_959);
or U6875 (N_6875,N_3183,N_4678);
and U6876 (N_6876,N_3049,N_3715);
nand U6877 (N_6877,N_1924,N_1217);
nor U6878 (N_6878,N_4286,N_239);
nor U6879 (N_6879,N_2063,N_3571);
nor U6880 (N_6880,N_4119,N_1809);
or U6881 (N_6881,N_3174,N_3760);
and U6882 (N_6882,N_4388,N_1069);
or U6883 (N_6883,N_3733,N_4380);
and U6884 (N_6884,N_2202,N_4849);
or U6885 (N_6885,N_4100,N_1928);
xnor U6886 (N_6886,N_2328,N_1689);
nor U6887 (N_6887,N_3027,N_3787);
xnor U6888 (N_6888,N_2465,N_941);
xnor U6889 (N_6889,N_1092,N_2941);
nor U6890 (N_6890,N_2600,N_3544);
or U6891 (N_6891,N_1063,N_3582);
nor U6892 (N_6892,N_2532,N_4007);
xor U6893 (N_6893,N_173,N_4195);
or U6894 (N_6894,N_3471,N_297);
or U6895 (N_6895,N_1595,N_3486);
nand U6896 (N_6896,N_3865,N_4313);
nand U6897 (N_6897,N_4386,N_3579);
nor U6898 (N_6898,N_4345,N_3306);
or U6899 (N_6899,N_798,N_4937);
nand U6900 (N_6900,N_186,N_4613);
nand U6901 (N_6901,N_1979,N_631);
nand U6902 (N_6902,N_1801,N_3201);
nor U6903 (N_6903,N_1270,N_1305);
or U6904 (N_6904,N_77,N_467);
nor U6905 (N_6905,N_492,N_746);
and U6906 (N_6906,N_2484,N_4252);
nand U6907 (N_6907,N_3498,N_4996);
nand U6908 (N_6908,N_4514,N_1345);
xnor U6909 (N_6909,N_3748,N_2281);
nand U6910 (N_6910,N_2081,N_1134);
or U6911 (N_6911,N_94,N_4553);
or U6912 (N_6912,N_3092,N_459);
nand U6913 (N_6913,N_1431,N_844);
xnor U6914 (N_6914,N_1409,N_634);
nand U6915 (N_6915,N_747,N_3150);
nor U6916 (N_6916,N_1793,N_4576);
or U6917 (N_6917,N_4659,N_1586);
or U6918 (N_6918,N_559,N_3717);
nand U6919 (N_6919,N_3610,N_3267);
nor U6920 (N_6920,N_1949,N_4423);
nor U6921 (N_6921,N_974,N_4180);
xnor U6922 (N_6922,N_4283,N_4732);
and U6923 (N_6923,N_585,N_1152);
or U6924 (N_6924,N_1125,N_2408);
or U6925 (N_6925,N_2828,N_2566);
nand U6926 (N_6926,N_2072,N_1007);
or U6927 (N_6927,N_3320,N_637);
xor U6928 (N_6928,N_2831,N_3569);
and U6929 (N_6929,N_4666,N_894);
and U6930 (N_6930,N_2252,N_198);
and U6931 (N_6931,N_2297,N_1299);
nand U6932 (N_6932,N_931,N_3835);
xor U6933 (N_6933,N_2954,N_396);
nand U6934 (N_6934,N_830,N_3090);
nand U6935 (N_6935,N_1204,N_3667);
or U6936 (N_6936,N_1118,N_1516);
xnor U6937 (N_6937,N_4392,N_3976);
nand U6938 (N_6938,N_2798,N_1615);
xnor U6939 (N_6939,N_1050,N_2840);
nand U6940 (N_6940,N_984,N_534);
or U6941 (N_6941,N_4749,N_3239);
or U6942 (N_6942,N_3249,N_3915);
nor U6943 (N_6943,N_2924,N_3425);
xnor U6944 (N_6944,N_4410,N_1665);
xor U6945 (N_6945,N_2056,N_1749);
nor U6946 (N_6946,N_1830,N_802);
and U6947 (N_6947,N_2626,N_4559);
xnor U6948 (N_6948,N_679,N_743);
xor U6949 (N_6949,N_2657,N_1998);
or U6950 (N_6950,N_600,N_1258);
nor U6951 (N_6951,N_156,N_3534);
or U6952 (N_6952,N_896,N_516);
nor U6953 (N_6953,N_2895,N_3050);
nor U6954 (N_6954,N_3848,N_2309);
nor U6955 (N_6955,N_2026,N_2433);
nor U6956 (N_6956,N_1348,N_1931);
or U6957 (N_6957,N_1682,N_3107);
and U6958 (N_6958,N_1137,N_2330);
and U6959 (N_6959,N_1194,N_1337);
or U6960 (N_6960,N_2235,N_3238);
or U6961 (N_6961,N_4785,N_2128);
and U6962 (N_6962,N_1478,N_279);
and U6963 (N_6963,N_64,N_2356);
nor U6964 (N_6964,N_4715,N_2734);
xnor U6965 (N_6965,N_768,N_2337);
and U6966 (N_6966,N_3043,N_1794);
xor U6967 (N_6967,N_4130,N_868);
and U6968 (N_6968,N_521,N_4887);
nand U6969 (N_6969,N_2548,N_3847);
and U6970 (N_6970,N_2088,N_653);
xor U6971 (N_6971,N_4900,N_575);
or U6972 (N_6972,N_1549,N_2627);
or U6973 (N_6973,N_3046,N_3432);
nor U6974 (N_6974,N_204,N_2413);
nor U6975 (N_6975,N_4510,N_2339);
xor U6976 (N_6976,N_1024,N_4837);
nand U6977 (N_6977,N_3731,N_258);
nor U6978 (N_6978,N_4271,N_2754);
xnor U6979 (N_6979,N_4288,N_252);
xnor U6980 (N_6980,N_3778,N_909);
and U6981 (N_6981,N_3602,N_4444);
nor U6982 (N_6982,N_1618,N_1660);
and U6983 (N_6983,N_2733,N_3302);
nor U6984 (N_6984,N_4480,N_63);
xnor U6985 (N_6985,N_4434,N_4506);
nand U6986 (N_6986,N_4956,N_1093);
or U6987 (N_6987,N_1527,N_331);
and U6988 (N_6988,N_2435,N_1268);
and U6989 (N_6989,N_2322,N_3264);
xor U6990 (N_6990,N_4190,N_2524);
and U6991 (N_6991,N_215,N_4896);
nor U6992 (N_6992,N_2790,N_2375);
xor U6993 (N_6993,N_4898,N_907);
and U6994 (N_6994,N_4684,N_1013);
nor U6995 (N_6995,N_772,N_1976);
nor U6996 (N_6996,N_2327,N_4969);
nand U6997 (N_6997,N_1981,N_2064);
nand U6998 (N_6998,N_2182,N_4527);
nor U6999 (N_6999,N_92,N_4712);
nor U7000 (N_7000,N_3332,N_2711);
nand U7001 (N_7001,N_1835,N_136);
xnor U7002 (N_7002,N_2634,N_4624);
and U7003 (N_7003,N_3586,N_2366);
and U7004 (N_7004,N_3819,N_1328);
or U7005 (N_7005,N_615,N_4255);
and U7006 (N_7006,N_2504,N_4595);
xnor U7007 (N_7007,N_586,N_290);
nand U7008 (N_7008,N_2307,N_3537);
nand U7009 (N_7009,N_4047,N_3811);
nand U7010 (N_7010,N_1518,N_663);
and U7011 (N_7011,N_665,N_2508);
and U7012 (N_7012,N_2968,N_3886);
nor U7013 (N_7013,N_2229,N_309);
nand U7014 (N_7014,N_1441,N_2430);
xor U7015 (N_7015,N_3478,N_294);
and U7016 (N_7016,N_4509,N_2415);
nor U7017 (N_7017,N_17,N_3597);
xor U7018 (N_7018,N_3373,N_4957);
nor U7019 (N_7019,N_321,N_4107);
nand U7020 (N_7020,N_310,N_164);
nand U7021 (N_7021,N_1344,N_4340);
xor U7022 (N_7022,N_1224,N_2077);
or U7023 (N_7023,N_488,N_2659);
nand U7024 (N_7024,N_749,N_899);
nor U7025 (N_7025,N_4750,N_58);
and U7026 (N_7026,N_4039,N_4745);
nand U7027 (N_7027,N_3421,N_2387);
xor U7028 (N_7028,N_2868,N_597);
xnor U7029 (N_7029,N_2619,N_2180);
and U7030 (N_7030,N_313,N_699);
nand U7031 (N_7031,N_996,N_2065);
xor U7032 (N_7032,N_4498,N_1210);
nand U7033 (N_7033,N_948,N_4006);
xor U7034 (N_7034,N_4414,N_340);
or U7035 (N_7035,N_2193,N_647);
nor U7036 (N_7036,N_3528,N_4892);
nor U7037 (N_7037,N_3773,N_3281);
and U7038 (N_7038,N_1626,N_2313);
xor U7039 (N_7039,N_2738,N_4452);
nand U7040 (N_7040,N_1386,N_3383);
nand U7041 (N_7041,N_2545,N_2234);
nand U7042 (N_7042,N_4389,N_4652);
xnor U7043 (N_7043,N_2760,N_4958);
nor U7044 (N_7044,N_3832,N_730);
nand U7045 (N_7045,N_2370,N_3337);
nor U7046 (N_7046,N_1729,N_855);
and U7047 (N_7047,N_2476,N_233);
nand U7048 (N_7048,N_1557,N_4460);
or U7049 (N_7049,N_4,N_2925);
nand U7050 (N_7050,N_891,N_3252);
or U7051 (N_7051,N_3591,N_4005);
xnor U7052 (N_7052,N_1983,N_1903);
and U7053 (N_7053,N_4901,N_1459);
xor U7054 (N_7054,N_2684,N_2736);
or U7055 (N_7055,N_1001,N_86);
nand U7056 (N_7056,N_2276,N_2767);
xor U7057 (N_7057,N_3032,N_2636);
and U7058 (N_7058,N_879,N_3546);
or U7059 (N_7059,N_1827,N_4167);
xnor U7060 (N_7060,N_2669,N_4023);
nor U7061 (N_7061,N_3203,N_2746);
or U7062 (N_7062,N_2661,N_4492);
and U7063 (N_7063,N_3754,N_4202);
nor U7064 (N_7064,N_965,N_2428);
or U7065 (N_7065,N_1852,N_1186);
nand U7066 (N_7066,N_315,N_1310);
nand U7067 (N_7067,N_2326,N_1632);
xor U7068 (N_7068,N_3210,N_3607);
or U7069 (N_7069,N_2934,N_2499);
nor U7070 (N_7070,N_4698,N_2725);
nor U7071 (N_7071,N_2488,N_4644);
or U7072 (N_7072,N_4072,N_3815);
xnor U7073 (N_7073,N_2290,N_3843);
or U7074 (N_7074,N_4681,N_783);
nand U7075 (N_7075,N_1946,N_1847);
nand U7076 (N_7076,N_2222,N_1921);
and U7077 (N_7077,N_212,N_831);
xor U7078 (N_7078,N_2039,N_2795);
nor U7079 (N_7079,N_3683,N_4367);
or U7080 (N_7080,N_4106,N_4512);
nand U7081 (N_7081,N_2473,N_4566);
or U7082 (N_7082,N_3279,N_1451);
nand U7083 (N_7083,N_1433,N_3038);
and U7084 (N_7084,N_1568,N_4784);
nand U7085 (N_7085,N_73,N_2972);
or U7086 (N_7086,N_2475,N_274);
or U7087 (N_7087,N_1776,N_99);
xor U7088 (N_7088,N_3991,N_4010);
or U7089 (N_7089,N_1282,N_3966);
nand U7090 (N_7090,N_4117,N_4963);
nand U7091 (N_7091,N_4535,N_1836);
xor U7092 (N_7092,N_31,N_3604);
and U7093 (N_7093,N_2021,N_327);
nand U7094 (N_7094,N_1645,N_3213);
xor U7095 (N_7095,N_423,N_4303);
and U7096 (N_7096,N_3300,N_2751);
nand U7097 (N_7097,N_2945,N_2463);
or U7098 (N_7098,N_985,N_27);
or U7099 (N_7099,N_1739,N_3580);
nand U7100 (N_7100,N_1691,N_2776);
xor U7101 (N_7101,N_1098,N_1952);
and U7102 (N_7102,N_797,N_1294);
or U7103 (N_7103,N_1600,N_1220);
and U7104 (N_7104,N_1252,N_945);
xor U7105 (N_7105,N_622,N_3322);
or U7106 (N_7106,N_4730,N_1631);
xnor U7107 (N_7107,N_3100,N_3929);
and U7108 (N_7108,N_4124,N_3194);
and U7109 (N_7109,N_1199,N_1608);
xor U7110 (N_7110,N_21,N_296);
and U7111 (N_7111,N_4299,N_2995);
and U7112 (N_7112,N_4024,N_527);
and U7113 (N_7113,N_3412,N_3263);
nor U7114 (N_7114,N_914,N_3808);
xnor U7115 (N_7115,N_1883,N_3047);
nand U7116 (N_7116,N_3048,N_4456);
xor U7117 (N_7117,N_4775,N_4710);
nand U7118 (N_7118,N_3370,N_4029);
nor U7119 (N_7119,N_678,N_1238);
nand U7120 (N_7120,N_2422,N_4403);
xor U7121 (N_7121,N_4653,N_344);
and U7122 (N_7122,N_3963,N_4426);
xnor U7123 (N_7123,N_1799,N_4800);
xnor U7124 (N_7124,N_4308,N_4267);
nor U7125 (N_7125,N_3086,N_2480);
nor U7126 (N_7126,N_4412,N_4597);
nand U7127 (N_7127,N_2799,N_3476);
and U7128 (N_7128,N_1489,N_3389);
or U7129 (N_7129,N_1581,N_341);
or U7130 (N_7130,N_3656,N_4474);
or U7131 (N_7131,N_3477,N_373);
nand U7132 (N_7132,N_2731,N_3192);
or U7133 (N_7133,N_2090,N_477);
xnor U7134 (N_7134,N_2390,N_392);
nor U7135 (N_7135,N_794,N_2692);
xnor U7136 (N_7136,N_2253,N_1173);
and U7137 (N_7137,N_125,N_1844);
or U7138 (N_7138,N_264,N_1536);
and U7139 (N_7139,N_2624,N_4752);
xor U7140 (N_7140,N_2722,N_3260);
and U7141 (N_7141,N_4347,N_501);
and U7142 (N_7142,N_128,N_3646);
xnor U7143 (N_7143,N_4689,N_4126);
and U7144 (N_7144,N_34,N_2102);
nor U7145 (N_7145,N_1905,N_2635);
nand U7146 (N_7146,N_2986,N_4708);
nand U7147 (N_7147,N_3323,N_4668);
nor U7148 (N_7148,N_4805,N_4147);
nand U7149 (N_7149,N_765,N_1544);
nand U7150 (N_7150,N_2912,N_2406);
nand U7151 (N_7151,N_2296,N_2471);
or U7152 (N_7152,N_1808,N_2173);
xor U7153 (N_7153,N_88,N_1948);
or U7154 (N_7154,N_2315,N_2353);
xor U7155 (N_7155,N_3780,N_1543);
nand U7156 (N_7156,N_4953,N_3697);
xor U7157 (N_7157,N_1219,N_721);
nor U7158 (N_7158,N_4131,N_4757);
and U7159 (N_7159,N_1890,N_4955);
or U7160 (N_7160,N_3638,N_3723);
nor U7161 (N_7161,N_2495,N_2961);
and U7162 (N_7162,N_1604,N_3163);
xnor U7163 (N_7163,N_3988,N_1131);
and U7164 (N_7164,N_4930,N_2928);
nand U7165 (N_7165,N_2643,N_4155);
and U7166 (N_7166,N_2185,N_4546);
or U7167 (N_7167,N_2444,N_970);
nor U7168 (N_7168,N_491,N_3619);
and U7169 (N_7169,N_1276,N_2850);
nand U7170 (N_7170,N_1902,N_1109);
and U7171 (N_7171,N_3328,N_4764);
nand U7172 (N_7172,N_3513,N_2948);
nand U7173 (N_7173,N_1066,N_8);
nand U7174 (N_7174,N_2060,N_655);
nor U7175 (N_7175,N_2041,N_4439);
nand U7176 (N_7176,N_3489,N_3846);
nand U7177 (N_7177,N_3666,N_1551);
and U7178 (N_7178,N_3417,N_4705);
or U7179 (N_7179,N_241,N_1406);
nand U7180 (N_7180,N_3222,N_1169);
nor U7181 (N_7181,N_2675,N_1465);
nand U7182 (N_7182,N_2117,N_2749);
or U7183 (N_7183,N_1837,N_3018);
or U7184 (N_7184,N_2539,N_3728);
or U7185 (N_7185,N_719,N_3235);
and U7186 (N_7186,N_1470,N_2233);
nand U7187 (N_7187,N_4711,N_1741);
or U7188 (N_7188,N_2893,N_262);
or U7189 (N_7189,N_238,N_4987);
xor U7190 (N_7190,N_3823,N_3076);
or U7191 (N_7191,N_1368,N_3407);
or U7192 (N_7192,N_888,N_3360);
xor U7193 (N_7193,N_4102,N_3212);
or U7194 (N_7194,N_2958,N_2875);
or U7195 (N_7195,N_3593,N_2025);
or U7196 (N_7196,N_949,N_4453);
and U7197 (N_7197,N_2766,N_530);
nand U7198 (N_7198,N_3695,N_80);
nand U7199 (N_7199,N_1493,N_1051);
nor U7200 (N_7200,N_1341,N_2818);
and U7201 (N_7201,N_2286,N_2861);
or U7202 (N_7202,N_2985,N_1788);
and U7203 (N_7203,N_1393,N_2466);
or U7204 (N_7204,N_1494,N_3901);
and U7205 (N_7205,N_3872,N_4009);
nor U7206 (N_7206,N_3448,N_2987);
and U7207 (N_7207,N_4058,N_1685);
nor U7208 (N_7208,N_4935,N_920);
or U7209 (N_7209,N_4733,N_160);
nand U7210 (N_7210,N_1246,N_2393);
and U7211 (N_7211,N_2049,N_591);
nor U7212 (N_7212,N_3567,N_4159);
xnor U7213 (N_7213,N_3228,N_153);
nor U7214 (N_7214,N_4813,N_876);
nor U7215 (N_7215,N_771,N_3844);
and U7216 (N_7216,N_1978,N_69);
nor U7217 (N_7217,N_1725,N_2386);
nand U7218 (N_7218,N_234,N_3452);
and U7219 (N_7219,N_1381,N_1571);
nand U7220 (N_7220,N_4366,N_323);
nand U7221 (N_7221,N_2681,N_4448);
or U7222 (N_7222,N_445,N_4967);
xnor U7223 (N_7223,N_3061,N_692);
xnor U7224 (N_7224,N_4926,N_3909);
or U7225 (N_7225,N_1955,N_4933);
nor U7226 (N_7226,N_2947,N_1874);
xor U7227 (N_7227,N_3999,N_4744);
nand U7228 (N_7228,N_2481,N_3140);
and U7229 (N_7229,N_4680,N_1229);
nor U7230 (N_7230,N_799,N_3995);
xor U7231 (N_7231,N_3817,N_4173);
xnor U7232 (N_7232,N_1533,N_1845);
nand U7233 (N_7233,N_1514,N_809);
xnor U7234 (N_7234,N_3555,N_4801);
or U7235 (N_7235,N_1986,N_3469);
nor U7236 (N_7236,N_2249,N_2118);
nand U7237 (N_7237,N_1475,N_884);
and U7238 (N_7238,N_2631,N_936);
or U7239 (N_7239,N_3256,N_3305);
nor U7240 (N_7240,N_1920,N_1548);
nor U7241 (N_7241,N_2735,N_3674);
xnor U7242 (N_7242,N_1947,N_3367);
xnor U7243 (N_7243,N_3797,N_1869);
nor U7244 (N_7244,N_2198,N_4256);
and U7245 (N_7245,N_1666,N_3694);
or U7246 (N_7246,N_288,N_2782);
nor U7247 (N_7247,N_1446,N_3965);
nor U7248 (N_7248,N_4001,N_2974);
nand U7249 (N_7249,N_1995,N_2973);
xor U7250 (N_7250,N_4247,N_3149);
nor U7251 (N_7251,N_832,N_3948);
nand U7252 (N_7252,N_2205,N_4026);
nor U7253 (N_7253,N_2583,N_505);
nor U7254 (N_7254,N_718,N_4638);
or U7255 (N_7255,N_3261,N_2288);
xor U7256 (N_7256,N_229,N_1612);
or U7257 (N_7257,N_2598,N_1712);
nand U7258 (N_7258,N_778,N_2105);
or U7259 (N_7259,N_3896,N_938);
or U7260 (N_7260,N_3529,N_3505);
nand U7261 (N_7261,N_319,N_734);
or U7262 (N_7262,N_1091,N_4909);
or U7263 (N_7263,N_693,N_3143);
and U7264 (N_7264,N_3852,N_3378);
xor U7265 (N_7265,N_3930,N_2238);
or U7266 (N_7266,N_4362,N_3919);
xor U7267 (N_7267,N_2204,N_1427);
nand U7268 (N_7268,N_2510,N_2119);
or U7269 (N_7269,N_2220,N_1428);
and U7270 (N_7270,N_2821,N_3341);
or U7271 (N_7271,N_3675,N_4121);
xnor U7272 (N_7272,N_3446,N_1190);
nor U7273 (N_7273,N_3974,N_2377);
or U7274 (N_7274,N_4220,N_3250);
nor U7275 (N_7275,N_46,N_2576);
nor U7276 (N_7276,N_636,N_1765);
or U7277 (N_7277,N_336,N_1096);
nand U7278 (N_7278,N_1810,N_1162);
nand U7279 (N_7279,N_3232,N_4050);
nor U7280 (N_7280,N_4275,N_553);
or U7281 (N_7281,N_2409,N_4992);
nor U7282 (N_7282,N_629,N_2450);
and U7283 (N_7283,N_481,N_3167);
or U7284 (N_7284,N_4599,N_618);
or U7285 (N_7285,N_4693,N_2015);
nand U7286 (N_7286,N_2442,N_4781);
nor U7287 (N_7287,N_2651,N_2368);
and U7288 (N_7288,N_2365,N_2917);
or U7289 (N_7289,N_2780,N_4459);
or U7290 (N_7290,N_4168,N_1245);
and U7291 (N_7291,N_1773,N_444);
or U7292 (N_7292,N_2956,N_1812);
nand U7293 (N_7293,N_1375,N_2768);
nor U7294 (N_7294,N_1147,N_4844);
xor U7295 (N_7295,N_4127,N_403);
and U7296 (N_7296,N_2648,N_2217);
nand U7297 (N_7297,N_4134,N_384);
or U7298 (N_7298,N_2535,N_1248);
nand U7299 (N_7299,N_3379,N_1892);
and U7300 (N_7300,N_2835,N_1889);
nand U7301 (N_7301,N_3516,N_2155);
xor U7302 (N_7302,N_2601,N_3737);
or U7303 (N_7303,N_2147,N_4866);
and U7304 (N_7304,N_2967,N_4051);
and U7305 (N_7305,N_795,N_3433);
nand U7306 (N_7306,N_2236,N_1962);
nand U7307 (N_7307,N_3902,N_435);
nand U7308 (N_7308,N_2245,N_1107);
or U7309 (N_7309,N_1343,N_812);
or U7310 (N_7310,N_1659,N_1335);
nor U7311 (N_7311,N_3890,N_556);
or U7312 (N_7312,N_862,N_4502);
and U7313 (N_7313,N_1695,N_594);
nor U7314 (N_7314,N_4329,N_3363);
or U7315 (N_7315,N_4135,N_145);
or U7316 (N_7316,N_4443,N_397);
nor U7317 (N_7317,N_3458,N_1647);
xor U7318 (N_7318,N_3681,N_2024);
nor U7319 (N_7319,N_1538,N_1686);
xor U7320 (N_7320,N_2399,N_4761);
nor U7321 (N_7321,N_1999,N_1657);
xor U7322 (N_7322,N_674,N_1079);
and U7323 (N_7323,N_2525,N_2348);
and U7324 (N_7324,N_44,N_4348);
or U7325 (N_7325,N_3402,N_1744);
nand U7326 (N_7326,N_3839,N_1811);
or U7327 (N_7327,N_1457,N_4394);
xnor U7328 (N_7328,N_2688,N_3782);
and U7329 (N_7329,N_159,N_2699);
xor U7330 (N_7330,N_4924,N_4911);
xnor U7331 (N_7331,N_1872,N_4661);
xor U7332 (N_7332,N_4908,N_3509);
and U7333 (N_7333,N_2083,N_1404);
nand U7334 (N_7334,N_875,N_2000);
and U7335 (N_7335,N_4059,N_4445);
nor U7336 (N_7336,N_437,N_4501);
nor U7337 (N_7337,N_1991,N_1038);
and U7338 (N_7338,N_751,N_1885);
or U7339 (N_7339,N_4184,N_4619);
nand U7340 (N_7340,N_4451,N_3128);
or U7341 (N_7341,N_2244,N_1399);
xnor U7342 (N_7342,N_295,N_3767);
nand U7343 (N_7343,N_3888,N_2550);
nand U7344 (N_7344,N_2569,N_2232);
nand U7345 (N_7345,N_4095,N_3716);
or U7346 (N_7346,N_1207,N_3286);
nor U7347 (N_7347,N_2454,N_2073);
or U7348 (N_7348,N_3411,N_3026);
xnor U7349 (N_7349,N_1526,N_4154);
nand U7350 (N_7350,N_1239,N_4114);
nor U7351 (N_7351,N_4358,N_1225);
nor U7352 (N_7352,N_3739,N_2523);
nand U7353 (N_7353,N_2656,N_4191);
or U7354 (N_7354,N_2613,N_2876);
or U7355 (N_7355,N_1624,N_41);
nor U7356 (N_7356,N_4428,N_2325);
and U7357 (N_7357,N_398,N_775);
nor U7358 (N_7358,N_2565,N_1086);
nand U7359 (N_7359,N_3318,N_118);
xnor U7360 (N_7360,N_4494,N_2517);
or U7361 (N_7361,N_2515,N_2003);
nand U7362 (N_7362,N_1643,N_1300);
xor U7363 (N_7363,N_412,N_1251);
xnor U7364 (N_7364,N_4590,N_3444);
nand U7365 (N_7365,N_2774,N_3669);
or U7366 (N_7366,N_2937,N_1458);
xnor U7367 (N_7367,N_3487,N_4682);
nand U7368 (N_7368,N_2777,N_1349);
and U7369 (N_7369,N_785,N_2179);
nand U7370 (N_7370,N_2447,N_2144);
or U7371 (N_7371,N_4259,N_4706);
nand U7372 (N_7372,N_682,N_954);
nor U7373 (N_7373,N_1366,N_2394);
and U7374 (N_7374,N_3524,N_589);
nor U7375 (N_7375,N_951,N_687);
and U7376 (N_7376,N_1308,N_1116);
xor U7377 (N_7377,N_1352,N_3009);
or U7378 (N_7378,N_4402,N_3060);
and U7379 (N_7379,N_4643,N_1552);
nand U7380 (N_7380,N_2616,N_2231);
nor U7381 (N_7381,N_619,N_3304);
nor U7382 (N_7382,N_2251,N_1782);
xnor U7383 (N_7383,N_2513,N_4913);
and U7384 (N_7384,N_2882,N_2706);
and U7385 (N_7385,N_1980,N_1742);
nand U7386 (N_7386,N_2014,N_3557);
or U7387 (N_7387,N_4690,N_103);
xor U7388 (N_7388,N_4847,N_1383);
nand U7389 (N_7389,N_2306,N_3523);
or U7390 (N_7390,N_2462,N_433);
or U7391 (N_7391,N_1302,N_390);
nor U7392 (N_7392,N_3951,N_4079);
xnor U7393 (N_7393,N_671,N_1807);
xor U7394 (N_7394,N_670,N_3506);
xnor U7395 (N_7395,N_3157,N_2261);
xnor U7396 (N_7396,N_2427,N_2880);
and U7397 (N_7397,N_881,N_1718);
xor U7398 (N_7398,N_1378,N_2698);
or U7399 (N_7399,N_613,N_3178);
or U7400 (N_7400,N_1285,N_3735);
nor U7401 (N_7401,N_3907,N_683);
or U7402 (N_7402,N_163,N_1480);
or U7403 (N_7403,N_4713,N_4111);
nor U7404 (N_7404,N_4922,N_1678);
and U7405 (N_7405,N_3434,N_558);
or U7406 (N_7406,N_1336,N_930);
or U7407 (N_7407,N_2300,N_1023);
nand U7408 (N_7408,N_2341,N_265);
and U7409 (N_7409,N_3810,N_1623);
nor U7410 (N_7410,N_353,N_2870);
xnor U7411 (N_7411,N_107,N_3296);
or U7412 (N_7412,N_490,N_356);
nor U7413 (N_7413,N_1058,N_1189);
nor U7414 (N_7414,N_2606,N_1846);
or U7415 (N_7415,N_2927,N_201);
xnor U7416 (N_7416,N_2457,N_4929);
nand U7417 (N_7417,N_1779,N_3307);
nor U7418 (N_7418,N_3240,N_639);
nor U7419 (N_7419,N_4152,N_328);
nand U7420 (N_7420,N_1327,N_3160);
nor U7421 (N_7421,N_237,N_3314);
or U7422 (N_7422,N_4156,N_84);
nor U7423 (N_7423,N_1022,N_2521);
xnor U7424 (N_7424,N_93,N_3520);
nor U7425 (N_7425,N_3548,N_2562);
or U7426 (N_7426,N_3335,N_3431);
or U7427 (N_7427,N_3358,N_4962);
and U7428 (N_7428,N_50,N_476);
and U7429 (N_7429,N_1637,N_4068);
xor U7430 (N_7430,N_2556,N_4091);
nor U7431 (N_7431,N_372,N_4738);
xnor U7432 (N_7432,N_867,N_1212);
nor U7433 (N_7433,N_599,N_766);
and U7434 (N_7434,N_1539,N_2748);
nor U7435 (N_7435,N_3629,N_3702);
and U7436 (N_7436,N_4122,N_2195);
xnor U7437 (N_7437,N_1144,N_2509);
or U7438 (N_7438,N_3111,N_2257);
nor U7439 (N_7439,N_2519,N_447);
nor U7440 (N_7440,N_4086,N_866);
nor U7441 (N_7441,N_3641,N_3499);
and U7442 (N_7442,N_3628,N_2747);
xor U7443 (N_7443,N_2852,N_2211);
xnor U7444 (N_7444,N_102,N_269);
and U7445 (N_7445,N_1254,N_1411);
nor U7446 (N_7446,N_4497,N_1233);
and U7447 (N_7447,N_3906,N_3857);
nor U7448 (N_7448,N_320,N_393);
and U7449 (N_7449,N_2874,N_3000);
nor U7450 (N_7450,N_2042,N_2660);
or U7451 (N_7451,N_2167,N_3408);
xnor U7452 (N_7452,N_4133,N_3224);
nand U7453 (N_7453,N_4153,N_3836);
nor U7454 (N_7454,N_3211,N_4253);
xnor U7455 (N_7455,N_2610,N_2862);
nand U7456 (N_7456,N_4545,N_3708);
nor U7457 (N_7457,N_3243,N_208);
or U7458 (N_7458,N_1214,N_217);
nand U7459 (N_7459,N_3348,N_939);
xnor U7460 (N_7460,N_4234,N_975);
nand U7461 (N_7461,N_3351,N_280);
nor U7462 (N_7462,N_2599,N_1157);
and U7463 (N_7463,N_1584,N_2572);
xnor U7464 (N_7464,N_4894,N_3870);
and U7465 (N_7465,N_3112,N_1074);
nand U7466 (N_7466,N_4008,N_4756);
nor U7467 (N_7467,N_281,N_405);
xor U7468 (N_7468,N_2966,N_1356);
nor U7469 (N_7469,N_1002,N_4123);
nor U7470 (N_7470,N_3441,N_854);
xor U7471 (N_7471,N_1434,N_2490);
xnor U7472 (N_7472,N_657,N_3786);
and U7473 (N_7473,N_2857,N_196);
nand U7474 (N_7474,N_4189,N_1633);
xor U7475 (N_7475,N_3121,N_1146);
and U7476 (N_7476,N_3581,N_3289);
and U7477 (N_7477,N_2975,N_4877);
and U7478 (N_7478,N_2129,N_2752);
and U7479 (N_7479,N_3916,N_2166);
and U7480 (N_7480,N_1569,N_105);
nor U7481 (N_7481,N_3473,N_703);
nor U7482 (N_7482,N_1821,N_4462);
nor U7483 (N_7483,N_3861,N_1629);
or U7484 (N_7484,N_3877,N_2157);
xor U7485 (N_7485,N_1653,N_3627);
nor U7486 (N_7486,N_1227,N_4305);
nor U7487 (N_7487,N_1085,N_2542);
and U7488 (N_7488,N_1528,N_3917);
xnor U7489 (N_7489,N_1913,N_2115);
nand U7490 (N_7490,N_1142,N_3532);
nor U7491 (N_7491,N_4138,N_187);
or U7492 (N_7492,N_4397,N_3700);
xnor U7493 (N_7493,N_1105,N_2148);
xor U7494 (N_7494,N_332,N_4802);
or U7495 (N_7495,N_1197,N_2530);
or U7496 (N_7496,N_1256,N_2696);
nor U7497 (N_7497,N_3151,N_1550);
nor U7498 (N_7498,N_242,N_3216);
and U7499 (N_7499,N_967,N_1722);
or U7500 (N_7500,N_4566,N_4282);
nand U7501 (N_7501,N_2376,N_895);
nor U7502 (N_7502,N_1604,N_4612);
nor U7503 (N_7503,N_3902,N_136);
nand U7504 (N_7504,N_2851,N_897);
or U7505 (N_7505,N_2952,N_3519);
nor U7506 (N_7506,N_2515,N_319);
or U7507 (N_7507,N_4113,N_2985);
nor U7508 (N_7508,N_901,N_4561);
nor U7509 (N_7509,N_2459,N_1626);
nor U7510 (N_7510,N_4441,N_2874);
and U7511 (N_7511,N_927,N_3241);
or U7512 (N_7512,N_3334,N_4102);
and U7513 (N_7513,N_44,N_981);
and U7514 (N_7514,N_4503,N_4966);
nand U7515 (N_7515,N_3073,N_1168);
nand U7516 (N_7516,N_2584,N_1877);
nand U7517 (N_7517,N_297,N_98);
and U7518 (N_7518,N_668,N_2865);
or U7519 (N_7519,N_90,N_3480);
nand U7520 (N_7520,N_4891,N_3571);
and U7521 (N_7521,N_699,N_470);
or U7522 (N_7522,N_72,N_805);
nand U7523 (N_7523,N_4314,N_4819);
or U7524 (N_7524,N_1813,N_699);
and U7525 (N_7525,N_4463,N_3551);
or U7526 (N_7526,N_1177,N_2917);
nand U7527 (N_7527,N_4697,N_4246);
xnor U7528 (N_7528,N_4483,N_2725);
xnor U7529 (N_7529,N_3162,N_4088);
nand U7530 (N_7530,N_2740,N_3095);
or U7531 (N_7531,N_1134,N_1101);
nand U7532 (N_7532,N_560,N_1);
nand U7533 (N_7533,N_4224,N_4955);
nor U7534 (N_7534,N_3520,N_2172);
xnor U7535 (N_7535,N_166,N_516);
nor U7536 (N_7536,N_4505,N_2713);
nor U7537 (N_7537,N_474,N_4350);
nand U7538 (N_7538,N_51,N_3553);
nand U7539 (N_7539,N_728,N_3);
and U7540 (N_7540,N_1946,N_1229);
nor U7541 (N_7541,N_4839,N_3436);
xnor U7542 (N_7542,N_2116,N_3121);
nor U7543 (N_7543,N_201,N_3964);
or U7544 (N_7544,N_648,N_3184);
nor U7545 (N_7545,N_1435,N_1869);
nand U7546 (N_7546,N_1949,N_4728);
and U7547 (N_7547,N_100,N_4399);
and U7548 (N_7548,N_2891,N_4129);
nand U7549 (N_7549,N_4116,N_3331);
or U7550 (N_7550,N_958,N_997);
nand U7551 (N_7551,N_1159,N_3626);
and U7552 (N_7552,N_4334,N_2539);
and U7553 (N_7553,N_3795,N_1881);
nor U7554 (N_7554,N_3934,N_2807);
or U7555 (N_7555,N_4589,N_1051);
nand U7556 (N_7556,N_1921,N_2698);
or U7557 (N_7557,N_4940,N_4201);
and U7558 (N_7558,N_4647,N_2910);
nand U7559 (N_7559,N_2459,N_4304);
nand U7560 (N_7560,N_4153,N_2469);
or U7561 (N_7561,N_4353,N_3017);
or U7562 (N_7562,N_4977,N_3520);
and U7563 (N_7563,N_4626,N_1448);
xor U7564 (N_7564,N_4084,N_2740);
and U7565 (N_7565,N_1638,N_1994);
xor U7566 (N_7566,N_645,N_1143);
or U7567 (N_7567,N_926,N_3158);
nand U7568 (N_7568,N_2263,N_240);
nor U7569 (N_7569,N_626,N_4469);
xor U7570 (N_7570,N_1166,N_2680);
and U7571 (N_7571,N_869,N_4357);
nor U7572 (N_7572,N_1448,N_3005);
nand U7573 (N_7573,N_3772,N_2431);
nor U7574 (N_7574,N_103,N_4098);
nand U7575 (N_7575,N_2189,N_4974);
or U7576 (N_7576,N_1199,N_2856);
or U7577 (N_7577,N_3655,N_4943);
nand U7578 (N_7578,N_600,N_4939);
nor U7579 (N_7579,N_3932,N_2386);
or U7580 (N_7580,N_3050,N_2827);
xor U7581 (N_7581,N_3268,N_3313);
xnor U7582 (N_7582,N_3940,N_709);
and U7583 (N_7583,N_2445,N_2332);
xnor U7584 (N_7584,N_2906,N_317);
or U7585 (N_7585,N_3217,N_817);
and U7586 (N_7586,N_2198,N_4981);
nor U7587 (N_7587,N_1954,N_4829);
or U7588 (N_7588,N_945,N_891);
nor U7589 (N_7589,N_2606,N_1042);
and U7590 (N_7590,N_3976,N_943);
nand U7591 (N_7591,N_803,N_640);
nor U7592 (N_7592,N_4492,N_1385);
xor U7593 (N_7593,N_2277,N_3369);
and U7594 (N_7594,N_3885,N_501);
or U7595 (N_7595,N_2903,N_831);
xnor U7596 (N_7596,N_1075,N_12);
xnor U7597 (N_7597,N_1129,N_3036);
and U7598 (N_7598,N_1798,N_4919);
and U7599 (N_7599,N_4613,N_1088);
nor U7600 (N_7600,N_136,N_2483);
xor U7601 (N_7601,N_833,N_3989);
nor U7602 (N_7602,N_1045,N_1272);
or U7603 (N_7603,N_2465,N_3098);
nand U7604 (N_7604,N_4076,N_1218);
xor U7605 (N_7605,N_3042,N_2751);
nor U7606 (N_7606,N_3309,N_4602);
or U7607 (N_7607,N_1371,N_3498);
nor U7608 (N_7608,N_1405,N_4725);
or U7609 (N_7609,N_3041,N_564);
and U7610 (N_7610,N_1918,N_1344);
xor U7611 (N_7611,N_3896,N_671);
nor U7612 (N_7612,N_4543,N_1632);
xor U7613 (N_7613,N_1077,N_2274);
nor U7614 (N_7614,N_1445,N_2329);
nand U7615 (N_7615,N_2472,N_1533);
xor U7616 (N_7616,N_2411,N_1820);
xnor U7617 (N_7617,N_4340,N_2913);
or U7618 (N_7618,N_1460,N_3218);
nor U7619 (N_7619,N_2660,N_1308);
nor U7620 (N_7620,N_949,N_587);
and U7621 (N_7621,N_4511,N_2113);
xor U7622 (N_7622,N_4546,N_2162);
and U7623 (N_7623,N_3862,N_373);
nor U7624 (N_7624,N_3937,N_4455);
xor U7625 (N_7625,N_4013,N_1504);
nor U7626 (N_7626,N_2455,N_172);
or U7627 (N_7627,N_493,N_4898);
and U7628 (N_7628,N_4653,N_3494);
and U7629 (N_7629,N_1812,N_247);
nand U7630 (N_7630,N_4730,N_530);
or U7631 (N_7631,N_2371,N_1844);
and U7632 (N_7632,N_1204,N_4695);
nor U7633 (N_7633,N_2030,N_188);
xor U7634 (N_7634,N_169,N_2868);
or U7635 (N_7635,N_1641,N_4689);
or U7636 (N_7636,N_1472,N_4882);
and U7637 (N_7637,N_1362,N_2429);
xor U7638 (N_7638,N_3302,N_3864);
and U7639 (N_7639,N_3714,N_2546);
nor U7640 (N_7640,N_3122,N_189);
xnor U7641 (N_7641,N_4291,N_1999);
xor U7642 (N_7642,N_1472,N_747);
and U7643 (N_7643,N_4062,N_3220);
xnor U7644 (N_7644,N_1712,N_1524);
nor U7645 (N_7645,N_967,N_4734);
or U7646 (N_7646,N_4844,N_3884);
xor U7647 (N_7647,N_1573,N_578);
xnor U7648 (N_7648,N_1476,N_39);
or U7649 (N_7649,N_2765,N_4556);
nor U7650 (N_7650,N_4984,N_526);
or U7651 (N_7651,N_3506,N_2815);
nor U7652 (N_7652,N_2278,N_2532);
nand U7653 (N_7653,N_159,N_4818);
xnor U7654 (N_7654,N_3745,N_527);
and U7655 (N_7655,N_1560,N_3442);
and U7656 (N_7656,N_3110,N_3039);
and U7657 (N_7657,N_1417,N_663);
and U7658 (N_7658,N_3613,N_1438);
nor U7659 (N_7659,N_2511,N_4987);
xor U7660 (N_7660,N_3793,N_578);
nand U7661 (N_7661,N_757,N_1960);
or U7662 (N_7662,N_4729,N_963);
nor U7663 (N_7663,N_1962,N_2920);
and U7664 (N_7664,N_2052,N_2839);
or U7665 (N_7665,N_2319,N_2143);
or U7666 (N_7666,N_2991,N_4022);
and U7667 (N_7667,N_2949,N_2273);
xor U7668 (N_7668,N_4482,N_4166);
nor U7669 (N_7669,N_3420,N_435);
and U7670 (N_7670,N_2917,N_2424);
nor U7671 (N_7671,N_602,N_574);
xor U7672 (N_7672,N_597,N_1980);
xor U7673 (N_7673,N_4089,N_1286);
nand U7674 (N_7674,N_3764,N_4490);
and U7675 (N_7675,N_897,N_1219);
xnor U7676 (N_7676,N_1681,N_3847);
or U7677 (N_7677,N_4914,N_2378);
and U7678 (N_7678,N_661,N_1178);
and U7679 (N_7679,N_3556,N_485);
nor U7680 (N_7680,N_4029,N_3076);
nand U7681 (N_7681,N_723,N_2528);
nand U7682 (N_7682,N_1425,N_4153);
or U7683 (N_7683,N_3499,N_2697);
xor U7684 (N_7684,N_1678,N_4480);
and U7685 (N_7685,N_165,N_2472);
nand U7686 (N_7686,N_3087,N_2669);
xnor U7687 (N_7687,N_1772,N_2025);
nand U7688 (N_7688,N_3368,N_802);
xor U7689 (N_7689,N_958,N_3145);
nor U7690 (N_7690,N_4313,N_3269);
or U7691 (N_7691,N_2933,N_1453);
and U7692 (N_7692,N_2325,N_4842);
or U7693 (N_7693,N_3540,N_553);
nor U7694 (N_7694,N_4052,N_2879);
xor U7695 (N_7695,N_473,N_3130);
and U7696 (N_7696,N_3030,N_861);
xor U7697 (N_7697,N_1396,N_1225);
xor U7698 (N_7698,N_1996,N_593);
and U7699 (N_7699,N_1096,N_4675);
or U7700 (N_7700,N_4900,N_2493);
xnor U7701 (N_7701,N_3111,N_3156);
or U7702 (N_7702,N_3154,N_2229);
or U7703 (N_7703,N_587,N_3742);
xnor U7704 (N_7704,N_3703,N_1613);
xor U7705 (N_7705,N_558,N_3491);
nand U7706 (N_7706,N_118,N_3941);
xnor U7707 (N_7707,N_1602,N_1915);
xnor U7708 (N_7708,N_3163,N_2265);
nand U7709 (N_7709,N_4766,N_4096);
xor U7710 (N_7710,N_4453,N_3849);
or U7711 (N_7711,N_3797,N_3751);
nand U7712 (N_7712,N_1665,N_197);
or U7713 (N_7713,N_2803,N_3604);
nand U7714 (N_7714,N_3498,N_398);
nand U7715 (N_7715,N_135,N_2309);
nor U7716 (N_7716,N_3680,N_1769);
xnor U7717 (N_7717,N_1687,N_1798);
xor U7718 (N_7718,N_3697,N_3369);
xnor U7719 (N_7719,N_4244,N_2629);
nor U7720 (N_7720,N_100,N_4027);
xnor U7721 (N_7721,N_4016,N_3534);
and U7722 (N_7722,N_3607,N_3042);
nor U7723 (N_7723,N_1445,N_3587);
nand U7724 (N_7724,N_1854,N_3426);
xor U7725 (N_7725,N_4131,N_2934);
nor U7726 (N_7726,N_2116,N_2855);
nor U7727 (N_7727,N_3283,N_1286);
nand U7728 (N_7728,N_4845,N_3060);
nand U7729 (N_7729,N_4642,N_2623);
nor U7730 (N_7730,N_2399,N_2017);
and U7731 (N_7731,N_399,N_948);
nand U7732 (N_7732,N_4886,N_2965);
or U7733 (N_7733,N_2579,N_4894);
and U7734 (N_7734,N_2380,N_3944);
xor U7735 (N_7735,N_869,N_1676);
or U7736 (N_7736,N_3671,N_1297);
and U7737 (N_7737,N_515,N_4);
xor U7738 (N_7738,N_4442,N_338);
nor U7739 (N_7739,N_2010,N_3746);
nand U7740 (N_7740,N_4942,N_3524);
xor U7741 (N_7741,N_4819,N_2977);
nor U7742 (N_7742,N_3603,N_2663);
or U7743 (N_7743,N_113,N_66);
xor U7744 (N_7744,N_4549,N_47);
nand U7745 (N_7745,N_4973,N_4489);
xor U7746 (N_7746,N_151,N_1505);
and U7747 (N_7747,N_679,N_2466);
xor U7748 (N_7748,N_2174,N_4849);
and U7749 (N_7749,N_3312,N_1251);
nand U7750 (N_7750,N_1814,N_3762);
xnor U7751 (N_7751,N_2276,N_335);
nand U7752 (N_7752,N_2539,N_4259);
xnor U7753 (N_7753,N_1751,N_4203);
and U7754 (N_7754,N_4230,N_4222);
and U7755 (N_7755,N_985,N_4378);
or U7756 (N_7756,N_3139,N_679);
nor U7757 (N_7757,N_4403,N_436);
nor U7758 (N_7758,N_377,N_2893);
nand U7759 (N_7759,N_2747,N_2060);
xor U7760 (N_7760,N_4467,N_2832);
and U7761 (N_7761,N_1914,N_676);
nor U7762 (N_7762,N_953,N_2445);
nand U7763 (N_7763,N_2269,N_1346);
and U7764 (N_7764,N_519,N_4156);
nor U7765 (N_7765,N_269,N_501);
xor U7766 (N_7766,N_4320,N_2463);
and U7767 (N_7767,N_743,N_2912);
or U7768 (N_7768,N_4026,N_995);
nand U7769 (N_7769,N_3198,N_1335);
or U7770 (N_7770,N_1416,N_1036);
nand U7771 (N_7771,N_4984,N_4445);
or U7772 (N_7772,N_2933,N_268);
nor U7773 (N_7773,N_4827,N_1971);
xnor U7774 (N_7774,N_1094,N_2284);
xor U7775 (N_7775,N_3857,N_927);
xnor U7776 (N_7776,N_4026,N_1596);
nor U7777 (N_7777,N_3026,N_3075);
xor U7778 (N_7778,N_231,N_4356);
xnor U7779 (N_7779,N_4996,N_4587);
nor U7780 (N_7780,N_4547,N_609);
nor U7781 (N_7781,N_4821,N_2037);
and U7782 (N_7782,N_2360,N_4475);
or U7783 (N_7783,N_944,N_2334);
and U7784 (N_7784,N_284,N_4503);
or U7785 (N_7785,N_191,N_4935);
nand U7786 (N_7786,N_282,N_1768);
or U7787 (N_7787,N_1265,N_458);
and U7788 (N_7788,N_1741,N_1756);
or U7789 (N_7789,N_905,N_878);
nand U7790 (N_7790,N_2500,N_4546);
xnor U7791 (N_7791,N_3807,N_1248);
nor U7792 (N_7792,N_1549,N_3305);
nor U7793 (N_7793,N_374,N_2237);
or U7794 (N_7794,N_2407,N_3338);
nor U7795 (N_7795,N_1768,N_1401);
nor U7796 (N_7796,N_1393,N_4232);
or U7797 (N_7797,N_1243,N_4543);
nor U7798 (N_7798,N_3689,N_1184);
nor U7799 (N_7799,N_865,N_4957);
or U7800 (N_7800,N_4308,N_4064);
or U7801 (N_7801,N_4093,N_2850);
or U7802 (N_7802,N_466,N_1942);
nor U7803 (N_7803,N_2623,N_3168);
or U7804 (N_7804,N_2863,N_2838);
nor U7805 (N_7805,N_3528,N_1541);
or U7806 (N_7806,N_2773,N_3251);
nand U7807 (N_7807,N_1944,N_4992);
or U7808 (N_7808,N_2409,N_4886);
and U7809 (N_7809,N_2788,N_4110);
xor U7810 (N_7810,N_4589,N_2291);
xnor U7811 (N_7811,N_4092,N_2041);
xor U7812 (N_7812,N_65,N_1203);
or U7813 (N_7813,N_1291,N_1209);
xor U7814 (N_7814,N_1372,N_1110);
nand U7815 (N_7815,N_1635,N_2894);
nor U7816 (N_7816,N_3338,N_320);
and U7817 (N_7817,N_359,N_3107);
and U7818 (N_7818,N_2587,N_4991);
or U7819 (N_7819,N_2522,N_2917);
xor U7820 (N_7820,N_3293,N_307);
or U7821 (N_7821,N_3357,N_3959);
nor U7822 (N_7822,N_3464,N_2555);
or U7823 (N_7823,N_4674,N_3008);
nand U7824 (N_7824,N_3291,N_1079);
nand U7825 (N_7825,N_393,N_2343);
or U7826 (N_7826,N_4669,N_1821);
or U7827 (N_7827,N_4126,N_1451);
or U7828 (N_7828,N_4031,N_2054);
nor U7829 (N_7829,N_4503,N_378);
and U7830 (N_7830,N_3109,N_2546);
and U7831 (N_7831,N_4656,N_2309);
xor U7832 (N_7832,N_2772,N_53);
nor U7833 (N_7833,N_2441,N_1048);
and U7834 (N_7834,N_552,N_1698);
and U7835 (N_7835,N_669,N_2008);
or U7836 (N_7836,N_2556,N_4585);
xnor U7837 (N_7837,N_1900,N_2664);
xnor U7838 (N_7838,N_1777,N_4910);
or U7839 (N_7839,N_3558,N_4336);
xnor U7840 (N_7840,N_4543,N_4176);
xor U7841 (N_7841,N_4655,N_4654);
xnor U7842 (N_7842,N_3085,N_1269);
xnor U7843 (N_7843,N_147,N_1597);
xor U7844 (N_7844,N_4454,N_467);
nor U7845 (N_7845,N_3763,N_784);
xor U7846 (N_7846,N_667,N_3844);
nand U7847 (N_7847,N_2020,N_1582);
and U7848 (N_7848,N_4223,N_3948);
or U7849 (N_7849,N_2402,N_782);
and U7850 (N_7850,N_3676,N_1242);
nor U7851 (N_7851,N_2950,N_2467);
xor U7852 (N_7852,N_1730,N_3358);
nand U7853 (N_7853,N_3993,N_4024);
or U7854 (N_7854,N_1909,N_2082);
nor U7855 (N_7855,N_2922,N_3334);
nand U7856 (N_7856,N_1204,N_1023);
and U7857 (N_7857,N_1352,N_1234);
xor U7858 (N_7858,N_4939,N_2616);
or U7859 (N_7859,N_27,N_2644);
and U7860 (N_7860,N_4117,N_2135);
nand U7861 (N_7861,N_575,N_4521);
or U7862 (N_7862,N_2105,N_4714);
xnor U7863 (N_7863,N_3018,N_4892);
xor U7864 (N_7864,N_3313,N_129);
nand U7865 (N_7865,N_3973,N_1879);
and U7866 (N_7866,N_2930,N_57);
nand U7867 (N_7867,N_2777,N_1282);
nor U7868 (N_7868,N_3766,N_1635);
and U7869 (N_7869,N_1575,N_1033);
nor U7870 (N_7870,N_4286,N_3949);
nor U7871 (N_7871,N_1034,N_4430);
xor U7872 (N_7872,N_608,N_4766);
or U7873 (N_7873,N_4283,N_4684);
or U7874 (N_7874,N_1829,N_4403);
or U7875 (N_7875,N_4802,N_78);
and U7876 (N_7876,N_1557,N_4706);
nand U7877 (N_7877,N_734,N_468);
or U7878 (N_7878,N_571,N_836);
nor U7879 (N_7879,N_1884,N_2501);
and U7880 (N_7880,N_4052,N_4468);
and U7881 (N_7881,N_2926,N_1840);
nor U7882 (N_7882,N_3423,N_1916);
or U7883 (N_7883,N_2360,N_820);
and U7884 (N_7884,N_2657,N_1301);
nand U7885 (N_7885,N_183,N_2069);
and U7886 (N_7886,N_3982,N_212);
nor U7887 (N_7887,N_2769,N_4369);
xnor U7888 (N_7888,N_2385,N_3534);
xnor U7889 (N_7889,N_2067,N_2013);
nor U7890 (N_7890,N_4790,N_2131);
or U7891 (N_7891,N_1982,N_487);
and U7892 (N_7892,N_4445,N_3864);
and U7893 (N_7893,N_116,N_330);
nor U7894 (N_7894,N_2579,N_2804);
nand U7895 (N_7895,N_1893,N_90);
nor U7896 (N_7896,N_2802,N_4369);
or U7897 (N_7897,N_4668,N_222);
nand U7898 (N_7898,N_4220,N_338);
or U7899 (N_7899,N_2867,N_3423);
nor U7900 (N_7900,N_3528,N_4160);
nor U7901 (N_7901,N_1954,N_4278);
xnor U7902 (N_7902,N_2783,N_2816);
xnor U7903 (N_7903,N_2816,N_552);
xnor U7904 (N_7904,N_4135,N_4767);
and U7905 (N_7905,N_1349,N_1053);
or U7906 (N_7906,N_2345,N_4963);
or U7907 (N_7907,N_4685,N_2715);
and U7908 (N_7908,N_4010,N_3585);
or U7909 (N_7909,N_3939,N_3820);
xnor U7910 (N_7910,N_4167,N_2429);
nand U7911 (N_7911,N_630,N_3505);
and U7912 (N_7912,N_4802,N_698);
nand U7913 (N_7913,N_3812,N_4418);
xor U7914 (N_7914,N_3724,N_1507);
and U7915 (N_7915,N_237,N_2491);
or U7916 (N_7916,N_783,N_4216);
xor U7917 (N_7917,N_184,N_2313);
and U7918 (N_7918,N_4322,N_4414);
or U7919 (N_7919,N_2156,N_1548);
and U7920 (N_7920,N_3874,N_1316);
nand U7921 (N_7921,N_812,N_2819);
nor U7922 (N_7922,N_713,N_2255);
and U7923 (N_7923,N_3475,N_4219);
nor U7924 (N_7924,N_1919,N_3270);
and U7925 (N_7925,N_4132,N_1996);
nand U7926 (N_7926,N_3933,N_2526);
nand U7927 (N_7927,N_2287,N_1969);
nor U7928 (N_7928,N_1714,N_3985);
xnor U7929 (N_7929,N_4970,N_4843);
or U7930 (N_7930,N_37,N_1340);
nand U7931 (N_7931,N_742,N_2411);
xor U7932 (N_7932,N_4764,N_316);
or U7933 (N_7933,N_2335,N_748);
nand U7934 (N_7934,N_4375,N_3711);
or U7935 (N_7935,N_91,N_3569);
nand U7936 (N_7936,N_1754,N_2283);
xnor U7937 (N_7937,N_3658,N_1888);
nor U7938 (N_7938,N_1990,N_4574);
nand U7939 (N_7939,N_328,N_1490);
and U7940 (N_7940,N_2438,N_4264);
xnor U7941 (N_7941,N_1027,N_2807);
xnor U7942 (N_7942,N_698,N_1420);
and U7943 (N_7943,N_1472,N_2557);
or U7944 (N_7944,N_1504,N_2977);
and U7945 (N_7945,N_3495,N_2743);
and U7946 (N_7946,N_2914,N_2150);
nor U7947 (N_7947,N_2340,N_3558);
and U7948 (N_7948,N_1302,N_614);
and U7949 (N_7949,N_555,N_3911);
nand U7950 (N_7950,N_1305,N_3698);
nor U7951 (N_7951,N_390,N_3244);
or U7952 (N_7952,N_4101,N_2198);
nand U7953 (N_7953,N_3063,N_1505);
or U7954 (N_7954,N_4884,N_4771);
or U7955 (N_7955,N_404,N_595);
nor U7956 (N_7956,N_2976,N_1710);
nor U7957 (N_7957,N_2538,N_1266);
nor U7958 (N_7958,N_1317,N_4233);
xor U7959 (N_7959,N_4188,N_2992);
and U7960 (N_7960,N_4840,N_2532);
and U7961 (N_7961,N_1126,N_4477);
and U7962 (N_7962,N_1705,N_3371);
xnor U7963 (N_7963,N_546,N_3533);
or U7964 (N_7964,N_2912,N_1708);
nand U7965 (N_7965,N_3211,N_1157);
nor U7966 (N_7966,N_96,N_170);
and U7967 (N_7967,N_3977,N_2660);
xnor U7968 (N_7968,N_926,N_4284);
nor U7969 (N_7969,N_4878,N_2453);
and U7970 (N_7970,N_4664,N_3179);
xnor U7971 (N_7971,N_581,N_4595);
xnor U7972 (N_7972,N_2514,N_1780);
nor U7973 (N_7973,N_3455,N_4466);
nor U7974 (N_7974,N_3326,N_1913);
and U7975 (N_7975,N_3243,N_3253);
xor U7976 (N_7976,N_1465,N_2747);
nand U7977 (N_7977,N_2966,N_1758);
xnor U7978 (N_7978,N_74,N_4258);
or U7979 (N_7979,N_1272,N_1059);
xnor U7980 (N_7980,N_602,N_953);
or U7981 (N_7981,N_850,N_3853);
nand U7982 (N_7982,N_2805,N_2149);
nand U7983 (N_7983,N_4289,N_3017);
nand U7984 (N_7984,N_3583,N_2673);
or U7985 (N_7985,N_1998,N_89);
nand U7986 (N_7986,N_1454,N_4647);
and U7987 (N_7987,N_1831,N_4599);
and U7988 (N_7988,N_3795,N_2567);
nor U7989 (N_7989,N_3374,N_1227);
and U7990 (N_7990,N_4542,N_787);
nor U7991 (N_7991,N_1948,N_4662);
nand U7992 (N_7992,N_1663,N_487);
or U7993 (N_7993,N_4157,N_587);
nor U7994 (N_7994,N_1720,N_295);
or U7995 (N_7995,N_85,N_3418);
xnor U7996 (N_7996,N_2370,N_4603);
xor U7997 (N_7997,N_119,N_1949);
nand U7998 (N_7998,N_4899,N_840);
nor U7999 (N_7999,N_4393,N_1033);
nor U8000 (N_8000,N_4424,N_1174);
and U8001 (N_8001,N_1896,N_508);
and U8002 (N_8002,N_2753,N_1085);
nor U8003 (N_8003,N_4287,N_880);
or U8004 (N_8004,N_1976,N_1607);
xor U8005 (N_8005,N_4057,N_3298);
and U8006 (N_8006,N_749,N_1116);
or U8007 (N_8007,N_4534,N_418);
nand U8008 (N_8008,N_2988,N_18);
xor U8009 (N_8009,N_4656,N_1831);
and U8010 (N_8010,N_1604,N_2084);
nor U8011 (N_8011,N_1205,N_1017);
xor U8012 (N_8012,N_362,N_263);
nand U8013 (N_8013,N_3920,N_4196);
nor U8014 (N_8014,N_3093,N_916);
and U8015 (N_8015,N_1619,N_4934);
and U8016 (N_8016,N_3550,N_1751);
nor U8017 (N_8017,N_1311,N_1014);
xor U8018 (N_8018,N_2376,N_4450);
or U8019 (N_8019,N_1206,N_382);
nand U8020 (N_8020,N_1943,N_1968);
nor U8021 (N_8021,N_3497,N_2104);
nand U8022 (N_8022,N_1791,N_1767);
or U8023 (N_8023,N_616,N_3781);
nor U8024 (N_8024,N_123,N_2426);
xnor U8025 (N_8025,N_410,N_569);
xnor U8026 (N_8026,N_4065,N_866);
and U8027 (N_8027,N_4308,N_682);
or U8028 (N_8028,N_3913,N_4007);
and U8029 (N_8029,N_4629,N_1453);
nor U8030 (N_8030,N_4833,N_3687);
or U8031 (N_8031,N_1321,N_3771);
nor U8032 (N_8032,N_1279,N_3396);
and U8033 (N_8033,N_2627,N_820);
nor U8034 (N_8034,N_2827,N_2532);
nand U8035 (N_8035,N_2101,N_3658);
or U8036 (N_8036,N_2780,N_2829);
nand U8037 (N_8037,N_4558,N_1307);
xor U8038 (N_8038,N_326,N_4923);
nor U8039 (N_8039,N_608,N_4500);
or U8040 (N_8040,N_4211,N_1892);
or U8041 (N_8041,N_4449,N_537);
or U8042 (N_8042,N_180,N_2866);
or U8043 (N_8043,N_2369,N_4250);
xnor U8044 (N_8044,N_4160,N_352);
and U8045 (N_8045,N_380,N_295);
or U8046 (N_8046,N_4377,N_3765);
or U8047 (N_8047,N_1798,N_3150);
nor U8048 (N_8048,N_1320,N_3337);
and U8049 (N_8049,N_1091,N_649);
xnor U8050 (N_8050,N_3285,N_496);
nor U8051 (N_8051,N_2490,N_3751);
nor U8052 (N_8052,N_2418,N_4831);
nor U8053 (N_8053,N_2333,N_2998);
nor U8054 (N_8054,N_3159,N_2795);
nor U8055 (N_8055,N_3867,N_94);
nand U8056 (N_8056,N_4633,N_1272);
nand U8057 (N_8057,N_4375,N_596);
nand U8058 (N_8058,N_2610,N_27);
and U8059 (N_8059,N_710,N_560);
nor U8060 (N_8060,N_869,N_2576);
nor U8061 (N_8061,N_2148,N_1473);
or U8062 (N_8062,N_4109,N_1251);
or U8063 (N_8063,N_670,N_881);
and U8064 (N_8064,N_540,N_3232);
nand U8065 (N_8065,N_3666,N_2320);
nand U8066 (N_8066,N_148,N_3301);
xnor U8067 (N_8067,N_2855,N_3626);
xnor U8068 (N_8068,N_4263,N_2494);
or U8069 (N_8069,N_3450,N_2374);
or U8070 (N_8070,N_3716,N_3611);
and U8071 (N_8071,N_1714,N_2551);
nand U8072 (N_8072,N_2656,N_1541);
nand U8073 (N_8073,N_2749,N_580);
xnor U8074 (N_8074,N_518,N_3434);
or U8075 (N_8075,N_623,N_2137);
xor U8076 (N_8076,N_1849,N_415);
xor U8077 (N_8077,N_4432,N_4497);
nand U8078 (N_8078,N_2433,N_3152);
or U8079 (N_8079,N_780,N_248);
and U8080 (N_8080,N_2819,N_1999);
or U8081 (N_8081,N_1859,N_4080);
and U8082 (N_8082,N_3977,N_4242);
xor U8083 (N_8083,N_3721,N_3375);
and U8084 (N_8084,N_2672,N_2098);
and U8085 (N_8085,N_71,N_147);
nor U8086 (N_8086,N_1963,N_978);
nor U8087 (N_8087,N_2977,N_2146);
and U8088 (N_8088,N_4366,N_3734);
and U8089 (N_8089,N_3006,N_3403);
or U8090 (N_8090,N_3738,N_3439);
or U8091 (N_8091,N_730,N_2941);
xor U8092 (N_8092,N_1868,N_3677);
nand U8093 (N_8093,N_4185,N_849);
and U8094 (N_8094,N_1190,N_2471);
xnor U8095 (N_8095,N_1486,N_3257);
nand U8096 (N_8096,N_3934,N_1657);
xnor U8097 (N_8097,N_4024,N_2483);
and U8098 (N_8098,N_4736,N_533);
xor U8099 (N_8099,N_3219,N_747);
nor U8100 (N_8100,N_3845,N_567);
xnor U8101 (N_8101,N_1789,N_1883);
or U8102 (N_8102,N_2839,N_2949);
xnor U8103 (N_8103,N_3876,N_1658);
and U8104 (N_8104,N_3795,N_622);
and U8105 (N_8105,N_1607,N_1448);
and U8106 (N_8106,N_16,N_1560);
or U8107 (N_8107,N_4507,N_664);
nand U8108 (N_8108,N_905,N_3132);
and U8109 (N_8109,N_4225,N_3807);
nor U8110 (N_8110,N_3367,N_510);
or U8111 (N_8111,N_1382,N_3746);
and U8112 (N_8112,N_2103,N_1383);
nand U8113 (N_8113,N_161,N_2993);
xor U8114 (N_8114,N_4415,N_2659);
xnor U8115 (N_8115,N_1462,N_3853);
nor U8116 (N_8116,N_4184,N_1222);
nand U8117 (N_8117,N_2894,N_4245);
nand U8118 (N_8118,N_4791,N_4257);
or U8119 (N_8119,N_1018,N_3902);
nor U8120 (N_8120,N_339,N_4826);
nor U8121 (N_8121,N_1526,N_3257);
nor U8122 (N_8122,N_2992,N_3316);
or U8123 (N_8123,N_4795,N_2067);
and U8124 (N_8124,N_1783,N_3383);
nand U8125 (N_8125,N_2947,N_3587);
or U8126 (N_8126,N_2902,N_1948);
xnor U8127 (N_8127,N_2673,N_4199);
nor U8128 (N_8128,N_4756,N_3707);
xor U8129 (N_8129,N_296,N_4188);
or U8130 (N_8130,N_605,N_3169);
or U8131 (N_8131,N_4245,N_1398);
nand U8132 (N_8132,N_4798,N_3654);
or U8133 (N_8133,N_2330,N_1867);
and U8134 (N_8134,N_3397,N_2802);
or U8135 (N_8135,N_2945,N_3051);
xor U8136 (N_8136,N_2972,N_1905);
and U8137 (N_8137,N_3853,N_1620);
nor U8138 (N_8138,N_4845,N_4239);
and U8139 (N_8139,N_1209,N_228);
nand U8140 (N_8140,N_4331,N_2410);
and U8141 (N_8141,N_3823,N_3863);
and U8142 (N_8142,N_3648,N_3292);
nor U8143 (N_8143,N_3493,N_2786);
nand U8144 (N_8144,N_1199,N_1700);
nor U8145 (N_8145,N_4768,N_3162);
nor U8146 (N_8146,N_4169,N_4699);
xor U8147 (N_8147,N_779,N_4769);
nand U8148 (N_8148,N_476,N_3856);
and U8149 (N_8149,N_3465,N_2295);
nand U8150 (N_8150,N_3886,N_2864);
and U8151 (N_8151,N_4532,N_4662);
nand U8152 (N_8152,N_931,N_4946);
nand U8153 (N_8153,N_2442,N_1391);
xnor U8154 (N_8154,N_967,N_91);
xnor U8155 (N_8155,N_3807,N_1516);
or U8156 (N_8156,N_1894,N_3682);
nor U8157 (N_8157,N_3132,N_2579);
and U8158 (N_8158,N_851,N_893);
nor U8159 (N_8159,N_3854,N_4997);
xnor U8160 (N_8160,N_829,N_2171);
nand U8161 (N_8161,N_919,N_1141);
xnor U8162 (N_8162,N_702,N_854);
nor U8163 (N_8163,N_1650,N_3959);
and U8164 (N_8164,N_2933,N_3241);
xnor U8165 (N_8165,N_1088,N_3499);
and U8166 (N_8166,N_822,N_2333);
nor U8167 (N_8167,N_4753,N_3459);
nor U8168 (N_8168,N_4862,N_3417);
nor U8169 (N_8169,N_3235,N_2574);
and U8170 (N_8170,N_1050,N_1338);
nand U8171 (N_8171,N_1442,N_2292);
and U8172 (N_8172,N_94,N_3733);
or U8173 (N_8173,N_4910,N_3703);
and U8174 (N_8174,N_2768,N_82);
nand U8175 (N_8175,N_2143,N_1254);
nand U8176 (N_8176,N_4966,N_2751);
or U8177 (N_8177,N_2426,N_4698);
nor U8178 (N_8178,N_3598,N_986);
and U8179 (N_8179,N_1259,N_4908);
nor U8180 (N_8180,N_4578,N_4101);
and U8181 (N_8181,N_3942,N_1630);
and U8182 (N_8182,N_4790,N_4723);
or U8183 (N_8183,N_1545,N_3994);
and U8184 (N_8184,N_1287,N_767);
nand U8185 (N_8185,N_806,N_2574);
nand U8186 (N_8186,N_4045,N_4328);
nor U8187 (N_8187,N_4084,N_4140);
or U8188 (N_8188,N_4031,N_1978);
nand U8189 (N_8189,N_4021,N_3016);
nor U8190 (N_8190,N_3423,N_2486);
or U8191 (N_8191,N_1067,N_664);
or U8192 (N_8192,N_994,N_1332);
or U8193 (N_8193,N_4482,N_814);
and U8194 (N_8194,N_2921,N_2911);
and U8195 (N_8195,N_4361,N_636);
nor U8196 (N_8196,N_182,N_2235);
nor U8197 (N_8197,N_1743,N_1914);
nor U8198 (N_8198,N_3579,N_4087);
and U8199 (N_8199,N_2369,N_4047);
xnor U8200 (N_8200,N_3336,N_2794);
nand U8201 (N_8201,N_4072,N_1815);
or U8202 (N_8202,N_1237,N_821);
or U8203 (N_8203,N_4947,N_4374);
nand U8204 (N_8204,N_388,N_4742);
nor U8205 (N_8205,N_1245,N_2257);
nor U8206 (N_8206,N_197,N_3911);
nor U8207 (N_8207,N_1014,N_3014);
nor U8208 (N_8208,N_123,N_2749);
nor U8209 (N_8209,N_1597,N_173);
nor U8210 (N_8210,N_890,N_2056);
or U8211 (N_8211,N_966,N_3341);
and U8212 (N_8212,N_461,N_2668);
and U8213 (N_8213,N_318,N_500);
nand U8214 (N_8214,N_4522,N_1612);
or U8215 (N_8215,N_1504,N_1025);
or U8216 (N_8216,N_1045,N_2264);
or U8217 (N_8217,N_1928,N_585);
nor U8218 (N_8218,N_851,N_2627);
or U8219 (N_8219,N_4248,N_3630);
nor U8220 (N_8220,N_917,N_1107);
xor U8221 (N_8221,N_4248,N_1508);
xor U8222 (N_8222,N_1880,N_1853);
nand U8223 (N_8223,N_665,N_1888);
nor U8224 (N_8224,N_713,N_1537);
and U8225 (N_8225,N_2265,N_578);
or U8226 (N_8226,N_4149,N_2612);
nor U8227 (N_8227,N_2124,N_2950);
and U8228 (N_8228,N_2424,N_1163);
and U8229 (N_8229,N_121,N_2783);
and U8230 (N_8230,N_842,N_2644);
and U8231 (N_8231,N_2156,N_4838);
nand U8232 (N_8232,N_1102,N_4886);
or U8233 (N_8233,N_4995,N_2039);
xnor U8234 (N_8234,N_1791,N_1535);
and U8235 (N_8235,N_512,N_3179);
nor U8236 (N_8236,N_2297,N_4022);
nand U8237 (N_8237,N_3879,N_1688);
xnor U8238 (N_8238,N_49,N_4243);
nand U8239 (N_8239,N_792,N_3620);
and U8240 (N_8240,N_385,N_2985);
and U8241 (N_8241,N_476,N_817);
or U8242 (N_8242,N_1932,N_1083);
or U8243 (N_8243,N_4233,N_1037);
nor U8244 (N_8244,N_2365,N_1475);
nand U8245 (N_8245,N_2796,N_439);
or U8246 (N_8246,N_4583,N_310);
xor U8247 (N_8247,N_4201,N_3661);
or U8248 (N_8248,N_3183,N_1028);
xnor U8249 (N_8249,N_1735,N_739);
and U8250 (N_8250,N_1161,N_558);
or U8251 (N_8251,N_3635,N_1578);
nor U8252 (N_8252,N_630,N_3179);
xor U8253 (N_8253,N_1894,N_1749);
nor U8254 (N_8254,N_1269,N_4099);
xnor U8255 (N_8255,N_3053,N_926);
xor U8256 (N_8256,N_2673,N_1871);
xor U8257 (N_8257,N_4840,N_2058);
nor U8258 (N_8258,N_4355,N_904);
and U8259 (N_8259,N_1654,N_2749);
or U8260 (N_8260,N_4905,N_4065);
or U8261 (N_8261,N_30,N_3955);
xnor U8262 (N_8262,N_260,N_561);
xor U8263 (N_8263,N_777,N_3495);
xnor U8264 (N_8264,N_1256,N_2513);
and U8265 (N_8265,N_2392,N_4932);
xnor U8266 (N_8266,N_3667,N_2473);
xor U8267 (N_8267,N_107,N_1926);
nand U8268 (N_8268,N_2659,N_1501);
xor U8269 (N_8269,N_1686,N_3710);
or U8270 (N_8270,N_4054,N_988);
or U8271 (N_8271,N_1844,N_847);
xnor U8272 (N_8272,N_1237,N_1928);
xor U8273 (N_8273,N_2956,N_4318);
nand U8274 (N_8274,N_1269,N_3523);
nand U8275 (N_8275,N_3793,N_3233);
and U8276 (N_8276,N_2005,N_1141);
and U8277 (N_8277,N_2759,N_2856);
or U8278 (N_8278,N_195,N_4031);
and U8279 (N_8279,N_3705,N_1523);
xor U8280 (N_8280,N_4510,N_3642);
xor U8281 (N_8281,N_4761,N_1930);
and U8282 (N_8282,N_724,N_863);
nor U8283 (N_8283,N_800,N_1410);
xnor U8284 (N_8284,N_2407,N_3370);
and U8285 (N_8285,N_2107,N_3101);
nor U8286 (N_8286,N_1077,N_80);
nor U8287 (N_8287,N_4088,N_3308);
xor U8288 (N_8288,N_2729,N_1440);
xnor U8289 (N_8289,N_1674,N_583);
nand U8290 (N_8290,N_3381,N_3218);
xnor U8291 (N_8291,N_4451,N_2456);
xnor U8292 (N_8292,N_174,N_836);
nor U8293 (N_8293,N_4241,N_3965);
nand U8294 (N_8294,N_3099,N_4459);
nand U8295 (N_8295,N_3916,N_426);
nand U8296 (N_8296,N_1092,N_486);
and U8297 (N_8297,N_3764,N_3882);
and U8298 (N_8298,N_1280,N_3313);
nand U8299 (N_8299,N_213,N_3184);
nand U8300 (N_8300,N_4567,N_4893);
and U8301 (N_8301,N_2878,N_2074);
or U8302 (N_8302,N_605,N_3099);
and U8303 (N_8303,N_1282,N_3928);
nor U8304 (N_8304,N_2840,N_4742);
or U8305 (N_8305,N_1168,N_4929);
or U8306 (N_8306,N_1853,N_4933);
nor U8307 (N_8307,N_296,N_4805);
or U8308 (N_8308,N_560,N_849);
or U8309 (N_8309,N_149,N_173);
nand U8310 (N_8310,N_3390,N_1512);
nor U8311 (N_8311,N_2545,N_1347);
or U8312 (N_8312,N_53,N_1523);
nor U8313 (N_8313,N_4071,N_1171);
or U8314 (N_8314,N_4530,N_3097);
nand U8315 (N_8315,N_1386,N_3992);
and U8316 (N_8316,N_2032,N_3357);
and U8317 (N_8317,N_695,N_189);
xor U8318 (N_8318,N_641,N_2050);
nor U8319 (N_8319,N_188,N_3478);
nand U8320 (N_8320,N_2006,N_2535);
nand U8321 (N_8321,N_2568,N_4802);
and U8322 (N_8322,N_4294,N_103);
nor U8323 (N_8323,N_344,N_1983);
xor U8324 (N_8324,N_1344,N_3584);
nand U8325 (N_8325,N_1088,N_1889);
and U8326 (N_8326,N_1820,N_4554);
and U8327 (N_8327,N_4066,N_1763);
or U8328 (N_8328,N_627,N_2817);
and U8329 (N_8329,N_3801,N_801);
xor U8330 (N_8330,N_2799,N_4129);
xnor U8331 (N_8331,N_1565,N_763);
and U8332 (N_8332,N_689,N_4244);
and U8333 (N_8333,N_53,N_4920);
and U8334 (N_8334,N_4743,N_3240);
or U8335 (N_8335,N_4400,N_3274);
or U8336 (N_8336,N_2903,N_1897);
xnor U8337 (N_8337,N_827,N_3560);
nor U8338 (N_8338,N_2695,N_3281);
nor U8339 (N_8339,N_2284,N_3691);
nor U8340 (N_8340,N_1556,N_3277);
and U8341 (N_8341,N_3888,N_3125);
nand U8342 (N_8342,N_3357,N_928);
or U8343 (N_8343,N_4927,N_2328);
xnor U8344 (N_8344,N_60,N_722);
nand U8345 (N_8345,N_1899,N_500);
or U8346 (N_8346,N_3742,N_4233);
nor U8347 (N_8347,N_1444,N_211);
nand U8348 (N_8348,N_167,N_1223);
and U8349 (N_8349,N_2754,N_701);
and U8350 (N_8350,N_9,N_244);
nand U8351 (N_8351,N_1754,N_2721);
nand U8352 (N_8352,N_1023,N_1166);
xnor U8353 (N_8353,N_2808,N_4267);
and U8354 (N_8354,N_270,N_2804);
or U8355 (N_8355,N_1173,N_4645);
and U8356 (N_8356,N_1531,N_1077);
xnor U8357 (N_8357,N_2100,N_4055);
nor U8358 (N_8358,N_4281,N_1739);
nor U8359 (N_8359,N_3495,N_4483);
nand U8360 (N_8360,N_1493,N_2038);
nor U8361 (N_8361,N_4387,N_2055);
nor U8362 (N_8362,N_688,N_4532);
and U8363 (N_8363,N_251,N_4689);
nor U8364 (N_8364,N_43,N_3075);
nor U8365 (N_8365,N_2466,N_1981);
nand U8366 (N_8366,N_4322,N_4535);
xor U8367 (N_8367,N_3255,N_1720);
nand U8368 (N_8368,N_854,N_1812);
xnor U8369 (N_8369,N_4033,N_3614);
or U8370 (N_8370,N_1575,N_282);
xor U8371 (N_8371,N_1834,N_468);
or U8372 (N_8372,N_3941,N_2482);
nand U8373 (N_8373,N_21,N_4704);
and U8374 (N_8374,N_263,N_38);
and U8375 (N_8375,N_4657,N_2430);
xnor U8376 (N_8376,N_3032,N_630);
nor U8377 (N_8377,N_3436,N_709);
or U8378 (N_8378,N_1619,N_4782);
and U8379 (N_8379,N_4441,N_4890);
nand U8380 (N_8380,N_2637,N_386);
xnor U8381 (N_8381,N_911,N_0);
nand U8382 (N_8382,N_4659,N_1024);
nor U8383 (N_8383,N_3027,N_418);
nor U8384 (N_8384,N_4866,N_121);
nor U8385 (N_8385,N_33,N_4965);
nor U8386 (N_8386,N_2265,N_432);
xor U8387 (N_8387,N_1795,N_2261);
xnor U8388 (N_8388,N_3937,N_1301);
xnor U8389 (N_8389,N_1154,N_62);
xor U8390 (N_8390,N_4488,N_2430);
nor U8391 (N_8391,N_3251,N_188);
or U8392 (N_8392,N_1931,N_3654);
or U8393 (N_8393,N_3620,N_2371);
and U8394 (N_8394,N_2860,N_4835);
and U8395 (N_8395,N_4879,N_3280);
or U8396 (N_8396,N_1741,N_213);
xor U8397 (N_8397,N_4497,N_862);
and U8398 (N_8398,N_1727,N_2570);
nor U8399 (N_8399,N_2604,N_824);
or U8400 (N_8400,N_4144,N_4779);
nand U8401 (N_8401,N_2430,N_2799);
nand U8402 (N_8402,N_3683,N_2809);
and U8403 (N_8403,N_385,N_510);
nand U8404 (N_8404,N_1576,N_670);
and U8405 (N_8405,N_1614,N_4084);
nor U8406 (N_8406,N_908,N_2969);
nor U8407 (N_8407,N_739,N_1636);
or U8408 (N_8408,N_1583,N_963);
and U8409 (N_8409,N_2535,N_3324);
and U8410 (N_8410,N_138,N_1660);
xor U8411 (N_8411,N_4351,N_2272);
nor U8412 (N_8412,N_4966,N_1127);
and U8413 (N_8413,N_4158,N_4805);
xnor U8414 (N_8414,N_1528,N_46);
nor U8415 (N_8415,N_3300,N_28);
or U8416 (N_8416,N_4989,N_3468);
and U8417 (N_8417,N_3820,N_1535);
or U8418 (N_8418,N_2568,N_2514);
nor U8419 (N_8419,N_1320,N_3400);
and U8420 (N_8420,N_1167,N_4408);
nand U8421 (N_8421,N_2591,N_3785);
nand U8422 (N_8422,N_1196,N_2702);
and U8423 (N_8423,N_3057,N_2287);
and U8424 (N_8424,N_500,N_427);
and U8425 (N_8425,N_3433,N_2312);
nand U8426 (N_8426,N_3846,N_3268);
and U8427 (N_8427,N_1348,N_33);
or U8428 (N_8428,N_2710,N_2018);
and U8429 (N_8429,N_1566,N_848);
xnor U8430 (N_8430,N_4172,N_3252);
and U8431 (N_8431,N_4013,N_4934);
nor U8432 (N_8432,N_3768,N_3619);
nor U8433 (N_8433,N_2635,N_3534);
nand U8434 (N_8434,N_1376,N_33);
nor U8435 (N_8435,N_1651,N_485);
and U8436 (N_8436,N_2602,N_3806);
and U8437 (N_8437,N_4973,N_4578);
or U8438 (N_8438,N_1841,N_1129);
or U8439 (N_8439,N_2151,N_1250);
nand U8440 (N_8440,N_3669,N_283);
xnor U8441 (N_8441,N_6,N_1275);
nand U8442 (N_8442,N_2186,N_156);
xnor U8443 (N_8443,N_2501,N_2385);
nand U8444 (N_8444,N_2584,N_3473);
nor U8445 (N_8445,N_4142,N_828);
nor U8446 (N_8446,N_1636,N_4141);
nand U8447 (N_8447,N_3496,N_4303);
nand U8448 (N_8448,N_301,N_3152);
or U8449 (N_8449,N_1601,N_4191);
xor U8450 (N_8450,N_3993,N_246);
nor U8451 (N_8451,N_1641,N_2967);
or U8452 (N_8452,N_1970,N_2757);
and U8453 (N_8453,N_3706,N_2943);
nor U8454 (N_8454,N_1591,N_71);
and U8455 (N_8455,N_3523,N_783);
nand U8456 (N_8456,N_4622,N_3262);
and U8457 (N_8457,N_4033,N_2520);
nor U8458 (N_8458,N_3863,N_3084);
xor U8459 (N_8459,N_1287,N_2168);
nor U8460 (N_8460,N_1778,N_213);
or U8461 (N_8461,N_3716,N_2342);
nor U8462 (N_8462,N_4208,N_4986);
nand U8463 (N_8463,N_4329,N_3584);
xor U8464 (N_8464,N_4540,N_1305);
or U8465 (N_8465,N_256,N_992);
and U8466 (N_8466,N_1559,N_990);
nand U8467 (N_8467,N_284,N_2543);
nand U8468 (N_8468,N_3375,N_1574);
nand U8469 (N_8469,N_2818,N_2101);
or U8470 (N_8470,N_4911,N_2513);
xor U8471 (N_8471,N_1210,N_1216);
xor U8472 (N_8472,N_1833,N_4686);
or U8473 (N_8473,N_2632,N_2128);
xnor U8474 (N_8474,N_2861,N_1903);
or U8475 (N_8475,N_531,N_3002);
and U8476 (N_8476,N_3028,N_4164);
and U8477 (N_8477,N_2605,N_2642);
or U8478 (N_8478,N_3906,N_1983);
and U8479 (N_8479,N_4281,N_3229);
nand U8480 (N_8480,N_3619,N_4200);
or U8481 (N_8481,N_805,N_820);
nor U8482 (N_8482,N_2178,N_617);
or U8483 (N_8483,N_2139,N_3104);
nor U8484 (N_8484,N_302,N_1897);
nor U8485 (N_8485,N_4623,N_3757);
xor U8486 (N_8486,N_2903,N_1599);
and U8487 (N_8487,N_3037,N_1468);
nor U8488 (N_8488,N_574,N_1569);
and U8489 (N_8489,N_1075,N_4943);
and U8490 (N_8490,N_1106,N_1911);
nand U8491 (N_8491,N_962,N_174);
nor U8492 (N_8492,N_3995,N_841);
and U8493 (N_8493,N_2858,N_1524);
xor U8494 (N_8494,N_1772,N_3061);
xnor U8495 (N_8495,N_3048,N_1496);
or U8496 (N_8496,N_160,N_4329);
and U8497 (N_8497,N_1939,N_4166);
xor U8498 (N_8498,N_1662,N_537);
xor U8499 (N_8499,N_3769,N_3461);
xor U8500 (N_8500,N_4450,N_1673);
or U8501 (N_8501,N_3365,N_4864);
xor U8502 (N_8502,N_3504,N_3805);
nor U8503 (N_8503,N_2234,N_4931);
nand U8504 (N_8504,N_1801,N_4002);
and U8505 (N_8505,N_2530,N_2193);
nor U8506 (N_8506,N_2605,N_3898);
xor U8507 (N_8507,N_3951,N_2894);
xnor U8508 (N_8508,N_551,N_4397);
nand U8509 (N_8509,N_760,N_3017);
xnor U8510 (N_8510,N_1163,N_3444);
and U8511 (N_8511,N_786,N_4667);
and U8512 (N_8512,N_3621,N_3458);
nand U8513 (N_8513,N_2059,N_1441);
and U8514 (N_8514,N_34,N_1991);
or U8515 (N_8515,N_1006,N_4657);
xnor U8516 (N_8516,N_4016,N_2815);
nand U8517 (N_8517,N_123,N_1756);
and U8518 (N_8518,N_4539,N_3015);
or U8519 (N_8519,N_294,N_1474);
nor U8520 (N_8520,N_3037,N_4337);
nor U8521 (N_8521,N_1793,N_4905);
nand U8522 (N_8522,N_98,N_820);
xor U8523 (N_8523,N_1556,N_2769);
and U8524 (N_8524,N_3319,N_421);
nand U8525 (N_8525,N_2855,N_297);
xor U8526 (N_8526,N_439,N_3494);
nor U8527 (N_8527,N_3002,N_4080);
xnor U8528 (N_8528,N_416,N_1339);
nor U8529 (N_8529,N_419,N_737);
nor U8530 (N_8530,N_4041,N_4792);
nand U8531 (N_8531,N_827,N_1551);
nor U8532 (N_8532,N_2906,N_1476);
nand U8533 (N_8533,N_3690,N_4490);
xnor U8534 (N_8534,N_1237,N_2410);
or U8535 (N_8535,N_4037,N_1057);
nor U8536 (N_8536,N_3877,N_4764);
xnor U8537 (N_8537,N_3534,N_2823);
nand U8538 (N_8538,N_2223,N_1552);
nor U8539 (N_8539,N_3254,N_2685);
and U8540 (N_8540,N_1997,N_2358);
xor U8541 (N_8541,N_2503,N_1361);
nor U8542 (N_8542,N_3522,N_4089);
or U8543 (N_8543,N_3873,N_3031);
nor U8544 (N_8544,N_3256,N_3959);
xor U8545 (N_8545,N_890,N_584);
or U8546 (N_8546,N_148,N_3157);
and U8547 (N_8547,N_2029,N_144);
and U8548 (N_8548,N_232,N_2670);
nand U8549 (N_8549,N_3509,N_4505);
or U8550 (N_8550,N_2337,N_4982);
nor U8551 (N_8551,N_1580,N_1540);
nor U8552 (N_8552,N_2711,N_765);
or U8553 (N_8553,N_1400,N_3164);
nand U8554 (N_8554,N_1144,N_3195);
xnor U8555 (N_8555,N_2570,N_4772);
xor U8556 (N_8556,N_4125,N_360);
or U8557 (N_8557,N_1429,N_2864);
xor U8558 (N_8558,N_1807,N_356);
and U8559 (N_8559,N_2986,N_3718);
or U8560 (N_8560,N_2803,N_1506);
or U8561 (N_8561,N_4846,N_2869);
xor U8562 (N_8562,N_4892,N_896);
nor U8563 (N_8563,N_2596,N_1586);
or U8564 (N_8564,N_3688,N_1003);
nor U8565 (N_8565,N_3340,N_1193);
and U8566 (N_8566,N_2196,N_2016);
xor U8567 (N_8567,N_1440,N_2960);
xor U8568 (N_8568,N_10,N_2199);
and U8569 (N_8569,N_3216,N_4993);
and U8570 (N_8570,N_3742,N_3620);
and U8571 (N_8571,N_3670,N_4031);
and U8572 (N_8572,N_2241,N_2731);
and U8573 (N_8573,N_4425,N_2708);
and U8574 (N_8574,N_4758,N_3145);
or U8575 (N_8575,N_1594,N_4634);
and U8576 (N_8576,N_807,N_3089);
nor U8577 (N_8577,N_4060,N_722);
nor U8578 (N_8578,N_3114,N_2912);
xnor U8579 (N_8579,N_289,N_4507);
xnor U8580 (N_8580,N_1918,N_372);
or U8581 (N_8581,N_1658,N_3134);
and U8582 (N_8582,N_1491,N_3317);
nand U8583 (N_8583,N_431,N_3321);
or U8584 (N_8584,N_245,N_4892);
nand U8585 (N_8585,N_2943,N_1232);
nand U8586 (N_8586,N_414,N_167);
nand U8587 (N_8587,N_3868,N_4897);
and U8588 (N_8588,N_2024,N_2608);
and U8589 (N_8589,N_2631,N_979);
nor U8590 (N_8590,N_818,N_4189);
or U8591 (N_8591,N_3904,N_3894);
or U8592 (N_8592,N_4879,N_2232);
nor U8593 (N_8593,N_2670,N_177);
nor U8594 (N_8594,N_2942,N_4952);
nor U8595 (N_8595,N_2013,N_4756);
nor U8596 (N_8596,N_415,N_3894);
xor U8597 (N_8597,N_2147,N_1365);
or U8598 (N_8598,N_2256,N_4770);
xor U8599 (N_8599,N_2334,N_4023);
and U8600 (N_8600,N_2561,N_172);
xor U8601 (N_8601,N_2095,N_4705);
nand U8602 (N_8602,N_4839,N_1982);
and U8603 (N_8603,N_453,N_928);
or U8604 (N_8604,N_323,N_3402);
xor U8605 (N_8605,N_218,N_4955);
and U8606 (N_8606,N_3231,N_680);
or U8607 (N_8607,N_4150,N_4933);
xor U8608 (N_8608,N_4491,N_633);
nor U8609 (N_8609,N_2052,N_1379);
and U8610 (N_8610,N_1069,N_4118);
xnor U8611 (N_8611,N_2027,N_1144);
xnor U8612 (N_8612,N_2950,N_2038);
or U8613 (N_8613,N_4298,N_4989);
and U8614 (N_8614,N_4946,N_260);
or U8615 (N_8615,N_3539,N_2336);
xnor U8616 (N_8616,N_3297,N_4789);
or U8617 (N_8617,N_1186,N_617);
nor U8618 (N_8618,N_1112,N_3147);
and U8619 (N_8619,N_2081,N_4097);
nand U8620 (N_8620,N_3359,N_2610);
nor U8621 (N_8621,N_1025,N_4023);
nand U8622 (N_8622,N_4911,N_2152);
nor U8623 (N_8623,N_2179,N_4660);
or U8624 (N_8624,N_2085,N_3149);
nand U8625 (N_8625,N_4871,N_4455);
or U8626 (N_8626,N_2385,N_4046);
nand U8627 (N_8627,N_3445,N_2093);
xor U8628 (N_8628,N_199,N_842);
or U8629 (N_8629,N_2088,N_2906);
xor U8630 (N_8630,N_997,N_2847);
xor U8631 (N_8631,N_3591,N_1082);
nand U8632 (N_8632,N_2292,N_173);
xnor U8633 (N_8633,N_2546,N_1318);
nand U8634 (N_8634,N_997,N_920);
nand U8635 (N_8635,N_2210,N_4542);
or U8636 (N_8636,N_2598,N_854);
and U8637 (N_8637,N_2789,N_737);
nand U8638 (N_8638,N_2704,N_378);
nor U8639 (N_8639,N_1064,N_3413);
nand U8640 (N_8640,N_4793,N_1039);
nand U8641 (N_8641,N_340,N_3024);
nor U8642 (N_8642,N_2623,N_1654);
nand U8643 (N_8643,N_2472,N_3067);
xnor U8644 (N_8644,N_3628,N_4385);
nor U8645 (N_8645,N_4170,N_382);
nand U8646 (N_8646,N_1689,N_3108);
xnor U8647 (N_8647,N_2974,N_4844);
xnor U8648 (N_8648,N_4364,N_3062);
nor U8649 (N_8649,N_2582,N_2522);
and U8650 (N_8650,N_2660,N_2425);
or U8651 (N_8651,N_4879,N_1504);
and U8652 (N_8652,N_3786,N_2060);
or U8653 (N_8653,N_4361,N_2001);
nand U8654 (N_8654,N_3586,N_2672);
nand U8655 (N_8655,N_3757,N_1455);
nor U8656 (N_8656,N_1797,N_176);
nand U8657 (N_8657,N_3034,N_897);
and U8658 (N_8658,N_4323,N_4812);
nand U8659 (N_8659,N_3454,N_3335);
nand U8660 (N_8660,N_1214,N_2548);
or U8661 (N_8661,N_1189,N_4650);
or U8662 (N_8662,N_3937,N_2241);
and U8663 (N_8663,N_4340,N_1797);
nand U8664 (N_8664,N_1546,N_1650);
or U8665 (N_8665,N_4255,N_4119);
nand U8666 (N_8666,N_1797,N_2962);
nor U8667 (N_8667,N_3844,N_1104);
xor U8668 (N_8668,N_4620,N_3843);
xor U8669 (N_8669,N_3339,N_1676);
xnor U8670 (N_8670,N_4276,N_983);
xnor U8671 (N_8671,N_2294,N_4231);
and U8672 (N_8672,N_3922,N_4948);
nor U8673 (N_8673,N_3412,N_2203);
nor U8674 (N_8674,N_1226,N_3093);
nand U8675 (N_8675,N_3239,N_2950);
nor U8676 (N_8676,N_3011,N_3753);
xor U8677 (N_8677,N_1813,N_3230);
nor U8678 (N_8678,N_3380,N_4235);
xor U8679 (N_8679,N_3162,N_4291);
nor U8680 (N_8680,N_4041,N_2082);
or U8681 (N_8681,N_2474,N_2626);
xnor U8682 (N_8682,N_3294,N_3338);
and U8683 (N_8683,N_1917,N_4851);
nor U8684 (N_8684,N_4789,N_529);
nor U8685 (N_8685,N_4638,N_3769);
nand U8686 (N_8686,N_3872,N_2045);
and U8687 (N_8687,N_3349,N_2163);
nor U8688 (N_8688,N_640,N_485);
nor U8689 (N_8689,N_2677,N_3852);
or U8690 (N_8690,N_1608,N_2849);
xor U8691 (N_8691,N_2580,N_1580);
and U8692 (N_8692,N_2357,N_281);
and U8693 (N_8693,N_2617,N_2465);
nand U8694 (N_8694,N_2978,N_3223);
nand U8695 (N_8695,N_338,N_3233);
and U8696 (N_8696,N_2224,N_3015);
or U8697 (N_8697,N_1265,N_1911);
nor U8698 (N_8698,N_962,N_2248);
nand U8699 (N_8699,N_3284,N_419);
nand U8700 (N_8700,N_1224,N_2996);
and U8701 (N_8701,N_1332,N_3123);
nand U8702 (N_8702,N_3862,N_2816);
nor U8703 (N_8703,N_2639,N_922);
nor U8704 (N_8704,N_4323,N_3430);
and U8705 (N_8705,N_4399,N_896);
nor U8706 (N_8706,N_2728,N_3348);
nor U8707 (N_8707,N_1041,N_1573);
nand U8708 (N_8708,N_1470,N_3996);
or U8709 (N_8709,N_2739,N_1883);
or U8710 (N_8710,N_622,N_485);
xor U8711 (N_8711,N_2623,N_573);
or U8712 (N_8712,N_254,N_1388);
xor U8713 (N_8713,N_972,N_302);
xor U8714 (N_8714,N_4204,N_3173);
and U8715 (N_8715,N_2017,N_2762);
and U8716 (N_8716,N_3509,N_1821);
nand U8717 (N_8717,N_1736,N_3904);
xor U8718 (N_8718,N_4759,N_1440);
nand U8719 (N_8719,N_4350,N_2177);
xnor U8720 (N_8720,N_2012,N_1829);
xor U8721 (N_8721,N_2330,N_3686);
or U8722 (N_8722,N_3600,N_3772);
or U8723 (N_8723,N_1831,N_3630);
and U8724 (N_8724,N_4563,N_4850);
and U8725 (N_8725,N_1816,N_4310);
nor U8726 (N_8726,N_480,N_333);
and U8727 (N_8727,N_1765,N_4165);
or U8728 (N_8728,N_3291,N_4050);
nand U8729 (N_8729,N_456,N_2517);
nor U8730 (N_8730,N_1275,N_922);
xor U8731 (N_8731,N_3116,N_2330);
nand U8732 (N_8732,N_1456,N_3116);
nor U8733 (N_8733,N_342,N_4685);
or U8734 (N_8734,N_3128,N_4043);
nand U8735 (N_8735,N_4124,N_2792);
or U8736 (N_8736,N_2127,N_2481);
and U8737 (N_8737,N_803,N_4726);
xnor U8738 (N_8738,N_834,N_1696);
and U8739 (N_8739,N_1524,N_2308);
and U8740 (N_8740,N_3498,N_3828);
or U8741 (N_8741,N_3537,N_2579);
xnor U8742 (N_8742,N_1258,N_4300);
xnor U8743 (N_8743,N_1436,N_2667);
or U8744 (N_8744,N_2417,N_1552);
and U8745 (N_8745,N_4235,N_775);
xor U8746 (N_8746,N_1609,N_479);
and U8747 (N_8747,N_2154,N_1665);
xor U8748 (N_8748,N_4876,N_4323);
nand U8749 (N_8749,N_3845,N_2072);
or U8750 (N_8750,N_2049,N_1777);
nand U8751 (N_8751,N_2244,N_3565);
xnor U8752 (N_8752,N_1785,N_1932);
nor U8753 (N_8753,N_4464,N_4086);
nor U8754 (N_8754,N_3315,N_3394);
nor U8755 (N_8755,N_2403,N_2284);
nor U8756 (N_8756,N_187,N_2888);
and U8757 (N_8757,N_305,N_3325);
nand U8758 (N_8758,N_2140,N_2245);
nand U8759 (N_8759,N_1972,N_598);
nor U8760 (N_8760,N_1382,N_1232);
nor U8761 (N_8761,N_116,N_1604);
xor U8762 (N_8762,N_1246,N_3791);
and U8763 (N_8763,N_1609,N_1608);
or U8764 (N_8764,N_97,N_3890);
xnor U8765 (N_8765,N_2909,N_613);
and U8766 (N_8766,N_3877,N_2128);
or U8767 (N_8767,N_1185,N_3922);
and U8768 (N_8768,N_3711,N_3008);
nand U8769 (N_8769,N_1879,N_4239);
nor U8770 (N_8770,N_70,N_1117);
xnor U8771 (N_8771,N_1684,N_2070);
nand U8772 (N_8772,N_4837,N_95);
and U8773 (N_8773,N_4136,N_641);
nor U8774 (N_8774,N_3490,N_2998);
xnor U8775 (N_8775,N_452,N_611);
xnor U8776 (N_8776,N_270,N_3768);
or U8777 (N_8777,N_1002,N_4932);
and U8778 (N_8778,N_4966,N_925);
nor U8779 (N_8779,N_1250,N_240);
or U8780 (N_8780,N_4502,N_3566);
nand U8781 (N_8781,N_2063,N_4469);
nand U8782 (N_8782,N_2678,N_2670);
nor U8783 (N_8783,N_3971,N_1402);
and U8784 (N_8784,N_587,N_1020);
nand U8785 (N_8785,N_3117,N_4724);
and U8786 (N_8786,N_1797,N_1200);
xor U8787 (N_8787,N_3464,N_1312);
xor U8788 (N_8788,N_2781,N_2141);
nand U8789 (N_8789,N_893,N_2638);
nand U8790 (N_8790,N_2155,N_4035);
nand U8791 (N_8791,N_4993,N_3131);
nor U8792 (N_8792,N_292,N_48);
xnor U8793 (N_8793,N_1059,N_86);
xor U8794 (N_8794,N_597,N_768);
and U8795 (N_8795,N_2187,N_808);
and U8796 (N_8796,N_4245,N_1584);
nor U8797 (N_8797,N_1396,N_2877);
or U8798 (N_8798,N_2008,N_571);
or U8799 (N_8799,N_4966,N_795);
and U8800 (N_8800,N_273,N_581);
nor U8801 (N_8801,N_694,N_984);
and U8802 (N_8802,N_1719,N_583);
and U8803 (N_8803,N_652,N_538);
and U8804 (N_8804,N_2122,N_4544);
nor U8805 (N_8805,N_4555,N_182);
nor U8806 (N_8806,N_2120,N_917);
or U8807 (N_8807,N_3237,N_3699);
nor U8808 (N_8808,N_3287,N_4237);
xnor U8809 (N_8809,N_3236,N_4268);
nand U8810 (N_8810,N_1378,N_1201);
nor U8811 (N_8811,N_1348,N_3493);
or U8812 (N_8812,N_53,N_1959);
nand U8813 (N_8813,N_2453,N_3861);
nor U8814 (N_8814,N_2381,N_4187);
or U8815 (N_8815,N_838,N_1366);
and U8816 (N_8816,N_77,N_307);
nor U8817 (N_8817,N_1359,N_316);
xnor U8818 (N_8818,N_943,N_319);
or U8819 (N_8819,N_2528,N_2010);
and U8820 (N_8820,N_4406,N_814);
nand U8821 (N_8821,N_3415,N_2489);
nor U8822 (N_8822,N_3826,N_2369);
and U8823 (N_8823,N_3909,N_2463);
or U8824 (N_8824,N_1581,N_4389);
or U8825 (N_8825,N_2962,N_235);
nand U8826 (N_8826,N_1065,N_2371);
nor U8827 (N_8827,N_3063,N_2536);
or U8828 (N_8828,N_4932,N_3511);
nand U8829 (N_8829,N_1725,N_1626);
nand U8830 (N_8830,N_2798,N_3017);
nor U8831 (N_8831,N_1050,N_1125);
xnor U8832 (N_8832,N_1648,N_4698);
or U8833 (N_8833,N_2748,N_4095);
or U8834 (N_8834,N_2225,N_2018);
nor U8835 (N_8835,N_2582,N_390);
and U8836 (N_8836,N_2930,N_2457);
nand U8837 (N_8837,N_4401,N_996);
or U8838 (N_8838,N_2233,N_4733);
xor U8839 (N_8839,N_2799,N_652);
xor U8840 (N_8840,N_4159,N_3735);
and U8841 (N_8841,N_4349,N_2998);
and U8842 (N_8842,N_3770,N_4955);
or U8843 (N_8843,N_4749,N_3458);
nand U8844 (N_8844,N_1069,N_4795);
or U8845 (N_8845,N_3131,N_4773);
xor U8846 (N_8846,N_1735,N_2302);
xor U8847 (N_8847,N_4921,N_1919);
nand U8848 (N_8848,N_1313,N_2262);
nand U8849 (N_8849,N_477,N_921);
xnor U8850 (N_8850,N_3648,N_3676);
nor U8851 (N_8851,N_983,N_1667);
nand U8852 (N_8852,N_1852,N_1589);
and U8853 (N_8853,N_3338,N_2234);
xor U8854 (N_8854,N_1227,N_3215);
nor U8855 (N_8855,N_1690,N_4840);
xnor U8856 (N_8856,N_4850,N_4441);
nor U8857 (N_8857,N_1070,N_4484);
nor U8858 (N_8858,N_2538,N_857);
and U8859 (N_8859,N_4881,N_1936);
nand U8860 (N_8860,N_649,N_4490);
xor U8861 (N_8861,N_2641,N_596);
and U8862 (N_8862,N_4257,N_3258);
and U8863 (N_8863,N_2721,N_913);
and U8864 (N_8864,N_1525,N_457);
or U8865 (N_8865,N_1542,N_950);
xnor U8866 (N_8866,N_3374,N_247);
nand U8867 (N_8867,N_2269,N_4811);
nand U8868 (N_8868,N_854,N_4847);
xnor U8869 (N_8869,N_3362,N_1060);
and U8870 (N_8870,N_2642,N_4813);
nor U8871 (N_8871,N_105,N_394);
and U8872 (N_8872,N_3018,N_1678);
nor U8873 (N_8873,N_3096,N_2208);
nor U8874 (N_8874,N_3843,N_3378);
nand U8875 (N_8875,N_2718,N_3685);
and U8876 (N_8876,N_2728,N_726);
nor U8877 (N_8877,N_1621,N_2180);
and U8878 (N_8878,N_3365,N_1460);
nand U8879 (N_8879,N_641,N_2629);
nand U8880 (N_8880,N_2693,N_4193);
and U8881 (N_8881,N_399,N_2712);
xnor U8882 (N_8882,N_1163,N_3252);
xor U8883 (N_8883,N_3431,N_4111);
or U8884 (N_8884,N_2440,N_3727);
and U8885 (N_8885,N_341,N_1772);
nand U8886 (N_8886,N_2378,N_4476);
and U8887 (N_8887,N_3356,N_3732);
and U8888 (N_8888,N_43,N_253);
nand U8889 (N_8889,N_4458,N_1079);
nor U8890 (N_8890,N_2229,N_2123);
or U8891 (N_8891,N_3066,N_3567);
xor U8892 (N_8892,N_4459,N_1843);
nand U8893 (N_8893,N_3632,N_4434);
or U8894 (N_8894,N_2987,N_2599);
xor U8895 (N_8895,N_834,N_2994);
xnor U8896 (N_8896,N_2272,N_2125);
and U8897 (N_8897,N_2827,N_3733);
nor U8898 (N_8898,N_4964,N_3703);
nor U8899 (N_8899,N_1962,N_3581);
and U8900 (N_8900,N_4032,N_3172);
nor U8901 (N_8901,N_2435,N_1252);
or U8902 (N_8902,N_1042,N_4620);
and U8903 (N_8903,N_1635,N_4475);
xnor U8904 (N_8904,N_3299,N_277);
xor U8905 (N_8905,N_1746,N_411);
xnor U8906 (N_8906,N_4996,N_4054);
or U8907 (N_8907,N_4823,N_2164);
or U8908 (N_8908,N_2860,N_3020);
xnor U8909 (N_8909,N_1373,N_4462);
nand U8910 (N_8910,N_2840,N_4377);
or U8911 (N_8911,N_4423,N_2137);
and U8912 (N_8912,N_1478,N_3826);
or U8913 (N_8913,N_3943,N_3374);
nor U8914 (N_8914,N_2603,N_142);
nand U8915 (N_8915,N_980,N_330);
nand U8916 (N_8916,N_2528,N_4700);
or U8917 (N_8917,N_2772,N_329);
nand U8918 (N_8918,N_414,N_1958);
and U8919 (N_8919,N_4171,N_1962);
nand U8920 (N_8920,N_3015,N_2638);
xnor U8921 (N_8921,N_1642,N_768);
and U8922 (N_8922,N_4252,N_3800);
nor U8923 (N_8923,N_4140,N_1679);
nor U8924 (N_8924,N_4125,N_2517);
nand U8925 (N_8925,N_2620,N_4110);
xor U8926 (N_8926,N_3620,N_3253);
xnor U8927 (N_8927,N_1367,N_1404);
or U8928 (N_8928,N_753,N_2751);
xnor U8929 (N_8929,N_3510,N_2593);
or U8930 (N_8930,N_1131,N_4318);
xnor U8931 (N_8931,N_340,N_3610);
nand U8932 (N_8932,N_3588,N_1696);
and U8933 (N_8933,N_1549,N_2241);
xor U8934 (N_8934,N_1094,N_1485);
xor U8935 (N_8935,N_196,N_3591);
nor U8936 (N_8936,N_3500,N_927);
or U8937 (N_8937,N_2239,N_883);
nand U8938 (N_8938,N_3336,N_3016);
nand U8939 (N_8939,N_1498,N_1127);
xnor U8940 (N_8940,N_1071,N_2640);
xnor U8941 (N_8941,N_515,N_2217);
and U8942 (N_8942,N_4633,N_1285);
and U8943 (N_8943,N_586,N_590);
xnor U8944 (N_8944,N_3426,N_1489);
nor U8945 (N_8945,N_1958,N_2779);
nor U8946 (N_8946,N_1414,N_3844);
nor U8947 (N_8947,N_4461,N_3029);
xor U8948 (N_8948,N_3685,N_4528);
nor U8949 (N_8949,N_2632,N_1392);
or U8950 (N_8950,N_1087,N_2364);
nor U8951 (N_8951,N_889,N_3862);
or U8952 (N_8952,N_4429,N_3762);
xnor U8953 (N_8953,N_4429,N_2715);
xnor U8954 (N_8954,N_1398,N_2060);
or U8955 (N_8955,N_3668,N_2638);
or U8956 (N_8956,N_4863,N_4867);
xnor U8957 (N_8957,N_780,N_3858);
and U8958 (N_8958,N_4603,N_2714);
xnor U8959 (N_8959,N_382,N_1953);
or U8960 (N_8960,N_4561,N_59);
nor U8961 (N_8961,N_2425,N_1675);
nor U8962 (N_8962,N_3762,N_146);
nor U8963 (N_8963,N_1477,N_4910);
and U8964 (N_8964,N_2191,N_2124);
or U8965 (N_8965,N_4463,N_3194);
and U8966 (N_8966,N_1967,N_247);
nand U8967 (N_8967,N_4109,N_4153);
and U8968 (N_8968,N_83,N_3135);
or U8969 (N_8969,N_2903,N_2740);
xor U8970 (N_8970,N_4410,N_4605);
nor U8971 (N_8971,N_3644,N_2504);
xor U8972 (N_8972,N_404,N_335);
xor U8973 (N_8973,N_4178,N_3320);
nand U8974 (N_8974,N_2776,N_4022);
and U8975 (N_8975,N_3785,N_1320);
nand U8976 (N_8976,N_3195,N_4591);
nand U8977 (N_8977,N_3693,N_1035);
and U8978 (N_8978,N_3787,N_400);
xor U8979 (N_8979,N_1044,N_3798);
nand U8980 (N_8980,N_4169,N_2270);
and U8981 (N_8981,N_6,N_4090);
or U8982 (N_8982,N_4525,N_2598);
and U8983 (N_8983,N_50,N_149);
xor U8984 (N_8984,N_2733,N_3451);
nor U8985 (N_8985,N_1669,N_134);
xnor U8986 (N_8986,N_494,N_1490);
and U8987 (N_8987,N_644,N_2997);
and U8988 (N_8988,N_1819,N_897);
or U8989 (N_8989,N_4407,N_840);
nand U8990 (N_8990,N_3570,N_562);
nand U8991 (N_8991,N_1937,N_3725);
nor U8992 (N_8992,N_2534,N_1867);
xnor U8993 (N_8993,N_3863,N_1697);
nor U8994 (N_8994,N_2360,N_3440);
nand U8995 (N_8995,N_2818,N_3643);
and U8996 (N_8996,N_3562,N_3698);
nor U8997 (N_8997,N_1273,N_3632);
or U8998 (N_8998,N_4796,N_841);
or U8999 (N_8999,N_2375,N_3053);
or U9000 (N_9000,N_3602,N_1117);
nor U9001 (N_9001,N_747,N_4573);
nor U9002 (N_9002,N_1282,N_4378);
and U9003 (N_9003,N_4761,N_3830);
nor U9004 (N_9004,N_2753,N_10);
and U9005 (N_9005,N_2557,N_646);
and U9006 (N_9006,N_4779,N_745);
nand U9007 (N_9007,N_2144,N_4649);
nand U9008 (N_9008,N_2008,N_3043);
and U9009 (N_9009,N_2909,N_125);
nor U9010 (N_9010,N_4216,N_4283);
or U9011 (N_9011,N_2772,N_1335);
or U9012 (N_9012,N_128,N_3471);
nand U9013 (N_9013,N_1921,N_3290);
nor U9014 (N_9014,N_1929,N_4576);
nand U9015 (N_9015,N_2242,N_2773);
xnor U9016 (N_9016,N_345,N_4681);
xor U9017 (N_9017,N_43,N_869);
and U9018 (N_9018,N_2212,N_1350);
nor U9019 (N_9019,N_4697,N_1447);
xor U9020 (N_9020,N_2064,N_2058);
xor U9021 (N_9021,N_1438,N_4849);
and U9022 (N_9022,N_2439,N_3884);
nor U9023 (N_9023,N_295,N_3086);
xnor U9024 (N_9024,N_3438,N_3595);
or U9025 (N_9025,N_3418,N_1070);
and U9026 (N_9026,N_3391,N_1611);
nand U9027 (N_9027,N_1221,N_4248);
nor U9028 (N_9028,N_1675,N_765);
and U9029 (N_9029,N_1768,N_756);
xnor U9030 (N_9030,N_2086,N_4797);
or U9031 (N_9031,N_3935,N_7);
or U9032 (N_9032,N_2012,N_2208);
nor U9033 (N_9033,N_2473,N_2322);
and U9034 (N_9034,N_4696,N_641);
nor U9035 (N_9035,N_4832,N_1194);
xor U9036 (N_9036,N_2386,N_2900);
or U9037 (N_9037,N_101,N_3128);
xor U9038 (N_9038,N_4362,N_2252);
xor U9039 (N_9039,N_2595,N_1635);
nor U9040 (N_9040,N_2826,N_1643);
or U9041 (N_9041,N_3243,N_72);
xor U9042 (N_9042,N_3511,N_4876);
and U9043 (N_9043,N_333,N_4195);
or U9044 (N_9044,N_3277,N_3567);
xnor U9045 (N_9045,N_3277,N_1570);
or U9046 (N_9046,N_3092,N_47);
xor U9047 (N_9047,N_3028,N_1058);
nor U9048 (N_9048,N_3449,N_1791);
xnor U9049 (N_9049,N_1278,N_3882);
nand U9050 (N_9050,N_1926,N_595);
nand U9051 (N_9051,N_1431,N_4998);
and U9052 (N_9052,N_3832,N_4061);
nor U9053 (N_9053,N_2702,N_2994);
nor U9054 (N_9054,N_4711,N_540);
nand U9055 (N_9055,N_2209,N_43);
nor U9056 (N_9056,N_1070,N_380);
xnor U9057 (N_9057,N_1448,N_2725);
xor U9058 (N_9058,N_2597,N_1465);
or U9059 (N_9059,N_1628,N_2920);
xor U9060 (N_9060,N_4835,N_1790);
xor U9061 (N_9061,N_2139,N_2706);
and U9062 (N_9062,N_1251,N_1564);
or U9063 (N_9063,N_1344,N_4348);
nand U9064 (N_9064,N_1921,N_3246);
and U9065 (N_9065,N_730,N_1256);
xor U9066 (N_9066,N_4619,N_2151);
and U9067 (N_9067,N_3414,N_2791);
and U9068 (N_9068,N_3213,N_3578);
xnor U9069 (N_9069,N_2035,N_359);
and U9070 (N_9070,N_2734,N_147);
nor U9071 (N_9071,N_2982,N_2004);
xnor U9072 (N_9072,N_573,N_4171);
or U9073 (N_9073,N_1786,N_3980);
nand U9074 (N_9074,N_2009,N_1911);
nor U9075 (N_9075,N_3271,N_83);
nor U9076 (N_9076,N_3392,N_2848);
xnor U9077 (N_9077,N_2284,N_4865);
or U9078 (N_9078,N_2838,N_2065);
and U9079 (N_9079,N_4110,N_3879);
xnor U9080 (N_9080,N_970,N_3278);
and U9081 (N_9081,N_974,N_1091);
xor U9082 (N_9082,N_923,N_4369);
xnor U9083 (N_9083,N_1792,N_3184);
or U9084 (N_9084,N_797,N_4182);
nand U9085 (N_9085,N_1274,N_3742);
xor U9086 (N_9086,N_3344,N_4755);
nor U9087 (N_9087,N_3533,N_2330);
or U9088 (N_9088,N_3049,N_1867);
nor U9089 (N_9089,N_4147,N_265);
or U9090 (N_9090,N_2333,N_1901);
nand U9091 (N_9091,N_2515,N_4917);
and U9092 (N_9092,N_4656,N_3434);
or U9093 (N_9093,N_2161,N_4666);
nand U9094 (N_9094,N_4732,N_433);
nand U9095 (N_9095,N_530,N_2683);
nor U9096 (N_9096,N_183,N_1810);
nand U9097 (N_9097,N_4423,N_3777);
xor U9098 (N_9098,N_3140,N_4985);
xor U9099 (N_9099,N_3130,N_377);
nand U9100 (N_9100,N_4012,N_4754);
nor U9101 (N_9101,N_3644,N_1483);
xor U9102 (N_9102,N_1394,N_1003);
or U9103 (N_9103,N_490,N_533);
nor U9104 (N_9104,N_293,N_1874);
nand U9105 (N_9105,N_1616,N_4951);
or U9106 (N_9106,N_3408,N_2206);
xnor U9107 (N_9107,N_104,N_3082);
or U9108 (N_9108,N_2084,N_1330);
nand U9109 (N_9109,N_3126,N_3453);
and U9110 (N_9110,N_810,N_3408);
nand U9111 (N_9111,N_3815,N_1756);
nand U9112 (N_9112,N_2217,N_4221);
or U9113 (N_9113,N_3309,N_2842);
nand U9114 (N_9114,N_3631,N_2274);
and U9115 (N_9115,N_3527,N_3263);
and U9116 (N_9116,N_3449,N_840);
and U9117 (N_9117,N_2824,N_3500);
nand U9118 (N_9118,N_3108,N_4560);
or U9119 (N_9119,N_3198,N_2186);
and U9120 (N_9120,N_2082,N_2605);
or U9121 (N_9121,N_4990,N_3184);
and U9122 (N_9122,N_608,N_4781);
nor U9123 (N_9123,N_4122,N_3691);
xnor U9124 (N_9124,N_4188,N_2938);
or U9125 (N_9125,N_4860,N_3414);
nor U9126 (N_9126,N_4475,N_3369);
xnor U9127 (N_9127,N_427,N_107);
nor U9128 (N_9128,N_3437,N_1145);
and U9129 (N_9129,N_869,N_2876);
xor U9130 (N_9130,N_924,N_4738);
and U9131 (N_9131,N_4690,N_441);
xnor U9132 (N_9132,N_1519,N_1601);
nand U9133 (N_9133,N_4833,N_3860);
nor U9134 (N_9134,N_240,N_4381);
xnor U9135 (N_9135,N_132,N_542);
xnor U9136 (N_9136,N_19,N_241);
nand U9137 (N_9137,N_2201,N_1935);
nand U9138 (N_9138,N_2816,N_3013);
nor U9139 (N_9139,N_2176,N_3929);
nand U9140 (N_9140,N_4073,N_2798);
or U9141 (N_9141,N_4858,N_4697);
nand U9142 (N_9142,N_1821,N_1311);
and U9143 (N_9143,N_1360,N_3465);
nor U9144 (N_9144,N_4852,N_338);
nand U9145 (N_9145,N_4367,N_4275);
nand U9146 (N_9146,N_1191,N_2458);
nor U9147 (N_9147,N_2367,N_4333);
and U9148 (N_9148,N_2906,N_3040);
or U9149 (N_9149,N_765,N_3729);
xnor U9150 (N_9150,N_1289,N_4376);
nand U9151 (N_9151,N_267,N_795);
nor U9152 (N_9152,N_1005,N_1143);
nor U9153 (N_9153,N_1482,N_4941);
xor U9154 (N_9154,N_2829,N_4988);
and U9155 (N_9155,N_2757,N_2933);
xnor U9156 (N_9156,N_221,N_4316);
or U9157 (N_9157,N_2172,N_2672);
nand U9158 (N_9158,N_4786,N_3320);
xnor U9159 (N_9159,N_1911,N_4015);
nor U9160 (N_9160,N_1428,N_4474);
or U9161 (N_9161,N_2720,N_2548);
xnor U9162 (N_9162,N_185,N_2729);
xor U9163 (N_9163,N_1011,N_2552);
nor U9164 (N_9164,N_915,N_1079);
or U9165 (N_9165,N_1052,N_2772);
nand U9166 (N_9166,N_1873,N_827);
nand U9167 (N_9167,N_3224,N_2866);
nor U9168 (N_9168,N_4691,N_4255);
nand U9169 (N_9169,N_1670,N_4593);
xnor U9170 (N_9170,N_2876,N_378);
or U9171 (N_9171,N_3123,N_433);
nand U9172 (N_9172,N_3169,N_4484);
nand U9173 (N_9173,N_147,N_4189);
or U9174 (N_9174,N_611,N_37);
nand U9175 (N_9175,N_1471,N_594);
nor U9176 (N_9176,N_2124,N_712);
and U9177 (N_9177,N_982,N_2486);
or U9178 (N_9178,N_1531,N_554);
xnor U9179 (N_9179,N_3779,N_947);
xor U9180 (N_9180,N_1899,N_941);
nor U9181 (N_9181,N_2682,N_4616);
or U9182 (N_9182,N_4487,N_2563);
nor U9183 (N_9183,N_2110,N_4093);
or U9184 (N_9184,N_275,N_3567);
nor U9185 (N_9185,N_1533,N_2711);
nor U9186 (N_9186,N_814,N_3344);
or U9187 (N_9187,N_2903,N_277);
xor U9188 (N_9188,N_3500,N_999);
or U9189 (N_9189,N_3599,N_4349);
xnor U9190 (N_9190,N_2592,N_632);
nor U9191 (N_9191,N_3478,N_1272);
or U9192 (N_9192,N_3403,N_2701);
xnor U9193 (N_9193,N_4053,N_585);
xor U9194 (N_9194,N_2930,N_593);
xor U9195 (N_9195,N_4121,N_1749);
xnor U9196 (N_9196,N_641,N_3345);
and U9197 (N_9197,N_4809,N_3534);
nor U9198 (N_9198,N_4890,N_2404);
xor U9199 (N_9199,N_3328,N_4921);
nand U9200 (N_9200,N_3241,N_2732);
nor U9201 (N_9201,N_1997,N_689);
and U9202 (N_9202,N_4639,N_266);
nor U9203 (N_9203,N_4796,N_4734);
or U9204 (N_9204,N_4910,N_4590);
or U9205 (N_9205,N_1343,N_4354);
nor U9206 (N_9206,N_4765,N_2377);
or U9207 (N_9207,N_1254,N_3729);
and U9208 (N_9208,N_2199,N_801);
and U9209 (N_9209,N_4845,N_4260);
or U9210 (N_9210,N_3960,N_2109);
and U9211 (N_9211,N_2525,N_2482);
xnor U9212 (N_9212,N_215,N_1226);
nand U9213 (N_9213,N_2970,N_575);
xor U9214 (N_9214,N_2164,N_4296);
and U9215 (N_9215,N_1691,N_2919);
xnor U9216 (N_9216,N_2799,N_3654);
nor U9217 (N_9217,N_461,N_54);
nor U9218 (N_9218,N_1675,N_4259);
nand U9219 (N_9219,N_4275,N_1298);
nor U9220 (N_9220,N_60,N_4289);
or U9221 (N_9221,N_882,N_1306);
and U9222 (N_9222,N_2662,N_2489);
nand U9223 (N_9223,N_1364,N_103);
nand U9224 (N_9224,N_4231,N_3657);
or U9225 (N_9225,N_2777,N_3021);
and U9226 (N_9226,N_3101,N_1265);
nand U9227 (N_9227,N_1454,N_1156);
nor U9228 (N_9228,N_3053,N_4182);
nor U9229 (N_9229,N_2650,N_3659);
or U9230 (N_9230,N_110,N_1314);
and U9231 (N_9231,N_920,N_2633);
or U9232 (N_9232,N_1415,N_3744);
xnor U9233 (N_9233,N_3839,N_3478);
or U9234 (N_9234,N_2123,N_28);
and U9235 (N_9235,N_4381,N_1858);
and U9236 (N_9236,N_1141,N_1266);
nand U9237 (N_9237,N_3751,N_3323);
or U9238 (N_9238,N_2344,N_4222);
and U9239 (N_9239,N_1663,N_2380);
nand U9240 (N_9240,N_2511,N_2436);
nor U9241 (N_9241,N_3574,N_891);
nor U9242 (N_9242,N_500,N_1755);
nor U9243 (N_9243,N_2965,N_3504);
nand U9244 (N_9244,N_4883,N_1914);
xnor U9245 (N_9245,N_2820,N_2925);
nor U9246 (N_9246,N_3681,N_3793);
xnor U9247 (N_9247,N_4048,N_1405);
nand U9248 (N_9248,N_3789,N_2321);
or U9249 (N_9249,N_1573,N_306);
or U9250 (N_9250,N_3452,N_3593);
and U9251 (N_9251,N_4361,N_1171);
xnor U9252 (N_9252,N_4901,N_3742);
or U9253 (N_9253,N_3667,N_4700);
or U9254 (N_9254,N_4314,N_2514);
or U9255 (N_9255,N_2394,N_3409);
and U9256 (N_9256,N_1159,N_4182);
or U9257 (N_9257,N_4206,N_653);
nand U9258 (N_9258,N_146,N_239);
and U9259 (N_9259,N_1336,N_344);
nand U9260 (N_9260,N_3419,N_170);
nand U9261 (N_9261,N_1876,N_2073);
and U9262 (N_9262,N_3785,N_1620);
or U9263 (N_9263,N_2234,N_542);
xnor U9264 (N_9264,N_1359,N_3224);
xor U9265 (N_9265,N_1496,N_222);
nor U9266 (N_9266,N_279,N_2583);
and U9267 (N_9267,N_876,N_2866);
xor U9268 (N_9268,N_4129,N_62);
nor U9269 (N_9269,N_409,N_2151);
xor U9270 (N_9270,N_1968,N_1774);
xnor U9271 (N_9271,N_3987,N_3345);
nand U9272 (N_9272,N_587,N_3831);
nand U9273 (N_9273,N_3198,N_2599);
xor U9274 (N_9274,N_404,N_3671);
and U9275 (N_9275,N_4325,N_1335);
and U9276 (N_9276,N_2868,N_116);
nor U9277 (N_9277,N_3432,N_4730);
nor U9278 (N_9278,N_3360,N_836);
nor U9279 (N_9279,N_4764,N_2197);
nand U9280 (N_9280,N_2083,N_3790);
nand U9281 (N_9281,N_3497,N_2732);
or U9282 (N_9282,N_3264,N_3560);
xor U9283 (N_9283,N_4203,N_4776);
or U9284 (N_9284,N_3797,N_2259);
xnor U9285 (N_9285,N_2339,N_2608);
nor U9286 (N_9286,N_3643,N_1089);
nor U9287 (N_9287,N_3122,N_3580);
or U9288 (N_9288,N_1878,N_1797);
or U9289 (N_9289,N_4671,N_4024);
and U9290 (N_9290,N_3266,N_2853);
or U9291 (N_9291,N_3482,N_1406);
nand U9292 (N_9292,N_312,N_1761);
and U9293 (N_9293,N_2562,N_3017);
xor U9294 (N_9294,N_1041,N_3749);
nor U9295 (N_9295,N_3437,N_999);
nor U9296 (N_9296,N_4612,N_1284);
nor U9297 (N_9297,N_1558,N_4910);
nor U9298 (N_9298,N_1107,N_4187);
xnor U9299 (N_9299,N_1580,N_1614);
nand U9300 (N_9300,N_47,N_2972);
nor U9301 (N_9301,N_3355,N_1358);
xnor U9302 (N_9302,N_4013,N_1222);
or U9303 (N_9303,N_1870,N_663);
nor U9304 (N_9304,N_4259,N_4089);
or U9305 (N_9305,N_2336,N_311);
xor U9306 (N_9306,N_3964,N_174);
nand U9307 (N_9307,N_1521,N_1383);
or U9308 (N_9308,N_4446,N_2130);
nor U9309 (N_9309,N_4360,N_2677);
and U9310 (N_9310,N_902,N_3284);
nor U9311 (N_9311,N_4998,N_1176);
nor U9312 (N_9312,N_3486,N_4882);
and U9313 (N_9313,N_705,N_3541);
nor U9314 (N_9314,N_3707,N_822);
xor U9315 (N_9315,N_4070,N_3362);
xnor U9316 (N_9316,N_1337,N_143);
or U9317 (N_9317,N_2926,N_1822);
nand U9318 (N_9318,N_3269,N_818);
or U9319 (N_9319,N_4377,N_1165);
nor U9320 (N_9320,N_29,N_1071);
and U9321 (N_9321,N_284,N_4817);
and U9322 (N_9322,N_4074,N_1860);
or U9323 (N_9323,N_238,N_3032);
nand U9324 (N_9324,N_4217,N_2071);
nor U9325 (N_9325,N_1159,N_1879);
nand U9326 (N_9326,N_528,N_443);
or U9327 (N_9327,N_1446,N_1514);
and U9328 (N_9328,N_3417,N_2446);
nor U9329 (N_9329,N_1156,N_4760);
nor U9330 (N_9330,N_1059,N_2113);
nand U9331 (N_9331,N_3196,N_1349);
xor U9332 (N_9332,N_4053,N_2034);
nor U9333 (N_9333,N_3704,N_4291);
xor U9334 (N_9334,N_1245,N_2892);
or U9335 (N_9335,N_2605,N_4348);
xor U9336 (N_9336,N_3866,N_443);
nor U9337 (N_9337,N_1409,N_4552);
nor U9338 (N_9338,N_3034,N_4195);
nand U9339 (N_9339,N_2605,N_3854);
nand U9340 (N_9340,N_3136,N_3688);
or U9341 (N_9341,N_167,N_2269);
and U9342 (N_9342,N_4889,N_4343);
nor U9343 (N_9343,N_3243,N_29);
nand U9344 (N_9344,N_808,N_3728);
xnor U9345 (N_9345,N_3117,N_1071);
or U9346 (N_9346,N_3355,N_3139);
and U9347 (N_9347,N_1938,N_4164);
nand U9348 (N_9348,N_2659,N_4309);
or U9349 (N_9349,N_2183,N_2601);
nand U9350 (N_9350,N_4702,N_3352);
or U9351 (N_9351,N_1829,N_1571);
nor U9352 (N_9352,N_4537,N_3663);
or U9353 (N_9353,N_4321,N_4727);
xnor U9354 (N_9354,N_44,N_1033);
nor U9355 (N_9355,N_428,N_2195);
and U9356 (N_9356,N_4506,N_108);
and U9357 (N_9357,N_651,N_4310);
or U9358 (N_9358,N_3380,N_4493);
and U9359 (N_9359,N_4278,N_449);
nor U9360 (N_9360,N_2022,N_4152);
nor U9361 (N_9361,N_259,N_1126);
nand U9362 (N_9362,N_1142,N_4311);
xnor U9363 (N_9363,N_4642,N_2478);
nor U9364 (N_9364,N_1414,N_2873);
and U9365 (N_9365,N_4726,N_4238);
and U9366 (N_9366,N_1123,N_3489);
nor U9367 (N_9367,N_3663,N_1774);
nor U9368 (N_9368,N_1918,N_2731);
nor U9369 (N_9369,N_3697,N_4735);
and U9370 (N_9370,N_2798,N_1670);
nor U9371 (N_9371,N_3076,N_2067);
nand U9372 (N_9372,N_3812,N_2221);
or U9373 (N_9373,N_2327,N_3417);
nand U9374 (N_9374,N_1767,N_1533);
nand U9375 (N_9375,N_2104,N_300);
nand U9376 (N_9376,N_565,N_505);
and U9377 (N_9377,N_4719,N_1471);
xnor U9378 (N_9378,N_2007,N_2863);
and U9379 (N_9379,N_1041,N_4822);
nor U9380 (N_9380,N_205,N_2673);
nand U9381 (N_9381,N_4938,N_1719);
and U9382 (N_9382,N_4668,N_2147);
and U9383 (N_9383,N_841,N_3816);
or U9384 (N_9384,N_1006,N_4600);
and U9385 (N_9385,N_1845,N_3399);
or U9386 (N_9386,N_1915,N_4508);
nand U9387 (N_9387,N_1991,N_1697);
and U9388 (N_9388,N_2676,N_3244);
or U9389 (N_9389,N_3798,N_1917);
xnor U9390 (N_9390,N_3403,N_3432);
and U9391 (N_9391,N_1620,N_838);
and U9392 (N_9392,N_3359,N_4619);
and U9393 (N_9393,N_2464,N_3737);
nor U9394 (N_9394,N_2729,N_2588);
and U9395 (N_9395,N_4360,N_1598);
nor U9396 (N_9396,N_3975,N_4229);
xnor U9397 (N_9397,N_2929,N_4546);
nor U9398 (N_9398,N_67,N_2496);
xnor U9399 (N_9399,N_288,N_2914);
or U9400 (N_9400,N_2625,N_3524);
and U9401 (N_9401,N_1740,N_3778);
xnor U9402 (N_9402,N_4778,N_2200);
or U9403 (N_9403,N_1835,N_667);
and U9404 (N_9404,N_4350,N_4629);
nor U9405 (N_9405,N_922,N_409);
nor U9406 (N_9406,N_40,N_2088);
xor U9407 (N_9407,N_1199,N_3267);
and U9408 (N_9408,N_3240,N_1870);
or U9409 (N_9409,N_650,N_2811);
and U9410 (N_9410,N_3059,N_95);
nor U9411 (N_9411,N_207,N_4177);
nor U9412 (N_9412,N_3684,N_303);
xnor U9413 (N_9413,N_152,N_3128);
nor U9414 (N_9414,N_4933,N_1036);
and U9415 (N_9415,N_151,N_1001);
xnor U9416 (N_9416,N_71,N_646);
xor U9417 (N_9417,N_4175,N_4476);
nand U9418 (N_9418,N_893,N_1195);
and U9419 (N_9419,N_4626,N_928);
nand U9420 (N_9420,N_4550,N_2174);
nand U9421 (N_9421,N_4698,N_4482);
and U9422 (N_9422,N_109,N_4016);
nor U9423 (N_9423,N_324,N_295);
nor U9424 (N_9424,N_2260,N_3494);
nand U9425 (N_9425,N_4981,N_4266);
xor U9426 (N_9426,N_1097,N_752);
nor U9427 (N_9427,N_2961,N_2341);
xor U9428 (N_9428,N_1678,N_2170);
or U9429 (N_9429,N_4504,N_3873);
nand U9430 (N_9430,N_2164,N_1668);
and U9431 (N_9431,N_4680,N_72);
and U9432 (N_9432,N_4612,N_1484);
nor U9433 (N_9433,N_4746,N_22);
nand U9434 (N_9434,N_2753,N_3731);
or U9435 (N_9435,N_4033,N_4294);
or U9436 (N_9436,N_2970,N_356);
xor U9437 (N_9437,N_1136,N_4652);
or U9438 (N_9438,N_1290,N_845);
and U9439 (N_9439,N_3242,N_1911);
or U9440 (N_9440,N_1060,N_4152);
and U9441 (N_9441,N_4386,N_2074);
or U9442 (N_9442,N_3154,N_1111);
nand U9443 (N_9443,N_3210,N_2842);
nor U9444 (N_9444,N_1950,N_2073);
nand U9445 (N_9445,N_2528,N_2623);
nand U9446 (N_9446,N_475,N_3727);
xor U9447 (N_9447,N_1712,N_481);
or U9448 (N_9448,N_2986,N_3456);
and U9449 (N_9449,N_4078,N_3911);
or U9450 (N_9450,N_210,N_4054);
xor U9451 (N_9451,N_1522,N_2936);
or U9452 (N_9452,N_493,N_458);
xor U9453 (N_9453,N_4100,N_1280);
and U9454 (N_9454,N_3474,N_1238);
xor U9455 (N_9455,N_294,N_4103);
xnor U9456 (N_9456,N_2102,N_748);
nor U9457 (N_9457,N_985,N_79);
xnor U9458 (N_9458,N_2541,N_3357);
and U9459 (N_9459,N_4292,N_1794);
xnor U9460 (N_9460,N_1201,N_3581);
nand U9461 (N_9461,N_3663,N_2090);
and U9462 (N_9462,N_3196,N_2642);
or U9463 (N_9463,N_1466,N_2125);
or U9464 (N_9464,N_2763,N_4312);
nor U9465 (N_9465,N_2575,N_3508);
nor U9466 (N_9466,N_2911,N_1236);
nor U9467 (N_9467,N_2866,N_1784);
xnor U9468 (N_9468,N_2846,N_3592);
and U9469 (N_9469,N_1597,N_2924);
or U9470 (N_9470,N_1453,N_1917);
nand U9471 (N_9471,N_2165,N_2535);
nor U9472 (N_9472,N_3338,N_4432);
nand U9473 (N_9473,N_1869,N_976);
and U9474 (N_9474,N_208,N_2524);
xor U9475 (N_9475,N_1133,N_881);
nand U9476 (N_9476,N_3568,N_377);
and U9477 (N_9477,N_1431,N_16);
nand U9478 (N_9478,N_687,N_2299);
nor U9479 (N_9479,N_2092,N_517);
and U9480 (N_9480,N_1338,N_4877);
and U9481 (N_9481,N_4231,N_336);
and U9482 (N_9482,N_318,N_2763);
nor U9483 (N_9483,N_3278,N_2957);
nand U9484 (N_9484,N_4186,N_3183);
and U9485 (N_9485,N_2929,N_1579);
or U9486 (N_9486,N_2327,N_492);
nor U9487 (N_9487,N_1827,N_286);
nor U9488 (N_9488,N_2276,N_3785);
xor U9489 (N_9489,N_2237,N_502);
or U9490 (N_9490,N_2417,N_3214);
and U9491 (N_9491,N_4506,N_3057);
nor U9492 (N_9492,N_4395,N_3118);
xnor U9493 (N_9493,N_4028,N_1971);
nand U9494 (N_9494,N_4509,N_3408);
xnor U9495 (N_9495,N_4725,N_976);
nor U9496 (N_9496,N_1777,N_2706);
nand U9497 (N_9497,N_4832,N_1541);
or U9498 (N_9498,N_367,N_2086);
nor U9499 (N_9499,N_3073,N_3730);
and U9500 (N_9500,N_4235,N_3365);
or U9501 (N_9501,N_1147,N_3297);
nor U9502 (N_9502,N_1127,N_2711);
nand U9503 (N_9503,N_3101,N_4953);
or U9504 (N_9504,N_4520,N_2889);
nand U9505 (N_9505,N_3723,N_1879);
xor U9506 (N_9506,N_3868,N_4206);
nor U9507 (N_9507,N_39,N_3925);
or U9508 (N_9508,N_2206,N_2282);
xnor U9509 (N_9509,N_2935,N_3548);
nand U9510 (N_9510,N_713,N_3399);
nand U9511 (N_9511,N_4419,N_1279);
nand U9512 (N_9512,N_2996,N_696);
xnor U9513 (N_9513,N_3055,N_3711);
nand U9514 (N_9514,N_1590,N_4705);
xor U9515 (N_9515,N_2864,N_4828);
xnor U9516 (N_9516,N_4471,N_3179);
xnor U9517 (N_9517,N_4456,N_183);
nand U9518 (N_9518,N_3454,N_1801);
nand U9519 (N_9519,N_752,N_943);
nand U9520 (N_9520,N_4343,N_472);
and U9521 (N_9521,N_9,N_769);
xnor U9522 (N_9522,N_800,N_3087);
xnor U9523 (N_9523,N_4101,N_2478);
xor U9524 (N_9524,N_2451,N_428);
xor U9525 (N_9525,N_3311,N_377);
or U9526 (N_9526,N_191,N_2419);
nand U9527 (N_9527,N_2912,N_4527);
nor U9528 (N_9528,N_286,N_1355);
nand U9529 (N_9529,N_2920,N_3169);
or U9530 (N_9530,N_4534,N_4913);
xor U9531 (N_9531,N_3357,N_4072);
nor U9532 (N_9532,N_184,N_2597);
nand U9533 (N_9533,N_2444,N_3451);
nor U9534 (N_9534,N_2387,N_3400);
nand U9535 (N_9535,N_1780,N_3037);
nor U9536 (N_9536,N_1655,N_4778);
and U9537 (N_9537,N_675,N_2048);
xnor U9538 (N_9538,N_720,N_2947);
and U9539 (N_9539,N_2151,N_2403);
or U9540 (N_9540,N_3365,N_1680);
nand U9541 (N_9541,N_2467,N_4554);
xnor U9542 (N_9542,N_3846,N_40);
xor U9543 (N_9543,N_1439,N_1738);
nand U9544 (N_9544,N_2648,N_1418);
and U9545 (N_9545,N_4906,N_587);
nor U9546 (N_9546,N_915,N_116);
xnor U9547 (N_9547,N_861,N_3596);
xor U9548 (N_9548,N_4937,N_688);
and U9549 (N_9549,N_1755,N_1206);
or U9550 (N_9550,N_2129,N_2982);
or U9551 (N_9551,N_2368,N_3738);
and U9552 (N_9552,N_4795,N_284);
xnor U9553 (N_9553,N_3869,N_97);
nor U9554 (N_9554,N_3873,N_1128);
nor U9555 (N_9555,N_761,N_3394);
or U9556 (N_9556,N_2689,N_2998);
or U9557 (N_9557,N_393,N_3155);
and U9558 (N_9558,N_4996,N_3153);
xnor U9559 (N_9559,N_1898,N_2524);
nor U9560 (N_9560,N_2892,N_1183);
or U9561 (N_9561,N_2705,N_4025);
and U9562 (N_9562,N_2324,N_120);
or U9563 (N_9563,N_785,N_4059);
and U9564 (N_9564,N_4784,N_3950);
and U9565 (N_9565,N_2838,N_1868);
xnor U9566 (N_9566,N_1718,N_4063);
nand U9567 (N_9567,N_4407,N_2732);
nor U9568 (N_9568,N_3310,N_2407);
xor U9569 (N_9569,N_4936,N_1386);
nand U9570 (N_9570,N_275,N_4614);
nand U9571 (N_9571,N_2631,N_3273);
nor U9572 (N_9572,N_1710,N_821);
nor U9573 (N_9573,N_4777,N_1262);
nor U9574 (N_9574,N_594,N_2098);
nor U9575 (N_9575,N_4447,N_3807);
and U9576 (N_9576,N_1361,N_3193);
nand U9577 (N_9577,N_4971,N_477);
and U9578 (N_9578,N_4098,N_1645);
nor U9579 (N_9579,N_1054,N_3495);
nand U9580 (N_9580,N_3270,N_1480);
xnor U9581 (N_9581,N_1489,N_1876);
nor U9582 (N_9582,N_2150,N_3966);
xnor U9583 (N_9583,N_4129,N_4324);
and U9584 (N_9584,N_3675,N_1717);
or U9585 (N_9585,N_979,N_1744);
nor U9586 (N_9586,N_1943,N_4951);
nor U9587 (N_9587,N_2313,N_2739);
or U9588 (N_9588,N_3356,N_462);
nor U9589 (N_9589,N_2422,N_3915);
nor U9590 (N_9590,N_1915,N_2813);
xnor U9591 (N_9591,N_4744,N_1887);
xnor U9592 (N_9592,N_3791,N_4178);
xnor U9593 (N_9593,N_1608,N_2880);
and U9594 (N_9594,N_3069,N_2807);
or U9595 (N_9595,N_1973,N_4303);
xor U9596 (N_9596,N_4813,N_4741);
nor U9597 (N_9597,N_115,N_4637);
nor U9598 (N_9598,N_3877,N_1047);
or U9599 (N_9599,N_3997,N_3015);
xor U9600 (N_9600,N_4603,N_4181);
nor U9601 (N_9601,N_298,N_2703);
nor U9602 (N_9602,N_1609,N_4227);
nor U9603 (N_9603,N_4274,N_220);
and U9604 (N_9604,N_3621,N_163);
nor U9605 (N_9605,N_1666,N_2851);
nor U9606 (N_9606,N_2408,N_4613);
nor U9607 (N_9607,N_4836,N_82);
or U9608 (N_9608,N_2927,N_4945);
and U9609 (N_9609,N_600,N_4551);
nand U9610 (N_9610,N_1720,N_4653);
or U9611 (N_9611,N_399,N_2070);
nand U9612 (N_9612,N_2588,N_1239);
or U9613 (N_9613,N_1439,N_3005);
nor U9614 (N_9614,N_3282,N_3791);
or U9615 (N_9615,N_2503,N_4409);
and U9616 (N_9616,N_1774,N_2426);
xor U9617 (N_9617,N_2897,N_3805);
and U9618 (N_9618,N_3018,N_353);
xnor U9619 (N_9619,N_1613,N_1973);
nand U9620 (N_9620,N_3464,N_2615);
nor U9621 (N_9621,N_882,N_1328);
nor U9622 (N_9622,N_625,N_2560);
and U9623 (N_9623,N_1549,N_1669);
and U9624 (N_9624,N_3298,N_4651);
nand U9625 (N_9625,N_4188,N_3462);
nand U9626 (N_9626,N_233,N_3354);
nor U9627 (N_9627,N_3856,N_2380);
xor U9628 (N_9628,N_3315,N_1989);
xor U9629 (N_9629,N_4145,N_2246);
nor U9630 (N_9630,N_1457,N_4887);
nand U9631 (N_9631,N_3300,N_3607);
xnor U9632 (N_9632,N_1926,N_4379);
nand U9633 (N_9633,N_1742,N_4265);
xor U9634 (N_9634,N_2478,N_3416);
nand U9635 (N_9635,N_2699,N_757);
xor U9636 (N_9636,N_284,N_117);
nor U9637 (N_9637,N_3068,N_540);
and U9638 (N_9638,N_435,N_2828);
xnor U9639 (N_9639,N_3678,N_3886);
and U9640 (N_9640,N_2402,N_4676);
or U9641 (N_9641,N_3408,N_1477);
xor U9642 (N_9642,N_4376,N_636);
and U9643 (N_9643,N_408,N_2552);
or U9644 (N_9644,N_1121,N_2583);
nor U9645 (N_9645,N_3058,N_4349);
or U9646 (N_9646,N_4362,N_1953);
nand U9647 (N_9647,N_338,N_1829);
xor U9648 (N_9648,N_4085,N_2851);
and U9649 (N_9649,N_1120,N_1191);
nor U9650 (N_9650,N_4161,N_750);
xnor U9651 (N_9651,N_4091,N_1259);
or U9652 (N_9652,N_15,N_2142);
nand U9653 (N_9653,N_168,N_796);
and U9654 (N_9654,N_398,N_1873);
xnor U9655 (N_9655,N_1432,N_1715);
and U9656 (N_9656,N_3303,N_3150);
and U9657 (N_9657,N_4365,N_2785);
xnor U9658 (N_9658,N_4444,N_1064);
nand U9659 (N_9659,N_165,N_1328);
and U9660 (N_9660,N_1431,N_1863);
nand U9661 (N_9661,N_3958,N_3166);
or U9662 (N_9662,N_4092,N_1648);
xor U9663 (N_9663,N_305,N_347);
nand U9664 (N_9664,N_4796,N_3281);
and U9665 (N_9665,N_4877,N_2694);
nand U9666 (N_9666,N_464,N_4446);
and U9667 (N_9667,N_2666,N_972);
nand U9668 (N_9668,N_2471,N_2261);
xnor U9669 (N_9669,N_3601,N_1930);
nor U9670 (N_9670,N_720,N_1934);
and U9671 (N_9671,N_2741,N_534);
or U9672 (N_9672,N_200,N_1962);
or U9673 (N_9673,N_2146,N_2205);
nor U9674 (N_9674,N_2355,N_1313);
or U9675 (N_9675,N_2303,N_1292);
and U9676 (N_9676,N_263,N_3931);
xnor U9677 (N_9677,N_3591,N_664);
xnor U9678 (N_9678,N_4269,N_1371);
nand U9679 (N_9679,N_1412,N_462);
nand U9680 (N_9680,N_1276,N_2841);
and U9681 (N_9681,N_1358,N_2240);
xnor U9682 (N_9682,N_65,N_4933);
or U9683 (N_9683,N_3981,N_913);
nor U9684 (N_9684,N_4897,N_1260);
or U9685 (N_9685,N_1997,N_1841);
or U9686 (N_9686,N_3156,N_2198);
nand U9687 (N_9687,N_2367,N_4703);
nand U9688 (N_9688,N_2395,N_1065);
xnor U9689 (N_9689,N_4303,N_917);
xor U9690 (N_9690,N_4677,N_2721);
or U9691 (N_9691,N_1981,N_1121);
nand U9692 (N_9692,N_559,N_2279);
nor U9693 (N_9693,N_1400,N_2473);
nor U9694 (N_9694,N_1344,N_1326);
or U9695 (N_9695,N_4754,N_3551);
nand U9696 (N_9696,N_665,N_1520);
nor U9697 (N_9697,N_1978,N_2640);
or U9698 (N_9698,N_2695,N_2359);
xnor U9699 (N_9699,N_1517,N_1961);
nand U9700 (N_9700,N_4534,N_118);
or U9701 (N_9701,N_127,N_4947);
and U9702 (N_9702,N_4646,N_4179);
and U9703 (N_9703,N_251,N_1017);
nand U9704 (N_9704,N_818,N_3752);
nor U9705 (N_9705,N_4421,N_4742);
nand U9706 (N_9706,N_1676,N_219);
xor U9707 (N_9707,N_1949,N_3426);
nand U9708 (N_9708,N_1586,N_2858);
nand U9709 (N_9709,N_4612,N_3623);
and U9710 (N_9710,N_2251,N_2180);
nor U9711 (N_9711,N_2268,N_3868);
or U9712 (N_9712,N_2567,N_945);
nand U9713 (N_9713,N_2338,N_3849);
or U9714 (N_9714,N_1373,N_1225);
nor U9715 (N_9715,N_4069,N_4812);
or U9716 (N_9716,N_1173,N_1561);
or U9717 (N_9717,N_3197,N_724);
nand U9718 (N_9718,N_2399,N_2959);
nor U9719 (N_9719,N_144,N_2071);
and U9720 (N_9720,N_3636,N_4906);
nor U9721 (N_9721,N_1088,N_3165);
xnor U9722 (N_9722,N_519,N_4613);
and U9723 (N_9723,N_3225,N_3478);
xor U9724 (N_9724,N_4456,N_3123);
xnor U9725 (N_9725,N_436,N_4346);
nor U9726 (N_9726,N_3308,N_704);
or U9727 (N_9727,N_1688,N_3362);
nand U9728 (N_9728,N_1699,N_214);
and U9729 (N_9729,N_591,N_4733);
nor U9730 (N_9730,N_3044,N_3552);
nand U9731 (N_9731,N_1444,N_4540);
xnor U9732 (N_9732,N_2231,N_369);
or U9733 (N_9733,N_4280,N_3201);
xnor U9734 (N_9734,N_2678,N_119);
xnor U9735 (N_9735,N_4732,N_222);
nor U9736 (N_9736,N_877,N_1628);
nand U9737 (N_9737,N_4699,N_752);
xor U9738 (N_9738,N_1241,N_2533);
nand U9739 (N_9739,N_2668,N_2274);
or U9740 (N_9740,N_21,N_4767);
nand U9741 (N_9741,N_4476,N_4270);
or U9742 (N_9742,N_3366,N_4535);
and U9743 (N_9743,N_4783,N_4059);
nand U9744 (N_9744,N_2519,N_1065);
and U9745 (N_9745,N_4788,N_724);
xnor U9746 (N_9746,N_781,N_154);
nor U9747 (N_9747,N_781,N_2607);
xor U9748 (N_9748,N_4115,N_469);
nand U9749 (N_9749,N_3359,N_1256);
and U9750 (N_9750,N_4973,N_4733);
and U9751 (N_9751,N_3675,N_3180);
or U9752 (N_9752,N_250,N_2061);
or U9753 (N_9753,N_59,N_4260);
xnor U9754 (N_9754,N_1385,N_1276);
or U9755 (N_9755,N_4051,N_4357);
and U9756 (N_9756,N_2334,N_3848);
or U9757 (N_9757,N_4260,N_1079);
or U9758 (N_9758,N_1009,N_290);
xor U9759 (N_9759,N_3672,N_505);
nand U9760 (N_9760,N_749,N_3934);
and U9761 (N_9761,N_3558,N_1988);
or U9762 (N_9762,N_737,N_1532);
xor U9763 (N_9763,N_747,N_600);
or U9764 (N_9764,N_310,N_38);
nor U9765 (N_9765,N_2042,N_4495);
nor U9766 (N_9766,N_3569,N_757);
xnor U9767 (N_9767,N_2774,N_4716);
or U9768 (N_9768,N_418,N_4309);
xor U9769 (N_9769,N_2818,N_2149);
nand U9770 (N_9770,N_4862,N_2080);
nand U9771 (N_9771,N_1001,N_788);
and U9772 (N_9772,N_4722,N_1269);
nand U9773 (N_9773,N_1943,N_2748);
or U9774 (N_9774,N_3094,N_3758);
nand U9775 (N_9775,N_3479,N_2186);
xor U9776 (N_9776,N_3705,N_249);
nor U9777 (N_9777,N_3051,N_3146);
nand U9778 (N_9778,N_1252,N_4862);
and U9779 (N_9779,N_4982,N_3497);
or U9780 (N_9780,N_4205,N_4295);
or U9781 (N_9781,N_1609,N_4420);
and U9782 (N_9782,N_2274,N_3724);
or U9783 (N_9783,N_3759,N_4381);
xnor U9784 (N_9784,N_2103,N_50);
or U9785 (N_9785,N_2483,N_232);
xor U9786 (N_9786,N_2725,N_3758);
xor U9787 (N_9787,N_2882,N_2676);
xor U9788 (N_9788,N_1180,N_3131);
xor U9789 (N_9789,N_2475,N_1238);
xnor U9790 (N_9790,N_3979,N_4961);
or U9791 (N_9791,N_778,N_657);
nor U9792 (N_9792,N_1947,N_2606);
and U9793 (N_9793,N_786,N_2398);
nor U9794 (N_9794,N_2655,N_2729);
nand U9795 (N_9795,N_3367,N_2452);
nor U9796 (N_9796,N_3606,N_4778);
and U9797 (N_9797,N_4024,N_1698);
nand U9798 (N_9798,N_1003,N_4123);
nor U9799 (N_9799,N_1974,N_4389);
nand U9800 (N_9800,N_1337,N_4341);
xor U9801 (N_9801,N_184,N_2898);
xor U9802 (N_9802,N_4386,N_1371);
or U9803 (N_9803,N_3924,N_2056);
nor U9804 (N_9804,N_95,N_3383);
nand U9805 (N_9805,N_3712,N_4459);
and U9806 (N_9806,N_4640,N_4875);
nand U9807 (N_9807,N_93,N_4809);
xnor U9808 (N_9808,N_1875,N_3799);
nand U9809 (N_9809,N_506,N_4536);
nor U9810 (N_9810,N_3740,N_2354);
nor U9811 (N_9811,N_3029,N_1492);
xor U9812 (N_9812,N_3115,N_4124);
nand U9813 (N_9813,N_653,N_3695);
xor U9814 (N_9814,N_94,N_1837);
xnor U9815 (N_9815,N_4320,N_277);
or U9816 (N_9816,N_566,N_3709);
and U9817 (N_9817,N_29,N_3039);
xor U9818 (N_9818,N_3573,N_1917);
and U9819 (N_9819,N_3164,N_4399);
nor U9820 (N_9820,N_7,N_3902);
and U9821 (N_9821,N_771,N_2551);
nand U9822 (N_9822,N_2326,N_1137);
nand U9823 (N_9823,N_1078,N_3681);
or U9824 (N_9824,N_245,N_519);
xor U9825 (N_9825,N_1309,N_3294);
nor U9826 (N_9826,N_1734,N_4634);
or U9827 (N_9827,N_2282,N_618);
nor U9828 (N_9828,N_1720,N_2138);
nand U9829 (N_9829,N_3695,N_4811);
xnor U9830 (N_9830,N_23,N_3223);
and U9831 (N_9831,N_4109,N_199);
nor U9832 (N_9832,N_3186,N_4123);
nor U9833 (N_9833,N_199,N_3926);
nor U9834 (N_9834,N_708,N_4371);
and U9835 (N_9835,N_1345,N_1652);
and U9836 (N_9836,N_1444,N_1508);
or U9837 (N_9837,N_3007,N_3737);
nand U9838 (N_9838,N_2967,N_1354);
nand U9839 (N_9839,N_1257,N_3116);
and U9840 (N_9840,N_3183,N_129);
or U9841 (N_9841,N_2697,N_965);
nand U9842 (N_9842,N_711,N_4837);
nor U9843 (N_9843,N_1767,N_3246);
xnor U9844 (N_9844,N_2237,N_4316);
or U9845 (N_9845,N_3667,N_143);
nand U9846 (N_9846,N_4123,N_3266);
or U9847 (N_9847,N_252,N_3309);
xnor U9848 (N_9848,N_2923,N_4629);
nand U9849 (N_9849,N_836,N_3578);
nor U9850 (N_9850,N_3547,N_2246);
xnor U9851 (N_9851,N_3203,N_943);
and U9852 (N_9852,N_586,N_1648);
xnor U9853 (N_9853,N_605,N_3714);
nand U9854 (N_9854,N_781,N_1203);
xor U9855 (N_9855,N_1550,N_2908);
nor U9856 (N_9856,N_449,N_2342);
or U9857 (N_9857,N_2261,N_1382);
nand U9858 (N_9858,N_2645,N_2306);
xor U9859 (N_9859,N_295,N_2113);
nand U9860 (N_9860,N_1245,N_3084);
nor U9861 (N_9861,N_4086,N_4942);
nand U9862 (N_9862,N_2306,N_291);
or U9863 (N_9863,N_1001,N_2486);
xnor U9864 (N_9864,N_4207,N_149);
nor U9865 (N_9865,N_1130,N_3518);
xor U9866 (N_9866,N_580,N_2571);
nor U9867 (N_9867,N_319,N_4056);
and U9868 (N_9868,N_1067,N_3477);
xnor U9869 (N_9869,N_2516,N_1809);
or U9870 (N_9870,N_4265,N_1769);
nand U9871 (N_9871,N_2711,N_518);
and U9872 (N_9872,N_208,N_237);
xor U9873 (N_9873,N_786,N_2575);
xnor U9874 (N_9874,N_1644,N_4366);
or U9875 (N_9875,N_1872,N_4381);
xnor U9876 (N_9876,N_3915,N_1737);
nor U9877 (N_9877,N_4197,N_4518);
or U9878 (N_9878,N_1965,N_219);
nor U9879 (N_9879,N_134,N_1453);
or U9880 (N_9880,N_3680,N_4364);
nand U9881 (N_9881,N_3704,N_2869);
and U9882 (N_9882,N_3933,N_4072);
xnor U9883 (N_9883,N_4746,N_4569);
xnor U9884 (N_9884,N_4034,N_1557);
nor U9885 (N_9885,N_685,N_4371);
xor U9886 (N_9886,N_977,N_404);
nor U9887 (N_9887,N_313,N_1453);
xor U9888 (N_9888,N_1048,N_64);
nand U9889 (N_9889,N_3228,N_3501);
xor U9890 (N_9890,N_456,N_2784);
nand U9891 (N_9891,N_4596,N_3214);
nand U9892 (N_9892,N_740,N_3199);
xnor U9893 (N_9893,N_42,N_561);
or U9894 (N_9894,N_3197,N_294);
nor U9895 (N_9895,N_1632,N_2750);
nand U9896 (N_9896,N_4225,N_4235);
nand U9897 (N_9897,N_3120,N_4035);
or U9898 (N_9898,N_4481,N_216);
nor U9899 (N_9899,N_999,N_2556);
xor U9900 (N_9900,N_1677,N_3615);
nor U9901 (N_9901,N_2451,N_759);
or U9902 (N_9902,N_872,N_518);
or U9903 (N_9903,N_4788,N_1946);
and U9904 (N_9904,N_4702,N_2762);
and U9905 (N_9905,N_1759,N_1284);
or U9906 (N_9906,N_4639,N_2088);
xnor U9907 (N_9907,N_3552,N_3447);
or U9908 (N_9908,N_4320,N_4317);
nand U9909 (N_9909,N_157,N_4978);
xor U9910 (N_9910,N_4534,N_4336);
xnor U9911 (N_9911,N_3366,N_4910);
nand U9912 (N_9912,N_4765,N_438);
and U9913 (N_9913,N_2343,N_3720);
nor U9914 (N_9914,N_1649,N_3733);
nor U9915 (N_9915,N_2634,N_516);
nand U9916 (N_9916,N_2880,N_2966);
nor U9917 (N_9917,N_791,N_4172);
nor U9918 (N_9918,N_3821,N_1015);
and U9919 (N_9919,N_475,N_4185);
and U9920 (N_9920,N_1718,N_4731);
nand U9921 (N_9921,N_2425,N_1146);
xnor U9922 (N_9922,N_2664,N_699);
xor U9923 (N_9923,N_4914,N_2395);
and U9924 (N_9924,N_583,N_3535);
nand U9925 (N_9925,N_4781,N_1201);
xnor U9926 (N_9926,N_1191,N_4393);
nand U9927 (N_9927,N_2386,N_1664);
or U9928 (N_9928,N_2895,N_391);
and U9929 (N_9929,N_1348,N_2558);
and U9930 (N_9930,N_3736,N_2015);
nand U9931 (N_9931,N_2925,N_3092);
xnor U9932 (N_9932,N_2800,N_1822);
nand U9933 (N_9933,N_940,N_805);
xnor U9934 (N_9934,N_4826,N_2012);
or U9935 (N_9935,N_1489,N_4712);
nor U9936 (N_9936,N_4576,N_1898);
and U9937 (N_9937,N_1884,N_4088);
xor U9938 (N_9938,N_2065,N_1090);
nand U9939 (N_9939,N_759,N_4581);
nand U9940 (N_9940,N_2837,N_3073);
xor U9941 (N_9941,N_3139,N_4288);
nor U9942 (N_9942,N_4627,N_48);
and U9943 (N_9943,N_1407,N_1834);
nor U9944 (N_9944,N_2788,N_2365);
nand U9945 (N_9945,N_2596,N_4190);
or U9946 (N_9946,N_4155,N_1059);
xnor U9947 (N_9947,N_3603,N_4118);
nand U9948 (N_9948,N_2311,N_4630);
and U9949 (N_9949,N_2757,N_3784);
nor U9950 (N_9950,N_132,N_4690);
or U9951 (N_9951,N_3499,N_3211);
nor U9952 (N_9952,N_4822,N_4849);
nor U9953 (N_9953,N_4855,N_2425);
xnor U9954 (N_9954,N_3498,N_2115);
nor U9955 (N_9955,N_4015,N_412);
nand U9956 (N_9956,N_4045,N_3084);
nand U9957 (N_9957,N_3504,N_2062);
and U9958 (N_9958,N_4054,N_225);
nor U9959 (N_9959,N_3593,N_4262);
or U9960 (N_9960,N_2655,N_4260);
nor U9961 (N_9961,N_825,N_2066);
xnor U9962 (N_9962,N_2227,N_2231);
or U9963 (N_9963,N_1699,N_2864);
nand U9964 (N_9964,N_4833,N_4730);
nand U9965 (N_9965,N_2522,N_4138);
or U9966 (N_9966,N_3048,N_974);
nor U9967 (N_9967,N_2863,N_341);
nand U9968 (N_9968,N_4288,N_2626);
xnor U9969 (N_9969,N_4059,N_2055);
nand U9970 (N_9970,N_511,N_4178);
and U9971 (N_9971,N_3494,N_685);
nor U9972 (N_9972,N_4261,N_1949);
and U9973 (N_9973,N_319,N_4981);
and U9974 (N_9974,N_4723,N_4195);
and U9975 (N_9975,N_2828,N_3523);
and U9976 (N_9976,N_4474,N_1733);
xor U9977 (N_9977,N_1937,N_770);
xnor U9978 (N_9978,N_3127,N_2611);
xnor U9979 (N_9979,N_1286,N_4665);
nand U9980 (N_9980,N_631,N_4475);
xnor U9981 (N_9981,N_3860,N_2006);
or U9982 (N_9982,N_1562,N_2688);
or U9983 (N_9983,N_1344,N_1787);
xnor U9984 (N_9984,N_230,N_2214);
nor U9985 (N_9985,N_809,N_4872);
nand U9986 (N_9986,N_4794,N_3253);
nor U9987 (N_9987,N_4206,N_1209);
xor U9988 (N_9988,N_4054,N_4024);
xor U9989 (N_9989,N_3751,N_2990);
xor U9990 (N_9990,N_1595,N_1179);
nor U9991 (N_9991,N_23,N_2698);
nand U9992 (N_9992,N_2938,N_349);
and U9993 (N_9993,N_3176,N_1266);
or U9994 (N_9994,N_200,N_4787);
or U9995 (N_9995,N_2432,N_1235);
xor U9996 (N_9996,N_3342,N_2401);
or U9997 (N_9997,N_1367,N_4243);
xnor U9998 (N_9998,N_93,N_1198);
or U9999 (N_9999,N_2958,N_2988);
nand UO_0 (O_0,N_6753,N_5021);
xnor UO_1 (O_1,N_9548,N_8419);
or UO_2 (O_2,N_5548,N_9482);
nor UO_3 (O_3,N_9701,N_6404);
or UO_4 (O_4,N_7945,N_5527);
or UO_5 (O_5,N_8351,N_8235);
nor UO_6 (O_6,N_9216,N_6090);
xor UO_7 (O_7,N_7811,N_7166);
or UO_8 (O_8,N_5278,N_9159);
nand UO_9 (O_9,N_5448,N_7459);
xnor UO_10 (O_10,N_7899,N_9348);
nand UO_11 (O_11,N_7887,N_5765);
xor UO_12 (O_12,N_7044,N_8829);
xor UO_13 (O_13,N_8137,N_7408);
nor UO_14 (O_14,N_8818,N_7805);
nand UO_15 (O_15,N_9615,N_8900);
nand UO_16 (O_16,N_7971,N_7313);
or UO_17 (O_17,N_6385,N_7630);
nor UO_18 (O_18,N_9625,N_8110);
nor UO_19 (O_19,N_8053,N_7696);
or UO_20 (O_20,N_8260,N_9765);
nand UO_21 (O_21,N_9783,N_7417);
and UO_22 (O_22,N_8734,N_9359);
xor UO_23 (O_23,N_5734,N_9374);
and UO_24 (O_24,N_8198,N_5222);
xor UO_25 (O_25,N_5204,N_9023);
nor UO_26 (O_26,N_6507,N_5939);
nor UO_27 (O_27,N_6713,N_9954);
nand UO_28 (O_28,N_5687,N_9907);
nand UO_29 (O_29,N_5434,N_7826);
nor UO_30 (O_30,N_9455,N_6030);
xnor UO_31 (O_31,N_8787,N_6707);
or UO_32 (O_32,N_9798,N_5975);
nand UO_33 (O_33,N_6551,N_8625);
or UO_34 (O_34,N_5624,N_9763);
nand UO_35 (O_35,N_5809,N_5369);
or UO_36 (O_36,N_5449,N_9600);
nand UO_37 (O_37,N_5184,N_5927);
xnor UO_38 (O_38,N_6122,N_6828);
xnor UO_39 (O_39,N_6422,N_5641);
nand UO_40 (O_40,N_9900,N_7588);
or UO_41 (O_41,N_7854,N_6176);
and UO_42 (O_42,N_8706,N_6668);
nand UO_43 (O_43,N_8055,N_7908);
xnor UO_44 (O_44,N_6718,N_6793);
nor UO_45 (O_45,N_9397,N_7426);
nand UO_46 (O_46,N_9779,N_6307);
and UO_47 (O_47,N_6169,N_5318);
nor UO_48 (O_48,N_7086,N_7098);
nor UO_49 (O_49,N_9093,N_9597);
and UO_50 (O_50,N_5831,N_8909);
nor UO_51 (O_51,N_8214,N_6313);
nand UO_52 (O_52,N_8553,N_6000);
and UO_53 (O_53,N_7866,N_5938);
or UO_54 (O_54,N_5471,N_8381);
and UO_55 (O_55,N_8789,N_7194);
xnor UO_56 (O_56,N_7285,N_8398);
xor UO_57 (O_57,N_5494,N_9363);
and UO_58 (O_58,N_7025,N_5428);
and UO_59 (O_59,N_6990,N_8317);
xnor UO_60 (O_60,N_8019,N_8643);
nor UO_61 (O_61,N_9380,N_8512);
or UO_62 (O_62,N_9558,N_8938);
nor UO_63 (O_63,N_5403,N_6433);
or UO_64 (O_64,N_9022,N_5165);
nand UO_65 (O_65,N_5045,N_5245);
and UO_66 (O_66,N_9098,N_8997);
nor UO_67 (O_67,N_6518,N_8407);
nor UO_68 (O_68,N_6391,N_6912);
or UO_69 (O_69,N_6850,N_9471);
nand UO_70 (O_70,N_7967,N_8362);
nand UO_71 (O_71,N_6006,N_9107);
nor UO_72 (O_72,N_7453,N_7316);
nor UO_73 (O_73,N_6166,N_9044);
nor UO_74 (O_74,N_6631,N_6460);
nand UO_75 (O_75,N_8896,N_6808);
and UO_76 (O_76,N_7160,N_5489);
and UO_77 (O_77,N_9459,N_5712);
and UO_78 (O_78,N_6800,N_6175);
nand UO_79 (O_79,N_8437,N_6361);
xor UO_80 (O_80,N_9028,N_7537);
and UO_81 (O_81,N_6048,N_6854);
xor UO_82 (O_82,N_6539,N_8733);
nor UO_83 (O_83,N_9539,N_9543);
or UO_84 (O_84,N_8810,N_9187);
nor UO_85 (O_85,N_5729,N_7363);
or UO_86 (O_86,N_9852,N_5492);
and UO_87 (O_87,N_9723,N_8422);
xor UO_88 (O_88,N_8729,N_7484);
nor UO_89 (O_89,N_9727,N_8052);
or UO_90 (O_90,N_6229,N_6192);
or UO_91 (O_91,N_5460,N_9859);
and UO_92 (O_92,N_5363,N_5518);
or UO_93 (O_93,N_7578,N_5197);
or UO_94 (O_94,N_8468,N_5886);
and UO_95 (O_95,N_7419,N_9583);
or UO_96 (O_96,N_7250,N_7172);
nor UO_97 (O_97,N_5968,N_7163);
xnor UO_98 (O_98,N_6418,N_5964);
nand UO_99 (O_99,N_6237,N_9752);
and UO_100 (O_100,N_6240,N_6023);
nand UO_101 (O_101,N_5485,N_7557);
or UO_102 (O_102,N_7847,N_6680);
and UO_103 (O_103,N_7757,N_5237);
nor UO_104 (O_104,N_7970,N_7850);
or UO_105 (O_105,N_9520,N_7657);
and UO_106 (O_106,N_9010,N_7185);
nand UO_107 (O_107,N_9166,N_5782);
nand UO_108 (O_108,N_7010,N_7526);
nand UO_109 (O_109,N_7771,N_5093);
and UO_110 (O_110,N_7695,N_7931);
nor UO_111 (O_111,N_9799,N_9608);
xnor UO_112 (O_112,N_5496,N_8460);
and UO_113 (O_113,N_8825,N_6232);
xnor UO_114 (O_114,N_9386,N_9494);
xor UO_115 (O_115,N_7183,N_9104);
nor UO_116 (O_116,N_5678,N_6403);
and UO_117 (O_117,N_9729,N_5118);
xor UO_118 (O_118,N_8673,N_5436);
nand UO_119 (O_119,N_8305,N_7164);
and UO_120 (O_120,N_8324,N_6630);
nor UO_121 (O_121,N_7875,N_6665);
or UO_122 (O_122,N_8543,N_7294);
nor UO_123 (O_123,N_5216,N_8363);
xor UO_124 (O_124,N_5928,N_9913);
xor UO_125 (O_125,N_6210,N_6413);
nand UO_126 (O_126,N_5064,N_5374);
and UO_127 (O_127,N_5498,N_5913);
nor UO_128 (O_128,N_9559,N_9129);
nand UO_129 (O_129,N_6788,N_8794);
nand UO_130 (O_130,N_5648,N_6969);
nor UO_131 (O_131,N_9309,N_7404);
and UO_132 (O_132,N_8336,N_8975);
and UO_133 (O_133,N_6435,N_6448);
and UO_134 (O_134,N_9510,N_5901);
and UO_135 (O_135,N_6659,N_5852);
or UO_136 (O_136,N_6271,N_6544);
or UO_137 (O_137,N_6339,N_5589);
nand UO_138 (O_138,N_9694,N_9419);
xor UO_139 (O_139,N_8385,N_9972);
or UO_140 (O_140,N_6337,N_9434);
or UO_141 (O_141,N_6841,N_5880);
and UO_142 (O_142,N_9285,N_5283);
nor UO_143 (O_143,N_9432,N_8780);
or UO_144 (O_144,N_7990,N_8189);
nor UO_145 (O_145,N_5170,N_6524);
and UO_146 (O_146,N_7151,N_7447);
or UO_147 (O_147,N_6728,N_8840);
and UO_148 (O_148,N_7056,N_6195);
nand UO_149 (O_149,N_7838,N_5607);
xor UO_150 (O_150,N_6615,N_6469);
xor UO_151 (O_151,N_6264,N_6275);
and UO_152 (O_152,N_8387,N_6720);
nand UO_153 (O_153,N_8392,N_6744);
or UO_154 (O_154,N_7514,N_5080);
nand UO_155 (O_155,N_7964,N_5925);
nor UO_156 (O_156,N_8708,N_7753);
nand UO_157 (O_157,N_5583,N_7744);
nand UO_158 (O_158,N_7018,N_7522);
nor UO_159 (O_159,N_5579,N_9998);
nor UO_160 (O_160,N_7431,N_8233);
nor UO_161 (O_161,N_9130,N_8481);
nor UO_162 (O_162,N_6031,N_8891);
and UO_163 (O_163,N_6203,N_5704);
nor UO_164 (O_164,N_6407,N_8890);
and UO_165 (O_165,N_5644,N_9986);
or UO_166 (O_166,N_9127,N_7305);
or UO_167 (O_167,N_8692,N_9938);
and UO_168 (O_168,N_6278,N_7125);
and UO_169 (O_169,N_8131,N_7535);
and UO_170 (O_170,N_7690,N_9525);
nor UO_171 (O_171,N_6400,N_8998);
xor UO_172 (O_172,N_8848,N_8372);
and UO_173 (O_173,N_7254,N_6346);
or UO_174 (O_174,N_9619,N_8313);
nor UO_175 (O_175,N_7807,N_6709);
nor UO_176 (O_176,N_7033,N_7400);
xor UO_177 (O_177,N_8176,N_5793);
xnor UO_178 (O_178,N_7533,N_5025);
or UO_179 (O_179,N_7213,N_9496);
and UO_180 (O_180,N_7559,N_7774);
nand UO_181 (O_181,N_5352,N_7874);
nand UO_182 (O_182,N_8161,N_9326);
xor UO_183 (O_183,N_6129,N_8528);
xor UO_184 (O_184,N_7984,N_5185);
nor UO_185 (O_185,N_5625,N_5999);
nor UO_186 (O_186,N_7245,N_9706);
xor UO_187 (O_187,N_8653,N_6685);
xnor UO_188 (O_188,N_9086,N_6671);
nor UO_189 (O_189,N_9606,N_8803);
and UO_190 (O_190,N_7653,N_9826);
and UO_191 (O_191,N_7820,N_7269);
or UO_192 (O_192,N_9568,N_7693);
nor UO_193 (O_193,N_6780,N_9320);
nor UO_194 (O_194,N_6170,N_5157);
or UO_195 (O_195,N_5982,N_5102);
nor UO_196 (O_196,N_9111,N_7237);
xor UO_197 (O_197,N_6927,N_5243);
nand UO_198 (O_198,N_7336,N_5385);
nor UO_199 (O_199,N_8159,N_7819);
nor UO_200 (O_200,N_8472,N_8112);
and UO_201 (O_201,N_5382,N_9045);
nand UO_202 (O_202,N_7692,N_9810);
xnor UO_203 (O_203,N_7446,N_7745);
or UO_204 (O_204,N_6660,N_9056);
xor UO_205 (O_205,N_8406,N_6546);
nand UO_206 (O_206,N_9709,N_8217);
or UO_207 (O_207,N_6576,N_6078);
and UO_208 (O_208,N_5890,N_6714);
and UO_209 (O_209,N_8784,N_8330);
nor UO_210 (O_210,N_7620,N_9161);
and UO_211 (O_211,N_9750,N_7528);
and UO_212 (O_212,N_8255,N_8199);
xor UO_213 (O_213,N_9470,N_5394);
and UO_214 (O_214,N_7199,N_6255);
xor UO_215 (O_215,N_9435,N_6848);
nand UO_216 (O_216,N_8721,N_8854);
nor UO_217 (O_217,N_8990,N_8246);
or UO_218 (O_218,N_6590,N_9152);
nand UO_219 (O_219,N_6749,N_9576);
nand UO_220 (O_220,N_5662,N_5430);
nor UO_221 (O_221,N_9282,N_8124);
or UO_222 (O_222,N_7794,N_9401);
xnor UO_223 (O_223,N_6710,N_6269);
nand UO_224 (O_224,N_5787,N_8169);
or UO_225 (O_225,N_5346,N_8262);
xor UO_226 (O_226,N_6062,N_7302);
or UO_227 (O_227,N_9231,N_8088);
nor UO_228 (O_228,N_9399,N_9812);
or UO_229 (O_229,N_8428,N_9295);
xor UO_230 (O_230,N_9145,N_7561);
and UO_231 (O_231,N_8004,N_6751);
nand UO_232 (O_232,N_6624,N_7165);
and UO_233 (O_233,N_7715,N_8342);
xnor UO_234 (O_234,N_6620,N_6135);
nor UO_235 (O_235,N_8257,N_9180);
and UO_236 (O_236,N_7995,N_9719);
xor UO_237 (O_237,N_6980,N_9513);
and UO_238 (O_238,N_5072,N_5701);
and UO_239 (O_239,N_5384,N_6046);
and UO_240 (O_240,N_8267,N_8357);
and UO_241 (O_241,N_6790,N_6627);
nand UO_242 (O_242,N_8878,N_6016);
nor UO_243 (O_243,N_8598,N_8704);
and UO_244 (O_244,N_8805,N_6686);
or UO_245 (O_245,N_6251,N_6938);
xor UO_246 (O_246,N_6497,N_5275);
or UO_247 (O_247,N_7109,N_9444);
xnor UO_248 (O_248,N_7047,N_9317);
nand UO_249 (O_249,N_5029,N_7394);
or UO_250 (O_250,N_9906,N_9036);
nor UO_251 (O_251,N_6849,N_6243);
and UO_252 (O_252,N_7116,N_9741);
nand UO_253 (O_253,N_5280,N_7441);
or UO_254 (O_254,N_6944,N_5424);
and UO_255 (O_255,N_6430,N_8005);
xnor UO_256 (O_256,N_7925,N_7677);
xnor UO_257 (O_257,N_9410,N_7396);
or UO_258 (O_258,N_5177,N_7576);
and UO_259 (O_259,N_8326,N_8648);
nor UO_260 (O_260,N_7065,N_8630);
nor UO_261 (O_261,N_8226,N_5180);
nor UO_262 (O_262,N_6677,N_6410);
nand UO_263 (O_263,N_6646,N_8934);
and UO_264 (O_264,N_8722,N_7597);
xor UO_265 (O_265,N_9966,N_5561);
or UO_266 (O_266,N_7052,N_8663);
or UO_267 (O_267,N_9668,N_8957);
nand UO_268 (O_268,N_7287,N_6241);
nor UO_269 (O_269,N_7729,N_5876);
or UO_270 (O_270,N_6412,N_6272);
nand UO_271 (O_271,N_9041,N_7023);
nor UO_272 (O_272,N_5164,N_6569);
nand UO_273 (O_273,N_6520,N_5877);
nand UO_274 (O_274,N_5539,N_5077);
nand UO_275 (O_275,N_8929,N_9464);
nand UO_276 (O_276,N_7439,N_7747);
or UO_277 (O_277,N_6058,N_5910);
or UO_278 (O_278,N_9047,N_7605);
nor UO_279 (O_279,N_7594,N_6308);
xor UO_280 (O_280,N_5630,N_9638);
xor UO_281 (O_281,N_8259,N_9404);
nand UO_282 (O_282,N_9795,N_8290);
xor UO_283 (O_283,N_7349,N_9774);
and UO_284 (O_284,N_8056,N_7144);
nor UO_285 (O_285,N_6020,N_9903);
and UO_286 (O_286,N_7223,N_9015);
and UO_287 (O_287,N_5688,N_6597);
and UO_288 (O_288,N_6865,N_9509);
xnor UO_289 (O_289,N_7765,N_9845);
and UO_290 (O_290,N_8429,N_6312);
nand UO_291 (O_291,N_9552,N_9014);
xor UO_292 (O_292,N_8862,N_9521);
or UO_293 (O_293,N_5673,N_6343);
or UO_294 (O_294,N_9681,N_7529);
nor UO_295 (O_295,N_5882,N_7937);
or UO_296 (O_296,N_9495,N_9195);
nor UO_297 (O_297,N_7095,N_7618);
or UO_298 (O_298,N_6155,N_7226);
and UO_299 (O_299,N_6739,N_6476);
and UO_300 (O_300,N_5138,N_8827);
and UO_301 (O_301,N_9655,N_6536);
or UO_302 (O_302,N_7062,N_5404);
xnor UO_303 (O_303,N_7872,N_6740);
nor UO_304 (O_304,N_9112,N_9124);
nor UO_305 (O_305,N_6970,N_6113);
or UO_306 (O_306,N_6382,N_6557);
xnor UO_307 (O_307,N_8390,N_9956);
nor UO_308 (O_308,N_6178,N_6010);
nor UO_309 (O_309,N_8048,N_9987);
and UO_310 (O_310,N_7545,N_5103);
nor UO_311 (O_311,N_9125,N_6880);
and UO_312 (O_312,N_8602,N_8699);
nand UO_313 (O_313,N_8339,N_5005);
and UO_314 (O_314,N_6570,N_7092);
nand UO_315 (O_315,N_5270,N_9747);
xnor UO_316 (O_316,N_5349,N_5050);
xnor UO_317 (O_317,N_5807,N_6366);
and UO_318 (O_318,N_6165,N_5848);
and UO_319 (O_319,N_5051,N_6290);
xor UO_320 (O_320,N_8358,N_5996);
nor UO_321 (O_321,N_5450,N_5043);
and UO_322 (O_322,N_9880,N_8254);
nor UO_323 (O_323,N_5918,N_6877);
nand UO_324 (O_324,N_6561,N_7943);
nor UO_325 (O_325,N_6652,N_6015);
and UO_326 (O_326,N_5653,N_9220);
or UO_327 (O_327,N_9665,N_6563);
xnor UO_328 (O_328,N_8637,N_8686);
xnor UO_329 (O_329,N_5954,N_8828);
and UO_330 (O_330,N_9328,N_5730);
and UO_331 (O_331,N_5841,N_5140);
or UO_332 (O_332,N_7667,N_5895);
xor UO_333 (O_333,N_7880,N_5778);
nand UO_334 (O_334,N_6644,N_6289);
nand UO_335 (O_335,N_6138,N_6968);
nor UO_336 (O_336,N_6967,N_6260);
nand UO_337 (O_337,N_7391,N_9275);
nor UO_338 (O_338,N_6383,N_8202);
nand UO_339 (O_339,N_6765,N_7112);
or UO_340 (O_340,N_5401,N_5478);
nand UO_341 (O_341,N_5231,N_9685);
xnor UO_342 (O_342,N_7768,N_5547);
xnor UO_343 (O_343,N_8936,N_9153);
nand UO_344 (O_344,N_5297,N_7057);
nor UO_345 (O_345,N_7622,N_7737);
xor UO_346 (O_346,N_7562,N_7048);
nand UO_347 (O_347,N_7483,N_7784);
xor UO_348 (O_348,N_8774,N_8824);
nor UO_349 (O_349,N_6319,N_6835);
nor UO_350 (O_350,N_6108,N_9265);
and UO_351 (O_351,N_9267,N_5720);
xor UO_352 (O_352,N_9114,N_9433);
or UO_353 (O_353,N_5463,N_5637);
nand UO_354 (O_354,N_6784,N_9686);
and UO_355 (O_355,N_5402,N_6691);
nand UO_356 (O_356,N_7389,N_6654);
xor UO_357 (O_357,N_9514,N_9310);
and UO_358 (O_358,N_9942,N_6089);
or UO_359 (O_359,N_7403,N_6249);
nand UO_360 (O_360,N_5405,N_7468);
or UO_361 (O_361,N_8961,N_6045);
or UO_362 (O_362,N_8670,N_6589);
and UO_363 (O_363,N_9883,N_9322);
and UO_364 (O_364,N_6099,N_9416);
and UO_365 (O_365,N_7688,N_5748);
nand UO_366 (O_366,N_9622,N_7407);
and UO_367 (O_367,N_8083,N_6294);
or UO_368 (O_368,N_9203,N_9738);
and UO_369 (O_369,N_7708,N_7944);
nand UO_370 (O_370,N_7210,N_9664);
xnor UO_371 (O_371,N_8477,N_6106);
nand UO_372 (O_372,N_6945,N_9767);
or UO_373 (O_373,N_7006,N_7523);
nor UO_374 (O_374,N_6256,N_6925);
xor UO_375 (O_375,N_6226,N_7954);
or UO_376 (O_376,N_9991,N_5221);
nand UO_377 (O_377,N_6457,N_8695);
nand UO_378 (O_378,N_5309,N_7186);
or UO_379 (O_379,N_7131,N_5879);
nand UO_380 (O_380,N_5109,N_5024);
and UO_381 (O_381,N_9882,N_8748);
or UO_382 (O_382,N_9189,N_7184);
or UO_383 (O_383,N_9780,N_8109);
and UO_384 (O_384,N_5040,N_6986);
or UO_385 (O_385,N_8714,N_5266);
nor UO_386 (O_386,N_5422,N_5065);
nor UO_387 (O_387,N_8937,N_6059);
nor UO_388 (O_388,N_8133,N_9209);
and UO_389 (O_389,N_6284,N_6856);
or UO_390 (O_390,N_7938,N_5739);
or UO_391 (O_391,N_5702,N_6658);
nor UO_392 (O_392,N_9451,N_8591);
and UO_393 (O_393,N_8275,N_9029);
and UO_394 (O_394,N_9052,N_8902);
nor UO_395 (O_395,N_8544,N_5724);
nand UO_396 (O_396,N_7904,N_6712);
nor UO_397 (O_397,N_5151,N_7743);
xnor UO_398 (O_398,N_7359,N_9946);
or UO_399 (O_399,N_5731,N_8893);
or UO_400 (O_400,N_9092,N_9866);
or UO_401 (O_401,N_5257,N_9289);
nor UO_402 (O_402,N_5797,N_5055);
and UO_403 (O_403,N_9895,N_6748);
nand UO_404 (O_404,N_9488,N_5059);
nand UO_405 (O_405,N_8626,N_9612);
nand UO_406 (O_406,N_8302,N_8979);
or UO_407 (O_407,N_9672,N_5903);
xor UO_408 (O_408,N_5282,N_9137);
xor UO_409 (O_409,N_9313,N_9553);
xnor UO_410 (O_410,N_6891,N_8730);
or UO_411 (O_411,N_5792,N_8234);
and UO_412 (O_412,N_6973,N_9039);
or UO_413 (O_413,N_5290,N_5885);
nand UO_414 (O_414,N_8391,N_9575);
nor UO_415 (O_415,N_9393,N_7353);
xor UO_416 (O_416,N_7783,N_6322);
and UO_417 (O_417,N_7267,N_8981);
xor UO_418 (O_418,N_9046,N_7542);
xnor UO_419 (O_419,N_6745,N_9083);
xor UO_420 (O_420,N_7883,N_6074);
and UO_421 (O_421,N_8657,N_8839);
nor UO_422 (O_422,N_9985,N_8098);
nor UO_423 (O_423,N_8037,N_8329);
nor UO_424 (O_424,N_8930,N_8006);
nor UO_425 (O_425,N_6838,N_7231);
nand UO_426 (O_426,N_8823,N_8622);
and UO_427 (O_427,N_5443,N_6224);
and UO_428 (O_428,N_5468,N_5322);
or UO_429 (O_429,N_5054,N_6402);
and UO_430 (O_430,N_8366,N_6505);
xor UO_431 (O_431,N_5336,N_5671);
or UO_432 (O_432,N_9332,N_7437);
nand UO_433 (O_433,N_7694,N_5114);
or UO_434 (O_434,N_7700,N_6217);
xor UO_435 (O_435,N_7332,N_9994);
xor UO_436 (O_436,N_5616,N_6140);
xor UO_437 (O_437,N_9218,N_9409);
and UO_438 (O_438,N_7648,N_5839);
xnor UO_439 (O_439,N_8015,N_9272);
or UO_440 (O_440,N_6755,N_7728);
nor UO_441 (O_441,N_5212,N_7501);
or UO_442 (O_442,N_9276,N_5191);
or UO_443 (O_443,N_7546,N_6928);
nor UO_444 (O_444,N_9394,N_7096);
nand UO_445 (O_445,N_5285,N_8779);
nor UO_446 (O_446,N_9214,N_6191);
nor UO_447 (O_447,N_7107,N_7779);
nand UO_448 (O_448,N_7666,N_7449);
nor UO_449 (O_449,N_5602,N_5715);
and UO_450 (O_450,N_6768,N_8550);
and UO_451 (O_451,N_9869,N_5914);
xnor UO_452 (O_452,N_8338,N_7998);
nor UO_453 (O_453,N_6786,N_7380);
or UO_454 (O_454,N_9116,N_6349);
nand UO_455 (O_455,N_6263,N_9556);
or UO_456 (O_456,N_6116,N_6818);
and UO_457 (O_457,N_7433,N_6351);
xor UO_458 (O_458,N_5718,N_8987);
and UO_459 (O_459,N_9939,N_6262);
xor UO_460 (O_460,N_5504,N_8238);
xnor UO_461 (O_461,N_8050,N_6423);
xnor UO_462 (O_462,N_8568,N_7721);
nor UO_463 (O_463,N_8194,N_7504);
nor UO_464 (O_464,N_8442,N_8315);
or UO_465 (O_465,N_7822,N_5523);
nor UO_466 (O_466,N_6297,N_9336);
and UO_467 (O_467,N_9354,N_8152);
and UO_468 (O_468,N_6245,N_5274);
xor UO_469 (O_469,N_8031,N_5654);
nand UO_470 (O_470,N_8826,N_7462);
or UO_471 (O_471,N_8959,N_6607);
nor UO_472 (O_472,N_9157,N_5159);
or UO_473 (O_473,N_6963,N_9621);
xnor UO_474 (O_474,N_8907,N_6481);
nand UO_475 (O_475,N_5915,N_6398);
or UO_476 (O_476,N_8371,N_9031);
or UO_477 (O_477,N_9926,N_5305);
nand UO_478 (O_478,N_6592,N_9245);
and UO_479 (O_479,N_7993,N_9609);
and UO_480 (O_480,N_9238,N_8287);
nand UO_481 (O_481,N_8737,N_8410);
or UO_482 (O_482,N_9851,N_9632);
nand UO_483 (O_483,N_9797,N_5052);
and UO_484 (O_484,N_9301,N_8311);
and UO_485 (O_485,N_6444,N_5823);
xnor UO_486 (O_486,N_5853,N_6440);
xnor UO_487 (O_487,N_7451,N_7631);
nor UO_488 (O_488,N_9696,N_9785);
or UO_489 (O_489,N_7179,N_7049);
nand UO_490 (O_490,N_9649,N_6425);
xor UO_491 (O_491,N_6216,N_7516);
nor UO_492 (O_492,N_9261,N_7673);
and UO_493 (O_493,N_6189,N_5020);
xor UO_494 (O_494,N_6606,N_8843);
or UO_495 (O_495,N_5551,N_6729);
and UO_496 (O_496,N_5166,N_8815);
xnor UO_497 (O_497,N_6844,N_9202);
xor UO_498 (O_498,N_6862,N_9519);
xnor UO_499 (O_499,N_6213,N_6377);
nor UO_500 (O_500,N_8856,N_7283);
nand UO_501 (O_501,N_9381,N_7600);
xor UO_502 (O_502,N_7173,N_7063);
nand UO_503 (O_503,N_8582,N_8456);
or UO_504 (O_504,N_9887,N_8640);
nor UO_505 (O_505,N_7777,N_9147);
or UO_506 (O_506,N_8349,N_6737);
and UO_507 (O_507,N_5855,N_7896);
xnor UO_508 (O_508,N_5240,N_9139);
xnor UO_509 (O_509,N_5868,N_7797);
nand UO_510 (O_510,N_5135,N_5912);
xor UO_511 (O_511,N_9874,N_9570);
nor UO_512 (O_512,N_9338,N_7640);
or UO_513 (O_513,N_6453,N_5563);
and UO_514 (O_514,N_9075,N_5026);
nand UO_515 (O_515,N_6814,N_5431);
and UO_516 (O_516,N_8180,N_9825);
xor UO_517 (O_517,N_7864,N_6875);
nand UO_518 (O_518,N_6750,N_9735);
nor UO_519 (O_519,N_9217,N_8726);
and UO_520 (O_520,N_9746,N_6564);
and UO_521 (O_521,N_8101,N_7352);
xor UO_522 (O_522,N_8960,N_6942);
or UO_523 (O_523,N_9551,N_5788);
nor UO_524 (O_524,N_8136,N_9915);
or UO_525 (O_525,N_5962,N_8636);
nor UO_526 (O_526,N_8178,N_7040);
and UO_527 (O_527,N_5453,N_8239);
xnor UO_528 (O_528,N_5172,N_6301);
nand UO_529 (O_529,N_9910,N_7758);
and UO_530 (O_530,N_7334,N_5519);
nand UO_531 (O_531,N_6125,N_6162);
nor UO_532 (O_532,N_7382,N_5032);
or UO_533 (O_533,N_5836,N_7705);
xor UO_534 (O_534,N_8483,N_5949);
or UO_535 (O_535,N_5126,N_5267);
or UO_536 (O_536,N_9542,N_7189);
or UO_537 (O_537,N_8514,N_9096);
and UO_538 (O_538,N_8157,N_9955);
nand UO_539 (O_539,N_8849,N_8207);
and UO_540 (O_540,N_5427,N_7961);
nor UO_541 (O_541,N_7152,N_9383);
nor UO_542 (O_542,N_7548,N_8117);
and UO_543 (O_543,N_8078,N_6039);
or UO_544 (O_544,N_7339,N_8033);
or UO_545 (O_545,N_6367,N_9760);
or UO_546 (O_546,N_7570,N_7795);
nand UO_547 (O_547,N_8768,N_6399);
and UO_548 (O_548,N_8139,N_8841);
nor UO_549 (O_549,N_9478,N_6114);
or UO_550 (O_550,N_6575,N_9856);
or UO_551 (O_551,N_6932,N_5844);
nor UO_552 (O_552,N_8396,N_9912);
nor UO_553 (O_553,N_5219,N_5441);
nand UO_554 (O_554,N_5312,N_5664);
or UO_555 (O_555,N_8731,N_7190);
nand UO_556 (O_556,N_5134,N_8590);
nand UO_557 (O_557,N_5575,N_7326);
nor UO_558 (O_558,N_5601,N_5473);
or UO_559 (O_559,N_5012,N_6510);
nand UO_560 (O_560,N_8360,N_6882);
nand UO_561 (O_561,N_7710,N_5584);
xor UO_562 (O_562,N_5357,N_5038);
xnor UO_563 (O_563,N_7727,N_6997);
nor UO_564 (O_564,N_7916,N_7634);
nand UO_565 (O_565,N_7225,N_9921);
nor UO_566 (O_566,N_8921,N_5414);
xnor UO_567 (O_567,N_6663,N_6234);
nand UO_568 (O_568,N_8873,N_8476);
or UO_569 (O_569,N_6461,N_5037);
xor UO_570 (O_570,N_5719,N_7773);
or UO_571 (O_571,N_9088,N_7736);
xnor UO_572 (O_572,N_9932,N_9654);
and UO_573 (O_573,N_5079,N_9389);
or UO_574 (O_574,N_7503,N_9362);
nand UO_575 (O_575,N_8447,N_7985);
nor UO_576 (O_576,N_9422,N_5178);
or UO_577 (O_577,N_5085,N_7881);
nor UO_578 (O_578,N_7701,N_7676);
and UO_579 (O_579,N_8096,N_6077);
nand UO_580 (O_580,N_6252,N_5000);
xnor UO_581 (O_581,N_7538,N_9003);
nor UO_582 (O_582,N_5393,N_7005);
or UO_583 (O_583,N_5565,N_6019);
nor UO_584 (O_584,N_6206,N_6535);
nor UO_585 (O_585,N_8836,N_8982);
nor UO_586 (O_586,N_9624,N_6054);
xnor UO_587 (O_587,N_7374,N_5753);
nor UO_588 (O_588,N_8316,N_7473);
and UO_589 (O_589,N_9271,N_8263);
nor UO_590 (O_590,N_6360,N_6025);
or UO_591 (O_591,N_5746,N_8503);
nor UO_592 (O_592,N_7463,N_6581);
or UO_593 (O_593,N_5301,N_7498);
or UO_594 (O_594,N_7497,N_5727);
nand UO_595 (O_595,N_6764,N_7256);
and UO_596 (O_596,N_6182,N_6013);
and UO_597 (O_597,N_8184,N_5499);
nor UO_598 (O_598,N_7253,N_8696);
and UO_599 (O_599,N_5476,N_7198);
or UO_600 (O_600,N_7135,N_5263);
nand UO_601 (O_601,N_6080,N_7209);
and UO_602 (O_602,N_6104,N_7215);
xnor UO_603 (O_603,N_5774,N_5825);
nor UO_604 (O_604,N_7815,N_9992);
xor UO_605 (O_605,N_8635,N_5130);
xor UO_606 (O_606,N_5789,N_7384);
and UO_607 (O_607,N_6207,N_5062);
nand UO_608 (O_608,N_5929,N_7139);
nand UO_609 (O_609,N_7411,N_6598);
nor UO_610 (O_610,N_6111,N_6157);
and UO_611 (O_611,N_6259,N_5586);
xor UO_612 (O_612,N_8495,N_6345);
nand UO_613 (O_613,N_6359,N_7928);
nor UO_614 (O_614,N_6458,N_5295);
or UO_615 (O_615,N_8173,N_8735);
nor UO_616 (O_616,N_5722,N_8949);
xnor UO_617 (O_617,N_7030,N_7831);
nand UO_618 (O_618,N_9717,N_6148);
xnor UO_619 (O_619,N_5771,N_9640);
or UO_620 (O_620,N_9977,N_5764);
or UO_621 (O_621,N_8872,N_6601);
or UO_622 (O_622,N_7238,N_8868);
nand UO_623 (O_623,N_5375,N_8148);
nor UO_624 (O_624,N_9610,N_8664);
and UO_625 (O_625,N_7665,N_5517);
nor UO_626 (O_626,N_8386,N_6840);
and UO_627 (O_627,N_7786,N_9820);
and UO_628 (O_628,N_9983,N_8596);
and UO_629 (O_629,N_7518,N_9281);
or UO_630 (O_630,N_5508,N_9791);
nor UO_631 (O_631,N_6199,N_8681);
or UO_632 (O_632,N_5101,N_5952);
xnor UO_633 (O_633,N_5086,N_7639);
nand UO_634 (O_634,N_8002,N_5669);
or UO_635 (O_635,N_8853,N_9138);
and UO_636 (O_636,N_9567,N_5148);
and UO_637 (O_637,N_5482,N_6146);
xor UO_638 (O_638,N_9303,N_5193);
nand UO_639 (O_639,N_6910,N_8395);
and UO_640 (O_640,N_5091,N_7685);
and UO_641 (O_641,N_5286,N_6661);
and UO_642 (O_642,N_7965,N_7461);
and UO_643 (O_643,N_8200,N_7992);
and UO_644 (O_644,N_7951,N_9160);
nor UO_645 (O_645,N_7958,N_5646);
nor UO_646 (O_646,N_9150,N_9627);
or UO_647 (O_647,N_5249,N_6117);
nand UO_648 (O_648,N_5544,N_7950);
nor UO_649 (O_649,N_7780,N_7193);
xnor UO_650 (O_650,N_6977,N_6679);
or UO_651 (O_651,N_5509,N_8382);
nor UO_652 (O_652,N_7479,N_8284);
or UO_653 (O_653,N_7115,N_8658);
and UO_654 (O_654,N_8996,N_7926);
and UO_655 (O_655,N_6975,N_9616);
and UO_656 (O_656,N_7983,N_7493);
and UO_657 (O_657,N_6285,N_6758);
and UO_658 (O_658,N_6500,N_8029);
nor UO_659 (O_659,N_7742,N_9530);
or UO_660 (O_660,N_6949,N_5919);
and UO_661 (O_661,N_6323,N_8307);
xor UO_662 (O_662,N_6296,N_6858);
and UO_663 (O_663,N_6277,N_5516);
nor UO_664 (O_664,N_8361,N_7001);
or UO_665 (O_665,N_6976,N_5036);
nor UO_666 (O_666,N_7974,N_7034);
and UO_667 (O_667,N_7796,N_8611);
nor UO_668 (O_668,N_8044,N_8266);
nand UO_669 (O_669,N_8415,N_7686);
nand UO_670 (O_670,N_8132,N_8253);
xnor UO_671 (O_671,N_5495,N_8623);
nand UO_672 (O_672,N_5735,N_7553);
xor UO_673 (O_673,N_9103,N_7947);
nand UO_674 (O_674,N_9589,N_7920);
xnor UO_675 (O_675,N_7606,N_9771);
and UO_676 (O_676,N_9582,N_6585);
and UO_677 (O_677,N_6254,N_5804);
nand UO_678 (O_678,N_6057,N_9439);
and UO_679 (O_679,N_8163,N_7420);
nand UO_680 (O_680,N_9207,N_8822);
nand UO_681 (O_681,N_9605,N_6807);
nand UO_682 (O_682,N_6139,N_6027);
xor UO_683 (O_683,N_6890,N_9574);
xor UO_684 (O_684,N_5104,N_8587);
and UO_685 (O_685,N_8245,N_8291);
and UO_686 (O_686,N_5260,N_5578);
nor UO_687 (O_687,N_9904,N_7706);
and UO_688 (O_688,N_6246,N_5215);
xor UO_689 (O_689,N_8847,N_9192);
xnor UO_690 (O_690,N_7785,N_9140);
nor UO_691 (O_691,N_6935,N_9670);
xor UO_692 (O_692,N_9865,N_8225);
xnor UO_693 (O_693,N_5820,N_7644);
xnor UO_694 (O_694,N_8314,N_8669);
or UO_695 (O_695,N_8420,N_7169);
and UO_696 (O_696,N_8745,N_5082);
and UO_697 (O_697,N_9013,N_9549);
or UO_698 (O_698,N_6003,N_5951);
and UO_699 (O_699,N_5995,N_7973);
and UO_700 (O_700,N_8130,N_9536);
xor UO_701 (O_701,N_6044,N_9241);
nor UO_702 (O_702,N_8268,N_7722);
and UO_703 (O_703,N_5007,N_6708);
nor UO_704 (O_704,N_9288,N_8995);
nand UO_705 (O_705,N_5597,N_9888);
and UO_706 (O_706,N_8516,N_6358);
or UO_707 (O_707,N_8106,N_7026);
nand UO_708 (O_708,N_9755,N_6047);
nand UO_709 (O_709,N_8436,N_7309);
and UO_710 (O_710,N_8344,N_5773);
xor UO_711 (O_711,N_5832,N_5988);
xor UO_712 (O_712,N_7412,N_7752);
xnor UO_713 (O_713,N_7176,N_8604);
and UO_714 (O_714,N_8935,N_9940);
or UO_715 (O_715,N_5781,N_5311);
nor UO_716 (O_716,N_6761,N_9984);
or UO_717 (O_717,N_8676,N_8923);
or UO_718 (O_718,N_6868,N_6061);
xnor UO_719 (O_719,N_6110,N_6280);
and UO_720 (O_720,N_8801,N_9102);
and UO_721 (O_721,N_8113,N_9355);
nand UO_722 (O_722,N_9834,N_9569);
nor UO_723 (O_723,N_9931,N_6937);
or UO_724 (O_724,N_9961,N_5033);
nor UO_725 (O_725,N_9595,N_8484);
nor UO_726 (O_726,N_7556,N_5902);
xnor UO_727 (O_727,N_8188,N_9803);
nor UO_728 (O_728,N_7378,N_9831);
nand UO_729 (O_729,N_6372,N_7599);
or UO_730 (O_730,N_9815,N_7311);
and UO_731 (O_731,N_7731,N_6778);
nor UO_732 (O_732,N_7734,N_9870);
xor UO_733 (O_733,N_7319,N_5537);
and UO_734 (O_734,N_9266,N_9629);
nand UO_735 (O_735,N_8286,N_7855);
nor UO_736 (O_736,N_5073,N_8761);
nand UO_737 (O_737,N_6552,N_9441);
and UO_738 (O_738,N_6070,N_7580);
nand UO_739 (O_739,N_9119,N_6562);
or UO_740 (O_740,N_6068,N_6455);
or UO_741 (O_741,N_8864,N_5078);
xnor UO_742 (O_742,N_6149,N_7242);
nand UO_743 (O_743,N_6636,N_8066);
nor UO_744 (O_744,N_7405,N_9480);
or UO_745 (O_745,N_5153,N_7957);
xor UO_746 (O_746,N_6055,N_6008);
xnor UO_747 (O_747,N_5056,N_6917);
nand UO_748 (O_748,N_7635,N_9848);
and UO_749 (O_749,N_5176,N_6987);
or UO_750 (O_750,N_7680,N_6943);
xnor UO_751 (O_751,N_9533,N_9033);
and UO_752 (O_752,N_9639,N_8288);
xor UO_753 (O_753,N_6266,N_9695);
and UO_754 (O_754,N_6286,N_6496);
nor UO_755 (O_755,N_7655,N_8081);
or UO_756 (O_756,N_6075,N_8943);
nor UO_757 (O_757,N_8906,N_9485);
nand UO_758 (O_758,N_7628,N_8687);
xnor UO_759 (O_759,N_5110,N_9177);
xor UO_760 (O_760,N_5603,N_6409);
xnor UO_761 (O_761,N_5745,N_8128);
or UO_762 (O_762,N_5195,N_7905);
or UO_763 (O_763,N_6951,N_6159);
xnor UO_764 (O_764,N_7475,N_9531);
xor UO_765 (O_765,N_9715,N_9342);
xor UO_766 (O_766,N_9920,N_8911);
nor UO_767 (O_767,N_9270,N_5845);
xor UO_768 (O_768,N_8962,N_6401);
or UO_769 (O_769,N_7290,N_5829);
xor UO_770 (O_770,N_9239,N_6493);
or UO_771 (O_771,N_7813,N_9631);
xor UO_772 (O_772,N_7279,N_9975);
nor UO_773 (O_773,N_5506,N_5145);
nor UO_774 (O_774,N_7110,N_8355);
and UO_775 (O_775,N_8616,N_5887);
nand UO_776 (O_776,N_6329,N_9460);
nand UO_777 (O_777,N_8915,N_5122);
and UO_778 (O_778,N_9314,N_9390);
nand UO_779 (O_779,N_7330,N_9970);
and UO_780 (O_780,N_7293,N_5941);
nor UO_781 (O_781,N_7003,N_7681);
or UO_782 (O_782,N_5761,N_8455);
or UO_783 (O_783,N_9429,N_9969);
xor UO_784 (O_784,N_8972,N_8759);
and UO_785 (O_785,N_7366,N_7608);
nor UO_786 (O_786,N_8448,N_7289);
nor UO_787 (O_787,N_8926,N_8369);
nand UO_788 (O_788,N_6017,N_6222);
nand UO_789 (O_789,N_9507,N_5553);
nand UO_790 (O_790,N_6188,N_8816);
nand UO_791 (O_791,N_9804,N_6655);
nor UO_792 (O_792,N_6876,N_5980);
nand UO_793 (O_793,N_6861,N_9564);
and UO_794 (O_794,N_9042,N_8129);
or UO_795 (O_795,N_6186,N_8861);
nand UO_796 (O_796,N_9693,N_7387);
and UO_797 (O_797,N_7834,N_8684);
nor UO_798 (O_798,N_6669,N_9171);
nand UO_799 (O_799,N_6355,N_8179);
or UO_800 (O_800,N_8914,N_9502);
nand UO_801 (O_801,N_5802,N_6035);
xnor UO_802 (O_802,N_8845,N_7167);
or UO_803 (O_803,N_8322,N_7358);
or UO_804 (O_804,N_5027,N_8649);
nand UO_805 (O_805,N_8256,N_9280);
and UO_806 (O_806,N_9080,N_8499);
nor UO_807 (O_807,N_8769,N_5979);
nor UO_808 (O_808,N_8897,N_8003);
or UO_809 (O_809,N_5333,N_8479);
or UO_810 (O_810,N_6806,N_8485);
nand UO_811 (O_811,N_9764,N_8919);
nor UO_812 (O_812,N_8585,N_8517);
nand UO_813 (O_813,N_8494,N_8782);
and UO_814 (O_814,N_9068,N_9713);
or UO_815 (O_815,N_6537,N_5533);
or UO_816 (O_816,N_8474,N_7170);
and UO_817 (O_817,N_9772,N_9908);
xnor UO_818 (O_818,N_6726,N_6549);
or UO_819 (O_819,N_6781,N_9635);
nand UO_820 (O_820,N_9135,N_6236);
and UO_821 (O_821,N_7381,N_5777);
nor UO_822 (O_822,N_5505,N_6049);
nor UO_823 (O_823,N_8857,N_8384);
nand UO_824 (O_824,N_6531,N_6397);
nor UO_825 (O_825,N_9573,N_9557);
nand UO_826 (O_826,N_9945,N_8655);
xor UO_827 (O_827,N_6832,N_5115);
nor UO_828 (O_828,N_7566,N_7914);
or UO_829 (O_829,N_6738,N_9193);
xor UO_830 (O_830,N_8505,N_5181);
or UO_831 (O_831,N_5423,N_7486);
nor UO_832 (O_832,N_6743,N_6414);
nand UO_833 (O_833,N_7424,N_9334);
nand UO_834 (O_834,N_9671,N_5354);
xor UO_835 (O_835,N_6704,N_8804);
xnor UO_836 (O_836,N_7104,N_5298);
and UO_837 (O_837,N_7792,N_6543);
and UO_838 (O_838,N_5679,N_8538);
nor UO_839 (O_839,N_6805,N_6992);
xor UO_840 (O_840,N_9846,N_5030);
or UO_841 (O_841,N_9614,N_6130);
xnor UO_842 (O_842,N_6647,N_5389);
and UO_843 (O_843,N_9273,N_9324);
and UO_844 (O_844,N_8531,N_8540);
xor UO_845 (O_845,N_6198,N_9993);
xnor UO_846 (O_846,N_6833,N_9873);
nand UO_847 (O_847,N_8628,N_6909);
and UO_848 (O_848,N_9306,N_8082);
nor UO_849 (O_849,N_5131,N_8166);
nand UO_850 (O_850,N_6097,N_8205);
and UO_851 (O_851,N_8045,N_9943);
and UO_852 (O_852,N_6109,N_7915);
xnor UO_853 (O_853,N_5545,N_7067);
nand UO_854 (O_854,N_9368,N_5315);
and UO_855 (O_855,N_5306,N_5350);
nand UO_856 (O_856,N_9544,N_5750);
nor UO_857 (O_857,N_6863,N_5214);
or UO_858 (O_858,N_7552,N_5009);
nor UO_859 (O_859,N_7499,N_5943);
nor UO_860 (O_860,N_7717,N_8563);
xor UO_861 (O_861,N_8511,N_9391);
and UO_862 (O_862,N_9151,N_5502);
xor UO_863 (O_863,N_9449,N_7849);
xnor UO_864 (O_864,N_9437,N_8244);
xor UO_865 (O_865,N_9365,N_6676);
nand UO_866 (O_866,N_6554,N_7949);
and UO_867 (O_867,N_9547,N_9898);
xor UO_868 (O_868,N_6567,N_7614);
nor UO_869 (O_869,N_9794,N_6364);
or UO_870 (O_870,N_5179,N_5364);
or UO_871 (O_871,N_8783,N_6041);
nor UO_872 (O_872,N_6167,N_9517);
or UO_873 (O_873,N_8837,N_9251);
nor UO_874 (O_874,N_7341,N_5273);
nor UO_875 (O_875,N_9742,N_9066);
xor UO_876 (O_876,N_8162,N_8312);
nand UO_877 (O_877,N_7856,N_6258);
nor UO_878 (O_878,N_8013,N_5786);
and UO_879 (O_879,N_9369,N_8892);
and UO_880 (O_880,N_6279,N_6757);
or UO_881 (O_881,N_6292,N_6211);
or UO_882 (O_882,N_9828,N_5898);
and UO_883 (O_883,N_8341,N_7851);
and UO_884 (O_884,N_5933,N_9000);
xor UO_885 (O_885,N_5152,N_8913);
or UO_886 (O_886,N_7278,N_6929);
nand UO_887 (O_887,N_5705,N_8527);
xnor UO_888 (O_888,N_9406,N_8834);
nand UO_889 (O_889,N_6185,N_8076);
xnor UO_890 (O_890,N_8325,N_9469);
and UO_891 (O_891,N_9653,N_6642);
nand UO_892 (O_892,N_6171,N_5330);
or UO_893 (O_893,N_7769,N_5838);
nand UO_894 (O_894,N_9698,N_6042);
or UO_895 (O_895,N_6924,N_5592);
and UO_896 (O_896,N_9002,N_8647);
xor UO_897 (O_897,N_6860,N_9094);
nor UO_898 (O_898,N_5570,N_5634);
nand UO_899 (O_899,N_6719,N_5906);
nand UO_900 (O_900,N_9476,N_6160);
or UO_901 (O_901,N_9952,N_7455);
xor UO_902 (O_902,N_8007,N_7900);
xor UO_903 (O_903,N_7678,N_5368);
nand UO_904 (O_904,N_8592,N_5612);
xnor UO_905 (O_905,N_6956,N_6640);
and UO_906 (O_906,N_9219,N_5136);
and UO_907 (O_907,N_9400,N_8501);
nor UO_908 (O_908,N_8927,N_7195);
nand UO_909 (O_909,N_7019,N_9360);
or UO_910 (O_910,N_7724,N_7321);
nand UO_911 (O_911,N_5967,N_7365);
nor UO_912 (O_912,N_6273,N_9782);
nor UO_913 (O_913,N_5108,N_5899);
xor UO_914 (O_914,N_5946,N_6001);
or UO_915 (O_915,N_6599,N_6767);
xnor UO_916 (O_916,N_5757,N_5944);
nand UO_917 (O_917,N_7071,N_7082);
and UO_918 (O_918,N_7260,N_7853);
nand UO_919 (O_919,N_9754,N_5672);
and UO_920 (O_920,N_9586,N_7373);
and UO_921 (O_921,N_9229,N_5479);
nand UO_922 (O_922,N_9661,N_5359);
nor UO_923 (O_923,N_5271,N_8881);
and UO_924 (O_924,N_9879,N_7607);
nor UO_925 (O_925,N_5139,N_9117);
and UO_926 (O_926,N_9647,N_6920);
nand UO_927 (O_927,N_5335,N_8762);
nand UO_928 (O_928,N_9630,N_5628);
and UO_929 (O_929,N_9446,N_8126);
nor UO_930 (O_930,N_7418,N_8174);
or UO_931 (O_931,N_5503,N_8547);
and UO_932 (O_932,N_5560,N_8282);
and UO_933 (O_933,N_5916,N_9149);
xnor UO_934 (O_934,N_7643,N_5317);
nand UO_935 (O_935,N_8171,N_6827);
and UO_936 (O_936,N_8755,N_6888);
xnor UO_937 (O_937,N_6325,N_6846);
nand UO_938 (O_938,N_9953,N_5486);
or UO_939 (O_939,N_5429,N_9816);
nand UO_940 (O_940,N_8738,N_6005);
nand UO_941 (O_941,N_5034,N_8791);
nor UO_942 (O_942,N_8100,N_7756);
nor UO_943 (O_943,N_8662,N_8446);
nand UO_944 (O_944,N_5875,N_7511);
xor UO_945 (O_945,N_7624,N_7862);
or UO_946 (O_946,N_7331,N_8457);
nand UO_947 (O_947,N_6571,N_7204);
or UO_948 (O_948,N_7346,N_7547);
or UO_949 (O_949,N_8231,N_8863);
nand UO_950 (O_950,N_7824,N_6079);
or UO_951 (O_951,N_9951,N_8170);
xnor UO_952 (O_952,N_7296,N_6420);
and UO_953 (O_953,N_5324,N_9550);
or UO_954 (O_954,N_5358,N_9431);
xnor UO_955 (O_955,N_9705,N_5233);
nor UO_956 (O_956,N_8380,N_8426);
and UO_957 (O_957,N_7425,N_9864);
and UO_958 (O_958,N_5651,N_7651);
xor UO_959 (O_959,N_7812,N_7997);
xor UO_960 (O_960,N_5432,N_7129);
xnor UO_961 (O_961,N_5511,N_5883);
nand UO_962 (O_962,N_8928,N_8744);
nand UO_963 (O_963,N_9889,N_7897);
or UO_964 (O_964,N_6475,N_5873);
and UO_965 (O_965,N_6682,N_5783);
nand UO_966 (O_966,N_6871,N_9960);
xnor UO_967 (O_967,N_6995,N_7817);
nand UO_968 (O_968,N_6299,N_7869);
nor UO_969 (O_969,N_9402,N_9704);
and UO_970 (O_970,N_5459,N_5937);
and UO_971 (O_971,N_5573,N_9677);
nor UO_972 (O_972,N_9877,N_5314);
nor UO_973 (O_973,N_7085,N_5733);
nor UO_974 (O_974,N_8111,N_6651);
xor UO_975 (O_975,N_9728,N_7572);
and UO_976 (O_976,N_6094,N_9108);
nor UO_977 (O_977,N_8773,N_9579);
nand UO_978 (O_978,N_7297,N_9430);
and UO_979 (O_979,N_5019,N_8883);
and UO_980 (O_980,N_6907,N_8417);
nand UO_981 (O_981,N_9134,N_8992);
xor UO_982 (O_982,N_6683,N_9071);
or UO_983 (O_983,N_9053,N_9329);
and UO_984 (O_984,N_7761,N_5035);
or UO_985 (O_985,N_9319,N_9292);
or UO_986 (O_986,N_6066,N_8222);
nand UO_987 (O_987,N_8149,N_8175);
and UO_988 (O_988,N_8724,N_7652);
or UO_989 (O_989,N_5811,N_5284);
nor UO_990 (O_990,N_7452,N_8792);
nor UO_991 (O_991,N_7591,N_5737);
nor UO_992 (O_992,N_9268,N_7976);
nand UO_993 (O_993,N_7800,N_9759);
xnor UO_994 (O_994,N_8869,N_7216);
and UO_995 (O_995,N_9857,N_5893);
nor UO_996 (O_996,N_7118,N_9461);
and UO_997 (O_997,N_7793,N_9540);
xnor UO_998 (O_998,N_7952,N_5144);
xor UO_999 (O_999,N_9645,N_9162);
nor UO_1000 (O_1000,N_5296,N_5749);
xnor UO_1001 (O_1001,N_6416,N_8973);
xor UO_1002 (O_1002,N_5420,N_8812);
and UO_1003 (O_1003,N_8966,N_8621);
xor UO_1004 (O_1004,N_7691,N_5186);
or UO_1005 (O_1005,N_9957,N_8434);
xnor UO_1006 (O_1006,N_8102,N_9225);
and UO_1007 (O_1007,N_6454,N_7064);
and UO_1008 (O_1008,N_9049,N_6614);
nand UO_1009 (O_1009,N_7153,N_7055);
nand UO_1010 (O_1010,N_8888,N_7595);
and UO_1011 (O_1011,N_5963,N_5044);
and UO_1012 (O_1012,N_8802,N_6887);
and UO_1013 (O_1013,N_7932,N_6295);
and UO_1014 (O_1014,N_5058,N_6161);
and UO_1015 (O_1015,N_9132,N_7432);
nor UO_1016 (O_1016,N_8838,N_6120);
or UO_1017 (O_1017,N_5590,N_8364);
and UO_1018 (O_1018,N_5629,N_6142);
xor UO_1019 (O_1019,N_8435,N_9305);
nor UO_1020 (O_1020,N_8707,N_6596);
and UO_1021 (O_1021,N_5571,N_8813);
xor UO_1022 (O_1022,N_9364,N_7629);
xor UO_1023 (O_1023,N_5627,N_7298);
or UO_1024 (O_1024,N_7568,N_6587);
and UO_1025 (O_1025,N_9486,N_5677);
and UO_1026 (O_1026,N_5613,N_6002);
xnor UO_1027 (O_1027,N_7645,N_5626);
or UO_1028 (O_1028,N_6107,N_9026);
and UO_1029 (O_1029,N_8425,N_8835);
nor UO_1030 (O_1030,N_8855,N_7436);
xor UO_1031 (O_1031,N_7270,N_8867);
nand UO_1032 (O_1032,N_9318,N_9702);
nor UO_1033 (O_1033,N_7579,N_8910);
and UO_1034 (O_1034,N_5095,N_5167);
xor UO_1035 (O_1035,N_8359,N_9934);
xnor UO_1036 (O_1036,N_8970,N_6930);
and UO_1037 (O_1037,N_8504,N_5074);
xor UO_1038 (O_1038,N_7852,N_6487);
nand UO_1039 (O_1039,N_9861,N_7763);
xor UO_1040 (O_1040,N_5692,N_5418);
nor UO_1041 (O_1041,N_7515,N_9473);
xor UO_1042 (O_1042,N_5226,N_5779);
nor UO_1043 (O_1043,N_6612,N_9532);
xor UO_1044 (O_1044,N_9426,N_8831);
or UO_1045 (O_1045,N_6633,N_7117);
xnor UO_1046 (O_1046,N_7549,N_9376);
nor UO_1047 (O_1047,N_7340,N_9274);
nand UO_1048 (O_1048,N_6513,N_6427);
and UO_1049 (O_1049,N_6204,N_5894);
and UO_1050 (O_1050,N_6388,N_8510);
nand UO_1051 (O_1051,N_6819,N_8025);
xnor UO_1052 (O_1052,N_7480,N_7832);
or UO_1053 (O_1053,N_8345,N_8140);
xor UO_1054 (O_1054,N_8922,N_9024);
xnor UO_1055 (O_1055,N_8042,N_9974);
and UO_1056 (O_1056,N_5986,N_8610);
or UO_1057 (O_1057,N_6479,N_5341);
nand UO_1058 (O_1058,N_9577,N_9454);
nand UO_1059 (O_1059,N_7471,N_9944);
and UO_1060 (O_1060,N_9427,N_5667);
or UO_1061 (O_1061,N_7228,N_7968);
nand UO_1062 (O_1062,N_9447,N_9414);
xor UO_1063 (O_1063,N_7142,N_9516);
xnor UO_1064 (O_1064,N_8705,N_5959);
and UO_1065 (O_1065,N_9346,N_7702);
nor UO_1066 (O_1066,N_7288,N_9142);
and UO_1067 (O_1067,N_5235,N_5611);
xnor UO_1068 (O_1068,N_8518,N_7094);
xnor UO_1069 (O_1069,N_8467,N_5255);
xnor UO_1070 (O_1070,N_7929,N_8400);
nand UO_1071 (O_1071,N_6283,N_5089);
nand UO_1072 (O_1072,N_5048,N_7069);
and UO_1073 (O_1073,N_6884,N_7650);
and UO_1074 (O_1074,N_5365,N_9981);
and UO_1075 (O_1075,N_5327,N_8480);
or UO_1076 (O_1076,N_8945,N_6328);
or UO_1077 (O_1077,N_7161,N_5161);
nand UO_1078 (O_1078,N_6556,N_5814);
nor UO_1079 (O_1079,N_9465,N_5289);
nand UO_1080 (O_1080,N_6515,N_8427);
xor UO_1081 (O_1081,N_5281,N_5480);
nand UO_1082 (O_1082,N_8946,N_6522);
nor UO_1083 (O_1083,N_5413,N_8580);
nand UO_1084 (O_1084,N_8879,N_7000);
nand UO_1085 (O_1085,N_7004,N_5610);
and UO_1086 (O_1086,N_7924,N_9133);
nor UO_1087 (O_1087,N_9652,N_6506);
xnor UO_1088 (O_1088,N_8319,N_6550);
nand UO_1089 (O_1089,N_6775,N_5948);
xor UO_1090 (O_1090,N_5300,N_8230);
and UO_1091 (O_1091,N_6072,N_7638);
and UO_1092 (O_1092,N_5061,N_8589);
and UO_1093 (O_1093,N_5554,N_5320);
nor UO_1094 (O_1094,N_9724,N_8564);
nand UO_1095 (O_1095,N_9325,N_7898);
xor UO_1096 (O_1096,N_9786,N_8874);
and UO_1097 (O_1097,N_5810,N_6378);
nand UO_1098 (O_1098,N_8432,N_8561);
and UO_1099 (O_1099,N_6795,N_7362);
nand UO_1100 (O_1100,N_8227,N_9333);
nor UO_1101 (O_1101,N_7224,N_8090);
nand UO_1102 (O_1102,N_9012,N_7187);
nor UO_1103 (O_1103,N_6306,N_5003);
and UO_1104 (O_1104,N_6594,N_6696);
nor UO_1105 (O_1105,N_6314,N_5299);
nor UO_1106 (O_1106,N_7310,N_7286);
nand UO_1107 (O_1107,N_6417,N_5111);
or UO_1108 (O_1108,N_6983,N_5752);
and UO_1109 (O_1109,N_5985,N_6348);
xor UO_1110 (O_1110,N_6268,N_6342);
and UO_1111 (O_1111,N_5097,N_8584);
or UO_1112 (O_1112,N_8572,N_7841);
or UO_1113 (O_1113,N_9257,N_9836);
or UO_1114 (O_1114,N_9204,N_6387);
or UO_1115 (O_1115,N_7140,N_9179);
or UO_1116 (O_1116,N_8009,N_5577);
nand UO_1117 (O_1117,N_6353,N_9323);
xnor UO_1118 (O_1118,N_8700,N_6584);
and UO_1119 (O_1119,N_5690,N_6291);
or UO_1120 (O_1120,N_8279,N_7830);
nor UO_1121 (O_1121,N_7723,N_9248);
xnor UO_1122 (O_1122,N_5433,N_9300);
nand UO_1123 (O_1123,N_9173,N_6699);
nor UO_1124 (O_1124,N_6449,N_8182);
or UO_1125 (O_1125,N_6974,N_6093);
nor UO_1126 (O_1126,N_6756,N_9999);
xnor UO_1127 (O_1127,N_8285,N_5238);
or UO_1128 (O_1128,N_7100,N_7143);
and UO_1129 (O_1129,N_5355,N_6831);
nand UO_1130 (O_1130,N_9817,N_5717);
or UO_1131 (O_1131,N_7156,N_6318);
and UO_1132 (O_1132,N_6443,N_5371);
or UO_1133 (O_1133,N_9628,N_6434);
or UO_1134 (O_1134,N_9829,N_9143);
xor UO_1135 (O_1135,N_9996,N_5469);
and UO_1136 (O_1136,N_6386,N_8741);
nand UO_1137 (O_1137,N_9105,N_7214);
nand UO_1138 (O_1138,N_5092,N_8583);
and UO_1139 (O_1139,N_8846,N_5854);
nor UO_1140 (O_1140,N_5316,N_6373);
and UO_1141 (O_1141,N_9894,N_5840);
xor UO_1142 (O_1142,N_7804,N_5201);
or UO_1143 (O_1143,N_6528,N_7370);
nand UO_1144 (O_1144,N_6864,N_5824);
xor UO_1145 (O_1145,N_5529,N_7922);
and UO_1146 (O_1146,N_8968,N_7258);
nand UO_1147 (O_1147,N_7371,N_9237);
nand UO_1148 (O_1148,N_8151,N_8603);
and UO_1149 (O_1149,N_6218,N_6267);
and UO_1150 (O_1150,N_5978,N_5512);
xor UO_1151 (O_1151,N_6036,N_6131);
or UO_1152 (O_1152,N_9169,N_6270);
nor UO_1153 (O_1153,N_5961,N_6989);
xnor UO_1154 (O_1154,N_5361,N_9467);
or UO_1155 (O_1155,N_7084,N_8627);
nand UO_1156 (O_1156,N_9809,N_6052);
and UO_1157 (O_1157,N_9197,N_8870);
xor UO_1158 (O_1158,N_6934,N_7699);
nand UO_1159 (O_1159,N_6244,N_8588);
or UO_1160 (O_1160,N_7659,N_6424);
xnor UO_1161 (O_1161,N_8743,N_5276);
nand UO_1162 (O_1162,N_6485,N_9294);
nand UO_1163 (O_1163,N_8720,N_8296);
and UO_1164 (O_1164,N_9534,N_7658);
nor UO_1165 (O_1165,N_7725,N_9853);
or UO_1166 (O_1166,N_8051,N_6489);
nand UO_1167 (O_1167,N_8213,N_5288);
xor UO_1168 (O_1168,N_6577,N_8795);
xor UO_1169 (O_1169,N_9634,N_5721);
or UO_1170 (O_1170,N_8001,N_5224);
xnor UO_1171 (O_1171,N_6852,N_6834);
or UO_1172 (O_1172,N_5068,N_5911);
xnor UO_1173 (O_1173,N_8389,N_5817);
nand UO_1174 (O_1174,N_7911,N_7939);
xnor UO_1175 (O_1175,N_6331,N_5174);
nand UO_1176 (O_1176,N_5326,N_5780);
or UO_1177 (O_1177,N_7888,N_7963);
or UO_1178 (O_1178,N_5342,N_9442);
nor UO_1179 (O_1179,N_5815,N_7910);
or UO_1180 (O_1180,N_8950,N_8292);
nor UO_1181 (O_1181,N_8065,N_6700);
and UO_1182 (O_1182,N_8709,N_6684);
nor UO_1183 (O_1183,N_5856,N_9126);
or UO_1184 (O_1184,N_5741,N_6100);
nor UO_1185 (O_1185,N_7519,N_8811);
or UO_1186 (O_1186,N_8127,N_8633);
and UO_1187 (O_1187,N_6486,N_6802);
and UO_1188 (O_1188,N_9922,N_7975);
nor UO_1189 (O_1189,N_6732,N_6134);
xnor UO_1190 (O_1190,N_7512,N_9382);
nand UO_1191 (O_1191,N_8321,N_9811);
and UO_1192 (O_1192,N_6124,N_9278);
nor UO_1193 (O_1193,N_8814,N_5120);
xnor UO_1194 (O_1194,N_5225,N_6442);
nor UO_1195 (O_1195,N_9923,N_5606);
nor UO_1196 (O_1196,N_9475,N_5264);
xnor UO_1197 (O_1197,N_7233,N_5100);
nor UO_1198 (O_1198,N_6678,N_6183);
and UO_1199 (O_1199,N_7377,N_8778);
xor UO_1200 (O_1200,N_8408,N_9379);
xnor UO_1201 (O_1201,N_7790,N_7174);
xor UO_1202 (O_1202,N_6916,N_5531);
xnor UO_1203 (O_1203,N_8221,N_9736);
or UO_1204 (O_1204,N_6098,N_9885);
and UO_1205 (O_1205,N_7206,N_7772);
xor UO_1206 (O_1206,N_6602,N_9343);
nor UO_1207 (O_1207,N_7750,N_5905);
nand UO_1208 (O_1208,N_6069,N_6541);
nand UO_1209 (O_1209,N_7509,N_9555);
xnor UO_1210 (O_1210,N_5541,N_8125);
or UO_1211 (O_1211,N_9578,N_5292);
and UO_1212 (O_1212,N_9312,N_8020);
xor UO_1213 (O_1213,N_8115,N_8566);
xnor UO_1214 (O_1214,N_5747,N_8350);
nand UO_1215 (O_1215,N_6219,N_7646);
nand UO_1216 (O_1216,N_7764,N_8771);
and UO_1217 (O_1217,N_5546,N_6445);
and UO_1218 (O_1218,N_6302,N_9247);
xnor UO_1219 (O_1219,N_9059,N_5572);
and UO_1220 (O_1220,N_8452,N_5362);
and UO_1221 (O_1221,N_6533,N_7809);
nand UO_1222 (O_1222,N_9598,N_6274);
or UO_1223 (O_1223,N_9425,N_7490);
nor UO_1224 (O_1224,N_8609,N_5989);
or UO_1225 (O_1225,N_7581,N_6759);
xor UO_1226 (O_1226,N_5955,N_7138);
xnor UO_1227 (O_1227,N_6923,N_7121);
or UO_1228 (O_1228,N_7457,N_7754);
and UO_1229 (O_1229,N_9566,N_5888);
and UO_1230 (O_1230,N_6803,N_5376);
or UO_1231 (O_1231,N_5754,N_6304);
or UO_1232 (O_1232,N_5594,N_9919);
nor UO_1233 (O_1233,N_8237,N_7837);
xor UO_1234 (O_1234,N_7859,N_7741);
nor UO_1235 (O_1235,N_8310,N_6558);
nand UO_1236 (O_1236,N_8620,N_6096);
and UO_1237 (O_1237,N_5084,N_8466);
or UO_1238 (O_1238,N_6664,N_5470);
or UO_1239 (O_1239,N_5147,N_9814);
nand UO_1240 (O_1240,N_7672,N_5399);
nand UO_1241 (O_1241,N_6354,N_9587);
and UO_1242 (O_1242,N_5417,N_5707);
xor UO_1243 (O_1243,N_9249,N_9321);
xnor UO_1244 (O_1244,N_7299,N_7836);
nor UO_1245 (O_1245,N_9172,N_6879);
xnor UO_1246 (O_1246,N_8776,N_8193);
and UO_1247 (O_1247,N_7399,N_7303);
or UO_1248 (O_1248,N_6894,N_7192);
nor UO_1249 (O_1249,N_5784,N_5609);
nand UO_1250 (O_1250,N_9110,N_5387);
nand UO_1251 (O_1251,N_6248,N_6645);
xor UO_1252 (O_1252,N_5960,N_7415);
nand UO_1253 (O_1253,N_5514,N_6812);
and UO_1254 (O_1254,N_8320,N_9020);
nand UO_1255 (O_1255,N_6504,N_5338);
nor UO_1256 (O_1256,N_9716,N_6648);
and UO_1257 (O_1257,N_5332,N_5670);
or UO_1258 (O_1258,N_9935,N_5904);
and UO_1259 (O_1259,N_6711,N_8819);
nor UO_1260 (O_1260,N_9656,N_9122);
xnor UO_1261 (O_1261,N_7087,N_6893);
or UO_1262 (O_1262,N_6611,N_6463);
nor UO_1263 (O_1263,N_7738,N_9308);
or UO_1264 (O_1264,N_9452,N_7347);
or UO_1265 (O_1265,N_9311,N_8866);
nand UO_1266 (O_1266,N_5442,N_8750);
nand UO_1267 (O_1267,N_5790,N_9648);
and UO_1268 (O_1268,N_8016,N_8513);
or UO_1269 (O_1269,N_6591,N_5259);
nor UO_1270 (O_1270,N_5994,N_5953);
nor UO_1271 (O_1271,N_5760,N_8600);
xnor UO_1272 (O_1272,N_7392,N_6901);
and UO_1273 (O_1273,N_9412,N_8218);
nor UO_1274 (O_1274,N_8443,N_9571);
or UO_1275 (O_1275,N_7861,N_6499);
xnor UO_1276 (O_1276,N_8070,N_9037);
nor UO_1277 (O_1277,N_7041,N_9155);
nor UO_1278 (O_1278,N_8061,N_7390);
or UO_1279 (O_1279,N_7980,N_7393);
or UO_1280 (O_1280,N_7799,N_9211);
and UO_1281 (O_1281,N_6484,N_9076);
or UO_1282 (O_1282,N_6822,N_6084);
nand UO_1283 (O_1283,N_5957,N_6649);
nor UO_1284 (O_1284,N_9048,N_7202);
nand UO_1285 (O_1285,N_9165,N_6026);
nor UO_1286 (O_1286,N_5057,N_7781);
xor UO_1287 (O_1287,N_7182,N_5892);
and UO_1288 (O_1288,N_5256,N_8715);
nand UO_1289 (O_1289,N_9298,N_7625);
nor UO_1290 (O_1290,N_8375,N_8850);
nor UO_1291 (O_1291,N_5155,N_8397);
nor UO_1292 (O_1292,N_6836,N_9594);
nor UO_1293 (O_1293,N_8248,N_6395);
xor UO_1294 (O_1294,N_7923,N_9838);
nor UO_1295 (O_1295,N_9184,N_7664);
nor UO_1296 (O_1296,N_9777,N_7329);
or UO_1297 (O_1297,N_5550,N_9500);
xnor UO_1298 (O_1298,N_5500,N_9331);
and UO_1299 (O_1299,N_7843,N_8767);
nand UO_1300 (O_1300,N_7180,N_9067);
nor UO_1301 (O_1301,N_6752,N_9843);
xor UO_1302 (O_1302,N_8441,N_5791);
xor UO_1303 (O_1303,N_8014,N_8728);
xnor UO_1304 (O_1304,N_8356,N_9156);
nor UO_1305 (O_1305,N_8971,N_6731);
and UO_1306 (O_1306,N_5515,N_7960);
xnor UO_1307 (O_1307,N_8354,N_7398);
xnor UO_1308 (O_1308,N_9588,N_6451);
nand UO_1309 (O_1309,N_6579,N_7936);
xor UO_1310 (O_1310,N_6958,N_9118);
nand UO_1311 (O_1311,N_9604,N_6144);
and UO_1312 (O_1312,N_5827,N_5658);
xnor UO_1313 (O_1313,N_8252,N_9768);
and UO_1314 (O_1314,N_7402,N_6282);
nand UO_1315 (O_1315,N_9339,N_8421);
xnor UO_1316 (O_1316,N_7369,N_6872);
nor UO_1317 (O_1317,N_6889,N_9722);
and UO_1318 (O_1318,N_8764,N_8492);
nand UO_1319 (O_1319,N_5762,N_7842);
nor UO_1320 (O_1320,N_8146,N_7262);
nand UO_1321 (O_1321,N_7301,N_7083);
nand UO_1322 (O_1322,N_8073,N_6817);
or UO_1323 (O_1323,N_9976,N_9388);
xnor UO_1324 (O_1324,N_5635,N_9659);
nand UO_1325 (O_1325,N_8405,N_6540);
nand UO_1326 (O_1326,N_7481,N_9403);
nor UO_1327 (O_1327,N_8377,N_9607);
xor UO_1328 (O_1328,N_8858,N_8549);
nand UO_1329 (O_1329,N_5767,N_7379);
and UO_1330 (O_1330,N_7766,N_8095);
nor UO_1331 (O_1331,N_6091,N_7364);
or UO_1332 (O_1332,N_7272,N_7130);
nand UO_1333 (O_1333,N_9537,N_8925);
and UO_1334 (O_1334,N_9526,N_7821);
xnor UO_1335 (O_1335,N_8535,N_6529);
xnor UO_1336 (O_1336,N_8594,N_9749);
or UO_1337 (O_1337,N_9483,N_9185);
nor UO_1338 (O_1338,N_6979,N_5706);
nand UO_1339 (O_1339,N_9618,N_9194);
or UO_1340 (O_1340,N_8860,N_9929);
and UO_1341 (O_1341,N_7406,N_6641);
xnor UO_1342 (O_1342,N_7917,N_5416);
xor UO_1343 (O_1343,N_5261,N_8035);
nand UO_1344 (O_1344,N_8677,N_6600);
nor UO_1345 (O_1345,N_6948,N_7212);
and UO_1346 (O_1346,N_5313,N_5487);
nand UO_1347 (O_1347,N_6369,N_6919);
or UO_1348 (O_1348,N_5936,N_5016);
xnor UO_1349 (O_1349,N_7586,N_9038);
nor UO_1350 (O_1350,N_6940,N_9458);
nor UO_1351 (O_1351,N_7531,N_8409);
nand UO_1352 (O_1352,N_8204,N_5076);
and UO_1353 (O_1353,N_5198,N_9373);
and UO_1354 (O_1354,N_9827,N_7906);
nor UO_1355 (O_1355,N_8463,N_7611);
and UO_1356 (O_1356,N_5623,N_6490);
nor UO_1357 (O_1357,N_9603,N_7076);
or UO_1358 (O_1358,N_7767,N_8470);
or UO_1359 (O_1359,N_8097,N_8639);
nor UO_1360 (O_1360,N_5621,N_6152);
and UO_1361 (O_1361,N_5974,N_5896);
xnor UO_1362 (O_1362,N_9775,N_6874);
and UO_1363 (O_1363,N_7927,N_5826);
xnor UO_1364 (O_1364,N_5232,N_5328);
and UO_1365 (O_1365,N_6374,N_7814);
xnor UO_1366 (O_1366,N_6867,N_8757);
and UO_1367 (O_1367,N_8209,N_5655);
or UO_1368 (O_1368,N_6899,N_8261);
or UO_1369 (O_1369,N_5337,N_8093);
xnor UO_1370 (O_1370,N_5755,N_6411);
or UO_1371 (O_1371,N_9087,N_6467);
and UO_1372 (O_1372,N_6993,N_7328);
nor UO_1373 (O_1373,N_7091,N_7895);
or UO_1374 (O_1374,N_8586,N_8464);
and UO_1375 (O_1375,N_9148,N_8023);
nor UO_1376 (O_1376,N_7848,N_5370);
xor UO_1377 (O_1377,N_5540,N_9050);
xor UO_1378 (O_1378,N_9515,N_8089);
nor UO_1379 (O_1379,N_7709,N_7320);
or UO_1380 (O_1380,N_6081,N_7261);
and UO_1381 (O_1381,N_9361,N_8251);
or UO_1382 (O_1382,N_8471,N_7941);
nor UO_1383 (O_1383,N_5437,N_5977);
nor UO_1384 (O_1384,N_8608,N_6961);
or UO_1385 (O_1385,N_8920,N_6136);
nor UO_1386 (O_1386,N_5461,N_9784);
nor UO_1387 (O_1387,N_8490,N_6181);
xnor UO_1388 (O_1388,N_7460,N_5168);
and UO_1389 (O_1389,N_7903,N_6896);
and UO_1390 (O_1390,N_6673,N_5857);
and UO_1391 (O_1391,N_9893,N_7884);
nor UO_1392 (O_1392,N_9847,N_5588);
or UO_1393 (O_1393,N_6441,N_5390);
xnor UO_1394 (O_1394,N_9523,N_9689);
or UO_1395 (O_1395,N_9641,N_9854);
xor UO_1396 (O_1396,N_8618,N_9120);
xnor UO_1397 (O_1397,N_8431,N_9007);
nand UO_1398 (O_1398,N_9881,N_8026);
and UO_1399 (O_1399,N_8012,N_6921);
and UO_1400 (O_1400,N_5558,N_9174);
nor UO_1401 (O_1401,N_6230,N_6900);
nor UO_1402 (O_1402,N_6043,N_6735);
nor UO_1403 (O_1403,N_7953,N_8736);
or UO_1404 (O_1404,N_5379,N_6902);
nand UO_1405 (O_1405,N_5822,N_8220);
nand UO_1406 (O_1406,N_6126,N_7221);
and UO_1407 (O_1407,N_8597,N_8028);
xnor UO_1408 (O_1408,N_9296,N_8059);
or UO_1409 (O_1409,N_5758,N_7988);
nand UO_1410 (O_1410,N_8958,N_5383);
and UO_1411 (O_1411,N_7584,N_7996);
nand UO_1412 (O_1412,N_7567,N_9658);
xor UO_1413 (O_1413,N_8624,N_6053);
or UO_1414 (O_1414,N_6392,N_9708);
nor UO_1415 (O_1415,N_6127,N_6356);
or UO_1416 (O_1416,N_5415,N_8552);
or UO_1417 (O_1417,N_5169,N_7890);
nand UO_1418 (O_1418,N_6205,N_9958);
nor UO_1419 (O_1419,N_9563,N_5493);
xnor UO_1420 (O_1420,N_9546,N_7227);
nand UO_1421 (O_1421,N_6813,N_8763);
nor UO_1422 (O_1422,N_5381,N_5250);
or UO_1423 (O_1423,N_9538,N_6634);
or UO_1424 (O_1424,N_6470,N_5213);
or UO_1425 (O_1425,N_5206,N_9611);
xnor UO_1426 (O_1426,N_7808,N_8348);
or UO_1427 (O_1427,N_8916,N_6239);
nand UO_1428 (O_1428,N_5121,N_5142);
or UO_1429 (O_1429,N_9844,N_5010);
nand UO_1430 (O_1430,N_7240,N_5921);
and UO_1431 (O_1431,N_6734,N_9917);
nand UO_1432 (O_1432,N_7409,N_8680);
nor UO_1433 (O_1433,N_5668,N_5008);
nor UO_1434 (O_1434,N_8808,N_7704);
or UO_1435 (O_1435,N_8799,N_5220);
nor UO_1436 (O_1436,N_5150,N_6617);
nand UO_1437 (O_1437,N_5287,N_7590);
or UO_1438 (O_1438,N_9078,N_9697);
or UO_1439 (O_1439,N_5218,N_6772);
nor UO_1440 (O_1440,N_5236,N_5966);
nand UO_1441 (O_1441,N_8086,N_9506);
nand UO_1442 (O_1442,N_6773,N_8754);
nor UO_1443 (O_1443,N_9637,N_8414);
nand UO_1444 (O_1444,N_8063,N_8951);
and UO_1445 (O_1445,N_6164,N_7017);
xor UO_1446 (O_1446,N_9269,N_7661);
or UO_1447 (O_1447,N_8424,N_7430);
or UO_1448 (O_1448,N_6966,N_7844);
nor UO_1449 (O_1449,N_7090,N_9800);
xor UO_1450 (O_1450,N_5650,N_8833);
nand UO_1451 (O_1451,N_8614,N_7829);
or UO_1452 (O_1452,N_9808,N_8402);
nand UO_1453 (O_1453,N_9392,N_8327);
nand UO_1454 (O_1454,N_8667,N_6798);
nand UO_1455 (O_1455,N_9581,N_5046);
xnor UO_1456 (O_1456,N_6666,N_5087);
nor UO_1457 (O_1457,N_8107,N_6300);
or UO_1458 (O_1458,N_9131,N_6746);
and UO_1459 (O_1459,N_7103,N_8942);
nand UO_1460 (O_1460,N_8228,N_5970);
nor UO_1461 (O_1461,N_6717,N_7492);
nand UO_1462 (O_1462,N_7558,N_8690);
nand UO_1463 (O_1463,N_9372,N_5576);
and UO_1464 (O_1464,N_8376,N_9901);
or UO_1465 (O_1465,N_6674,N_5549);
nor UO_1466 (O_1466,N_6492,N_5188);
or UO_1467 (O_1467,N_8340,N_8691);
or UO_1468 (O_1468,N_7507,N_7050);
nor UO_1469 (O_1469,N_8451,N_7282);
nor UO_1470 (O_1470,N_5520,N_9387);
nor UO_1471 (O_1471,N_9565,N_9186);
or UO_1472 (O_1472,N_9034,N_7582);
and UO_1473 (O_1473,N_8788,N_7440);
nand UO_1474 (O_1474,N_5392,N_9352);
or UO_1475 (O_1475,N_8530,N_7058);
xor UO_1476 (O_1476,N_7870,N_9617);
and UO_1477 (O_1477,N_6150,N_6672);
or UO_1478 (O_1478,N_7775,N_5521);
and UO_1479 (O_1479,N_6984,N_8075);
xor UO_1480 (O_1480,N_7141,N_7036);
and UO_1481 (O_1481,N_7656,N_9657);
and UO_1482 (O_1482,N_9613,N_7427);
and UO_1483 (O_1483,N_6897,N_8264);
nand UO_1484 (O_1484,N_7252,N_7268);
or UO_1485 (O_1485,N_6545,N_9503);
nand UO_1486 (O_1486,N_5128,N_5776);
nor UO_1487 (O_1487,N_6578,N_7886);
and UO_1488 (O_1488,N_8956,N_6532);
or UO_1489 (O_1489,N_5849,N_7150);
xor UO_1490 (O_1490,N_5397,N_7257);
nor UO_1491 (O_1491,N_5908,N_8886);
nand UO_1492 (O_1492,N_8877,N_9440);
nor UO_1493 (O_1493,N_8947,N_6933);
nor UO_1494 (O_1494,N_8884,N_7337);
and UO_1495 (O_1495,N_9450,N_8186);
and UO_1496 (O_1496,N_8697,N_7367);
and UO_1497 (O_1497,N_5837,N_5636);
nor UO_1498 (O_1498,N_7577,N_8727);
or UO_1499 (O_1499,N_7818,N_9371);
endmodule