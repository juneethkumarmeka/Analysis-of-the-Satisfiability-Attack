module basic_1500_15000_2000_20_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_1362,In_900);
nand U1 (N_1,In_673,In_1235);
and U2 (N_2,In_1497,In_1240);
or U3 (N_3,In_908,In_1450);
nor U4 (N_4,In_1239,In_944);
nor U5 (N_5,In_391,In_478);
or U6 (N_6,In_203,In_77);
and U7 (N_7,In_335,In_287);
and U8 (N_8,In_1356,In_680);
or U9 (N_9,In_1165,In_244);
nor U10 (N_10,In_19,In_1255);
and U11 (N_11,In_1457,In_42);
or U12 (N_12,In_1327,In_1387);
nor U13 (N_13,In_1144,In_109);
or U14 (N_14,In_1238,In_1424);
nand U15 (N_15,In_884,In_1147);
nand U16 (N_16,In_426,In_1376);
nand U17 (N_17,In_828,In_1146);
nor U18 (N_18,In_877,In_738);
and U19 (N_19,In_855,In_1080);
or U20 (N_20,In_916,In_1474);
nor U21 (N_21,In_220,In_577);
or U22 (N_22,In_312,In_52);
and U23 (N_23,In_1445,In_556);
nand U24 (N_24,In_1477,In_1053);
nand U25 (N_25,In_274,In_982);
and U26 (N_26,In_1315,In_509);
or U27 (N_27,In_392,In_943);
or U28 (N_28,In_231,In_461);
and U29 (N_29,In_119,In_1451);
nand U30 (N_30,In_585,In_182);
or U31 (N_31,In_1429,In_258);
or U32 (N_32,In_242,In_554);
and U33 (N_33,In_394,In_713);
and U34 (N_34,In_471,In_1493);
or U35 (N_35,In_78,In_747);
and U36 (N_36,In_282,In_882);
nand U37 (N_37,In_261,In_1321);
and U38 (N_38,In_911,In_887);
nor U39 (N_39,In_278,In_474);
nor U40 (N_40,In_1231,In_12);
nor U41 (N_41,In_237,In_311);
or U42 (N_42,In_739,In_522);
nor U43 (N_43,In_752,In_997);
nand U44 (N_44,In_567,In_1126);
nor U45 (N_45,In_1192,In_1464);
nand U46 (N_46,In_219,In_682);
nand U47 (N_47,In_571,In_1314);
nand U48 (N_48,In_117,In_1041);
nand U49 (N_49,In_1408,In_634);
nand U50 (N_50,In_616,In_61);
or U51 (N_51,In_318,In_569);
and U52 (N_52,In_580,In_1128);
nor U53 (N_53,In_90,In_1068);
nand U54 (N_54,In_385,In_243);
and U55 (N_55,In_1092,In_198);
nand U56 (N_56,In_288,In_351);
or U57 (N_57,In_53,In_443);
nor U58 (N_58,In_24,In_126);
nand U59 (N_59,In_349,In_1027);
or U60 (N_60,In_775,In_500);
or U61 (N_61,In_625,In_130);
or U62 (N_62,In_423,In_446);
or U63 (N_63,In_240,In_1453);
nand U64 (N_64,In_1189,In_912);
nand U65 (N_65,In_1130,In_1182);
nand U66 (N_66,In_1277,In_1166);
and U67 (N_67,In_1466,In_910);
and U68 (N_68,In_1329,In_995);
nor U69 (N_69,In_812,In_1361);
and U70 (N_70,In_473,In_742);
nor U71 (N_71,In_1295,In_330);
or U72 (N_72,In_846,In_743);
nor U73 (N_73,In_783,In_353);
and U74 (N_74,In_544,In_133);
nor U75 (N_75,In_989,In_934);
nand U76 (N_76,In_451,In_487);
xor U77 (N_77,In_786,In_355);
nor U78 (N_78,In_1310,In_142);
nand U79 (N_79,In_650,In_1218);
or U80 (N_80,In_456,In_1434);
xnor U81 (N_81,In_976,In_1495);
nand U82 (N_82,In_578,In_1412);
nor U83 (N_83,In_396,In_284);
nand U84 (N_84,In_5,In_1286);
nand U85 (N_85,In_429,In_1015);
and U86 (N_86,In_1026,In_896);
or U87 (N_87,In_960,In_346);
and U88 (N_88,In_1479,In_922);
nand U89 (N_89,In_1004,In_407);
and U90 (N_90,In_1208,In_1273);
and U91 (N_91,In_157,In_513);
or U92 (N_92,In_457,In_29);
nor U93 (N_93,In_1317,In_476);
nor U94 (N_94,In_728,In_1485);
and U95 (N_95,In_602,In_1148);
nand U96 (N_96,In_361,In_1161);
nor U97 (N_97,In_520,In_290);
or U98 (N_98,In_668,In_86);
nand U99 (N_99,In_95,In_956);
nand U100 (N_100,In_804,In_1331);
nor U101 (N_101,In_1037,In_450);
xnor U102 (N_102,In_377,In_654);
or U103 (N_103,In_1051,In_606);
nand U104 (N_104,In_608,In_901);
or U105 (N_105,In_372,In_99);
nor U106 (N_106,In_1186,In_1256);
nand U107 (N_107,In_1353,In_563);
nand U108 (N_108,In_712,In_735);
or U109 (N_109,In_892,In_579);
or U110 (N_110,In_204,In_414);
nor U111 (N_111,In_135,In_310);
nand U112 (N_112,In_401,In_406);
or U113 (N_113,In_954,In_951);
nand U114 (N_114,In_1355,In_350);
or U115 (N_115,In_762,In_547);
or U116 (N_116,In_605,In_837);
nand U117 (N_117,In_723,In_1202);
nor U118 (N_118,In_525,In_1222);
nand U119 (N_119,In_811,In_48);
and U120 (N_120,In_440,In_1123);
or U121 (N_121,In_207,In_768);
or U122 (N_122,In_316,In_695);
or U123 (N_123,In_941,In_67);
nand U124 (N_124,In_868,In_766);
and U125 (N_125,In_949,In_25);
nand U126 (N_126,In_131,In_212);
and U127 (N_127,In_245,In_193);
or U128 (N_128,In_100,In_1122);
or U129 (N_129,In_1458,In_1253);
xor U130 (N_130,In_800,In_62);
and U131 (N_131,In_1334,In_570);
nor U132 (N_132,In_851,In_1431);
nor U133 (N_133,In_797,In_388);
nand U134 (N_134,In_1280,In_600);
or U135 (N_135,In_1430,In_1216);
and U136 (N_136,In_792,In_915);
nand U137 (N_137,In_81,In_291);
nor U138 (N_138,In_590,In_1022);
or U139 (N_139,In_151,In_345);
nor U140 (N_140,In_686,In_1496);
nor U141 (N_141,In_348,In_799);
nand U142 (N_142,In_1013,In_468);
or U143 (N_143,In_1044,In_44);
or U144 (N_144,In_187,In_1440);
or U145 (N_145,In_70,In_987);
and U146 (N_146,In_1030,In_1196);
and U147 (N_147,In_189,In_526);
or U148 (N_148,In_410,In_1211);
nand U149 (N_149,In_1336,In_58);
and U150 (N_150,In_1384,In_301);
or U151 (N_151,In_1061,In_517);
nand U152 (N_152,In_1489,In_558);
or U153 (N_153,In_55,In_455);
or U154 (N_154,In_999,In_645);
and U155 (N_155,In_232,In_1008);
or U156 (N_156,In_110,In_1108);
nand U157 (N_157,In_438,In_906);
or U158 (N_158,In_1323,In_1276);
nor U159 (N_159,In_787,In_420);
nand U160 (N_160,In_706,In_818);
nand U161 (N_161,In_338,In_913);
nor U162 (N_162,In_34,In_541);
nand U163 (N_163,In_950,In_59);
and U164 (N_164,In_11,In_635);
nor U165 (N_165,In_293,In_186);
or U166 (N_166,In_1324,In_166);
nand U167 (N_167,In_1404,In_94);
nor U168 (N_168,In_872,In_337);
nand U169 (N_169,In_753,In_694);
and U170 (N_170,In_856,In_741);
nor U171 (N_171,In_1330,In_924);
and U172 (N_172,In_121,In_134);
and U173 (N_173,In_754,In_1419);
nor U174 (N_174,In_617,In_619);
and U175 (N_175,In_128,In_1220);
or U176 (N_176,In_442,In_586);
nand U177 (N_177,In_1272,In_1198);
and U178 (N_178,In_1193,In_796);
or U179 (N_179,In_1071,In_1268);
nand U180 (N_180,In_1116,In_1232);
or U181 (N_181,In_444,In_241);
and U182 (N_182,In_160,In_519);
nand U183 (N_183,In_749,In_1195);
and U184 (N_184,In_909,In_1215);
and U185 (N_185,In_1019,In_795);
or U186 (N_186,In_501,In_632);
xor U187 (N_187,In_638,In_225);
or U188 (N_188,In_830,In_808);
or U189 (N_189,In_174,In_294);
nand U190 (N_190,In_1152,In_430);
nand U191 (N_191,In_1390,In_983);
or U192 (N_192,In_1149,In_1398);
or U193 (N_193,In_1210,In_1368);
and U194 (N_194,In_827,In_188);
and U195 (N_195,In_314,In_1476);
or U196 (N_196,In_1133,In_1306);
nand U197 (N_197,In_660,In_1075);
and U198 (N_198,In_737,In_593);
and U199 (N_199,In_1085,In_651);
and U200 (N_200,In_199,In_352);
or U201 (N_201,In_1074,In_824);
nor U202 (N_202,In_631,In_175);
and U203 (N_203,In_1005,In_1176);
nor U204 (N_204,In_698,In_1389);
or U205 (N_205,In_113,In_13);
and U206 (N_206,In_957,In_1400);
and U207 (N_207,In_953,In_1112);
and U208 (N_208,In_1246,In_163);
and U209 (N_209,In_1313,In_1098);
and U210 (N_210,In_14,In_197);
nor U211 (N_211,In_666,In_1282);
and U212 (N_212,In_507,In_412);
nand U213 (N_213,In_946,In_482);
or U214 (N_214,In_1170,In_530);
or U215 (N_215,In_1304,In_1339);
and U216 (N_216,In_1251,In_1415);
nor U217 (N_217,In_255,In_453);
nor U218 (N_218,In_1499,In_1179);
or U219 (N_219,In_432,In_20);
nand U220 (N_220,In_705,In_1183);
or U221 (N_221,In_497,In_825);
or U222 (N_222,In_503,In_143);
nor U223 (N_223,In_49,In_1250);
nand U224 (N_224,In_1248,In_1349);
and U225 (N_225,In_889,In_38);
or U226 (N_226,In_1145,In_209);
and U227 (N_227,In_445,In_1197);
or U228 (N_228,In_897,In_248);
nand U229 (N_229,In_68,In_138);
nor U230 (N_230,In_1350,In_21);
nand U231 (N_231,In_648,In_1254);
nor U232 (N_232,In_76,In_1088);
or U233 (N_233,In_1288,In_683);
nor U234 (N_234,In_144,In_535);
or U235 (N_235,In_1494,In_879);
nor U236 (N_236,In_1020,In_1000);
nand U237 (N_237,In_1091,In_79);
and U238 (N_238,In_793,In_1498);
or U239 (N_239,In_620,In_1343);
or U240 (N_240,In_192,In_782);
and U241 (N_241,In_974,In_433);
nor U242 (N_242,In_758,In_181);
and U243 (N_243,In_1120,In_623);
nor U244 (N_244,In_1100,In_779);
nand U245 (N_245,In_159,In_145);
nor U246 (N_246,In_120,In_930);
or U247 (N_247,In_228,In_331);
nor U248 (N_248,In_611,In_1438);
nand U249 (N_249,In_1229,In_194);
or U250 (N_250,In_104,In_527);
and U251 (N_251,In_85,In_1160);
nand U252 (N_252,In_1372,In_167);
nor U253 (N_253,In_1206,In_1351);
nand U254 (N_254,In_1473,In_176);
or U255 (N_255,In_780,In_376);
nand U256 (N_256,In_514,In_1094);
and U257 (N_257,In_1131,In_932);
and U258 (N_258,In_477,In_1428);
nand U259 (N_259,In_777,In_277);
nand U260 (N_260,In_1059,In_566);
and U261 (N_261,In_905,In_734);
nor U262 (N_262,In_458,In_844);
nand U263 (N_263,In_1433,In_454);
or U264 (N_264,In_172,In_1043);
xnor U265 (N_265,In_760,In_923);
and U266 (N_266,In_564,In_744);
nand U267 (N_267,In_729,In_424);
nand U268 (N_268,In_273,In_858);
and U269 (N_269,In_1337,In_1150);
nor U270 (N_270,In_494,In_1326);
and U271 (N_271,In_1153,In_836);
nand U272 (N_272,In_1490,In_367);
or U273 (N_273,In_82,In_899);
nor U274 (N_274,In_1487,In_389);
and U275 (N_275,In_480,In_853);
or U276 (N_276,In_1471,In_1032);
nand U277 (N_277,In_1348,In_1352);
nand U278 (N_278,In_1249,In_153);
and U279 (N_279,In_437,In_379);
or U280 (N_280,In_1258,In_1174);
nand U281 (N_281,In_1262,In_1180);
xor U282 (N_282,In_340,In_1111);
or U283 (N_283,In_693,In_127);
and U284 (N_284,In_832,In_1260);
nor U285 (N_285,In_546,In_411);
or U286 (N_286,In_746,In_572);
and U287 (N_287,In_1163,In_1296);
or U288 (N_288,In_628,In_1006);
and U289 (N_289,In_1184,In_1328);
or U290 (N_290,In_1157,In_765);
and U291 (N_291,In_1357,In_1118);
nor U292 (N_292,In_1492,In_537);
and U293 (N_293,In_971,In_17);
and U294 (N_294,In_1344,In_96);
nor U295 (N_295,In_1200,In_603);
or U296 (N_296,In_1454,In_1138);
nor U297 (N_297,In_977,In_1046);
or U298 (N_298,In_902,In_561);
and U299 (N_299,In_289,In_10);
nand U300 (N_300,In_1342,In_584);
nand U301 (N_301,In_1127,In_1391);
nand U302 (N_302,In_612,In_1385);
nand U303 (N_303,In_1265,In_576);
nor U304 (N_304,In_227,In_745);
and U305 (N_305,In_465,In_226);
nor U306 (N_306,In_607,In_1055);
or U307 (N_307,In_45,In_813);
nor U308 (N_308,In_557,In_1312);
and U309 (N_309,In_286,In_156);
and U310 (N_310,In_327,In_652);
nand U311 (N_311,In_663,In_534);
and U312 (N_312,In_1036,In_862);
nor U313 (N_313,In_1459,In_1099);
or U314 (N_314,In_1219,In_724);
or U315 (N_315,In_610,In_518);
and U316 (N_316,In_1468,In_1311);
nand U317 (N_317,In_1335,In_1201);
and U318 (N_318,In_402,In_472);
or U319 (N_319,In_89,In_1264);
or U320 (N_320,In_821,In_1093);
nor U321 (N_321,In_173,In_436);
or U322 (N_322,In_1395,In_646);
nand U323 (N_323,In_328,In_1401);
and U324 (N_324,In_1050,In_843);
or U325 (N_325,In_1345,In_926);
nor U326 (N_326,In_249,In_1114);
and U327 (N_327,In_1137,In_772);
nor U328 (N_328,In_727,In_667);
and U329 (N_329,In_806,In_1141);
or U330 (N_330,In_1241,In_116);
and U331 (N_331,In_1370,In_550);
nor U332 (N_332,In_931,In_368);
or U333 (N_333,In_103,In_1081);
nor U334 (N_334,In_581,In_1284);
or U335 (N_335,In_993,In_929);
nor U336 (N_336,In_904,In_553);
and U337 (N_337,In_1488,In_15);
nor U338 (N_338,In_770,In_1301);
nand U339 (N_339,In_1325,In_1191);
and U340 (N_340,In_803,In_84);
and U341 (N_341,In_861,In_279);
nand U342 (N_342,In_1411,In_1378);
and U343 (N_343,In_0,In_57);
and U344 (N_344,In_894,In_1244);
and U345 (N_345,In_1432,In_115);
nor U346 (N_346,In_4,In_1447);
nor U347 (N_347,In_303,In_1217);
and U348 (N_348,In_658,In_1441);
nand U349 (N_349,In_35,In_1084);
or U350 (N_350,In_604,In_191);
nor U351 (N_351,In_914,In_1397);
nor U352 (N_352,In_405,In_398);
and U353 (N_353,In_381,In_1230);
or U354 (N_354,In_1333,In_873);
and U355 (N_355,In_1076,In_994);
or U356 (N_356,In_1267,In_875);
and U357 (N_357,In_309,In_344);
nand U358 (N_358,In_515,In_1456);
and U359 (N_359,In_205,In_467);
nand U360 (N_360,In_141,In_1417);
nand U361 (N_361,In_1406,In_1279);
xor U362 (N_362,In_1444,In_63);
or U363 (N_363,In_92,In_991);
and U364 (N_364,In_774,In_164);
and U365 (N_365,In_216,In_492);
and U366 (N_366,In_215,In_702);
nand U367 (N_367,In_1382,In_626);
and U368 (N_368,In_1436,In_998);
nor U369 (N_369,In_699,In_326);
and U370 (N_370,In_1278,In_51);
and U371 (N_371,In_1380,In_955);
nor U372 (N_372,In_397,In_1448);
nor U373 (N_373,In_1105,In_1309);
or U374 (N_374,In_1205,In_980);
nor U375 (N_375,In_1287,In_814);
nor U376 (N_376,In_413,In_302);
nand U377 (N_377,In_1181,In_246);
nor U378 (N_378,In_575,In_489);
and U379 (N_379,In_1117,In_637);
and U380 (N_380,In_716,In_1);
nand U381 (N_381,In_1082,In_452);
nand U382 (N_382,In_1300,In_360);
or U383 (N_383,In_269,In_485);
nor U384 (N_384,In_1060,In_945);
nor U385 (N_385,In_1156,In_1292);
or U386 (N_386,In_973,In_685);
and U387 (N_387,In_921,In_859);
nor U388 (N_388,In_447,In_621);
nor U389 (N_389,In_664,In_395);
or U390 (N_390,In_486,In_137);
nor U391 (N_391,In_757,In_701);
or U392 (N_392,In_1318,In_1274);
or U393 (N_393,In_677,In_270);
nand U394 (N_394,In_74,In_1035);
and U395 (N_395,In_1143,In_601);
or U396 (N_396,In_523,In_1298);
nor U397 (N_397,In_988,In_1207);
or U398 (N_398,In_996,In_1307);
or U399 (N_399,In_107,In_823);
and U400 (N_400,In_1106,In_545);
nand U401 (N_401,In_937,In_463);
nand U402 (N_402,In_481,In_711);
nor U403 (N_403,In_236,In_629);
and U404 (N_404,In_1154,In_907);
nor U405 (N_405,In_1426,In_573);
nor U406 (N_406,In_959,In_97);
and U407 (N_407,In_657,In_1346);
or U408 (N_408,In_1052,In_551);
nor U409 (N_409,In_1394,In_948);
and U410 (N_410,In_30,In_435);
nor U411 (N_411,In_27,In_1285);
nor U412 (N_412,In_1422,In_1188);
nor U413 (N_413,In_252,In_891);
nand U414 (N_414,In_1119,In_850);
and U415 (N_415,In_408,In_674);
or U416 (N_416,In_177,In_1172);
nand U417 (N_417,In_1402,In_895);
nor U418 (N_418,In_365,In_506);
nand U419 (N_419,In_1469,In_649);
nand U420 (N_420,In_1365,In_597);
nand U421 (N_421,In_158,In_1129);
nand U422 (N_422,In_106,In_794);
nand U423 (N_423,In_1332,In_9);
nand U424 (N_424,In_785,In_155);
and U425 (N_425,In_1340,In_259);
nand U426 (N_426,In_816,In_967);
or U427 (N_427,In_280,In_149);
nor U428 (N_428,In_1449,In_118);
or U429 (N_429,In_721,In_1281);
nand U430 (N_430,In_1047,In_964);
nand U431 (N_431,In_75,In_919);
and U432 (N_432,In_562,In_1486);
nor U433 (N_433,In_1416,In_88);
nand U434 (N_434,In_829,In_1242);
or U435 (N_435,In_1101,In_317);
nand U436 (N_436,In_210,In_696);
and U437 (N_437,In_1113,In_1057);
nand U438 (N_438,In_334,In_1257);
and U439 (N_439,In_1104,In_356);
xnor U440 (N_440,In_1347,In_970);
and U441 (N_441,In_697,In_733);
or U442 (N_442,In_479,In_196);
nor U443 (N_443,In_18,In_1413);
or U444 (N_444,In_596,In_633);
and U445 (N_445,In_1109,In_588);
nand U446 (N_446,In_320,In_565);
or U447 (N_447,In_1374,In_1090);
nor U448 (N_448,In_1029,In_1140);
nor U449 (N_449,In_1173,In_615);
nand U450 (N_450,In_935,In_1168);
nand U451 (N_451,In_1031,In_874);
nor U452 (N_452,In_917,In_253);
nor U453 (N_453,In_112,In_1002);
nor U454 (N_454,In_152,In_1021);
nand U455 (N_455,In_1316,In_315);
or U456 (N_456,In_1442,In_548);
nor U457 (N_457,In_150,In_33);
nand U458 (N_458,In_920,In_965);
nor U459 (N_459,In_539,In_893);
nor U460 (N_460,In_325,In_703);
nor U461 (N_461,In_422,In_234);
nand U462 (N_462,In_574,In_1463);
nor U463 (N_463,In_1236,In_559);
or U464 (N_464,In_1465,In_213);
nor U465 (N_465,In_1245,In_1294);
nor U466 (N_466,In_878,In_1018);
or U467 (N_467,In_1283,In_162);
nor U468 (N_468,In_751,In_8);
nand U469 (N_469,In_1322,In_1012);
and U470 (N_470,In_329,In_475);
nand U471 (N_471,In_781,In_1199);
or U472 (N_472,In_139,In_1293);
nor U473 (N_473,In_3,In_528);
or U474 (N_474,In_459,In_979);
or U475 (N_475,In_984,In_1270);
and U476 (N_476,In_1048,In_502);
or U477 (N_477,In_613,In_1227);
nand U478 (N_478,In_470,In_885);
nor U479 (N_479,In_687,In_653);
nor U480 (N_480,In_1393,In_809);
and U481 (N_481,In_28,In_918);
nand U482 (N_482,In_594,In_549);
or U483 (N_483,In_1159,In_122);
nor U484 (N_484,In_400,In_516);
nand U485 (N_485,In_1096,In_540);
nor U486 (N_486,In_942,In_359);
or U487 (N_487,In_434,In_202);
nand U488 (N_488,In_750,In_1034);
or U489 (N_489,In_393,In_609);
or U490 (N_490,In_582,In_952);
and U491 (N_491,In_854,In_80);
or U492 (N_492,In_985,In_364);
nor U493 (N_493,In_986,In_272);
nor U494 (N_494,In_321,In_1399);
and U495 (N_495,In_1107,In_769);
or U496 (N_496,In_60,In_890);
nor U497 (N_497,In_807,In_449);
or U498 (N_498,In_676,In_1001);
or U499 (N_499,In_256,In_464);
nor U500 (N_500,In_238,In_690);
and U501 (N_501,In_1461,In_938);
and U502 (N_502,In_661,In_730);
and U503 (N_503,In_498,In_838);
xnor U504 (N_504,In_267,In_700);
nand U505 (N_505,In_1042,In_692);
and U506 (N_506,In_647,In_788);
nor U507 (N_507,In_1011,In_47);
nor U508 (N_508,In_23,In_1437);
nor U509 (N_509,In_627,In_1483);
nand U510 (N_510,In_441,In_656);
and U511 (N_511,In_1388,In_390);
nand U512 (N_512,In_732,In_857);
nand U513 (N_513,In_111,In_681);
nand U514 (N_514,In_409,In_867);
or U515 (N_515,In_493,In_1478);
or U516 (N_516,In_380,In_298);
or U517 (N_517,In_1407,In_1049);
nand U518 (N_518,In_250,In_383);
or U519 (N_519,In_200,In_266);
and U520 (N_520,In_46,In_927);
nor U521 (N_521,In_834,In_260);
nand U522 (N_522,In_1269,In_598);
or U523 (N_523,In_966,In_715);
and U524 (N_524,In_36,In_399);
and U525 (N_525,In_179,In_98);
and U526 (N_526,In_1110,In_140);
or U527 (N_527,In_132,In_839);
or U528 (N_528,In_333,In_925);
or U529 (N_529,In_1360,In_275);
nor U530 (N_530,In_1225,In_852);
and U531 (N_531,In_521,In_1097);
or U532 (N_532,In_1308,In_254);
and U533 (N_533,In_1291,In_771);
nand U534 (N_534,In_171,In_251);
nand U535 (N_535,In_866,In_387);
nor U536 (N_536,In_841,In_93);
and U537 (N_537,In_659,In_1358);
nand U538 (N_538,In_1421,In_524);
nand U539 (N_539,In_371,In_169);
nand U540 (N_540,In_431,In_1373);
nor U541 (N_541,In_840,In_759);
nor U542 (N_542,In_496,In_101);
nor U543 (N_543,In_1066,In_560);
or U544 (N_544,In_789,In_714);
nor U545 (N_545,In_835,In_65);
nor U546 (N_546,In_1009,In_1087);
nand U547 (N_547,In_1275,In_849);
nand U548 (N_548,In_871,In_1095);
and U549 (N_549,In_1045,In_1014);
nor U550 (N_550,In_1386,In_1243);
nand U551 (N_551,In_1038,In_1289);
or U552 (N_552,In_833,In_801);
nor U553 (N_553,In_972,In_1169);
or U554 (N_554,In_322,In_161);
nor U555 (N_555,In_1425,In_384);
and U556 (N_556,In_587,In_6);
nand U557 (N_557,In_589,In_168);
nor U558 (N_558,In_1132,In_817);
and U559 (N_559,In_1023,In_1016);
and U560 (N_560,In_936,In_642);
nor U561 (N_561,In_1266,In_1420);
nor U562 (N_562,In_1303,In_798);
nand U563 (N_563,In_1039,In_968);
or U564 (N_564,In_1366,In_704);
and U565 (N_565,In_981,In_1054);
nand U566 (N_566,In_1369,In_1263);
nand U567 (N_567,In_876,In_1379);
or U568 (N_568,In_102,In_1377);
nor U569 (N_569,In_323,In_211);
nand U570 (N_570,In_1079,In_1418);
and U571 (N_571,In_129,In_490);
nor U572 (N_572,In_555,In_510);
nor U573 (N_573,In_595,In_439);
nand U574 (N_574,In_1151,In_1410);
nor U575 (N_575,In_1375,In_764);
or U576 (N_576,In_183,In_416);
or U577 (N_577,In_1299,In_644);
nand U578 (N_578,In_722,In_417);
nor U579 (N_579,In_108,In_1142);
and U580 (N_580,In_136,In_1209);
or U581 (N_581,In_1136,In_427);
nand U582 (N_582,In_791,In_1063);
nand U583 (N_583,In_688,In_347);
or U584 (N_584,In_512,In_1115);
nand U585 (N_585,In_883,In_1024);
nor U586 (N_586,In_1072,In_975);
nor U587 (N_587,In_1363,In_418);
or U588 (N_588,In_1237,In_2);
nor U589 (N_589,In_1185,In_1452);
nand U590 (N_590,In_369,In_820);
or U591 (N_591,In_542,In_271);
and U592 (N_592,In_31,In_684);
or U593 (N_593,In_1077,In_1359);
and U594 (N_594,In_1446,In_614);
or U595 (N_595,In_1354,In_1396);
or U596 (N_596,In_1073,In_324);
nand U597 (N_597,In_425,In_1271);
nand U598 (N_598,In_1341,In_147);
nor U599 (N_599,In_933,In_357);
nor U600 (N_600,In_146,In_784);
and U601 (N_601,In_170,In_217);
and U602 (N_602,In_707,In_552);
nand U603 (N_603,In_87,In_662);
nor U604 (N_604,In_184,In_1070);
nand U605 (N_605,In_1083,In_748);
nand U606 (N_606,In_466,In_718);
and U607 (N_607,In_1252,In_1069);
or U608 (N_608,In_1134,In_1203);
nand U609 (N_609,In_448,In_1214);
and U610 (N_610,In_880,In_224);
nor U611 (N_611,In_1228,In_263);
nor U612 (N_612,In_214,In_1302);
nand U613 (N_613,In_16,In_374);
nand U614 (N_614,In_230,In_462);
nand U615 (N_615,In_283,In_1367);
or U616 (N_616,In_469,In_495);
or U617 (N_617,In_736,In_32);
or U618 (N_618,In_1439,In_947);
and U619 (N_619,In_1194,In_1423);
and U620 (N_620,In_1089,In_624);
or U621 (N_621,In_1187,In_1121);
nor U622 (N_622,In_306,In_708);
nor U623 (N_623,In_810,In_940);
and U624 (N_624,In_533,In_1204);
or U625 (N_625,In_190,In_56);
or U626 (N_626,In_148,In_591);
nor U627 (N_627,In_689,In_1058);
nor U628 (N_628,In_848,In_847);
nand U629 (N_629,In_1086,In_805);
nand U630 (N_630,In_543,In_71);
nand U631 (N_631,In_1234,In_990);
nand U632 (N_632,In_125,In_710);
nor U633 (N_633,In_778,In_292);
or U634 (N_634,In_358,In_819);
nor U635 (N_635,In_415,In_717);
or U636 (N_636,In_505,In_300);
nand U637 (N_637,In_257,In_903);
nor U638 (N_638,In_504,In_767);
or U639 (N_639,In_265,In_643);
nand U640 (N_640,In_756,In_1139);
nor U641 (N_641,In_460,In_341);
or U642 (N_642,In_1167,In_1247);
nor U643 (N_643,In_178,In_826);
and U644 (N_644,In_307,In_1040);
nand U645 (N_645,In_233,In_1409);
nor U646 (N_646,In_532,In_404);
nor U647 (N_647,In_709,In_1164);
and U648 (N_648,In_296,In_978);
or U649 (N_649,In_262,In_1427);
and U650 (N_650,In_961,In_881);
nor U651 (N_651,In_1135,In_1371);
or U652 (N_652,In_105,In_488);
or U653 (N_653,In_1482,In_1480);
and U654 (N_654,In_529,In_7);
nor U655 (N_655,In_869,In_428);
nand U656 (N_656,In_285,In_1158);
nand U657 (N_657,In_1364,In_221);
nand U658 (N_658,In_870,In_41);
and U659 (N_659,In_1297,In_1033);
and U660 (N_660,In_842,In_222);
or U661 (N_661,In_1025,In_1338);
and U662 (N_662,In_776,In_154);
and U663 (N_663,In_1305,In_1467);
and U664 (N_664,In_1383,In_672);
nand U665 (N_665,In_1472,In_304);
and U666 (N_666,In_264,In_1226);
nor U667 (N_667,In_740,In_790);
nand U668 (N_668,In_1484,In_1125);
or U669 (N_669,In_568,In_484);
and U670 (N_670,In_1470,In_731);
nand U671 (N_671,In_308,In_622);
and U672 (N_672,In_22,In_276);
or U673 (N_673,In_37,In_123);
nand U674 (N_674,In_1224,In_185);
or U675 (N_675,In_319,In_382);
or U676 (N_676,In_863,In_636);
nand U677 (N_677,In_339,In_1065);
nor U678 (N_678,In_332,In_1221);
nor U679 (N_679,In_508,In_1064);
nor U680 (N_680,In_726,In_1261);
or U681 (N_681,In_1190,In_1178);
nand U682 (N_682,In_538,In_1460);
and U683 (N_683,In_802,In_992);
and U684 (N_684,In_247,In_83);
nand U685 (N_685,In_342,In_618);
nand U686 (N_686,In_297,In_1320);
and U687 (N_687,In_822,In_958);
nor U688 (N_688,In_1062,In_640);
nor U689 (N_689,In_1481,In_40);
or U690 (N_690,In_1403,In_39);
nor U691 (N_691,In_218,In_229);
nor U692 (N_692,In_386,In_1010);
nor U693 (N_693,In_865,In_536);
nor U694 (N_694,In_50,In_375);
and U695 (N_695,In_419,In_669);
or U696 (N_696,In_1381,In_1491);
and U697 (N_697,In_1175,In_655);
or U698 (N_698,In_1124,In_354);
nor U699 (N_699,In_928,In_223);
nand U700 (N_700,In_763,In_678);
nor U701 (N_701,In_1475,In_1414);
nor U702 (N_702,In_1162,In_43);
xor U703 (N_703,In_1103,In_362);
nor U704 (N_704,In_64,In_26);
or U705 (N_705,In_343,In_755);
nand U706 (N_706,In_378,In_671);
and U707 (N_707,In_1102,In_268);
and U708 (N_708,In_583,In_691);
or U709 (N_709,In_1212,In_665);
nor U710 (N_710,In_1017,In_670);
nand U711 (N_711,In_675,In_720);
or U712 (N_712,In_124,In_511);
or U713 (N_713,In_373,In_421);
or U714 (N_714,In_1443,In_773);
nor U715 (N_715,In_239,In_1259);
nor U716 (N_716,In_295,In_1405);
and U717 (N_717,In_1171,In_888);
nor U718 (N_718,In_180,In_592);
nor U719 (N_719,In_639,In_363);
or U720 (N_720,In_165,In_403);
and U721 (N_721,In_531,In_630);
or U722 (N_722,In_69,In_860);
nor U723 (N_723,In_1177,In_1155);
nand U724 (N_724,In_1319,In_66);
nand U725 (N_725,In_864,In_1435);
and U726 (N_726,In_72,In_114);
or U727 (N_727,In_1078,In_898);
nor U728 (N_728,In_962,In_499);
and U729 (N_729,In_886,In_366);
or U730 (N_730,In_845,In_54);
nand U731 (N_731,In_1007,In_1462);
and U732 (N_732,In_336,In_599);
nand U733 (N_733,In_725,In_208);
nor U734 (N_734,In_195,In_73);
and U735 (N_735,In_641,In_1223);
or U736 (N_736,In_1028,In_1213);
nor U737 (N_737,In_815,In_305);
nand U738 (N_738,In_91,In_1392);
nand U739 (N_739,In_1056,In_831);
or U740 (N_740,In_761,In_963);
nand U741 (N_741,In_201,In_939);
nor U742 (N_742,In_1067,In_491);
nand U743 (N_743,In_719,In_206);
and U744 (N_744,In_969,In_235);
nand U745 (N_745,In_1233,In_1290);
or U746 (N_746,In_299,In_370);
and U747 (N_747,In_313,In_1003);
and U748 (N_748,In_1455,In_679);
and U749 (N_749,In_483,In_281);
or U750 (N_750,N_191,N_150);
nor U751 (N_751,N_537,N_529);
and U752 (N_752,N_551,N_700);
or U753 (N_753,N_454,N_379);
nand U754 (N_754,N_267,N_686);
and U755 (N_755,N_162,N_350);
or U756 (N_756,N_421,N_61);
and U757 (N_757,N_603,N_93);
nor U758 (N_758,N_546,N_221);
nor U759 (N_759,N_688,N_247);
nor U760 (N_760,N_97,N_527);
nand U761 (N_761,N_129,N_196);
or U762 (N_762,N_400,N_244);
and U763 (N_763,N_301,N_654);
and U764 (N_764,N_638,N_586);
nand U765 (N_765,N_538,N_134);
and U766 (N_766,N_572,N_189);
and U767 (N_767,N_10,N_656);
and U768 (N_768,N_45,N_288);
xor U769 (N_769,N_582,N_352);
or U770 (N_770,N_290,N_458);
nand U771 (N_771,N_506,N_100);
and U772 (N_772,N_73,N_67);
nor U773 (N_773,N_396,N_148);
nor U774 (N_774,N_530,N_9);
nor U775 (N_775,N_622,N_228);
nor U776 (N_776,N_147,N_659);
and U777 (N_777,N_377,N_20);
nor U778 (N_778,N_417,N_615);
and U779 (N_779,N_619,N_625);
and U780 (N_780,N_683,N_532);
or U781 (N_781,N_208,N_503);
nor U782 (N_782,N_57,N_704);
and U783 (N_783,N_88,N_299);
nand U784 (N_784,N_736,N_497);
nand U785 (N_785,N_416,N_660);
and U786 (N_786,N_263,N_284);
nand U787 (N_787,N_607,N_91);
and U788 (N_788,N_663,N_117);
or U789 (N_789,N_307,N_262);
and U790 (N_790,N_163,N_64);
nor U791 (N_791,N_116,N_87);
nand U792 (N_792,N_576,N_200);
nand U793 (N_793,N_701,N_174);
or U794 (N_794,N_329,N_110);
nand U795 (N_795,N_748,N_278);
nand U796 (N_796,N_337,N_351);
or U797 (N_797,N_606,N_171);
or U798 (N_798,N_491,N_697);
or U799 (N_799,N_685,N_154);
and U800 (N_800,N_480,N_369);
and U801 (N_801,N_399,N_453);
nor U802 (N_802,N_353,N_362);
nor U803 (N_803,N_627,N_408);
nand U804 (N_804,N_401,N_38);
nor U805 (N_805,N_469,N_272);
nand U806 (N_806,N_344,N_260);
nand U807 (N_807,N_501,N_520);
and U808 (N_808,N_695,N_270);
nor U809 (N_809,N_160,N_470);
or U810 (N_810,N_678,N_462);
and U811 (N_811,N_600,N_342);
nand U812 (N_812,N_133,N_511);
nand U813 (N_813,N_742,N_339);
and U814 (N_814,N_620,N_249);
and U815 (N_815,N_314,N_21);
or U816 (N_816,N_113,N_304);
or U817 (N_817,N_450,N_335);
nand U818 (N_818,N_223,N_481);
nor U819 (N_819,N_541,N_16);
or U820 (N_820,N_348,N_407);
nor U821 (N_821,N_598,N_673);
nand U822 (N_822,N_112,N_550);
nor U823 (N_823,N_323,N_166);
nor U824 (N_824,N_41,N_645);
or U825 (N_825,N_92,N_489);
nand U826 (N_826,N_526,N_563);
nand U827 (N_827,N_361,N_11);
nor U828 (N_828,N_302,N_53);
and U829 (N_829,N_6,N_712);
nor U830 (N_830,N_635,N_676);
or U831 (N_831,N_24,N_218);
and U832 (N_832,N_643,N_202);
and U833 (N_833,N_680,N_443);
or U834 (N_834,N_592,N_2);
or U835 (N_835,N_731,N_324);
or U836 (N_836,N_193,N_78);
and U837 (N_837,N_231,N_617);
nand U838 (N_838,N_601,N_207);
nand U839 (N_839,N_583,N_521);
and U840 (N_840,N_178,N_297);
or U841 (N_841,N_562,N_15);
and U842 (N_842,N_464,N_440);
and U843 (N_843,N_152,N_613);
nor U844 (N_844,N_226,N_54);
or U845 (N_845,N_512,N_35);
or U846 (N_846,N_98,N_80);
and U847 (N_847,N_315,N_292);
or U848 (N_848,N_32,N_291);
nor U849 (N_849,N_406,N_439);
or U850 (N_850,N_665,N_460);
nand U851 (N_851,N_390,N_664);
nand U852 (N_852,N_410,N_199);
and U853 (N_853,N_423,N_545);
nand U854 (N_854,N_146,N_611);
or U855 (N_855,N_373,N_326);
nand U856 (N_856,N_588,N_385);
and U857 (N_857,N_142,N_436);
nand U858 (N_858,N_571,N_658);
or U859 (N_859,N_246,N_310);
or U860 (N_860,N_60,N_52);
or U861 (N_861,N_43,N_79);
or U862 (N_862,N_415,N_340);
nand U863 (N_863,N_457,N_623);
nor U864 (N_864,N_283,N_599);
xor U865 (N_865,N_119,N_306);
and U866 (N_866,N_238,N_181);
nand U867 (N_867,N_99,N_426);
and U868 (N_868,N_186,N_381);
or U869 (N_869,N_641,N_220);
nand U870 (N_870,N_182,N_509);
or U871 (N_871,N_372,N_251);
and U872 (N_872,N_504,N_714);
nand U873 (N_873,N_203,N_420);
nand U874 (N_874,N_466,N_311);
or U875 (N_875,N_394,N_380);
or U876 (N_876,N_37,N_227);
or U877 (N_877,N_271,N_187);
nor U878 (N_878,N_4,N_636);
and U879 (N_879,N_371,N_253);
and U880 (N_880,N_528,N_281);
or U881 (N_881,N_725,N_575);
nand U882 (N_882,N_22,N_156);
or U883 (N_883,N_3,N_298);
or U884 (N_884,N_412,N_488);
nand U885 (N_885,N_386,N_157);
nor U886 (N_886,N_183,N_286);
nand U887 (N_887,N_492,N_188);
or U888 (N_888,N_455,N_164);
and U889 (N_889,N_698,N_86);
or U890 (N_890,N_734,N_82);
and U891 (N_891,N_513,N_425);
or U892 (N_892,N_68,N_233);
and U893 (N_893,N_728,N_1);
nand U894 (N_894,N_137,N_414);
nor U895 (N_895,N_320,N_39);
or U896 (N_896,N_89,N_424);
nor U897 (N_897,N_405,N_105);
or U898 (N_898,N_608,N_579);
and U899 (N_899,N_94,N_493);
nor U900 (N_900,N_544,N_723);
and U901 (N_901,N_367,N_177);
nand U902 (N_902,N_63,N_397);
or U903 (N_903,N_382,N_138);
and U904 (N_904,N_366,N_313);
nand U905 (N_905,N_479,N_168);
nand U906 (N_906,N_71,N_411);
and U907 (N_907,N_642,N_336);
and U908 (N_908,N_543,N_595);
or U909 (N_909,N_467,N_126);
nor U910 (N_910,N_248,N_490);
or U911 (N_911,N_27,N_487);
or U912 (N_912,N_590,N_328);
nor U913 (N_913,N_355,N_661);
nor U914 (N_914,N_523,N_709);
or U915 (N_915,N_327,N_525);
nor U916 (N_916,N_671,N_567);
nor U917 (N_917,N_437,N_631);
and U918 (N_918,N_215,N_732);
nand U919 (N_919,N_201,N_726);
nand U920 (N_920,N_713,N_46);
or U921 (N_921,N_741,N_596);
or U922 (N_922,N_17,N_19);
or U923 (N_923,N_710,N_42);
or U924 (N_924,N_357,N_427);
nor U925 (N_925,N_456,N_419);
and U926 (N_926,N_574,N_50);
nand U927 (N_927,N_114,N_743);
nor U928 (N_928,N_375,N_224);
nand U929 (N_929,N_31,N_681);
nor U930 (N_930,N_468,N_345);
nand U931 (N_931,N_475,N_719);
nor U932 (N_932,N_185,N_715);
and U933 (N_933,N_280,N_12);
nor U934 (N_934,N_747,N_522);
and U935 (N_935,N_438,N_29);
and U936 (N_936,N_593,N_165);
nand U937 (N_937,N_237,N_265);
nand U938 (N_938,N_36,N_121);
and U939 (N_939,N_359,N_261);
nand U940 (N_940,N_161,N_51);
nand U941 (N_941,N_618,N_5);
and U942 (N_942,N_616,N_358);
and U943 (N_943,N_295,N_275);
nor U944 (N_944,N_277,N_531);
nand U945 (N_945,N_318,N_395);
nand U946 (N_946,N_604,N_646);
and U947 (N_947,N_703,N_705);
and U948 (N_948,N_442,N_749);
and U949 (N_949,N_540,N_392);
and U950 (N_950,N_677,N_632);
or U951 (N_951,N_49,N_364);
nand U952 (N_952,N_136,N_431);
or U953 (N_953,N_384,N_149);
and U954 (N_954,N_95,N_533);
nand U955 (N_955,N_445,N_463);
and U956 (N_956,N_624,N_103);
nand U957 (N_957,N_172,N_552);
or U958 (N_958,N_192,N_518);
nor U959 (N_959,N_474,N_535);
nand U960 (N_960,N_34,N_140);
nor U961 (N_961,N_145,N_484);
or U962 (N_962,N_733,N_213);
and U963 (N_963,N_669,N_486);
and U964 (N_964,N_115,N_499);
nor U965 (N_965,N_626,N_374);
nand U966 (N_966,N_668,N_151);
nor U967 (N_967,N_347,N_609);
nor U968 (N_968,N_96,N_338);
or U969 (N_969,N_334,N_255);
and U970 (N_970,N_180,N_679);
nand U971 (N_971,N_434,N_158);
or U972 (N_972,N_670,N_430);
nor U973 (N_973,N_498,N_47);
nand U974 (N_974,N_81,N_691);
nor U975 (N_975,N_211,N_478);
nand U976 (N_976,N_252,N_124);
nand U977 (N_977,N_243,N_630);
nor U978 (N_978,N_418,N_745);
or U979 (N_979,N_0,N_516);
or U980 (N_980,N_305,N_730);
nor U981 (N_981,N_30,N_312);
or U982 (N_982,N_273,N_428);
and U983 (N_983,N_476,N_90);
and U984 (N_984,N_222,N_666);
nor U985 (N_985,N_234,N_122);
and U986 (N_986,N_413,N_610);
and U987 (N_987,N_109,N_628);
nor U988 (N_988,N_471,N_319);
nor U989 (N_989,N_648,N_66);
nand U990 (N_990,N_65,N_432);
or U991 (N_991,N_689,N_706);
or U992 (N_992,N_637,N_132);
nor U993 (N_993,N_155,N_331);
nor U994 (N_994,N_107,N_33);
and U995 (N_995,N_690,N_694);
nor U996 (N_996,N_507,N_120);
nand U997 (N_997,N_657,N_217);
nand U998 (N_998,N_106,N_287);
or U999 (N_999,N_317,N_111);
nor U1000 (N_1000,N_40,N_495);
nand U1001 (N_1001,N_118,N_303);
or U1002 (N_1002,N_716,N_274);
nor U1003 (N_1003,N_472,N_553);
and U1004 (N_1004,N_190,N_587);
nand U1005 (N_1005,N_449,N_614);
and U1006 (N_1006,N_18,N_542);
nand U1007 (N_1007,N_236,N_547);
and U1008 (N_1008,N_26,N_266);
or U1009 (N_1009,N_7,N_219);
nor U1010 (N_1010,N_707,N_360);
or U1011 (N_1011,N_605,N_232);
nor U1012 (N_1012,N_585,N_702);
or U1013 (N_1013,N_170,N_195);
nor U1014 (N_1014,N_308,N_591);
or U1015 (N_1015,N_565,N_564);
or U1016 (N_1016,N_139,N_56);
nand U1017 (N_1017,N_452,N_101);
nor U1018 (N_1018,N_74,N_108);
nand U1019 (N_1019,N_655,N_58);
nand U1020 (N_1020,N_556,N_722);
or U1021 (N_1021,N_578,N_241);
and U1022 (N_1022,N_104,N_404);
nor U1023 (N_1023,N_514,N_212);
or U1024 (N_1024,N_184,N_197);
or U1025 (N_1025,N_216,N_444);
nor U1026 (N_1026,N_433,N_293);
nand U1027 (N_1027,N_568,N_69);
or U1028 (N_1028,N_744,N_446);
or U1029 (N_1029,N_746,N_534);
nand U1030 (N_1030,N_354,N_387);
nand U1031 (N_1031,N_621,N_718);
nand U1032 (N_1032,N_173,N_692);
nand U1033 (N_1033,N_176,N_653);
or U1034 (N_1034,N_584,N_483);
or U1035 (N_1035,N_370,N_48);
or U1036 (N_1036,N_59,N_235);
and U1037 (N_1037,N_639,N_737);
and U1038 (N_1038,N_684,N_194);
nand U1039 (N_1039,N_332,N_602);
and U1040 (N_1040,N_256,N_515);
nor U1041 (N_1041,N_209,N_346);
and U1042 (N_1042,N_672,N_539);
nand U1043 (N_1043,N_740,N_496);
and U1044 (N_1044,N_210,N_77);
nor U1045 (N_1045,N_519,N_289);
or U1046 (N_1046,N_393,N_76);
and U1047 (N_1047,N_735,N_368);
and U1048 (N_1048,N_242,N_296);
nor U1049 (N_1049,N_465,N_720);
or U1050 (N_1050,N_125,N_28);
and U1051 (N_1051,N_153,N_557);
nand U1052 (N_1052,N_365,N_13);
and U1053 (N_1053,N_502,N_102);
nor U1054 (N_1054,N_383,N_693);
or U1055 (N_1055,N_240,N_581);
xor U1056 (N_1056,N_500,N_250);
nand U1057 (N_1057,N_577,N_687);
nor U1058 (N_1058,N_245,N_403);
nand U1059 (N_1059,N_205,N_640);
or U1060 (N_1060,N_198,N_555);
or U1061 (N_1061,N_179,N_388);
or U1062 (N_1062,N_536,N_135);
or U1063 (N_1063,N_389,N_727);
and U1064 (N_1064,N_675,N_651);
or U1065 (N_1065,N_300,N_333);
xor U1066 (N_1066,N_682,N_44);
or U1067 (N_1067,N_448,N_141);
nor U1068 (N_1068,N_508,N_696);
nand U1069 (N_1069,N_398,N_409);
or U1070 (N_1070,N_269,N_356);
and U1071 (N_1071,N_127,N_14);
nand U1072 (N_1072,N_634,N_322);
or U1073 (N_1073,N_451,N_229);
and U1074 (N_1074,N_662,N_285);
nand U1075 (N_1075,N_343,N_282);
nor U1076 (N_1076,N_128,N_667);
and U1077 (N_1077,N_376,N_309);
nand U1078 (N_1078,N_649,N_699);
and U1079 (N_1079,N_55,N_131);
and U1080 (N_1080,N_402,N_724);
nor U1081 (N_1081,N_70,N_321);
nand U1082 (N_1082,N_279,N_589);
nor U1083 (N_1083,N_633,N_62);
nor U1084 (N_1084,N_23,N_721);
and U1085 (N_1085,N_477,N_554);
nor U1086 (N_1086,N_349,N_558);
nor U1087 (N_1087,N_167,N_341);
nand U1088 (N_1088,N_144,N_594);
nor U1089 (N_1089,N_650,N_257);
or U1090 (N_1090,N_580,N_629);
or U1091 (N_1091,N_524,N_738);
nand U1092 (N_1092,N_214,N_83);
nor U1093 (N_1093,N_169,N_435);
and U1094 (N_1094,N_708,N_461);
nand U1095 (N_1095,N_473,N_597);
nor U1096 (N_1096,N_225,N_549);
and U1097 (N_1097,N_325,N_517);
nand U1098 (N_1098,N_276,N_561);
nor U1099 (N_1099,N_391,N_363);
or U1100 (N_1100,N_130,N_559);
and U1101 (N_1101,N_573,N_548);
nor U1102 (N_1102,N_75,N_510);
or U1103 (N_1103,N_644,N_316);
nand U1104 (N_1104,N_674,N_143);
and U1105 (N_1105,N_570,N_230);
nand U1106 (N_1106,N_441,N_485);
or U1107 (N_1107,N_239,N_717);
and U1108 (N_1108,N_294,N_206);
nor U1109 (N_1109,N_378,N_566);
nor U1110 (N_1110,N_560,N_123);
or U1111 (N_1111,N_729,N_505);
nand U1112 (N_1112,N_652,N_739);
and U1113 (N_1113,N_175,N_447);
xnor U1114 (N_1114,N_8,N_264);
nand U1115 (N_1115,N_429,N_612);
or U1116 (N_1116,N_459,N_422);
nor U1117 (N_1117,N_72,N_647);
nand U1118 (N_1118,N_268,N_84);
nand U1119 (N_1119,N_330,N_259);
nand U1120 (N_1120,N_258,N_569);
nor U1121 (N_1121,N_494,N_711);
nand U1122 (N_1122,N_204,N_25);
or U1123 (N_1123,N_254,N_85);
nor U1124 (N_1124,N_159,N_482);
or U1125 (N_1125,N_307,N_186);
or U1126 (N_1126,N_13,N_107);
nand U1127 (N_1127,N_471,N_197);
nand U1128 (N_1128,N_170,N_287);
or U1129 (N_1129,N_106,N_487);
and U1130 (N_1130,N_511,N_245);
nor U1131 (N_1131,N_610,N_370);
nor U1132 (N_1132,N_499,N_23);
nor U1133 (N_1133,N_469,N_376);
and U1134 (N_1134,N_622,N_692);
and U1135 (N_1135,N_493,N_632);
nor U1136 (N_1136,N_402,N_529);
nand U1137 (N_1137,N_122,N_534);
nor U1138 (N_1138,N_195,N_289);
or U1139 (N_1139,N_198,N_118);
nand U1140 (N_1140,N_135,N_616);
or U1141 (N_1141,N_21,N_216);
nor U1142 (N_1142,N_99,N_568);
and U1143 (N_1143,N_546,N_672);
nor U1144 (N_1144,N_269,N_632);
or U1145 (N_1145,N_112,N_554);
and U1146 (N_1146,N_632,N_514);
and U1147 (N_1147,N_435,N_261);
or U1148 (N_1148,N_184,N_668);
or U1149 (N_1149,N_318,N_723);
or U1150 (N_1150,N_495,N_129);
and U1151 (N_1151,N_308,N_700);
nor U1152 (N_1152,N_696,N_401);
nand U1153 (N_1153,N_736,N_91);
or U1154 (N_1154,N_399,N_417);
nand U1155 (N_1155,N_180,N_547);
and U1156 (N_1156,N_430,N_130);
and U1157 (N_1157,N_599,N_692);
or U1158 (N_1158,N_520,N_740);
or U1159 (N_1159,N_367,N_389);
nand U1160 (N_1160,N_375,N_461);
and U1161 (N_1161,N_669,N_683);
nand U1162 (N_1162,N_552,N_65);
and U1163 (N_1163,N_209,N_290);
nand U1164 (N_1164,N_237,N_693);
or U1165 (N_1165,N_696,N_579);
nor U1166 (N_1166,N_137,N_276);
and U1167 (N_1167,N_589,N_471);
and U1168 (N_1168,N_299,N_544);
and U1169 (N_1169,N_537,N_641);
and U1170 (N_1170,N_104,N_345);
nand U1171 (N_1171,N_381,N_680);
nor U1172 (N_1172,N_62,N_324);
nand U1173 (N_1173,N_59,N_287);
and U1174 (N_1174,N_444,N_441);
nand U1175 (N_1175,N_309,N_418);
nor U1176 (N_1176,N_137,N_127);
or U1177 (N_1177,N_620,N_183);
nor U1178 (N_1178,N_536,N_721);
or U1179 (N_1179,N_481,N_344);
or U1180 (N_1180,N_123,N_82);
nand U1181 (N_1181,N_48,N_295);
and U1182 (N_1182,N_721,N_438);
nor U1183 (N_1183,N_261,N_237);
nand U1184 (N_1184,N_124,N_549);
nor U1185 (N_1185,N_690,N_547);
and U1186 (N_1186,N_117,N_205);
nand U1187 (N_1187,N_280,N_619);
nand U1188 (N_1188,N_678,N_373);
and U1189 (N_1189,N_32,N_734);
or U1190 (N_1190,N_557,N_543);
xor U1191 (N_1191,N_159,N_469);
nor U1192 (N_1192,N_196,N_314);
nand U1193 (N_1193,N_591,N_748);
nand U1194 (N_1194,N_376,N_595);
or U1195 (N_1195,N_715,N_275);
nand U1196 (N_1196,N_293,N_79);
nand U1197 (N_1197,N_512,N_178);
nand U1198 (N_1198,N_144,N_277);
nand U1199 (N_1199,N_124,N_26);
or U1200 (N_1200,N_603,N_591);
or U1201 (N_1201,N_422,N_515);
or U1202 (N_1202,N_627,N_682);
nand U1203 (N_1203,N_634,N_386);
and U1204 (N_1204,N_107,N_705);
nand U1205 (N_1205,N_428,N_457);
and U1206 (N_1206,N_475,N_213);
or U1207 (N_1207,N_432,N_729);
nand U1208 (N_1208,N_248,N_158);
nor U1209 (N_1209,N_43,N_147);
nand U1210 (N_1210,N_473,N_523);
and U1211 (N_1211,N_515,N_288);
or U1212 (N_1212,N_579,N_338);
nor U1213 (N_1213,N_555,N_497);
nand U1214 (N_1214,N_718,N_435);
nor U1215 (N_1215,N_139,N_164);
xnor U1216 (N_1216,N_677,N_260);
nor U1217 (N_1217,N_329,N_466);
nor U1218 (N_1218,N_245,N_2);
nor U1219 (N_1219,N_254,N_737);
and U1220 (N_1220,N_272,N_491);
nor U1221 (N_1221,N_66,N_324);
and U1222 (N_1222,N_47,N_542);
nor U1223 (N_1223,N_50,N_144);
or U1224 (N_1224,N_262,N_622);
nand U1225 (N_1225,N_101,N_213);
nand U1226 (N_1226,N_151,N_564);
and U1227 (N_1227,N_466,N_327);
nand U1228 (N_1228,N_330,N_325);
nor U1229 (N_1229,N_388,N_649);
and U1230 (N_1230,N_316,N_699);
or U1231 (N_1231,N_645,N_637);
nand U1232 (N_1232,N_58,N_251);
nor U1233 (N_1233,N_0,N_101);
and U1234 (N_1234,N_357,N_217);
or U1235 (N_1235,N_6,N_551);
or U1236 (N_1236,N_178,N_94);
nand U1237 (N_1237,N_379,N_423);
nand U1238 (N_1238,N_399,N_737);
nand U1239 (N_1239,N_649,N_558);
nand U1240 (N_1240,N_123,N_68);
or U1241 (N_1241,N_722,N_713);
nor U1242 (N_1242,N_388,N_673);
or U1243 (N_1243,N_355,N_668);
and U1244 (N_1244,N_747,N_598);
and U1245 (N_1245,N_653,N_113);
or U1246 (N_1246,N_88,N_82);
and U1247 (N_1247,N_638,N_53);
or U1248 (N_1248,N_348,N_664);
and U1249 (N_1249,N_556,N_28);
and U1250 (N_1250,N_611,N_405);
and U1251 (N_1251,N_123,N_580);
nand U1252 (N_1252,N_259,N_205);
nand U1253 (N_1253,N_42,N_530);
or U1254 (N_1254,N_75,N_356);
nor U1255 (N_1255,N_416,N_405);
and U1256 (N_1256,N_395,N_156);
or U1257 (N_1257,N_253,N_673);
or U1258 (N_1258,N_395,N_734);
nor U1259 (N_1259,N_293,N_458);
nand U1260 (N_1260,N_203,N_110);
nand U1261 (N_1261,N_680,N_8);
and U1262 (N_1262,N_167,N_161);
nor U1263 (N_1263,N_5,N_245);
nor U1264 (N_1264,N_295,N_196);
or U1265 (N_1265,N_474,N_485);
and U1266 (N_1266,N_434,N_192);
nor U1267 (N_1267,N_293,N_740);
or U1268 (N_1268,N_143,N_396);
and U1269 (N_1269,N_730,N_493);
nand U1270 (N_1270,N_635,N_358);
nand U1271 (N_1271,N_508,N_136);
nand U1272 (N_1272,N_231,N_677);
and U1273 (N_1273,N_430,N_526);
and U1274 (N_1274,N_280,N_666);
nand U1275 (N_1275,N_319,N_189);
nor U1276 (N_1276,N_673,N_432);
nor U1277 (N_1277,N_263,N_223);
and U1278 (N_1278,N_274,N_82);
and U1279 (N_1279,N_309,N_435);
nand U1280 (N_1280,N_434,N_543);
and U1281 (N_1281,N_497,N_304);
nand U1282 (N_1282,N_566,N_111);
or U1283 (N_1283,N_224,N_647);
and U1284 (N_1284,N_280,N_637);
nand U1285 (N_1285,N_313,N_340);
nand U1286 (N_1286,N_279,N_675);
nand U1287 (N_1287,N_553,N_577);
and U1288 (N_1288,N_165,N_187);
or U1289 (N_1289,N_39,N_387);
and U1290 (N_1290,N_241,N_359);
nor U1291 (N_1291,N_252,N_386);
nand U1292 (N_1292,N_92,N_108);
and U1293 (N_1293,N_699,N_341);
and U1294 (N_1294,N_160,N_724);
nand U1295 (N_1295,N_133,N_672);
and U1296 (N_1296,N_695,N_527);
nor U1297 (N_1297,N_520,N_458);
nand U1298 (N_1298,N_13,N_603);
nor U1299 (N_1299,N_148,N_309);
or U1300 (N_1300,N_366,N_723);
and U1301 (N_1301,N_530,N_112);
nand U1302 (N_1302,N_217,N_462);
or U1303 (N_1303,N_124,N_664);
nand U1304 (N_1304,N_54,N_140);
nor U1305 (N_1305,N_512,N_118);
and U1306 (N_1306,N_0,N_443);
nand U1307 (N_1307,N_88,N_714);
nor U1308 (N_1308,N_271,N_370);
and U1309 (N_1309,N_36,N_663);
or U1310 (N_1310,N_455,N_303);
nor U1311 (N_1311,N_672,N_323);
nor U1312 (N_1312,N_212,N_131);
nand U1313 (N_1313,N_29,N_580);
nor U1314 (N_1314,N_63,N_563);
or U1315 (N_1315,N_102,N_645);
nand U1316 (N_1316,N_287,N_83);
or U1317 (N_1317,N_335,N_512);
nand U1318 (N_1318,N_257,N_167);
nand U1319 (N_1319,N_127,N_341);
nor U1320 (N_1320,N_608,N_346);
nand U1321 (N_1321,N_658,N_334);
and U1322 (N_1322,N_469,N_579);
or U1323 (N_1323,N_606,N_305);
or U1324 (N_1324,N_620,N_653);
and U1325 (N_1325,N_252,N_280);
or U1326 (N_1326,N_205,N_280);
nor U1327 (N_1327,N_81,N_285);
nor U1328 (N_1328,N_288,N_281);
nor U1329 (N_1329,N_49,N_166);
or U1330 (N_1330,N_683,N_335);
nor U1331 (N_1331,N_496,N_462);
or U1332 (N_1332,N_488,N_201);
and U1333 (N_1333,N_284,N_14);
nand U1334 (N_1334,N_266,N_2);
nand U1335 (N_1335,N_160,N_726);
or U1336 (N_1336,N_78,N_120);
nand U1337 (N_1337,N_321,N_408);
nor U1338 (N_1338,N_409,N_665);
and U1339 (N_1339,N_326,N_618);
and U1340 (N_1340,N_10,N_189);
nand U1341 (N_1341,N_273,N_223);
nand U1342 (N_1342,N_258,N_66);
nor U1343 (N_1343,N_749,N_627);
nand U1344 (N_1344,N_511,N_508);
and U1345 (N_1345,N_726,N_11);
or U1346 (N_1346,N_315,N_648);
nand U1347 (N_1347,N_52,N_740);
nor U1348 (N_1348,N_407,N_105);
and U1349 (N_1349,N_262,N_550);
and U1350 (N_1350,N_178,N_399);
nand U1351 (N_1351,N_676,N_35);
nand U1352 (N_1352,N_29,N_710);
or U1353 (N_1353,N_112,N_579);
or U1354 (N_1354,N_46,N_236);
or U1355 (N_1355,N_569,N_359);
and U1356 (N_1356,N_375,N_218);
or U1357 (N_1357,N_17,N_328);
or U1358 (N_1358,N_174,N_234);
and U1359 (N_1359,N_488,N_698);
nor U1360 (N_1360,N_384,N_610);
xor U1361 (N_1361,N_402,N_429);
nand U1362 (N_1362,N_381,N_129);
or U1363 (N_1363,N_538,N_66);
nor U1364 (N_1364,N_696,N_66);
and U1365 (N_1365,N_92,N_452);
and U1366 (N_1366,N_557,N_40);
nor U1367 (N_1367,N_571,N_118);
nor U1368 (N_1368,N_82,N_643);
nor U1369 (N_1369,N_583,N_0);
nor U1370 (N_1370,N_629,N_469);
nand U1371 (N_1371,N_506,N_627);
nor U1372 (N_1372,N_332,N_158);
or U1373 (N_1373,N_604,N_527);
or U1374 (N_1374,N_649,N_713);
or U1375 (N_1375,N_192,N_733);
nand U1376 (N_1376,N_483,N_42);
and U1377 (N_1377,N_682,N_492);
nor U1378 (N_1378,N_414,N_280);
nor U1379 (N_1379,N_636,N_160);
and U1380 (N_1380,N_548,N_288);
and U1381 (N_1381,N_226,N_174);
nor U1382 (N_1382,N_191,N_25);
nor U1383 (N_1383,N_159,N_582);
nand U1384 (N_1384,N_361,N_669);
nor U1385 (N_1385,N_638,N_245);
nand U1386 (N_1386,N_694,N_337);
nand U1387 (N_1387,N_84,N_216);
nor U1388 (N_1388,N_223,N_20);
nor U1389 (N_1389,N_464,N_399);
nor U1390 (N_1390,N_131,N_23);
nand U1391 (N_1391,N_363,N_541);
nor U1392 (N_1392,N_542,N_690);
nand U1393 (N_1393,N_369,N_656);
or U1394 (N_1394,N_28,N_474);
xnor U1395 (N_1395,N_678,N_713);
or U1396 (N_1396,N_566,N_5);
or U1397 (N_1397,N_405,N_635);
or U1398 (N_1398,N_673,N_707);
and U1399 (N_1399,N_224,N_257);
or U1400 (N_1400,N_510,N_544);
and U1401 (N_1401,N_435,N_306);
nand U1402 (N_1402,N_473,N_125);
and U1403 (N_1403,N_561,N_11);
nor U1404 (N_1404,N_593,N_537);
or U1405 (N_1405,N_157,N_383);
and U1406 (N_1406,N_574,N_607);
or U1407 (N_1407,N_367,N_12);
nand U1408 (N_1408,N_180,N_570);
nand U1409 (N_1409,N_722,N_60);
or U1410 (N_1410,N_712,N_234);
nand U1411 (N_1411,N_63,N_713);
or U1412 (N_1412,N_507,N_521);
or U1413 (N_1413,N_620,N_186);
nor U1414 (N_1414,N_737,N_89);
nand U1415 (N_1415,N_157,N_434);
and U1416 (N_1416,N_497,N_419);
nand U1417 (N_1417,N_398,N_364);
or U1418 (N_1418,N_738,N_737);
nand U1419 (N_1419,N_75,N_495);
nor U1420 (N_1420,N_133,N_582);
or U1421 (N_1421,N_72,N_650);
nor U1422 (N_1422,N_74,N_445);
and U1423 (N_1423,N_71,N_599);
and U1424 (N_1424,N_611,N_206);
nor U1425 (N_1425,N_469,N_37);
and U1426 (N_1426,N_168,N_245);
nor U1427 (N_1427,N_415,N_408);
nor U1428 (N_1428,N_599,N_418);
or U1429 (N_1429,N_28,N_640);
nor U1430 (N_1430,N_680,N_467);
nand U1431 (N_1431,N_443,N_84);
nor U1432 (N_1432,N_115,N_728);
nor U1433 (N_1433,N_339,N_441);
or U1434 (N_1434,N_594,N_27);
or U1435 (N_1435,N_156,N_155);
nand U1436 (N_1436,N_708,N_16);
nand U1437 (N_1437,N_5,N_502);
or U1438 (N_1438,N_429,N_333);
nor U1439 (N_1439,N_583,N_672);
nand U1440 (N_1440,N_656,N_249);
and U1441 (N_1441,N_574,N_440);
xor U1442 (N_1442,N_445,N_477);
nand U1443 (N_1443,N_215,N_97);
or U1444 (N_1444,N_270,N_520);
nand U1445 (N_1445,N_357,N_665);
nor U1446 (N_1446,N_281,N_406);
or U1447 (N_1447,N_368,N_139);
nand U1448 (N_1448,N_556,N_360);
nand U1449 (N_1449,N_624,N_490);
and U1450 (N_1450,N_72,N_669);
nand U1451 (N_1451,N_493,N_371);
nand U1452 (N_1452,N_191,N_629);
nor U1453 (N_1453,N_147,N_162);
and U1454 (N_1454,N_418,N_307);
or U1455 (N_1455,N_80,N_653);
and U1456 (N_1456,N_712,N_622);
nand U1457 (N_1457,N_523,N_581);
and U1458 (N_1458,N_221,N_418);
or U1459 (N_1459,N_647,N_362);
nor U1460 (N_1460,N_41,N_251);
nor U1461 (N_1461,N_551,N_615);
nand U1462 (N_1462,N_681,N_449);
nand U1463 (N_1463,N_720,N_636);
nor U1464 (N_1464,N_226,N_621);
nor U1465 (N_1465,N_579,N_583);
nand U1466 (N_1466,N_145,N_717);
and U1467 (N_1467,N_69,N_335);
nor U1468 (N_1468,N_577,N_123);
nor U1469 (N_1469,N_205,N_643);
nor U1470 (N_1470,N_98,N_539);
nor U1471 (N_1471,N_625,N_532);
and U1472 (N_1472,N_377,N_210);
or U1473 (N_1473,N_164,N_168);
nand U1474 (N_1474,N_245,N_142);
nor U1475 (N_1475,N_588,N_617);
nor U1476 (N_1476,N_215,N_44);
nor U1477 (N_1477,N_665,N_170);
and U1478 (N_1478,N_447,N_559);
and U1479 (N_1479,N_26,N_4);
and U1480 (N_1480,N_207,N_81);
or U1481 (N_1481,N_262,N_596);
and U1482 (N_1482,N_162,N_90);
or U1483 (N_1483,N_279,N_255);
and U1484 (N_1484,N_245,N_176);
nor U1485 (N_1485,N_221,N_657);
and U1486 (N_1486,N_369,N_639);
or U1487 (N_1487,N_212,N_355);
and U1488 (N_1488,N_50,N_222);
nor U1489 (N_1489,N_288,N_214);
nor U1490 (N_1490,N_521,N_640);
nor U1491 (N_1491,N_358,N_318);
and U1492 (N_1492,N_289,N_592);
nor U1493 (N_1493,N_226,N_661);
or U1494 (N_1494,N_408,N_668);
nor U1495 (N_1495,N_133,N_411);
nand U1496 (N_1496,N_49,N_99);
or U1497 (N_1497,N_361,N_116);
nor U1498 (N_1498,N_242,N_633);
nor U1499 (N_1499,N_155,N_436);
nand U1500 (N_1500,N_1397,N_1496);
nand U1501 (N_1501,N_1040,N_898);
nand U1502 (N_1502,N_1141,N_1183);
nand U1503 (N_1503,N_821,N_1333);
and U1504 (N_1504,N_1453,N_836);
nor U1505 (N_1505,N_864,N_1030);
nand U1506 (N_1506,N_876,N_1317);
nand U1507 (N_1507,N_886,N_920);
nand U1508 (N_1508,N_1407,N_1176);
and U1509 (N_1509,N_1203,N_1196);
nor U1510 (N_1510,N_914,N_1236);
nor U1511 (N_1511,N_1483,N_1089);
nor U1512 (N_1512,N_1171,N_751);
and U1513 (N_1513,N_1271,N_1231);
nor U1514 (N_1514,N_1081,N_1104);
nor U1515 (N_1515,N_1480,N_1395);
or U1516 (N_1516,N_799,N_925);
and U1517 (N_1517,N_1447,N_750);
or U1518 (N_1518,N_1027,N_1157);
nor U1519 (N_1519,N_1432,N_957);
nor U1520 (N_1520,N_1458,N_1002);
or U1521 (N_1521,N_1034,N_1044);
nor U1522 (N_1522,N_1289,N_1019);
nor U1523 (N_1523,N_1206,N_1495);
and U1524 (N_1524,N_1435,N_867);
or U1525 (N_1525,N_973,N_1471);
nand U1526 (N_1526,N_1046,N_1308);
nor U1527 (N_1527,N_1076,N_1360);
or U1528 (N_1528,N_827,N_1217);
nand U1529 (N_1529,N_934,N_1350);
nand U1530 (N_1530,N_1120,N_1390);
and U1531 (N_1531,N_767,N_849);
nor U1532 (N_1532,N_1187,N_1109);
or U1533 (N_1533,N_1466,N_1182);
nor U1534 (N_1534,N_978,N_875);
or U1535 (N_1535,N_912,N_814);
or U1536 (N_1536,N_882,N_1079);
nor U1537 (N_1537,N_972,N_951);
nor U1538 (N_1538,N_945,N_1322);
or U1539 (N_1539,N_1420,N_791);
or U1540 (N_1540,N_1055,N_1335);
and U1541 (N_1541,N_1169,N_1052);
and U1542 (N_1542,N_952,N_900);
and U1543 (N_1543,N_1123,N_771);
or U1544 (N_1544,N_1393,N_913);
and U1545 (N_1545,N_1475,N_1355);
or U1546 (N_1546,N_1073,N_872);
nor U1547 (N_1547,N_1313,N_1020);
and U1548 (N_1548,N_1150,N_1151);
nand U1549 (N_1549,N_996,N_1143);
nor U1550 (N_1550,N_1290,N_757);
nand U1551 (N_1551,N_1107,N_1400);
nand U1552 (N_1552,N_1232,N_1048);
or U1553 (N_1553,N_1374,N_1170);
and U1554 (N_1554,N_1037,N_1427);
or U1555 (N_1555,N_1383,N_1245);
nand U1556 (N_1556,N_1460,N_1185);
or U1557 (N_1557,N_1237,N_950);
nor U1558 (N_1558,N_1018,N_1003);
and U1559 (N_1559,N_1470,N_878);
nor U1560 (N_1560,N_1178,N_760);
nor U1561 (N_1561,N_933,N_1438);
and U1562 (N_1562,N_1340,N_793);
and U1563 (N_1563,N_1316,N_1474);
nor U1564 (N_1564,N_1106,N_1063);
or U1565 (N_1565,N_853,N_1184);
nor U1566 (N_1566,N_870,N_896);
nor U1567 (N_1567,N_1159,N_1090);
nand U1568 (N_1568,N_1315,N_1175);
and U1569 (N_1569,N_1416,N_923);
or U1570 (N_1570,N_1112,N_764);
nor U1571 (N_1571,N_982,N_852);
nor U1572 (N_1572,N_877,N_861);
or U1573 (N_1573,N_1299,N_1023);
nand U1574 (N_1574,N_1302,N_1325);
and U1575 (N_1575,N_924,N_761);
and U1576 (N_1576,N_850,N_974);
and U1577 (N_1577,N_819,N_956);
or U1578 (N_1578,N_1481,N_828);
nand U1579 (N_1579,N_1386,N_1300);
and U1580 (N_1580,N_1050,N_1225);
nor U1581 (N_1581,N_1147,N_879);
nor U1582 (N_1582,N_789,N_1411);
or U1583 (N_1583,N_797,N_1437);
nand U1584 (N_1584,N_1220,N_1005);
or U1585 (N_1585,N_1174,N_869);
nor U1586 (N_1586,N_1301,N_773);
or U1587 (N_1587,N_1028,N_1465);
or U1588 (N_1588,N_801,N_1281);
nor U1589 (N_1589,N_1066,N_1093);
nand U1590 (N_1590,N_1482,N_1263);
or U1591 (N_1591,N_860,N_863);
or U1592 (N_1592,N_755,N_1130);
nor U1593 (N_1593,N_1348,N_840);
or U1594 (N_1594,N_880,N_871);
or U1595 (N_1595,N_955,N_1469);
nand U1596 (N_1596,N_1294,N_780);
and U1597 (N_1597,N_1058,N_1456);
nor U1598 (N_1598,N_813,N_1221);
or U1599 (N_1599,N_1140,N_883);
nand U1600 (N_1600,N_784,N_833);
or U1601 (N_1601,N_901,N_1153);
nor U1602 (N_1602,N_774,N_1202);
nand U1603 (N_1603,N_1376,N_1423);
nand U1604 (N_1604,N_1372,N_1097);
or U1605 (N_1605,N_855,N_1062);
nor U1606 (N_1606,N_893,N_1015);
and U1607 (N_1607,N_1488,N_965);
nor U1608 (N_1608,N_1406,N_1408);
and U1609 (N_1609,N_1189,N_1096);
nor U1610 (N_1610,N_1441,N_1402);
and U1611 (N_1611,N_1233,N_1379);
nor U1612 (N_1612,N_1207,N_1007);
nor U1613 (N_1613,N_1000,N_1259);
and U1614 (N_1614,N_917,N_1378);
or U1615 (N_1615,N_1387,N_1158);
or U1616 (N_1616,N_936,N_987);
nand U1617 (N_1617,N_859,N_1428);
nand U1618 (N_1618,N_1454,N_809);
and U1619 (N_1619,N_1424,N_1381);
nor U1620 (N_1620,N_1014,N_1293);
and U1621 (N_1621,N_1326,N_1067);
or U1622 (N_1622,N_1247,N_1163);
or U1623 (N_1623,N_1074,N_1119);
nor U1624 (N_1624,N_1328,N_902);
and U1625 (N_1625,N_1056,N_975);
nand U1626 (N_1626,N_899,N_1115);
nand U1627 (N_1627,N_1144,N_1262);
nand U1628 (N_1628,N_1364,N_1190);
or U1629 (N_1629,N_765,N_788);
nand U1630 (N_1630,N_1138,N_1256);
or U1631 (N_1631,N_1330,N_1165);
or U1632 (N_1632,N_1219,N_1468);
nor U1633 (N_1633,N_1223,N_986);
nand U1634 (N_1634,N_1426,N_1270);
nor U1635 (N_1635,N_792,N_1195);
nor U1636 (N_1636,N_1113,N_1312);
nor U1637 (N_1637,N_1446,N_762);
nand U1638 (N_1638,N_1298,N_868);
nand U1639 (N_1639,N_1320,N_1248);
and U1640 (N_1640,N_1227,N_903);
and U1641 (N_1641,N_1108,N_829);
or U1642 (N_1642,N_752,N_817);
nand U1643 (N_1643,N_1442,N_775);
and U1644 (N_1644,N_1467,N_1425);
or U1645 (N_1645,N_1354,N_1486);
nand U1646 (N_1646,N_1384,N_874);
nor U1647 (N_1647,N_1489,N_769);
or U1648 (N_1648,N_1125,N_1049);
nand U1649 (N_1649,N_776,N_1356);
or U1650 (N_1650,N_1345,N_1297);
and U1651 (N_1651,N_781,N_1336);
nor U1652 (N_1652,N_1026,N_1121);
nand U1653 (N_1653,N_1092,N_1273);
nand U1654 (N_1654,N_1021,N_1373);
nor U1655 (N_1655,N_1314,N_783);
or U1656 (N_1656,N_1200,N_1082);
and U1657 (N_1657,N_1129,N_1124);
nand U1658 (N_1658,N_1095,N_824);
nand U1659 (N_1659,N_1332,N_842);
nor U1660 (N_1660,N_1351,N_910);
and U1661 (N_1661,N_1162,N_1116);
nand U1662 (N_1662,N_831,N_1161);
nand U1663 (N_1663,N_1166,N_1472);
or U1664 (N_1664,N_1088,N_1292);
xor U1665 (N_1665,N_1367,N_1168);
or U1666 (N_1666,N_1252,N_997);
nor U1667 (N_1667,N_1272,N_889);
nor U1668 (N_1668,N_1324,N_1417);
nor U1669 (N_1669,N_963,N_1181);
or U1670 (N_1670,N_1041,N_1327);
and U1671 (N_1671,N_1346,N_1286);
or U1672 (N_1672,N_1464,N_991);
nand U1673 (N_1673,N_835,N_888);
and U1674 (N_1674,N_1385,N_1392);
or U1675 (N_1675,N_1499,N_805);
or U1676 (N_1676,N_1053,N_949);
nor U1677 (N_1677,N_804,N_854);
nand U1678 (N_1678,N_1306,N_1337);
or U1679 (N_1679,N_895,N_1068);
nor U1680 (N_1680,N_873,N_1114);
nand U1681 (N_1681,N_1380,N_1004);
and U1682 (N_1682,N_1061,N_810);
nand U1683 (N_1683,N_1180,N_1016);
nand U1684 (N_1684,N_959,N_1038);
nand U1685 (N_1685,N_919,N_1358);
nand U1686 (N_1686,N_1216,N_967);
and U1687 (N_1687,N_1191,N_1445);
nand U1688 (N_1688,N_1264,N_998);
and U1689 (N_1689,N_1494,N_1008);
and U1690 (N_1690,N_1042,N_1398);
nand U1691 (N_1691,N_964,N_1269);
or U1692 (N_1692,N_1127,N_1208);
nand U1693 (N_1693,N_812,N_1085);
or U1694 (N_1694,N_1266,N_1137);
nand U1695 (N_1695,N_938,N_1031);
nor U1696 (N_1696,N_756,N_1421);
or U1697 (N_1697,N_848,N_931);
or U1698 (N_1698,N_1414,N_1497);
nor U1699 (N_1699,N_770,N_1257);
or U1700 (N_1700,N_946,N_918);
and U1701 (N_1701,N_1439,N_1403);
nor U1702 (N_1702,N_1240,N_1173);
or U1703 (N_1703,N_1246,N_1135);
and U1704 (N_1704,N_1131,N_795);
or U1705 (N_1705,N_922,N_1431);
and U1706 (N_1706,N_1152,N_1280);
nor U1707 (N_1707,N_1006,N_1359);
nor U1708 (N_1708,N_1283,N_1084);
nor U1709 (N_1709,N_1087,N_1122);
nand U1710 (N_1710,N_897,N_994);
or U1711 (N_1711,N_939,N_1487);
and U1712 (N_1712,N_1422,N_1224);
or U1713 (N_1713,N_1111,N_1249);
nand U1714 (N_1714,N_1405,N_1410);
and U1715 (N_1715,N_1197,N_823);
nor U1716 (N_1716,N_1349,N_846);
nor U1717 (N_1717,N_1440,N_1479);
or U1718 (N_1718,N_908,N_796);
nand U1719 (N_1719,N_865,N_1303);
nand U1720 (N_1720,N_1434,N_1267);
nand U1721 (N_1721,N_1103,N_807);
nand U1722 (N_1722,N_1274,N_1078);
or U1723 (N_1723,N_1241,N_1209);
and U1724 (N_1724,N_989,N_1101);
and U1725 (N_1725,N_1341,N_1244);
nand U1726 (N_1726,N_834,N_1370);
or U1727 (N_1727,N_794,N_1211);
nand U1728 (N_1728,N_1110,N_944);
nand U1729 (N_1729,N_932,N_826);
or U1730 (N_1730,N_1369,N_1279);
nand U1731 (N_1731,N_1133,N_1253);
nand U1732 (N_1732,N_1455,N_1357);
or U1733 (N_1733,N_1205,N_811);
or U1734 (N_1734,N_1099,N_1419);
nor U1735 (N_1735,N_1477,N_1045);
and U1736 (N_1736,N_927,N_1117);
and U1737 (N_1737,N_1134,N_1478);
or U1738 (N_1738,N_1156,N_970);
and U1739 (N_1739,N_1094,N_1035);
and U1740 (N_1740,N_1011,N_856);
or U1741 (N_1741,N_929,N_942);
and U1742 (N_1742,N_1484,N_1362);
and U1743 (N_1743,N_1275,N_984);
nor U1744 (N_1744,N_1091,N_977);
or U1745 (N_1745,N_1389,N_1155);
or U1746 (N_1746,N_1430,N_921);
or U1747 (N_1747,N_937,N_768);
or U1748 (N_1748,N_892,N_1366);
nor U1749 (N_1749,N_1083,N_1167);
nand U1750 (N_1750,N_1025,N_1451);
nor U1751 (N_1751,N_759,N_1188);
nand U1752 (N_1752,N_962,N_1295);
and U1753 (N_1753,N_862,N_980);
nor U1754 (N_1754,N_1001,N_1060);
and U1755 (N_1755,N_1069,N_1309);
nor U1756 (N_1756,N_1228,N_1010);
and U1757 (N_1757,N_1365,N_1457);
or U1758 (N_1758,N_841,N_930);
nor U1759 (N_1759,N_1287,N_1258);
nor U1760 (N_1760,N_1070,N_1282);
nand U1761 (N_1761,N_1118,N_995);
nor U1762 (N_1762,N_1239,N_881);
or U1763 (N_1763,N_985,N_1098);
or U1764 (N_1764,N_926,N_843);
nor U1765 (N_1765,N_1329,N_1210);
and U1766 (N_1766,N_753,N_1250);
nor U1767 (N_1767,N_1235,N_1319);
nand U1768 (N_1768,N_1450,N_1473);
or U1769 (N_1769,N_971,N_1128);
and U1770 (N_1770,N_1305,N_847);
and U1771 (N_1771,N_891,N_778);
and U1772 (N_1772,N_1436,N_1243);
nor U1773 (N_1773,N_1142,N_825);
nor U1774 (N_1774,N_818,N_1388);
and U1775 (N_1775,N_1218,N_911);
and U1776 (N_1776,N_1490,N_1404);
or U1777 (N_1777,N_885,N_1277);
nor U1778 (N_1778,N_906,N_1371);
and U1779 (N_1779,N_1036,N_1032);
and U1780 (N_1780,N_1375,N_1377);
nor U1781 (N_1781,N_1399,N_1164);
and U1782 (N_1782,N_1214,N_858);
or U1783 (N_1783,N_1304,N_1276);
or U1784 (N_1784,N_1194,N_993);
nor U1785 (N_1785,N_1201,N_1462);
or U1786 (N_1786,N_1353,N_1444);
and U1787 (N_1787,N_1017,N_1260);
and U1788 (N_1788,N_844,N_1461);
or U1789 (N_1789,N_968,N_787);
nand U1790 (N_1790,N_851,N_1051);
nand U1791 (N_1791,N_1285,N_1343);
or U1792 (N_1792,N_832,N_1009);
nor U1793 (N_1793,N_1323,N_1334);
or U1794 (N_1794,N_941,N_887);
nand U1795 (N_1795,N_943,N_1054);
nand U1796 (N_1796,N_894,N_1352);
or U1797 (N_1797,N_969,N_866);
nand U1798 (N_1798,N_800,N_816);
nor U1799 (N_1799,N_1064,N_890);
nand U1800 (N_1800,N_958,N_857);
nand U1801 (N_1801,N_1132,N_798);
or U1802 (N_1802,N_1013,N_1029);
nand U1803 (N_1803,N_1363,N_1251);
or U1804 (N_1804,N_1077,N_1459);
nor U1805 (N_1805,N_1296,N_1047);
nand U1806 (N_1806,N_1215,N_1492);
nor U1807 (N_1807,N_1476,N_1255);
and U1808 (N_1808,N_1493,N_1254);
or U1809 (N_1809,N_961,N_1012);
nand U1810 (N_1810,N_1149,N_1139);
and U1811 (N_1811,N_915,N_1172);
nand U1812 (N_1812,N_990,N_1086);
nor U1813 (N_1813,N_1284,N_1136);
nor U1814 (N_1814,N_960,N_1412);
nor U1815 (N_1815,N_1072,N_1193);
nand U1816 (N_1816,N_1105,N_839);
nor U1817 (N_1817,N_905,N_1198);
xnor U1818 (N_1818,N_909,N_1415);
and U1819 (N_1819,N_988,N_1368);
nand U1820 (N_1820,N_1059,N_779);
and U1821 (N_1821,N_1102,N_837);
and U1822 (N_1822,N_966,N_940);
or U1823 (N_1823,N_1033,N_1039);
or U1824 (N_1824,N_1022,N_1307);
or U1825 (N_1825,N_803,N_954);
or U1826 (N_1826,N_947,N_1278);
and U1827 (N_1827,N_1321,N_1242);
nor U1828 (N_1828,N_786,N_1331);
or U1829 (N_1829,N_1268,N_754);
or U1830 (N_1830,N_1145,N_1443);
or U1831 (N_1831,N_1212,N_1452);
and U1832 (N_1832,N_979,N_1261);
nand U1833 (N_1833,N_1288,N_1186);
nand U1834 (N_1834,N_1126,N_1265);
nor U1835 (N_1835,N_1222,N_806);
or U1836 (N_1836,N_1394,N_838);
nand U1837 (N_1837,N_1199,N_1146);
nand U1838 (N_1838,N_1485,N_1179);
or U1839 (N_1839,N_928,N_1361);
nand U1840 (N_1840,N_1449,N_758);
and U1841 (N_1841,N_1418,N_992);
or U1842 (N_1842,N_884,N_904);
nor U1843 (N_1843,N_1229,N_1382);
and U1844 (N_1844,N_916,N_1148);
and U1845 (N_1845,N_1413,N_830);
or U1846 (N_1846,N_1409,N_785);
or U1847 (N_1847,N_1230,N_1498);
and U1848 (N_1848,N_1043,N_1396);
or U1849 (N_1849,N_1226,N_1318);
and U1850 (N_1850,N_1154,N_790);
nor U1851 (N_1851,N_1491,N_777);
and U1852 (N_1852,N_1338,N_845);
and U1853 (N_1853,N_763,N_1448);
xor U1854 (N_1854,N_1100,N_1057);
or U1855 (N_1855,N_999,N_802);
xor U1856 (N_1856,N_1160,N_766);
nand U1857 (N_1857,N_953,N_820);
or U1858 (N_1858,N_1463,N_1311);
or U1859 (N_1859,N_948,N_1433);
or U1860 (N_1860,N_1344,N_1339);
and U1861 (N_1861,N_1347,N_1204);
and U1862 (N_1862,N_1310,N_1234);
or U1863 (N_1863,N_1192,N_815);
or U1864 (N_1864,N_1024,N_1080);
and U1865 (N_1865,N_1429,N_1075);
or U1866 (N_1866,N_1291,N_782);
nand U1867 (N_1867,N_976,N_1065);
or U1868 (N_1868,N_1177,N_1342);
nor U1869 (N_1869,N_822,N_1391);
nor U1870 (N_1870,N_808,N_1213);
or U1871 (N_1871,N_981,N_1071);
nand U1872 (N_1872,N_935,N_1401);
and U1873 (N_1873,N_983,N_907);
nand U1874 (N_1874,N_772,N_1238);
nand U1875 (N_1875,N_806,N_1243);
nor U1876 (N_1876,N_933,N_1221);
nor U1877 (N_1877,N_1096,N_1460);
and U1878 (N_1878,N_1176,N_1158);
nor U1879 (N_1879,N_922,N_1146);
and U1880 (N_1880,N_1418,N_794);
and U1881 (N_1881,N_785,N_1498);
or U1882 (N_1882,N_1441,N_1066);
or U1883 (N_1883,N_1498,N_1299);
or U1884 (N_1884,N_1469,N_1426);
or U1885 (N_1885,N_1146,N_1181);
and U1886 (N_1886,N_917,N_1439);
or U1887 (N_1887,N_1214,N_937);
and U1888 (N_1888,N_1328,N_1369);
or U1889 (N_1889,N_1088,N_827);
nand U1890 (N_1890,N_1463,N_902);
nor U1891 (N_1891,N_1071,N_1464);
or U1892 (N_1892,N_992,N_1278);
and U1893 (N_1893,N_1064,N_781);
nand U1894 (N_1894,N_1039,N_1145);
and U1895 (N_1895,N_1223,N_1228);
nand U1896 (N_1896,N_819,N_1057);
or U1897 (N_1897,N_935,N_1160);
or U1898 (N_1898,N_991,N_904);
and U1899 (N_1899,N_864,N_1123);
or U1900 (N_1900,N_925,N_1321);
and U1901 (N_1901,N_1091,N_795);
nand U1902 (N_1902,N_1457,N_937);
and U1903 (N_1903,N_1064,N_1259);
or U1904 (N_1904,N_1272,N_1006);
and U1905 (N_1905,N_1017,N_1163);
nor U1906 (N_1906,N_818,N_1478);
nor U1907 (N_1907,N_1396,N_1041);
and U1908 (N_1908,N_1328,N_848);
nor U1909 (N_1909,N_911,N_1337);
nor U1910 (N_1910,N_1493,N_1308);
and U1911 (N_1911,N_1273,N_1284);
and U1912 (N_1912,N_1418,N_1211);
nor U1913 (N_1913,N_1285,N_1178);
and U1914 (N_1914,N_1328,N_898);
or U1915 (N_1915,N_1233,N_1447);
or U1916 (N_1916,N_972,N_841);
or U1917 (N_1917,N_855,N_824);
nand U1918 (N_1918,N_908,N_1080);
nor U1919 (N_1919,N_1008,N_1478);
and U1920 (N_1920,N_1280,N_1250);
nand U1921 (N_1921,N_1266,N_1209);
or U1922 (N_1922,N_826,N_931);
and U1923 (N_1923,N_1252,N_1125);
nor U1924 (N_1924,N_1357,N_785);
or U1925 (N_1925,N_1164,N_1091);
and U1926 (N_1926,N_805,N_1351);
nor U1927 (N_1927,N_886,N_898);
nand U1928 (N_1928,N_1283,N_1460);
and U1929 (N_1929,N_1187,N_1163);
nand U1930 (N_1930,N_967,N_825);
and U1931 (N_1931,N_1418,N_1465);
nand U1932 (N_1932,N_1454,N_1257);
and U1933 (N_1933,N_1463,N_1319);
nand U1934 (N_1934,N_1389,N_1195);
or U1935 (N_1935,N_1493,N_789);
and U1936 (N_1936,N_1407,N_1154);
or U1937 (N_1937,N_852,N_1212);
and U1938 (N_1938,N_1107,N_1237);
nor U1939 (N_1939,N_831,N_1031);
or U1940 (N_1940,N_1266,N_1341);
nand U1941 (N_1941,N_1174,N_1336);
nand U1942 (N_1942,N_899,N_1239);
nor U1943 (N_1943,N_1343,N_1048);
or U1944 (N_1944,N_1097,N_1287);
nand U1945 (N_1945,N_997,N_1307);
nand U1946 (N_1946,N_797,N_1433);
and U1947 (N_1947,N_814,N_1121);
or U1948 (N_1948,N_1155,N_1109);
or U1949 (N_1949,N_1438,N_1015);
or U1950 (N_1950,N_1007,N_1217);
nand U1951 (N_1951,N_1495,N_998);
or U1952 (N_1952,N_1014,N_1100);
nor U1953 (N_1953,N_909,N_1490);
and U1954 (N_1954,N_1259,N_1496);
nor U1955 (N_1955,N_1217,N_1269);
nand U1956 (N_1956,N_1499,N_935);
and U1957 (N_1957,N_1077,N_954);
nand U1958 (N_1958,N_1345,N_1181);
or U1959 (N_1959,N_840,N_817);
or U1960 (N_1960,N_1201,N_989);
nor U1961 (N_1961,N_1498,N_1255);
or U1962 (N_1962,N_987,N_800);
nand U1963 (N_1963,N_1306,N_1316);
or U1964 (N_1964,N_1244,N_944);
nand U1965 (N_1965,N_1022,N_1318);
and U1966 (N_1966,N_927,N_1132);
and U1967 (N_1967,N_788,N_960);
nor U1968 (N_1968,N_1387,N_1083);
nand U1969 (N_1969,N_860,N_771);
nor U1970 (N_1970,N_905,N_1046);
nand U1971 (N_1971,N_1208,N_977);
nor U1972 (N_1972,N_953,N_1394);
or U1973 (N_1973,N_1317,N_964);
or U1974 (N_1974,N_1407,N_1331);
nor U1975 (N_1975,N_783,N_1286);
and U1976 (N_1976,N_1436,N_1271);
or U1977 (N_1977,N_886,N_987);
nor U1978 (N_1978,N_852,N_1258);
or U1979 (N_1979,N_1223,N_1420);
nand U1980 (N_1980,N_1429,N_929);
nor U1981 (N_1981,N_832,N_774);
nand U1982 (N_1982,N_1019,N_1131);
nand U1983 (N_1983,N_892,N_1257);
nand U1984 (N_1984,N_1023,N_783);
nor U1985 (N_1985,N_1273,N_1155);
nor U1986 (N_1986,N_1366,N_1361);
and U1987 (N_1987,N_1359,N_979);
and U1988 (N_1988,N_1327,N_1174);
and U1989 (N_1989,N_811,N_1287);
nand U1990 (N_1990,N_1005,N_779);
nor U1991 (N_1991,N_1062,N_1096);
and U1992 (N_1992,N_1369,N_1332);
or U1993 (N_1993,N_1284,N_1458);
and U1994 (N_1994,N_940,N_1185);
and U1995 (N_1995,N_1469,N_912);
xor U1996 (N_1996,N_806,N_1257);
and U1997 (N_1997,N_815,N_929);
nor U1998 (N_1998,N_1045,N_935);
nor U1999 (N_1999,N_1334,N_814);
nor U2000 (N_2000,N_1430,N_758);
or U2001 (N_2001,N_958,N_1338);
or U2002 (N_2002,N_881,N_1020);
and U2003 (N_2003,N_1340,N_1343);
nor U2004 (N_2004,N_1055,N_751);
nand U2005 (N_2005,N_1166,N_1297);
and U2006 (N_2006,N_1244,N_829);
nor U2007 (N_2007,N_1215,N_1300);
nand U2008 (N_2008,N_1378,N_1202);
nor U2009 (N_2009,N_1183,N_1380);
or U2010 (N_2010,N_777,N_911);
nor U2011 (N_2011,N_1036,N_920);
or U2012 (N_2012,N_1362,N_1381);
and U2013 (N_2013,N_752,N_1468);
and U2014 (N_2014,N_1468,N_1005);
nand U2015 (N_2015,N_1435,N_834);
nand U2016 (N_2016,N_1029,N_1253);
or U2017 (N_2017,N_830,N_1023);
or U2018 (N_2018,N_901,N_1457);
nand U2019 (N_2019,N_1045,N_1329);
nand U2020 (N_2020,N_1089,N_877);
nor U2021 (N_2021,N_1045,N_1317);
nand U2022 (N_2022,N_1265,N_1445);
or U2023 (N_2023,N_1487,N_984);
and U2024 (N_2024,N_1091,N_857);
nor U2025 (N_2025,N_1441,N_1357);
and U2026 (N_2026,N_787,N_988);
or U2027 (N_2027,N_1016,N_817);
nand U2028 (N_2028,N_1028,N_1333);
or U2029 (N_2029,N_1483,N_875);
and U2030 (N_2030,N_799,N_1224);
and U2031 (N_2031,N_930,N_993);
and U2032 (N_2032,N_1235,N_1068);
nor U2033 (N_2033,N_1066,N_1435);
xor U2034 (N_2034,N_1044,N_1461);
nor U2035 (N_2035,N_1262,N_1282);
nand U2036 (N_2036,N_1192,N_885);
nand U2037 (N_2037,N_1355,N_1233);
and U2038 (N_2038,N_1376,N_1463);
nand U2039 (N_2039,N_1490,N_1382);
nor U2040 (N_2040,N_1026,N_1278);
or U2041 (N_2041,N_798,N_1457);
xor U2042 (N_2042,N_1274,N_1445);
and U2043 (N_2043,N_1422,N_1359);
or U2044 (N_2044,N_1094,N_1167);
and U2045 (N_2045,N_1041,N_900);
or U2046 (N_2046,N_766,N_874);
nand U2047 (N_2047,N_1307,N_1145);
and U2048 (N_2048,N_1129,N_1035);
or U2049 (N_2049,N_1074,N_1090);
or U2050 (N_2050,N_1489,N_1145);
nand U2051 (N_2051,N_1155,N_1431);
and U2052 (N_2052,N_892,N_871);
nand U2053 (N_2053,N_1423,N_1444);
nor U2054 (N_2054,N_881,N_1081);
and U2055 (N_2055,N_1063,N_1477);
and U2056 (N_2056,N_1108,N_1076);
nor U2057 (N_2057,N_759,N_1027);
or U2058 (N_2058,N_1300,N_1131);
and U2059 (N_2059,N_1338,N_997);
nand U2060 (N_2060,N_1412,N_847);
and U2061 (N_2061,N_1276,N_935);
and U2062 (N_2062,N_931,N_1113);
and U2063 (N_2063,N_769,N_1273);
nand U2064 (N_2064,N_1037,N_924);
nand U2065 (N_2065,N_999,N_781);
and U2066 (N_2066,N_1218,N_850);
and U2067 (N_2067,N_1121,N_1434);
and U2068 (N_2068,N_1444,N_1107);
nand U2069 (N_2069,N_808,N_1224);
nor U2070 (N_2070,N_1097,N_1141);
or U2071 (N_2071,N_962,N_1289);
or U2072 (N_2072,N_820,N_1073);
nor U2073 (N_2073,N_939,N_1412);
or U2074 (N_2074,N_1456,N_1356);
and U2075 (N_2075,N_967,N_1186);
or U2076 (N_2076,N_1255,N_1231);
nand U2077 (N_2077,N_1433,N_1170);
nor U2078 (N_2078,N_945,N_1088);
nor U2079 (N_2079,N_1207,N_821);
and U2080 (N_2080,N_1484,N_1338);
nor U2081 (N_2081,N_1188,N_969);
nor U2082 (N_2082,N_1192,N_1101);
or U2083 (N_2083,N_1297,N_1262);
or U2084 (N_2084,N_1398,N_1048);
or U2085 (N_2085,N_1005,N_774);
nor U2086 (N_2086,N_1017,N_1480);
nand U2087 (N_2087,N_1207,N_1332);
and U2088 (N_2088,N_936,N_1118);
or U2089 (N_2089,N_785,N_1331);
and U2090 (N_2090,N_1267,N_810);
or U2091 (N_2091,N_1106,N_1183);
nand U2092 (N_2092,N_1458,N_1168);
nand U2093 (N_2093,N_1294,N_1123);
and U2094 (N_2094,N_933,N_1277);
and U2095 (N_2095,N_1163,N_1264);
nand U2096 (N_2096,N_1313,N_1042);
or U2097 (N_2097,N_1268,N_990);
or U2098 (N_2098,N_1338,N_1081);
nor U2099 (N_2099,N_1387,N_823);
nand U2100 (N_2100,N_1221,N_1247);
and U2101 (N_2101,N_1464,N_870);
nor U2102 (N_2102,N_1030,N_1170);
nand U2103 (N_2103,N_1208,N_794);
nor U2104 (N_2104,N_1079,N_793);
and U2105 (N_2105,N_815,N_1256);
or U2106 (N_2106,N_1180,N_911);
or U2107 (N_2107,N_845,N_1284);
and U2108 (N_2108,N_1155,N_818);
and U2109 (N_2109,N_832,N_1361);
or U2110 (N_2110,N_1308,N_945);
or U2111 (N_2111,N_935,N_1124);
and U2112 (N_2112,N_876,N_1083);
nor U2113 (N_2113,N_995,N_1089);
nand U2114 (N_2114,N_1438,N_1130);
or U2115 (N_2115,N_1191,N_1016);
nor U2116 (N_2116,N_1144,N_922);
nand U2117 (N_2117,N_838,N_951);
nand U2118 (N_2118,N_803,N_1401);
or U2119 (N_2119,N_1037,N_1362);
or U2120 (N_2120,N_1102,N_1346);
and U2121 (N_2121,N_1101,N_823);
nand U2122 (N_2122,N_843,N_1107);
nand U2123 (N_2123,N_1441,N_1454);
nand U2124 (N_2124,N_878,N_1207);
nand U2125 (N_2125,N_1295,N_1025);
and U2126 (N_2126,N_1287,N_1182);
nor U2127 (N_2127,N_1168,N_1283);
or U2128 (N_2128,N_951,N_872);
or U2129 (N_2129,N_1244,N_929);
or U2130 (N_2130,N_1029,N_1069);
and U2131 (N_2131,N_1400,N_1439);
or U2132 (N_2132,N_751,N_1022);
xor U2133 (N_2133,N_1085,N_1107);
or U2134 (N_2134,N_920,N_1056);
nor U2135 (N_2135,N_1242,N_964);
and U2136 (N_2136,N_1091,N_1140);
and U2137 (N_2137,N_1231,N_1273);
nor U2138 (N_2138,N_1436,N_973);
nand U2139 (N_2139,N_827,N_826);
nor U2140 (N_2140,N_764,N_847);
and U2141 (N_2141,N_771,N_1395);
nor U2142 (N_2142,N_1217,N_1484);
nor U2143 (N_2143,N_764,N_1003);
nor U2144 (N_2144,N_1485,N_1167);
or U2145 (N_2145,N_958,N_764);
and U2146 (N_2146,N_934,N_1101);
nand U2147 (N_2147,N_1335,N_1106);
nand U2148 (N_2148,N_1183,N_1350);
and U2149 (N_2149,N_1222,N_1188);
nor U2150 (N_2150,N_1159,N_912);
and U2151 (N_2151,N_1317,N_1216);
or U2152 (N_2152,N_1171,N_1408);
and U2153 (N_2153,N_928,N_1070);
nand U2154 (N_2154,N_770,N_1337);
and U2155 (N_2155,N_1125,N_1398);
nand U2156 (N_2156,N_1236,N_1099);
nor U2157 (N_2157,N_1499,N_898);
or U2158 (N_2158,N_1238,N_853);
or U2159 (N_2159,N_963,N_1179);
nand U2160 (N_2160,N_1036,N_1082);
and U2161 (N_2161,N_1100,N_1188);
and U2162 (N_2162,N_1117,N_1242);
and U2163 (N_2163,N_995,N_790);
nor U2164 (N_2164,N_1171,N_1212);
and U2165 (N_2165,N_1042,N_934);
or U2166 (N_2166,N_882,N_1212);
nand U2167 (N_2167,N_1022,N_925);
nor U2168 (N_2168,N_1210,N_866);
xor U2169 (N_2169,N_1422,N_1109);
nand U2170 (N_2170,N_825,N_1175);
nor U2171 (N_2171,N_1132,N_1403);
nand U2172 (N_2172,N_1262,N_787);
or U2173 (N_2173,N_1034,N_1078);
nand U2174 (N_2174,N_1172,N_1285);
nand U2175 (N_2175,N_1112,N_1280);
nor U2176 (N_2176,N_759,N_1231);
nor U2177 (N_2177,N_1067,N_1492);
or U2178 (N_2178,N_1332,N_1028);
and U2179 (N_2179,N_1354,N_1430);
and U2180 (N_2180,N_1476,N_1403);
nand U2181 (N_2181,N_1212,N_1179);
nor U2182 (N_2182,N_1470,N_1081);
and U2183 (N_2183,N_1192,N_953);
and U2184 (N_2184,N_1189,N_1403);
or U2185 (N_2185,N_1091,N_1315);
and U2186 (N_2186,N_1332,N_880);
and U2187 (N_2187,N_1243,N_897);
nor U2188 (N_2188,N_1215,N_1041);
nor U2189 (N_2189,N_958,N_901);
and U2190 (N_2190,N_1028,N_1274);
nand U2191 (N_2191,N_1230,N_992);
and U2192 (N_2192,N_1024,N_779);
nor U2193 (N_2193,N_1309,N_842);
nand U2194 (N_2194,N_1309,N_1039);
nand U2195 (N_2195,N_786,N_1135);
nor U2196 (N_2196,N_1141,N_1464);
nor U2197 (N_2197,N_999,N_1039);
nand U2198 (N_2198,N_1156,N_1279);
and U2199 (N_2199,N_1467,N_805);
and U2200 (N_2200,N_1296,N_1337);
nor U2201 (N_2201,N_823,N_1261);
or U2202 (N_2202,N_1484,N_1365);
nor U2203 (N_2203,N_1200,N_1236);
nor U2204 (N_2204,N_957,N_1127);
and U2205 (N_2205,N_943,N_1179);
nor U2206 (N_2206,N_1152,N_867);
or U2207 (N_2207,N_1310,N_1181);
nand U2208 (N_2208,N_1425,N_1217);
or U2209 (N_2209,N_784,N_994);
nor U2210 (N_2210,N_1485,N_1367);
or U2211 (N_2211,N_1059,N_1230);
and U2212 (N_2212,N_1146,N_871);
nor U2213 (N_2213,N_1303,N_886);
and U2214 (N_2214,N_1108,N_1112);
nor U2215 (N_2215,N_1422,N_1391);
nor U2216 (N_2216,N_1321,N_1462);
or U2217 (N_2217,N_1032,N_1026);
nand U2218 (N_2218,N_1404,N_1392);
and U2219 (N_2219,N_1136,N_1377);
and U2220 (N_2220,N_1063,N_1348);
nor U2221 (N_2221,N_1309,N_1222);
or U2222 (N_2222,N_1108,N_1359);
or U2223 (N_2223,N_1259,N_938);
and U2224 (N_2224,N_865,N_1480);
nor U2225 (N_2225,N_1211,N_1344);
nand U2226 (N_2226,N_841,N_1345);
or U2227 (N_2227,N_828,N_1366);
nor U2228 (N_2228,N_952,N_1041);
or U2229 (N_2229,N_1007,N_1069);
nand U2230 (N_2230,N_778,N_1001);
and U2231 (N_2231,N_1322,N_1021);
and U2232 (N_2232,N_1398,N_1310);
nand U2233 (N_2233,N_977,N_1343);
or U2234 (N_2234,N_1128,N_815);
nand U2235 (N_2235,N_1237,N_1024);
or U2236 (N_2236,N_1025,N_983);
and U2237 (N_2237,N_1107,N_1183);
and U2238 (N_2238,N_1452,N_1410);
and U2239 (N_2239,N_1300,N_1028);
nor U2240 (N_2240,N_894,N_1167);
nand U2241 (N_2241,N_1013,N_1361);
or U2242 (N_2242,N_1131,N_1333);
and U2243 (N_2243,N_1484,N_1334);
and U2244 (N_2244,N_1415,N_1405);
or U2245 (N_2245,N_1497,N_1483);
or U2246 (N_2246,N_947,N_932);
or U2247 (N_2247,N_945,N_805);
nor U2248 (N_2248,N_1346,N_786);
xnor U2249 (N_2249,N_1436,N_823);
or U2250 (N_2250,N_1923,N_2020);
nand U2251 (N_2251,N_1704,N_1677);
and U2252 (N_2252,N_1547,N_1861);
nor U2253 (N_2253,N_2104,N_1659);
nand U2254 (N_2254,N_1919,N_1734);
and U2255 (N_2255,N_1959,N_2058);
nand U2256 (N_2256,N_1789,N_2093);
or U2257 (N_2257,N_1618,N_1864);
and U2258 (N_2258,N_1599,N_2076);
or U2259 (N_2259,N_2150,N_2206);
nand U2260 (N_2260,N_2047,N_1961);
or U2261 (N_2261,N_2231,N_2078);
nand U2262 (N_2262,N_1716,N_1684);
nand U2263 (N_2263,N_1715,N_1780);
nor U2264 (N_2264,N_1649,N_1916);
nor U2265 (N_2265,N_1774,N_1543);
nand U2266 (N_2266,N_1823,N_1576);
and U2267 (N_2267,N_1933,N_2062);
nor U2268 (N_2268,N_1759,N_1730);
nor U2269 (N_2269,N_2011,N_1900);
or U2270 (N_2270,N_1676,N_2130);
and U2271 (N_2271,N_2173,N_2181);
and U2272 (N_2272,N_1924,N_2180);
nand U2273 (N_2273,N_2057,N_1697);
and U2274 (N_2274,N_1714,N_2039);
nand U2275 (N_2275,N_1564,N_1891);
nand U2276 (N_2276,N_2029,N_1520);
nor U2277 (N_2277,N_2228,N_1904);
nor U2278 (N_2278,N_1703,N_2131);
and U2279 (N_2279,N_2146,N_2242);
nor U2280 (N_2280,N_1765,N_1633);
or U2281 (N_2281,N_2209,N_2051);
or U2282 (N_2282,N_1687,N_1932);
nand U2283 (N_2283,N_1507,N_2063);
or U2284 (N_2284,N_2036,N_2077);
or U2285 (N_2285,N_2249,N_1748);
nor U2286 (N_2286,N_2100,N_1770);
and U2287 (N_2287,N_1978,N_1808);
nand U2288 (N_2288,N_1784,N_2159);
nor U2289 (N_2289,N_1629,N_2184);
nor U2290 (N_2290,N_1558,N_2061);
or U2291 (N_2291,N_1859,N_1824);
nor U2292 (N_2292,N_1550,N_1971);
and U2293 (N_2293,N_1631,N_1837);
and U2294 (N_2294,N_1614,N_1554);
or U2295 (N_2295,N_2141,N_1605);
nor U2296 (N_2296,N_2232,N_1723);
nor U2297 (N_2297,N_1858,N_1999);
or U2298 (N_2298,N_1525,N_1907);
nand U2299 (N_2299,N_1947,N_1513);
nor U2300 (N_2300,N_1753,N_1918);
nor U2301 (N_2301,N_1777,N_1805);
nand U2302 (N_2302,N_2056,N_2118);
nor U2303 (N_2303,N_1583,N_1533);
nor U2304 (N_2304,N_2119,N_1559);
or U2305 (N_2305,N_1630,N_1580);
nand U2306 (N_2306,N_1701,N_1811);
and U2307 (N_2307,N_1693,N_1601);
or U2308 (N_2308,N_2114,N_1809);
nor U2309 (N_2309,N_2064,N_2136);
and U2310 (N_2310,N_1528,N_1556);
nand U2311 (N_2311,N_1835,N_2230);
and U2312 (N_2312,N_1813,N_1762);
or U2313 (N_2313,N_1840,N_1941);
or U2314 (N_2314,N_2109,N_1851);
nor U2315 (N_2315,N_1839,N_1742);
nor U2316 (N_2316,N_1934,N_2185);
or U2317 (N_2317,N_2144,N_2208);
or U2318 (N_2318,N_1775,N_1983);
nand U2319 (N_2319,N_2154,N_1738);
nand U2320 (N_2320,N_2068,N_2031);
nand U2321 (N_2321,N_2237,N_1761);
or U2322 (N_2322,N_1963,N_1731);
and U2323 (N_2323,N_1820,N_1663);
nor U2324 (N_2324,N_2045,N_2121);
and U2325 (N_2325,N_1910,N_1812);
nand U2326 (N_2326,N_1588,N_2112);
nand U2327 (N_2327,N_1653,N_2129);
nor U2328 (N_2328,N_2215,N_1591);
nor U2329 (N_2329,N_1587,N_1682);
nand U2330 (N_2330,N_2040,N_1966);
or U2331 (N_2331,N_1509,N_2001);
xnor U2332 (N_2332,N_1551,N_2101);
nor U2333 (N_2333,N_1594,N_1893);
or U2334 (N_2334,N_1981,N_1819);
nor U2335 (N_2335,N_1827,N_1897);
nor U2336 (N_2336,N_2070,N_1647);
nor U2337 (N_2337,N_2096,N_1935);
and U2338 (N_2338,N_1740,N_2134);
and U2339 (N_2339,N_1838,N_1561);
or U2340 (N_2340,N_1767,N_1688);
nor U2341 (N_2341,N_1937,N_1913);
or U2342 (N_2342,N_1843,N_2190);
and U2343 (N_2343,N_1706,N_1834);
or U2344 (N_2344,N_1832,N_2165);
nand U2345 (N_2345,N_2082,N_2226);
nand U2346 (N_2346,N_1787,N_2053);
nor U2347 (N_2347,N_1628,N_2167);
and U2348 (N_2348,N_1709,N_1720);
nor U2349 (N_2349,N_1865,N_1725);
nor U2350 (N_2350,N_2140,N_1890);
or U2351 (N_2351,N_1931,N_2059);
or U2352 (N_2352,N_1661,N_1726);
nor U2353 (N_2353,N_1846,N_2193);
nor U2354 (N_2354,N_2103,N_1712);
xor U2355 (N_2355,N_2015,N_2018);
or U2356 (N_2356,N_1721,N_1841);
nand U2357 (N_2357,N_1750,N_1847);
nand U2358 (N_2358,N_1560,N_1566);
nand U2359 (N_2359,N_1786,N_1960);
nand U2360 (N_2360,N_1732,N_1584);
nor U2361 (N_2361,N_1680,N_1648);
nand U2362 (N_2362,N_2002,N_1806);
and U2363 (N_2363,N_1691,N_2128);
nor U2364 (N_2364,N_1878,N_2201);
nand U2365 (N_2365,N_2156,N_1579);
nand U2366 (N_2366,N_1894,N_1848);
and U2367 (N_2367,N_1939,N_1764);
nor U2368 (N_2368,N_2044,N_1517);
or U2369 (N_2369,N_1973,N_2194);
and U2370 (N_2370,N_1545,N_1822);
and U2371 (N_2371,N_2046,N_1796);
and U2372 (N_2372,N_2037,N_1927);
and U2373 (N_2373,N_2160,N_2089);
nand U2374 (N_2374,N_1527,N_2041);
nor U2375 (N_2375,N_1906,N_1968);
and U2376 (N_2376,N_2176,N_1536);
and U2377 (N_2377,N_2217,N_1953);
and U2378 (N_2378,N_2229,N_1756);
or U2379 (N_2379,N_1917,N_1791);
nor U2380 (N_2380,N_1785,N_1850);
and U2381 (N_2381,N_2214,N_1623);
nand U2382 (N_2382,N_1698,N_1657);
and U2383 (N_2383,N_1581,N_2090);
nor U2384 (N_2384,N_2097,N_1853);
nand U2385 (N_2385,N_2221,N_2245);
and U2386 (N_2386,N_2021,N_1674);
nand U2387 (N_2387,N_1728,N_1644);
or U2388 (N_2388,N_2182,N_1825);
nor U2389 (N_2389,N_1793,N_1708);
and U2390 (N_2390,N_1747,N_2205);
and U2391 (N_2391,N_1678,N_2014);
nor U2392 (N_2392,N_1699,N_1922);
and U2393 (N_2393,N_2172,N_1617);
nor U2394 (N_2394,N_2009,N_1634);
or U2395 (N_2395,N_1802,N_1982);
and U2396 (N_2396,N_1842,N_2080);
or U2397 (N_2397,N_1997,N_1673);
or U2398 (N_2398,N_1943,N_1899);
xnor U2399 (N_2399,N_1860,N_1719);
nor U2400 (N_2400,N_2196,N_1537);
nand U2401 (N_2401,N_1570,N_2177);
and U2402 (N_2402,N_2149,N_1951);
nor U2403 (N_2403,N_1988,N_2148);
and U2404 (N_2404,N_1552,N_1669);
and U2405 (N_2405,N_1529,N_2025);
nand U2406 (N_2406,N_1615,N_2017);
nand U2407 (N_2407,N_2162,N_2010);
and U2408 (N_2408,N_1912,N_2246);
xnor U2409 (N_2409,N_1626,N_1553);
and U2410 (N_2410,N_1741,N_2052);
nand U2411 (N_2411,N_2116,N_2042);
nand U2412 (N_2412,N_2235,N_2030);
or U2413 (N_2413,N_1778,N_2222);
nor U2414 (N_2414,N_2098,N_1514);
nor U2415 (N_2415,N_1745,N_1755);
and U2416 (N_2416,N_1586,N_1737);
nand U2417 (N_2417,N_2111,N_2123);
nand U2418 (N_2418,N_1883,N_1672);
nand U2419 (N_2419,N_2024,N_1974);
and U2420 (N_2420,N_1854,N_1915);
nand U2421 (N_2421,N_1585,N_1855);
or U2422 (N_2422,N_2127,N_1751);
or U2423 (N_2423,N_1925,N_1926);
nand U2424 (N_2424,N_1980,N_2079);
and U2425 (N_2425,N_1727,N_1569);
nand U2426 (N_2426,N_1975,N_1690);
nor U2427 (N_2427,N_2092,N_1549);
nand U2428 (N_2428,N_1722,N_1643);
and U2429 (N_2429,N_2216,N_2126);
nand U2430 (N_2430,N_1621,N_1743);
nand U2431 (N_2431,N_2223,N_1944);
nor U2432 (N_2432,N_1606,N_1700);
nand U2433 (N_2433,N_1895,N_1574);
and U2434 (N_2434,N_1871,N_2087);
or U2435 (N_2435,N_1818,N_1531);
nor U2436 (N_2436,N_2213,N_2153);
nor U2437 (N_2437,N_1582,N_2005);
and U2438 (N_2438,N_1689,N_1686);
and U2439 (N_2439,N_1645,N_1639);
or U2440 (N_2440,N_1942,N_2197);
and U2441 (N_2441,N_1636,N_1754);
nand U2442 (N_2442,N_1746,N_1831);
nor U2443 (N_2443,N_1989,N_1870);
and U2444 (N_2444,N_2048,N_2094);
nand U2445 (N_2445,N_2147,N_1646);
and U2446 (N_2446,N_1613,N_2202);
or U2447 (N_2447,N_1996,N_2236);
nor U2448 (N_2448,N_1724,N_1692);
nor U2449 (N_2449,N_1856,N_1874);
and U2450 (N_2450,N_1936,N_2075);
or U2451 (N_2451,N_1664,N_1945);
and U2452 (N_2452,N_1660,N_2050);
nor U2453 (N_2453,N_2085,N_1985);
or U2454 (N_2454,N_1665,N_1521);
and U2455 (N_2455,N_2171,N_1984);
nand U2456 (N_2456,N_1679,N_2241);
nand U2457 (N_2457,N_1972,N_2038);
nor U2458 (N_2458,N_2218,N_1694);
or U2459 (N_2459,N_2027,N_1766);
and U2460 (N_2460,N_2032,N_2195);
nor U2461 (N_2461,N_2207,N_1844);
or U2462 (N_2462,N_1577,N_1530);
nor U2463 (N_2463,N_1501,N_2248);
and U2464 (N_2464,N_1565,N_1651);
or U2465 (N_2465,N_1640,N_2174);
nor U2466 (N_2466,N_1888,N_2161);
and U2467 (N_2467,N_1776,N_1597);
nand U2468 (N_2468,N_1881,N_2233);
and U2469 (N_2469,N_1535,N_1656);
or U2470 (N_2470,N_2212,N_1826);
nand U2471 (N_2471,N_1506,N_1779);
or U2472 (N_2472,N_2105,N_1572);
nor U2473 (N_2473,N_1970,N_1515);
or U2474 (N_2474,N_1901,N_2175);
nor U2475 (N_2475,N_1814,N_2224);
nand U2476 (N_2476,N_1772,N_2168);
or U2477 (N_2477,N_2227,N_1683);
nand U2478 (N_2478,N_1800,N_2091);
nor U2479 (N_2479,N_1799,N_1781);
nand U2480 (N_2480,N_2124,N_1829);
nand U2481 (N_2481,N_1548,N_1713);
and U2482 (N_2482,N_2012,N_1739);
nand U2483 (N_2483,N_2074,N_1769);
nor U2484 (N_2484,N_2151,N_1862);
nand U2485 (N_2485,N_2211,N_1868);
or U2486 (N_2486,N_1782,N_1620);
xor U2487 (N_2487,N_1886,N_1685);
and U2488 (N_2488,N_1675,N_2244);
and U2489 (N_2489,N_2204,N_2135);
or U2490 (N_2490,N_1619,N_1794);
and U2491 (N_2491,N_1598,N_2225);
nand U2492 (N_2492,N_1538,N_2164);
or U2493 (N_2493,N_1804,N_1500);
nand U2494 (N_2494,N_2155,N_1938);
or U2495 (N_2495,N_2139,N_1607);
nand U2496 (N_2496,N_1611,N_1807);
nand U2497 (N_2497,N_2083,N_1578);
or U2498 (N_2498,N_1830,N_1532);
nor U2499 (N_2499,N_1986,N_2188);
nand U2500 (N_2500,N_1892,N_1879);
nand U2501 (N_2501,N_2187,N_1994);
and U2502 (N_2502,N_1872,N_1958);
or U2503 (N_2503,N_1608,N_2192);
or U2504 (N_2504,N_1711,N_1758);
and U2505 (N_2505,N_1662,N_1749);
or U2506 (N_2506,N_1610,N_1705);
and U2507 (N_2507,N_2023,N_1815);
nor U2508 (N_2508,N_2183,N_2071);
nor U2509 (N_2509,N_2219,N_1666);
nor U2510 (N_2510,N_2152,N_2035);
nor U2511 (N_2511,N_1992,N_1519);
xnor U2512 (N_2512,N_1542,N_1696);
and U2513 (N_2513,N_2125,N_1849);
and U2514 (N_2514,N_2170,N_1863);
or U2515 (N_2515,N_1876,N_1757);
or U2516 (N_2516,N_2189,N_2006);
nor U2517 (N_2517,N_1512,N_1949);
or U2518 (N_2518,N_1921,N_1967);
nor U2519 (N_2519,N_2234,N_2138);
nand U2520 (N_2520,N_2106,N_1671);
nor U2521 (N_2521,N_1510,N_2043);
nor U2522 (N_2522,N_1801,N_1718);
nand U2523 (N_2523,N_1555,N_2199);
nand U2524 (N_2524,N_1638,N_1571);
nand U2525 (N_2525,N_2210,N_1568);
and U2526 (N_2526,N_1867,N_2133);
or U2527 (N_2527,N_1768,N_1956);
and U2528 (N_2528,N_1518,N_2069);
nor U2529 (N_2529,N_1710,N_1505);
nand U2530 (N_2530,N_1624,N_2200);
nand U2531 (N_2531,N_1852,N_1788);
or U2532 (N_2532,N_1914,N_1845);
nand U2533 (N_2533,N_1695,N_1828);
and U2534 (N_2534,N_1652,N_1817);
or U2535 (N_2535,N_1744,N_1504);
or U2536 (N_2536,N_1522,N_1523);
nand U2537 (N_2537,N_2084,N_1733);
nor U2538 (N_2538,N_2003,N_1987);
and U2539 (N_2539,N_2072,N_2060);
or U2540 (N_2540,N_1625,N_1516);
or U2541 (N_2541,N_1736,N_1962);
or U2542 (N_2542,N_2115,N_2137);
nand U2543 (N_2543,N_1979,N_1905);
nor U2544 (N_2544,N_1763,N_1946);
nand U2545 (N_2545,N_1790,N_1642);
or U2546 (N_2546,N_1795,N_1908);
nand U2547 (N_2547,N_2086,N_1909);
nand U2548 (N_2548,N_2247,N_2198);
or U2549 (N_2549,N_2004,N_1540);
nor U2550 (N_2550,N_1600,N_1637);
nand U2551 (N_2551,N_1735,N_1627);
and U2552 (N_2552,N_1882,N_2007);
nand U2553 (N_2553,N_1575,N_1641);
and U2554 (N_2554,N_1590,N_1792);
or U2555 (N_2555,N_1650,N_2026);
or U2556 (N_2556,N_1898,N_2120);
nand U2557 (N_2557,N_1596,N_1667);
nand U2558 (N_2558,N_2220,N_1612);
nand U2559 (N_2559,N_1632,N_2067);
nor U2560 (N_2560,N_1911,N_1873);
nand U2561 (N_2561,N_1573,N_1903);
nand U2562 (N_2562,N_1503,N_2107);
nor U2563 (N_2563,N_1998,N_1885);
and U2564 (N_2564,N_2122,N_1880);
nor U2565 (N_2565,N_1977,N_1681);
and U2566 (N_2566,N_2008,N_1592);
and U2567 (N_2567,N_2113,N_1810);
nor U2568 (N_2568,N_1976,N_1995);
and U2569 (N_2569,N_1544,N_2019);
nor U2570 (N_2570,N_1508,N_1821);
and U2571 (N_2571,N_2033,N_1920);
and U2572 (N_2572,N_2166,N_1866);
or U2573 (N_2573,N_1557,N_1887);
nor U2574 (N_2574,N_1950,N_1589);
nor U2575 (N_2575,N_1511,N_2158);
or U2576 (N_2576,N_1954,N_1797);
nor U2577 (N_2577,N_1869,N_1524);
nor U2578 (N_2578,N_1990,N_1833);
or U2579 (N_2579,N_2049,N_1526);
or U2580 (N_2580,N_2191,N_1670);
and U2581 (N_2581,N_1896,N_1803);
nor U2582 (N_2582,N_1609,N_1604);
nor U2583 (N_2583,N_1539,N_1729);
or U2584 (N_2584,N_1616,N_1567);
and U2585 (N_2585,N_1964,N_1702);
and U2586 (N_2586,N_1857,N_1595);
nand U2587 (N_2587,N_2117,N_1993);
and U2588 (N_2588,N_1889,N_1534);
or U2589 (N_2589,N_1654,N_2243);
or U2590 (N_2590,N_1760,N_1798);
or U2591 (N_2591,N_2132,N_2099);
or U2592 (N_2592,N_2088,N_2095);
and U2593 (N_2593,N_1752,N_2110);
nand U2594 (N_2594,N_1603,N_1717);
and U2595 (N_2595,N_2145,N_1658);
and U2596 (N_2596,N_1875,N_2179);
nand U2597 (N_2597,N_2054,N_2066);
or U2598 (N_2598,N_2203,N_2186);
or U2599 (N_2599,N_2055,N_2073);
nand U2600 (N_2600,N_1655,N_1902);
and U2601 (N_2601,N_1562,N_2081);
nor U2602 (N_2602,N_1816,N_1965);
nor U2603 (N_2603,N_1541,N_1930);
nor U2604 (N_2604,N_1593,N_2240);
nand U2605 (N_2605,N_2016,N_1502);
or U2606 (N_2606,N_2000,N_2163);
nand U2607 (N_2607,N_2238,N_1948);
and U2608 (N_2608,N_1929,N_1957);
nand U2609 (N_2609,N_1940,N_2108);
nand U2610 (N_2610,N_2034,N_2013);
nor U2611 (N_2611,N_1563,N_1546);
or U2612 (N_2612,N_1884,N_2239);
nand U2613 (N_2613,N_2143,N_1707);
nor U2614 (N_2614,N_1602,N_2142);
or U2615 (N_2615,N_2157,N_1668);
nand U2616 (N_2616,N_1928,N_1877);
nand U2617 (N_2617,N_1836,N_2065);
and U2618 (N_2618,N_1771,N_2028);
and U2619 (N_2619,N_1991,N_1635);
nand U2620 (N_2620,N_1952,N_1955);
or U2621 (N_2621,N_1622,N_2169);
and U2622 (N_2622,N_1783,N_1969);
or U2623 (N_2623,N_2102,N_2178);
and U2624 (N_2624,N_2022,N_1773);
or U2625 (N_2625,N_2013,N_1954);
nand U2626 (N_2626,N_1698,N_2146);
or U2627 (N_2627,N_2095,N_2045);
or U2628 (N_2628,N_2153,N_2247);
or U2629 (N_2629,N_2055,N_1852);
and U2630 (N_2630,N_1504,N_1651);
and U2631 (N_2631,N_1799,N_1612);
and U2632 (N_2632,N_1688,N_1916);
and U2633 (N_2633,N_2105,N_1938);
and U2634 (N_2634,N_1987,N_1826);
or U2635 (N_2635,N_2052,N_1539);
and U2636 (N_2636,N_1722,N_1928);
and U2637 (N_2637,N_2054,N_1683);
nand U2638 (N_2638,N_1502,N_2033);
nor U2639 (N_2639,N_2219,N_2203);
and U2640 (N_2640,N_1801,N_1677);
nand U2641 (N_2641,N_2239,N_1980);
and U2642 (N_2642,N_2155,N_1927);
nand U2643 (N_2643,N_1870,N_1771);
and U2644 (N_2644,N_1560,N_1642);
or U2645 (N_2645,N_1600,N_1516);
nor U2646 (N_2646,N_1846,N_2004);
and U2647 (N_2647,N_1643,N_1538);
nand U2648 (N_2648,N_1544,N_1905);
nand U2649 (N_2649,N_2100,N_1521);
nor U2650 (N_2650,N_2008,N_2063);
and U2651 (N_2651,N_1528,N_1580);
and U2652 (N_2652,N_2248,N_1739);
nor U2653 (N_2653,N_1736,N_1894);
nor U2654 (N_2654,N_1767,N_1655);
or U2655 (N_2655,N_1637,N_1525);
nand U2656 (N_2656,N_1871,N_1632);
nand U2657 (N_2657,N_1628,N_2191);
and U2658 (N_2658,N_1830,N_1832);
and U2659 (N_2659,N_2230,N_1534);
nor U2660 (N_2660,N_1993,N_1834);
nand U2661 (N_2661,N_2057,N_1612);
nand U2662 (N_2662,N_1703,N_1561);
or U2663 (N_2663,N_1940,N_1766);
nor U2664 (N_2664,N_1964,N_1910);
or U2665 (N_2665,N_2107,N_1685);
nor U2666 (N_2666,N_1964,N_1735);
or U2667 (N_2667,N_2216,N_2120);
nand U2668 (N_2668,N_2032,N_1520);
nor U2669 (N_2669,N_2100,N_1999);
nand U2670 (N_2670,N_1940,N_1977);
nand U2671 (N_2671,N_2208,N_2137);
nand U2672 (N_2672,N_1723,N_1604);
and U2673 (N_2673,N_1901,N_1674);
or U2674 (N_2674,N_1874,N_1625);
nand U2675 (N_2675,N_1731,N_2083);
or U2676 (N_2676,N_1607,N_1762);
and U2677 (N_2677,N_2044,N_1667);
xor U2678 (N_2678,N_1612,N_2204);
xor U2679 (N_2679,N_2103,N_1845);
and U2680 (N_2680,N_2203,N_1703);
or U2681 (N_2681,N_1723,N_1571);
and U2682 (N_2682,N_1652,N_1529);
nand U2683 (N_2683,N_2106,N_1540);
or U2684 (N_2684,N_2047,N_1622);
and U2685 (N_2685,N_1955,N_1659);
nand U2686 (N_2686,N_1860,N_2026);
or U2687 (N_2687,N_1817,N_2114);
xnor U2688 (N_2688,N_1957,N_1946);
nand U2689 (N_2689,N_1841,N_1842);
nand U2690 (N_2690,N_1777,N_1719);
and U2691 (N_2691,N_2224,N_1601);
or U2692 (N_2692,N_2041,N_2224);
and U2693 (N_2693,N_1826,N_1905);
nor U2694 (N_2694,N_1913,N_1807);
or U2695 (N_2695,N_1565,N_2019);
nand U2696 (N_2696,N_1940,N_2021);
nand U2697 (N_2697,N_1805,N_1669);
nor U2698 (N_2698,N_2115,N_1705);
nor U2699 (N_2699,N_2208,N_2212);
and U2700 (N_2700,N_1726,N_2090);
and U2701 (N_2701,N_1702,N_1752);
nor U2702 (N_2702,N_1871,N_1691);
nor U2703 (N_2703,N_2131,N_2188);
and U2704 (N_2704,N_1668,N_2189);
or U2705 (N_2705,N_1755,N_1738);
nor U2706 (N_2706,N_2021,N_1562);
and U2707 (N_2707,N_1551,N_1788);
and U2708 (N_2708,N_1712,N_2086);
nand U2709 (N_2709,N_1727,N_2025);
nor U2710 (N_2710,N_1636,N_1697);
nor U2711 (N_2711,N_2060,N_2053);
nor U2712 (N_2712,N_2184,N_1983);
nand U2713 (N_2713,N_1889,N_1977);
or U2714 (N_2714,N_1732,N_2193);
nor U2715 (N_2715,N_1714,N_1751);
nor U2716 (N_2716,N_1864,N_2190);
xnor U2717 (N_2717,N_2232,N_1711);
and U2718 (N_2718,N_2197,N_1857);
and U2719 (N_2719,N_1794,N_1545);
and U2720 (N_2720,N_1569,N_1696);
or U2721 (N_2721,N_2116,N_1984);
nor U2722 (N_2722,N_1529,N_1671);
or U2723 (N_2723,N_1519,N_1568);
nand U2724 (N_2724,N_2150,N_1837);
nand U2725 (N_2725,N_1937,N_1876);
nor U2726 (N_2726,N_1996,N_1766);
nor U2727 (N_2727,N_1579,N_1537);
nor U2728 (N_2728,N_2022,N_1995);
nor U2729 (N_2729,N_1562,N_2235);
or U2730 (N_2730,N_2132,N_1619);
and U2731 (N_2731,N_1748,N_2051);
or U2732 (N_2732,N_1862,N_1915);
or U2733 (N_2733,N_1566,N_1612);
xor U2734 (N_2734,N_1677,N_1837);
nand U2735 (N_2735,N_2027,N_2087);
or U2736 (N_2736,N_2141,N_2012);
and U2737 (N_2737,N_1897,N_2053);
or U2738 (N_2738,N_1873,N_1642);
nand U2739 (N_2739,N_2147,N_1982);
nor U2740 (N_2740,N_1590,N_2146);
or U2741 (N_2741,N_2181,N_2184);
nand U2742 (N_2742,N_1754,N_1911);
or U2743 (N_2743,N_1565,N_1753);
and U2744 (N_2744,N_1968,N_2072);
nand U2745 (N_2745,N_1867,N_1952);
or U2746 (N_2746,N_1757,N_2156);
nor U2747 (N_2747,N_1708,N_1545);
or U2748 (N_2748,N_2108,N_1677);
nor U2749 (N_2749,N_1735,N_1803);
nand U2750 (N_2750,N_1673,N_2237);
nand U2751 (N_2751,N_1767,N_1648);
nor U2752 (N_2752,N_2035,N_1869);
nor U2753 (N_2753,N_1854,N_2212);
or U2754 (N_2754,N_1937,N_2056);
nor U2755 (N_2755,N_2053,N_1813);
and U2756 (N_2756,N_1539,N_2045);
or U2757 (N_2757,N_2030,N_1862);
or U2758 (N_2758,N_1544,N_2036);
or U2759 (N_2759,N_2081,N_1640);
and U2760 (N_2760,N_1534,N_1765);
or U2761 (N_2761,N_1946,N_2011);
or U2762 (N_2762,N_1836,N_1530);
nand U2763 (N_2763,N_2108,N_2194);
and U2764 (N_2764,N_1848,N_1621);
or U2765 (N_2765,N_1822,N_1769);
nor U2766 (N_2766,N_2105,N_1700);
or U2767 (N_2767,N_1673,N_1565);
nor U2768 (N_2768,N_1777,N_1641);
nor U2769 (N_2769,N_1770,N_2095);
or U2770 (N_2770,N_2223,N_1507);
or U2771 (N_2771,N_2121,N_2148);
nor U2772 (N_2772,N_2134,N_1842);
nor U2773 (N_2773,N_1726,N_1568);
or U2774 (N_2774,N_1958,N_1731);
nor U2775 (N_2775,N_1651,N_1763);
nor U2776 (N_2776,N_1659,N_1595);
or U2777 (N_2777,N_2164,N_2171);
or U2778 (N_2778,N_2173,N_1678);
or U2779 (N_2779,N_1700,N_1772);
or U2780 (N_2780,N_2052,N_1987);
nor U2781 (N_2781,N_1594,N_1829);
nor U2782 (N_2782,N_2118,N_1860);
or U2783 (N_2783,N_2236,N_2103);
and U2784 (N_2784,N_1527,N_1907);
and U2785 (N_2785,N_2128,N_1507);
and U2786 (N_2786,N_1876,N_1769);
xnor U2787 (N_2787,N_2148,N_1667);
and U2788 (N_2788,N_2178,N_1857);
nor U2789 (N_2789,N_1773,N_1734);
or U2790 (N_2790,N_1846,N_1997);
and U2791 (N_2791,N_1729,N_1688);
nor U2792 (N_2792,N_2162,N_1714);
nor U2793 (N_2793,N_1968,N_2039);
nand U2794 (N_2794,N_1515,N_1881);
or U2795 (N_2795,N_2006,N_1733);
or U2796 (N_2796,N_1515,N_1935);
nor U2797 (N_2797,N_1847,N_2229);
nand U2798 (N_2798,N_1747,N_1655);
and U2799 (N_2799,N_1915,N_1614);
or U2800 (N_2800,N_1946,N_2140);
or U2801 (N_2801,N_2052,N_1646);
and U2802 (N_2802,N_1762,N_1982);
and U2803 (N_2803,N_2149,N_2199);
and U2804 (N_2804,N_1963,N_1504);
or U2805 (N_2805,N_2233,N_1681);
and U2806 (N_2806,N_1997,N_1566);
or U2807 (N_2807,N_2040,N_2025);
nand U2808 (N_2808,N_1741,N_2094);
or U2809 (N_2809,N_1795,N_2210);
nor U2810 (N_2810,N_1836,N_1759);
nand U2811 (N_2811,N_1539,N_1661);
nand U2812 (N_2812,N_2025,N_2049);
or U2813 (N_2813,N_1682,N_2183);
and U2814 (N_2814,N_1550,N_1997);
and U2815 (N_2815,N_1651,N_1935);
and U2816 (N_2816,N_1962,N_1805);
nand U2817 (N_2817,N_1814,N_1658);
and U2818 (N_2818,N_2055,N_1798);
nand U2819 (N_2819,N_2175,N_2008);
or U2820 (N_2820,N_1763,N_1980);
and U2821 (N_2821,N_2153,N_1660);
nand U2822 (N_2822,N_1758,N_1786);
nand U2823 (N_2823,N_1914,N_1771);
nand U2824 (N_2824,N_1790,N_1972);
nor U2825 (N_2825,N_1684,N_1807);
and U2826 (N_2826,N_1628,N_1743);
and U2827 (N_2827,N_1625,N_1641);
nor U2828 (N_2828,N_2233,N_1588);
and U2829 (N_2829,N_1907,N_1928);
or U2830 (N_2830,N_2012,N_2171);
nand U2831 (N_2831,N_2185,N_2214);
and U2832 (N_2832,N_1966,N_1742);
or U2833 (N_2833,N_2133,N_1544);
and U2834 (N_2834,N_1922,N_1688);
and U2835 (N_2835,N_1555,N_1733);
and U2836 (N_2836,N_1790,N_2181);
nor U2837 (N_2837,N_2179,N_1721);
nor U2838 (N_2838,N_1654,N_2239);
or U2839 (N_2839,N_1652,N_1767);
nor U2840 (N_2840,N_2018,N_1541);
nor U2841 (N_2841,N_1669,N_2169);
and U2842 (N_2842,N_2161,N_1608);
or U2843 (N_2843,N_1855,N_1801);
or U2844 (N_2844,N_2041,N_1805);
or U2845 (N_2845,N_1832,N_2180);
nor U2846 (N_2846,N_1950,N_1541);
or U2847 (N_2847,N_1804,N_1700);
and U2848 (N_2848,N_2240,N_1993);
nand U2849 (N_2849,N_1974,N_2020);
nor U2850 (N_2850,N_1915,N_1684);
nor U2851 (N_2851,N_2180,N_1508);
nand U2852 (N_2852,N_2098,N_1872);
nand U2853 (N_2853,N_1918,N_1869);
nand U2854 (N_2854,N_2045,N_2081);
or U2855 (N_2855,N_2036,N_2140);
or U2856 (N_2856,N_2015,N_1687);
or U2857 (N_2857,N_2138,N_2060);
nor U2858 (N_2858,N_2093,N_1506);
and U2859 (N_2859,N_2158,N_2144);
nand U2860 (N_2860,N_1997,N_1919);
nand U2861 (N_2861,N_1667,N_1548);
and U2862 (N_2862,N_1779,N_1856);
nor U2863 (N_2863,N_2229,N_1944);
nand U2864 (N_2864,N_2226,N_1837);
nand U2865 (N_2865,N_1951,N_1748);
nor U2866 (N_2866,N_2228,N_1984);
nor U2867 (N_2867,N_1823,N_1651);
or U2868 (N_2868,N_1931,N_2247);
nand U2869 (N_2869,N_2240,N_2144);
and U2870 (N_2870,N_1776,N_1540);
nand U2871 (N_2871,N_1939,N_2035);
and U2872 (N_2872,N_2049,N_2159);
or U2873 (N_2873,N_1716,N_1599);
or U2874 (N_2874,N_1862,N_1557);
or U2875 (N_2875,N_1932,N_1698);
and U2876 (N_2876,N_1527,N_1603);
nand U2877 (N_2877,N_1868,N_1965);
or U2878 (N_2878,N_2152,N_1702);
and U2879 (N_2879,N_1579,N_1654);
or U2880 (N_2880,N_1537,N_1534);
or U2881 (N_2881,N_1850,N_2188);
or U2882 (N_2882,N_1711,N_1660);
nand U2883 (N_2883,N_1656,N_1899);
or U2884 (N_2884,N_1662,N_2080);
nand U2885 (N_2885,N_1555,N_2097);
nand U2886 (N_2886,N_1897,N_1752);
nor U2887 (N_2887,N_1742,N_2069);
or U2888 (N_2888,N_1611,N_2034);
or U2889 (N_2889,N_1756,N_1818);
nand U2890 (N_2890,N_1778,N_2164);
nor U2891 (N_2891,N_1565,N_1648);
nor U2892 (N_2892,N_1685,N_2135);
or U2893 (N_2893,N_1558,N_1783);
and U2894 (N_2894,N_2044,N_1942);
nor U2895 (N_2895,N_1975,N_2131);
or U2896 (N_2896,N_1510,N_1550);
nor U2897 (N_2897,N_2148,N_1803);
nor U2898 (N_2898,N_1873,N_1788);
and U2899 (N_2899,N_1826,N_1859);
nand U2900 (N_2900,N_1983,N_1788);
nor U2901 (N_2901,N_2245,N_1937);
nand U2902 (N_2902,N_1987,N_2132);
nand U2903 (N_2903,N_2054,N_2018);
nor U2904 (N_2904,N_1596,N_1920);
nor U2905 (N_2905,N_2093,N_1905);
xnor U2906 (N_2906,N_2188,N_1749);
or U2907 (N_2907,N_2125,N_1939);
nand U2908 (N_2908,N_1922,N_2092);
and U2909 (N_2909,N_2095,N_1917);
or U2910 (N_2910,N_1954,N_2176);
nor U2911 (N_2911,N_2164,N_2026);
and U2912 (N_2912,N_1854,N_2203);
nor U2913 (N_2913,N_1526,N_2060);
nand U2914 (N_2914,N_1869,N_1981);
or U2915 (N_2915,N_2213,N_2174);
nand U2916 (N_2916,N_1570,N_1940);
and U2917 (N_2917,N_1971,N_2155);
or U2918 (N_2918,N_2040,N_2143);
nand U2919 (N_2919,N_1527,N_2058);
and U2920 (N_2920,N_1951,N_1783);
and U2921 (N_2921,N_1664,N_1683);
nand U2922 (N_2922,N_1719,N_1776);
and U2923 (N_2923,N_1523,N_1869);
and U2924 (N_2924,N_1838,N_1604);
nand U2925 (N_2925,N_1541,N_2188);
and U2926 (N_2926,N_1895,N_2055);
or U2927 (N_2927,N_1828,N_1764);
nand U2928 (N_2928,N_2193,N_2068);
nor U2929 (N_2929,N_2008,N_1842);
nand U2930 (N_2930,N_2179,N_1555);
nand U2931 (N_2931,N_1900,N_2159);
or U2932 (N_2932,N_1630,N_1878);
or U2933 (N_2933,N_2058,N_1931);
or U2934 (N_2934,N_1722,N_1511);
nand U2935 (N_2935,N_1769,N_1863);
and U2936 (N_2936,N_1540,N_1977);
and U2937 (N_2937,N_1979,N_2107);
or U2938 (N_2938,N_1646,N_1500);
or U2939 (N_2939,N_2004,N_2177);
or U2940 (N_2940,N_1812,N_1803);
nor U2941 (N_2941,N_2003,N_2155);
nand U2942 (N_2942,N_2042,N_1670);
or U2943 (N_2943,N_1605,N_2167);
or U2944 (N_2944,N_2119,N_1671);
and U2945 (N_2945,N_1828,N_2009);
nor U2946 (N_2946,N_1836,N_2145);
and U2947 (N_2947,N_1873,N_1714);
or U2948 (N_2948,N_2195,N_1659);
and U2949 (N_2949,N_2041,N_1515);
and U2950 (N_2950,N_2009,N_2143);
nand U2951 (N_2951,N_1661,N_2133);
nor U2952 (N_2952,N_1684,N_2087);
nor U2953 (N_2953,N_1775,N_2067);
nor U2954 (N_2954,N_1837,N_1950);
or U2955 (N_2955,N_2007,N_2040);
nand U2956 (N_2956,N_2107,N_1549);
nand U2957 (N_2957,N_1862,N_1839);
nand U2958 (N_2958,N_2246,N_1505);
and U2959 (N_2959,N_1847,N_1698);
and U2960 (N_2960,N_2187,N_2188);
or U2961 (N_2961,N_1962,N_2230);
nor U2962 (N_2962,N_1865,N_1545);
nand U2963 (N_2963,N_1943,N_2180);
nor U2964 (N_2964,N_1936,N_2086);
nor U2965 (N_2965,N_2076,N_1877);
or U2966 (N_2966,N_1624,N_2064);
nand U2967 (N_2967,N_1690,N_2064);
nor U2968 (N_2968,N_2044,N_1924);
nand U2969 (N_2969,N_1708,N_1711);
nor U2970 (N_2970,N_1737,N_1961);
nor U2971 (N_2971,N_2181,N_2089);
and U2972 (N_2972,N_1989,N_1902);
and U2973 (N_2973,N_1752,N_2207);
nand U2974 (N_2974,N_2186,N_2120);
nand U2975 (N_2975,N_2227,N_1777);
and U2976 (N_2976,N_2118,N_1848);
nand U2977 (N_2977,N_2068,N_2120);
nor U2978 (N_2978,N_2187,N_1756);
nor U2979 (N_2979,N_2060,N_2010);
nor U2980 (N_2980,N_2003,N_2032);
nand U2981 (N_2981,N_1653,N_1721);
nand U2982 (N_2982,N_1917,N_2032);
nand U2983 (N_2983,N_2122,N_1996);
or U2984 (N_2984,N_2085,N_1997);
or U2985 (N_2985,N_1926,N_1842);
xnor U2986 (N_2986,N_2038,N_1914);
nand U2987 (N_2987,N_1978,N_1560);
nand U2988 (N_2988,N_1684,N_2093);
or U2989 (N_2989,N_1560,N_1969);
and U2990 (N_2990,N_1715,N_1921);
nand U2991 (N_2991,N_1720,N_2072);
or U2992 (N_2992,N_1905,N_1879);
or U2993 (N_2993,N_1508,N_2060);
or U2994 (N_2994,N_1949,N_1988);
nand U2995 (N_2995,N_1987,N_2217);
nor U2996 (N_2996,N_2237,N_2131);
nor U2997 (N_2997,N_1771,N_1625);
or U2998 (N_2998,N_1505,N_1649);
or U2999 (N_2999,N_1749,N_1532);
nand U3000 (N_3000,N_2642,N_2397);
nor U3001 (N_3001,N_2437,N_2580);
and U3002 (N_3002,N_2393,N_2812);
nand U3003 (N_3003,N_2528,N_2276);
nor U3004 (N_3004,N_2763,N_2932);
nor U3005 (N_3005,N_2966,N_2895);
or U3006 (N_3006,N_2367,N_2949);
nand U3007 (N_3007,N_2554,N_2770);
nor U3008 (N_3008,N_2680,N_2700);
or U3009 (N_3009,N_2382,N_2446);
nor U3010 (N_3010,N_2352,N_2704);
or U3011 (N_3011,N_2284,N_2725);
nor U3012 (N_3012,N_2432,N_2458);
or U3013 (N_3013,N_2481,N_2830);
nor U3014 (N_3014,N_2594,N_2761);
or U3015 (N_3015,N_2597,N_2961);
nor U3016 (N_3016,N_2869,N_2493);
nand U3017 (N_3017,N_2614,N_2996);
nor U3018 (N_3018,N_2719,N_2428);
or U3019 (N_3019,N_2688,N_2671);
nor U3020 (N_3020,N_2933,N_2484);
and U3021 (N_3021,N_2709,N_2308);
nor U3022 (N_3022,N_2569,N_2563);
and U3023 (N_3023,N_2997,N_2400);
nand U3024 (N_3024,N_2645,N_2426);
or U3025 (N_3025,N_2943,N_2486);
nor U3026 (N_3026,N_2867,N_2390);
nand U3027 (N_3027,N_2937,N_2440);
or U3028 (N_3028,N_2621,N_2553);
nor U3029 (N_3029,N_2463,N_2386);
nand U3030 (N_3030,N_2275,N_2282);
and U3031 (N_3031,N_2847,N_2336);
and U3032 (N_3032,N_2615,N_2695);
and U3033 (N_3033,N_2376,N_2502);
or U3034 (N_3034,N_2514,N_2371);
or U3035 (N_3035,N_2547,N_2473);
nor U3036 (N_3036,N_2756,N_2622);
or U3037 (N_3037,N_2431,N_2441);
or U3038 (N_3038,N_2470,N_2329);
or U3039 (N_3039,N_2721,N_2824);
nand U3040 (N_3040,N_2968,N_2505);
and U3041 (N_3041,N_2658,N_2504);
nand U3042 (N_3042,N_2288,N_2909);
or U3043 (N_3043,N_2723,N_2457);
nand U3044 (N_3044,N_2634,N_2627);
nor U3045 (N_3045,N_2903,N_2277);
or U3046 (N_3046,N_2900,N_2586);
and U3047 (N_3047,N_2632,N_2734);
xor U3048 (N_3048,N_2380,N_2831);
and U3049 (N_3049,N_2482,N_2777);
and U3050 (N_3050,N_2731,N_2808);
or U3051 (N_3051,N_2445,N_2970);
nor U3052 (N_3052,N_2814,N_2990);
or U3053 (N_3053,N_2999,N_2471);
nor U3054 (N_3054,N_2507,N_2617);
nor U3055 (N_3055,N_2759,N_2938);
nor U3056 (N_3056,N_2822,N_2994);
nor U3057 (N_3057,N_2844,N_2414);
nand U3058 (N_3058,N_2604,N_2885);
or U3059 (N_3059,N_2828,N_2792);
or U3060 (N_3060,N_2332,N_2760);
and U3061 (N_3061,N_2601,N_2785);
and U3062 (N_3062,N_2716,N_2732);
and U3063 (N_3063,N_2897,N_2356);
nand U3064 (N_3064,N_2550,N_2372);
or U3065 (N_3065,N_2772,N_2341);
or U3066 (N_3066,N_2442,N_2941);
or U3067 (N_3067,N_2268,N_2264);
nor U3068 (N_3068,N_2764,N_2659);
nor U3069 (N_3069,N_2748,N_2524);
and U3070 (N_3070,N_2637,N_2730);
and U3071 (N_3071,N_2720,N_2931);
nand U3072 (N_3072,N_2703,N_2889);
and U3073 (N_3073,N_2269,N_2670);
or U3074 (N_3074,N_2453,N_2657);
or U3075 (N_3075,N_2892,N_2508);
and U3076 (N_3076,N_2790,N_2874);
or U3077 (N_3077,N_2684,N_2973);
nor U3078 (N_3078,N_2599,N_2667);
and U3079 (N_3079,N_2404,N_2510);
or U3080 (N_3080,N_2354,N_2965);
and U3081 (N_3081,N_2837,N_2656);
nor U3082 (N_3082,N_2767,N_2575);
or U3083 (N_3083,N_2856,N_2836);
and U3084 (N_3084,N_2364,N_2727);
nor U3085 (N_3085,N_2906,N_2689);
and U3086 (N_3086,N_2713,N_2302);
nor U3087 (N_3087,N_2497,N_2363);
nand U3088 (N_3088,N_2663,N_2698);
and U3089 (N_3089,N_2461,N_2818);
and U3090 (N_3090,N_2624,N_2494);
or U3091 (N_3091,N_2829,N_2773);
and U3092 (N_3092,N_2564,N_2983);
xor U3093 (N_3093,N_2595,N_2786);
and U3094 (N_3094,N_2464,N_2883);
nor U3095 (N_3095,N_2537,N_2304);
or U3096 (N_3096,N_2661,N_2876);
nor U3097 (N_3097,N_2384,N_2751);
nor U3098 (N_3098,N_2291,N_2718);
nand U3099 (N_3099,N_2693,N_2349);
nand U3100 (N_3100,N_2333,N_2838);
nand U3101 (N_3101,N_2603,N_2289);
or U3102 (N_3102,N_2697,N_2478);
or U3103 (N_3103,N_2678,N_2285);
and U3104 (N_3104,N_2823,N_2607);
or U3105 (N_3105,N_2496,N_2520);
or U3106 (N_3106,N_2472,N_2981);
and U3107 (N_3107,N_2303,N_2944);
nand U3108 (N_3108,N_2438,N_2577);
nand U3109 (N_3109,N_2585,N_2287);
nand U3110 (N_3110,N_2758,N_2745);
nor U3111 (N_3111,N_2958,N_2884);
nor U3112 (N_3112,N_2369,N_2702);
or U3113 (N_3113,N_2503,N_2561);
or U3114 (N_3114,N_2439,N_2640);
nor U3115 (N_3115,N_2253,N_2323);
or U3116 (N_3116,N_2858,N_2696);
or U3117 (N_3117,N_2715,N_2297);
nor U3118 (N_3118,N_2655,N_2930);
or U3119 (N_3119,N_2406,N_2747);
or U3120 (N_3120,N_2392,N_2705);
xnor U3121 (N_3121,N_2257,N_2669);
nand U3122 (N_3122,N_2330,N_2972);
or U3123 (N_3123,N_2467,N_2851);
or U3124 (N_3124,N_2648,N_2625);
or U3125 (N_3125,N_2988,N_2784);
or U3126 (N_3126,N_2879,N_2572);
or U3127 (N_3127,N_2489,N_2396);
and U3128 (N_3128,N_2600,N_2950);
nor U3129 (N_3129,N_2629,N_2827);
nor U3130 (N_3130,N_2385,N_2525);
and U3131 (N_3131,N_2281,N_2339);
and U3132 (N_3132,N_2992,N_2807);
nand U3133 (N_3133,N_2509,N_2421);
nand U3134 (N_3134,N_2989,N_2571);
nor U3135 (N_3135,N_2861,N_2279);
nand U3136 (N_3136,N_2724,N_2845);
nor U3137 (N_3137,N_2608,N_2865);
and U3138 (N_3138,N_2312,N_2955);
or U3139 (N_3139,N_2616,N_2351);
nand U3140 (N_3140,N_2910,N_2849);
and U3141 (N_3141,N_2299,N_2839);
nand U3142 (N_3142,N_2868,N_2541);
nand U3143 (N_3143,N_2819,N_2915);
nand U3144 (N_3144,N_2841,N_2305);
or U3145 (N_3145,N_2899,N_2956);
nand U3146 (N_3146,N_2840,N_2511);
or U3147 (N_3147,N_2787,N_2320);
or U3148 (N_3148,N_2630,N_2982);
and U3149 (N_3149,N_2871,N_2775);
nand U3150 (N_3150,N_2523,N_2654);
or U3151 (N_3151,N_2602,N_2945);
and U3152 (N_3152,N_2912,N_2324);
and U3153 (N_3153,N_2412,N_2391);
nand U3154 (N_3154,N_2902,N_2638);
and U3155 (N_3155,N_2605,N_2581);
and U3156 (N_3156,N_2480,N_2898);
nand U3157 (N_3157,N_2863,N_2250);
nor U3158 (N_3158,N_2801,N_2576);
nor U3159 (N_3159,N_2306,N_2820);
nand U3160 (N_3160,N_2410,N_2971);
nand U3161 (N_3161,N_2984,N_2368);
xnor U3162 (N_3162,N_2854,N_2596);
or U3163 (N_3163,N_2610,N_2833);
and U3164 (N_3164,N_2987,N_2766);
nor U3165 (N_3165,N_2474,N_2832);
nor U3166 (N_3166,N_2907,N_2942);
nor U3167 (N_3167,N_2318,N_2717);
nor U3168 (N_3168,N_2534,N_2298);
or U3169 (N_3169,N_2701,N_2444);
nand U3170 (N_3170,N_2813,N_2325);
nand U3171 (N_3171,N_2462,N_2940);
and U3172 (N_3172,N_2405,N_2797);
or U3173 (N_3173,N_2952,N_2455);
nand U3174 (N_3174,N_2925,N_2749);
and U3175 (N_3175,N_2890,N_2682);
and U3176 (N_3176,N_2995,N_2559);
nor U3177 (N_3177,N_2451,N_2527);
and U3178 (N_3178,N_2694,N_2460);
or U3179 (N_3179,N_2935,N_2360);
or U3180 (N_3180,N_2450,N_2652);
or U3181 (N_3181,N_2789,N_2321);
or U3182 (N_3182,N_2769,N_2755);
nor U3183 (N_3183,N_2788,N_2567);
and U3184 (N_3184,N_2492,N_2345);
xnor U3185 (N_3185,N_2980,N_2864);
nand U3186 (N_3186,N_2799,N_2293);
nor U3187 (N_3187,N_2531,N_2860);
or U3188 (N_3188,N_2469,N_2370);
or U3189 (N_3189,N_2389,N_2737);
nand U3190 (N_3190,N_2315,N_2562);
nand U3191 (N_3191,N_2733,N_2641);
nand U3192 (N_3192,N_2795,N_2873);
nor U3193 (N_3193,N_2353,N_2378);
nor U3194 (N_3194,N_2835,N_2476);
nor U3195 (N_3195,N_2948,N_2639);
and U3196 (N_3196,N_2361,N_2373);
nand U3197 (N_3197,N_2251,N_2643);
or U3198 (N_3198,N_2452,N_2752);
nor U3199 (N_3199,N_2928,N_2875);
or U3200 (N_3200,N_2398,N_2313);
nand U3201 (N_3201,N_2342,N_2316);
nand U3202 (N_3202,N_2675,N_2843);
or U3203 (N_3203,N_2454,N_2294);
or U3204 (N_3204,N_2905,N_2475);
nor U3205 (N_3205,N_2417,N_2252);
and U3206 (N_3206,N_2340,N_2636);
nand U3207 (N_3207,N_2783,N_2816);
nor U3208 (N_3208,N_2708,N_2436);
and U3209 (N_3209,N_2687,N_2456);
or U3210 (N_3210,N_2379,N_2591);
nor U3211 (N_3211,N_2401,N_2495);
nand U3212 (N_3212,N_2485,N_2913);
or U3213 (N_3213,N_2626,N_2362);
nand U3214 (N_3214,N_2939,N_2753);
and U3215 (N_3215,N_2631,N_2549);
nor U3216 (N_3216,N_2544,N_2292);
and U3217 (N_3217,N_2628,N_2842);
nor U3218 (N_3218,N_2326,N_2374);
or U3219 (N_3219,N_2501,N_2490);
and U3220 (N_3220,N_2934,N_2366);
nor U3221 (N_3221,N_2878,N_2757);
nor U3222 (N_3222,N_2668,N_2853);
or U3223 (N_3223,N_2821,N_2533);
nor U3224 (N_3224,N_2781,N_2515);
nand U3225 (N_3225,N_2848,N_2741);
nand U3226 (N_3226,N_2740,N_2746);
nand U3227 (N_3227,N_2692,N_2590);
or U3228 (N_3228,N_2300,N_2826);
nor U3229 (N_3229,N_2258,N_2548);
nor U3230 (N_3230,N_2811,N_2262);
and U3231 (N_3231,N_2809,N_2271);
nor U3232 (N_3232,N_2424,N_2407);
or U3233 (N_3233,N_2953,N_2402);
or U3234 (N_3234,N_2573,N_2295);
nand U3235 (N_3235,N_2466,N_2993);
nor U3236 (N_3236,N_2518,N_2739);
and U3237 (N_3237,N_2375,N_2346);
nand U3238 (N_3238,N_2646,N_2660);
and U3239 (N_3239,N_2918,N_2261);
and U3240 (N_3240,N_2539,N_2729);
and U3241 (N_3241,N_2403,N_2334);
or U3242 (N_3242,N_2557,N_2435);
or U3243 (N_3243,N_2974,N_2443);
nand U3244 (N_3244,N_2806,N_2635);
and U3245 (N_3245,N_2613,N_2714);
nor U3246 (N_3246,N_2556,N_2348);
nand U3247 (N_3247,N_2662,N_2255);
and U3248 (N_3248,N_2513,N_2399);
or U3249 (N_3249,N_2620,N_2433);
nand U3250 (N_3250,N_2338,N_2872);
and U3251 (N_3251,N_2387,N_2947);
and U3252 (N_3252,N_2774,N_2270);
and U3253 (N_3253,N_2619,N_2896);
nor U3254 (N_3254,N_2653,N_2771);
and U3255 (N_3255,N_2975,N_2543);
nor U3256 (N_3256,N_2422,N_2290);
nand U3257 (N_3257,N_2582,N_2377);
or U3258 (N_3258,N_2711,N_2256);
nor U3259 (N_3259,N_2791,N_2560);
and U3260 (N_3260,N_2780,N_2921);
or U3261 (N_3261,N_2592,N_2852);
nand U3262 (N_3262,N_2690,N_2565);
or U3263 (N_3263,N_2327,N_2491);
nand U3264 (N_3264,N_2691,N_2859);
nand U3265 (N_3265,N_2350,N_2584);
nand U3266 (N_3266,N_2926,N_2483);
nor U3267 (N_3267,N_2611,N_2459);
nand U3268 (N_3268,N_2286,N_2959);
and U3269 (N_3269,N_2914,N_2522);
and U3270 (N_3270,N_2516,N_2416);
and U3271 (N_3271,N_2280,N_2985);
nor U3272 (N_3272,N_2259,N_2882);
nand U3273 (N_3273,N_2673,N_2347);
and U3274 (N_3274,N_2328,N_2920);
nand U3275 (N_3275,N_2969,N_2609);
or U3276 (N_3276,N_2672,N_2978);
nor U3277 (N_3277,N_2744,N_2587);
nor U3278 (N_3278,N_2893,N_2535);
or U3279 (N_3279,N_2960,N_2862);
nand U3280 (N_3280,N_2650,N_2310);
or U3281 (N_3281,N_2381,N_2888);
nand U3282 (N_3282,N_2908,N_2963);
nand U3283 (N_3283,N_2357,N_2736);
or U3284 (N_3284,N_2344,N_2521);
or U3285 (N_3285,N_2612,N_2337);
and U3286 (N_3286,N_2425,N_2274);
nand U3287 (N_3287,N_2589,N_2707);
and U3288 (N_3288,N_2499,N_2904);
nand U3289 (N_3289,N_2506,N_2886);
or U3290 (N_3290,N_2726,N_2911);
nand U3291 (N_3291,N_2877,N_2924);
nand U3292 (N_3292,N_2916,N_2644);
nor U3293 (N_3293,N_2706,N_2681);
nor U3294 (N_3294,N_2815,N_2468);
or U3295 (N_3295,N_2578,N_2779);
nor U3296 (N_3296,N_2583,N_2278);
nor U3297 (N_3297,N_2359,N_2388);
or U3298 (N_3298,N_2817,N_2296);
nand U3299 (N_3299,N_2283,N_2551);
nand U3300 (N_3300,N_2409,N_2800);
or U3301 (N_3301,N_2802,N_2686);
nor U3302 (N_3302,N_2568,N_2427);
or U3303 (N_3303,N_2919,N_2570);
and U3304 (N_3304,N_2343,N_2793);
and U3305 (N_3305,N_2530,N_2383);
nor U3306 (N_3306,N_2618,N_2936);
and U3307 (N_3307,N_2804,N_2488);
nor U3308 (N_3308,N_2880,N_2498);
nor U3309 (N_3309,N_2976,N_2319);
and U3310 (N_3310,N_2998,N_2487);
nand U3311 (N_3311,N_2810,N_2986);
nand U3312 (N_3312,N_2272,N_2420);
and U3313 (N_3313,N_2665,N_2517);
or U3314 (N_3314,N_2750,N_2754);
and U3315 (N_3315,N_2267,N_2664);
nand U3316 (N_3316,N_2307,N_2927);
or U3317 (N_3317,N_2434,N_2846);
and U3318 (N_3318,N_2712,N_2649);
or U3319 (N_3319,N_2891,N_2623);
nor U3320 (N_3320,N_2738,N_2532);
nand U3321 (N_3321,N_2633,N_2542);
nor U3322 (N_3322,N_2957,N_2666);
nand U3323 (N_3323,N_2449,N_2574);
or U3324 (N_3324,N_2710,N_2796);
or U3325 (N_3325,N_2699,N_2870);
and U3326 (N_3326,N_2894,N_2263);
nor U3327 (N_3327,N_2552,N_2423);
and U3328 (N_3328,N_2606,N_2429);
nand U3329 (N_3329,N_2685,N_2355);
nand U3330 (N_3330,N_2545,N_2415);
nor U3331 (N_3331,N_2260,N_2728);
or U3332 (N_3332,N_2266,N_2954);
or U3333 (N_3333,N_2776,N_2677);
nand U3334 (N_3334,N_2546,N_2419);
and U3335 (N_3335,N_2322,N_2762);
nand U3336 (N_3336,N_2866,N_2477);
or U3337 (N_3337,N_2448,N_2679);
and U3338 (N_3338,N_2538,N_2465);
nand U3339 (N_3339,N_2651,N_2536);
or U3340 (N_3340,N_2555,N_2418);
and U3341 (N_3341,N_2529,N_2977);
and U3342 (N_3342,N_2834,N_2803);
nand U3343 (N_3343,N_2265,N_2991);
nand U3344 (N_3344,N_2273,N_2923);
nand U3345 (N_3345,N_2331,N_2722);
and U3346 (N_3346,N_2558,N_2794);
nand U3347 (N_3347,N_2519,N_2742);
xor U3348 (N_3348,N_2311,N_2479);
and U3349 (N_3349,N_2901,N_2579);
nor U3350 (N_3350,N_2964,N_2768);
nor U3351 (N_3351,N_2526,N_2674);
and U3352 (N_3352,N_2540,N_2855);
and U3353 (N_3353,N_2798,N_2314);
or U3354 (N_3354,N_2887,N_2301);
or U3355 (N_3355,N_2782,N_2805);
nand U3356 (N_3356,N_2254,N_2778);
and U3357 (N_3357,N_2317,N_2647);
or U3358 (N_3358,N_2951,N_2309);
and U3359 (N_3359,N_2512,N_2588);
or U3360 (N_3360,N_2946,N_2358);
and U3361 (N_3361,N_2395,N_2683);
and U3362 (N_3362,N_2743,N_2447);
and U3363 (N_3363,N_2857,N_2411);
and U3364 (N_3364,N_2413,N_2962);
and U3365 (N_3365,N_2430,N_2850);
nand U3366 (N_3366,N_2735,N_2922);
and U3367 (N_3367,N_2765,N_2676);
nand U3368 (N_3368,N_2917,N_2825);
and U3369 (N_3369,N_2967,N_2365);
and U3370 (N_3370,N_2566,N_2500);
nand U3371 (N_3371,N_2881,N_2394);
or U3372 (N_3372,N_2979,N_2408);
or U3373 (N_3373,N_2593,N_2598);
and U3374 (N_3374,N_2335,N_2929);
or U3375 (N_3375,N_2483,N_2974);
or U3376 (N_3376,N_2717,N_2562);
nand U3377 (N_3377,N_2999,N_2434);
nand U3378 (N_3378,N_2293,N_2784);
and U3379 (N_3379,N_2635,N_2750);
nor U3380 (N_3380,N_2637,N_2528);
nor U3381 (N_3381,N_2446,N_2566);
or U3382 (N_3382,N_2435,N_2687);
and U3383 (N_3383,N_2581,N_2299);
nor U3384 (N_3384,N_2810,N_2969);
or U3385 (N_3385,N_2447,N_2376);
nand U3386 (N_3386,N_2933,N_2280);
nor U3387 (N_3387,N_2342,N_2604);
and U3388 (N_3388,N_2773,N_2673);
or U3389 (N_3389,N_2933,N_2393);
and U3390 (N_3390,N_2919,N_2933);
or U3391 (N_3391,N_2954,N_2865);
or U3392 (N_3392,N_2761,N_2919);
nor U3393 (N_3393,N_2429,N_2976);
nor U3394 (N_3394,N_2965,N_2332);
nand U3395 (N_3395,N_2627,N_2582);
and U3396 (N_3396,N_2654,N_2434);
or U3397 (N_3397,N_2843,N_2781);
or U3398 (N_3398,N_2693,N_2541);
or U3399 (N_3399,N_2538,N_2992);
nor U3400 (N_3400,N_2792,N_2280);
nand U3401 (N_3401,N_2325,N_2513);
and U3402 (N_3402,N_2426,N_2680);
and U3403 (N_3403,N_2648,N_2331);
nand U3404 (N_3404,N_2313,N_2571);
or U3405 (N_3405,N_2668,N_2824);
and U3406 (N_3406,N_2796,N_2298);
and U3407 (N_3407,N_2852,N_2943);
or U3408 (N_3408,N_2736,N_2588);
xnor U3409 (N_3409,N_2810,N_2851);
or U3410 (N_3410,N_2886,N_2457);
nand U3411 (N_3411,N_2343,N_2462);
or U3412 (N_3412,N_2967,N_2508);
nor U3413 (N_3413,N_2614,N_2700);
or U3414 (N_3414,N_2969,N_2558);
or U3415 (N_3415,N_2969,N_2340);
and U3416 (N_3416,N_2679,N_2437);
or U3417 (N_3417,N_2787,N_2445);
nand U3418 (N_3418,N_2309,N_2608);
or U3419 (N_3419,N_2832,N_2795);
nor U3420 (N_3420,N_2856,N_2701);
nor U3421 (N_3421,N_2762,N_2401);
or U3422 (N_3422,N_2272,N_2444);
or U3423 (N_3423,N_2281,N_2932);
nor U3424 (N_3424,N_2731,N_2327);
nand U3425 (N_3425,N_2364,N_2603);
nand U3426 (N_3426,N_2746,N_2419);
nand U3427 (N_3427,N_2979,N_2992);
nand U3428 (N_3428,N_2847,N_2494);
and U3429 (N_3429,N_2738,N_2744);
or U3430 (N_3430,N_2605,N_2402);
or U3431 (N_3431,N_2260,N_2484);
nand U3432 (N_3432,N_2556,N_2773);
nor U3433 (N_3433,N_2770,N_2358);
and U3434 (N_3434,N_2844,N_2708);
nor U3435 (N_3435,N_2593,N_2385);
nor U3436 (N_3436,N_2309,N_2613);
nand U3437 (N_3437,N_2405,N_2716);
xor U3438 (N_3438,N_2461,N_2636);
and U3439 (N_3439,N_2373,N_2602);
and U3440 (N_3440,N_2824,N_2352);
nor U3441 (N_3441,N_2670,N_2288);
nand U3442 (N_3442,N_2705,N_2696);
and U3443 (N_3443,N_2675,N_2468);
nand U3444 (N_3444,N_2485,N_2917);
or U3445 (N_3445,N_2683,N_2874);
or U3446 (N_3446,N_2549,N_2503);
or U3447 (N_3447,N_2459,N_2785);
nor U3448 (N_3448,N_2930,N_2941);
and U3449 (N_3449,N_2982,N_2313);
or U3450 (N_3450,N_2439,N_2493);
nand U3451 (N_3451,N_2372,N_2264);
and U3452 (N_3452,N_2331,N_2528);
nand U3453 (N_3453,N_2962,N_2403);
or U3454 (N_3454,N_2814,N_2727);
nor U3455 (N_3455,N_2930,N_2572);
nor U3456 (N_3456,N_2779,N_2297);
and U3457 (N_3457,N_2798,N_2298);
nor U3458 (N_3458,N_2360,N_2812);
nor U3459 (N_3459,N_2516,N_2689);
nor U3460 (N_3460,N_2768,N_2542);
nor U3461 (N_3461,N_2391,N_2736);
nor U3462 (N_3462,N_2452,N_2419);
and U3463 (N_3463,N_2724,N_2953);
or U3464 (N_3464,N_2966,N_2715);
nand U3465 (N_3465,N_2255,N_2683);
and U3466 (N_3466,N_2967,N_2505);
nor U3467 (N_3467,N_2408,N_2990);
nor U3468 (N_3468,N_2324,N_2524);
nor U3469 (N_3469,N_2397,N_2886);
or U3470 (N_3470,N_2965,N_2759);
and U3471 (N_3471,N_2310,N_2645);
nand U3472 (N_3472,N_2727,N_2834);
or U3473 (N_3473,N_2305,N_2823);
or U3474 (N_3474,N_2696,N_2404);
nand U3475 (N_3475,N_2589,N_2632);
and U3476 (N_3476,N_2762,N_2267);
nand U3477 (N_3477,N_2837,N_2830);
nor U3478 (N_3478,N_2396,N_2412);
nor U3479 (N_3479,N_2961,N_2377);
xnor U3480 (N_3480,N_2753,N_2778);
or U3481 (N_3481,N_2253,N_2297);
or U3482 (N_3482,N_2281,N_2945);
or U3483 (N_3483,N_2300,N_2988);
or U3484 (N_3484,N_2687,N_2909);
and U3485 (N_3485,N_2561,N_2568);
nor U3486 (N_3486,N_2984,N_2473);
and U3487 (N_3487,N_2274,N_2752);
or U3488 (N_3488,N_2983,N_2270);
and U3489 (N_3489,N_2792,N_2794);
and U3490 (N_3490,N_2550,N_2522);
and U3491 (N_3491,N_2728,N_2369);
nor U3492 (N_3492,N_2977,N_2353);
and U3493 (N_3493,N_2384,N_2823);
and U3494 (N_3494,N_2781,N_2291);
nor U3495 (N_3495,N_2354,N_2339);
nand U3496 (N_3496,N_2469,N_2760);
nor U3497 (N_3497,N_2824,N_2627);
and U3498 (N_3498,N_2358,N_2590);
nand U3499 (N_3499,N_2762,N_2282);
nor U3500 (N_3500,N_2908,N_2336);
nor U3501 (N_3501,N_2853,N_2841);
or U3502 (N_3502,N_2823,N_2654);
and U3503 (N_3503,N_2563,N_2847);
nand U3504 (N_3504,N_2251,N_2609);
nand U3505 (N_3505,N_2578,N_2780);
and U3506 (N_3506,N_2587,N_2376);
nand U3507 (N_3507,N_2928,N_2910);
nand U3508 (N_3508,N_2938,N_2783);
nand U3509 (N_3509,N_2517,N_2369);
nor U3510 (N_3510,N_2417,N_2265);
nor U3511 (N_3511,N_2632,N_2894);
nand U3512 (N_3512,N_2772,N_2727);
or U3513 (N_3513,N_2885,N_2631);
nor U3514 (N_3514,N_2335,N_2497);
nor U3515 (N_3515,N_2589,N_2794);
nand U3516 (N_3516,N_2271,N_2346);
and U3517 (N_3517,N_2696,N_2793);
nand U3518 (N_3518,N_2625,N_2266);
or U3519 (N_3519,N_2659,N_2519);
and U3520 (N_3520,N_2919,N_2789);
nor U3521 (N_3521,N_2403,N_2950);
xnor U3522 (N_3522,N_2452,N_2463);
and U3523 (N_3523,N_2800,N_2379);
and U3524 (N_3524,N_2298,N_2657);
nor U3525 (N_3525,N_2650,N_2783);
nand U3526 (N_3526,N_2731,N_2973);
nand U3527 (N_3527,N_2998,N_2273);
xnor U3528 (N_3528,N_2649,N_2539);
xnor U3529 (N_3529,N_2509,N_2851);
nand U3530 (N_3530,N_2905,N_2654);
nand U3531 (N_3531,N_2589,N_2848);
and U3532 (N_3532,N_2937,N_2739);
and U3533 (N_3533,N_2339,N_2379);
nor U3534 (N_3534,N_2595,N_2934);
xor U3535 (N_3535,N_2517,N_2356);
or U3536 (N_3536,N_2643,N_2696);
nand U3537 (N_3537,N_2995,N_2732);
and U3538 (N_3538,N_2498,N_2442);
or U3539 (N_3539,N_2619,N_2312);
nor U3540 (N_3540,N_2828,N_2750);
nand U3541 (N_3541,N_2390,N_2290);
nand U3542 (N_3542,N_2391,N_2467);
and U3543 (N_3543,N_2580,N_2926);
and U3544 (N_3544,N_2572,N_2884);
nand U3545 (N_3545,N_2407,N_2372);
nand U3546 (N_3546,N_2279,N_2506);
nor U3547 (N_3547,N_2714,N_2495);
or U3548 (N_3548,N_2284,N_2839);
nor U3549 (N_3549,N_2787,N_2739);
nand U3550 (N_3550,N_2835,N_2709);
or U3551 (N_3551,N_2324,N_2961);
nor U3552 (N_3552,N_2377,N_2358);
nand U3553 (N_3553,N_2325,N_2699);
nand U3554 (N_3554,N_2975,N_2748);
nand U3555 (N_3555,N_2828,N_2798);
nand U3556 (N_3556,N_2601,N_2340);
nor U3557 (N_3557,N_2621,N_2411);
xnor U3558 (N_3558,N_2898,N_2366);
nor U3559 (N_3559,N_2557,N_2540);
or U3560 (N_3560,N_2598,N_2686);
nand U3561 (N_3561,N_2253,N_2845);
and U3562 (N_3562,N_2782,N_2412);
or U3563 (N_3563,N_2947,N_2977);
nor U3564 (N_3564,N_2803,N_2436);
or U3565 (N_3565,N_2996,N_2710);
and U3566 (N_3566,N_2731,N_2682);
nor U3567 (N_3567,N_2849,N_2673);
nand U3568 (N_3568,N_2260,N_2412);
or U3569 (N_3569,N_2633,N_2532);
and U3570 (N_3570,N_2382,N_2658);
nand U3571 (N_3571,N_2550,N_2476);
or U3572 (N_3572,N_2397,N_2914);
or U3573 (N_3573,N_2800,N_2953);
and U3574 (N_3574,N_2525,N_2853);
or U3575 (N_3575,N_2481,N_2802);
nor U3576 (N_3576,N_2636,N_2496);
or U3577 (N_3577,N_2250,N_2346);
nor U3578 (N_3578,N_2810,N_2781);
nand U3579 (N_3579,N_2538,N_2578);
nor U3580 (N_3580,N_2267,N_2858);
nor U3581 (N_3581,N_2856,N_2412);
or U3582 (N_3582,N_2887,N_2799);
nand U3583 (N_3583,N_2913,N_2690);
or U3584 (N_3584,N_2607,N_2936);
and U3585 (N_3585,N_2992,N_2915);
and U3586 (N_3586,N_2267,N_2695);
or U3587 (N_3587,N_2936,N_2854);
and U3588 (N_3588,N_2769,N_2277);
and U3589 (N_3589,N_2651,N_2364);
or U3590 (N_3590,N_2369,N_2493);
nand U3591 (N_3591,N_2631,N_2374);
nor U3592 (N_3592,N_2328,N_2326);
and U3593 (N_3593,N_2334,N_2641);
and U3594 (N_3594,N_2524,N_2269);
nand U3595 (N_3595,N_2776,N_2882);
or U3596 (N_3596,N_2545,N_2830);
and U3597 (N_3597,N_2424,N_2439);
nand U3598 (N_3598,N_2783,N_2894);
nor U3599 (N_3599,N_2484,N_2587);
nor U3600 (N_3600,N_2883,N_2706);
or U3601 (N_3601,N_2303,N_2611);
nor U3602 (N_3602,N_2674,N_2310);
or U3603 (N_3603,N_2409,N_2961);
and U3604 (N_3604,N_2918,N_2562);
nor U3605 (N_3605,N_2905,N_2852);
nor U3606 (N_3606,N_2984,N_2374);
and U3607 (N_3607,N_2308,N_2635);
xnor U3608 (N_3608,N_2425,N_2470);
and U3609 (N_3609,N_2531,N_2436);
and U3610 (N_3610,N_2949,N_2510);
or U3611 (N_3611,N_2343,N_2803);
nor U3612 (N_3612,N_2370,N_2929);
nand U3613 (N_3613,N_2354,N_2531);
and U3614 (N_3614,N_2612,N_2289);
or U3615 (N_3615,N_2364,N_2957);
nand U3616 (N_3616,N_2986,N_2947);
or U3617 (N_3617,N_2757,N_2398);
or U3618 (N_3618,N_2439,N_2762);
nand U3619 (N_3619,N_2935,N_2948);
nand U3620 (N_3620,N_2300,N_2570);
nor U3621 (N_3621,N_2618,N_2881);
or U3622 (N_3622,N_2713,N_2469);
or U3623 (N_3623,N_2823,N_2840);
and U3624 (N_3624,N_2326,N_2914);
or U3625 (N_3625,N_2779,N_2363);
nand U3626 (N_3626,N_2823,N_2420);
or U3627 (N_3627,N_2736,N_2757);
or U3628 (N_3628,N_2780,N_2776);
and U3629 (N_3629,N_2294,N_2718);
nand U3630 (N_3630,N_2688,N_2660);
and U3631 (N_3631,N_2272,N_2376);
nor U3632 (N_3632,N_2266,N_2392);
nand U3633 (N_3633,N_2389,N_2837);
nor U3634 (N_3634,N_2417,N_2290);
nand U3635 (N_3635,N_2336,N_2482);
and U3636 (N_3636,N_2317,N_2394);
or U3637 (N_3637,N_2260,N_2731);
or U3638 (N_3638,N_2346,N_2751);
nor U3639 (N_3639,N_2553,N_2759);
and U3640 (N_3640,N_2700,N_2437);
xor U3641 (N_3641,N_2404,N_2927);
nand U3642 (N_3642,N_2321,N_2714);
nor U3643 (N_3643,N_2413,N_2557);
or U3644 (N_3644,N_2896,N_2438);
nand U3645 (N_3645,N_2290,N_2549);
or U3646 (N_3646,N_2384,N_2945);
nor U3647 (N_3647,N_2592,N_2755);
nand U3648 (N_3648,N_2380,N_2996);
or U3649 (N_3649,N_2942,N_2645);
nor U3650 (N_3650,N_2624,N_2846);
nand U3651 (N_3651,N_2771,N_2744);
and U3652 (N_3652,N_2931,N_2678);
nand U3653 (N_3653,N_2714,N_2827);
nor U3654 (N_3654,N_2617,N_2586);
nand U3655 (N_3655,N_2695,N_2698);
nand U3656 (N_3656,N_2292,N_2751);
or U3657 (N_3657,N_2540,N_2613);
nand U3658 (N_3658,N_2744,N_2791);
nor U3659 (N_3659,N_2555,N_2585);
nand U3660 (N_3660,N_2503,N_2860);
or U3661 (N_3661,N_2872,N_2786);
and U3662 (N_3662,N_2658,N_2618);
and U3663 (N_3663,N_2521,N_2653);
nor U3664 (N_3664,N_2748,N_2762);
nand U3665 (N_3665,N_2337,N_2301);
and U3666 (N_3666,N_2691,N_2833);
and U3667 (N_3667,N_2508,N_2978);
and U3668 (N_3668,N_2770,N_2461);
or U3669 (N_3669,N_2373,N_2583);
xnor U3670 (N_3670,N_2865,N_2977);
nor U3671 (N_3671,N_2684,N_2361);
or U3672 (N_3672,N_2959,N_2598);
nand U3673 (N_3673,N_2835,N_2634);
and U3674 (N_3674,N_2769,N_2318);
nor U3675 (N_3675,N_2862,N_2715);
and U3676 (N_3676,N_2935,N_2877);
or U3677 (N_3677,N_2551,N_2378);
nand U3678 (N_3678,N_2330,N_2417);
nor U3679 (N_3679,N_2876,N_2768);
and U3680 (N_3680,N_2748,N_2441);
nor U3681 (N_3681,N_2718,N_2280);
nor U3682 (N_3682,N_2592,N_2534);
nand U3683 (N_3683,N_2995,N_2940);
nor U3684 (N_3684,N_2569,N_2714);
nor U3685 (N_3685,N_2546,N_2763);
nor U3686 (N_3686,N_2404,N_2484);
nor U3687 (N_3687,N_2412,N_2615);
and U3688 (N_3688,N_2762,N_2595);
nand U3689 (N_3689,N_2884,N_2983);
or U3690 (N_3690,N_2717,N_2448);
and U3691 (N_3691,N_2792,N_2956);
or U3692 (N_3692,N_2250,N_2749);
and U3693 (N_3693,N_2735,N_2517);
nand U3694 (N_3694,N_2351,N_2526);
or U3695 (N_3695,N_2862,N_2500);
nand U3696 (N_3696,N_2582,N_2937);
or U3697 (N_3697,N_2574,N_2906);
and U3698 (N_3698,N_2399,N_2875);
nor U3699 (N_3699,N_2460,N_2757);
and U3700 (N_3700,N_2545,N_2735);
nor U3701 (N_3701,N_2789,N_2631);
nor U3702 (N_3702,N_2333,N_2827);
nor U3703 (N_3703,N_2632,N_2853);
and U3704 (N_3704,N_2683,N_2776);
or U3705 (N_3705,N_2787,N_2549);
and U3706 (N_3706,N_2351,N_2938);
and U3707 (N_3707,N_2727,N_2465);
or U3708 (N_3708,N_2705,N_2708);
or U3709 (N_3709,N_2834,N_2820);
nand U3710 (N_3710,N_2383,N_2535);
and U3711 (N_3711,N_2466,N_2862);
nor U3712 (N_3712,N_2709,N_2524);
nand U3713 (N_3713,N_2318,N_2809);
xor U3714 (N_3714,N_2902,N_2946);
or U3715 (N_3715,N_2632,N_2391);
and U3716 (N_3716,N_2968,N_2425);
nand U3717 (N_3717,N_2956,N_2883);
or U3718 (N_3718,N_2502,N_2954);
nor U3719 (N_3719,N_2265,N_2554);
or U3720 (N_3720,N_2315,N_2250);
or U3721 (N_3721,N_2279,N_2749);
and U3722 (N_3722,N_2860,N_2456);
and U3723 (N_3723,N_2554,N_2557);
nand U3724 (N_3724,N_2465,N_2765);
nor U3725 (N_3725,N_2906,N_2551);
or U3726 (N_3726,N_2528,N_2458);
and U3727 (N_3727,N_2512,N_2877);
and U3728 (N_3728,N_2712,N_2828);
and U3729 (N_3729,N_2746,N_2381);
nand U3730 (N_3730,N_2566,N_2518);
nand U3731 (N_3731,N_2406,N_2308);
nand U3732 (N_3732,N_2639,N_2608);
nor U3733 (N_3733,N_2785,N_2847);
nor U3734 (N_3734,N_2464,N_2497);
nor U3735 (N_3735,N_2391,N_2766);
nor U3736 (N_3736,N_2851,N_2338);
and U3737 (N_3737,N_2752,N_2971);
and U3738 (N_3738,N_2686,N_2258);
and U3739 (N_3739,N_2631,N_2392);
and U3740 (N_3740,N_2501,N_2886);
nor U3741 (N_3741,N_2563,N_2556);
nor U3742 (N_3742,N_2334,N_2716);
or U3743 (N_3743,N_2397,N_2328);
and U3744 (N_3744,N_2545,N_2316);
or U3745 (N_3745,N_2919,N_2868);
or U3746 (N_3746,N_2437,N_2826);
nor U3747 (N_3747,N_2413,N_2523);
nor U3748 (N_3748,N_2587,N_2997);
nand U3749 (N_3749,N_2329,N_2881);
nor U3750 (N_3750,N_3392,N_3296);
or U3751 (N_3751,N_3334,N_3206);
or U3752 (N_3752,N_3199,N_3132);
nor U3753 (N_3753,N_3650,N_3431);
nor U3754 (N_3754,N_3578,N_3530);
and U3755 (N_3755,N_3406,N_3268);
and U3756 (N_3756,N_3173,N_3124);
nand U3757 (N_3757,N_3463,N_3198);
and U3758 (N_3758,N_3653,N_3277);
or U3759 (N_3759,N_3086,N_3708);
nor U3760 (N_3760,N_3117,N_3218);
and U3761 (N_3761,N_3420,N_3271);
nor U3762 (N_3762,N_3372,N_3022);
or U3763 (N_3763,N_3287,N_3395);
nand U3764 (N_3764,N_3566,N_3721);
xor U3765 (N_3765,N_3599,N_3148);
nand U3766 (N_3766,N_3363,N_3348);
or U3767 (N_3767,N_3010,N_3492);
nor U3768 (N_3768,N_3454,N_3353);
or U3769 (N_3769,N_3172,N_3633);
and U3770 (N_3770,N_3498,N_3582);
and U3771 (N_3771,N_3478,N_3640);
nor U3772 (N_3772,N_3565,N_3562);
or U3773 (N_3773,N_3641,N_3228);
nor U3774 (N_3774,N_3432,N_3627);
or U3775 (N_3775,N_3476,N_3371);
nand U3776 (N_3776,N_3488,N_3546);
and U3777 (N_3777,N_3682,N_3396);
and U3778 (N_3778,N_3734,N_3731);
nand U3779 (N_3779,N_3591,N_3009);
or U3780 (N_3780,N_3075,N_3030);
nand U3781 (N_3781,N_3312,N_3537);
or U3782 (N_3782,N_3303,N_3114);
and U3783 (N_3783,N_3725,N_3288);
nor U3784 (N_3784,N_3576,N_3036);
and U3785 (N_3785,N_3624,N_3350);
nor U3786 (N_3786,N_3068,N_3096);
nand U3787 (N_3787,N_3084,N_3062);
and U3788 (N_3788,N_3176,N_3186);
or U3789 (N_3789,N_3158,N_3361);
nand U3790 (N_3790,N_3364,N_3581);
and U3791 (N_3791,N_3729,N_3482);
nor U3792 (N_3792,N_3259,N_3143);
and U3793 (N_3793,N_3024,N_3294);
nor U3794 (N_3794,N_3090,N_3458);
nand U3795 (N_3795,N_3051,N_3033);
or U3796 (N_3796,N_3233,N_3203);
or U3797 (N_3797,N_3025,N_3265);
nor U3798 (N_3798,N_3178,N_3179);
and U3799 (N_3799,N_3521,N_3315);
and U3800 (N_3800,N_3246,N_3106);
or U3801 (N_3801,N_3507,N_3144);
or U3802 (N_3802,N_3526,N_3425);
nand U3803 (N_3803,N_3192,N_3103);
or U3804 (N_3804,N_3409,N_3029);
or U3805 (N_3805,N_3436,N_3673);
nor U3806 (N_3806,N_3380,N_3485);
nor U3807 (N_3807,N_3672,N_3517);
nor U3808 (N_3808,N_3428,N_3523);
nor U3809 (N_3809,N_3214,N_3719);
nor U3810 (N_3810,N_3330,N_3568);
or U3811 (N_3811,N_3127,N_3706);
nand U3812 (N_3812,N_3157,N_3621);
nor U3813 (N_3813,N_3477,N_3328);
nor U3814 (N_3814,N_3669,N_3710);
and U3815 (N_3815,N_3610,N_3461);
nor U3816 (N_3816,N_3447,N_3366);
nor U3817 (N_3817,N_3159,N_3067);
and U3818 (N_3818,N_3389,N_3598);
nand U3819 (N_3819,N_3049,N_3320);
nor U3820 (N_3820,N_3619,N_3560);
nand U3821 (N_3821,N_3405,N_3234);
nand U3822 (N_3822,N_3702,N_3063);
and U3823 (N_3823,N_3381,N_3607);
and U3824 (N_3824,N_3401,N_3243);
nor U3825 (N_3825,N_3065,N_3635);
xor U3826 (N_3826,N_3441,N_3700);
nor U3827 (N_3827,N_3433,N_3440);
or U3828 (N_3828,N_3491,N_3301);
or U3829 (N_3829,N_3168,N_3101);
and U3830 (N_3830,N_3429,N_3166);
nor U3831 (N_3831,N_3612,N_3533);
nand U3832 (N_3832,N_3443,N_3462);
and U3833 (N_3833,N_3365,N_3539);
and U3834 (N_3834,N_3455,N_3021);
and U3835 (N_3835,N_3535,N_3514);
or U3836 (N_3836,N_3654,N_3239);
nor U3837 (N_3837,N_3648,N_3577);
nor U3838 (N_3838,N_3270,N_3260);
nand U3839 (N_3839,N_3129,N_3616);
xnor U3840 (N_3840,N_3674,N_3709);
and U3841 (N_3841,N_3235,N_3087);
nand U3842 (N_3842,N_3304,N_3745);
xor U3843 (N_3843,N_3080,N_3574);
nor U3844 (N_3844,N_3076,N_3722);
nor U3845 (N_3845,N_3370,N_3630);
and U3846 (N_3846,N_3314,N_3368);
nor U3847 (N_3847,N_3543,N_3164);
or U3848 (N_3848,N_3445,N_3601);
nor U3849 (N_3849,N_3605,N_3085);
or U3850 (N_3850,N_3554,N_3423);
and U3851 (N_3851,N_3329,N_3412);
nor U3852 (N_3852,N_3019,N_3319);
nor U3853 (N_3853,N_3050,N_3707);
or U3854 (N_3854,N_3230,N_3390);
and U3855 (N_3855,N_3376,N_3267);
and U3856 (N_3856,N_3394,N_3603);
nand U3857 (N_3857,N_3494,N_3358);
nand U3858 (N_3858,N_3446,N_3538);
nor U3859 (N_3859,N_3404,N_3282);
nand U3860 (N_3860,N_3520,N_3109);
nand U3861 (N_3861,N_3338,N_3094);
nor U3862 (N_3862,N_3182,N_3400);
xnor U3863 (N_3863,N_3074,N_3584);
nand U3864 (N_3864,N_3378,N_3006);
and U3865 (N_3865,N_3480,N_3295);
nand U3866 (N_3866,N_3437,N_3592);
nand U3867 (N_3867,N_3023,N_3043);
nand U3868 (N_3868,N_3205,N_3618);
and U3869 (N_3869,N_3735,N_3647);
or U3870 (N_3870,N_3570,N_3118);
or U3871 (N_3871,N_3138,N_3548);
nand U3872 (N_3872,N_3519,N_3013);
and U3873 (N_3873,N_3232,N_3174);
and U3874 (N_3874,N_3667,N_3306);
and U3875 (N_3875,N_3196,N_3684);
and U3876 (N_3876,N_3016,N_3649);
nor U3877 (N_3877,N_3511,N_3726);
or U3878 (N_3878,N_3435,N_3339);
and U3879 (N_3879,N_3430,N_3255);
nor U3880 (N_3880,N_3217,N_3718);
nor U3881 (N_3881,N_3559,N_3397);
and U3882 (N_3882,N_3279,N_3170);
or U3883 (N_3883,N_3620,N_3595);
nor U3884 (N_3884,N_3007,N_3048);
nor U3885 (N_3885,N_3438,N_3623);
or U3886 (N_3886,N_3497,N_3202);
nor U3887 (N_3887,N_3383,N_3208);
nand U3888 (N_3888,N_3356,N_3183);
xor U3889 (N_3889,N_3632,N_3008);
nand U3890 (N_3890,N_3678,N_3626);
or U3891 (N_3891,N_3308,N_3716);
or U3892 (N_3892,N_3072,N_3163);
nor U3893 (N_3893,N_3453,N_3345);
nor U3894 (N_3894,N_3439,N_3490);
or U3895 (N_3895,N_3026,N_3189);
nand U3896 (N_3896,N_3427,N_3225);
nor U3897 (N_3897,N_3272,N_3638);
and U3898 (N_3898,N_3387,N_3139);
nor U3899 (N_3899,N_3506,N_3666);
nand U3900 (N_3900,N_3073,N_3108);
nor U3901 (N_3901,N_3130,N_3622);
nand U3902 (N_3902,N_3015,N_3256);
nor U3903 (N_3903,N_3317,N_3579);
nand U3904 (N_3904,N_3466,N_3407);
nand U3905 (N_3905,N_3529,N_3692);
nand U3906 (N_3906,N_3054,N_3421);
or U3907 (N_3907,N_3664,N_3374);
nor U3908 (N_3908,N_3585,N_3422);
nand U3909 (N_3909,N_3167,N_3083);
or U3910 (N_3910,N_3588,N_3059);
nand U3911 (N_3911,N_3636,N_3698);
nor U3912 (N_3912,N_3711,N_3242);
and U3913 (N_3913,N_3112,N_3379);
nand U3914 (N_3914,N_3160,N_3424);
nor U3915 (N_3915,N_3691,N_3133);
and U3916 (N_3916,N_3123,N_3657);
and U3917 (N_3917,N_3609,N_3697);
and U3918 (N_3918,N_3012,N_3060);
or U3919 (N_3919,N_3194,N_3252);
and U3920 (N_3920,N_3216,N_3683);
nand U3921 (N_3921,N_3212,N_3528);
nor U3922 (N_3922,N_3237,N_3495);
nor U3923 (N_3923,N_3651,N_3525);
or U3924 (N_3924,N_3058,N_3644);
and U3925 (N_3925,N_3316,N_3590);
or U3926 (N_3926,N_3318,N_3020);
nand U3927 (N_3927,N_3249,N_3555);
nor U3928 (N_3928,N_3699,N_3238);
and U3929 (N_3929,N_3587,N_3081);
and U3930 (N_3930,N_3696,N_3193);
and U3931 (N_3931,N_3248,N_3542);
nand U3932 (N_3932,N_3518,N_3322);
nor U3933 (N_3933,N_3355,N_3274);
nand U3934 (N_3934,N_3126,N_3418);
nor U3935 (N_3935,N_3034,N_3403);
or U3936 (N_3936,N_3694,N_3503);
nand U3937 (N_3937,N_3111,N_3464);
and U3938 (N_3938,N_3136,N_3035);
and U3939 (N_3939,N_3145,N_3197);
or U3940 (N_3940,N_3335,N_3135);
nand U3941 (N_3941,N_3093,N_3089);
or U3942 (N_3942,N_3276,N_3465);
or U3943 (N_3943,N_3662,N_3028);
nand U3944 (N_3944,N_3434,N_3448);
or U3945 (N_3945,N_3741,N_3646);
and U3946 (N_3946,N_3597,N_3540);
and U3947 (N_3947,N_3367,N_3291);
nand U3948 (N_3948,N_3341,N_3410);
nor U3949 (N_3949,N_3298,N_3483);
nand U3950 (N_3950,N_3047,N_3629);
or U3951 (N_3951,N_3137,N_3689);
or U3952 (N_3952,N_3037,N_3385);
and U3953 (N_3953,N_3284,N_3125);
nor U3954 (N_3954,N_3705,N_3146);
nor U3955 (N_3955,N_3739,N_3349);
or U3956 (N_3956,N_3169,N_3408);
nand U3957 (N_3957,N_3285,N_3375);
or U3958 (N_3958,N_3305,N_3512);
or U3959 (N_3959,N_3082,N_3141);
nor U3960 (N_3960,N_3444,N_3567);
nand U3961 (N_3961,N_3343,N_3088);
and U3962 (N_3962,N_3027,N_3631);
and U3963 (N_3963,N_3289,N_3606);
or U3964 (N_3964,N_3634,N_3474);
or U3965 (N_3965,N_3360,N_3263);
nor U3966 (N_3966,N_3241,N_3748);
and U3967 (N_3967,N_3323,N_3541);
and U3968 (N_3968,N_3362,N_3264);
nor U3969 (N_3969,N_3665,N_3275);
and U3970 (N_3970,N_3617,N_3704);
and U3971 (N_3971,N_3253,N_3128);
nand U3972 (N_3972,N_3740,N_3254);
or U3973 (N_3973,N_3229,N_3737);
nand U3974 (N_3974,N_3652,N_3701);
nand U3975 (N_3975,N_3044,N_3642);
and U3976 (N_3976,N_3031,N_3457);
nor U3977 (N_3977,N_3245,N_3278);
nand U3978 (N_3978,N_3715,N_3614);
and U3979 (N_3979,N_3207,N_3219);
nand U3980 (N_3980,N_3100,N_3593);
nor U3981 (N_3981,N_3723,N_3104);
xor U3982 (N_3982,N_3057,N_3484);
and U3983 (N_3983,N_3663,N_3052);
or U3984 (N_3984,N_3185,N_3602);
or U3985 (N_3985,N_3105,N_3177);
nand U3986 (N_3986,N_3116,N_3502);
xnor U3987 (N_3987,N_3522,N_3534);
nand U3988 (N_3988,N_3501,N_3014);
and U3989 (N_3989,N_3107,N_3442);
nand U3990 (N_3990,N_3677,N_3213);
nand U3991 (N_3991,N_3600,N_3188);
nand U3992 (N_3992,N_3744,N_3551);
nand U3993 (N_3993,N_3262,N_3352);
nor U3994 (N_3994,N_3120,N_3680);
or U3995 (N_3995,N_3738,N_3300);
xor U3996 (N_3996,N_3038,N_3505);
nor U3997 (N_3997,N_3190,N_3215);
or U3998 (N_3998,N_3414,N_3149);
and U3999 (N_3999,N_3563,N_3005);
or U4000 (N_4000,N_3211,N_3569);
nor U4001 (N_4001,N_3281,N_3515);
nor U4002 (N_4002,N_3098,N_3686);
or U4003 (N_4003,N_3717,N_3359);
or U4004 (N_4004,N_3299,N_3573);
nor U4005 (N_4005,N_3327,N_3449);
or U4006 (N_4006,N_3628,N_3504);
nor U4007 (N_4007,N_3655,N_3175);
nand U4008 (N_4008,N_3223,N_3187);
and U4009 (N_4009,N_3313,N_3733);
nor U4010 (N_4010,N_3589,N_3344);
nor U4011 (N_4011,N_3184,N_3416);
nor U4012 (N_4012,N_3377,N_3459);
and U4013 (N_4013,N_3415,N_3333);
nand U4014 (N_4014,N_3531,N_3625);
nand U4015 (N_4015,N_3549,N_3419);
and U4016 (N_4016,N_3712,N_3045);
or U4017 (N_4017,N_3002,N_3236);
nand U4018 (N_4018,N_3131,N_3496);
or U4019 (N_4019,N_3309,N_3095);
nand U4020 (N_4020,N_3000,N_3608);
xnor U4021 (N_4021,N_3347,N_3283);
nor U4022 (N_4022,N_3643,N_3055);
nand U4023 (N_4023,N_3572,N_3042);
nand U4024 (N_4024,N_3473,N_3292);
nor U4025 (N_4025,N_3056,N_3749);
and U4026 (N_4026,N_3645,N_3247);
and U4027 (N_4027,N_3398,N_3261);
and U4028 (N_4028,N_3687,N_3671);
nor U4029 (N_4029,N_3544,N_3451);
or U4030 (N_4030,N_3204,N_3547);
and U4031 (N_4031,N_3475,N_3553);
nand U4032 (N_4032,N_3388,N_3332);
or U4033 (N_4033,N_3516,N_3311);
nand U4034 (N_4034,N_3097,N_3201);
and U4035 (N_4035,N_3596,N_3018);
nor U4036 (N_4036,N_3724,N_3180);
nand U4037 (N_4037,N_3659,N_3558);
nor U4038 (N_4038,N_3594,N_3615);
or U4039 (N_4039,N_3269,N_3121);
nand U4040 (N_4040,N_3658,N_3685);
nand U4041 (N_4041,N_3670,N_3011);
and U4042 (N_4042,N_3140,N_3102);
nor U4043 (N_4043,N_3639,N_3061);
nand U4044 (N_4044,N_3077,N_3720);
and U4045 (N_4045,N_3452,N_3152);
nand U4046 (N_4046,N_3142,N_3460);
and U4047 (N_4047,N_3550,N_3342);
and U4048 (N_4048,N_3417,N_3017);
nor U4049 (N_4049,N_3280,N_3310);
and U4050 (N_4050,N_3536,N_3070);
or U4051 (N_4051,N_3171,N_3064);
and U4052 (N_4052,N_3250,N_3134);
nand U4053 (N_4053,N_3742,N_3181);
and U4054 (N_4054,N_3003,N_3393);
or U4055 (N_4055,N_3220,N_3331);
nor U4056 (N_4056,N_3115,N_3747);
or U4057 (N_4057,N_3325,N_3481);
or U4058 (N_4058,N_3471,N_3732);
nor U4059 (N_4059,N_3557,N_3221);
or U4060 (N_4060,N_3561,N_3676);
nand U4061 (N_4061,N_3091,N_3346);
and U4062 (N_4062,N_3730,N_3426);
nor U4063 (N_4063,N_3266,N_3326);
or U4064 (N_4064,N_3545,N_3079);
and U4065 (N_4065,N_3119,N_3373);
or U4066 (N_4066,N_3611,N_3524);
nand U4067 (N_4067,N_3222,N_3532);
nor U4068 (N_4068,N_3575,N_3604);
nor U4069 (N_4069,N_3487,N_3357);
nor U4070 (N_4070,N_3244,N_3258);
nand U4071 (N_4071,N_3110,N_3069);
nand U4072 (N_4072,N_3470,N_3195);
xnor U4073 (N_4073,N_3210,N_3154);
nand U4074 (N_4074,N_3382,N_3399);
nor U4075 (N_4075,N_3302,N_3209);
nor U4076 (N_4076,N_3099,N_3571);
and U4077 (N_4077,N_3469,N_3656);
or U4078 (N_4078,N_3078,N_3564);
or U4079 (N_4079,N_3307,N_3369);
xor U4080 (N_4080,N_3402,N_3290);
nor U4081 (N_4081,N_3714,N_3113);
nand U4082 (N_4082,N_3411,N_3675);
nand U4083 (N_4083,N_3486,N_3191);
nor U4084 (N_4084,N_3257,N_3668);
or U4085 (N_4085,N_3150,N_3324);
xnor U4086 (N_4086,N_3001,N_3552);
nand U4087 (N_4087,N_3231,N_3153);
nand U4088 (N_4088,N_3489,N_3472);
nand U4089 (N_4089,N_3041,N_3240);
nor U4090 (N_4090,N_3391,N_3556);
nor U4091 (N_4091,N_3336,N_3092);
or U4092 (N_4092,N_3746,N_3467);
nand U4093 (N_4093,N_3613,N_3527);
and U4094 (N_4094,N_3450,N_3122);
nor U4095 (N_4095,N_3040,N_3583);
nand U4096 (N_4096,N_3354,N_3273);
nand U4097 (N_4097,N_3703,N_3661);
or U4098 (N_4098,N_3200,N_3499);
and U4099 (N_4099,N_3147,N_3337);
nand U4100 (N_4100,N_3046,N_3162);
nor U4101 (N_4101,N_3510,N_3713);
nor U4102 (N_4102,N_3321,N_3580);
or U4103 (N_4103,N_3293,N_3681);
or U4104 (N_4104,N_3468,N_3004);
nand U4105 (N_4105,N_3032,N_3508);
nand U4106 (N_4106,N_3340,N_3513);
or U4107 (N_4107,N_3456,N_3727);
and U4108 (N_4108,N_3743,N_3637);
nor U4109 (N_4109,N_3493,N_3156);
nand U4110 (N_4110,N_3693,N_3039);
or U4111 (N_4111,N_3660,N_3286);
or U4112 (N_4112,N_3351,N_3690);
nand U4113 (N_4113,N_3155,N_3695);
nor U4114 (N_4114,N_3384,N_3224);
nand U4115 (N_4115,N_3251,N_3297);
or U4116 (N_4116,N_3736,N_3728);
or U4117 (N_4117,N_3509,N_3386);
nand U4118 (N_4118,N_3688,N_3500);
nor U4119 (N_4119,N_3165,N_3586);
nand U4120 (N_4120,N_3413,N_3053);
or U4121 (N_4121,N_3226,N_3679);
nor U4122 (N_4122,N_3151,N_3161);
nor U4123 (N_4123,N_3071,N_3066);
and U4124 (N_4124,N_3479,N_3227);
nand U4125 (N_4125,N_3138,N_3702);
nor U4126 (N_4126,N_3346,N_3030);
nand U4127 (N_4127,N_3248,N_3709);
nand U4128 (N_4128,N_3162,N_3366);
or U4129 (N_4129,N_3692,N_3175);
or U4130 (N_4130,N_3543,N_3711);
nand U4131 (N_4131,N_3526,N_3650);
and U4132 (N_4132,N_3101,N_3274);
and U4133 (N_4133,N_3485,N_3449);
or U4134 (N_4134,N_3397,N_3275);
and U4135 (N_4135,N_3637,N_3327);
nand U4136 (N_4136,N_3603,N_3699);
nand U4137 (N_4137,N_3399,N_3625);
and U4138 (N_4138,N_3416,N_3421);
or U4139 (N_4139,N_3596,N_3605);
and U4140 (N_4140,N_3100,N_3562);
and U4141 (N_4141,N_3413,N_3212);
nand U4142 (N_4142,N_3022,N_3027);
or U4143 (N_4143,N_3147,N_3289);
and U4144 (N_4144,N_3579,N_3139);
nor U4145 (N_4145,N_3421,N_3493);
nand U4146 (N_4146,N_3343,N_3316);
nand U4147 (N_4147,N_3149,N_3693);
and U4148 (N_4148,N_3609,N_3458);
nand U4149 (N_4149,N_3086,N_3384);
and U4150 (N_4150,N_3543,N_3222);
nor U4151 (N_4151,N_3530,N_3162);
or U4152 (N_4152,N_3360,N_3165);
nand U4153 (N_4153,N_3449,N_3732);
or U4154 (N_4154,N_3438,N_3677);
nor U4155 (N_4155,N_3097,N_3716);
nor U4156 (N_4156,N_3697,N_3549);
nor U4157 (N_4157,N_3398,N_3360);
nor U4158 (N_4158,N_3243,N_3387);
or U4159 (N_4159,N_3572,N_3200);
nor U4160 (N_4160,N_3232,N_3359);
nand U4161 (N_4161,N_3430,N_3707);
and U4162 (N_4162,N_3598,N_3514);
nand U4163 (N_4163,N_3412,N_3286);
or U4164 (N_4164,N_3197,N_3157);
nor U4165 (N_4165,N_3433,N_3490);
nand U4166 (N_4166,N_3482,N_3173);
and U4167 (N_4167,N_3167,N_3163);
or U4168 (N_4168,N_3447,N_3665);
and U4169 (N_4169,N_3021,N_3266);
and U4170 (N_4170,N_3490,N_3187);
nor U4171 (N_4171,N_3026,N_3601);
and U4172 (N_4172,N_3563,N_3192);
or U4173 (N_4173,N_3614,N_3102);
nand U4174 (N_4174,N_3428,N_3327);
xnor U4175 (N_4175,N_3336,N_3103);
and U4176 (N_4176,N_3638,N_3065);
or U4177 (N_4177,N_3715,N_3718);
nor U4178 (N_4178,N_3651,N_3322);
nor U4179 (N_4179,N_3520,N_3172);
nand U4180 (N_4180,N_3114,N_3179);
nor U4181 (N_4181,N_3286,N_3226);
and U4182 (N_4182,N_3097,N_3075);
and U4183 (N_4183,N_3506,N_3391);
or U4184 (N_4184,N_3107,N_3018);
or U4185 (N_4185,N_3537,N_3254);
and U4186 (N_4186,N_3722,N_3184);
and U4187 (N_4187,N_3621,N_3351);
or U4188 (N_4188,N_3355,N_3738);
nand U4189 (N_4189,N_3168,N_3191);
or U4190 (N_4190,N_3179,N_3542);
or U4191 (N_4191,N_3261,N_3526);
nand U4192 (N_4192,N_3027,N_3176);
and U4193 (N_4193,N_3693,N_3273);
xnor U4194 (N_4194,N_3551,N_3038);
nor U4195 (N_4195,N_3540,N_3740);
xnor U4196 (N_4196,N_3285,N_3644);
nor U4197 (N_4197,N_3118,N_3256);
nand U4198 (N_4198,N_3534,N_3215);
nor U4199 (N_4199,N_3706,N_3722);
nand U4200 (N_4200,N_3544,N_3560);
and U4201 (N_4201,N_3345,N_3357);
nor U4202 (N_4202,N_3002,N_3082);
nor U4203 (N_4203,N_3697,N_3730);
nor U4204 (N_4204,N_3004,N_3281);
or U4205 (N_4205,N_3537,N_3026);
or U4206 (N_4206,N_3162,N_3229);
nor U4207 (N_4207,N_3544,N_3157);
or U4208 (N_4208,N_3714,N_3031);
and U4209 (N_4209,N_3168,N_3544);
nand U4210 (N_4210,N_3487,N_3366);
and U4211 (N_4211,N_3097,N_3155);
or U4212 (N_4212,N_3293,N_3214);
nor U4213 (N_4213,N_3468,N_3638);
and U4214 (N_4214,N_3272,N_3245);
and U4215 (N_4215,N_3584,N_3305);
nor U4216 (N_4216,N_3399,N_3388);
nor U4217 (N_4217,N_3356,N_3170);
nor U4218 (N_4218,N_3036,N_3219);
and U4219 (N_4219,N_3112,N_3366);
and U4220 (N_4220,N_3302,N_3614);
nand U4221 (N_4221,N_3152,N_3680);
or U4222 (N_4222,N_3215,N_3050);
and U4223 (N_4223,N_3262,N_3042);
nor U4224 (N_4224,N_3524,N_3426);
nand U4225 (N_4225,N_3027,N_3127);
and U4226 (N_4226,N_3201,N_3563);
and U4227 (N_4227,N_3068,N_3463);
nand U4228 (N_4228,N_3455,N_3249);
nand U4229 (N_4229,N_3711,N_3608);
xor U4230 (N_4230,N_3458,N_3276);
and U4231 (N_4231,N_3015,N_3686);
nor U4232 (N_4232,N_3173,N_3718);
or U4233 (N_4233,N_3267,N_3412);
nand U4234 (N_4234,N_3583,N_3085);
nor U4235 (N_4235,N_3144,N_3101);
and U4236 (N_4236,N_3412,N_3670);
and U4237 (N_4237,N_3667,N_3212);
nand U4238 (N_4238,N_3344,N_3215);
and U4239 (N_4239,N_3217,N_3516);
nand U4240 (N_4240,N_3671,N_3431);
xor U4241 (N_4241,N_3291,N_3012);
and U4242 (N_4242,N_3531,N_3034);
nor U4243 (N_4243,N_3659,N_3646);
or U4244 (N_4244,N_3579,N_3614);
and U4245 (N_4245,N_3546,N_3472);
and U4246 (N_4246,N_3279,N_3456);
nor U4247 (N_4247,N_3206,N_3452);
nand U4248 (N_4248,N_3725,N_3375);
nor U4249 (N_4249,N_3272,N_3257);
or U4250 (N_4250,N_3465,N_3337);
or U4251 (N_4251,N_3186,N_3721);
or U4252 (N_4252,N_3209,N_3200);
nand U4253 (N_4253,N_3074,N_3492);
and U4254 (N_4254,N_3083,N_3276);
or U4255 (N_4255,N_3634,N_3552);
nor U4256 (N_4256,N_3392,N_3748);
and U4257 (N_4257,N_3566,N_3355);
and U4258 (N_4258,N_3169,N_3229);
and U4259 (N_4259,N_3374,N_3515);
xor U4260 (N_4260,N_3529,N_3435);
and U4261 (N_4261,N_3221,N_3546);
or U4262 (N_4262,N_3564,N_3641);
or U4263 (N_4263,N_3530,N_3352);
nor U4264 (N_4264,N_3421,N_3098);
or U4265 (N_4265,N_3292,N_3467);
nor U4266 (N_4266,N_3558,N_3453);
nor U4267 (N_4267,N_3162,N_3385);
or U4268 (N_4268,N_3506,N_3286);
nand U4269 (N_4269,N_3335,N_3388);
nor U4270 (N_4270,N_3496,N_3298);
and U4271 (N_4271,N_3458,N_3611);
and U4272 (N_4272,N_3134,N_3056);
nand U4273 (N_4273,N_3568,N_3557);
nor U4274 (N_4274,N_3709,N_3356);
or U4275 (N_4275,N_3309,N_3607);
nor U4276 (N_4276,N_3747,N_3496);
and U4277 (N_4277,N_3719,N_3341);
xor U4278 (N_4278,N_3714,N_3422);
and U4279 (N_4279,N_3521,N_3107);
nand U4280 (N_4280,N_3560,N_3512);
and U4281 (N_4281,N_3392,N_3080);
nor U4282 (N_4282,N_3379,N_3323);
nand U4283 (N_4283,N_3475,N_3605);
nor U4284 (N_4284,N_3715,N_3261);
nand U4285 (N_4285,N_3251,N_3385);
nor U4286 (N_4286,N_3731,N_3475);
nor U4287 (N_4287,N_3712,N_3475);
nor U4288 (N_4288,N_3422,N_3139);
and U4289 (N_4289,N_3307,N_3437);
and U4290 (N_4290,N_3415,N_3163);
or U4291 (N_4291,N_3668,N_3546);
nor U4292 (N_4292,N_3176,N_3597);
nand U4293 (N_4293,N_3485,N_3265);
nand U4294 (N_4294,N_3362,N_3003);
and U4295 (N_4295,N_3170,N_3684);
or U4296 (N_4296,N_3728,N_3066);
and U4297 (N_4297,N_3007,N_3665);
and U4298 (N_4298,N_3508,N_3341);
and U4299 (N_4299,N_3081,N_3079);
and U4300 (N_4300,N_3487,N_3297);
nand U4301 (N_4301,N_3392,N_3562);
or U4302 (N_4302,N_3075,N_3185);
nor U4303 (N_4303,N_3525,N_3393);
or U4304 (N_4304,N_3295,N_3059);
and U4305 (N_4305,N_3107,N_3304);
and U4306 (N_4306,N_3444,N_3583);
nand U4307 (N_4307,N_3122,N_3501);
nand U4308 (N_4308,N_3518,N_3362);
and U4309 (N_4309,N_3375,N_3207);
or U4310 (N_4310,N_3239,N_3395);
nand U4311 (N_4311,N_3285,N_3716);
and U4312 (N_4312,N_3354,N_3175);
nand U4313 (N_4313,N_3585,N_3438);
nor U4314 (N_4314,N_3672,N_3675);
or U4315 (N_4315,N_3459,N_3694);
nand U4316 (N_4316,N_3626,N_3506);
nand U4317 (N_4317,N_3146,N_3045);
nand U4318 (N_4318,N_3300,N_3103);
nor U4319 (N_4319,N_3519,N_3483);
and U4320 (N_4320,N_3115,N_3641);
and U4321 (N_4321,N_3068,N_3203);
nor U4322 (N_4322,N_3157,N_3217);
nor U4323 (N_4323,N_3482,N_3359);
or U4324 (N_4324,N_3219,N_3234);
nor U4325 (N_4325,N_3641,N_3487);
nand U4326 (N_4326,N_3069,N_3185);
nand U4327 (N_4327,N_3634,N_3641);
and U4328 (N_4328,N_3582,N_3000);
nand U4329 (N_4329,N_3360,N_3185);
nand U4330 (N_4330,N_3478,N_3003);
or U4331 (N_4331,N_3458,N_3319);
nor U4332 (N_4332,N_3021,N_3178);
and U4333 (N_4333,N_3716,N_3289);
nand U4334 (N_4334,N_3668,N_3256);
nor U4335 (N_4335,N_3536,N_3651);
and U4336 (N_4336,N_3478,N_3141);
nor U4337 (N_4337,N_3264,N_3704);
nor U4338 (N_4338,N_3684,N_3161);
xor U4339 (N_4339,N_3359,N_3350);
or U4340 (N_4340,N_3333,N_3545);
or U4341 (N_4341,N_3459,N_3381);
nand U4342 (N_4342,N_3180,N_3019);
nor U4343 (N_4343,N_3047,N_3372);
nand U4344 (N_4344,N_3026,N_3334);
nand U4345 (N_4345,N_3428,N_3153);
or U4346 (N_4346,N_3714,N_3064);
nor U4347 (N_4347,N_3706,N_3040);
nand U4348 (N_4348,N_3232,N_3482);
nand U4349 (N_4349,N_3491,N_3168);
and U4350 (N_4350,N_3218,N_3100);
or U4351 (N_4351,N_3154,N_3346);
and U4352 (N_4352,N_3107,N_3067);
nand U4353 (N_4353,N_3008,N_3391);
nor U4354 (N_4354,N_3575,N_3186);
or U4355 (N_4355,N_3742,N_3737);
and U4356 (N_4356,N_3360,N_3201);
or U4357 (N_4357,N_3143,N_3093);
or U4358 (N_4358,N_3131,N_3291);
or U4359 (N_4359,N_3705,N_3168);
nor U4360 (N_4360,N_3126,N_3472);
nand U4361 (N_4361,N_3542,N_3010);
nor U4362 (N_4362,N_3592,N_3574);
nand U4363 (N_4363,N_3373,N_3650);
nand U4364 (N_4364,N_3468,N_3695);
nand U4365 (N_4365,N_3663,N_3571);
nand U4366 (N_4366,N_3470,N_3115);
and U4367 (N_4367,N_3547,N_3262);
nand U4368 (N_4368,N_3107,N_3019);
or U4369 (N_4369,N_3420,N_3251);
nor U4370 (N_4370,N_3729,N_3029);
and U4371 (N_4371,N_3489,N_3740);
nor U4372 (N_4372,N_3277,N_3477);
and U4373 (N_4373,N_3509,N_3715);
or U4374 (N_4374,N_3497,N_3215);
nor U4375 (N_4375,N_3018,N_3166);
and U4376 (N_4376,N_3610,N_3406);
or U4377 (N_4377,N_3425,N_3330);
and U4378 (N_4378,N_3191,N_3496);
nor U4379 (N_4379,N_3434,N_3660);
nand U4380 (N_4380,N_3347,N_3356);
nor U4381 (N_4381,N_3162,N_3340);
nor U4382 (N_4382,N_3121,N_3038);
nor U4383 (N_4383,N_3050,N_3570);
or U4384 (N_4384,N_3380,N_3647);
or U4385 (N_4385,N_3019,N_3101);
nand U4386 (N_4386,N_3528,N_3409);
and U4387 (N_4387,N_3608,N_3084);
nor U4388 (N_4388,N_3108,N_3151);
nand U4389 (N_4389,N_3487,N_3096);
nand U4390 (N_4390,N_3559,N_3036);
nor U4391 (N_4391,N_3070,N_3187);
and U4392 (N_4392,N_3035,N_3031);
or U4393 (N_4393,N_3615,N_3242);
nand U4394 (N_4394,N_3484,N_3577);
or U4395 (N_4395,N_3389,N_3083);
and U4396 (N_4396,N_3380,N_3746);
nand U4397 (N_4397,N_3078,N_3002);
nor U4398 (N_4398,N_3280,N_3742);
nand U4399 (N_4399,N_3384,N_3494);
or U4400 (N_4400,N_3101,N_3520);
nand U4401 (N_4401,N_3244,N_3515);
and U4402 (N_4402,N_3008,N_3039);
and U4403 (N_4403,N_3217,N_3721);
and U4404 (N_4404,N_3737,N_3468);
nor U4405 (N_4405,N_3744,N_3213);
nor U4406 (N_4406,N_3370,N_3434);
nor U4407 (N_4407,N_3233,N_3287);
nand U4408 (N_4408,N_3697,N_3671);
nand U4409 (N_4409,N_3714,N_3745);
nor U4410 (N_4410,N_3715,N_3696);
and U4411 (N_4411,N_3562,N_3654);
and U4412 (N_4412,N_3059,N_3442);
or U4413 (N_4413,N_3131,N_3477);
nand U4414 (N_4414,N_3698,N_3701);
and U4415 (N_4415,N_3552,N_3110);
or U4416 (N_4416,N_3464,N_3365);
nand U4417 (N_4417,N_3242,N_3114);
nand U4418 (N_4418,N_3462,N_3480);
or U4419 (N_4419,N_3152,N_3621);
and U4420 (N_4420,N_3293,N_3191);
nand U4421 (N_4421,N_3472,N_3564);
nand U4422 (N_4422,N_3124,N_3727);
and U4423 (N_4423,N_3513,N_3061);
nand U4424 (N_4424,N_3510,N_3617);
or U4425 (N_4425,N_3724,N_3224);
nand U4426 (N_4426,N_3144,N_3513);
nor U4427 (N_4427,N_3165,N_3494);
nor U4428 (N_4428,N_3017,N_3007);
and U4429 (N_4429,N_3451,N_3716);
and U4430 (N_4430,N_3573,N_3231);
and U4431 (N_4431,N_3212,N_3442);
nor U4432 (N_4432,N_3124,N_3167);
nor U4433 (N_4433,N_3238,N_3704);
and U4434 (N_4434,N_3098,N_3558);
and U4435 (N_4435,N_3404,N_3505);
nand U4436 (N_4436,N_3296,N_3092);
or U4437 (N_4437,N_3006,N_3363);
nand U4438 (N_4438,N_3601,N_3103);
xnor U4439 (N_4439,N_3231,N_3214);
and U4440 (N_4440,N_3072,N_3245);
nor U4441 (N_4441,N_3166,N_3217);
nand U4442 (N_4442,N_3142,N_3507);
or U4443 (N_4443,N_3139,N_3671);
or U4444 (N_4444,N_3040,N_3328);
nor U4445 (N_4445,N_3614,N_3112);
or U4446 (N_4446,N_3299,N_3428);
nor U4447 (N_4447,N_3465,N_3600);
nand U4448 (N_4448,N_3559,N_3023);
nor U4449 (N_4449,N_3300,N_3195);
or U4450 (N_4450,N_3576,N_3629);
or U4451 (N_4451,N_3404,N_3615);
nor U4452 (N_4452,N_3299,N_3282);
nor U4453 (N_4453,N_3741,N_3544);
and U4454 (N_4454,N_3577,N_3672);
nand U4455 (N_4455,N_3232,N_3636);
nand U4456 (N_4456,N_3016,N_3419);
and U4457 (N_4457,N_3658,N_3245);
xor U4458 (N_4458,N_3747,N_3182);
and U4459 (N_4459,N_3729,N_3399);
or U4460 (N_4460,N_3671,N_3649);
and U4461 (N_4461,N_3376,N_3203);
or U4462 (N_4462,N_3511,N_3084);
or U4463 (N_4463,N_3742,N_3304);
and U4464 (N_4464,N_3084,N_3193);
and U4465 (N_4465,N_3651,N_3421);
nor U4466 (N_4466,N_3412,N_3724);
nand U4467 (N_4467,N_3369,N_3713);
nor U4468 (N_4468,N_3643,N_3251);
or U4469 (N_4469,N_3530,N_3713);
or U4470 (N_4470,N_3281,N_3168);
nor U4471 (N_4471,N_3547,N_3692);
and U4472 (N_4472,N_3228,N_3240);
or U4473 (N_4473,N_3401,N_3392);
nor U4474 (N_4474,N_3302,N_3250);
nor U4475 (N_4475,N_3032,N_3276);
and U4476 (N_4476,N_3109,N_3645);
or U4477 (N_4477,N_3412,N_3011);
nor U4478 (N_4478,N_3102,N_3008);
nor U4479 (N_4479,N_3154,N_3385);
xnor U4480 (N_4480,N_3333,N_3010);
and U4481 (N_4481,N_3098,N_3620);
nor U4482 (N_4482,N_3013,N_3113);
nor U4483 (N_4483,N_3349,N_3007);
nand U4484 (N_4484,N_3189,N_3221);
nand U4485 (N_4485,N_3215,N_3059);
nand U4486 (N_4486,N_3589,N_3104);
or U4487 (N_4487,N_3419,N_3448);
or U4488 (N_4488,N_3575,N_3696);
or U4489 (N_4489,N_3419,N_3650);
nand U4490 (N_4490,N_3165,N_3581);
and U4491 (N_4491,N_3633,N_3351);
and U4492 (N_4492,N_3638,N_3353);
and U4493 (N_4493,N_3218,N_3713);
nand U4494 (N_4494,N_3394,N_3369);
or U4495 (N_4495,N_3603,N_3000);
or U4496 (N_4496,N_3304,N_3711);
and U4497 (N_4497,N_3111,N_3452);
nand U4498 (N_4498,N_3432,N_3451);
nand U4499 (N_4499,N_3312,N_3137);
nor U4500 (N_4500,N_3984,N_3950);
or U4501 (N_4501,N_3999,N_4152);
nor U4502 (N_4502,N_3762,N_3935);
and U4503 (N_4503,N_4106,N_3894);
nand U4504 (N_4504,N_4038,N_3995);
nand U4505 (N_4505,N_4217,N_3771);
nor U4506 (N_4506,N_3873,N_4225);
nor U4507 (N_4507,N_3792,N_4272);
and U4508 (N_4508,N_3842,N_4119);
and U4509 (N_4509,N_4389,N_4252);
nand U4510 (N_4510,N_4329,N_4056);
nor U4511 (N_4511,N_4428,N_3912);
or U4512 (N_4512,N_4249,N_4216);
nor U4513 (N_4513,N_3848,N_4312);
and U4514 (N_4514,N_3907,N_4009);
or U4515 (N_4515,N_3952,N_4087);
and U4516 (N_4516,N_4364,N_3899);
and U4517 (N_4517,N_3858,N_4221);
nor U4518 (N_4518,N_4324,N_3925);
and U4519 (N_4519,N_4308,N_4295);
nand U4520 (N_4520,N_3875,N_4450);
nor U4521 (N_4521,N_3835,N_4292);
nor U4522 (N_4522,N_4062,N_3856);
and U4523 (N_4523,N_4394,N_3754);
nand U4524 (N_4524,N_3919,N_4229);
nor U4525 (N_4525,N_4403,N_4137);
and U4526 (N_4526,N_4071,N_4391);
nand U4527 (N_4527,N_4343,N_4218);
and U4528 (N_4528,N_3906,N_4165);
nor U4529 (N_4529,N_3819,N_4412);
or U4530 (N_4530,N_4069,N_4478);
or U4531 (N_4531,N_4299,N_4141);
or U4532 (N_4532,N_4184,N_4427);
or U4533 (N_4533,N_4273,N_3934);
nand U4534 (N_4534,N_3964,N_4086);
and U4535 (N_4535,N_4396,N_3868);
nand U4536 (N_4536,N_3854,N_4146);
and U4537 (N_4537,N_4489,N_3800);
and U4538 (N_4538,N_3755,N_4493);
nand U4539 (N_4539,N_4468,N_4352);
or U4540 (N_4540,N_3832,N_4175);
nand U4541 (N_4541,N_4193,N_4134);
nor U4542 (N_4542,N_4104,N_4109);
nor U4543 (N_4543,N_3824,N_4178);
or U4544 (N_4544,N_4487,N_3917);
and U4545 (N_4545,N_4154,N_4199);
or U4546 (N_4546,N_3987,N_3794);
nand U4547 (N_4547,N_3852,N_3847);
or U4548 (N_4548,N_3797,N_4264);
nand U4549 (N_4549,N_4317,N_4397);
or U4550 (N_4550,N_3833,N_4390);
and U4551 (N_4551,N_4017,N_4052);
or U4552 (N_4552,N_4213,N_4328);
nand U4553 (N_4553,N_3876,N_4441);
or U4554 (N_4554,N_4307,N_4118);
nand U4555 (N_4555,N_3905,N_3983);
and U4556 (N_4556,N_4383,N_4142);
and U4557 (N_4557,N_4456,N_3978);
and U4558 (N_4558,N_4274,N_3838);
and U4559 (N_4559,N_3979,N_4382);
or U4560 (N_4560,N_3877,N_4262);
and U4561 (N_4561,N_3770,N_4344);
nand U4562 (N_4562,N_4325,N_4004);
nand U4563 (N_4563,N_3805,N_4173);
nor U4564 (N_4564,N_4475,N_4244);
nor U4565 (N_4565,N_3924,N_4181);
xor U4566 (N_4566,N_3760,N_4305);
or U4567 (N_4567,N_3844,N_4153);
nor U4568 (N_4568,N_4018,N_4346);
nand U4569 (N_4569,N_4138,N_4198);
or U4570 (N_4570,N_4445,N_3765);
nand U4571 (N_4571,N_3779,N_4319);
nor U4572 (N_4572,N_3926,N_3892);
nand U4573 (N_4573,N_4304,N_4446);
nor U4574 (N_4574,N_4415,N_4437);
nor U4575 (N_4575,N_3870,N_4379);
and U4576 (N_4576,N_4370,N_4356);
nand U4577 (N_4577,N_4406,N_3915);
nand U4578 (N_4578,N_4032,N_3809);
or U4579 (N_4579,N_3993,N_3871);
nor U4580 (N_4580,N_3862,N_4014);
nor U4581 (N_4581,N_4250,N_3831);
or U4582 (N_4582,N_4296,N_4030);
and U4583 (N_4583,N_3956,N_4191);
xor U4584 (N_4584,N_4372,N_3945);
or U4585 (N_4585,N_4036,N_4245);
nand U4586 (N_4586,N_3961,N_4349);
nand U4587 (N_4587,N_4484,N_3982);
nor U4588 (N_4588,N_4368,N_4340);
or U4589 (N_4589,N_4101,N_4151);
nand U4590 (N_4590,N_4290,N_4347);
and U4591 (N_4591,N_3895,N_4341);
or U4592 (N_4592,N_3752,N_3767);
nand U4593 (N_4593,N_4462,N_4410);
nand U4594 (N_4594,N_3949,N_4012);
nand U4595 (N_4595,N_3773,N_4129);
nand U4596 (N_4596,N_4298,N_4265);
nand U4597 (N_4597,N_4208,N_4465);
and U4598 (N_4598,N_4123,N_4496);
or U4599 (N_4599,N_4192,N_4070);
nor U4600 (N_4600,N_4238,N_3841);
nor U4601 (N_4601,N_3750,N_4337);
and U4602 (N_4602,N_4385,N_4286);
nor U4603 (N_4603,N_4327,N_4477);
nand U4604 (N_4604,N_4033,N_4490);
or U4605 (N_4605,N_4065,N_4015);
nor U4606 (N_4606,N_3859,N_3953);
or U4607 (N_4607,N_3867,N_4078);
nor U4608 (N_4608,N_3929,N_4331);
nand U4609 (N_4609,N_4064,N_3944);
nand U4610 (N_4610,N_3855,N_4203);
nor U4611 (N_4611,N_3843,N_3786);
nor U4612 (N_4612,N_4001,N_4114);
and U4613 (N_4613,N_4499,N_3845);
nand U4614 (N_4614,N_4369,N_4016);
or U4615 (N_4615,N_4103,N_3897);
nand U4616 (N_4616,N_4417,N_4281);
nor U4617 (N_4617,N_3849,N_4285);
nand U4618 (N_4618,N_3946,N_4117);
nor U4619 (N_4619,N_4342,N_3942);
nor U4620 (N_4620,N_3814,N_4357);
xor U4621 (N_4621,N_4059,N_4149);
and U4622 (N_4622,N_4425,N_3801);
nand U4623 (N_4623,N_4194,N_3902);
nor U4624 (N_4624,N_4419,N_4276);
and U4625 (N_4625,N_4362,N_3903);
nor U4626 (N_4626,N_4201,N_4143);
nand U4627 (N_4627,N_4454,N_4429);
nand U4628 (N_4628,N_4474,N_4303);
or U4629 (N_4629,N_4091,N_3866);
and U4630 (N_4630,N_4309,N_4237);
or U4631 (N_4631,N_4387,N_4377);
nor U4632 (N_4632,N_4183,N_3980);
and U4633 (N_4633,N_4472,N_3932);
nor U4634 (N_4634,N_4310,N_4363);
or U4635 (N_4635,N_4093,N_4076);
nand U4636 (N_4636,N_3766,N_4224);
and U4637 (N_4637,N_3799,N_3783);
and U4638 (N_4638,N_4270,N_4266);
nand U4639 (N_4639,N_4359,N_4081);
nor U4640 (N_4640,N_3985,N_4409);
nor U4641 (N_4641,N_4322,N_4414);
or U4642 (N_4642,N_3850,N_3857);
nor U4643 (N_4643,N_4162,N_4278);
or U4644 (N_4644,N_3840,N_4302);
nor U4645 (N_4645,N_4133,N_4206);
nand U4646 (N_4646,N_4088,N_4044);
and U4647 (N_4647,N_4443,N_4430);
nand U4648 (N_4648,N_4063,N_4455);
nor U4649 (N_4649,N_3878,N_4386);
nand U4650 (N_4650,N_4200,N_3991);
and U4651 (N_4651,N_3827,N_4046);
nand U4652 (N_4652,N_3764,N_3986);
or U4653 (N_4653,N_4355,N_3828);
nand U4654 (N_4654,N_3921,N_4147);
nand U4655 (N_4655,N_3811,N_3763);
or U4656 (N_4656,N_4043,N_3933);
and U4657 (N_4657,N_3943,N_4228);
and U4658 (N_4658,N_3768,N_4116);
nand U4659 (N_4659,N_3772,N_4318);
nand U4660 (N_4660,N_3791,N_4057);
nand U4661 (N_4661,N_3777,N_3804);
or U4662 (N_4662,N_4140,N_4423);
nor U4663 (N_4663,N_4073,N_3774);
nand U4664 (N_4664,N_4395,N_4246);
nand U4665 (N_4665,N_4452,N_4481);
and U4666 (N_4666,N_4447,N_4282);
or U4667 (N_4667,N_3911,N_4061);
nand U4668 (N_4668,N_4314,N_4189);
nand U4669 (N_4669,N_3822,N_3884);
and U4670 (N_4670,N_3969,N_4185);
or U4671 (N_4671,N_4321,N_4239);
and U4672 (N_4672,N_3853,N_4156);
nor U4673 (N_4673,N_3893,N_4361);
nor U4674 (N_4674,N_4060,N_4011);
and U4675 (N_4675,N_3823,N_4214);
or U4676 (N_4676,N_3837,N_4433);
nand U4677 (N_4677,N_3789,N_4035);
or U4678 (N_4678,N_4451,N_4345);
or U4679 (N_4679,N_4127,N_4440);
and U4680 (N_4680,N_3780,N_4074);
and U4681 (N_4681,N_4072,N_4420);
or U4682 (N_4682,N_4082,N_4145);
and U4683 (N_4683,N_4393,N_4097);
and U4684 (N_4684,N_3756,N_3790);
nor U4685 (N_4685,N_4180,N_4126);
and U4686 (N_4686,N_3761,N_4461);
nor U4687 (N_4687,N_4411,N_4005);
and U4688 (N_4688,N_4269,N_4223);
nor U4689 (N_4689,N_3890,N_4172);
nor U4690 (N_4690,N_4486,N_4373);
nand U4691 (N_4691,N_4287,N_4247);
nor U4692 (N_4692,N_4381,N_4111);
nand U4693 (N_4693,N_3927,N_4029);
nor U4694 (N_4694,N_4048,N_4431);
and U4695 (N_4695,N_4444,N_4332);
nand U4696 (N_4696,N_3839,N_4421);
nand U4697 (N_4697,N_4339,N_4284);
nand U4698 (N_4698,N_3948,N_4166);
and U4699 (N_4699,N_4459,N_4148);
or U4700 (N_4700,N_4100,N_3990);
and U4701 (N_4701,N_4460,N_4248);
and U4702 (N_4702,N_4023,N_3796);
and U4703 (N_4703,N_4480,N_4350);
or U4704 (N_4704,N_4034,N_4055);
nand U4705 (N_4705,N_3975,N_4215);
nand U4706 (N_4706,N_4089,N_4066);
or U4707 (N_4707,N_4413,N_3938);
nor U4708 (N_4708,N_4333,N_4279);
or U4709 (N_4709,N_4259,N_4235);
nor U4710 (N_4710,N_4358,N_3787);
nand U4711 (N_4711,N_4476,N_3834);
and U4712 (N_4712,N_4351,N_4267);
nand U4713 (N_4713,N_4027,N_3775);
and U4714 (N_4714,N_3863,N_3989);
or U4715 (N_4715,N_4187,N_3886);
or U4716 (N_4716,N_4316,N_3898);
and U4717 (N_4717,N_4054,N_4376);
or U4718 (N_4718,N_3996,N_4040);
nor U4719 (N_4719,N_3782,N_4367);
nand U4720 (N_4720,N_4479,N_3891);
or U4721 (N_4721,N_4320,N_4261);
nand U4722 (N_4722,N_4079,N_4050);
nand U4723 (N_4723,N_3883,N_3901);
nor U4724 (N_4724,N_3920,N_3807);
xnor U4725 (N_4725,N_4045,N_4485);
nor U4726 (N_4726,N_3810,N_4469);
and U4727 (N_4727,N_4232,N_4186);
nor U4728 (N_4728,N_4159,N_4300);
nor U4729 (N_4729,N_4330,N_4039);
and U4730 (N_4730,N_4492,N_4360);
nand U4731 (N_4731,N_3851,N_4157);
or U4732 (N_4732,N_4418,N_4006);
nand U4733 (N_4733,N_4084,N_4002);
and U4734 (N_4734,N_4466,N_4301);
nand U4735 (N_4735,N_4135,N_4242);
nand U4736 (N_4736,N_3923,N_4399);
nor U4737 (N_4737,N_4098,N_4096);
or U4738 (N_4738,N_4435,N_4068);
or U4739 (N_4739,N_4121,N_4392);
and U4740 (N_4740,N_4222,N_3882);
nand U4741 (N_4741,N_4306,N_4113);
or U4742 (N_4742,N_3815,N_4211);
nand U4743 (N_4743,N_4275,N_3812);
nor U4744 (N_4744,N_3928,N_4384);
nand U4745 (N_4745,N_4220,N_4230);
or U4746 (N_4746,N_4488,N_4007);
nand U4747 (N_4747,N_3997,N_4110);
or U4748 (N_4748,N_4402,N_3861);
nor U4749 (N_4749,N_4075,N_4263);
or U4750 (N_4750,N_4058,N_4374);
or U4751 (N_4751,N_3830,N_4457);
nand U4752 (N_4752,N_3802,N_3860);
nand U4753 (N_4753,N_4227,N_4254);
and U4754 (N_4754,N_4095,N_4464);
nor U4755 (N_4755,N_4131,N_4080);
and U4756 (N_4756,N_3962,N_4139);
nor U4757 (N_4757,N_3785,N_3806);
and U4758 (N_4758,N_3931,N_3872);
and U4759 (N_4759,N_4171,N_4000);
and U4760 (N_4760,N_4256,N_4439);
or U4761 (N_4761,N_4371,N_4378);
and U4762 (N_4762,N_4196,N_4416);
nand U4763 (N_4763,N_4102,N_3798);
and U4764 (N_4764,N_3971,N_3753);
or U4765 (N_4765,N_3821,N_4204);
or U4766 (N_4766,N_3769,N_3900);
and U4767 (N_4767,N_4335,N_4195);
and U4768 (N_4768,N_4354,N_4260);
nand U4769 (N_4769,N_3817,N_3820);
nand U4770 (N_4770,N_4231,N_4280);
nor U4771 (N_4771,N_3757,N_4164);
and U4772 (N_4772,N_3930,N_3960);
nor U4773 (N_4773,N_3947,N_3973);
nand U4774 (N_4774,N_3788,N_4365);
nand U4775 (N_4775,N_4255,N_4241);
nor U4776 (N_4776,N_4253,N_4041);
or U4777 (N_4777,N_4473,N_3951);
nor U4778 (N_4778,N_4449,N_3992);
or U4779 (N_4779,N_4167,N_3776);
or U4780 (N_4780,N_3808,N_3887);
and U4781 (N_4781,N_4202,N_4179);
nand U4782 (N_4782,N_4190,N_4083);
nor U4783 (N_4783,N_4122,N_3869);
nand U4784 (N_4784,N_4026,N_3977);
and U4785 (N_4785,N_4283,N_4426);
or U4786 (N_4786,N_3998,N_4010);
and U4787 (N_4787,N_4277,N_3888);
nor U4788 (N_4788,N_3988,N_4037);
and U4789 (N_4789,N_3994,N_4482);
or U4790 (N_4790,N_4442,N_4471);
or U4791 (N_4791,N_4182,N_4257);
and U4792 (N_4792,N_3959,N_4051);
or U4793 (N_4793,N_3829,N_3758);
and U4794 (N_4794,N_4019,N_4107);
and U4795 (N_4795,N_4125,N_3965);
or U4796 (N_4796,N_4049,N_4353);
and U4797 (N_4797,N_4483,N_4124);
nor U4798 (N_4798,N_4021,N_4132);
and U4799 (N_4799,N_4115,N_3864);
or U4800 (N_4800,N_4470,N_3881);
nor U4801 (N_4801,N_3968,N_4174);
or U4802 (N_4802,N_4158,N_4022);
nor U4803 (N_4803,N_4348,N_4020);
and U4804 (N_4804,N_4226,N_4336);
nand U4805 (N_4805,N_4494,N_4047);
nor U4806 (N_4806,N_3913,N_4144);
or U4807 (N_4807,N_4099,N_3922);
and U4808 (N_4808,N_4407,N_3937);
nand U4809 (N_4809,N_4130,N_4497);
nor U4810 (N_4810,N_3910,N_4294);
nand U4811 (N_4811,N_3879,N_4150);
nand U4812 (N_4812,N_4170,N_4366);
nor U4813 (N_4813,N_4268,N_3936);
nand U4814 (N_4814,N_4326,N_4271);
nor U4815 (N_4815,N_4094,N_4067);
nand U4816 (N_4816,N_4013,N_4297);
or U4817 (N_4817,N_4219,N_4334);
nor U4818 (N_4818,N_3974,N_4236);
nand U4819 (N_4819,N_4136,N_4053);
and U4820 (N_4820,N_4205,N_3751);
nand U4821 (N_4821,N_3958,N_3889);
and U4822 (N_4822,N_4498,N_3826);
nor U4823 (N_4823,N_4212,N_4008);
and U4824 (N_4824,N_4042,N_4400);
and U4825 (N_4825,N_3954,N_4380);
and U4826 (N_4826,N_4176,N_4491);
nand U4827 (N_4827,N_4240,N_3904);
nand U4828 (N_4828,N_4338,N_4289);
and U4829 (N_4829,N_4436,N_3909);
nor U4830 (N_4830,N_3836,N_3976);
or U4831 (N_4831,N_4120,N_4168);
nand U4832 (N_4832,N_4243,N_4422);
nand U4833 (N_4833,N_4405,N_4424);
nor U4834 (N_4834,N_4288,N_4209);
nor U4835 (N_4835,N_3781,N_3880);
or U4836 (N_4836,N_3963,N_3865);
xnor U4837 (N_4837,N_4434,N_4432);
or U4838 (N_4838,N_4177,N_4258);
and U4839 (N_4839,N_4251,N_4105);
xnor U4840 (N_4840,N_3896,N_4090);
and U4841 (N_4841,N_3955,N_4025);
and U4842 (N_4842,N_4453,N_3966);
nor U4843 (N_4843,N_3813,N_3972);
and U4844 (N_4844,N_4401,N_4315);
and U4845 (N_4845,N_3981,N_3825);
and U4846 (N_4846,N_4323,N_4311);
and U4847 (N_4847,N_3940,N_3967);
and U4848 (N_4848,N_3957,N_3914);
nor U4849 (N_4849,N_4404,N_4388);
or U4850 (N_4850,N_4112,N_3939);
and U4851 (N_4851,N_3970,N_4234);
and U4852 (N_4852,N_3908,N_4207);
nor U4853 (N_4853,N_3795,N_3846);
or U4854 (N_4854,N_3784,N_4161);
or U4855 (N_4855,N_4291,N_3941);
nor U4856 (N_4856,N_4210,N_4458);
nand U4857 (N_4857,N_3818,N_4375);
or U4858 (N_4858,N_3793,N_4438);
and U4859 (N_4859,N_4408,N_3874);
and U4860 (N_4860,N_4233,N_4092);
and U4861 (N_4861,N_4160,N_4031);
nor U4862 (N_4862,N_3778,N_4028);
nor U4863 (N_4863,N_4108,N_4003);
or U4864 (N_4864,N_4188,N_4128);
and U4865 (N_4865,N_3803,N_3916);
and U4866 (N_4866,N_4169,N_4197);
or U4867 (N_4867,N_4313,N_4495);
and U4868 (N_4868,N_4398,N_4293);
nor U4869 (N_4869,N_4077,N_4463);
or U4870 (N_4870,N_3918,N_3816);
and U4871 (N_4871,N_4163,N_4024);
nor U4872 (N_4872,N_3885,N_3759);
or U4873 (N_4873,N_4155,N_4448);
nand U4874 (N_4874,N_4085,N_4467);
and U4875 (N_4875,N_4161,N_3931);
or U4876 (N_4876,N_3910,N_4202);
nand U4877 (N_4877,N_4026,N_3819);
or U4878 (N_4878,N_4182,N_4238);
nor U4879 (N_4879,N_4100,N_4389);
nor U4880 (N_4880,N_4273,N_4182);
and U4881 (N_4881,N_4287,N_4339);
nor U4882 (N_4882,N_4184,N_4239);
nand U4883 (N_4883,N_4490,N_4109);
and U4884 (N_4884,N_4168,N_4169);
or U4885 (N_4885,N_4081,N_3759);
or U4886 (N_4886,N_4262,N_4466);
nand U4887 (N_4887,N_3768,N_4387);
or U4888 (N_4888,N_4201,N_3831);
and U4889 (N_4889,N_4261,N_3856);
nor U4890 (N_4890,N_3915,N_3965);
nor U4891 (N_4891,N_4150,N_3959);
and U4892 (N_4892,N_4207,N_4336);
and U4893 (N_4893,N_4017,N_4330);
nor U4894 (N_4894,N_3780,N_3997);
or U4895 (N_4895,N_4459,N_3932);
and U4896 (N_4896,N_4464,N_4128);
nand U4897 (N_4897,N_4314,N_3822);
nand U4898 (N_4898,N_4498,N_4215);
and U4899 (N_4899,N_4054,N_3960);
and U4900 (N_4900,N_3854,N_4270);
nor U4901 (N_4901,N_4179,N_3800);
nand U4902 (N_4902,N_4257,N_4362);
and U4903 (N_4903,N_3884,N_3847);
and U4904 (N_4904,N_4450,N_4433);
or U4905 (N_4905,N_4038,N_4421);
and U4906 (N_4906,N_3837,N_4365);
and U4907 (N_4907,N_4230,N_3849);
and U4908 (N_4908,N_4194,N_3853);
nor U4909 (N_4909,N_4182,N_3760);
nor U4910 (N_4910,N_4226,N_4129);
and U4911 (N_4911,N_4429,N_3955);
nand U4912 (N_4912,N_3888,N_3880);
or U4913 (N_4913,N_3804,N_4453);
and U4914 (N_4914,N_4319,N_4177);
nand U4915 (N_4915,N_4354,N_4075);
nor U4916 (N_4916,N_4324,N_4499);
or U4917 (N_4917,N_4480,N_3796);
nor U4918 (N_4918,N_3981,N_4168);
nor U4919 (N_4919,N_3873,N_4035);
nand U4920 (N_4920,N_4111,N_4089);
nor U4921 (N_4921,N_3952,N_4471);
or U4922 (N_4922,N_3782,N_4044);
nor U4923 (N_4923,N_3862,N_4197);
xor U4924 (N_4924,N_4410,N_4478);
and U4925 (N_4925,N_3957,N_4141);
nand U4926 (N_4926,N_4439,N_4238);
or U4927 (N_4927,N_4158,N_4330);
and U4928 (N_4928,N_3913,N_4476);
nand U4929 (N_4929,N_4042,N_3858);
and U4930 (N_4930,N_4491,N_4041);
xnor U4931 (N_4931,N_4124,N_3938);
or U4932 (N_4932,N_4347,N_4206);
and U4933 (N_4933,N_3794,N_4236);
and U4934 (N_4934,N_3865,N_4306);
nand U4935 (N_4935,N_3779,N_3938);
or U4936 (N_4936,N_4394,N_4378);
or U4937 (N_4937,N_4188,N_4280);
and U4938 (N_4938,N_4004,N_4184);
nor U4939 (N_4939,N_4360,N_4154);
nor U4940 (N_4940,N_3818,N_4456);
nand U4941 (N_4941,N_4160,N_4084);
and U4942 (N_4942,N_3851,N_4062);
or U4943 (N_4943,N_3899,N_4114);
nand U4944 (N_4944,N_3821,N_3790);
nor U4945 (N_4945,N_4040,N_3769);
or U4946 (N_4946,N_3997,N_3902);
nor U4947 (N_4947,N_4129,N_3900);
nand U4948 (N_4948,N_3964,N_4360);
nor U4949 (N_4949,N_3827,N_4401);
and U4950 (N_4950,N_4384,N_3983);
or U4951 (N_4951,N_4023,N_4406);
or U4952 (N_4952,N_4180,N_4424);
nand U4953 (N_4953,N_4290,N_4475);
nor U4954 (N_4954,N_4404,N_4166);
nand U4955 (N_4955,N_4028,N_4374);
or U4956 (N_4956,N_4156,N_4102);
nand U4957 (N_4957,N_4257,N_4261);
nor U4958 (N_4958,N_4306,N_4441);
or U4959 (N_4959,N_3780,N_3943);
or U4960 (N_4960,N_4197,N_4087);
nor U4961 (N_4961,N_3892,N_4272);
or U4962 (N_4962,N_4113,N_3805);
or U4963 (N_4963,N_4331,N_4210);
or U4964 (N_4964,N_3778,N_3785);
nor U4965 (N_4965,N_4445,N_4314);
nand U4966 (N_4966,N_3889,N_3796);
and U4967 (N_4967,N_4244,N_4358);
nor U4968 (N_4968,N_3823,N_4237);
nand U4969 (N_4969,N_4284,N_3915);
nand U4970 (N_4970,N_4272,N_3982);
nand U4971 (N_4971,N_4240,N_4145);
nand U4972 (N_4972,N_3827,N_4342);
and U4973 (N_4973,N_4423,N_3979);
or U4974 (N_4974,N_4360,N_4393);
nand U4975 (N_4975,N_4195,N_4018);
or U4976 (N_4976,N_4446,N_4383);
nand U4977 (N_4977,N_4317,N_4192);
or U4978 (N_4978,N_4369,N_4298);
and U4979 (N_4979,N_3939,N_3856);
nor U4980 (N_4980,N_4475,N_3755);
nand U4981 (N_4981,N_3934,N_4436);
or U4982 (N_4982,N_3989,N_4083);
nor U4983 (N_4983,N_3894,N_3830);
xnor U4984 (N_4984,N_3892,N_4197);
and U4985 (N_4985,N_3759,N_4441);
nand U4986 (N_4986,N_4255,N_4387);
or U4987 (N_4987,N_4192,N_3863);
nand U4988 (N_4988,N_4129,N_3753);
and U4989 (N_4989,N_4374,N_4005);
and U4990 (N_4990,N_3787,N_3838);
nor U4991 (N_4991,N_3939,N_4027);
nor U4992 (N_4992,N_4262,N_3847);
and U4993 (N_4993,N_3755,N_4336);
or U4994 (N_4994,N_4036,N_3998);
nand U4995 (N_4995,N_4217,N_4048);
and U4996 (N_4996,N_4292,N_4408);
nand U4997 (N_4997,N_3936,N_4185);
and U4998 (N_4998,N_3829,N_3949);
nor U4999 (N_4999,N_4372,N_3761);
nor U5000 (N_5000,N_3764,N_4129);
or U5001 (N_5001,N_4184,N_3862);
nand U5002 (N_5002,N_3775,N_4378);
nand U5003 (N_5003,N_4350,N_4160);
or U5004 (N_5004,N_3758,N_3825);
nand U5005 (N_5005,N_4358,N_4004);
xor U5006 (N_5006,N_4348,N_4190);
and U5007 (N_5007,N_4221,N_3760);
nor U5008 (N_5008,N_4393,N_4084);
nand U5009 (N_5009,N_4021,N_4204);
or U5010 (N_5010,N_3937,N_4318);
and U5011 (N_5011,N_4167,N_4359);
nand U5012 (N_5012,N_3816,N_3825);
nand U5013 (N_5013,N_4340,N_4232);
or U5014 (N_5014,N_4212,N_3849);
and U5015 (N_5015,N_4004,N_4243);
or U5016 (N_5016,N_4450,N_4118);
or U5017 (N_5017,N_3941,N_4466);
nand U5018 (N_5018,N_3811,N_4357);
nor U5019 (N_5019,N_4366,N_3798);
nor U5020 (N_5020,N_4480,N_4340);
or U5021 (N_5021,N_4071,N_3755);
nand U5022 (N_5022,N_3916,N_3768);
or U5023 (N_5023,N_4265,N_4334);
or U5024 (N_5024,N_4444,N_4312);
nor U5025 (N_5025,N_3859,N_3813);
nand U5026 (N_5026,N_3848,N_3940);
nor U5027 (N_5027,N_4036,N_4166);
nand U5028 (N_5028,N_4091,N_3964);
nand U5029 (N_5029,N_4068,N_4477);
nand U5030 (N_5030,N_4287,N_4499);
nand U5031 (N_5031,N_3854,N_4425);
nor U5032 (N_5032,N_4032,N_4305);
nor U5033 (N_5033,N_4302,N_4008);
and U5034 (N_5034,N_4108,N_4417);
or U5035 (N_5035,N_4372,N_4358);
and U5036 (N_5036,N_4453,N_3790);
or U5037 (N_5037,N_4261,N_4253);
nor U5038 (N_5038,N_4137,N_4125);
or U5039 (N_5039,N_4232,N_3980);
nor U5040 (N_5040,N_4495,N_4366);
nand U5041 (N_5041,N_4205,N_3927);
nor U5042 (N_5042,N_4027,N_4070);
nor U5043 (N_5043,N_4011,N_4343);
or U5044 (N_5044,N_4441,N_3761);
nor U5045 (N_5045,N_4006,N_4331);
nor U5046 (N_5046,N_4228,N_3944);
nand U5047 (N_5047,N_4003,N_4370);
nand U5048 (N_5048,N_4016,N_3866);
xor U5049 (N_5049,N_4125,N_4073);
and U5050 (N_5050,N_4323,N_3974);
nand U5051 (N_5051,N_4100,N_4259);
and U5052 (N_5052,N_4354,N_3905);
and U5053 (N_5053,N_4341,N_3992);
nand U5054 (N_5054,N_3762,N_3818);
and U5055 (N_5055,N_4463,N_4044);
or U5056 (N_5056,N_3977,N_4359);
or U5057 (N_5057,N_4376,N_3910);
nand U5058 (N_5058,N_4495,N_3857);
nand U5059 (N_5059,N_4191,N_4210);
nor U5060 (N_5060,N_4349,N_4300);
and U5061 (N_5061,N_4012,N_3963);
or U5062 (N_5062,N_4342,N_3875);
nor U5063 (N_5063,N_4414,N_4181);
nor U5064 (N_5064,N_4106,N_3757);
nand U5065 (N_5065,N_4012,N_3868);
or U5066 (N_5066,N_4455,N_4070);
nand U5067 (N_5067,N_4037,N_3795);
nor U5068 (N_5068,N_4150,N_3866);
nor U5069 (N_5069,N_4317,N_4223);
and U5070 (N_5070,N_4123,N_4434);
nand U5071 (N_5071,N_3980,N_3856);
or U5072 (N_5072,N_3899,N_4138);
or U5073 (N_5073,N_4047,N_3784);
nor U5074 (N_5074,N_4412,N_4472);
or U5075 (N_5075,N_3912,N_3822);
and U5076 (N_5076,N_4165,N_4259);
or U5077 (N_5077,N_4326,N_4436);
and U5078 (N_5078,N_4445,N_4122);
and U5079 (N_5079,N_4229,N_4032);
or U5080 (N_5080,N_4090,N_4492);
and U5081 (N_5081,N_3871,N_4374);
nand U5082 (N_5082,N_4363,N_3889);
and U5083 (N_5083,N_4462,N_4060);
nand U5084 (N_5084,N_4445,N_3947);
nor U5085 (N_5085,N_4119,N_4449);
nor U5086 (N_5086,N_3953,N_3937);
and U5087 (N_5087,N_4292,N_4390);
nor U5088 (N_5088,N_4212,N_3778);
and U5089 (N_5089,N_4293,N_3815);
nand U5090 (N_5090,N_4405,N_3917);
nand U5091 (N_5091,N_4020,N_4290);
nand U5092 (N_5092,N_4439,N_3965);
or U5093 (N_5093,N_4364,N_4180);
and U5094 (N_5094,N_3980,N_4149);
nand U5095 (N_5095,N_4475,N_4302);
nor U5096 (N_5096,N_3819,N_4086);
nand U5097 (N_5097,N_3827,N_4490);
and U5098 (N_5098,N_4038,N_4466);
nand U5099 (N_5099,N_3976,N_4248);
nor U5100 (N_5100,N_3752,N_4142);
and U5101 (N_5101,N_4146,N_4428);
or U5102 (N_5102,N_4457,N_4024);
and U5103 (N_5103,N_4330,N_3781);
and U5104 (N_5104,N_4248,N_4087);
and U5105 (N_5105,N_3781,N_4031);
nand U5106 (N_5106,N_4197,N_3991);
and U5107 (N_5107,N_4238,N_4125);
or U5108 (N_5108,N_3814,N_4090);
and U5109 (N_5109,N_4350,N_4016);
or U5110 (N_5110,N_4062,N_3957);
and U5111 (N_5111,N_4201,N_3996);
or U5112 (N_5112,N_4287,N_4349);
and U5113 (N_5113,N_3816,N_4293);
nand U5114 (N_5114,N_4069,N_4273);
or U5115 (N_5115,N_4183,N_3761);
or U5116 (N_5116,N_4054,N_4415);
nand U5117 (N_5117,N_4397,N_3796);
nand U5118 (N_5118,N_3807,N_4121);
nor U5119 (N_5119,N_4218,N_4389);
and U5120 (N_5120,N_4482,N_4269);
nand U5121 (N_5121,N_3854,N_3961);
or U5122 (N_5122,N_4321,N_4315);
nand U5123 (N_5123,N_3957,N_3882);
or U5124 (N_5124,N_4197,N_4404);
and U5125 (N_5125,N_4117,N_3791);
nand U5126 (N_5126,N_3885,N_4403);
and U5127 (N_5127,N_4126,N_3902);
or U5128 (N_5128,N_3774,N_3835);
or U5129 (N_5129,N_3842,N_4492);
nor U5130 (N_5130,N_3775,N_3801);
or U5131 (N_5131,N_4314,N_3979);
nor U5132 (N_5132,N_3939,N_3969);
nor U5133 (N_5133,N_4424,N_4175);
nand U5134 (N_5134,N_4010,N_4475);
and U5135 (N_5135,N_4300,N_4322);
nor U5136 (N_5136,N_4350,N_3782);
nand U5137 (N_5137,N_4440,N_4326);
and U5138 (N_5138,N_3927,N_4376);
nor U5139 (N_5139,N_3868,N_3986);
nor U5140 (N_5140,N_4108,N_4457);
nor U5141 (N_5141,N_4025,N_3877);
nand U5142 (N_5142,N_4461,N_3978);
or U5143 (N_5143,N_4055,N_3965);
nor U5144 (N_5144,N_3986,N_4051);
nand U5145 (N_5145,N_4068,N_3754);
and U5146 (N_5146,N_3878,N_4498);
nor U5147 (N_5147,N_4362,N_3984);
nor U5148 (N_5148,N_3769,N_3985);
and U5149 (N_5149,N_3931,N_4330);
nor U5150 (N_5150,N_4365,N_3977);
or U5151 (N_5151,N_4337,N_4289);
nor U5152 (N_5152,N_4068,N_4023);
nand U5153 (N_5153,N_4221,N_4003);
or U5154 (N_5154,N_3961,N_4326);
and U5155 (N_5155,N_4024,N_3938);
nor U5156 (N_5156,N_4460,N_4126);
and U5157 (N_5157,N_4348,N_4182);
xor U5158 (N_5158,N_4260,N_4297);
nor U5159 (N_5159,N_3962,N_4491);
and U5160 (N_5160,N_3868,N_3859);
and U5161 (N_5161,N_3767,N_4434);
or U5162 (N_5162,N_4275,N_3975);
or U5163 (N_5163,N_4350,N_3916);
nor U5164 (N_5164,N_3939,N_3895);
nor U5165 (N_5165,N_4438,N_4314);
and U5166 (N_5166,N_3857,N_3918);
or U5167 (N_5167,N_4229,N_4154);
nor U5168 (N_5168,N_3901,N_3854);
or U5169 (N_5169,N_4358,N_4249);
nor U5170 (N_5170,N_4228,N_4139);
nor U5171 (N_5171,N_4465,N_4175);
or U5172 (N_5172,N_4106,N_4447);
nor U5173 (N_5173,N_4009,N_3918);
xnor U5174 (N_5174,N_3845,N_4097);
or U5175 (N_5175,N_3919,N_3947);
nand U5176 (N_5176,N_4166,N_3855);
nand U5177 (N_5177,N_4101,N_4324);
nor U5178 (N_5178,N_4082,N_3802);
nand U5179 (N_5179,N_4463,N_4180);
nand U5180 (N_5180,N_4047,N_4318);
or U5181 (N_5181,N_4383,N_4187);
nor U5182 (N_5182,N_4464,N_4472);
nand U5183 (N_5183,N_3883,N_4064);
nor U5184 (N_5184,N_4052,N_4086);
or U5185 (N_5185,N_4248,N_4320);
nor U5186 (N_5186,N_4289,N_4255);
nand U5187 (N_5187,N_4384,N_4093);
nor U5188 (N_5188,N_4159,N_4392);
or U5189 (N_5189,N_4277,N_4431);
or U5190 (N_5190,N_4073,N_3948);
or U5191 (N_5191,N_4478,N_3865);
or U5192 (N_5192,N_4209,N_4421);
xnor U5193 (N_5193,N_4016,N_3850);
and U5194 (N_5194,N_4245,N_4074);
or U5195 (N_5195,N_4451,N_3916);
or U5196 (N_5196,N_4087,N_4368);
and U5197 (N_5197,N_4290,N_4460);
or U5198 (N_5198,N_4339,N_4205);
or U5199 (N_5199,N_4455,N_4005);
and U5200 (N_5200,N_4035,N_3865);
or U5201 (N_5201,N_4491,N_4057);
or U5202 (N_5202,N_4130,N_4195);
and U5203 (N_5203,N_3753,N_4349);
or U5204 (N_5204,N_4189,N_4219);
nand U5205 (N_5205,N_3993,N_4414);
and U5206 (N_5206,N_4216,N_4071);
and U5207 (N_5207,N_3979,N_4186);
nor U5208 (N_5208,N_4099,N_4194);
nor U5209 (N_5209,N_4340,N_4141);
and U5210 (N_5210,N_4433,N_4432);
nor U5211 (N_5211,N_4294,N_4167);
or U5212 (N_5212,N_3993,N_4497);
or U5213 (N_5213,N_3799,N_4136);
or U5214 (N_5214,N_4394,N_4157);
or U5215 (N_5215,N_4157,N_4201);
nor U5216 (N_5216,N_4068,N_4495);
nand U5217 (N_5217,N_3922,N_4210);
nor U5218 (N_5218,N_4319,N_4287);
and U5219 (N_5219,N_3847,N_3785);
nor U5220 (N_5220,N_4425,N_3998);
and U5221 (N_5221,N_3887,N_4159);
or U5222 (N_5222,N_4048,N_3803);
nor U5223 (N_5223,N_4483,N_3941);
nand U5224 (N_5224,N_4048,N_4439);
nand U5225 (N_5225,N_4255,N_4356);
or U5226 (N_5226,N_4307,N_4120);
nor U5227 (N_5227,N_4387,N_4117);
or U5228 (N_5228,N_4332,N_4249);
or U5229 (N_5229,N_4456,N_4156);
or U5230 (N_5230,N_4404,N_3787);
nor U5231 (N_5231,N_4301,N_4035);
nand U5232 (N_5232,N_4378,N_4401);
or U5233 (N_5233,N_3857,N_4120);
nand U5234 (N_5234,N_3818,N_4341);
and U5235 (N_5235,N_3826,N_4241);
and U5236 (N_5236,N_4021,N_4390);
and U5237 (N_5237,N_4360,N_3999);
or U5238 (N_5238,N_3992,N_4097);
nand U5239 (N_5239,N_4424,N_4178);
and U5240 (N_5240,N_4406,N_3928);
nor U5241 (N_5241,N_3778,N_4463);
and U5242 (N_5242,N_4232,N_3997);
and U5243 (N_5243,N_3917,N_3752);
or U5244 (N_5244,N_3755,N_4488);
nor U5245 (N_5245,N_4332,N_4031);
or U5246 (N_5246,N_4114,N_3873);
nand U5247 (N_5247,N_4043,N_4431);
nand U5248 (N_5248,N_3929,N_3770);
and U5249 (N_5249,N_4356,N_3829);
and U5250 (N_5250,N_5203,N_5021);
nand U5251 (N_5251,N_5166,N_4740);
and U5252 (N_5252,N_4706,N_5053);
nor U5253 (N_5253,N_4925,N_5022);
or U5254 (N_5254,N_4796,N_4799);
and U5255 (N_5255,N_4910,N_5196);
nor U5256 (N_5256,N_5028,N_4697);
and U5257 (N_5257,N_5120,N_5115);
nor U5258 (N_5258,N_4755,N_5145);
or U5259 (N_5259,N_5118,N_4847);
and U5260 (N_5260,N_4524,N_4867);
nand U5261 (N_5261,N_4620,N_4977);
nand U5262 (N_5262,N_5225,N_4574);
and U5263 (N_5263,N_4961,N_4729);
and U5264 (N_5264,N_4721,N_5163);
nand U5265 (N_5265,N_4969,N_4835);
and U5266 (N_5266,N_4992,N_4905);
nor U5267 (N_5267,N_4749,N_5039);
nor U5268 (N_5268,N_5098,N_4887);
nand U5269 (N_5269,N_5151,N_5026);
or U5270 (N_5270,N_4991,N_4713);
and U5271 (N_5271,N_4743,N_4908);
nor U5272 (N_5272,N_4576,N_4568);
nor U5273 (N_5273,N_4757,N_4629);
and U5274 (N_5274,N_5070,N_5065);
and U5275 (N_5275,N_4946,N_5023);
nand U5276 (N_5276,N_4562,N_4644);
nand U5277 (N_5277,N_5057,N_5068);
or U5278 (N_5278,N_5035,N_4958);
nand U5279 (N_5279,N_4546,N_5034);
and U5280 (N_5280,N_4826,N_4722);
and U5281 (N_5281,N_4979,N_4781);
and U5282 (N_5282,N_5008,N_4968);
and U5283 (N_5283,N_5036,N_4636);
or U5284 (N_5284,N_5169,N_5159);
nand U5285 (N_5285,N_4681,N_4702);
nor U5286 (N_5286,N_4542,N_5173);
or U5287 (N_5287,N_4658,N_4807);
or U5288 (N_5288,N_5227,N_5217);
and U5289 (N_5289,N_5032,N_4824);
nand U5290 (N_5290,N_5071,N_4857);
xnor U5291 (N_5291,N_4858,N_4565);
nor U5292 (N_5292,N_4689,N_4733);
and U5293 (N_5293,N_4864,N_5238);
or U5294 (N_5294,N_4639,N_5056);
nor U5295 (N_5295,N_4547,N_4793);
and U5296 (N_5296,N_5042,N_4525);
and U5297 (N_5297,N_5067,N_4573);
nand U5298 (N_5298,N_4596,N_4570);
nand U5299 (N_5299,N_5155,N_5054);
or U5300 (N_5300,N_4594,N_5123);
xnor U5301 (N_5301,N_5104,N_4580);
nand U5302 (N_5302,N_5073,N_4764);
or U5303 (N_5303,N_4677,N_4708);
and U5304 (N_5304,N_4940,N_5185);
and U5305 (N_5305,N_5037,N_4543);
and U5306 (N_5306,N_5174,N_4919);
nand U5307 (N_5307,N_5214,N_4974);
and U5308 (N_5308,N_4667,N_5184);
nand U5309 (N_5309,N_4859,N_4759);
nand U5310 (N_5310,N_5016,N_4656);
nor U5311 (N_5311,N_4723,N_4627);
nor U5312 (N_5312,N_4558,N_4704);
and U5313 (N_5313,N_5153,N_4825);
nand U5314 (N_5314,N_4760,N_5136);
and U5315 (N_5315,N_4665,N_5130);
or U5316 (N_5316,N_4701,N_5033);
or U5317 (N_5317,N_4834,N_4775);
nand U5318 (N_5318,N_5210,N_4561);
or U5319 (N_5319,N_4690,N_4985);
nand U5320 (N_5320,N_4604,N_5051);
and U5321 (N_5321,N_4548,N_4720);
nand U5322 (N_5322,N_4763,N_5085);
and U5323 (N_5323,N_4805,N_4739);
nor U5324 (N_5324,N_5103,N_4592);
nand U5325 (N_5325,N_4886,N_4553);
and U5326 (N_5326,N_5055,N_4651);
or U5327 (N_5327,N_5087,N_4661);
and U5328 (N_5328,N_5079,N_5062);
or U5329 (N_5329,N_5193,N_4909);
nand U5330 (N_5330,N_4680,N_5011);
nand U5331 (N_5331,N_4798,N_5030);
or U5332 (N_5332,N_5243,N_4841);
nand U5333 (N_5333,N_4560,N_5232);
and U5334 (N_5334,N_5077,N_4972);
or U5335 (N_5335,N_4773,N_4995);
nor U5336 (N_5336,N_4581,N_4672);
and U5337 (N_5337,N_5190,N_4539);
and U5338 (N_5338,N_5179,N_4534);
or U5339 (N_5339,N_4682,N_5014);
nor U5340 (N_5340,N_4942,N_4555);
and U5341 (N_5341,N_4559,N_4950);
or U5342 (N_5342,N_5106,N_5082);
or U5343 (N_5343,N_4692,N_5048);
nor U5344 (N_5344,N_4820,N_4663);
nor U5345 (N_5345,N_4506,N_4753);
and U5346 (N_5346,N_5158,N_5201);
and U5347 (N_5347,N_4741,N_5245);
or U5348 (N_5348,N_4552,N_4920);
nand U5349 (N_5349,N_4626,N_4586);
or U5350 (N_5350,N_4612,N_5182);
nor U5351 (N_5351,N_4994,N_4971);
nor U5352 (N_5352,N_4997,N_4650);
nand U5353 (N_5353,N_5189,N_4711);
nand U5354 (N_5354,N_4698,N_4838);
nand U5355 (N_5355,N_4808,N_4615);
or U5356 (N_5356,N_5249,N_4556);
or U5357 (N_5357,N_5050,N_4707);
or U5358 (N_5358,N_4877,N_4715);
nand U5359 (N_5359,N_4765,N_4806);
or U5360 (N_5360,N_4873,N_4662);
or U5361 (N_5361,N_4771,N_5088);
nor U5362 (N_5362,N_4640,N_4926);
or U5363 (N_5363,N_4609,N_4976);
nand U5364 (N_5364,N_4549,N_4705);
or U5365 (N_5365,N_5094,N_5195);
and U5366 (N_5366,N_4571,N_5031);
nand U5367 (N_5367,N_5220,N_5059);
nand U5368 (N_5368,N_4579,N_4980);
nor U5369 (N_5369,N_4645,N_4693);
nor U5370 (N_5370,N_5187,N_4792);
nand U5371 (N_5371,N_4724,N_4929);
and U5372 (N_5372,N_4931,N_4914);
and U5373 (N_5373,N_5170,N_5208);
nand U5374 (N_5374,N_5224,N_4800);
and U5375 (N_5375,N_4769,N_5063);
nor U5376 (N_5376,N_4747,N_4633);
nor U5377 (N_5377,N_4881,N_4975);
nor U5378 (N_5378,N_4522,N_5186);
or U5379 (N_5379,N_4566,N_4554);
nand U5380 (N_5380,N_4801,N_5108);
or U5381 (N_5381,N_4718,N_4589);
and U5382 (N_5382,N_4660,N_4927);
or U5383 (N_5383,N_4903,N_4699);
nand U5384 (N_5384,N_5006,N_4694);
nor U5385 (N_5385,N_5119,N_4528);
and U5386 (N_5386,N_4954,N_5141);
and U5387 (N_5387,N_4578,N_5235);
nor U5388 (N_5388,N_5047,N_4804);
nor U5389 (N_5389,N_4537,N_4659);
nand U5390 (N_5390,N_5191,N_4517);
nand U5391 (N_5391,N_5194,N_4738);
nor U5392 (N_5392,N_4965,N_4744);
or U5393 (N_5393,N_4735,N_4829);
nand U5394 (N_5394,N_4737,N_5049);
nand U5395 (N_5395,N_5024,N_4736);
nand U5396 (N_5396,N_4840,N_4944);
and U5397 (N_5397,N_4683,N_4649);
and U5398 (N_5398,N_4898,N_4582);
or U5399 (N_5399,N_5124,N_4803);
nor U5400 (N_5400,N_4618,N_5212);
and U5401 (N_5401,N_5211,N_4684);
nand U5402 (N_5402,N_4595,N_4790);
and U5403 (N_5403,N_4606,N_4779);
nor U5404 (N_5404,N_5043,N_4623);
and U5405 (N_5405,N_5218,N_4508);
nand U5406 (N_5406,N_5020,N_5083);
nor U5407 (N_5407,N_4754,N_4782);
and U5408 (N_5408,N_4959,N_5114);
nand U5409 (N_5409,N_4628,N_4583);
nand U5410 (N_5410,N_4676,N_4742);
nor U5411 (N_5411,N_5164,N_4577);
nor U5412 (N_5412,N_4678,N_5204);
and U5413 (N_5413,N_4936,N_5197);
and U5414 (N_5414,N_4734,N_4605);
or U5415 (N_5415,N_4885,N_5125);
and U5416 (N_5416,N_5058,N_4732);
nand U5417 (N_5417,N_4511,N_4837);
or U5418 (N_5418,N_4527,N_4990);
nor U5419 (N_5419,N_4933,N_4624);
or U5420 (N_5420,N_4671,N_4756);
nor U5421 (N_5421,N_5157,N_4564);
or U5422 (N_5422,N_5112,N_5084);
nor U5423 (N_5423,N_5215,N_4584);
nor U5424 (N_5424,N_4501,N_4674);
and U5425 (N_5425,N_5241,N_4998);
or U5426 (N_5426,N_4865,N_5010);
and U5427 (N_5427,N_4861,N_5132);
and U5428 (N_5428,N_5202,N_4719);
and U5429 (N_5429,N_5207,N_4685);
and U5430 (N_5430,N_4823,N_4850);
and U5431 (N_5431,N_4730,N_4917);
nor U5432 (N_5432,N_5140,N_4949);
nand U5433 (N_5433,N_4621,N_5167);
nor U5434 (N_5434,N_4780,N_4745);
nand U5435 (N_5435,N_4852,N_5005);
nand U5436 (N_5436,N_5236,N_5240);
or U5437 (N_5437,N_4853,N_5052);
and U5438 (N_5438,N_4844,N_4669);
nor U5439 (N_5439,N_5229,N_4540);
and U5440 (N_5440,N_4777,N_4938);
and U5441 (N_5441,N_4599,N_5025);
nor U5442 (N_5442,N_4726,N_4842);
or U5443 (N_5443,N_4591,N_4934);
or U5444 (N_5444,N_4657,N_4695);
and U5445 (N_5445,N_4696,N_5038);
nor U5446 (N_5446,N_4987,N_5116);
nand U5447 (N_5447,N_5007,N_4758);
or U5448 (N_5448,N_4863,N_4809);
nor U5449 (N_5449,N_5209,N_4673);
or U5450 (N_5450,N_5081,N_4544);
nor U5451 (N_5451,N_4831,N_4523);
and U5452 (N_5452,N_5149,N_5213);
nand U5453 (N_5453,N_4794,N_4916);
nand U5454 (N_5454,N_4631,N_4608);
or U5455 (N_5455,N_4545,N_5064);
and U5456 (N_5456,N_5000,N_4960);
or U5457 (N_5457,N_4514,N_4891);
and U5458 (N_5458,N_5075,N_4637);
and U5459 (N_5459,N_5178,N_4846);
nand U5460 (N_5460,N_4984,N_4770);
and U5461 (N_5461,N_4569,N_5183);
or U5462 (N_5462,N_4830,N_4789);
nor U5463 (N_5463,N_5113,N_5198);
nor U5464 (N_5464,N_4983,N_4664);
and U5465 (N_5465,N_4797,N_4911);
nor U5466 (N_5466,N_4817,N_4996);
and U5467 (N_5467,N_4928,N_4956);
and U5468 (N_5468,N_5095,N_4783);
nor U5469 (N_5469,N_5107,N_4748);
and U5470 (N_5470,N_4646,N_4868);
or U5471 (N_5471,N_5041,N_5076);
or U5472 (N_5472,N_4505,N_5154);
or U5473 (N_5473,N_4879,N_5066);
nand U5474 (N_5474,N_5101,N_5069);
and U5475 (N_5475,N_4727,N_4828);
or U5476 (N_5476,N_4647,N_4746);
or U5477 (N_5477,N_4939,N_5138);
xor U5478 (N_5478,N_5003,N_4654);
nor U5479 (N_5479,N_4810,N_5102);
nand U5480 (N_5480,N_5040,N_5248);
and U5481 (N_5481,N_4526,N_4848);
and U5482 (N_5482,N_4688,N_4894);
and U5483 (N_5483,N_5131,N_4989);
and U5484 (N_5484,N_4507,N_5097);
nand U5485 (N_5485,N_5181,N_5015);
or U5486 (N_5486,N_5216,N_5091);
or U5487 (N_5487,N_5129,N_4888);
nor U5488 (N_5488,N_4981,N_4752);
or U5489 (N_5489,N_4768,N_4811);
and U5490 (N_5490,N_5176,N_5002);
and U5491 (N_5491,N_5009,N_5223);
nor U5492 (N_5492,N_4814,N_4890);
and U5493 (N_5493,N_5247,N_4788);
or U5494 (N_5494,N_4536,N_4832);
and U5495 (N_5495,N_4851,N_4686);
and U5496 (N_5496,N_4725,N_5146);
or U5497 (N_5497,N_4778,N_4625);
nor U5498 (N_5498,N_4786,N_4611);
nor U5499 (N_5499,N_4967,N_5027);
nand U5500 (N_5500,N_4907,N_4535);
and U5501 (N_5501,N_4839,N_4833);
and U5502 (N_5502,N_5019,N_5122);
nand U5503 (N_5503,N_4630,N_4856);
and U5504 (N_5504,N_4533,N_4632);
or U5505 (N_5505,N_4516,N_4973);
or U5506 (N_5506,N_4901,N_4716);
nor U5507 (N_5507,N_4550,N_4935);
and U5508 (N_5508,N_5099,N_4666);
or U5509 (N_5509,N_4870,N_4978);
and U5510 (N_5510,N_4691,N_4787);
nor U5511 (N_5511,N_5156,N_5222);
nor U5512 (N_5512,N_5221,N_4915);
and U5513 (N_5513,N_4590,N_5078);
or U5514 (N_5514,N_5239,N_4945);
nand U5515 (N_5515,N_5089,N_4648);
or U5516 (N_5516,N_4812,N_4731);
and U5517 (N_5517,N_4538,N_4947);
or U5518 (N_5518,N_4795,N_4670);
nand U5519 (N_5519,N_4512,N_4986);
nand U5520 (N_5520,N_4613,N_4948);
nor U5521 (N_5521,N_4588,N_5188);
and U5522 (N_5522,N_5139,N_4703);
and U5523 (N_5523,N_4531,N_4937);
nand U5524 (N_5524,N_4597,N_4880);
nand U5525 (N_5525,N_4515,N_5096);
or U5526 (N_5526,N_5162,N_4668);
nor U5527 (N_5527,N_4572,N_5160);
nor U5528 (N_5528,N_4862,N_4896);
nor U5529 (N_5529,N_4962,N_4988);
or U5530 (N_5530,N_4563,N_5012);
and U5531 (N_5531,N_4966,N_4772);
and U5532 (N_5532,N_4712,N_4871);
nand U5533 (N_5533,N_4529,N_4906);
or U5534 (N_5534,N_5171,N_5109);
or U5535 (N_5535,N_4893,N_4784);
nand U5536 (N_5536,N_4643,N_4816);
nand U5537 (N_5537,N_5144,N_4884);
nand U5538 (N_5538,N_5135,N_5080);
nor U5539 (N_5539,N_4855,N_4912);
nand U5540 (N_5540,N_5142,N_4819);
nor U5541 (N_5541,N_4895,N_4614);
nor U5542 (N_5542,N_4504,N_4774);
or U5543 (N_5543,N_4617,N_4675);
and U5544 (N_5544,N_4575,N_5100);
nor U5545 (N_5545,N_4883,N_4761);
nand U5546 (N_5546,N_4902,N_4642);
and U5547 (N_5547,N_5105,N_4509);
or U5548 (N_5548,N_4921,N_4875);
nor U5549 (N_5549,N_4941,N_4622);
and U5550 (N_5550,N_4776,N_4913);
nand U5551 (N_5551,N_4952,N_4963);
or U5552 (N_5552,N_4500,N_4930);
and U5553 (N_5553,N_4869,N_4943);
and U5554 (N_5554,N_4641,N_5205);
and U5555 (N_5555,N_4872,N_4815);
or U5556 (N_5556,N_4530,N_4503);
and U5557 (N_5557,N_5233,N_5092);
nor U5558 (N_5558,N_5126,N_4766);
nand U5559 (N_5559,N_5230,N_5228);
and U5560 (N_5560,N_4714,N_5086);
and U5561 (N_5561,N_5093,N_4892);
and U5562 (N_5562,N_5044,N_4951);
and U5563 (N_5563,N_4785,N_4845);
or U5564 (N_5564,N_5150,N_5137);
nor U5565 (N_5565,N_5180,N_5234);
nor U5566 (N_5566,N_4587,N_4932);
or U5567 (N_5567,N_4541,N_5127);
nand U5568 (N_5568,N_5206,N_4821);
and U5569 (N_5569,N_5165,N_4638);
nand U5570 (N_5570,N_4924,N_5117);
and U5571 (N_5571,N_4882,N_4557);
and U5572 (N_5572,N_4982,N_5237);
nor U5573 (N_5573,N_4818,N_4900);
or U5574 (N_5574,N_5200,N_5017);
nand U5575 (N_5575,N_5143,N_5244);
or U5576 (N_5576,N_4843,N_4717);
and U5577 (N_5577,N_4849,N_4953);
nand U5578 (N_5578,N_5147,N_5192);
or U5579 (N_5579,N_5172,N_4600);
or U5580 (N_5580,N_4874,N_5152);
or U5581 (N_5581,N_5060,N_5074);
nor U5582 (N_5582,N_4518,N_4700);
nor U5583 (N_5583,N_4679,N_5133);
and U5584 (N_5584,N_5161,N_4889);
nand U5585 (N_5585,N_5148,N_4634);
and U5586 (N_5586,N_4866,N_4635);
and U5587 (N_5587,N_4899,N_5231);
nor U5588 (N_5588,N_4602,N_5134);
nand U5589 (N_5589,N_5199,N_4918);
or U5590 (N_5590,N_4653,N_4762);
nor U5591 (N_5591,N_5013,N_4616);
nor U5592 (N_5592,N_4878,N_4619);
and U5593 (N_5593,N_5175,N_4593);
nand U5594 (N_5594,N_5177,N_4510);
nor U5595 (N_5595,N_4610,N_5111);
or U5596 (N_5596,N_5029,N_4750);
nand U5597 (N_5597,N_4802,N_4860);
nor U5598 (N_5598,N_4652,N_4827);
or U5599 (N_5599,N_4585,N_4607);
or U5600 (N_5600,N_4813,N_4767);
nor U5601 (N_5601,N_5045,N_4603);
nand U5602 (N_5602,N_4791,N_5246);
and U5603 (N_5603,N_4993,N_4521);
nand U5604 (N_5604,N_5061,N_5001);
or U5605 (N_5605,N_4520,N_4687);
and U5606 (N_5606,N_5168,N_4751);
and U5607 (N_5607,N_4822,N_5046);
or U5608 (N_5608,N_4904,N_4709);
or U5609 (N_5609,N_4999,N_4957);
and U5610 (N_5610,N_5128,N_5121);
or U5611 (N_5611,N_5004,N_4922);
or U5612 (N_5612,N_4551,N_4655);
and U5613 (N_5613,N_5072,N_5090);
or U5614 (N_5614,N_4964,N_4876);
nor U5615 (N_5615,N_4502,N_4710);
nand U5616 (N_5616,N_5226,N_5018);
nand U5617 (N_5617,N_5242,N_4567);
nor U5618 (N_5618,N_4923,N_4532);
and U5619 (N_5619,N_4955,N_4598);
and U5620 (N_5620,N_5110,N_4519);
nor U5621 (N_5621,N_4836,N_4728);
nor U5622 (N_5622,N_5219,N_4970);
nand U5623 (N_5623,N_4854,N_4601);
nand U5624 (N_5624,N_4897,N_4513);
or U5625 (N_5625,N_5040,N_4775);
and U5626 (N_5626,N_5129,N_5222);
nand U5627 (N_5627,N_5084,N_4804);
nand U5628 (N_5628,N_5044,N_4609);
nand U5629 (N_5629,N_4996,N_5083);
and U5630 (N_5630,N_5102,N_4948);
nor U5631 (N_5631,N_4636,N_4971);
and U5632 (N_5632,N_4988,N_4895);
nand U5633 (N_5633,N_4938,N_4929);
nand U5634 (N_5634,N_4536,N_4863);
nor U5635 (N_5635,N_4614,N_4798);
or U5636 (N_5636,N_4520,N_4934);
and U5637 (N_5637,N_4910,N_4962);
and U5638 (N_5638,N_4552,N_4659);
nor U5639 (N_5639,N_4546,N_5053);
and U5640 (N_5640,N_5025,N_5174);
nand U5641 (N_5641,N_4813,N_5143);
and U5642 (N_5642,N_4605,N_5157);
and U5643 (N_5643,N_4842,N_4869);
nand U5644 (N_5644,N_5184,N_4563);
nor U5645 (N_5645,N_4713,N_4986);
nand U5646 (N_5646,N_4764,N_4866);
or U5647 (N_5647,N_5077,N_5173);
and U5648 (N_5648,N_4634,N_4888);
nand U5649 (N_5649,N_4768,N_4889);
nor U5650 (N_5650,N_5118,N_4758);
or U5651 (N_5651,N_4641,N_5011);
nand U5652 (N_5652,N_5165,N_4767);
nand U5653 (N_5653,N_4863,N_4600);
or U5654 (N_5654,N_4902,N_5152);
and U5655 (N_5655,N_4541,N_5243);
and U5656 (N_5656,N_5129,N_4504);
and U5657 (N_5657,N_4575,N_4726);
and U5658 (N_5658,N_5248,N_4712);
nand U5659 (N_5659,N_4730,N_4791);
and U5660 (N_5660,N_5137,N_4714);
nor U5661 (N_5661,N_4833,N_5171);
and U5662 (N_5662,N_5107,N_4536);
nor U5663 (N_5663,N_4887,N_4557);
nor U5664 (N_5664,N_4876,N_4594);
or U5665 (N_5665,N_4764,N_4742);
or U5666 (N_5666,N_5176,N_4631);
or U5667 (N_5667,N_5233,N_5164);
xnor U5668 (N_5668,N_4995,N_5234);
and U5669 (N_5669,N_5189,N_5020);
and U5670 (N_5670,N_4750,N_5211);
xor U5671 (N_5671,N_5098,N_4740);
nand U5672 (N_5672,N_4946,N_4872);
nand U5673 (N_5673,N_4902,N_4596);
nand U5674 (N_5674,N_4526,N_5085);
and U5675 (N_5675,N_4961,N_4894);
and U5676 (N_5676,N_4685,N_5114);
nand U5677 (N_5677,N_4883,N_5107);
nand U5678 (N_5678,N_4615,N_4580);
nor U5679 (N_5679,N_4724,N_4910);
nor U5680 (N_5680,N_4721,N_4741);
and U5681 (N_5681,N_5001,N_4609);
or U5682 (N_5682,N_5010,N_5112);
xnor U5683 (N_5683,N_5184,N_5105);
nand U5684 (N_5684,N_4629,N_5020);
nor U5685 (N_5685,N_4747,N_5030);
and U5686 (N_5686,N_4646,N_4522);
nand U5687 (N_5687,N_4974,N_4568);
nor U5688 (N_5688,N_4555,N_4977);
or U5689 (N_5689,N_4642,N_4851);
nand U5690 (N_5690,N_5085,N_5136);
nor U5691 (N_5691,N_5035,N_5029);
nand U5692 (N_5692,N_4855,N_4789);
and U5693 (N_5693,N_5082,N_4759);
nand U5694 (N_5694,N_4583,N_5099);
or U5695 (N_5695,N_5115,N_5118);
nand U5696 (N_5696,N_4695,N_4914);
and U5697 (N_5697,N_4849,N_4706);
and U5698 (N_5698,N_4974,N_4875);
and U5699 (N_5699,N_5016,N_4789);
and U5700 (N_5700,N_4951,N_4539);
and U5701 (N_5701,N_5181,N_5065);
nor U5702 (N_5702,N_4687,N_5008);
or U5703 (N_5703,N_5140,N_4713);
or U5704 (N_5704,N_5233,N_4688);
nand U5705 (N_5705,N_5235,N_5080);
and U5706 (N_5706,N_4546,N_5064);
or U5707 (N_5707,N_5228,N_5128);
and U5708 (N_5708,N_5163,N_5116);
nor U5709 (N_5709,N_5102,N_5016);
nor U5710 (N_5710,N_4687,N_4854);
and U5711 (N_5711,N_5084,N_4515);
nand U5712 (N_5712,N_4964,N_5195);
or U5713 (N_5713,N_4625,N_4510);
nand U5714 (N_5714,N_5103,N_4807);
or U5715 (N_5715,N_5108,N_5248);
or U5716 (N_5716,N_4710,N_4545);
nand U5717 (N_5717,N_4604,N_5139);
and U5718 (N_5718,N_5065,N_5045);
or U5719 (N_5719,N_5223,N_5169);
or U5720 (N_5720,N_4615,N_4600);
and U5721 (N_5721,N_4512,N_5071);
and U5722 (N_5722,N_5086,N_5212);
nor U5723 (N_5723,N_5073,N_4596);
and U5724 (N_5724,N_4962,N_4980);
nand U5725 (N_5725,N_4930,N_4553);
and U5726 (N_5726,N_4528,N_4984);
nor U5727 (N_5727,N_4532,N_5037);
nand U5728 (N_5728,N_5181,N_4612);
nand U5729 (N_5729,N_4895,N_4616);
and U5730 (N_5730,N_4518,N_5124);
or U5731 (N_5731,N_4602,N_4996);
nand U5732 (N_5732,N_5089,N_5206);
or U5733 (N_5733,N_4916,N_4672);
and U5734 (N_5734,N_4926,N_4548);
or U5735 (N_5735,N_4681,N_4829);
or U5736 (N_5736,N_5149,N_5159);
nand U5737 (N_5737,N_4648,N_4546);
and U5738 (N_5738,N_4682,N_4611);
and U5739 (N_5739,N_4643,N_4756);
and U5740 (N_5740,N_4945,N_5209);
nand U5741 (N_5741,N_5107,N_4691);
nor U5742 (N_5742,N_4975,N_4992);
or U5743 (N_5743,N_4915,N_5157);
nand U5744 (N_5744,N_4708,N_5128);
or U5745 (N_5745,N_4966,N_4965);
nand U5746 (N_5746,N_5086,N_5104);
and U5747 (N_5747,N_4964,N_4505);
nand U5748 (N_5748,N_5242,N_4694);
nor U5749 (N_5749,N_5070,N_5082);
nand U5750 (N_5750,N_4690,N_4617);
and U5751 (N_5751,N_5093,N_5092);
and U5752 (N_5752,N_4837,N_4826);
nor U5753 (N_5753,N_5219,N_5156);
nand U5754 (N_5754,N_4710,N_4648);
nor U5755 (N_5755,N_4785,N_4550);
nor U5756 (N_5756,N_5183,N_4503);
nor U5757 (N_5757,N_4564,N_4800);
nand U5758 (N_5758,N_4648,N_4834);
and U5759 (N_5759,N_4879,N_5136);
and U5760 (N_5760,N_4680,N_4987);
and U5761 (N_5761,N_4835,N_5245);
and U5762 (N_5762,N_4872,N_4720);
nor U5763 (N_5763,N_4803,N_5115);
nor U5764 (N_5764,N_4728,N_4592);
or U5765 (N_5765,N_4510,N_5156);
nand U5766 (N_5766,N_4641,N_4901);
nand U5767 (N_5767,N_4606,N_4604);
nand U5768 (N_5768,N_5072,N_5162);
or U5769 (N_5769,N_4990,N_4849);
and U5770 (N_5770,N_4721,N_4695);
and U5771 (N_5771,N_4869,N_4890);
and U5772 (N_5772,N_5181,N_5127);
or U5773 (N_5773,N_4747,N_4711);
nand U5774 (N_5774,N_4506,N_4754);
or U5775 (N_5775,N_4743,N_4739);
or U5776 (N_5776,N_4778,N_4631);
and U5777 (N_5777,N_4712,N_5141);
and U5778 (N_5778,N_4970,N_4800);
nand U5779 (N_5779,N_5144,N_5178);
nand U5780 (N_5780,N_5153,N_4979);
nor U5781 (N_5781,N_4837,N_4543);
or U5782 (N_5782,N_5076,N_5132);
nand U5783 (N_5783,N_5211,N_4734);
or U5784 (N_5784,N_5094,N_4578);
or U5785 (N_5785,N_5113,N_4536);
or U5786 (N_5786,N_4540,N_4543);
or U5787 (N_5787,N_4587,N_4641);
nor U5788 (N_5788,N_4674,N_5211);
nor U5789 (N_5789,N_4903,N_4514);
nand U5790 (N_5790,N_4685,N_5084);
or U5791 (N_5791,N_4505,N_5206);
or U5792 (N_5792,N_4901,N_5249);
and U5793 (N_5793,N_4870,N_4584);
nand U5794 (N_5794,N_4789,N_4783);
and U5795 (N_5795,N_5070,N_5157);
nand U5796 (N_5796,N_5064,N_4857);
or U5797 (N_5797,N_5226,N_4865);
or U5798 (N_5798,N_4914,N_4932);
nand U5799 (N_5799,N_5088,N_5083);
nand U5800 (N_5800,N_4517,N_5210);
nand U5801 (N_5801,N_4566,N_5067);
or U5802 (N_5802,N_5127,N_4547);
nand U5803 (N_5803,N_5011,N_5221);
and U5804 (N_5804,N_5074,N_4706);
or U5805 (N_5805,N_4798,N_4671);
or U5806 (N_5806,N_4544,N_5137);
or U5807 (N_5807,N_4851,N_5207);
nand U5808 (N_5808,N_4721,N_4522);
or U5809 (N_5809,N_5024,N_4680);
nand U5810 (N_5810,N_4503,N_5080);
nand U5811 (N_5811,N_4791,N_4982);
and U5812 (N_5812,N_4696,N_5200);
nor U5813 (N_5813,N_5020,N_5237);
and U5814 (N_5814,N_4695,N_4577);
nand U5815 (N_5815,N_4974,N_4853);
nor U5816 (N_5816,N_4650,N_5231);
or U5817 (N_5817,N_5204,N_4561);
nand U5818 (N_5818,N_4838,N_4761);
or U5819 (N_5819,N_4558,N_5232);
and U5820 (N_5820,N_5245,N_4867);
or U5821 (N_5821,N_4989,N_5104);
nand U5822 (N_5822,N_4636,N_5201);
and U5823 (N_5823,N_4899,N_5216);
nor U5824 (N_5824,N_4904,N_5227);
nor U5825 (N_5825,N_5054,N_4753);
or U5826 (N_5826,N_5096,N_5070);
nor U5827 (N_5827,N_5180,N_5160);
and U5828 (N_5828,N_5089,N_4616);
or U5829 (N_5829,N_4625,N_4688);
or U5830 (N_5830,N_5202,N_5179);
nor U5831 (N_5831,N_4694,N_4949);
nor U5832 (N_5832,N_5233,N_4895);
nor U5833 (N_5833,N_5199,N_4798);
and U5834 (N_5834,N_5227,N_5080);
or U5835 (N_5835,N_4867,N_4914);
nand U5836 (N_5836,N_4692,N_5011);
nand U5837 (N_5837,N_4891,N_5128);
or U5838 (N_5838,N_4955,N_4970);
and U5839 (N_5839,N_4862,N_5198);
nand U5840 (N_5840,N_4970,N_4943);
nand U5841 (N_5841,N_4802,N_4903);
nand U5842 (N_5842,N_5241,N_4938);
nand U5843 (N_5843,N_5017,N_4989);
nor U5844 (N_5844,N_4799,N_4792);
nor U5845 (N_5845,N_4831,N_4782);
nor U5846 (N_5846,N_5098,N_5222);
and U5847 (N_5847,N_5116,N_5200);
nand U5848 (N_5848,N_4833,N_4571);
or U5849 (N_5849,N_4850,N_4980);
nand U5850 (N_5850,N_5030,N_5118);
nor U5851 (N_5851,N_5029,N_4663);
or U5852 (N_5852,N_4633,N_4522);
and U5853 (N_5853,N_4777,N_5019);
and U5854 (N_5854,N_4523,N_5040);
and U5855 (N_5855,N_4613,N_4866);
and U5856 (N_5856,N_4891,N_4670);
and U5857 (N_5857,N_4778,N_4516);
nand U5858 (N_5858,N_5003,N_4989);
nor U5859 (N_5859,N_5160,N_4704);
and U5860 (N_5860,N_4612,N_4532);
or U5861 (N_5861,N_5226,N_5211);
and U5862 (N_5862,N_4941,N_4545);
nand U5863 (N_5863,N_4946,N_4526);
nand U5864 (N_5864,N_5202,N_5054);
and U5865 (N_5865,N_4723,N_4726);
nand U5866 (N_5866,N_4537,N_4691);
xor U5867 (N_5867,N_5041,N_5090);
and U5868 (N_5868,N_4785,N_4805);
and U5869 (N_5869,N_5203,N_5169);
and U5870 (N_5870,N_4760,N_5078);
xnor U5871 (N_5871,N_4703,N_5237);
or U5872 (N_5872,N_4505,N_4863);
nor U5873 (N_5873,N_4947,N_4652);
nand U5874 (N_5874,N_5008,N_5118);
or U5875 (N_5875,N_4696,N_5209);
nor U5876 (N_5876,N_5161,N_5085);
and U5877 (N_5877,N_4780,N_5077);
and U5878 (N_5878,N_4630,N_4866);
and U5879 (N_5879,N_5182,N_4816);
nor U5880 (N_5880,N_4960,N_4863);
and U5881 (N_5881,N_4653,N_4631);
nand U5882 (N_5882,N_4649,N_4667);
nor U5883 (N_5883,N_5064,N_5149);
or U5884 (N_5884,N_4807,N_5039);
and U5885 (N_5885,N_4520,N_4783);
nor U5886 (N_5886,N_4643,N_4532);
and U5887 (N_5887,N_4566,N_4812);
and U5888 (N_5888,N_4536,N_5186);
or U5889 (N_5889,N_4915,N_4755);
nor U5890 (N_5890,N_4774,N_4602);
nor U5891 (N_5891,N_4858,N_5054);
nand U5892 (N_5892,N_4606,N_4930);
nor U5893 (N_5893,N_4971,N_4646);
or U5894 (N_5894,N_4659,N_5130);
or U5895 (N_5895,N_5218,N_4526);
or U5896 (N_5896,N_4696,N_5042);
and U5897 (N_5897,N_5062,N_4814);
or U5898 (N_5898,N_4702,N_5061);
nand U5899 (N_5899,N_4659,N_4573);
nand U5900 (N_5900,N_4983,N_4857);
and U5901 (N_5901,N_5096,N_4634);
nor U5902 (N_5902,N_5216,N_4690);
and U5903 (N_5903,N_4871,N_4727);
or U5904 (N_5904,N_4828,N_4614);
and U5905 (N_5905,N_4900,N_4735);
or U5906 (N_5906,N_4658,N_4659);
or U5907 (N_5907,N_5027,N_5218);
or U5908 (N_5908,N_5180,N_4726);
and U5909 (N_5909,N_4688,N_4830);
or U5910 (N_5910,N_5084,N_4510);
nand U5911 (N_5911,N_5097,N_4790);
nor U5912 (N_5912,N_5068,N_5130);
or U5913 (N_5913,N_5069,N_4778);
nand U5914 (N_5914,N_5209,N_4707);
or U5915 (N_5915,N_5069,N_5042);
nor U5916 (N_5916,N_4532,N_5192);
and U5917 (N_5917,N_4563,N_4707);
nor U5918 (N_5918,N_4593,N_4516);
nand U5919 (N_5919,N_5114,N_5117);
nor U5920 (N_5920,N_4923,N_4587);
and U5921 (N_5921,N_5248,N_4906);
nand U5922 (N_5922,N_4784,N_5175);
or U5923 (N_5923,N_4659,N_4889);
nor U5924 (N_5924,N_4986,N_5055);
nand U5925 (N_5925,N_5233,N_5095);
or U5926 (N_5926,N_4522,N_4897);
nor U5927 (N_5927,N_4823,N_4691);
nand U5928 (N_5928,N_4985,N_5026);
and U5929 (N_5929,N_4983,N_4855);
or U5930 (N_5930,N_5223,N_4518);
and U5931 (N_5931,N_4790,N_4600);
nor U5932 (N_5932,N_5209,N_4506);
nor U5933 (N_5933,N_5160,N_5120);
and U5934 (N_5934,N_5230,N_4901);
and U5935 (N_5935,N_5138,N_4520);
or U5936 (N_5936,N_4880,N_4790);
and U5937 (N_5937,N_5125,N_5046);
nand U5938 (N_5938,N_4959,N_4761);
and U5939 (N_5939,N_5035,N_4898);
nand U5940 (N_5940,N_5229,N_4637);
and U5941 (N_5941,N_4681,N_4826);
or U5942 (N_5942,N_4608,N_5079);
and U5943 (N_5943,N_4686,N_4794);
nor U5944 (N_5944,N_4670,N_5181);
xor U5945 (N_5945,N_4824,N_5222);
nand U5946 (N_5946,N_4555,N_4831);
and U5947 (N_5947,N_4885,N_4960);
or U5948 (N_5948,N_4862,N_4900);
nand U5949 (N_5949,N_4916,N_4744);
and U5950 (N_5950,N_5187,N_4896);
nor U5951 (N_5951,N_5028,N_4620);
nand U5952 (N_5952,N_4581,N_4834);
nor U5953 (N_5953,N_4717,N_5132);
nand U5954 (N_5954,N_4511,N_4692);
and U5955 (N_5955,N_4789,N_5098);
nor U5956 (N_5956,N_5135,N_4598);
nand U5957 (N_5957,N_4567,N_4585);
xor U5958 (N_5958,N_4833,N_4589);
or U5959 (N_5959,N_4663,N_4611);
and U5960 (N_5960,N_5087,N_4877);
nand U5961 (N_5961,N_4929,N_4598);
nand U5962 (N_5962,N_5235,N_5025);
nor U5963 (N_5963,N_4833,N_5109);
nand U5964 (N_5964,N_4520,N_5157);
and U5965 (N_5965,N_4526,N_4528);
or U5966 (N_5966,N_4791,N_5002);
nand U5967 (N_5967,N_4791,N_5000);
nand U5968 (N_5968,N_5120,N_4756);
or U5969 (N_5969,N_4732,N_4780);
and U5970 (N_5970,N_4783,N_5069);
nand U5971 (N_5971,N_5062,N_4638);
nand U5972 (N_5972,N_4848,N_4549);
nand U5973 (N_5973,N_4590,N_4816);
and U5974 (N_5974,N_5092,N_4680);
or U5975 (N_5975,N_4567,N_5128);
and U5976 (N_5976,N_4911,N_4506);
and U5977 (N_5977,N_5089,N_5136);
or U5978 (N_5978,N_5175,N_5243);
xnor U5979 (N_5979,N_4916,N_5104);
nand U5980 (N_5980,N_5101,N_4515);
or U5981 (N_5981,N_4520,N_5220);
and U5982 (N_5982,N_4817,N_4512);
and U5983 (N_5983,N_4786,N_5178);
or U5984 (N_5984,N_5111,N_4548);
nor U5985 (N_5985,N_4685,N_5000);
nor U5986 (N_5986,N_4706,N_4517);
xnor U5987 (N_5987,N_4765,N_4962);
or U5988 (N_5988,N_5109,N_5207);
and U5989 (N_5989,N_5137,N_5072);
nand U5990 (N_5990,N_5175,N_5104);
and U5991 (N_5991,N_4798,N_4667);
nor U5992 (N_5992,N_5016,N_5119);
nor U5993 (N_5993,N_4683,N_5168);
or U5994 (N_5994,N_4545,N_4803);
nand U5995 (N_5995,N_5064,N_5148);
or U5996 (N_5996,N_4824,N_4822);
nand U5997 (N_5997,N_4947,N_5144);
and U5998 (N_5998,N_4989,N_4751);
or U5999 (N_5999,N_5090,N_5203);
and U6000 (N_6000,N_5548,N_5499);
or U6001 (N_6001,N_5566,N_5629);
or U6002 (N_6002,N_5437,N_5380);
or U6003 (N_6003,N_5733,N_5607);
nand U6004 (N_6004,N_5891,N_5585);
and U6005 (N_6005,N_5333,N_5630);
and U6006 (N_6006,N_5800,N_5671);
nand U6007 (N_6007,N_5645,N_5513);
nand U6008 (N_6008,N_5668,N_5913);
nor U6009 (N_6009,N_5856,N_5572);
nor U6010 (N_6010,N_5732,N_5852);
or U6011 (N_6011,N_5392,N_5324);
nor U6012 (N_6012,N_5640,N_5610);
and U6013 (N_6013,N_5721,N_5446);
nand U6014 (N_6014,N_5745,N_5691);
or U6015 (N_6015,N_5811,N_5367);
nand U6016 (N_6016,N_5617,N_5754);
nand U6017 (N_6017,N_5942,N_5558);
nor U6018 (N_6018,N_5632,N_5991);
or U6019 (N_6019,N_5264,N_5330);
nor U6020 (N_6020,N_5878,N_5468);
and U6021 (N_6021,N_5717,N_5709);
or U6022 (N_6022,N_5426,N_5345);
and U6023 (N_6023,N_5821,N_5714);
nand U6024 (N_6024,N_5778,N_5809);
nor U6025 (N_6025,N_5712,N_5390);
or U6026 (N_6026,N_5934,N_5310);
nor U6027 (N_6027,N_5602,N_5600);
nor U6028 (N_6028,N_5883,N_5447);
nand U6029 (N_6029,N_5478,N_5995);
or U6030 (N_6030,N_5603,N_5452);
nor U6031 (N_6031,N_5419,N_5894);
and U6032 (N_6032,N_5787,N_5824);
or U6033 (N_6033,N_5764,N_5965);
and U6034 (N_6034,N_5615,N_5291);
nand U6035 (N_6035,N_5368,N_5693);
nor U6036 (N_6036,N_5501,N_5338);
and U6037 (N_6037,N_5592,N_5285);
nand U6038 (N_6038,N_5861,N_5805);
or U6039 (N_6039,N_5842,N_5837);
nand U6040 (N_6040,N_5850,N_5922);
nor U6041 (N_6041,N_5619,N_5540);
nor U6042 (N_6042,N_5797,N_5584);
nor U6043 (N_6043,N_5760,N_5502);
and U6044 (N_6044,N_5955,N_5892);
nand U6045 (N_6045,N_5986,N_5288);
and U6046 (N_6046,N_5876,N_5576);
and U6047 (N_6047,N_5959,N_5573);
nand U6048 (N_6048,N_5961,N_5574);
and U6049 (N_6049,N_5967,N_5661);
or U6050 (N_6050,N_5863,N_5460);
and U6051 (N_6051,N_5308,N_5870);
and U6052 (N_6052,N_5362,N_5461);
or U6053 (N_6053,N_5316,N_5329);
and U6054 (N_6054,N_5723,N_5365);
or U6055 (N_6055,N_5261,N_5512);
or U6056 (N_6056,N_5351,N_5289);
nand U6057 (N_6057,N_5425,N_5530);
and U6058 (N_6058,N_5653,N_5341);
or U6059 (N_6059,N_5579,N_5686);
nand U6060 (N_6060,N_5356,N_5253);
or U6061 (N_6061,N_5500,N_5747);
and U6062 (N_6062,N_5265,N_5947);
nor U6063 (N_6063,N_5780,N_5618);
or U6064 (N_6064,N_5560,N_5484);
or U6065 (N_6065,N_5458,N_5921);
nand U6066 (N_6066,N_5314,N_5533);
xor U6067 (N_6067,N_5940,N_5812);
and U6068 (N_6068,N_5660,N_5334);
nand U6069 (N_6069,N_5793,N_5542);
or U6070 (N_6070,N_5267,N_5552);
nand U6071 (N_6071,N_5422,N_5677);
and U6072 (N_6072,N_5923,N_5377);
and U6073 (N_6073,N_5424,N_5428);
and U6074 (N_6074,N_5399,N_5734);
and U6075 (N_6075,N_5514,N_5374);
or U6076 (N_6076,N_5725,N_5969);
nand U6077 (N_6077,N_5486,N_5873);
nor U6078 (N_6078,N_5381,N_5930);
nor U6079 (N_6079,N_5538,N_5252);
and U6080 (N_6080,N_5938,N_5694);
nor U6081 (N_6081,N_5667,N_5698);
nand U6082 (N_6082,N_5335,N_5565);
nor U6083 (N_6083,N_5866,N_5304);
nand U6084 (N_6084,N_5373,N_5358);
and U6085 (N_6085,N_5646,N_5864);
and U6086 (N_6086,N_5601,N_5407);
or U6087 (N_6087,N_5872,N_5492);
and U6088 (N_6088,N_5404,N_5716);
or U6089 (N_6089,N_5874,N_5744);
or U6090 (N_6090,N_5700,N_5774);
and U6091 (N_6091,N_5559,N_5944);
and U6092 (N_6092,N_5784,N_5675);
xnor U6093 (N_6093,N_5280,N_5976);
and U6094 (N_6094,N_5956,N_5846);
or U6095 (N_6095,N_5975,N_5755);
and U6096 (N_6096,N_5427,N_5665);
nand U6097 (N_6097,N_5349,N_5928);
nor U6098 (N_6098,N_5914,N_5283);
and U6099 (N_6099,N_5884,N_5912);
or U6100 (N_6100,N_5457,N_5357);
or U6101 (N_6101,N_5647,N_5806);
and U6102 (N_6102,N_5522,N_5897);
nand U6103 (N_6103,N_5266,N_5526);
or U6104 (N_6104,N_5933,N_5803);
nor U6105 (N_6105,N_5498,N_5997);
nand U6106 (N_6106,N_5529,N_5409);
nand U6107 (N_6107,N_5580,N_5752);
nor U6108 (N_6108,N_5871,N_5295);
or U6109 (N_6109,N_5282,N_5818);
nor U6110 (N_6110,N_5284,N_5463);
nand U6111 (N_6111,N_5383,N_5909);
and U6112 (N_6112,N_5396,N_5477);
and U6113 (N_6113,N_5702,N_5516);
nand U6114 (N_6114,N_5858,N_5844);
or U6115 (N_6115,N_5964,N_5379);
and U6116 (N_6116,N_5386,N_5773);
and U6117 (N_6117,N_5370,N_5624);
nor U6118 (N_6118,N_5342,N_5294);
and U6119 (N_6119,N_5493,N_5410);
or U6120 (N_6120,N_5465,N_5537);
nand U6121 (N_6121,N_5631,N_5801);
nor U6122 (N_6122,N_5766,N_5688);
nor U6123 (N_6123,N_5527,N_5518);
and U6124 (N_6124,N_5920,N_5826);
or U6125 (N_6125,N_5637,N_5550);
or U6126 (N_6126,N_5974,N_5697);
nand U6127 (N_6127,N_5577,N_5759);
nor U6128 (N_6128,N_5590,N_5785);
or U6129 (N_6129,N_5321,N_5328);
or U6130 (N_6130,N_5950,N_5937);
nor U6131 (N_6131,N_5347,N_5926);
and U6132 (N_6132,N_5534,N_5834);
or U6133 (N_6133,N_5730,N_5366);
and U6134 (N_6134,N_5751,N_5663);
nor U6135 (N_6135,N_5739,N_5385);
nand U6136 (N_6136,N_5907,N_5382);
and U6137 (N_6137,N_5886,N_5554);
nor U6138 (N_6138,N_5517,N_5925);
nand U6139 (N_6139,N_5839,N_5626);
or U6140 (N_6140,N_5319,N_5935);
nand U6141 (N_6141,N_5960,N_5911);
or U6142 (N_6142,N_5450,N_5662);
nor U6143 (N_6143,N_5757,N_5679);
xnor U6144 (N_6144,N_5337,N_5401);
nor U6145 (N_6145,N_5474,N_5491);
nor U6146 (N_6146,N_5352,N_5664);
or U6147 (N_6147,N_5256,N_5438);
nor U6148 (N_6148,N_5707,N_5482);
nand U6149 (N_6149,N_5808,N_5369);
nor U6150 (N_6150,N_5810,N_5682);
or U6151 (N_6151,N_5982,N_5855);
and U6152 (N_6152,N_5957,N_5887);
or U6153 (N_6153,N_5790,N_5741);
nor U6154 (N_6154,N_5900,N_5431);
nor U6155 (N_6155,N_5494,N_5789);
nand U6156 (N_6156,N_5623,N_5509);
or U6157 (N_6157,N_5555,N_5924);
and U6158 (N_6158,N_5731,N_5905);
nand U6159 (N_6159,N_5859,N_5633);
and U6160 (N_6160,N_5795,N_5339);
nand U6161 (N_6161,N_5670,N_5817);
nand U6162 (N_6162,N_5415,N_5588);
or U6163 (N_6163,N_5363,N_5454);
nor U6164 (N_6164,N_5881,N_5853);
or U6165 (N_6165,N_5849,N_5326);
nand U6166 (N_6166,N_5353,N_5860);
or U6167 (N_6167,N_5958,N_5567);
or U6168 (N_6168,N_5654,N_5348);
nor U6169 (N_6169,N_5388,N_5779);
nor U6170 (N_6170,N_5504,N_5292);
nand U6171 (N_6171,N_5830,N_5948);
or U6172 (N_6172,N_5286,N_5262);
nand U6173 (N_6173,N_5690,N_5656);
nand U6174 (N_6174,N_5359,N_5402);
and U6175 (N_6175,N_5740,N_5625);
and U6176 (N_6176,N_5543,N_5993);
and U6177 (N_6177,N_5609,N_5657);
and U6178 (N_6178,N_5479,N_5445);
nor U6179 (N_6179,N_5487,N_5398);
nand U6180 (N_6180,N_5258,N_5724);
nand U6181 (N_6181,N_5753,N_5704);
or U6182 (N_6182,N_5564,N_5932);
or U6183 (N_6183,N_5539,N_5776);
or U6184 (N_6184,N_5838,N_5756);
xor U6185 (N_6185,N_5476,N_5557);
nor U6186 (N_6186,N_5750,N_5836);
or U6187 (N_6187,N_5489,N_5765);
nor U6188 (N_6188,N_5520,N_5678);
nor U6189 (N_6189,N_5699,N_5620);
or U6190 (N_6190,N_5898,N_5815);
nand U6191 (N_6191,N_5762,N_5503);
or U6192 (N_6192,N_5880,N_5831);
and U6193 (N_6193,N_5825,N_5442);
and U6194 (N_6194,N_5397,N_5391);
or U6195 (N_6195,N_5984,N_5464);
or U6196 (N_6196,N_5648,N_5443);
nand U6197 (N_6197,N_5908,N_5655);
nand U6198 (N_6198,N_5346,N_5918);
nand U6199 (N_6199,N_5736,N_5738);
nand U6200 (N_6200,N_5775,N_5638);
nand U6201 (N_6201,N_5901,N_5593);
and U6202 (N_6202,N_5666,N_5250);
nor U6203 (N_6203,N_5395,N_5293);
nor U6204 (N_6204,N_5372,N_5435);
or U6205 (N_6205,N_5659,N_5720);
nor U6206 (N_6206,N_5695,N_5405);
nor U6207 (N_6207,N_5896,N_5783);
or U6208 (N_6208,N_5804,N_5416);
or U6209 (N_6209,N_5336,N_5862);
and U6210 (N_6210,N_5945,N_5962);
xnor U6211 (N_6211,N_5269,N_5432);
or U6212 (N_6212,N_5816,N_5758);
nor U6213 (N_6213,N_5641,N_5952);
or U6214 (N_6214,N_5763,N_5578);
nor U6215 (N_6215,N_5318,N_5701);
nor U6216 (N_6216,N_5888,N_5939);
or U6217 (N_6217,N_5551,N_5323);
or U6218 (N_6218,N_5541,N_5596);
nand U6219 (N_6219,N_5575,N_5469);
nor U6220 (N_6220,N_5389,N_5915);
or U6221 (N_6221,N_5545,N_5865);
nand U6222 (N_6222,N_5899,N_5384);
and U6223 (N_6223,N_5927,N_5473);
and U6224 (N_6224,N_5919,N_5378);
or U6225 (N_6225,N_5819,N_5355);
and U6226 (N_6226,N_5587,N_5260);
and U6227 (N_6227,N_5791,N_5583);
xnor U6228 (N_6228,N_5710,N_5510);
or U6229 (N_6229,N_5992,N_5544);
or U6230 (N_6230,N_5658,N_5413);
and U6231 (N_6231,N_5393,N_5561);
or U6232 (N_6232,N_5423,N_5715);
nor U6233 (N_6233,N_5488,N_5987);
nor U6234 (N_6234,N_5255,N_5718);
and U6235 (N_6235,N_5781,N_5794);
nor U6236 (N_6236,N_5951,N_5949);
nor U6237 (N_6237,N_5879,N_5418);
and U6238 (N_6238,N_5306,N_5331);
nor U6239 (N_6239,N_5279,N_5275);
nand U6240 (N_6240,N_5820,N_5594);
nand U6241 (N_6241,N_5867,N_5854);
and U6242 (N_6242,N_5636,N_5589);
nor U6243 (N_6243,N_5315,N_5614);
nand U6244 (N_6244,N_5851,N_5713);
nand U6245 (N_6245,N_5444,N_5521);
xnor U6246 (N_6246,N_5449,N_5400);
nor U6247 (N_6247,N_5728,N_5361);
and U6248 (N_6248,N_5711,N_5649);
nand U6249 (N_6249,N_5799,N_5508);
or U6250 (N_6250,N_5344,N_5971);
or U6251 (N_6251,N_5466,N_5953);
or U6252 (N_6252,N_5471,N_5313);
and U6253 (N_6253,N_5403,N_5340);
nor U6254 (N_6254,N_5273,N_5481);
or U6255 (N_6255,N_5563,N_5978);
nor U6256 (N_6256,N_5259,N_5505);
nand U6257 (N_6257,N_5582,N_5581);
nor U6258 (N_6258,N_5524,N_5606);
nand U6259 (N_6259,N_5634,N_5777);
or U6260 (N_6260,N_5515,N_5681);
nor U6261 (N_6261,N_5742,N_5767);
nor U6262 (N_6262,N_5868,N_5436);
or U6263 (N_6263,N_5893,N_5568);
nand U6264 (N_6264,N_5943,N_5470);
and U6265 (N_6265,N_5772,N_5475);
and U6266 (N_6266,N_5325,N_5414);
or U6267 (N_6267,N_5485,N_5983);
nand U6268 (N_6268,N_5299,N_5364);
nand U6269 (N_6269,N_5547,N_5727);
or U6270 (N_6270,N_5317,N_5985);
nand U6271 (N_6271,N_5535,N_5696);
nand U6272 (N_6272,N_5683,N_5546);
nand U6273 (N_6273,N_5743,N_5375);
and U6274 (N_6274,N_5954,N_5980);
and U6275 (N_6275,N_5376,N_5350);
xor U6276 (N_6276,N_5519,N_5703);
nand U6277 (N_6277,N_5902,N_5506);
or U6278 (N_6278,N_5309,N_5936);
or U6279 (N_6279,N_5495,N_5613);
nor U6280 (N_6280,N_5472,N_5343);
or U6281 (N_6281,N_5769,N_5684);
nor U6282 (N_6282,N_5611,N_5360);
or U6283 (N_6283,N_5672,N_5748);
or U6284 (N_6284,N_5977,N_5644);
or U6285 (N_6285,N_5455,N_5706);
nand U6286 (N_6286,N_5417,N_5796);
and U6287 (N_6287,N_5788,N_5798);
nor U6288 (N_6288,N_5483,N_5929);
or U6289 (N_6289,N_5628,N_5511);
or U6290 (N_6290,N_5467,N_5430);
or U6291 (N_6291,N_5999,N_5270);
nor U6292 (N_6292,N_5268,N_5412);
or U6293 (N_6293,N_5411,N_5642);
and U6294 (N_6294,N_5719,N_5332);
nand U6295 (N_6295,N_5296,N_5536);
or U6296 (N_6296,N_5271,N_5786);
or U6297 (N_6297,N_5705,N_5599);
and U6298 (N_6298,N_5674,N_5605);
and U6299 (N_6299,N_5327,N_5406);
and U6300 (N_6300,N_5746,N_5832);
nor U6301 (N_6301,N_5941,N_5591);
and U6302 (N_6302,N_5420,N_5301);
nor U6303 (N_6303,N_5440,N_5689);
nand U6304 (N_6304,N_5885,N_5278);
nand U6305 (N_6305,N_5973,N_5895);
and U6306 (N_6306,N_5737,N_5708);
or U6307 (N_6307,N_5595,N_5827);
nor U6308 (N_6308,N_5792,N_5312);
and U6309 (N_6309,N_5687,N_5889);
or U6310 (N_6310,N_5966,N_5290);
nor U6311 (N_6311,N_5835,N_5303);
nand U6312 (N_6312,N_5627,N_5571);
nor U6313 (N_6313,N_5990,N_5569);
nand U6314 (N_6314,N_5768,N_5612);
or U6315 (N_6315,N_5586,N_5823);
nor U6316 (N_6316,N_5525,N_5254);
nor U6317 (N_6317,N_5439,N_5813);
and U6318 (N_6318,N_5496,N_5877);
and U6319 (N_6319,N_5297,N_5770);
or U6320 (N_6320,N_5726,N_5875);
and U6321 (N_6321,N_5311,N_5643);
xor U6322 (N_6322,N_5639,N_5972);
nand U6323 (N_6323,N_5916,N_5685);
nand U6324 (N_6324,N_5998,N_5429);
or U6325 (N_6325,N_5621,N_5616);
or U6326 (N_6326,N_5300,N_5456);
nand U6327 (N_6327,N_5305,N_5845);
and U6328 (N_6328,N_5598,N_5970);
nand U6329 (N_6329,N_5833,N_5287);
nand U6330 (N_6330,N_5650,N_5729);
and U6331 (N_6331,N_5989,N_5570);
nor U6332 (N_6332,N_5652,N_5910);
xor U6333 (N_6333,N_5996,N_5302);
or U6334 (N_6334,N_5680,N_5994);
or U6335 (N_6335,N_5782,N_5807);
nand U6336 (N_6336,N_5276,N_5669);
and U6337 (N_6337,N_5433,N_5462);
or U6338 (N_6338,N_5274,N_5841);
and U6339 (N_6339,N_5840,N_5387);
nor U6340 (N_6340,N_5608,N_5802);
and U6341 (N_6341,N_5814,N_5394);
or U6342 (N_6342,N_5272,N_5277);
or U6343 (N_6343,N_5507,N_5263);
nand U6344 (N_6344,N_5981,N_5822);
or U6345 (N_6345,N_5553,N_5906);
or U6346 (N_6346,N_5979,N_5549);
or U6347 (N_6347,N_5408,N_5622);
nand U6348 (N_6348,N_5497,N_5651);
and U6349 (N_6349,N_5988,N_5869);
or U6350 (N_6350,N_5882,N_5917);
nor U6351 (N_6351,N_5890,N_5635);
nor U6352 (N_6352,N_5673,N_5857);
or U6353 (N_6353,N_5735,N_5421);
or U6354 (N_6354,N_5771,N_5298);
nor U6355 (N_6355,N_5453,N_5597);
and U6356 (N_6356,N_5904,N_5848);
nor U6357 (N_6357,N_5722,N_5843);
nor U6358 (N_6358,N_5281,N_5448);
and U6359 (N_6359,N_5354,N_5322);
nor U6360 (N_6360,N_5903,N_5441);
nor U6361 (N_6361,N_5968,N_5604);
and U6362 (N_6362,N_5562,N_5251);
nand U6363 (N_6363,N_5523,N_5761);
and U6364 (N_6364,N_5556,N_5829);
nor U6365 (N_6365,N_5528,N_5847);
and U6366 (N_6366,N_5828,N_5257);
nand U6367 (N_6367,N_5451,N_5490);
nor U6368 (N_6368,N_5531,N_5946);
nor U6369 (N_6369,N_5307,N_5692);
or U6370 (N_6370,N_5480,N_5676);
nor U6371 (N_6371,N_5371,N_5320);
nor U6372 (N_6372,N_5532,N_5963);
or U6373 (N_6373,N_5749,N_5931);
or U6374 (N_6374,N_5434,N_5459);
nor U6375 (N_6375,N_5568,N_5848);
and U6376 (N_6376,N_5302,N_5406);
and U6377 (N_6377,N_5861,N_5303);
nand U6378 (N_6378,N_5441,N_5427);
nand U6379 (N_6379,N_5744,N_5642);
and U6380 (N_6380,N_5373,N_5934);
nand U6381 (N_6381,N_5967,N_5614);
or U6382 (N_6382,N_5340,N_5353);
nand U6383 (N_6383,N_5812,N_5292);
or U6384 (N_6384,N_5922,N_5352);
nand U6385 (N_6385,N_5520,N_5650);
nand U6386 (N_6386,N_5287,N_5311);
nand U6387 (N_6387,N_5683,N_5283);
or U6388 (N_6388,N_5303,N_5837);
nand U6389 (N_6389,N_5264,N_5504);
and U6390 (N_6390,N_5676,N_5547);
and U6391 (N_6391,N_5610,N_5614);
and U6392 (N_6392,N_5731,N_5572);
nand U6393 (N_6393,N_5700,N_5975);
nor U6394 (N_6394,N_5527,N_5449);
nor U6395 (N_6395,N_5978,N_5501);
or U6396 (N_6396,N_5444,N_5743);
nand U6397 (N_6397,N_5685,N_5590);
nor U6398 (N_6398,N_5745,N_5306);
and U6399 (N_6399,N_5882,N_5802);
nand U6400 (N_6400,N_5952,N_5666);
nor U6401 (N_6401,N_5528,N_5456);
or U6402 (N_6402,N_5871,N_5328);
and U6403 (N_6403,N_5943,N_5337);
nor U6404 (N_6404,N_5840,N_5691);
and U6405 (N_6405,N_5686,N_5649);
nand U6406 (N_6406,N_5492,N_5585);
nand U6407 (N_6407,N_5978,N_5473);
nor U6408 (N_6408,N_5727,N_5518);
nor U6409 (N_6409,N_5922,N_5683);
nand U6410 (N_6410,N_5969,N_5960);
nor U6411 (N_6411,N_5807,N_5521);
and U6412 (N_6412,N_5864,N_5637);
nand U6413 (N_6413,N_5309,N_5566);
or U6414 (N_6414,N_5528,N_5722);
or U6415 (N_6415,N_5676,N_5608);
nor U6416 (N_6416,N_5710,N_5718);
and U6417 (N_6417,N_5549,N_5763);
nor U6418 (N_6418,N_5588,N_5675);
and U6419 (N_6419,N_5650,N_5922);
or U6420 (N_6420,N_5780,N_5844);
nor U6421 (N_6421,N_5776,N_5269);
and U6422 (N_6422,N_5753,N_5532);
nor U6423 (N_6423,N_5734,N_5414);
nor U6424 (N_6424,N_5760,N_5849);
or U6425 (N_6425,N_5679,N_5982);
and U6426 (N_6426,N_5426,N_5576);
nor U6427 (N_6427,N_5431,N_5619);
and U6428 (N_6428,N_5419,N_5890);
and U6429 (N_6429,N_5282,N_5618);
or U6430 (N_6430,N_5742,N_5476);
or U6431 (N_6431,N_5280,N_5888);
and U6432 (N_6432,N_5709,N_5646);
or U6433 (N_6433,N_5444,N_5259);
and U6434 (N_6434,N_5441,N_5251);
nor U6435 (N_6435,N_5541,N_5960);
and U6436 (N_6436,N_5264,N_5780);
and U6437 (N_6437,N_5446,N_5433);
or U6438 (N_6438,N_5652,N_5305);
nand U6439 (N_6439,N_5655,N_5768);
nand U6440 (N_6440,N_5954,N_5283);
nor U6441 (N_6441,N_5333,N_5292);
and U6442 (N_6442,N_5894,N_5388);
nor U6443 (N_6443,N_5506,N_5633);
or U6444 (N_6444,N_5521,N_5818);
nor U6445 (N_6445,N_5946,N_5851);
and U6446 (N_6446,N_5776,N_5373);
nor U6447 (N_6447,N_5963,N_5750);
nor U6448 (N_6448,N_5887,N_5580);
and U6449 (N_6449,N_5653,N_5776);
and U6450 (N_6450,N_5985,N_5612);
nor U6451 (N_6451,N_5766,N_5666);
or U6452 (N_6452,N_5506,N_5823);
and U6453 (N_6453,N_5315,N_5256);
nand U6454 (N_6454,N_5467,N_5471);
nor U6455 (N_6455,N_5365,N_5917);
nor U6456 (N_6456,N_5731,N_5308);
nand U6457 (N_6457,N_5554,N_5498);
nand U6458 (N_6458,N_5949,N_5414);
nand U6459 (N_6459,N_5424,N_5563);
or U6460 (N_6460,N_5351,N_5715);
or U6461 (N_6461,N_5779,N_5714);
nand U6462 (N_6462,N_5565,N_5269);
nand U6463 (N_6463,N_5795,N_5775);
nor U6464 (N_6464,N_5356,N_5837);
nand U6465 (N_6465,N_5608,N_5392);
nand U6466 (N_6466,N_5940,N_5671);
nand U6467 (N_6467,N_5862,N_5482);
nand U6468 (N_6468,N_5466,N_5736);
and U6469 (N_6469,N_5475,N_5527);
nor U6470 (N_6470,N_5897,N_5367);
or U6471 (N_6471,N_5840,N_5534);
and U6472 (N_6472,N_5812,N_5740);
nor U6473 (N_6473,N_5471,N_5262);
and U6474 (N_6474,N_5437,N_5416);
or U6475 (N_6475,N_5523,N_5987);
nor U6476 (N_6476,N_5912,N_5319);
nand U6477 (N_6477,N_5310,N_5816);
or U6478 (N_6478,N_5868,N_5283);
nor U6479 (N_6479,N_5406,N_5532);
or U6480 (N_6480,N_5940,N_5677);
and U6481 (N_6481,N_5394,N_5448);
nor U6482 (N_6482,N_5570,N_5561);
nand U6483 (N_6483,N_5953,N_5851);
or U6484 (N_6484,N_5727,N_5772);
nand U6485 (N_6485,N_5919,N_5426);
and U6486 (N_6486,N_5793,N_5292);
or U6487 (N_6487,N_5482,N_5663);
and U6488 (N_6488,N_5287,N_5776);
nand U6489 (N_6489,N_5293,N_5800);
nor U6490 (N_6490,N_5972,N_5702);
or U6491 (N_6491,N_5698,N_5682);
nor U6492 (N_6492,N_5685,N_5999);
nand U6493 (N_6493,N_5391,N_5629);
nor U6494 (N_6494,N_5524,N_5716);
or U6495 (N_6495,N_5735,N_5906);
nand U6496 (N_6496,N_5771,N_5310);
nor U6497 (N_6497,N_5898,N_5444);
and U6498 (N_6498,N_5374,N_5442);
and U6499 (N_6499,N_5313,N_5510);
and U6500 (N_6500,N_5938,N_5939);
nor U6501 (N_6501,N_5415,N_5768);
and U6502 (N_6502,N_5506,N_5576);
and U6503 (N_6503,N_5253,N_5976);
nor U6504 (N_6504,N_5963,N_5521);
nand U6505 (N_6505,N_5808,N_5393);
nor U6506 (N_6506,N_5373,N_5436);
and U6507 (N_6507,N_5999,N_5746);
or U6508 (N_6508,N_5325,N_5664);
and U6509 (N_6509,N_5501,N_5435);
nand U6510 (N_6510,N_5778,N_5776);
nand U6511 (N_6511,N_5528,N_5298);
and U6512 (N_6512,N_5544,N_5683);
nor U6513 (N_6513,N_5589,N_5686);
and U6514 (N_6514,N_5275,N_5764);
nor U6515 (N_6515,N_5644,N_5406);
nor U6516 (N_6516,N_5423,N_5912);
nor U6517 (N_6517,N_5912,N_5832);
nand U6518 (N_6518,N_5457,N_5513);
or U6519 (N_6519,N_5284,N_5954);
nor U6520 (N_6520,N_5860,N_5408);
and U6521 (N_6521,N_5618,N_5614);
nand U6522 (N_6522,N_5832,N_5876);
or U6523 (N_6523,N_5549,N_5627);
and U6524 (N_6524,N_5371,N_5755);
and U6525 (N_6525,N_5367,N_5673);
nand U6526 (N_6526,N_5427,N_5942);
nand U6527 (N_6527,N_5573,N_5942);
nor U6528 (N_6528,N_5943,N_5708);
nand U6529 (N_6529,N_5602,N_5850);
and U6530 (N_6530,N_5512,N_5493);
and U6531 (N_6531,N_5708,N_5270);
xnor U6532 (N_6532,N_5588,N_5719);
nor U6533 (N_6533,N_5515,N_5525);
nor U6534 (N_6534,N_5479,N_5361);
or U6535 (N_6535,N_5506,N_5303);
or U6536 (N_6536,N_5348,N_5766);
nand U6537 (N_6537,N_5581,N_5969);
and U6538 (N_6538,N_5426,N_5732);
or U6539 (N_6539,N_5566,N_5396);
nand U6540 (N_6540,N_5323,N_5298);
nand U6541 (N_6541,N_5449,N_5605);
nor U6542 (N_6542,N_5380,N_5577);
and U6543 (N_6543,N_5497,N_5881);
nor U6544 (N_6544,N_5890,N_5928);
and U6545 (N_6545,N_5676,N_5257);
and U6546 (N_6546,N_5574,N_5508);
nand U6547 (N_6547,N_5304,N_5336);
nor U6548 (N_6548,N_5649,N_5304);
or U6549 (N_6549,N_5374,N_5550);
and U6550 (N_6550,N_5698,N_5395);
nor U6551 (N_6551,N_5760,N_5356);
or U6552 (N_6552,N_5899,N_5726);
nand U6553 (N_6553,N_5434,N_5323);
and U6554 (N_6554,N_5729,N_5566);
nor U6555 (N_6555,N_5943,N_5880);
or U6556 (N_6556,N_5987,N_5875);
nand U6557 (N_6557,N_5924,N_5433);
nor U6558 (N_6558,N_5698,N_5428);
and U6559 (N_6559,N_5687,N_5971);
nor U6560 (N_6560,N_5924,N_5530);
nor U6561 (N_6561,N_5922,N_5265);
and U6562 (N_6562,N_5955,N_5906);
nand U6563 (N_6563,N_5632,N_5582);
or U6564 (N_6564,N_5813,N_5390);
nand U6565 (N_6565,N_5529,N_5833);
or U6566 (N_6566,N_5922,N_5663);
nand U6567 (N_6567,N_5843,N_5476);
and U6568 (N_6568,N_5844,N_5543);
and U6569 (N_6569,N_5926,N_5608);
nand U6570 (N_6570,N_5508,N_5461);
nand U6571 (N_6571,N_5369,N_5855);
or U6572 (N_6572,N_5502,N_5850);
or U6573 (N_6573,N_5695,N_5709);
nand U6574 (N_6574,N_5358,N_5439);
nand U6575 (N_6575,N_5945,N_5266);
and U6576 (N_6576,N_5472,N_5946);
nor U6577 (N_6577,N_5816,N_5558);
nor U6578 (N_6578,N_5508,N_5618);
nor U6579 (N_6579,N_5604,N_5466);
nand U6580 (N_6580,N_5920,N_5576);
nand U6581 (N_6581,N_5628,N_5633);
and U6582 (N_6582,N_5571,N_5893);
and U6583 (N_6583,N_5708,N_5441);
nand U6584 (N_6584,N_5251,N_5721);
or U6585 (N_6585,N_5696,N_5330);
and U6586 (N_6586,N_5507,N_5259);
nor U6587 (N_6587,N_5253,N_5886);
nand U6588 (N_6588,N_5697,N_5530);
nand U6589 (N_6589,N_5296,N_5392);
or U6590 (N_6590,N_5700,N_5525);
nor U6591 (N_6591,N_5714,N_5382);
or U6592 (N_6592,N_5733,N_5701);
nand U6593 (N_6593,N_5618,N_5395);
or U6594 (N_6594,N_5346,N_5488);
and U6595 (N_6595,N_5619,N_5746);
or U6596 (N_6596,N_5648,N_5378);
and U6597 (N_6597,N_5576,N_5371);
nor U6598 (N_6598,N_5366,N_5985);
nor U6599 (N_6599,N_5561,N_5833);
and U6600 (N_6600,N_5588,N_5396);
nor U6601 (N_6601,N_5594,N_5349);
nand U6602 (N_6602,N_5315,N_5645);
or U6603 (N_6603,N_5692,N_5551);
nand U6604 (N_6604,N_5792,N_5455);
nor U6605 (N_6605,N_5960,N_5533);
or U6606 (N_6606,N_5689,N_5944);
nor U6607 (N_6607,N_5933,N_5930);
nor U6608 (N_6608,N_5281,N_5340);
nand U6609 (N_6609,N_5300,N_5490);
or U6610 (N_6610,N_5628,N_5894);
or U6611 (N_6611,N_5280,N_5882);
or U6612 (N_6612,N_5977,N_5984);
nor U6613 (N_6613,N_5942,N_5526);
or U6614 (N_6614,N_5923,N_5903);
or U6615 (N_6615,N_5421,N_5491);
or U6616 (N_6616,N_5985,N_5265);
or U6617 (N_6617,N_5858,N_5390);
nor U6618 (N_6618,N_5924,N_5772);
nor U6619 (N_6619,N_5929,N_5926);
and U6620 (N_6620,N_5463,N_5451);
or U6621 (N_6621,N_5948,N_5667);
nand U6622 (N_6622,N_5874,N_5544);
xor U6623 (N_6623,N_5504,N_5748);
and U6624 (N_6624,N_5319,N_5889);
or U6625 (N_6625,N_5489,N_5964);
or U6626 (N_6626,N_5497,N_5536);
or U6627 (N_6627,N_5762,N_5333);
and U6628 (N_6628,N_5679,N_5607);
and U6629 (N_6629,N_5894,N_5844);
and U6630 (N_6630,N_5686,N_5517);
nor U6631 (N_6631,N_5401,N_5762);
nand U6632 (N_6632,N_5693,N_5525);
nor U6633 (N_6633,N_5748,N_5784);
nand U6634 (N_6634,N_5785,N_5366);
nor U6635 (N_6635,N_5366,N_5950);
nand U6636 (N_6636,N_5683,N_5627);
and U6637 (N_6637,N_5577,N_5715);
nand U6638 (N_6638,N_5393,N_5511);
or U6639 (N_6639,N_5330,N_5529);
nand U6640 (N_6640,N_5892,N_5836);
nand U6641 (N_6641,N_5785,N_5445);
nand U6642 (N_6642,N_5746,N_5346);
and U6643 (N_6643,N_5944,N_5252);
nor U6644 (N_6644,N_5680,N_5340);
nor U6645 (N_6645,N_5654,N_5880);
or U6646 (N_6646,N_5899,N_5503);
and U6647 (N_6647,N_5520,N_5400);
and U6648 (N_6648,N_5609,N_5713);
nand U6649 (N_6649,N_5792,N_5259);
or U6650 (N_6650,N_5268,N_5328);
nor U6651 (N_6651,N_5413,N_5448);
or U6652 (N_6652,N_5284,N_5660);
nand U6653 (N_6653,N_5706,N_5910);
or U6654 (N_6654,N_5341,N_5544);
nor U6655 (N_6655,N_5597,N_5497);
nor U6656 (N_6656,N_5804,N_5787);
nor U6657 (N_6657,N_5440,N_5751);
and U6658 (N_6658,N_5938,N_5848);
and U6659 (N_6659,N_5597,N_5306);
or U6660 (N_6660,N_5316,N_5650);
nor U6661 (N_6661,N_5835,N_5702);
and U6662 (N_6662,N_5330,N_5279);
or U6663 (N_6663,N_5560,N_5729);
nor U6664 (N_6664,N_5848,N_5886);
nand U6665 (N_6665,N_5616,N_5644);
and U6666 (N_6666,N_5388,N_5361);
nand U6667 (N_6667,N_5358,N_5409);
nand U6668 (N_6668,N_5845,N_5612);
nand U6669 (N_6669,N_5344,N_5829);
or U6670 (N_6670,N_5656,N_5415);
and U6671 (N_6671,N_5277,N_5449);
nor U6672 (N_6672,N_5597,N_5826);
or U6673 (N_6673,N_5554,N_5383);
and U6674 (N_6674,N_5541,N_5348);
nand U6675 (N_6675,N_5731,N_5559);
and U6676 (N_6676,N_5939,N_5770);
nor U6677 (N_6677,N_5297,N_5836);
or U6678 (N_6678,N_5397,N_5728);
nand U6679 (N_6679,N_5390,N_5323);
or U6680 (N_6680,N_5749,N_5901);
nand U6681 (N_6681,N_5579,N_5877);
nand U6682 (N_6682,N_5412,N_5346);
nor U6683 (N_6683,N_5364,N_5562);
nand U6684 (N_6684,N_5832,N_5722);
nand U6685 (N_6685,N_5482,N_5748);
nor U6686 (N_6686,N_5595,N_5559);
or U6687 (N_6687,N_5285,N_5327);
nor U6688 (N_6688,N_5547,N_5693);
or U6689 (N_6689,N_5619,N_5834);
or U6690 (N_6690,N_5289,N_5966);
or U6691 (N_6691,N_5994,N_5403);
nand U6692 (N_6692,N_5596,N_5395);
nor U6693 (N_6693,N_5783,N_5292);
nor U6694 (N_6694,N_5476,N_5615);
nand U6695 (N_6695,N_5412,N_5422);
or U6696 (N_6696,N_5855,N_5627);
or U6697 (N_6697,N_5806,N_5750);
nand U6698 (N_6698,N_5864,N_5480);
or U6699 (N_6699,N_5347,N_5972);
nand U6700 (N_6700,N_5250,N_5711);
nand U6701 (N_6701,N_5708,N_5823);
or U6702 (N_6702,N_5728,N_5839);
nor U6703 (N_6703,N_5658,N_5429);
nand U6704 (N_6704,N_5604,N_5804);
or U6705 (N_6705,N_5809,N_5629);
nand U6706 (N_6706,N_5822,N_5896);
xnor U6707 (N_6707,N_5310,N_5909);
nand U6708 (N_6708,N_5360,N_5523);
and U6709 (N_6709,N_5501,N_5317);
and U6710 (N_6710,N_5769,N_5900);
and U6711 (N_6711,N_5754,N_5843);
or U6712 (N_6712,N_5946,N_5326);
or U6713 (N_6713,N_5526,N_5514);
nor U6714 (N_6714,N_5411,N_5773);
or U6715 (N_6715,N_5608,N_5752);
nand U6716 (N_6716,N_5816,N_5786);
nand U6717 (N_6717,N_5547,N_5655);
and U6718 (N_6718,N_5463,N_5804);
nor U6719 (N_6719,N_5987,N_5653);
nand U6720 (N_6720,N_5904,N_5552);
and U6721 (N_6721,N_5308,N_5786);
nand U6722 (N_6722,N_5552,N_5871);
nor U6723 (N_6723,N_5532,N_5356);
nand U6724 (N_6724,N_5829,N_5526);
nor U6725 (N_6725,N_5369,N_5258);
and U6726 (N_6726,N_5848,N_5778);
and U6727 (N_6727,N_5584,N_5486);
or U6728 (N_6728,N_5994,N_5301);
nor U6729 (N_6729,N_5352,N_5322);
nand U6730 (N_6730,N_5980,N_5734);
nor U6731 (N_6731,N_5838,N_5426);
nand U6732 (N_6732,N_5714,N_5332);
or U6733 (N_6733,N_5771,N_5462);
nand U6734 (N_6734,N_5966,N_5404);
and U6735 (N_6735,N_5902,N_5991);
or U6736 (N_6736,N_5560,N_5544);
xnor U6737 (N_6737,N_5307,N_5827);
and U6738 (N_6738,N_5669,N_5366);
nand U6739 (N_6739,N_5598,N_5381);
nand U6740 (N_6740,N_5256,N_5648);
nor U6741 (N_6741,N_5317,N_5524);
or U6742 (N_6742,N_5868,N_5883);
nor U6743 (N_6743,N_5478,N_5808);
and U6744 (N_6744,N_5848,N_5832);
and U6745 (N_6745,N_5799,N_5692);
nand U6746 (N_6746,N_5475,N_5565);
nand U6747 (N_6747,N_5977,N_5258);
or U6748 (N_6748,N_5524,N_5278);
and U6749 (N_6749,N_5634,N_5878);
nor U6750 (N_6750,N_6260,N_6173);
nand U6751 (N_6751,N_6393,N_6674);
nand U6752 (N_6752,N_6680,N_6564);
nor U6753 (N_6753,N_6692,N_6205);
and U6754 (N_6754,N_6220,N_6481);
or U6755 (N_6755,N_6448,N_6523);
and U6756 (N_6756,N_6656,N_6585);
nor U6757 (N_6757,N_6050,N_6018);
nand U6758 (N_6758,N_6637,N_6199);
nor U6759 (N_6759,N_6715,N_6691);
nor U6760 (N_6760,N_6297,N_6302);
nor U6761 (N_6761,N_6693,N_6589);
or U6762 (N_6762,N_6280,N_6449);
nor U6763 (N_6763,N_6681,N_6417);
or U6764 (N_6764,N_6288,N_6643);
nor U6765 (N_6765,N_6093,N_6215);
and U6766 (N_6766,N_6565,N_6624);
and U6767 (N_6767,N_6248,N_6274);
nand U6768 (N_6768,N_6540,N_6476);
and U6769 (N_6769,N_6015,N_6272);
and U6770 (N_6770,N_6172,N_6039);
nor U6771 (N_6771,N_6709,N_6291);
or U6772 (N_6772,N_6223,N_6058);
and U6773 (N_6773,N_6703,N_6638);
or U6774 (N_6774,N_6433,N_6437);
nand U6775 (N_6775,N_6521,N_6002);
nor U6776 (N_6776,N_6699,N_6454);
and U6777 (N_6777,N_6456,N_6442);
and U6778 (N_6778,N_6701,N_6102);
nand U6779 (N_6779,N_6086,N_6380);
nor U6780 (N_6780,N_6636,N_6382);
nor U6781 (N_6781,N_6430,N_6561);
nand U6782 (N_6782,N_6211,N_6390);
or U6783 (N_6783,N_6101,N_6293);
or U6784 (N_6784,N_6295,N_6135);
or U6785 (N_6785,N_6161,N_6396);
nand U6786 (N_6786,N_6103,N_6661);
nor U6787 (N_6787,N_6096,N_6165);
nand U6788 (N_6788,N_6240,N_6076);
nor U6789 (N_6789,N_6209,N_6733);
nor U6790 (N_6790,N_6590,N_6458);
nor U6791 (N_6791,N_6163,N_6168);
nand U6792 (N_6792,N_6416,N_6089);
nand U6793 (N_6793,N_6330,N_6367);
or U6794 (N_6794,N_6016,N_6210);
or U6795 (N_6795,N_6517,N_6319);
nor U6796 (N_6796,N_6505,N_6546);
nand U6797 (N_6797,N_6337,N_6213);
nor U6798 (N_6798,N_6073,N_6418);
and U6799 (N_6799,N_6225,N_6035);
or U6800 (N_6800,N_6358,N_6524);
nand U6801 (N_6801,N_6542,N_6536);
and U6802 (N_6802,N_6728,N_6094);
or U6803 (N_6803,N_6494,N_6312);
nand U6804 (N_6804,N_6192,N_6239);
nand U6805 (N_6805,N_6045,N_6154);
nand U6806 (N_6806,N_6270,N_6510);
nor U6807 (N_6807,N_6645,N_6139);
and U6808 (N_6808,N_6175,N_6379);
and U6809 (N_6809,N_6028,N_6359);
or U6810 (N_6810,N_6164,N_6013);
and U6811 (N_6811,N_6356,N_6212);
or U6812 (N_6812,N_6233,N_6610);
or U6813 (N_6813,N_6552,N_6308);
and U6814 (N_6814,N_6608,N_6030);
or U6815 (N_6815,N_6554,N_6056);
or U6816 (N_6816,N_6112,N_6434);
nor U6817 (N_6817,N_6403,N_6227);
nand U6818 (N_6818,N_6604,N_6483);
nand U6819 (N_6819,N_6515,N_6612);
or U6820 (N_6820,N_6591,N_6653);
nor U6821 (N_6821,N_6189,N_6625);
nor U6822 (N_6822,N_6607,N_6644);
nor U6823 (N_6823,N_6063,N_6556);
nand U6824 (N_6824,N_6120,N_6547);
and U6825 (N_6825,N_6595,N_6660);
and U6826 (N_6826,N_6493,N_6374);
nor U6827 (N_6827,N_6115,N_6499);
nand U6828 (N_6828,N_6057,N_6593);
and U6829 (N_6829,N_6187,N_6679);
or U6830 (N_6830,N_6108,N_6221);
or U6831 (N_6831,N_6070,N_6560);
and U6832 (N_6832,N_6357,N_6282);
or U6833 (N_6833,N_6306,N_6052);
nor U6834 (N_6834,N_6512,N_6346);
and U6835 (N_6835,N_6329,N_6577);
or U6836 (N_6836,N_6235,N_6649);
or U6837 (N_6837,N_6271,N_6046);
nor U6838 (N_6838,N_6150,N_6324);
or U6839 (N_6839,N_6010,N_6498);
and U6840 (N_6840,N_6341,N_6415);
or U6841 (N_6841,N_6325,N_6311);
nor U6842 (N_6842,N_6659,N_6019);
and U6843 (N_6843,N_6368,N_6074);
nor U6844 (N_6844,N_6520,N_6605);
nand U6845 (N_6845,N_6746,N_6206);
or U6846 (N_6846,N_6229,N_6177);
or U6847 (N_6847,N_6237,N_6395);
nor U6848 (N_6848,N_6048,N_6640);
and U6849 (N_6849,N_6180,N_6409);
nor U6850 (N_6850,N_6726,N_6566);
or U6851 (N_6851,N_6158,N_6208);
nand U6852 (N_6852,N_6040,N_6735);
or U6853 (N_6853,N_6179,N_6686);
and U6854 (N_6854,N_6492,N_6252);
or U6855 (N_6855,N_6677,N_6570);
nand U6856 (N_6856,N_6537,N_6734);
or U6857 (N_6857,N_6062,N_6597);
nor U6858 (N_6858,N_6254,N_6087);
or U6859 (N_6859,N_6668,N_6317);
nand U6860 (N_6860,N_6632,N_6485);
or U6861 (N_6861,N_6472,N_6011);
or U6862 (N_6862,N_6279,N_6332);
or U6863 (N_6863,N_6557,N_6628);
nor U6864 (N_6864,N_6615,N_6569);
or U6865 (N_6865,N_6553,N_6104);
nor U6866 (N_6866,N_6447,N_6292);
nor U6867 (N_6867,N_6249,N_6082);
and U6868 (N_6868,N_6548,N_6479);
or U6869 (N_6869,N_6372,N_6322);
or U6870 (N_6870,N_6268,N_6061);
and U6871 (N_6871,N_6539,N_6344);
nand U6872 (N_6872,N_6331,N_6222);
xnor U6873 (N_6873,N_6694,N_6144);
and U6874 (N_6874,N_6360,N_6200);
or U6875 (N_6875,N_6670,N_6105);
nand U6876 (N_6876,N_6743,N_6214);
or U6877 (N_6877,N_6504,N_6256);
nand U6878 (N_6878,N_6518,N_6581);
or U6879 (N_6879,N_6353,N_6132);
or U6880 (N_6880,N_6054,N_6429);
or U6881 (N_6881,N_6246,N_6051);
or U6882 (N_6882,N_6722,N_6712);
and U6883 (N_6883,N_6174,N_6596);
nand U6884 (N_6884,N_6287,N_6384);
nor U6885 (N_6885,N_6592,N_6195);
nand U6886 (N_6886,N_6503,N_6606);
nor U6887 (N_6887,N_6435,N_6348);
nand U6888 (N_6888,N_6613,N_6444);
or U6889 (N_6889,N_6354,N_6113);
nand U6890 (N_6890,N_6641,N_6742);
and U6891 (N_6891,N_6497,N_6284);
nor U6892 (N_6892,N_6690,N_6029);
nor U6893 (N_6893,N_6309,N_6005);
nor U6894 (N_6894,N_6122,N_6041);
nand U6895 (N_6895,N_6190,N_6525);
nand U6896 (N_6896,N_6470,N_6304);
or U6897 (N_6897,N_6579,N_6068);
nor U6898 (N_6898,N_6488,N_6261);
xor U6899 (N_6899,N_6345,N_6738);
or U6900 (N_6900,N_6343,N_6391);
or U6901 (N_6901,N_6711,N_6529);
nand U6902 (N_6902,N_6106,N_6626);
and U6903 (N_6903,N_6737,N_6535);
nor U6904 (N_6904,N_6171,N_6355);
and U6905 (N_6905,N_6410,N_6658);
or U6906 (N_6906,N_6184,N_6020);
nand U6907 (N_6907,N_6422,N_6138);
nor U6908 (N_6908,N_6705,N_6662);
nand U6909 (N_6909,N_6037,N_6230);
nand U6910 (N_6910,N_6664,N_6559);
nand U6911 (N_6911,N_6185,N_6574);
nor U6912 (N_6912,N_6720,N_6477);
nor U6913 (N_6913,N_6397,N_6012);
or U6914 (N_6914,N_6219,N_6009);
or U6915 (N_6915,N_6032,N_6370);
nand U6916 (N_6916,N_6467,N_6134);
nor U6917 (N_6917,N_6081,N_6622);
nor U6918 (N_6918,N_6155,N_6080);
nand U6919 (N_6919,N_6003,N_6563);
nor U6920 (N_6920,N_6727,N_6069);
nand U6921 (N_6921,N_6310,N_6621);
nor U6922 (N_6922,N_6739,N_6299);
xnor U6923 (N_6923,N_6516,N_6001);
nand U6924 (N_6924,N_6716,N_6431);
nor U6925 (N_6925,N_6509,N_6474);
and U6926 (N_6926,N_6065,N_6111);
nor U6927 (N_6927,N_6684,N_6635);
nand U6928 (N_6928,N_6049,N_6421);
and U6929 (N_6929,N_6342,N_6339);
nor U6930 (N_6930,N_6313,N_6545);
nand U6931 (N_6931,N_6116,N_6673);
or U6932 (N_6932,N_6441,N_6480);
nand U6933 (N_6933,N_6736,N_6091);
xor U6934 (N_6934,N_6234,N_6501);
nor U6935 (N_6935,N_6623,N_6140);
and U6936 (N_6936,N_6486,N_6714);
nand U6937 (N_6937,N_6464,N_6603);
nor U6938 (N_6938,N_6098,N_6582);
nand U6939 (N_6939,N_6022,N_6698);
nor U6940 (N_6940,N_6267,N_6404);
or U6941 (N_6941,N_6126,N_6588);
and U6942 (N_6942,N_6201,N_6196);
and U6943 (N_6943,N_6601,N_6148);
or U6944 (N_6944,N_6482,N_6307);
and U6945 (N_6945,N_6289,N_6575);
nand U6946 (N_6946,N_6528,N_6451);
nand U6947 (N_6947,N_6713,N_6747);
nor U6948 (N_6948,N_6146,N_6576);
nand U6949 (N_6949,N_6176,N_6191);
or U6950 (N_6950,N_6696,N_6487);
and U6951 (N_6951,N_6710,N_6532);
nor U6952 (N_6952,N_6527,N_6262);
and U6953 (N_6953,N_6471,N_6259);
or U6954 (N_6954,N_6000,N_6303);
and U6955 (N_6955,N_6147,N_6149);
nor U6956 (N_6956,N_6241,N_6084);
and U6957 (N_6957,N_6064,N_6033);
or U6958 (N_6958,N_6247,N_6531);
nand U6959 (N_6959,N_6253,N_6700);
or U6960 (N_6960,N_6162,N_6478);
nand U6961 (N_6961,N_6425,N_6469);
and U6962 (N_6962,N_6169,N_6004);
nand U6963 (N_6963,N_6188,N_6055);
nand U6964 (N_6964,N_6408,N_6023);
and U6965 (N_6965,N_6182,N_6506);
and U6966 (N_6966,N_6017,N_6071);
xnor U6967 (N_6967,N_6678,N_6741);
and U6968 (N_6968,N_6630,N_6489);
or U6969 (N_6969,N_6450,N_6721);
or U6970 (N_6970,N_6669,N_6042);
nor U6971 (N_6971,N_6671,N_6377);
or U6972 (N_6972,N_6647,N_6465);
or U6973 (N_6973,N_6602,N_6530);
nor U6974 (N_6974,N_6336,N_6286);
or U6975 (N_6975,N_6301,N_6639);
and U6976 (N_6976,N_6383,N_6453);
and U6977 (N_6977,N_6133,N_6484);
nor U6978 (N_6978,N_6541,N_6060);
and U6979 (N_6979,N_6619,N_6092);
nor U6980 (N_6980,N_6142,N_6704);
nor U6981 (N_6981,N_6666,N_6723);
or U6982 (N_6982,N_6316,N_6683);
nor U6983 (N_6983,N_6244,N_6117);
or U6984 (N_6984,N_6347,N_6255);
nand U6985 (N_6985,N_6290,N_6014);
and U6986 (N_6986,N_6413,N_6202);
nor U6987 (N_6987,N_6567,N_6572);
nor U6988 (N_6988,N_6522,N_6651);
nor U6989 (N_6989,N_6036,N_6026);
nand U6990 (N_6990,N_6242,N_6587);
nor U6991 (N_6991,N_6243,N_6688);
nor U6992 (N_6992,N_6366,N_6405);
nand U6993 (N_6993,N_6538,N_6629);
nor U6994 (N_6994,N_6326,N_6167);
and U6995 (N_6995,N_6457,N_6131);
and U6996 (N_6996,N_6264,N_6654);
or U6997 (N_6997,N_6314,N_6077);
nor U6998 (N_6998,N_6697,N_6376);
and U6999 (N_6999,N_6725,N_6038);
or U7000 (N_7000,N_6152,N_6551);
nor U7001 (N_7001,N_6490,N_6695);
and U7002 (N_7002,N_6318,N_6406);
nor U7003 (N_7003,N_6034,N_6151);
nor U7004 (N_7004,N_6369,N_6315);
nand U7005 (N_7005,N_6729,N_6088);
and U7006 (N_7006,N_6207,N_6328);
and U7007 (N_7007,N_6047,N_6321);
xor U7008 (N_7008,N_6153,N_6466);
or U7009 (N_7009,N_6231,N_6507);
nor U7010 (N_7010,N_6266,N_6511);
nor U7011 (N_7011,N_6371,N_6333);
nor U7012 (N_7012,N_6238,N_6562);
nor U7013 (N_7013,N_6245,N_6351);
nand U7014 (N_7014,N_6285,N_6378);
and U7015 (N_7015,N_6445,N_6508);
nor U7016 (N_7016,N_6578,N_6276);
nand U7017 (N_7017,N_6526,N_6648);
nor U7018 (N_7018,N_6008,N_6475);
or U7019 (N_7019,N_6702,N_6443);
and U7020 (N_7020,N_6095,N_6110);
or U7021 (N_7021,N_6584,N_6394);
or U7022 (N_7022,N_6119,N_6228);
or U7023 (N_7023,N_6568,N_6534);
or U7024 (N_7024,N_6203,N_6611);
or U7025 (N_7025,N_6159,N_6634);
nand U7026 (N_7026,N_6197,N_6543);
or U7027 (N_7027,N_6412,N_6420);
and U7028 (N_7028,N_6294,N_6107);
and U7029 (N_7029,N_6125,N_6423);
nand U7030 (N_7030,N_6365,N_6401);
nand U7031 (N_7031,N_6387,N_6193);
nor U7032 (N_7032,N_6137,N_6687);
nor U7033 (N_7033,N_6599,N_6460);
and U7034 (N_7034,N_6426,N_6170);
or U7035 (N_7035,N_6263,N_6265);
and U7036 (N_7036,N_6439,N_6558);
xnor U7037 (N_7037,N_6078,N_6079);
nand U7038 (N_7038,N_6609,N_6657);
nand U7039 (N_7039,N_6427,N_6198);
or U7040 (N_7040,N_6514,N_6502);
nor U7041 (N_7041,N_6513,N_6281);
nor U7042 (N_7042,N_6130,N_6025);
nand U7043 (N_7043,N_6044,N_6118);
nor U7044 (N_7044,N_6186,N_6204);
nor U7045 (N_7045,N_6143,N_6226);
or U7046 (N_7046,N_6571,N_6500);
nor U7047 (N_7047,N_6685,N_6109);
nor U7048 (N_7048,N_6436,N_6361);
or U7049 (N_7049,N_6620,N_6349);
and U7050 (N_7050,N_6650,N_6402);
or U7051 (N_7051,N_6642,N_6617);
nor U7052 (N_7052,N_6682,N_6099);
nor U7053 (N_7053,N_6740,N_6128);
or U7054 (N_7054,N_6618,N_6006);
or U7055 (N_7055,N_6340,N_6224);
or U7056 (N_7056,N_6283,N_6352);
nand U7057 (N_7057,N_6550,N_6305);
nand U7058 (N_7058,N_6300,N_6533);
and U7059 (N_7059,N_6381,N_6127);
and U7060 (N_7060,N_6194,N_6021);
nand U7061 (N_7061,N_6440,N_6114);
or U7062 (N_7062,N_6446,N_6160);
nand U7063 (N_7063,N_6708,N_6549);
and U7064 (N_7064,N_6706,N_6277);
or U7065 (N_7065,N_6335,N_6491);
nand U7066 (N_7066,N_6166,N_6251);
nand U7067 (N_7067,N_6373,N_6217);
and U7068 (N_7068,N_6027,N_6375);
and U7069 (N_7069,N_6232,N_6555);
and U7070 (N_7070,N_6414,N_6675);
or U7071 (N_7071,N_6399,N_6544);
nor U7072 (N_7072,N_6072,N_6463);
and U7073 (N_7073,N_6236,N_6083);
nor U7074 (N_7074,N_6473,N_6633);
and U7075 (N_7075,N_6724,N_6419);
nand U7076 (N_7076,N_6455,N_6719);
and U7077 (N_7077,N_6327,N_6580);
and U7078 (N_7078,N_6136,N_6085);
nor U7079 (N_7079,N_6730,N_6732);
and U7080 (N_7080,N_6067,N_6438);
or U7081 (N_7081,N_6053,N_6689);
and U7082 (N_7082,N_6123,N_6278);
nand U7083 (N_7083,N_6461,N_6586);
nand U7084 (N_7084,N_6141,N_6655);
nor U7085 (N_7085,N_6178,N_6350);
nor U7086 (N_7086,N_6145,N_6432);
nand U7087 (N_7087,N_6424,N_6676);
and U7088 (N_7088,N_6667,N_6614);
nor U7089 (N_7089,N_6269,N_6124);
and U7090 (N_7090,N_6364,N_6257);
nor U7091 (N_7091,N_6388,N_6717);
and U7092 (N_7092,N_6452,N_6007);
nor U7093 (N_7093,N_6031,N_6400);
or U7094 (N_7094,N_6573,N_6298);
or U7095 (N_7095,N_6600,N_6672);
nor U7096 (N_7096,N_6459,N_6275);
or U7097 (N_7097,N_6258,N_6748);
and U7098 (N_7098,N_6129,N_6652);
nand U7099 (N_7099,N_6100,N_6273);
nand U7100 (N_7100,N_6090,N_6665);
and U7101 (N_7101,N_6392,N_6181);
or U7102 (N_7102,N_6462,N_6121);
and U7103 (N_7103,N_6744,N_6334);
nor U7104 (N_7104,N_6627,N_6646);
nor U7105 (N_7105,N_6594,N_6043);
or U7106 (N_7106,N_6183,N_6749);
or U7107 (N_7107,N_6157,N_6495);
or U7108 (N_7108,N_6216,N_6411);
nand U7109 (N_7109,N_6156,N_6598);
nand U7110 (N_7110,N_6616,N_6407);
nand U7111 (N_7111,N_6218,N_6362);
nand U7112 (N_7112,N_6323,N_6386);
and U7113 (N_7113,N_6663,N_6707);
or U7114 (N_7114,N_6583,N_6059);
and U7115 (N_7115,N_6468,N_6519);
nor U7116 (N_7116,N_6631,N_6363);
and U7117 (N_7117,N_6024,N_6097);
nand U7118 (N_7118,N_6718,N_6320);
or U7119 (N_7119,N_6731,N_6338);
or U7120 (N_7120,N_6250,N_6496);
or U7121 (N_7121,N_6296,N_6385);
and U7122 (N_7122,N_6389,N_6398);
nand U7123 (N_7123,N_6745,N_6066);
or U7124 (N_7124,N_6075,N_6428);
nor U7125 (N_7125,N_6034,N_6169);
and U7126 (N_7126,N_6020,N_6428);
and U7127 (N_7127,N_6520,N_6585);
or U7128 (N_7128,N_6098,N_6161);
and U7129 (N_7129,N_6603,N_6261);
nor U7130 (N_7130,N_6505,N_6266);
and U7131 (N_7131,N_6300,N_6651);
nand U7132 (N_7132,N_6747,N_6110);
nor U7133 (N_7133,N_6709,N_6491);
nand U7134 (N_7134,N_6110,N_6209);
and U7135 (N_7135,N_6031,N_6118);
and U7136 (N_7136,N_6570,N_6125);
xnor U7137 (N_7137,N_6371,N_6043);
or U7138 (N_7138,N_6456,N_6254);
nor U7139 (N_7139,N_6509,N_6324);
nor U7140 (N_7140,N_6209,N_6604);
or U7141 (N_7141,N_6609,N_6384);
nor U7142 (N_7142,N_6370,N_6727);
nor U7143 (N_7143,N_6472,N_6213);
nor U7144 (N_7144,N_6667,N_6408);
or U7145 (N_7145,N_6169,N_6610);
and U7146 (N_7146,N_6562,N_6364);
or U7147 (N_7147,N_6428,N_6315);
nor U7148 (N_7148,N_6006,N_6678);
and U7149 (N_7149,N_6634,N_6217);
nand U7150 (N_7150,N_6523,N_6227);
or U7151 (N_7151,N_6272,N_6441);
nand U7152 (N_7152,N_6326,N_6419);
and U7153 (N_7153,N_6545,N_6616);
and U7154 (N_7154,N_6447,N_6604);
nand U7155 (N_7155,N_6326,N_6039);
nand U7156 (N_7156,N_6731,N_6268);
nand U7157 (N_7157,N_6067,N_6031);
or U7158 (N_7158,N_6302,N_6460);
nor U7159 (N_7159,N_6453,N_6270);
and U7160 (N_7160,N_6516,N_6453);
nor U7161 (N_7161,N_6540,N_6483);
nor U7162 (N_7162,N_6604,N_6018);
or U7163 (N_7163,N_6610,N_6172);
nand U7164 (N_7164,N_6326,N_6088);
and U7165 (N_7165,N_6125,N_6498);
nand U7166 (N_7166,N_6513,N_6082);
or U7167 (N_7167,N_6472,N_6190);
nand U7168 (N_7168,N_6136,N_6036);
nor U7169 (N_7169,N_6589,N_6444);
or U7170 (N_7170,N_6560,N_6285);
or U7171 (N_7171,N_6231,N_6167);
nor U7172 (N_7172,N_6282,N_6525);
and U7173 (N_7173,N_6124,N_6384);
nand U7174 (N_7174,N_6369,N_6470);
or U7175 (N_7175,N_6326,N_6427);
or U7176 (N_7176,N_6481,N_6731);
or U7177 (N_7177,N_6347,N_6373);
or U7178 (N_7178,N_6292,N_6457);
nand U7179 (N_7179,N_6047,N_6204);
and U7180 (N_7180,N_6578,N_6523);
and U7181 (N_7181,N_6456,N_6534);
nand U7182 (N_7182,N_6501,N_6139);
and U7183 (N_7183,N_6207,N_6147);
and U7184 (N_7184,N_6555,N_6070);
and U7185 (N_7185,N_6583,N_6127);
nand U7186 (N_7186,N_6325,N_6655);
or U7187 (N_7187,N_6390,N_6278);
or U7188 (N_7188,N_6635,N_6016);
nand U7189 (N_7189,N_6262,N_6414);
and U7190 (N_7190,N_6063,N_6494);
nand U7191 (N_7191,N_6193,N_6076);
nand U7192 (N_7192,N_6394,N_6593);
nor U7193 (N_7193,N_6700,N_6627);
or U7194 (N_7194,N_6670,N_6725);
or U7195 (N_7195,N_6073,N_6396);
and U7196 (N_7196,N_6510,N_6633);
and U7197 (N_7197,N_6137,N_6406);
or U7198 (N_7198,N_6544,N_6369);
and U7199 (N_7199,N_6249,N_6747);
or U7200 (N_7200,N_6485,N_6541);
and U7201 (N_7201,N_6303,N_6419);
and U7202 (N_7202,N_6103,N_6674);
nor U7203 (N_7203,N_6292,N_6626);
or U7204 (N_7204,N_6144,N_6580);
and U7205 (N_7205,N_6228,N_6324);
or U7206 (N_7206,N_6618,N_6217);
and U7207 (N_7207,N_6595,N_6490);
nor U7208 (N_7208,N_6436,N_6486);
or U7209 (N_7209,N_6049,N_6524);
and U7210 (N_7210,N_6436,N_6543);
nand U7211 (N_7211,N_6070,N_6382);
or U7212 (N_7212,N_6021,N_6283);
nand U7213 (N_7213,N_6576,N_6673);
or U7214 (N_7214,N_6231,N_6015);
and U7215 (N_7215,N_6416,N_6485);
nand U7216 (N_7216,N_6211,N_6326);
and U7217 (N_7217,N_6503,N_6323);
xor U7218 (N_7218,N_6662,N_6336);
or U7219 (N_7219,N_6672,N_6028);
or U7220 (N_7220,N_6363,N_6000);
nor U7221 (N_7221,N_6079,N_6045);
or U7222 (N_7222,N_6489,N_6518);
and U7223 (N_7223,N_6611,N_6597);
or U7224 (N_7224,N_6242,N_6334);
nand U7225 (N_7225,N_6086,N_6432);
or U7226 (N_7226,N_6188,N_6184);
nand U7227 (N_7227,N_6017,N_6718);
and U7228 (N_7228,N_6634,N_6060);
and U7229 (N_7229,N_6636,N_6185);
and U7230 (N_7230,N_6303,N_6016);
or U7231 (N_7231,N_6729,N_6289);
and U7232 (N_7232,N_6395,N_6656);
nand U7233 (N_7233,N_6480,N_6023);
nor U7234 (N_7234,N_6223,N_6248);
and U7235 (N_7235,N_6619,N_6444);
nand U7236 (N_7236,N_6233,N_6292);
and U7237 (N_7237,N_6048,N_6293);
nor U7238 (N_7238,N_6704,N_6334);
nor U7239 (N_7239,N_6287,N_6719);
or U7240 (N_7240,N_6568,N_6243);
nand U7241 (N_7241,N_6717,N_6581);
nand U7242 (N_7242,N_6123,N_6191);
or U7243 (N_7243,N_6543,N_6110);
or U7244 (N_7244,N_6069,N_6416);
or U7245 (N_7245,N_6079,N_6238);
nand U7246 (N_7246,N_6662,N_6241);
and U7247 (N_7247,N_6402,N_6620);
or U7248 (N_7248,N_6010,N_6132);
nand U7249 (N_7249,N_6160,N_6059);
nand U7250 (N_7250,N_6009,N_6412);
or U7251 (N_7251,N_6326,N_6227);
nor U7252 (N_7252,N_6218,N_6150);
nand U7253 (N_7253,N_6445,N_6717);
or U7254 (N_7254,N_6050,N_6248);
and U7255 (N_7255,N_6730,N_6298);
nor U7256 (N_7256,N_6550,N_6509);
and U7257 (N_7257,N_6673,N_6505);
xnor U7258 (N_7258,N_6116,N_6526);
or U7259 (N_7259,N_6113,N_6150);
or U7260 (N_7260,N_6194,N_6436);
nor U7261 (N_7261,N_6099,N_6411);
nand U7262 (N_7262,N_6221,N_6706);
nor U7263 (N_7263,N_6261,N_6227);
nor U7264 (N_7264,N_6740,N_6049);
nor U7265 (N_7265,N_6030,N_6174);
nor U7266 (N_7266,N_6003,N_6505);
and U7267 (N_7267,N_6524,N_6685);
or U7268 (N_7268,N_6745,N_6729);
nor U7269 (N_7269,N_6232,N_6466);
nor U7270 (N_7270,N_6740,N_6117);
or U7271 (N_7271,N_6728,N_6137);
or U7272 (N_7272,N_6310,N_6401);
or U7273 (N_7273,N_6323,N_6112);
or U7274 (N_7274,N_6031,N_6191);
nor U7275 (N_7275,N_6138,N_6177);
or U7276 (N_7276,N_6740,N_6668);
nand U7277 (N_7277,N_6417,N_6159);
nor U7278 (N_7278,N_6549,N_6595);
and U7279 (N_7279,N_6050,N_6085);
nor U7280 (N_7280,N_6278,N_6654);
nand U7281 (N_7281,N_6138,N_6690);
or U7282 (N_7282,N_6228,N_6647);
and U7283 (N_7283,N_6235,N_6665);
nand U7284 (N_7284,N_6083,N_6574);
nor U7285 (N_7285,N_6126,N_6015);
or U7286 (N_7286,N_6561,N_6513);
or U7287 (N_7287,N_6190,N_6413);
or U7288 (N_7288,N_6602,N_6727);
or U7289 (N_7289,N_6317,N_6047);
nor U7290 (N_7290,N_6477,N_6412);
nand U7291 (N_7291,N_6716,N_6562);
nand U7292 (N_7292,N_6244,N_6589);
nor U7293 (N_7293,N_6605,N_6576);
or U7294 (N_7294,N_6100,N_6469);
and U7295 (N_7295,N_6429,N_6574);
nand U7296 (N_7296,N_6427,N_6355);
nand U7297 (N_7297,N_6503,N_6684);
nand U7298 (N_7298,N_6341,N_6722);
and U7299 (N_7299,N_6166,N_6745);
or U7300 (N_7300,N_6688,N_6042);
and U7301 (N_7301,N_6550,N_6633);
nand U7302 (N_7302,N_6162,N_6470);
and U7303 (N_7303,N_6022,N_6254);
and U7304 (N_7304,N_6553,N_6001);
and U7305 (N_7305,N_6480,N_6340);
or U7306 (N_7306,N_6265,N_6524);
and U7307 (N_7307,N_6231,N_6317);
nand U7308 (N_7308,N_6528,N_6061);
nor U7309 (N_7309,N_6506,N_6588);
or U7310 (N_7310,N_6495,N_6676);
or U7311 (N_7311,N_6687,N_6060);
nor U7312 (N_7312,N_6157,N_6603);
or U7313 (N_7313,N_6086,N_6172);
or U7314 (N_7314,N_6243,N_6086);
or U7315 (N_7315,N_6339,N_6116);
nand U7316 (N_7316,N_6383,N_6190);
and U7317 (N_7317,N_6376,N_6031);
and U7318 (N_7318,N_6387,N_6513);
or U7319 (N_7319,N_6004,N_6247);
nor U7320 (N_7320,N_6395,N_6467);
or U7321 (N_7321,N_6162,N_6342);
nand U7322 (N_7322,N_6324,N_6721);
nor U7323 (N_7323,N_6292,N_6365);
nor U7324 (N_7324,N_6520,N_6187);
or U7325 (N_7325,N_6725,N_6311);
and U7326 (N_7326,N_6048,N_6041);
and U7327 (N_7327,N_6496,N_6563);
nand U7328 (N_7328,N_6444,N_6665);
and U7329 (N_7329,N_6332,N_6429);
nor U7330 (N_7330,N_6481,N_6596);
nand U7331 (N_7331,N_6669,N_6722);
nor U7332 (N_7332,N_6687,N_6180);
nor U7333 (N_7333,N_6452,N_6462);
nor U7334 (N_7334,N_6511,N_6217);
or U7335 (N_7335,N_6590,N_6254);
or U7336 (N_7336,N_6521,N_6200);
nor U7337 (N_7337,N_6443,N_6585);
or U7338 (N_7338,N_6560,N_6241);
or U7339 (N_7339,N_6463,N_6390);
and U7340 (N_7340,N_6109,N_6329);
nand U7341 (N_7341,N_6337,N_6287);
or U7342 (N_7342,N_6731,N_6150);
nand U7343 (N_7343,N_6680,N_6236);
and U7344 (N_7344,N_6246,N_6442);
or U7345 (N_7345,N_6330,N_6093);
and U7346 (N_7346,N_6176,N_6279);
and U7347 (N_7347,N_6450,N_6657);
nand U7348 (N_7348,N_6089,N_6239);
and U7349 (N_7349,N_6613,N_6277);
and U7350 (N_7350,N_6316,N_6417);
or U7351 (N_7351,N_6299,N_6228);
nand U7352 (N_7352,N_6214,N_6643);
nor U7353 (N_7353,N_6591,N_6735);
nor U7354 (N_7354,N_6497,N_6214);
nor U7355 (N_7355,N_6365,N_6334);
or U7356 (N_7356,N_6511,N_6590);
or U7357 (N_7357,N_6422,N_6021);
or U7358 (N_7358,N_6534,N_6272);
or U7359 (N_7359,N_6387,N_6153);
or U7360 (N_7360,N_6580,N_6461);
xnor U7361 (N_7361,N_6590,N_6372);
and U7362 (N_7362,N_6278,N_6578);
or U7363 (N_7363,N_6142,N_6710);
or U7364 (N_7364,N_6535,N_6375);
or U7365 (N_7365,N_6061,N_6241);
nand U7366 (N_7366,N_6220,N_6302);
or U7367 (N_7367,N_6421,N_6119);
and U7368 (N_7368,N_6280,N_6573);
or U7369 (N_7369,N_6054,N_6389);
nor U7370 (N_7370,N_6552,N_6613);
nor U7371 (N_7371,N_6315,N_6486);
nor U7372 (N_7372,N_6530,N_6489);
nor U7373 (N_7373,N_6461,N_6318);
and U7374 (N_7374,N_6362,N_6683);
nor U7375 (N_7375,N_6705,N_6109);
or U7376 (N_7376,N_6292,N_6461);
and U7377 (N_7377,N_6300,N_6043);
nand U7378 (N_7378,N_6593,N_6636);
nand U7379 (N_7379,N_6690,N_6267);
nor U7380 (N_7380,N_6343,N_6427);
nand U7381 (N_7381,N_6124,N_6379);
or U7382 (N_7382,N_6328,N_6038);
nand U7383 (N_7383,N_6060,N_6633);
or U7384 (N_7384,N_6154,N_6183);
and U7385 (N_7385,N_6512,N_6384);
nand U7386 (N_7386,N_6520,N_6455);
or U7387 (N_7387,N_6721,N_6605);
or U7388 (N_7388,N_6284,N_6611);
and U7389 (N_7389,N_6585,N_6423);
nand U7390 (N_7390,N_6415,N_6146);
nand U7391 (N_7391,N_6073,N_6196);
nor U7392 (N_7392,N_6291,N_6450);
nand U7393 (N_7393,N_6585,N_6731);
and U7394 (N_7394,N_6697,N_6746);
and U7395 (N_7395,N_6237,N_6001);
and U7396 (N_7396,N_6399,N_6108);
nor U7397 (N_7397,N_6065,N_6147);
and U7398 (N_7398,N_6319,N_6217);
and U7399 (N_7399,N_6256,N_6268);
or U7400 (N_7400,N_6654,N_6582);
nor U7401 (N_7401,N_6617,N_6477);
nor U7402 (N_7402,N_6317,N_6736);
nand U7403 (N_7403,N_6554,N_6702);
or U7404 (N_7404,N_6574,N_6389);
or U7405 (N_7405,N_6294,N_6240);
nand U7406 (N_7406,N_6043,N_6076);
nand U7407 (N_7407,N_6247,N_6386);
or U7408 (N_7408,N_6459,N_6632);
nand U7409 (N_7409,N_6652,N_6142);
nand U7410 (N_7410,N_6731,N_6419);
nand U7411 (N_7411,N_6117,N_6123);
and U7412 (N_7412,N_6460,N_6567);
nand U7413 (N_7413,N_6689,N_6546);
nand U7414 (N_7414,N_6637,N_6583);
nor U7415 (N_7415,N_6675,N_6693);
nand U7416 (N_7416,N_6734,N_6693);
and U7417 (N_7417,N_6227,N_6011);
nand U7418 (N_7418,N_6255,N_6152);
nand U7419 (N_7419,N_6027,N_6232);
nand U7420 (N_7420,N_6498,N_6418);
nand U7421 (N_7421,N_6598,N_6017);
nor U7422 (N_7422,N_6052,N_6289);
and U7423 (N_7423,N_6051,N_6563);
or U7424 (N_7424,N_6195,N_6371);
nand U7425 (N_7425,N_6501,N_6070);
nor U7426 (N_7426,N_6424,N_6703);
nor U7427 (N_7427,N_6015,N_6447);
nor U7428 (N_7428,N_6283,N_6561);
and U7429 (N_7429,N_6299,N_6196);
or U7430 (N_7430,N_6432,N_6303);
nor U7431 (N_7431,N_6550,N_6304);
or U7432 (N_7432,N_6541,N_6172);
nand U7433 (N_7433,N_6267,N_6283);
nand U7434 (N_7434,N_6417,N_6270);
nor U7435 (N_7435,N_6398,N_6494);
or U7436 (N_7436,N_6100,N_6438);
nand U7437 (N_7437,N_6007,N_6037);
xnor U7438 (N_7438,N_6005,N_6332);
nand U7439 (N_7439,N_6475,N_6421);
and U7440 (N_7440,N_6529,N_6142);
and U7441 (N_7441,N_6707,N_6573);
or U7442 (N_7442,N_6658,N_6615);
nand U7443 (N_7443,N_6124,N_6140);
nor U7444 (N_7444,N_6584,N_6350);
nor U7445 (N_7445,N_6109,N_6053);
nand U7446 (N_7446,N_6708,N_6175);
or U7447 (N_7447,N_6681,N_6191);
nor U7448 (N_7448,N_6127,N_6116);
nor U7449 (N_7449,N_6147,N_6281);
nand U7450 (N_7450,N_6415,N_6531);
nand U7451 (N_7451,N_6023,N_6617);
or U7452 (N_7452,N_6573,N_6344);
nor U7453 (N_7453,N_6539,N_6717);
xnor U7454 (N_7454,N_6443,N_6408);
and U7455 (N_7455,N_6019,N_6383);
or U7456 (N_7456,N_6445,N_6190);
nand U7457 (N_7457,N_6103,N_6418);
and U7458 (N_7458,N_6074,N_6715);
and U7459 (N_7459,N_6166,N_6255);
nand U7460 (N_7460,N_6699,N_6011);
or U7461 (N_7461,N_6640,N_6081);
nor U7462 (N_7462,N_6335,N_6106);
or U7463 (N_7463,N_6036,N_6490);
or U7464 (N_7464,N_6227,N_6254);
nand U7465 (N_7465,N_6408,N_6095);
nand U7466 (N_7466,N_6588,N_6603);
and U7467 (N_7467,N_6609,N_6077);
and U7468 (N_7468,N_6556,N_6372);
nor U7469 (N_7469,N_6264,N_6272);
or U7470 (N_7470,N_6491,N_6444);
and U7471 (N_7471,N_6174,N_6398);
nand U7472 (N_7472,N_6100,N_6268);
nand U7473 (N_7473,N_6000,N_6017);
nand U7474 (N_7474,N_6109,N_6719);
nand U7475 (N_7475,N_6075,N_6483);
nand U7476 (N_7476,N_6086,N_6226);
and U7477 (N_7477,N_6489,N_6278);
or U7478 (N_7478,N_6470,N_6467);
nor U7479 (N_7479,N_6251,N_6719);
nand U7480 (N_7480,N_6063,N_6219);
or U7481 (N_7481,N_6338,N_6550);
nor U7482 (N_7482,N_6486,N_6461);
and U7483 (N_7483,N_6653,N_6574);
or U7484 (N_7484,N_6065,N_6100);
or U7485 (N_7485,N_6054,N_6197);
or U7486 (N_7486,N_6448,N_6378);
or U7487 (N_7487,N_6545,N_6559);
nor U7488 (N_7488,N_6708,N_6689);
and U7489 (N_7489,N_6163,N_6104);
or U7490 (N_7490,N_6565,N_6580);
nor U7491 (N_7491,N_6095,N_6024);
or U7492 (N_7492,N_6107,N_6005);
nor U7493 (N_7493,N_6008,N_6092);
or U7494 (N_7494,N_6269,N_6666);
xor U7495 (N_7495,N_6109,N_6172);
nor U7496 (N_7496,N_6089,N_6164);
and U7497 (N_7497,N_6387,N_6054);
nor U7498 (N_7498,N_6550,N_6602);
nor U7499 (N_7499,N_6081,N_6024);
nor U7500 (N_7500,N_7352,N_7481);
nand U7501 (N_7501,N_7019,N_7394);
or U7502 (N_7502,N_7034,N_7184);
xor U7503 (N_7503,N_6854,N_7053);
and U7504 (N_7504,N_6832,N_7334);
nor U7505 (N_7505,N_7423,N_7152);
or U7506 (N_7506,N_7122,N_7061);
nor U7507 (N_7507,N_7381,N_7302);
nor U7508 (N_7508,N_6821,N_7477);
or U7509 (N_7509,N_6971,N_6850);
and U7510 (N_7510,N_7223,N_7073);
nand U7511 (N_7511,N_6783,N_7375);
nor U7512 (N_7512,N_7157,N_6868);
nand U7513 (N_7513,N_6804,N_7487);
and U7514 (N_7514,N_7000,N_7208);
and U7515 (N_7515,N_6840,N_7028);
nor U7516 (N_7516,N_7046,N_6917);
or U7517 (N_7517,N_7438,N_7360);
or U7518 (N_7518,N_7368,N_6905);
or U7519 (N_7519,N_6772,N_7125);
and U7520 (N_7520,N_7175,N_6827);
and U7521 (N_7521,N_7387,N_7104);
nand U7522 (N_7522,N_7277,N_6959);
nand U7523 (N_7523,N_7221,N_6945);
nand U7524 (N_7524,N_7138,N_6752);
nor U7525 (N_7525,N_7301,N_7474);
and U7526 (N_7526,N_7244,N_6866);
or U7527 (N_7527,N_6870,N_7362);
nand U7528 (N_7528,N_7120,N_7101);
and U7529 (N_7529,N_7224,N_7432);
and U7530 (N_7530,N_7147,N_6873);
nand U7531 (N_7531,N_6967,N_7068);
nor U7532 (N_7532,N_7282,N_7412);
or U7533 (N_7533,N_6985,N_7317);
or U7534 (N_7534,N_7112,N_7306);
nor U7535 (N_7535,N_6876,N_6766);
and U7536 (N_7536,N_7022,N_7365);
or U7537 (N_7537,N_7257,N_7137);
and U7538 (N_7538,N_6970,N_7148);
or U7539 (N_7539,N_7009,N_6923);
nand U7540 (N_7540,N_6989,N_7176);
and U7541 (N_7541,N_6883,N_7256);
and U7542 (N_7542,N_7386,N_7410);
or U7543 (N_7543,N_7354,N_7070);
xnor U7544 (N_7544,N_7199,N_7107);
and U7545 (N_7545,N_6976,N_6913);
nand U7546 (N_7546,N_7151,N_7380);
xor U7547 (N_7547,N_7226,N_7027);
or U7548 (N_7548,N_7372,N_7088);
or U7549 (N_7549,N_6991,N_6891);
or U7550 (N_7550,N_7266,N_6920);
nand U7551 (N_7551,N_6927,N_6839);
nand U7552 (N_7552,N_7276,N_7333);
and U7553 (N_7553,N_6758,N_6911);
and U7554 (N_7554,N_6799,N_7461);
nor U7555 (N_7555,N_7204,N_7207);
nor U7556 (N_7556,N_7032,N_6784);
and U7557 (N_7557,N_6939,N_7210);
nor U7558 (N_7558,N_7076,N_7024);
or U7559 (N_7559,N_7241,N_7219);
and U7560 (N_7560,N_7469,N_6847);
and U7561 (N_7561,N_6879,N_6884);
nand U7562 (N_7562,N_7233,N_7440);
or U7563 (N_7563,N_7110,N_6836);
nor U7564 (N_7564,N_6788,N_7357);
or U7565 (N_7565,N_7012,N_6900);
and U7566 (N_7566,N_6816,N_7499);
and U7567 (N_7567,N_7332,N_6775);
nand U7568 (N_7568,N_7143,N_6830);
or U7569 (N_7569,N_7421,N_7154);
nor U7570 (N_7570,N_6929,N_6935);
nor U7571 (N_7571,N_7427,N_7265);
and U7572 (N_7572,N_7327,N_7488);
or U7573 (N_7573,N_7396,N_6793);
and U7574 (N_7574,N_7468,N_6969);
and U7575 (N_7575,N_7458,N_6898);
and U7576 (N_7576,N_6828,N_7038);
nand U7577 (N_7577,N_6776,N_7111);
or U7578 (N_7578,N_7393,N_7126);
or U7579 (N_7579,N_6755,N_7424);
nand U7580 (N_7580,N_7047,N_7344);
nand U7581 (N_7581,N_7132,N_6768);
nand U7582 (N_7582,N_6863,N_7462);
and U7583 (N_7583,N_7459,N_6994);
nor U7584 (N_7584,N_6813,N_7250);
or U7585 (N_7585,N_7338,N_6877);
nor U7586 (N_7586,N_6820,N_7051);
nand U7587 (N_7587,N_6983,N_7401);
nor U7588 (N_7588,N_7460,N_6947);
and U7589 (N_7589,N_7139,N_7081);
and U7590 (N_7590,N_7262,N_7272);
or U7591 (N_7591,N_7059,N_7379);
nor U7592 (N_7592,N_7418,N_6902);
or U7593 (N_7593,N_7407,N_7284);
nand U7594 (N_7594,N_7213,N_7229);
and U7595 (N_7595,N_7382,N_7405);
and U7596 (N_7596,N_6903,N_7491);
nor U7597 (N_7597,N_7194,N_7090);
nor U7598 (N_7598,N_7206,N_7473);
or U7599 (N_7599,N_6853,N_7013);
or U7600 (N_7600,N_7377,N_7337);
and U7601 (N_7601,N_7486,N_7039);
or U7602 (N_7602,N_6826,N_7245);
or U7603 (N_7603,N_7464,N_7158);
nand U7604 (N_7604,N_7323,N_6794);
nand U7605 (N_7605,N_7177,N_7066);
and U7606 (N_7606,N_7350,N_7355);
and U7607 (N_7607,N_7071,N_7456);
or U7608 (N_7608,N_6800,N_7325);
nor U7609 (N_7609,N_7005,N_6961);
nor U7610 (N_7610,N_6977,N_6882);
and U7611 (N_7611,N_6774,N_7397);
and U7612 (N_7612,N_7315,N_7050);
or U7613 (N_7613,N_7324,N_6978);
nand U7614 (N_7614,N_7293,N_7079);
nand U7615 (N_7615,N_6938,N_6823);
nor U7616 (N_7616,N_7170,N_6769);
nor U7617 (N_7617,N_7220,N_7471);
nor U7618 (N_7618,N_7114,N_7052);
nand U7619 (N_7619,N_7318,N_7239);
or U7620 (N_7620,N_7413,N_7203);
nand U7621 (N_7621,N_7135,N_7255);
and U7622 (N_7622,N_7014,N_7436);
nand U7623 (N_7623,N_6881,N_7341);
and U7624 (N_7624,N_7145,N_7298);
nand U7625 (N_7625,N_7231,N_6958);
nor U7626 (N_7626,N_7169,N_7096);
nor U7627 (N_7627,N_7197,N_7063);
xnor U7628 (N_7628,N_6846,N_6809);
nor U7629 (N_7629,N_7017,N_7236);
xor U7630 (N_7630,N_7035,N_7100);
and U7631 (N_7631,N_6915,N_6856);
nand U7632 (N_7632,N_7209,N_6932);
and U7633 (N_7633,N_6750,N_7055);
or U7634 (N_7634,N_6931,N_7041);
or U7635 (N_7635,N_7029,N_7190);
nor U7636 (N_7636,N_6950,N_7155);
or U7637 (N_7637,N_6965,N_7455);
and U7638 (N_7638,N_7191,N_7439);
or U7639 (N_7639,N_6770,N_6859);
nand U7640 (N_7640,N_6785,N_7275);
and U7641 (N_7641,N_6921,N_7165);
and U7642 (N_7642,N_7322,N_6764);
nand U7643 (N_7643,N_7217,N_6896);
or U7644 (N_7644,N_6999,N_6956);
or U7645 (N_7645,N_6963,N_7045);
nand U7646 (N_7646,N_7346,N_7215);
nand U7647 (N_7647,N_7127,N_6835);
and U7648 (N_7648,N_6778,N_7305);
nand U7649 (N_7649,N_6761,N_7105);
or U7650 (N_7650,N_7390,N_6937);
or U7651 (N_7651,N_7011,N_6781);
or U7652 (N_7652,N_7227,N_7482);
nand U7653 (N_7653,N_7330,N_6944);
or U7654 (N_7654,N_7278,N_7414);
or U7655 (N_7655,N_7251,N_7308);
or U7656 (N_7656,N_7367,N_7415);
nand U7657 (N_7657,N_6909,N_7263);
and U7658 (N_7658,N_7450,N_7311);
and U7659 (N_7659,N_7328,N_7296);
xor U7660 (N_7660,N_7335,N_7339);
and U7661 (N_7661,N_6875,N_7404);
nor U7662 (N_7662,N_6953,N_7358);
or U7663 (N_7663,N_7069,N_6998);
or U7664 (N_7664,N_7483,N_7159);
or U7665 (N_7665,N_7130,N_7202);
nand U7666 (N_7666,N_7168,N_6943);
or U7667 (N_7667,N_7285,N_7389);
or U7668 (N_7668,N_6845,N_7248);
or U7669 (N_7669,N_6771,N_7161);
xnor U7670 (N_7670,N_7188,N_6871);
or U7671 (N_7671,N_7102,N_7150);
and U7672 (N_7672,N_7467,N_7099);
and U7673 (N_7673,N_7270,N_6833);
nand U7674 (N_7674,N_7001,N_7428);
nand U7675 (N_7675,N_7097,N_6981);
or U7676 (N_7676,N_7268,N_7087);
xor U7677 (N_7677,N_6988,N_7292);
or U7678 (N_7678,N_6754,N_6806);
or U7679 (N_7679,N_7240,N_6791);
and U7680 (N_7680,N_7447,N_6808);
nor U7681 (N_7681,N_7426,N_7037);
and U7682 (N_7682,N_6810,N_7200);
and U7683 (N_7683,N_7319,N_6759);
nor U7684 (N_7684,N_7340,N_7373);
nand U7685 (N_7685,N_7134,N_7411);
and U7686 (N_7686,N_6760,N_7178);
or U7687 (N_7687,N_7273,N_7356);
and U7688 (N_7688,N_6992,N_6997);
and U7689 (N_7689,N_6777,N_7484);
or U7690 (N_7690,N_6841,N_7271);
nor U7691 (N_7691,N_7166,N_7383);
and U7692 (N_7692,N_7082,N_7092);
or U7693 (N_7693,N_7288,N_7205);
and U7694 (N_7694,N_6767,N_7406);
nor U7695 (N_7695,N_6897,N_6790);
nor U7696 (N_7696,N_6962,N_7131);
or U7697 (N_7697,N_6796,N_7181);
or U7698 (N_7698,N_6811,N_7472);
and U7699 (N_7699,N_7454,N_7281);
nor U7700 (N_7700,N_6893,N_7313);
and U7701 (N_7701,N_6795,N_7336);
nor U7702 (N_7702,N_6865,N_7289);
nor U7703 (N_7703,N_7149,N_6892);
and U7704 (N_7704,N_7212,N_7195);
and U7705 (N_7705,N_7291,N_6838);
nand U7706 (N_7706,N_7062,N_6818);
nand U7707 (N_7707,N_6812,N_7106);
nor U7708 (N_7708,N_6910,N_7253);
or U7709 (N_7709,N_6926,N_7025);
nand U7710 (N_7710,N_7093,N_7448);
nand U7711 (N_7711,N_6933,N_7043);
nor U7712 (N_7712,N_6878,N_7074);
nor U7713 (N_7713,N_6986,N_7048);
and U7714 (N_7714,N_7198,N_7264);
nor U7715 (N_7715,N_6973,N_6975);
nor U7716 (N_7716,N_6936,N_7123);
nand U7717 (N_7717,N_7441,N_7353);
nor U7718 (N_7718,N_6814,N_6894);
and U7719 (N_7719,N_6914,N_7067);
and U7720 (N_7720,N_7002,N_7077);
and U7721 (N_7721,N_6786,N_7031);
or U7722 (N_7722,N_6904,N_6889);
or U7723 (N_7723,N_7118,N_7321);
and U7724 (N_7724,N_7258,N_7044);
nand U7725 (N_7725,N_7167,N_6831);
nand U7726 (N_7726,N_7269,N_7451);
xor U7727 (N_7727,N_7314,N_7160);
nand U7728 (N_7728,N_7216,N_7442);
nand U7729 (N_7729,N_7449,N_7162);
nor U7730 (N_7730,N_7286,N_7156);
and U7731 (N_7731,N_7218,N_6844);
nand U7732 (N_7732,N_7098,N_6951);
or U7733 (N_7733,N_7008,N_6968);
and U7734 (N_7734,N_6890,N_6851);
nand U7735 (N_7735,N_7080,N_7054);
and U7736 (N_7736,N_7033,N_6887);
and U7737 (N_7737,N_7260,N_7299);
or U7738 (N_7738,N_7466,N_7128);
nand U7739 (N_7739,N_7417,N_7363);
nand U7740 (N_7740,N_7498,N_7247);
and U7741 (N_7741,N_7086,N_7084);
or U7742 (N_7742,N_7303,N_6919);
nand U7743 (N_7743,N_6980,N_6855);
nor U7744 (N_7744,N_7179,N_7429);
and U7745 (N_7745,N_6797,N_7189);
nand U7746 (N_7746,N_6906,N_7230);
nor U7747 (N_7747,N_6798,N_7402);
and U7748 (N_7748,N_7153,N_7476);
nand U7749 (N_7749,N_7295,N_7446);
nand U7750 (N_7750,N_7225,N_6972);
and U7751 (N_7751,N_6848,N_6773);
and U7752 (N_7752,N_6780,N_6957);
nor U7753 (N_7753,N_7117,N_6955);
or U7754 (N_7754,N_6817,N_7274);
nand U7755 (N_7755,N_7312,N_7408);
nor U7756 (N_7756,N_7015,N_6907);
or U7757 (N_7757,N_6899,N_7091);
nand U7758 (N_7758,N_7343,N_7246);
or U7759 (N_7759,N_6888,N_7495);
xnor U7760 (N_7760,N_7463,N_6843);
and U7761 (N_7761,N_7173,N_7108);
or U7762 (N_7762,N_7211,N_7234);
and U7763 (N_7763,N_7297,N_7261);
or U7764 (N_7764,N_7078,N_6842);
and U7765 (N_7765,N_6872,N_6805);
and U7766 (N_7766,N_7388,N_6979);
and U7767 (N_7767,N_7437,N_7490);
or U7768 (N_7768,N_6852,N_7119);
nor U7769 (N_7769,N_7243,N_6996);
or U7770 (N_7770,N_6787,N_7434);
nor U7771 (N_7771,N_7366,N_7349);
or U7772 (N_7772,N_7452,N_6869);
or U7773 (N_7773,N_7416,N_7026);
or U7774 (N_7774,N_6885,N_7058);
nand U7775 (N_7775,N_7196,N_7403);
or U7776 (N_7776,N_7140,N_7222);
nand U7777 (N_7777,N_7494,N_6765);
or U7778 (N_7778,N_7249,N_7385);
nand U7779 (N_7779,N_7420,N_7201);
and U7780 (N_7780,N_6837,N_7129);
nand U7781 (N_7781,N_7470,N_7398);
or U7782 (N_7782,N_7287,N_7391);
and U7783 (N_7783,N_7395,N_7095);
nand U7784 (N_7784,N_7182,N_6862);
nand U7785 (N_7785,N_7345,N_7040);
or U7786 (N_7786,N_6922,N_7072);
nand U7787 (N_7787,N_6949,N_7443);
nand U7788 (N_7788,N_6960,N_7023);
xnor U7789 (N_7789,N_6895,N_7478);
xor U7790 (N_7790,N_7364,N_6815);
or U7791 (N_7791,N_7259,N_6982);
or U7792 (N_7792,N_7103,N_7444);
nor U7793 (N_7793,N_6930,N_7171);
nand U7794 (N_7794,N_7307,N_7348);
or U7795 (N_7795,N_7018,N_6858);
or U7796 (N_7796,N_7267,N_6987);
nand U7797 (N_7797,N_6952,N_7400);
nand U7798 (N_7798,N_7290,N_7228);
and U7799 (N_7799,N_7174,N_7238);
nor U7800 (N_7800,N_6912,N_7342);
nand U7801 (N_7801,N_7370,N_7020);
nand U7802 (N_7802,N_7431,N_7142);
nand U7803 (N_7803,N_6918,N_7331);
and U7804 (N_7804,N_6886,N_7232);
and U7805 (N_7805,N_7146,N_7042);
nand U7806 (N_7806,N_7083,N_7280);
xor U7807 (N_7807,N_7049,N_7185);
nand U7808 (N_7808,N_6867,N_7214);
nor U7809 (N_7809,N_7254,N_7183);
nor U7810 (N_7810,N_7193,N_7309);
and U7811 (N_7811,N_6941,N_7113);
and U7812 (N_7812,N_7252,N_7430);
and U7813 (N_7813,N_6934,N_6802);
or U7814 (N_7814,N_7384,N_7116);
nor U7815 (N_7815,N_7347,N_7021);
and U7816 (N_7816,N_6948,N_7057);
nand U7817 (N_7817,N_7359,N_7453);
or U7818 (N_7818,N_7310,N_7361);
or U7819 (N_7819,N_7485,N_6928);
nand U7820 (N_7820,N_7326,N_6751);
nor U7821 (N_7821,N_6940,N_6901);
nor U7822 (N_7822,N_7056,N_7489);
nor U7823 (N_7823,N_7124,N_7492);
and U7824 (N_7824,N_7186,N_7399);
or U7825 (N_7825,N_6782,N_6864);
nand U7826 (N_7826,N_7065,N_7465);
or U7827 (N_7827,N_6874,N_6925);
nor U7828 (N_7828,N_7016,N_7320);
xnor U7829 (N_7829,N_7409,N_7294);
or U7830 (N_7830,N_6753,N_6789);
and U7831 (N_7831,N_7006,N_7004);
nor U7832 (N_7832,N_7094,N_7136);
nand U7833 (N_7833,N_7392,N_7164);
or U7834 (N_7834,N_7479,N_7374);
and U7835 (N_7835,N_7457,N_6974);
or U7836 (N_7836,N_6762,N_7237);
or U7837 (N_7837,N_6763,N_7187);
and U7838 (N_7838,N_7003,N_6807);
or U7839 (N_7839,N_7064,N_7007);
and U7840 (N_7840,N_6803,N_6860);
nor U7841 (N_7841,N_7141,N_7144);
nand U7842 (N_7842,N_7304,N_7422);
or U7843 (N_7843,N_7376,N_6990);
nor U7844 (N_7844,N_7279,N_7030);
and U7845 (N_7845,N_6779,N_7172);
nor U7846 (N_7846,N_7163,N_7475);
and U7847 (N_7847,N_7378,N_6954);
and U7848 (N_7848,N_7075,N_7351);
or U7849 (N_7849,N_6822,N_6824);
and U7850 (N_7850,N_7316,N_6942);
or U7851 (N_7851,N_7010,N_7300);
xnor U7852 (N_7852,N_6819,N_7445);
nor U7853 (N_7853,N_6792,N_6801);
or U7854 (N_7854,N_6861,N_7371);
and U7855 (N_7855,N_6995,N_6857);
and U7856 (N_7856,N_7115,N_7133);
nor U7857 (N_7857,N_7480,N_7085);
and U7858 (N_7858,N_7060,N_7369);
or U7859 (N_7859,N_7235,N_7493);
or U7860 (N_7860,N_7036,N_6964);
xnor U7861 (N_7861,N_6829,N_6825);
or U7862 (N_7862,N_7425,N_7435);
and U7863 (N_7863,N_7497,N_7433);
and U7864 (N_7864,N_6880,N_6993);
or U7865 (N_7865,N_6908,N_6757);
and U7866 (N_7866,N_6984,N_7121);
and U7867 (N_7867,N_7283,N_7242);
nand U7868 (N_7868,N_7419,N_6834);
and U7869 (N_7869,N_6966,N_6756);
nand U7870 (N_7870,N_7109,N_7180);
nand U7871 (N_7871,N_7496,N_6946);
nand U7872 (N_7872,N_7329,N_6916);
nand U7873 (N_7873,N_7192,N_6849);
nor U7874 (N_7874,N_7089,N_6924);
nor U7875 (N_7875,N_6822,N_7075);
or U7876 (N_7876,N_6764,N_7167);
nand U7877 (N_7877,N_7021,N_6952);
and U7878 (N_7878,N_7127,N_6774);
nand U7879 (N_7879,N_7395,N_7462);
or U7880 (N_7880,N_6942,N_6817);
nor U7881 (N_7881,N_7227,N_6863);
or U7882 (N_7882,N_6943,N_6797);
and U7883 (N_7883,N_6760,N_6908);
and U7884 (N_7884,N_7299,N_7182);
and U7885 (N_7885,N_6922,N_7462);
and U7886 (N_7886,N_7112,N_7063);
or U7887 (N_7887,N_6929,N_7045);
nor U7888 (N_7888,N_7103,N_7216);
nand U7889 (N_7889,N_7462,N_7235);
and U7890 (N_7890,N_6990,N_7308);
and U7891 (N_7891,N_7335,N_7477);
or U7892 (N_7892,N_6822,N_6752);
and U7893 (N_7893,N_7149,N_7236);
nor U7894 (N_7894,N_6924,N_6848);
nor U7895 (N_7895,N_7148,N_7172);
nand U7896 (N_7896,N_7463,N_6782);
nand U7897 (N_7897,N_7428,N_6896);
or U7898 (N_7898,N_7471,N_7318);
or U7899 (N_7899,N_7047,N_7496);
or U7900 (N_7900,N_7324,N_6896);
nor U7901 (N_7901,N_7272,N_6993);
nor U7902 (N_7902,N_7473,N_6943);
nor U7903 (N_7903,N_7289,N_7491);
nor U7904 (N_7904,N_7457,N_6885);
nor U7905 (N_7905,N_6986,N_7097);
nor U7906 (N_7906,N_6893,N_7032);
or U7907 (N_7907,N_6796,N_7454);
nor U7908 (N_7908,N_7172,N_7131);
or U7909 (N_7909,N_6791,N_7451);
nand U7910 (N_7910,N_7271,N_7032);
nor U7911 (N_7911,N_7069,N_7467);
and U7912 (N_7912,N_6960,N_7268);
nand U7913 (N_7913,N_7128,N_6903);
or U7914 (N_7914,N_6857,N_7109);
nand U7915 (N_7915,N_7020,N_7050);
nand U7916 (N_7916,N_7060,N_7473);
nor U7917 (N_7917,N_6883,N_6889);
and U7918 (N_7918,N_7301,N_7249);
and U7919 (N_7919,N_7013,N_7302);
nor U7920 (N_7920,N_7373,N_6783);
nor U7921 (N_7921,N_7288,N_6923);
nand U7922 (N_7922,N_6976,N_7043);
or U7923 (N_7923,N_6850,N_6878);
or U7924 (N_7924,N_6953,N_7373);
and U7925 (N_7925,N_7092,N_7498);
or U7926 (N_7926,N_7040,N_7373);
nand U7927 (N_7927,N_7313,N_7088);
and U7928 (N_7928,N_7272,N_7399);
and U7929 (N_7929,N_7111,N_6759);
and U7930 (N_7930,N_6901,N_7323);
nor U7931 (N_7931,N_7158,N_7037);
or U7932 (N_7932,N_7147,N_6863);
and U7933 (N_7933,N_7368,N_7101);
or U7934 (N_7934,N_7172,N_6951);
and U7935 (N_7935,N_7057,N_6943);
or U7936 (N_7936,N_7048,N_6946);
nor U7937 (N_7937,N_6963,N_6788);
nand U7938 (N_7938,N_6855,N_7156);
nor U7939 (N_7939,N_6809,N_7348);
nand U7940 (N_7940,N_6831,N_7166);
nand U7941 (N_7941,N_7126,N_7489);
or U7942 (N_7942,N_6986,N_7293);
or U7943 (N_7943,N_6970,N_6968);
and U7944 (N_7944,N_7297,N_7418);
nand U7945 (N_7945,N_7069,N_7267);
or U7946 (N_7946,N_7449,N_7474);
and U7947 (N_7947,N_7432,N_6821);
and U7948 (N_7948,N_7037,N_6970);
nor U7949 (N_7949,N_6953,N_7307);
nor U7950 (N_7950,N_7498,N_6824);
and U7951 (N_7951,N_7318,N_6977);
nand U7952 (N_7952,N_7328,N_7048);
and U7953 (N_7953,N_7329,N_7149);
nand U7954 (N_7954,N_7082,N_6858);
nand U7955 (N_7955,N_7067,N_7195);
and U7956 (N_7956,N_6870,N_6794);
and U7957 (N_7957,N_7015,N_7089);
nor U7958 (N_7958,N_7412,N_7403);
nand U7959 (N_7959,N_7383,N_6773);
nor U7960 (N_7960,N_7459,N_7016);
or U7961 (N_7961,N_6878,N_7263);
and U7962 (N_7962,N_7135,N_6788);
or U7963 (N_7963,N_7050,N_7239);
and U7964 (N_7964,N_6887,N_6923);
nor U7965 (N_7965,N_6863,N_6786);
nand U7966 (N_7966,N_7407,N_7242);
or U7967 (N_7967,N_6922,N_7169);
or U7968 (N_7968,N_7347,N_7239);
nand U7969 (N_7969,N_7440,N_6982);
nand U7970 (N_7970,N_7129,N_6886);
nand U7971 (N_7971,N_7163,N_7030);
nor U7972 (N_7972,N_6824,N_6787);
nand U7973 (N_7973,N_7495,N_7399);
and U7974 (N_7974,N_7091,N_6871);
nand U7975 (N_7975,N_7049,N_6790);
nand U7976 (N_7976,N_7038,N_7159);
and U7977 (N_7977,N_7036,N_6881);
and U7978 (N_7978,N_7469,N_7390);
and U7979 (N_7979,N_6857,N_7093);
nand U7980 (N_7980,N_7343,N_6897);
or U7981 (N_7981,N_7336,N_6976);
and U7982 (N_7982,N_6890,N_7446);
and U7983 (N_7983,N_7085,N_7440);
and U7984 (N_7984,N_6857,N_6870);
nor U7985 (N_7985,N_6895,N_6783);
nor U7986 (N_7986,N_7068,N_7268);
and U7987 (N_7987,N_7468,N_7262);
nand U7988 (N_7988,N_7260,N_7490);
and U7989 (N_7989,N_6882,N_7011);
nor U7990 (N_7990,N_6830,N_6901);
or U7991 (N_7991,N_7259,N_6790);
nor U7992 (N_7992,N_6805,N_6865);
and U7993 (N_7993,N_7134,N_6875);
and U7994 (N_7994,N_7277,N_7339);
and U7995 (N_7995,N_7055,N_7345);
and U7996 (N_7996,N_7220,N_7391);
or U7997 (N_7997,N_7320,N_7082);
nor U7998 (N_7998,N_7275,N_7388);
nand U7999 (N_7999,N_6766,N_7387);
or U8000 (N_8000,N_6994,N_6926);
or U8001 (N_8001,N_7377,N_7264);
nand U8002 (N_8002,N_7243,N_6887);
nor U8003 (N_8003,N_6949,N_7189);
or U8004 (N_8004,N_7462,N_7480);
and U8005 (N_8005,N_7149,N_7327);
nor U8006 (N_8006,N_6841,N_7441);
and U8007 (N_8007,N_7051,N_7366);
nand U8008 (N_8008,N_7364,N_6795);
and U8009 (N_8009,N_7328,N_6859);
or U8010 (N_8010,N_6961,N_6876);
or U8011 (N_8011,N_7135,N_7490);
nor U8012 (N_8012,N_7184,N_7447);
xnor U8013 (N_8013,N_7233,N_7014);
nor U8014 (N_8014,N_7089,N_7365);
nand U8015 (N_8015,N_7088,N_7415);
or U8016 (N_8016,N_7145,N_6950);
nand U8017 (N_8017,N_7388,N_6859);
nand U8018 (N_8018,N_7409,N_7139);
nor U8019 (N_8019,N_6797,N_7004);
and U8020 (N_8020,N_7399,N_7045);
nand U8021 (N_8021,N_7259,N_6793);
or U8022 (N_8022,N_7352,N_7289);
and U8023 (N_8023,N_7175,N_6907);
nor U8024 (N_8024,N_6866,N_6924);
or U8025 (N_8025,N_7046,N_7096);
and U8026 (N_8026,N_7484,N_7049);
and U8027 (N_8027,N_7474,N_6885);
and U8028 (N_8028,N_6945,N_6880);
nor U8029 (N_8029,N_7417,N_7183);
and U8030 (N_8030,N_6902,N_7161);
nand U8031 (N_8031,N_6986,N_6927);
and U8032 (N_8032,N_7463,N_7175);
or U8033 (N_8033,N_7452,N_7300);
nand U8034 (N_8034,N_7420,N_7299);
nand U8035 (N_8035,N_7057,N_7385);
and U8036 (N_8036,N_7169,N_7210);
and U8037 (N_8037,N_6803,N_6761);
nor U8038 (N_8038,N_6957,N_7193);
nor U8039 (N_8039,N_7117,N_7478);
and U8040 (N_8040,N_6787,N_6998);
xor U8041 (N_8041,N_7055,N_7318);
nor U8042 (N_8042,N_6787,N_6844);
and U8043 (N_8043,N_6863,N_6994);
or U8044 (N_8044,N_7422,N_6760);
or U8045 (N_8045,N_7279,N_6993);
nand U8046 (N_8046,N_7350,N_7320);
or U8047 (N_8047,N_6993,N_6807);
or U8048 (N_8048,N_7121,N_7091);
nand U8049 (N_8049,N_6828,N_7057);
and U8050 (N_8050,N_7300,N_7313);
and U8051 (N_8051,N_7452,N_6939);
nand U8052 (N_8052,N_7456,N_7337);
and U8053 (N_8053,N_7255,N_7394);
or U8054 (N_8054,N_6875,N_7120);
nor U8055 (N_8055,N_7118,N_6957);
nor U8056 (N_8056,N_7008,N_6957);
or U8057 (N_8057,N_6767,N_7453);
nand U8058 (N_8058,N_6870,N_7210);
nand U8059 (N_8059,N_6795,N_6972);
nand U8060 (N_8060,N_7290,N_7074);
nand U8061 (N_8061,N_7423,N_7466);
nand U8062 (N_8062,N_7484,N_7114);
and U8063 (N_8063,N_7183,N_7466);
or U8064 (N_8064,N_6984,N_7299);
or U8065 (N_8065,N_7018,N_7176);
nand U8066 (N_8066,N_7371,N_6962);
nand U8067 (N_8067,N_7327,N_7101);
nand U8068 (N_8068,N_7064,N_6829);
nor U8069 (N_8069,N_7154,N_7184);
nor U8070 (N_8070,N_7336,N_6934);
nor U8071 (N_8071,N_7072,N_7081);
or U8072 (N_8072,N_7345,N_6892);
or U8073 (N_8073,N_7036,N_7162);
and U8074 (N_8074,N_7150,N_7218);
nor U8075 (N_8075,N_6769,N_6757);
nor U8076 (N_8076,N_7210,N_7284);
nand U8077 (N_8077,N_6804,N_7364);
nor U8078 (N_8078,N_7185,N_7184);
and U8079 (N_8079,N_7084,N_7307);
and U8080 (N_8080,N_7052,N_6765);
and U8081 (N_8081,N_6762,N_6983);
and U8082 (N_8082,N_6863,N_7132);
nand U8083 (N_8083,N_6832,N_6940);
nor U8084 (N_8084,N_6813,N_6766);
or U8085 (N_8085,N_7179,N_7486);
or U8086 (N_8086,N_6777,N_6811);
nand U8087 (N_8087,N_7220,N_7276);
nor U8088 (N_8088,N_7193,N_6984);
and U8089 (N_8089,N_6949,N_7145);
and U8090 (N_8090,N_7462,N_7473);
or U8091 (N_8091,N_6776,N_6877);
and U8092 (N_8092,N_7221,N_7454);
nor U8093 (N_8093,N_7131,N_7205);
nand U8094 (N_8094,N_7461,N_7255);
nor U8095 (N_8095,N_6870,N_7159);
and U8096 (N_8096,N_7182,N_7265);
and U8097 (N_8097,N_7356,N_6887);
and U8098 (N_8098,N_7273,N_7442);
nand U8099 (N_8099,N_7320,N_7402);
nor U8100 (N_8100,N_6843,N_7473);
or U8101 (N_8101,N_6916,N_6778);
nand U8102 (N_8102,N_7074,N_7379);
or U8103 (N_8103,N_6809,N_7499);
and U8104 (N_8104,N_6896,N_7418);
nor U8105 (N_8105,N_6997,N_7472);
nand U8106 (N_8106,N_7077,N_7383);
nor U8107 (N_8107,N_7386,N_7448);
or U8108 (N_8108,N_6771,N_7196);
nor U8109 (N_8109,N_7193,N_7457);
or U8110 (N_8110,N_7075,N_6768);
nand U8111 (N_8111,N_7116,N_7010);
or U8112 (N_8112,N_7095,N_7233);
and U8113 (N_8113,N_7163,N_7197);
nand U8114 (N_8114,N_6914,N_7374);
and U8115 (N_8115,N_7245,N_7107);
and U8116 (N_8116,N_6791,N_6821);
nor U8117 (N_8117,N_7127,N_6967);
or U8118 (N_8118,N_7257,N_7465);
or U8119 (N_8119,N_7221,N_7116);
nor U8120 (N_8120,N_6824,N_6826);
nand U8121 (N_8121,N_6819,N_7256);
nor U8122 (N_8122,N_7406,N_7424);
nor U8123 (N_8123,N_7408,N_7102);
and U8124 (N_8124,N_7343,N_7161);
or U8125 (N_8125,N_7141,N_6772);
nor U8126 (N_8126,N_7182,N_6767);
and U8127 (N_8127,N_6860,N_6993);
or U8128 (N_8128,N_6950,N_6885);
nor U8129 (N_8129,N_7077,N_7385);
nor U8130 (N_8130,N_6826,N_7065);
nor U8131 (N_8131,N_7431,N_6845);
and U8132 (N_8132,N_7022,N_7008);
or U8133 (N_8133,N_6985,N_7219);
or U8134 (N_8134,N_6993,N_7141);
nand U8135 (N_8135,N_7077,N_6975);
nor U8136 (N_8136,N_7119,N_6838);
and U8137 (N_8137,N_6986,N_7444);
and U8138 (N_8138,N_7117,N_7169);
or U8139 (N_8139,N_6796,N_7120);
nand U8140 (N_8140,N_7175,N_7119);
and U8141 (N_8141,N_7265,N_7121);
nand U8142 (N_8142,N_6901,N_7322);
nand U8143 (N_8143,N_7073,N_7429);
nor U8144 (N_8144,N_7470,N_7044);
xor U8145 (N_8145,N_7355,N_6870);
nand U8146 (N_8146,N_7080,N_7078);
and U8147 (N_8147,N_6783,N_7361);
or U8148 (N_8148,N_7477,N_7349);
nand U8149 (N_8149,N_7035,N_7496);
nor U8150 (N_8150,N_7446,N_7045);
nand U8151 (N_8151,N_7042,N_6915);
nor U8152 (N_8152,N_7159,N_7330);
or U8153 (N_8153,N_6946,N_6845);
nand U8154 (N_8154,N_6900,N_7373);
nand U8155 (N_8155,N_6751,N_7397);
nor U8156 (N_8156,N_7073,N_7204);
and U8157 (N_8157,N_7423,N_7059);
or U8158 (N_8158,N_6986,N_7098);
nor U8159 (N_8159,N_7248,N_7218);
and U8160 (N_8160,N_7077,N_6859);
or U8161 (N_8161,N_7318,N_7340);
nor U8162 (N_8162,N_6951,N_6997);
nor U8163 (N_8163,N_6813,N_7437);
nand U8164 (N_8164,N_7022,N_7458);
and U8165 (N_8165,N_7370,N_7262);
nor U8166 (N_8166,N_7264,N_7060);
and U8167 (N_8167,N_6751,N_7285);
or U8168 (N_8168,N_7418,N_7359);
nor U8169 (N_8169,N_6868,N_6785);
nor U8170 (N_8170,N_7347,N_7319);
and U8171 (N_8171,N_6883,N_7399);
and U8172 (N_8172,N_7031,N_7034);
and U8173 (N_8173,N_6868,N_6931);
and U8174 (N_8174,N_6804,N_6863);
nor U8175 (N_8175,N_6820,N_6779);
or U8176 (N_8176,N_7383,N_6905);
nor U8177 (N_8177,N_7356,N_7188);
nor U8178 (N_8178,N_7121,N_7440);
or U8179 (N_8179,N_6854,N_7196);
and U8180 (N_8180,N_7103,N_7028);
nor U8181 (N_8181,N_7265,N_7282);
and U8182 (N_8182,N_6766,N_7311);
or U8183 (N_8183,N_7463,N_6914);
nand U8184 (N_8184,N_7383,N_6995);
and U8185 (N_8185,N_7073,N_7349);
or U8186 (N_8186,N_7314,N_7287);
and U8187 (N_8187,N_7270,N_7493);
nand U8188 (N_8188,N_7390,N_6800);
and U8189 (N_8189,N_7266,N_7079);
nand U8190 (N_8190,N_6865,N_7096);
nor U8191 (N_8191,N_6971,N_7204);
or U8192 (N_8192,N_7029,N_6883);
nor U8193 (N_8193,N_7035,N_6935);
and U8194 (N_8194,N_7176,N_6753);
nand U8195 (N_8195,N_7056,N_6970);
or U8196 (N_8196,N_7130,N_7194);
and U8197 (N_8197,N_7429,N_6946);
or U8198 (N_8198,N_7099,N_7144);
nand U8199 (N_8199,N_7139,N_7462);
nand U8200 (N_8200,N_6885,N_7196);
or U8201 (N_8201,N_6926,N_7207);
nand U8202 (N_8202,N_6772,N_7349);
nand U8203 (N_8203,N_7244,N_7422);
nand U8204 (N_8204,N_7254,N_7344);
and U8205 (N_8205,N_7020,N_7108);
nor U8206 (N_8206,N_6780,N_7185);
and U8207 (N_8207,N_7320,N_7318);
and U8208 (N_8208,N_6817,N_7309);
nand U8209 (N_8209,N_6883,N_7460);
nor U8210 (N_8210,N_6928,N_6805);
nand U8211 (N_8211,N_7176,N_7059);
or U8212 (N_8212,N_6837,N_7360);
or U8213 (N_8213,N_7267,N_7038);
and U8214 (N_8214,N_6992,N_6880);
nor U8215 (N_8215,N_7305,N_7388);
and U8216 (N_8216,N_6989,N_6931);
or U8217 (N_8217,N_7416,N_7490);
and U8218 (N_8218,N_7014,N_7030);
nand U8219 (N_8219,N_6863,N_7167);
nor U8220 (N_8220,N_7468,N_7142);
and U8221 (N_8221,N_7242,N_7394);
or U8222 (N_8222,N_6911,N_6780);
or U8223 (N_8223,N_7062,N_7356);
nand U8224 (N_8224,N_6817,N_6902);
nand U8225 (N_8225,N_6879,N_7107);
nand U8226 (N_8226,N_7210,N_7090);
nor U8227 (N_8227,N_7089,N_7255);
nand U8228 (N_8228,N_7098,N_7343);
nor U8229 (N_8229,N_7404,N_6853);
and U8230 (N_8230,N_6975,N_6818);
or U8231 (N_8231,N_6770,N_7204);
and U8232 (N_8232,N_6858,N_6808);
nand U8233 (N_8233,N_6998,N_7454);
nand U8234 (N_8234,N_7131,N_7246);
or U8235 (N_8235,N_7468,N_7058);
nor U8236 (N_8236,N_7338,N_7374);
nor U8237 (N_8237,N_7132,N_6857);
or U8238 (N_8238,N_6822,N_7286);
nand U8239 (N_8239,N_7048,N_7491);
or U8240 (N_8240,N_6865,N_7462);
nor U8241 (N_8241,N_7028,N_6893);
and U8242 (N_8242,N_6807,N_7181);
and U8243 (N_8243,N_6838,N_6903);
nor U8244 (N_8244,N_7458,N_7187);
and U8245 (N_8245,N_7293,N_7435);
nand U8246 (N_8246,N_6813,N_7492);
and U8247 (N_8247,N_6854,N_6984);
nand U8248 (N_8248,N_6778,N_7438);
nor U8249 (N_8249,N_6765,N_7429);
nor U8250 (N_8250,N_7910,N_7996);
nor U8251 (N_8251,N_7587,N_7824);
and U8252 (N_8252,N_8139,N_7892);
nand U8253 (N_8253,N_7985,N_7907);
xor U8254 (N_8254,N_7671,N_7518);
and U8255 (N_8255,N_7780,N_7505);
nand U8256 (N_8256,N_7622,N_7632);
or U8257 (N_8257,N_7995,N_8148);
nand U8258 (N_8258,N_8112,N_7576);
nand U8259 (N_8259,N_7945,N_8171);
nor U8260 (N_8260,N_7772,N_8189);
and U8261 (N_8261,N_7618,N_7514);
or U8262 (N_8262,N_8046,N_7957);
and U8263 (N_8263,N_7666,N_7800);
nor U8264 (N_8264,N_7675,N_7938);
and U8265 (N_8265,N_7887,N_7943);
or U8266 (N_8266,N_7695,N_7717);
nand U8267 (N_8267,N_8236,N_7734);
and U8268 (N_8268,N_7791,N_8237);
and U8269 (N_8269,N_7762,N_8161);
or U8270 (N_8270,N_8122,N_7889);
nand U8271 (N_8271,N_8177,N_7561);
nor U8272 (N_8272,N_7819,N_8095);
nand U8273 (N_8273,N_7669,N_7774);
nand U8274 (N_8274,N_8009,N_7592);
and U8275 (N_8275,N_8100,N_8153);
and U8276 (N_8276,N_8016,N_7535);
and U8277 (N_8277,N_8173,N_8049);
or U8278 (N_8278,N_7962,N_7710);
or U8279 (N_8279,N_7882,N_7832);
and U8280 (N_8280,N_8005,N_7683);
nand U8281 (N_8281,N_8142,N_7768);
and U8282 (N_8282,N_7950,N_8132);
nand U8283 (N_8283,N_7944,N_7672);
nor U8284 (N_8284,N_7853,N_7743);
and U8285 (N_8285,N_7828,N_8052);
nor U8286 (N_8286,N_7639,N_7811);
or U8287 (N_8287,N_7593,N_7658);
and U8288 (N_8288,N_8225,N_7504);
and U8289 (N_8289,N_7647,N_7611);
or U8290 (N_8290,N_7829,N_7685);
and U8291 (N_8291,N_7720,N_8240);
nand U8292 (N_8292,N_8223,N_7788);
nor U8293 (N_8293,N_7822,N_7506);
nor U8294 (N_8294,N_7702,N_7871);
or U8295 (N_8295,N_8040,N_7886);
nor U8296 (N_8296,N_8013,N_8056);
xnor U8297 (N_8297,N_7787,N_8008);
and U8298 (N_8298,N_7815,N_8012);
or U8299 (N_8299,N_7911,N_7559);
and U8300 (N_8300,N_8118,N_8160);
nor U8301 (N_8301,N_8107,N_7827);
nor U8302 (N_8302,N_7713,N_7967);
nand U8303 (N_8303,N_7877,N_8214);
and U8304 (N_8304,N_8217,N_7503);
nand U8305 (N_8305,N_7992,N_7607);
and U8306 (N_8306,N_8154,N_7541);
nor U8307 (N_8307,N_7784,N_8034);
nand U8308 (N_8308,N_8080,N_7854);
nand U8309 (N_8309,N_7746,N_7567);
or U8310 (N_8310,N_7530,N_7513);
or U8311 (N_8311,N_8014,N_8226);
nand U8312 (N_8312,N_8128,N_7659);
or U8313 (N_8313,N_7723,N_8174);
and U8314 (N_8314,N_7670,N_7821);
or U8315 (N_8315,N_7715,N_7709);
nand U8316 (N_8316,N_7764,N_7864);
or U8317 (N_8317,N_8001,N_8033);
and U8318 (N_8318,N_7726,N_7583);
or U8319 (N_8319,N_7874,N_7582);
nor U8320 (N_8320,N_8141,N_7870);
or U8321 (N_8321,N_8007,N_7668);
nor U8322 (N_8322,N_7727,N_7729);
and U8323 (N_8323,N_7794,N_8233);
nand U8324 (N_8324,N_7554,N_8029);
or U8325 (N_8325,N_8028,N_7572);
nand U8326 (N_8326,N_8098,N_7722);
or U8327 (N_8327,N_8144,N_8091);
or U8328 (N_8328,N_8081,N_7916);
nand U8329 (N_8329,N_8094,N_7703);
and U8330 (N_8330,N_7537,N_7981);
or U8331 (N_8331,N_7711,N_7744);
nor U8332 (N_8332,N_7975,N_8243);
nand U8333 (N_8333,N_7799,N_7553);
and U8334 (N_8334,N_8193,N_7570);
and U8335 (N_8335,N_8065,N_7620);
nand U8336 (N_8336,N_8210,N_8136);
nor U8337 (N_8337,N_8245,N_7516);
nor U8338 (N_8338,N_8050,N_8242);
nand U8339 (N_8339,N_7617,N_7951);
nand U8340 (N_8340,N_8010,N_8131);
or U8341 (N_8341,N_7804,N_7507);
nand U8342 (N_8342,N_7803,N_8085);
and U8343 (N_8343,N_8190,N_7602);
or U8344 (N_8344,N_7801,N_7624);
or U8345 (N_8345,N_8146,N_7777);
or U8346 (N_8346,N_8194,N_8077);
nand U8347 (N_8347,N_7594,N_7972);
nand U8348 (N_8348,N_7646,N_8062);
and U8349 (N_8349,N_7830,N_7562);
nand U8350 (N_8350,N_7919,N_7939);
and U8351 (N_8351,N_7536,N_7937);
and U8352 (N_8352,N_7529,N_7616);
and U8353 (N_8353,N_7866,N_7663);
or U8354 (N_8354,N_7809,N_7716);
nor U8355 (N_8355,N_7748,N_8045);
nor U8356 (N_8356,N_7896,N_7705);
nor U8357 (N_8357,N_8063,N_8069);
nor U8358 (N_8358,N_8249,N_8022);
nor U8359 (N_8359,N_8156,N_7863);
nand U8360 (N_8360,N_7608,N_7795);
and U8361 (N_8361,N_7545,N_8057);
and U8362 (N_8362,N_7501,N_7812);
or U8363 (N_8363,N_7750,N_7598);
nand U8364 (N_8364,N_8076,N_7596);
nor U8365 (N_8365,N_8186,N_7868);
or U8366 (N_8366,N_7857,N_7927);
nor U8367 (N_8367,N_7793,N_7802);
or U8368 (N_8368,N_7818,N_7942);
nand U8369 (N_8369,N_7925,N_8149);
or U8370 (N_8370,N_7585,N_8015);
or U8371 (N_8371,N_7767,N_7875);
nor U8372 (N_8372,N_7783,N_7965);
nand U8373 (N_8373,N_8230,N_8157);
and U8374 (N_8374,N_7573,N_7958);
and U8375 (N_8375,N_7991,N_7941);
xor U8376 (N_8376,N_8216,N_8143);
nor U8377 (N_8377,N_7527,N_7921);
nand U8378 (N_8378,N_7741,N_7796);
nand U8379 (N_8379,N_7934,N_7922);
and U8380 (N_8380,N_7844,N_7751);
or U8381 (N_8381,N_7964,N_8126);
and U8382 (N_8382,N_7888,N_7842);
nand U8383 (N_8383,N_8082,N_7660);
and U8384 (N_8384,N_7656,N_7610);
nand U8385 (N_8385,N_7881,N_7859);
and U8386 (N_8386,N_7528,N_7655);
and U8387 (N_8387,N_7901,N_7657);
nor U8388 (N_8388,N_7712,N_7953);
or U8389 (N_8389,N_8155,N_8244);
nand U8390 (N_8390,N_8133,N_7776);
or U8391 (N_8391,N_8169,N_7872);
or U8392 (N_8392,N_7766,N_7906);
nor U8393 (N_8393,N_8093,N_7867);
nor U8394 (N_8394,N_8168,N_8172);
and U8395 (N_8395,N_7786,N_7701);
nor U8396 (N_8396,N_8200,N_7990);
and U8397 (N_8397,N_8075,N_7736);
nand U8398 (N_8398,N_7539,N_7930);
nor U8399 (N_8399,N_7813,N_8058);
and U8400 (N_8400,N_8101,N_7989);
or U8401 (N_8401,N_8024,N_7644);
nor U8402 (N_8402,N_8211,N_7973);
or U8403 (N_8403,N_8231,N_7817);
and U8404 (N_8404,N_7974,N_7556);
or U8405 (N_8405,N_8039,N_7932);
nand U8406 (N_8406,N_8079,N_7725);
xnor U8407 (N_8407,N_7823,N_7933);
xor U8408 (N_8408,N_7918,N_7733);
and U8409 (N_8409,N_7532,N_8203);
nor U8410 (N_8410,N_7926,N_8130);
nor U8411 (N_8411,N_7970,N_7599);
nor U8412 (N_8412,N_8123,N_8195);
or U8413 (N_8413,N_7831,N_7667);
nand U8414 (N_8414,N_7763,N_8038);
nand U8415 (N_8415,N_8023,N_8191);
nor U8416 (N_8416,N_7577,N_7542);
nor U8417 (N_8417,N_7971,N_7861);
and U8418 (N_8418,N_7700,N_8002);
or U8419 (N_8419,N_7924,N_7770);
and U8420 (N_8420,N_7524,N_7952);
nor U8421 (N_8421,N_7778,N_7963);
nor U8422 (N_8422,N_8150,N_7628);
nor U8423 (N_8423,N_8119,N_8218);
and U8424 (N_8424,N_8113,N_7634);
and U8425 (N_8425,N_8111,N_8032);
or U8426 (N_8426,N_7902,N_7846);
nor U8427 (N_8427,N_7923,N_7841);
or U8428 (N_8428,N_8105,N_7909);
or U8429 (N_8429,N_8042,N_8247);
and U8430 (N_8430,N_7900,N_7614);
and U8431 (N_8431,N_7935,N_8178);
or U8432 (N_8432,N_7517,N_7531);
or U8433 (N_8433,N_8120,N_7961);
nand U8434 (N_8434,N_8213,N_8238);
nor U8435 (N_8435,N_8182,N_7597);
nor U8436 (N_8436,N_7931,N_8071);
and U8437 (N_8437,N_7714,N_8176);
or U8438 (N_8438,N_8006,N_7755);
nor U8439 (N_8439,N_7641,N_7645);
or U8440 (N_8440,N_7835,N_8000);
nand U8441 (N_8441,N_7903,N_7968);
and U8442 (N_8442,N_7775,N_7640);
nand U8443 (N_8443,N_8068,N_7581);
or U8444 (N_8444,N_7880,N_7651);
nand U8445 (N_8445,N_7643,N_7869);
or U8446 (N_8446,N_8165,N_8114);
and U8447 (N_8447,N_7563,N_7546);
nand U8448 (N_8448,N_8159,N_8031);
and U8449 (N_8449,N_8125,N_7500);
nand U8450 (N_8450,N_7836,N_8115);
and U8451 (N_8451,N_8212,N_7706);
and U8452 (N_8452,N_8152,N_7999);
nand U8453 (N_8453,N_7790,N_8180);
or U8454 (N_8454,N_7758,N_7834);
nor U8455 (N_8455,N_8110,N_7630);
or U8456 (N_8456,N_7913,N_7699);
or U8457 (N_8457,N_8064,N_8158);
or U8458 (N_8458,N_7908,N_7533);
and U8459 (N_8459,N_8078,N_7912);
nor U8460 (N_8460,N_8151,N_7591);
nand U8461 (N_8461,N_7543,N_7978);
or U8462 (N_8462,N_7749,N_8207);
or U8463 (N_8463,N_7635,N_7946);
or U8464 (N_8464,N_7740,N_8073);
and U8465 (N_8465,N_7688,N_7858);
and U8466 (N_8466,N_8219,N_7654);
or U8467 (N_8467,N_7947,N_7684);
and U8468 (N_8468,N_7724,N_7551);
or U8469 (N_8469,N_8026,N_7574);
nor U8470 (N_8470,N_7648,N_8067);
nand U8471 (N_8471,N_7986,N_7739);
and U8472 (N_8472,N_8030,N_8206);
nor U8473 (N_8473,N_8087,N_7826);
and U8474 (N_8474,N_7940,N_7865);
nor U8475 (N_8475,N_8145,N_7806);
and U8476 (N_8476,N_7730,N_8074);
and U8477 (N_8477,N_7689,N_7606);
nand U8478 (N_8478,N_7840,N_7633);
nand U8479 (N_8479,N_7627,N_7629);
nor U8480 (N_8480,N_7696,N_7549);
nand U8481 (N_8481,N_8072,N_7589);
nand U8482 (N_8482,N_7885,N_7509);
nor U8483 (N_8483,N_8228,N_8035);
nand U8484 (N_8484,N_7997,N_7984);
xor U8485 (N_8485,N_7816,N_7757);
or U8486 (N_8486,N_8248,N_8199);
and U8487 (N_8487,N_8048,N_8102);
nand U8488 (N_8488,N_7642,N_8175);
nand U8489 (N_8489,N_8044,N_7682);
nand U8490 (N_8490,N_7626,N_7955);
nor U8491 (N_8491,N_7580,N_7566);
or U8492 (N_8492,N_7928,N_7653);
and U8493 (N_8493,N_7686,N_7732);
nor U8494 (N_8494,N_7511,N_7852);
nor U8495 (N_8495,N_7987,N_7782);
or U8496 (N_8496,N_8066,N_8037);
nor U8497 (N_8497,N_8086,N_8090);
nor U8498 (N_8498,N_7609,N_8061);
nand U8499 (N_8499,N_8221,N_7693);
and U8500 (N_8500,N_7833,N_7704);
and U8501 (N_8501,N_7590,N_7756);
nand U8502 (N_8502,N_8204,N_8205);
nand U8503 (N_8503,N_7538,N_8192);
and U8504 (N_8504,N_7718,N_8116);
nand U8505 (N_8505,N_7521,N_7983);
nand U8506 (N_8506,N_8246,N_7891);
nor U8507 (N_8507,N_8092,N_8170);
or U8508 (N_8508,N_8222,N_7636);
or U8509 (N_8509,N_8018,N_8097);
nand U8510 (N_8510,N_8011,N_7754);
and U8511 (N_8511,N_8235,N_7638);
or U8512 (N_8512,N_8162,N_7547);
nor U8513 (N_8513,N_7707,N_7837);
nand U8514 (N_8514,N_7600,N_7855);
and U8515 (N_8515,N_7760,N_7747);
nor U8516 (N_8516,N_7555,N_8208);
and U8517 (N_8517,N_7649,N_7856);
nor U8518 (N_8518,N_7694,N_8229);
and U8519 (N_8519,N_7808,N_7860);
nand U8520 (N_8520,N_7584,N_8201);
or U8521 (N_8521,N_7510,N_7665);
and U8522 (N_8522,N_7998,N_7719);
or U8523 (N_8523,N_7613,N_7697);
nor U8524 (N_8524,N_8215,N_7548);
and U8525 (N_8525,N_7674,N_7915);
and U8526 (N_8526,N_7612,N_7637);
nor U8527 (N_8527,N_7769,N_8227);
nor U8528 (N_8528,N_7565,N_7738);
or U8529 (N_8529,N_8183,N_7621);
and U8530 (N_8530,N_7789,N_7752);
and U8531 (N_8531,N_7969,N_8020);
and U8532 (N_8532,N_7526,N_7523);
nor U8533 (N_8533,N_7745,N_7721);
nand U8534 (N_8534,N_7569,N_7650);
or U8535 (N_8535,N_7765,N_7557);
nand U8536 (N_8536,N_7792,N_8021);
and U8537 (N_8537,N_7728,N_7568);
xnor U8538 (N_8538,N_8239,N_7579);
nand U8539 (N_8539,N_7781,N_8185);
or U8540 (N_8540,N_7960,N_8129);
or U8541 (N_8541,N_7691,N_7623);
nand U8542 (N_8542,N_7515,N_8164);
and U8543 (N_8543,N_7508,N_8179);
or U8544 (N_8544,N_8121,N_8043);
and U8545 (N_8545,N_7615,N_8232);
or U8546 (N_8546,N_7878,N_7519);
or U8547 (N_8547,N_7993,N_7678);
nor U8548 (N_8548,N_7798,N_7771);
and U8549 (N_8549,N_8036,N_7692);
nand U8550 (N_8550,N_7605,N_8109);
and U8551 (N_8551,N_8025,N_7661);
nor U8552 (N_8552,N_7843,N_7550);
nor U8553 (N_8553,N_7679,N_7761);
nand U8554 (N_8554,N_8197,N_8184);
and U8555 (N_8555,N_8054,N_8198);
nor U8556 (N_8556,N_8209,N_8004);
nor U8557 (N_8557,N_8055,N_7673);
and U8558 (N_8558,N_7914,N_7540);
or U8559 (N_8559,N_7604,N_7936);
or U8560 (N_8560,N_7899,N_8220);
or U8561 (N_8561,N_7753,N_7807);
and U8562 (N_8562,N_7595,N_7884);
nor U8563 (N_8563,N_8103,N_7603);
nand U8564 (N_8564,N_8019,N_7731);
nor U8565 (N_8565,N_7779,N_8099);
nor U8566 (N_8566,N_7898,N_7980);
nand U8567 (N_8567,N_7625,N_7920);
nand U8568 (N_8568,N_8106,N_7797);
or U8569 (N_8569,N_7698,N_7820);
and U8570 (N_8570,N_7677,N_7904);
and U8571 (N_8571,N_7929,N_7680);
or U8572 (N_8572,N_8234,N_7814);
nand U8573 (N_8573,N_8187,N_7502);
nor U8574 (N_8574,N_7735,N_7851);
or U8575 (N_8575,N_7917,N_7966);
or U8576 (N_8576,N_7578,N_7839);
or U8577 (N_8577,N_8060,N_7571);
or U8578 (N_8578,N_8163,N_7785);
or U8579 (N_8579,N_7956,N_7976);
or U8580 (N_8580,N_7850,N_7552);
and U8581 (N_8581,N_7662,N_7979);
and U8582 (N_8582,N_7982,N_7948);
nor U8583 (N_8583,N_7586,N_8053);
and U8584 (N_8584,N_7879,N_7631);
and U8585 (N_8585,N_7905,N_7954);
nand U8586 (N_8586,N_7849,N_8104);
or U8587 (N_8587,N_7534,N_8070);
nor U8588 (N_8588,N_8181,N_8134);
and U8589 (N_8589,N_8084,N_7601);
nor U8590 (N_8590,N_7847,N_7522);
nor U8591 (N_8591,N_8138,N_8224);
or U8592 (N_8592,N_7564,N_8083);
or U8593 (N_8593,N_7897,N_8088);
nand U8594 (N_8594,N_8137,N_7588);
nor U8595 (N_8595,N_8241,N_8108);
nor U8596 (N_8596,N_7690,N_7805);
nand U8597 (N_8597,N_7773,N_8096);
nand U8598 (N_8598,N_7994,N_8188);
and U8599 (N_8599,N_8202,N_7558);
nor U8600 (N_8600,N_8196,N_7838);
and U8601 (N_8601,N_7845,N_7742);
or U8602 (N_8602,N_7825,N_8041);
nand U8603 (N_8603,N_7848,N_7737);
nand U8604 (N_8604,N_7619,N_7664);
nor U8605 (N_8605,N_7525,N_7873);
and U8606 (N_8606,N_7810,N_7687);
and U8607 (N_8607,N_7890,N_8017);
and U8608 (N_8608,N_8167,N_7949);
nor U8609 (N_8609,N_8059,N_8003);
or U8610 (N_8610,N_7560,N_8147);
and U8611 (N_8611,N_7893,N_8140);
or U8612 (N_8612,N_8135,N_8117);
or U8613 (N_8613,N_7512,N_7544);
nor U8614 (N_8614,N_7988,N_7959);
or U8615 (N_8615,N_7676,N_7894);
or U8616 (N_8616,N_7681,N_7977);
and U8617 (N_8617,N_7759,N_8127);
and U8618 (N_8618,N_7895,N_7862);
or U8619 (N_8619,N_7883,N_7708);
and U8620 (N_8620,N_8166,N_7520);
or U8621 (N_8621,N_7575,N_7652);
nand U8622 (N_8622,N_8027,N_8089);
nor U8623 (N_8623,N_8124,N_7876);
nand U8624 (N_8624,N_8047,N_8051);
or U8625 (N_8625,N_7826,N_8053);
or U8626 (N_8626,N_8022,N_7709);
or U8627 (N_8627,N_8162,N_8155);
nand U8628 (N_8628,N_8202,N_7711);
and U8629 (N_8629,N_7692,N_7582);
and U8630 (N_8630,N_7699,N_8072);
nor U8631 (N_8631,N_8152,N_8190);
nor U8632 (N_8632,N_8033,N_7657);
or U8633 (N_8633,N_7903,N_7951);
nor U8634 (N_8634,N_7708,N_8064);
and U8635 (N_8635,N_7590,N_7692);
and U8636 (N_8636,N_8109,N_7876);
xor U8637 (N_8637,N_7803,N_7927);
nor U8638 (N_8638,N_7800,N_8089);
xnor U8639 (N_8639,N_8058,N_8161);
or U8640 (N_8640,N_7824,N_7904);
nor U8641 (N_8641,N_8247,N_8052);
or U8642 (N_8642,N_7876,N_7547);
or U8643 (N_8643,N_7977,N_7968);
and U8644 (N_8644,N_8190,N_7668);
and U8645 (N_8645,N_8004,N_7831);
nor U8646 (N_8646,N_7687,N_7973);
nor U8647 (N_8647,N_8174,N_8243);
nor U8648 (N_8648,N_7800,N_7818);
and U8649 (N_8649,N_7833,N_7608);
nor U8650 (N_8650,N_7610,N_7882);
nand U8651 (N_8651,N_7594,N_7565);
nor U8652 (N_8652,N_7902,N_8049);
or U8653 (N_8653,N_8108,N_7673);
nand U8654 (N_8654,N_7685,N_8158);
nor U8655 (N_8655,N_8057,N_8244);
or U8656 (N_8656,N_7646,N_7643);
or U8657 (N_8657,N_8026,N_8033);
or U8658 (N_8658,N_7905,N_7681);
nor U8659 (N_8659,N_7939,N_7754);
nand U8660 (N_8660,N_8179,N_7765);
nand U8661 (N_8661,N_7653,N_7963);
nor U8662 (N_8662,N_7744,N_7965);
or U8663 (N_8663,N_7865,N_7870);
and U8664 (N_8664,N_8221,N_7697);
or U8665 (N_8665,N_7992,N_7714);
nand U8666 (N_8666,N_7924,N_7794);
and U8667 (N_8667,N_7562,N_7539);
and U8668 (N_8668,N_7581,N_8135);
nand U8669 (N_8669,N_7653,N_8052);
nand U8670 (N_8670,N_8246,N_8045);
and U8671 (N_8671,N_7883,N_7530);
nor U8672 (N_8672,N_7706,N_8036);
or U8673 (N_8673,N_7524,N_8044);
nor U8674 (N_8674,N_7881,N_7529);
xnor U8675 (N_8675,N_7846,N_8113);
or U8676 (N_8676,N_8008,N_8050);
and U8677 (N_8677,N_7996,N_7800);
nand U8678 (N_8678,N_7641,N_7614);
or U8679 (N_8679,N_8197,N_7718);
nand U8680 (N_8680,N_7542,N_8159);
nor U8681 (N_8681,N_8196,N_7622);
nand U8682 (N_8682,N_7508,N_7745);
and U8683 (N_8683,N_7779,N_7837);
or U8684 (N_8684,N_8097,N_7853);
nor U8685 (N_8685,N_7958,N_7902);
and U8686 (N_8686,N_7889,N_7674);
nand U8687 (N_8687,N_8098,N_7624);
and U8688 (N_8688,N_7825,N_7890);
nand U8689 (N_8689,N_8217,N_7935);
or U8690 (N_8690,N_7539,N_7588);
and U8691 (N_8691,N_7629,N_7560);
or U8692 (N_8692,N_7900,N_7506);
nand U8693 (N_8693,N_8047,N_7763);
nand U8694 (N_8694,N_7689,N_7994);
nand U8695 (N_8695,N_7639,N_7796);
and U8696 (N_8696,N_8123,N_7569);
nand U8697 (N_8697,N_7864,N_7805);
nor U8698 (N_8698,N_8224,N_7846);
and U8699 (N_8699,N_8193,N_7736);
nor U8700 (N_8700,N_7640,N_7928);
and U8701 (N_8701,N_7900,N_7716);
nor U8702 (N_8702,N_8035,N_7659);
or U8703 (N_8703,N_7871,N_8011);
and U8704 (N_8704,N_8208,N_7744);
nand U8705 (N_8705,N_7580,N_7554);
nand U8706 (N_8706,N_7597,N_7887);
or U8707 (N_8707,N_7854,N_7942);
or U8708 (N_8708,N_8233,N_8208);
nand U8709 (N_8709,N_8200,N_8237);
and U8710 (N_8710,N_7744,N_7720);
nand U8711 (N_8711,N_8041,N_7960);
or U8712 (N_8712,N_7662,N_7658);
nor U8713 (N_8713,N_7911,N_7707);
or U8714 (N_8714,N_7577,N_7936);
and U8715 (N_8715,N_7585,N_7767);
and U8716 (N_8716,N_7695,N_7988);
nand U8717 (N_8717,N_7748,N_8037);
nand U8718 (N_8718,N_8151,N_7578);
or U8719 (N_8719,N_7949,N_7677);
nand U8720 (N_8720,N_8138,N_8203);
nor U8721 (N_8721,N_7506,N_8196);
nand U8722 (N_8722,N_7721,N_7707);
and U8723 (N_8723,N_7817,N_7614);
and U8724 (N_8724,N_7574,N_7660);
or U8725 (N_8725,N_8190,N_7551);
nand U8726 (N_8726,N_7872,N_8055);
nand U8727 (N_8727,N_7716,N_7751);
and U8728 (N_8728,N_7740,N_7779);
and U8729 (N_8729,N_7970,N_7932);
and U8730 (N_8730,N_8037,N_8032);
and U8731 (N_8731,N_8221,N_8086);
and U8732 (N_8732,N_8035,N_7613);
or U8733 (N_8733,N_7517,N_7822);
nand U8734 (N_8734,N_7615,N_7710);
nor U8735 (N_8735,N_7848,N_8032);
nand U8736 (N_8736,N_7885,N_7733);
and U8737 (N_8737,N_7957,N_8166);
nor U8738 (N_8738,N_7628,N_8124);
and U8739 (N_8739,N_7940,N_7811);
nor U8740 (N_8740,N_7505,N_7697);
nand U8741 (N_8741,N_8152,N_8224);
or U8742 (N_8742,N_7774,N_7754);
xnor U8743 (N_8743,N_7688,N_7618);
nand U8744 (N_8744,N_7863,N_7891);
or U8745 (N_8745,N_8215,N_7933);
nor U8746 (N_8746,N_7598,N_7990);
or U8747 (N_8747,N_8195,N_7714);
nor U8748 (N_8748,N_7637,N_7724);
or U8749 (N_8749,N_7811,N_7609);
and U8750 (N_8750,N_7549,N_8181);
xnor U8751 (N_8751,N_8235,N_8226);
or U8752 (N_8752,N_8247,N_7730);
or U8753 (N_8753,N_7994,N_7693);
or U8754 (N_8754,N_7565,N_8229);
nand U8755 (N_8755,N_8162,N_8191);
or U8756 (N_8756,N_7704,N_8059);
nor U8757 (N_8757,N_7604,N_7804);
or U8758 (N_8758,N_7962,N_7744);
nor U8759 (N_8759,N_7775,N_8030);
nand U8760 (N_8760,N_7550,N_8043);
nor U8761 (N_8761,N_7671,N_7687);
nor U8762 (N_8762,N_8057,N_7531);
and U8763 (N_8763,N_7568,N_8099);
or U8764 (N_8764,N_7893,N_8182);
nor U8765 (N_8765,N_7605,N_8022);
or U8766 (N_8766,N_7915,N_7765);
nand U8767 (N_8767,N_8080,N_7982);
nand U8768 (N_8768,N_7503,N_8085);
or U8769 (N_8769,N_7591,N_8078);
nand U8770 (N_8770,N_7806,N_7874);
nand U8771 (N_8771,N_7864,N_7676);
or U8772 (N_8772,N_8160,N_8127);
and U8773 (N_8773,N_7645,N_7549);
nor U8774 (N_8774,N_8185,N_7758);
and U8775 (N_8775,N_8249,N_7521);
nor U8776 (N_8776,N_7974,N_7656);
nand U8777 (N_8777,N_7924,N_7646);
and U8778 (N_8778,N_8065,N_7883);
nand U8779 (N_8779,N_8096,N_7955);
and U8780 (N_8780,N_7847,N_8210);
and U8781 (N_8781,N_7759,N_8176);
and U8782 (N_8782,N_7529,N_7748);
or U8783 (N_8783,N_7989,N_7837);
or U8784 (N_8784,N_8063,N_8074);
nand U8785 (N_8785,N_7500,N_8135);
nor U8786 (N_8786,N_7975,N_7925);
or U8787 (N_8787,N_7839,N_7961);
nor U8788 (N_8788,N_7604,N_7542);
nor U8789 (N_8789,N_8099,N_7912);
nor U8790 (N_8790,N_7875,N_7844);
nand U8791 (N_8791,N_8243,N_7765);
nand U8792 (N_8792,N_8039,N_7717);
or U8793 (N_8793,N_7961,N_8133);
nor U8794 (N_8794,N_7583,N_7922);
nand U8795 (N_8795,N_8051,N_7792);
nor U8796 (N_8796,N_7823,N_7832);
nor U8797 (N_8797,N_7884,N_7566);
or U8798 (N_8798,N_8144,N_7529);
and U8799 (N_8799,N_8124,N_8232);
nor U8800 (N_8800,N_7898,N_8126);
nand U8801 (N_8801,N_7519,N_7594);
nand U8802 (N_8802,N_7791,N_7588);
nand U8803 (N_8803,N_7999,N_7657);
nand U8804 (N_8804,N_8007,N_7846);
nor U8805 (N_8805,N_7604,N_7559);
nand U8806 (N_8806,N_7775,N_7571);
or U8807 (N_8807,N_7905,N_8113);
and U8808 (N_8808,N_8079,N_7533);
or U8809 (N_8809,N_8248,N_7654);
nand U8810 (N_8810,N_7875,N_7878);
nand U8811 (N_8811,N_7808,N_8122);
nand U8812 (N_8812,N_7653,N_7623);
nor U8813 (N_8813,N_8007,N_7605);
nand U8814 (N_8814,N_8116,N_7579);
nand U8815 (N_8815,N_7999,N_7502);
nand U8816 (N_8816,N_7949,N_7589);
nor U8817 (N_8817,N_8188,N_8034);
nor U8818 (N_8818,N_8088,N_7875);
nor U8819 (N_8819,N_7609,N_7796);
xnor U8820 (N_8820,N_7784,N_7601);
and U8821 (N_8821,N_7903,N_8236);
nor U8822 (N_8822,N_8222,N_7644);
and U8823 (N_8823,N_7808,N_8192);
or U8824 (N_8824,N_7987,N_7734);
and U8825 (N_8825,N_7710,N_7665);
or U8826 (N_8826,N_7725,N_7984);
and U8827 (N_8827,N_8059,N_8222);
or U8828 (N_8828,N_7810,N_8200);
or U8829 (N_8829,N_7525,N_8031);
nor U8830 (N_8830,N_8106,N_7721);
or U8831 (N_8831,N_7517,N_8086);
nand U8832 (N_8832,N_8035,N_7716);
or U8833 (N_8833,N_7786,N_7587);
nor U8834 (N_8834,N_7754,N_8013);
nand U8835 (N_8835,N_7745,N_7604);
nand U8836 (N_8836,N_7562,N_8184);
or U8837 (N_8837,N_8126,N_8019);
nor U8838 (N_8838,N_8162,N_7955);
or U8839 (N_8839,N_8081,N_7935);
nand U8840 (N_8840,N_7595,N_7847);
nor U8841 (N_8841,N_8149,N_7878);
nand U8842 (N_8842,N_7992,N_7940);
and U8843 (N_8843,N_7672,N_7603);
and U8844 (N_8844,N_8203,N_8077);
nand U8845 (N_8845,N_7850,N_7990);
or U8846 (N_8846,N_8031,N_7835);
nor U8847 (N_8847,N_7670,N_7758);
or U8848 (N_8848,N_7973,N_7698);
nor U8849 (N_8849,N_7935,N_8052);
nand U8850 (N_8850,N_7726,N_7779);
or U8851 (N_8851,N_7562,N_7895);
nand U8852 (N_8852,N_7601,N_7551);
nand U8853 (N_8853,N_7697,N_8039);
or U8854 (N_8854,N_7669,N_8243);
nor U8855 (N_8855,N_7932,N_8073);
nand U8856 (N_8856,N_8007,N_7928);
and U8857 (N_8857,N_7637,N_8050);
nor U8858 (N_8858,N_8204,N_7716);
and U8859 (N_8859,N_8033,N_8162);
nor U8860 (N_8860,N_8224,N_7775);
and U8861 (N_8861,N_7722,N_7991);
nand U8862 (N_8862,N_8034,N_7645);
or U8863 (N_8863,N_7716,N_7547);
nand U8864 (N_8864,N_8153,N_8023);
nor U8865 (N_8865,N_8071,N_8049);
nor U8866 (N_8866,N_8187,N_7799);
nor U8867 (N_8867,N_7927,N_8234);
and U8868 (N_8868,N_8093,N_8238);
and U8869 (N_8869,N_7783,N_7949);
or U8870 (N_8870,N_7540,N_7547);
and U8871 (N_8871,N_7828,N_7865);
nand U8872 (N_8872,N_8016,N_7845);
nand U8873 (N_8873,N_8040,N_8229);
nand U8874 (N_8874,N_7992,N_7845);
nand U8875 (N_8875,N_8219,N_7792);
or U8876 (N_8876,N_7703,N_7958);
nor U8877 (N_8877,N_7673,N_7500);
nor U8878 (N_8878,N_8016,N_8196);
nor U8879 (N_8879,N_7870,N_7608);
or U8880 (N_8880,N_7594,N_7536);
and U8881 (N_8881,N_7881,N_7867);
nand U8882 (N_8882,N_7830,N_8111);
nor U8883 (N_8883,N_7681,N_8218);
nand U8884 (N_8884,N_8129,N_7698);
nor U8885 (N_8885,N_8077,N_8160);
nand U8886 (N_8886,N_7596,N_8054);
or U8887 (N_8887,N_8148,N_7647);
and U8888 (N_8888,N_8136,N_7834);
or U8889 (N_8889,N_7704,N_7662);
and U8890 (N_8890,N_8165,N_7649);
or U8891 (N_8891,N_7595,N_7852);
or U8892 (N_8892,N_8157,N_8177);
nor U8893 (N_8893,N_8070,N_8042);
and U8894 (N_8894,N_7731,N_7823);
nand U8895 (N_8895,N_8216,N_8123);
or U8896 (N_8896,N_8073,N_7580);
nand U8897 (N_8897,N_8031,N_7507);
and U8898 (N_8898,N_8171,N_7841);
nor U8899 (N_8899,N_7623,N_7811);
nor U8900 (N_8900,N_7725,N_7740);
nand U8901 (N_8901,N_7731,N_7545);
nor U8902 (N_8902,N_7716,N_7709);
nand U8903 (N_8903,N_8183,N_7887);
and U8904 (N_8904,N_7791,N_7859);
nor U8905 (N_8905,N_7616,N_7864);
nor U8906 (N_8906,N_8186,N_8171);
nor U8907 (N_8907,N_8051,N_7938);
nor U8908 (N_8908,N_7609,N_7522);
nor U8909 (N_8909,N_7747,N_7756);
xnor U8910 (N_8910,N_7590,N_7912);
nor U8911 (N_8911,N_7662,N_8041);
and U8912 (N_8912,N_7883,N_7742);
or U8913 (N_8913,N_8098,N_7552);
nand U8914 (N_8914,N_8082,N_7999);
and U8915 (N_8915,N_7554,N_8166);
or U8916 (N_8916,N_7629,N_8037);
or U8917 (N_8917,N_8153,N_7749);
or U8918 (N_8918,N_7836,N_7820);
and U8919 (N_8919,N_7782,N_8084);
and U8920 (N_8920,N_7759,N_7969);
and U8921 (N_8921,N_8087,N_8125);
and U8922 (N_8922,N_7519,N_7988);
and U8923 (N_8923,N_8006,N_7804);
nor U8924 (N_8924,N_7627,N_7865);
or U8925 (N_8925,N_8245,N_7994);
or U8926 (N_8926,N_7554,N_7875);
nand U8927 (N_8927,N_8175,N_8029);
or U8928 (N_8928,N_7938,N_8189);
nand U8929 (N_8929,N_8027,N_7513);
nand U8930 (N_8930,N_8166,N_7738);
and U8931 (N_8931,N_8239,N_8086);
nor U8932 (N_8932,N_7509,N_7930);
or U8933 (N_8933,N_7962,N_7938);
nor U8934 (N_8934,N_8035,N_7956);
nor U8935 (N_8935,N_7531,N_7581);
or U8936 (N_8936,N_7882,N_8244);
and U8937 (N_8937,N_8108,N_7559);
and U8938 (N_8938,N_7891,N_8137);
or U8939 (N_8939,N_8113,N_7744);
or U8940 (N_8940,N_7756,N_7898);
nand U8941 (N_8941,N_8076,N_7506);
nor U8942 (N_8942,N_8197,N_7988);
nand U8943 (N_8943,N_7726,N_8002);
and U8944 (N_8944,N_7642,N_7662);
or U8945 (N_8945,N_8126,N_7952);
or U8946 (N_8946,N_8145,N_7785);
nand U8947 (N_8947,N_7969,N_7652);
nand U8948 (N_8948,N_7688,N_8092);
nand U8949 (N_8949,N_7949,N_7930);
and U8950 (N_8950,N_8020,N_8086);
or U8951 (N_8951,N_7716,N_8070);
or U8952 (N_8952,N_8051,N_7742);
nor U8953 (N_8953,N_7742,N_7850);
or U8954 (N_8954,N_8062,N_7803);
nor U8955 (N_8955,N_7781,N_7882);
or U8956 (N_8956,N_7619,N_8063);
nor U8957 (N_8957,N_7508,N_7605);
and U8958 (N_8958,N_7657,N_8020);
nor U8959 (N_8959,N_8043,N_7834);
or U8960 (N_8960,N_7826,N_8232);
nor U8961 (N_8961,N_7776,N_8124);
and U8962 (N_8962,N_7618,N_7529);
nand U8963 (N_8963,N_7712,N_7809);
nand U8964 (N_8964,N_7980,N_8076);
nor U8965 (N_8965,N_7819,N_7668);
and U8966 (N_8966,N_7942,N_7848);
or U8967 (N_8967,N_8006,N_7590);
nor U8968 (N_8968,N_8118,N_7947);
nor U8969 (N_8969,N_7798,N_8153);
or U8970 (N_8970,N_8160,N_7593);
nor U8971 (N_8971,N_7536,N_7580);
or U8972 (N_8972,N_7695,N_7829);
or U8973 (N_8973,N_8003,N_8208);
and U8974 (N_8974,N_8136,N_7780);
nor U8975 (N_8975,N_7723,N_7616);
and U8976 (N_8976,N_7949,N_8202);
nor U8977 (N_8977,N_7709,N_8216);
and U8978 (N_8978,N_8051,N_7705);
or U8979 (N_8979,N_7818,N_8102);
nand U8980 (N_8980,N_8229,N_7617);
or U8981 (N_8981,N_7962,N_7600);
or U8982 (N_8982,N_7681,N_7580);
and U8983 (N_8983,N_7690,N_8087);
nand U8984 (N_8984,N_7774,N_7761);
and U8985 (N_8985,N_8160,N_7535);
and U8986 (N_8986,N_7705,N_7663);
or U8987 (N_8987,N_7974,N_8040);
nand U8988 (N_8988,N_7930,N_7752);
nand U8989 (N_8989,N_7721,N_8228);
or U8990 (N_8990,N_7942,N_7531);
and U8991 (N_8991,N_8198,N_7809);
nor U8992 (N_8992,N_7580,N_7909);
and U8993 (N_8993,N_7793,N_8241);
nor U8994 (N_8994,N_7912,N_7822);
nand U8995 (N_8995,N_7527,N_8040);
or U8996 (N_8996,N_8177,N_8047);
and U8997 (N_8997,N_8088,N_7871);
and U8998 (N_8998,N_7825,N_7617);
and U8999 (N_8999,N_8212,N_8169);
nand U9000 (N_9000,N_8568,N_8795);
and U9001 (N_9001,N_8834,N_8565);
or U9002 (N_9002,N_8672,N_8355);
or U9003 (N_9003,N_8490,N_8342);
or U9004 (N_9004,N_8854,N_8633);
and U9005 (N_9005,N_8442,N_8901);
or U9006 (N_9006,N_8932,N_8805);
and U9007 (N_9007,N_8474,N_8972);
nor U9008 (N_9008,N_8642,N_8439);
or U9009 (N_9009,N_8971,N_8992);
nor U9010 (N_9010,N_8626,N_8622);
and U9011 (N_9011,N_8542,N_8464);
or U9012 (N_9012,N_8373,N_8598);
and U9013 (N_9013,N_8462,N_8806);
nor U9014 (N_9014,N_8870,N_8552);
and U9015 (N_9015,N_8832,N_8758);
and U9016 (N_9016,N_8882,N_8554);
nor U9017 (N_9017,N_8619,N_8727);
or U9018 (N_9018,N_8657,N_8323);
or U9019 (N_9019,N_8859,N_8815);
nand U9020 (N_9020,N_8690,N_8850);
nor U9021 (N_9021,N_8989,N_8766);
nor U9022 (N_9022,N_8592,N_8845);
or U9023 (N_9023,N_8998,N_8943);
and U9024 (N_9024,N_8480,N_8441);
or U9025 (N_9025,N_8829,N_8278);
or U9026 (N_9026,N_8798,N_8713);
and U9027 (N_9027,N_8425,N_8652);
nor U9028 (N_9028,N_8849,N_8263);
and U9029 (N_9029,N_8863,N_8506);
or U9030 (N_9030,N_8827,N_8505);
nor U9031 (N_9031,N_8694,N_8327);
nand U9032 (N_9032,N_8538,N_8684);
and U9033 (N_9033,N_8299,N_8303);
nand U9034 (N_9034,N_8701,N_8584);
or U9035 (N_9035,N_8364,N_8520);
nand U9036 (N_9036,N_8985,N_8775);
and U9037 (N_9037,N_8774,N_8874);
nor U9038 (N_9038,N_8884,N_8852);
and U9039 (N_9039,N_8340,N_8422);
or U9040 (N_9040,N_8731,N_8498);
nor U9041 (N_9041,N_8939,N_8305);
nand U9042 (N_9042,N_8999,N_8277);
nor U9043 (N_9043,N_8463,N_8624);
or U9044 (N_9044,N_8281,N_8344);
nor U9045 (N_9045,N_8888,N_8258);
or U9046 (N_9046,N_8530,N_8679);
nor U9047 (N_9047,N_8458,N_8754);
nand U9048 (N_9048,N_8535,N_8778);
and U9049 (N_9049,N_8986,N_8401);
and U9050 (N_9050,N_8251,N_8508);
nor U9051 (N_9051,N_8447,N_8937);
and U9052 (N_9052,N_8362,N_8335);
and U9053 (N_9053,N_8322,N_8835);
nand U9054 (N_9054,N_8523,N_8651);
xnor U9055 (N_9055,N_8471,N_8454);
nand U9056 (N_9056,N_8744,N_8846);
nand U9057 (N_9057,N_8764,N_8519);
or U9058 (N_9058,N_8319,N_8430);
or U9059 (N_9059,N_8872,N_8759);
nor U9060 (N_9060,N_8638,N_8489);
nand U9061 (N_9061,N_8631,N_8532);
or U9062 (N_9062,N_8963,N_8976);
or U9063 (N_9063,N_8499,N_8749);
nand U9064 (N_9064,N_8708,N_8296);
or U9065 (N_9065,N_8867,N_8803);
nand U9066 (N_9066,N_8929,N_8644);
nor U9067 (N_9067,N_8515,N_8715);
and U9068 (N_9068,N_8533,N_8368);
and U9069 (N_9069,N_8830,N_8324);
and U9070 (N_9070,N_8625,N_8881);
and U9071 (N_9071,N_8583,N_8313);
nor U9072 (N_9072,N_8814,N_8421);
nand U9073 (N_9073,N_8397,N_8918);
and U9074 (N_9074,N_8593,N_8602);
nand U9075 (N_9075,N_8947,N_8733);
and U9076 (N_9076,N_8879,N_8496);
and U9077 (N_9077,N_8514,N_8351);
or U9078 (N_9078,N_8525,N_8370);
and U9079 (N_9079,N_8682,N_8786);
nor U9080 (N_9080,N_8561,N_8403);
nor U9081 (N_9081,N_8928,N_8777);
and U9082 (N_9082,N_8876,N_8391);
and U9083 (N_9083,N_8477,N_8383);
nand U9084 (N_9084,N_8767,N_8415);
nor U9085 (N_9085,N_8930,N_8635);
nor U9086 (N_9086,N_8276,N_8528);
nand U9087 (N_9087,N_8892,N_8321);
nand U9088 (N_9088,N_8800,N_8941);
or U9089 (N_9089,N_8910,N_8676);
or U9090 (N_9090,N_8659,N_8896);
nor U9091 (N_9091,N_8686,N_8261);
and U9092 (N_9092,N_8637,N_8265);
or U9093 (N_9093,N_8467,N_8497);
and U9094 (N_9094,N_8601,N_8495);
nor U9095 (N_9095,N_8577,N_8275);
nand U9096 (N_9096,N_8712,N_8536);
nor U9097 (N_9097,N_8377,N_8311);
nor U9098 (N_9098,N_8994,N_8997);
nor U9099 (N_9099,N_8649,N_8501);
nor U9100 (N_9100,N_8527,N_8360);
or U9101 (N_9101,N_8379,N_8504);
or U9102 (N_9102,N_8628,N_8309);
or U9103 (N_9103,N_8955,N_8529);
and U9104 (N_9104,N_8449,N_8641);
nor U9105 (N_9105,N_8558,N_8609);
or U9106 (N_9106,N_8952,N_8349);
nor U9107 (N_9107,N_8640,N_8469);
and U9108 (N_9108,N_8868,N_8297);
nand U9109 (N_9109,N_8616,N_8451);
or U9110 (N_9110,N_8877,N_8295);
nand U9111 (N_9111,N_8511,N_8329);
and U9112 (N_9112,N_8500,N_8889);
nor U9113 (N_9113,N_8596,N_8784);
nor U9114 (N_9114,N_8510,N_8747);
or U9115 (N_9115,N_8540,N_8376);
and U9116 (N_9116,N_8902,N_8424);
or U9117 (N_9117,N_8338,N_8613);
nor U9118 (N_9118,N_8267,N_8546);
or U9119 (N_9119,N_8770,N_8435);
nor U9120 (N_9120,N_8352,N_8799);
and U9121 (N_9121,N_8844,N_8785);
or U9122 (N_9122,N_8663,N_8954);
and U9123 (N_9123,N_8434,N_8361);
or U9124 (N_9124,N_8356,N_8250);
nand U9125 (N_9125,N_8949,N_8962);
or U9126 (N_9126,N_8757,N_8730);
or U9127 (N_9127,N_8919,N_8857);
nand U9128 (N_9128,N_8917,N_8860);
and U9129 (N_9129,N_8594,N_8861);
and U9130 (N_9130,N_8665,N_8869);
nor U9131 (N_9131,N_8559,N_8959);
and U9132 (N_9132,N_8936,N_8433);
nor U9133 (N_9133,N_8965,N_8550);
nor U9134 (N_9134,N_8746,N_8621);
nand U9135 (N_9135,N_8804,N_8655);
or U9136 (N_9136,N_8518,N_8371);
or U9137 (N_9137,N_8721,N_8466);
and U9138 (N_9138,N_8838,N_8560);
and U9139 (N_9139,N_8650,N_8308);
and U9140 (N_9140,N_8916,N_8906);
nor U9141 (N_9141,N_8951,N_8555);
or U9142 (N_9142,N_8871,N_8808);
or U9143 (N_9143,N_8534,N_8885);
and U9144 (N_9144,N_8571,N_8562);
or U9145 (N_9145,N_8851,N_8390);
or U9146 (N_9146,N_8891,N_8456);
and U9147 (N_9147,N_8410,N_8366);
or U9148 (N_9148,N_8790,N_8841);
or U9149 (N_9149,N_8807,N_8612);
or U9150 (N_9150,N_8703,N_8933);
xnor U9151 (N_9151,N_8605,N_8330);
nor U9152 (N_9152,N_8492,N_8938);
or U9153 (N_9153,N_8611,N_8387);
nand U9154 (N_9154,N_8465,N_8486);
nand U9155 (N_9155,N_8260,N_8942);
nand U9156 (N_9156,N_8292,N_8266);
nor U9157 (N_9157,N_8887,N_8911);
nand U9158 (N_9158,N_8796,N_8705);
nand U9159 (N_9159,N_8945,N_8252);
nand U9160 (N_9160,N_8283,N_8755);
nand U9161 (N_9161,N_8318,N_8468);
nand U9162 (N_9162,N_8895,N_8788);
and U9163 (N_9163,N_8839,N_8685);
or U9164 (N_9164,N_8543,N_8620);
nor U9165 (N_9165,N_8893,N_8446);
or U9166 (N_9166,N_8473,N_8566);
nand U9167 (N_9167,N_8697,N_8894);
nand U9168 (N_9168,N_8255,N_8926);
nor U9169 (N_9169,N_8953,N_8588);
nor U9170 (N_9170,N_8729,N_8950);
or U9171 (N_9171,N_8284,N_8981);
and U9172 (N_9172,N_8294,N_8946);
nor U9173 (N_9173,N_8873,N_8453);
nand U9174 (N_9174,N_8545,N_8964);
nand U9175 (N_9175,N_8481,N_8272);
nand U9176 (N_9176,N_8984,N_8334);
or U9177 (N_9177,N_8789,N_8833);
nor U9178 (N_9178,N_8580,N_8769);
nor U9179 (N_9179,N_8865,N_8810);
or U9180 (N_9180,N_8987,N_8494);
and U9181 (N_9181,N_8699,N_8760);
nor U9182 (N_9182,N_8812,N_8512);
or U9183 (N_9183,N_8380,N_8429);
nand U9184 (N_9184,N_8818,N_8956);
nand U9185 (N_9185,N_8483,N_8978);
nor U9186 (N_9186,N_8811,N_8742);
and U9187 (N_9187,N_8677,N_8793);
or U9188 (N_9188,N_8618,N_8670);
nand U9189 (N_9189,N_8801,N_8988);
and U9190 (N_9190,N_8979,N_8751);
and U9191 (N_9191,N_8488,N_8572);
or U9192 (N_9192,N_8634,N_8966);
and U9193 (N_9193,N_8343,N_8781);
nand U9194 (N_9194,N_8516,N_8413);
nor U9195 (N_9195,N_8678,N_8802);
and U9196 (N_9196,N_8734,N_8600);
and U9197 (N_9197,N_8502,N_8925);
nor U9198 (N_9198,N_8270,N_8521);
and U9199 (N_9199,N_8875,N_8432);
or U9200 (N_9200,N_8549,N_8898);
or U9201 (N_9201,N_8382,N_8688);
nand U9202 (N_9202,N_8262,N_8912);
nand U9203 (N_9203,N_8298,N_8569);
nor U9204 (N_9204,N_8743,N_8363);
nand U9205 (N_9205,N_8585,N_8900);
xnor U9206 (N_9206,N_8692,N_8689);
nor U9207 (N_9207,N_8791,N_8752);
or U9208 (N_9208,N_8470,N_8691);
or U9209 (N_9209,N_8687,N_8254);
nand U9210 (N_9210,N_8913,N_8408);
nor U9211 (N_9211,N_8597,N_8890);
or U9212 (N_9212,N_8444,N_8348);
or U9213 (N_9213,N_8967,N_8856);
nand U9214 (N_9214,N_8328,N_8886);
or U9215 (N_9215,N_8914,N_8287);
nor U9216 (N_9216,N_8960,N_8817);
or U9217 (N_9217,N_8438,N_8539);
nor U9218 (N_9218,N_8974,N_8393);
and U9219 (N_9219,N_8738,N_8279);
and U9220 (N_9220,N_8491,N_8595);
nand U9221 (N_9221,N_8915,N_8493);
xor U9222 (N_9222,N_8776,N_8656);
xor U9223 (N_9223,N_8668,N_8648);
and U9224 (N_9224,N_8357,N_8825);
and U9225 (N_9225,N_8828,N_8418);
nor U9226 (N_9226,N_8615,N_8768);
or U9227 (N_9227,N_8388,N_8337);
nor U9228 (N_9228,N_8878,N_8285);
or U9229 (N_9229,N_8840,N_8253);
or U9230 (N_9230,N_8700,N_8820);
and U9231 (N_9231,N_8460,N_8899);
nand U9232 (N_9232,N_8993,N_8765);
and U9233 (N_9233,N_8567,N_8923);
and U9234 (N_9234,N_8440,N_8780);
xnor U9235 (N_9235,N_8358,N_8478);
and U9236 (N_9236,N_8485,N_8405);
nor U9237 (N_9237,N_8632,N_8259);
and U9238 (N_9238,N_8931,N_8706);
or U9239 (N_9239,N_8763,N_8302);
or U9240 (N_9240,N_8718,N_8639);
nor U9241 (N_9241,N_8858,N_8646);
or U9242 (N_9242,N_8280,N_8375);
nand U9243 (N_9243,N_8369,N_8394);
nor U9244 (N_9244,N_8735,N_8842);
nor U9245 (N_9245,N_8853,N_8517);
or U9246 (N_9246,N_8395,N_8315);
nand U9247 (N_9247,N_8317,N_8737);
and U9248 (N_9248,N_8445,N_8924);
nor U9249 (N_9249,N_8675,N_8414);
nor U9250 (N_9250,N_8957,N_8599);
and U9251 (N_9251,N_8400,N_8771);
nor U9252 (N_9252,N_8389,N_8709);
nand U9253 (N_9253,N_8831,N_8437);
and U9254 (N_9254,N_8958,N_8617);
nand U9255 (N_9255,N_8983,N_8741);
nor U9256 (N_9256,N_8579,N_8381);
and U9257 (N_9257,N_8331,N_8669);
and U9258 (N_9258,N_8667,N_8479);
nor U9259 (N_9259,N_8787,N_8461);
nor U9260 (N_9260,N_8578,N_8431);
nand U9261 (N_9261,N_8384,N_8427);
nand U9262 (N_9262,N_8664,N_8702);
or U9263 (N_9263,N_8636,N_8392);
nand U9264 (N_9264,N_8608,N_8816);
or U9265 (N_9265,N_8575,N_8607);
or U9266 (N_9266,N_8264,N_8604);
xnor U9267 (N_9267,N_8783,N_8359);
or U9268 (N_9268,N_8563,N_8455);
nand U9269 (N_9269,N_8658,N_8995);
nor U9270 (N_9270,N_8704,N_8304);
nor U9271 (N_9271,N_8269,N_8336);
and U9272 (N_9272,N_8726,N_8472);
or U9273 (N_9273,N_8374,N_8969);
or U9274 (N_9274,N_8990,N_8794);
or U9275 (N_9275,N_8716,N_8541);
or U9276 (N_9276,N_8922,N_8696);
nor U9277 (N_9277,N_8531,N_8288);
nor U9278 (N_9278,N_8836,N_8711);
and U9279 (N_9279,N_8725,N_8772);
or U9280 (N_9280,N_8404,N_8920);
or U9281 (N_9281,N_8647,N_8293);
and U9282 (N_9282,N_8398,N_8551);
or U9283 (N_9283,N_8643,N_8409);
nand U9284 (N_9284,N_8367,N_8671);
nor U9285 (N_9285,N_8557,N_8779);
and U9286 (N_9286,N_8797,N_8407);
or U9287 (N_9287,N_8773,N_8666);
nand U9288 (N_9288,N_8864,N_8970);
or U9289 (N_9289,N_8847,N_8720);
and U9290 (N_9290,N_8286,N_8339);
or U9291 (N_9291,N_8333,N_8372);
and U9292 (N_9292,N_8544,N_8386);
and U9293 (N_9293,N_8904,N_8574);
or U9294 (N_9294,N_8547,N_8353);
nor U9295 (N_9295,N_8909,N_8312);
xnor U9296 (N_9296,N_8416,N_8385);
nand U9297 (N_9297,N_8487,N_8723);
nand U9298 (N_9298,N_8564,N_8450);
and U9299 (N_9299,N_8345,N_8587);
nand U9300 (N_9300,N_8623,N_8629);
or U9301 (N_9301,N_8509,N_8402);
nor U9302 (N_9302,N_8576,N_8883);
nor U9303 (N_9303,N_8822,N_8740);
and U9304 (N_9304,N_8761,N_8452);
and U9305 (N_9305,N_8843,N_8274);
and U9306 (N_9306,N_8428,N_8934);
nand U9307 (N_9307,N_8320,N_8683);
nor U9308 (N_9308,N_8762,N_8524);
and U9309 (N_9309,N_8426,N_8819);
xnor U9310 (N_9310,N_8714,N_8855);
and U9311 (N_9311,N_8282,N_8482);
or U9312 (N_9312,N_8717,N_8782);
or U9313 (N_9313,N_8821,N_8927);
and U9314 (N_9314,N_8346,N_8606);
or U9315 (N_9315,N_8419,N_8325);
and U9316 (N_9316,N_8589,N_8748);
or U9317 (N_9317,N_8753,N_8792);
nor U9318 (N_9318,N_8436,N_8695);
or U9319 (N_9319,N_8553,N_8739);
nor U9320 (N_9320,N_8399,N_8745);
or U9321 (N_9321,N_8586,N_8908);
and U9322 (N_9322,N_8314,N_8582);
nand U9323 (N_9323,N_8698,N_8907);
nand U9324 (N_9324,N_8291,N_8968);
nand U9325 (N_9325,N_8570,N_8719);
or U9326 (N_9326,N_8332,N_8866);
nor U9327 (N_9327,N_8905,N_8645);
and U9328 (N_9328,N_8289,N_8457);
or U9329 (N_9329,N_8290,N_8310);
xnor U9330 (N_9330,N_8459,N_8848);
and U9331 (N_9331,N_8680,N_8973);
and U9332 (N_9332,N_8903,N_8940);
and U9333 (N_9333,N_8823,N_8347);
xnor U9334 (N_9334,N_8354,N_8654);
and U9335 (N_9335,N_8996,N_8991);
or U9336 (N_9336,N_8476,N_8732);
and U9337 (N_9337,N_8824,N_8316);
and U9338 (N_9338,N_8548,N_8722);
nor U9339 (N_9339,N_8661,N_8660);
and U9340 (N_9340,N_8614,N_8307);
or U9341 (N_9341,N_8961,N_8880);
and U9342 (N_9342,N_8423,N_8977);
nand U9343 (N_9343,N_8948,N_8448);
and U9344 (N_9344,N_8378,N_8522);
or U9345 (N_9345,N_8556,N_8412);
nor U9346 (N_9346,N_8756,N_8300);
nor U9347 (N_9347,N_8503,N_8921);
and U9348 (N_9348,N_8365,N_8610);
and U9349 (N_9349,N_8982,N_8975);
nand U9350 (N_9350,N_8750,N_8630);
nor U9351 (N_9351,N_8980,N_8350);
and U9352 (N_9352,N_8326,N_8257);
nor U9353 (N_9353,N_8862,N_8537);
or U9354 (N_9354,N_8273,N_8673);
nand U9355 (N_9355,N_8724,N_8590);
or U9356 (N_9356,N_8443,N_8341);
and U9357 (N_9357,N_8406,N_8268);
and U9358 (N_9358,N_8710,N_8271);
or U9359 (N_9359,N_8591,N_8728);
nand U9360 (N_9360,N_8935,N_8826);
and U9361 (N_9361,N_8809,N_8653);
nor U9362 (N_9362,N_8681,N_8662);
nand U9363 (N_9363,N_8736,N_8674);
or U9364 (N_9364,N_8513,N_8693);
or U9365 (N_9365,N_8411,N_8301);
nand U9366 (N_9366,N_8420,N_8837);
xor U9367 (N_9367,N_8573,N_8526);
and U9368 (N_9368,N_8417,N_8627);
nand U9369 (N_9369,N_8603,N_8306);
or U9370 (N_9370,N_8897,N_8507);
or U9371 (N_9371,N_8813,N_8396);
nand U9372 (N_9372,N_8707,N_8581);
nor U9373 (N_9373,N_8484,N_8475);
or U9374 (N_9374,N_8944,N_8256);
xnor U9375 (N_9375,N_8971,N_8890);
and U9376 (N_9376,N_8394,N_8520);
nand U9377 (N_9377,N_8641,N_8984);
and U9378 (N_9378,N_8527,N_8261);
or U9379 (N_9379,N_8935,N_8798);
and U9380 (N_9380,N_8761,N_8536);
nand U9381 (N_9381,N_8702,N_8545);
nand U9382 (N_9382,N_8379,N_8344);
or U9383 (N_9383,N_8448,N_8807);
or U9384 (N_9384,N_8754,N_8281);
nor U9385 (N_9385,N_8765,N_8374);
and U9386 (N_9386,N_8996,N_8695);
nor U9387 (N_9387,N_8752,N_8770);
nand U9388 (N_9388,N_8559,N_8980);
and U9389 (N_9389,N_8385,N_8308);
nor U9390 (N_9390,N_8977,N_8350);
and U9391 (N_9391,N_8620,N_8662);
or U9392 (N_9392,N_8671,N_8877);
or U9393 (N_9393,N_8830,N_8436);
and U9394 (N_9394,N_8681,N_8993);
nor U9395 (N_9395,N_8716,N_8755);
nand U9396 (N_9396,N_8376,N_8557);
and U9397 (N_9397,N_8761,N_8991);
nand U9398 (N_9398,N_8398,N_8288);
or U9399 (N_9399,N_8720,N_8912);
and U9400 (N_9400,N_8438,N_8675);
nand U9401 (N_9401,N_8961,N_8577);
or U9402 (N_9402,N_8973,N_8374);
nand U9403 (N_9403,N_8952,N_8931);
nand U9404 (N_9404,N_8837,N_8697);
nand U9405 (N_9405,N_8337,N_8508);
nand U9406 (N_9406,N_8410,N_8588);
and U9407 (N_9407,N_8845,N_8928);
or U9408 (N_9408,N_8332,N_8583);
nor U9409 (N_9409,N_8626,N_8858);
nand U9410 (N_9410,N_8730,N_8538);
nand U9411 (N_9411,N_8597,N_8319);
or U9412 (N_9412,N_8468,N_8544);
and U9413 (N_9413,N_8277,N_8614);
nand U9414 (N_9414,N_8350,N_8688);
or U9415 (N_9415,N_8823,N_8704);
nand U9416 (N_9416,N_8699,N_8798);
or U9417 (N_9417,N_8393,N_8481);
or U9418 (N_9418,N_8769,N_8668);
and U9419 (N_9419,N_8720,N_8505);
nor U9420 (N_9420,N_8781,N_8520);
nor U9421 (N_9421,N_8822,N_8953);
nand U9422 (N_9422,N_8734,N_8712);
nor U9423 (N_9423,N_8698,N_8688);
nor U9424 (N_9424,N_8416,N_8524);
or U9425 (N_9425,N_8303,N_8594);
nor U9426 (N_9426,N_8971,N_8348);
and U9427 (N_9427,N_8970,N_8569);
and U9428 (N_9428,N_8843,N_8747);
nor U9429 (N_9429,N_8330,N_8743);
and U9430 (N_9430,N_8615,N_8545);
nand U9431 (N_9431,N_8778,N_8947);
and U9432 (N_9432,N_8823,N_8402);
nor U9433 (N_9433,N_8890,N_8438);
or U9434 (N_9434,N_8588,N_8908);
nand U9435 (N_9435,N_8860,N_8687);
and U9436 (N_9436,N_8754,N_8366);
nor U9437 (N_9437,N_8358,N_8406);
or U9438 (N_9438,N_8721,N_8449);
nor U9439 (N_9439,N_8574,N_8261);
and U9440 (N_9440,N_8418,N_8587);
and U9441 (N_9441,N_8291,N_8520);
and U9442 (N_9442,N_8319,N_8692);
nand U9443 (N_9443,N_8588,N_8989);
or U9444 (N_9444,N_8905,N_8336);
nor U9445 (N_9445,N_8803,N_8775);
and U9446 (N_9446,N_8251,N_8746);
and U9447 (N_9447,N_8496,N_8629);
and U9448 (N_9448,N_8774,N_8818);
nor U9449 (N_9449,N_8899,N_8821);
nor U9450 (N_9450,N_8346,N_8702);
or U9451 (N_9451,N_8605,N_8440);
and U9452 (N_9452,N_8955,N_8988);
and U9453 (N_9453,N_8959,N_8631);
or U9454 (N_9454,N_8895,N_8763);
or U9455 (N_9455,N_8894,N_8539);
nor U9456 (N_9456,N_8641,N_8868);
or U9457 (N_9457,N_8798,N_8431);
nand U9458 (N_9458,N_8910,N_8962);
nand U9459 (N_9459,N_8367,N_8460);
nand U9460 (N_9460,N_8722,N_8525);
nor U9461 (N_9461,N_8497,N_8594);
nand U9462 (N_9462,N_8418,N_8605);
and U9463 (N_9463,N_8986,N_8766);
nand U9464 (N_9464,N_8362,N_8445);
and U9465 (N_9465,N_8797,N_8307);
nand U9466 (N_9466,N_8338,N_8618);
nor U9467 (N_9467,N_8978,N_8523);
nor U9468 (N_9468,N_8343,N_8357);
or U9469 (N_9469,N_8556,N_8636);
nand U9470 (N_9470,N_8322,N_8436);
and U9471 (N_9471,N_8424,N_8591);
nand U9472 (N_9472,N_8488,N_8433);
and U9473 (N_9473,N_8450,N_8786);
nor U9474 (N_9474,N_8932,N_8561);
or U9475 (N_9475,N_8401,N_8770);
nor U9476 (N_9476,N_8367,N_8881);
nand U9477 (N_9477,N_8571,N_8881);
and U9478 (N_9478,N_8574,N_8455);
nand U9479 (N_9479,N_8722,N_8970);
or U9480 (N_9480,N_8354,N_8542);
or U9481 (N_9481,N_8371,N_8681);
nand U9482 (N_9482,N_8323,N_8466);
nor U9483 (N_9483,N_8931,N_8886);
nand U9484 (N_9484,N_8747,N_8716);
and U9485 (N_9485,N_8725,N_8849);
nor U9486 (N_9486,N_8261,N_8850);
or U9487 (N_9487,N_8372,N_8347);
or U9488 (N_9488,N_8309,N_8264);
nand U9489 (N_9489,N_8547,N_8521);
and U9490 (N_9490,N_8999,N_8752);
nor U9491 (N_9491,N_8270,N_8899);
or U9492 (N_9492,N_8736,N_8338);
nor U9493 (N_9493,N_8279,N_8533);
and U9494 (N_9494,N_8837,N_8726);
or U9495 (N_9495,N_8757,N_8462);
nor U9496 (N_9496,N_8380,N_8363);
and U9497 (N_9497,N_8315,N_8530);
nand U9498 (N_9498,N_8665,N_8593);
and U9499 (N_9499,N_8579,N_8670);
or U9500 (N_9500,N_8416,N_8660);
nor U9501 (N_9501,N_8901,N_8595);
nand U9502 (N_9502,N_8578,N_8474);
or U9503 (N_9503,N_8345,N_8543);
nand U9504 (N_9504,N_8550,N_8733);
or U9505 (N_9505,N_8286,N_8290);
nor U9506 (N_9506,N_8377,N_8437);
nand U9507 (N_9507,N_8936,N_8599);
nand U9508 (N_9508,N_8609,N_8472);
or U9509 (N_9509,N_8801,N_8750);
and U9510 (N_9510,N_8566,N_8435);
and U9511 (N_9511,N_8625,N_8912);
nor U9512 (N_9512,N_8817,N_8271);
and U9513 (N_9513,N_8736,N_8462);
and U9514 (N_9514,N_8406,N_8555);
nand U9515 (N_9515,N_8910,N_8694);
and U9516 (N_9516,N_8355,N_8698);
nand U9517 (N_9517,N_8892,N_8479);
and U9518 (N_9518,N_8526,N_8925);
and U9519 (N_9519,N_8398,N_8289);
or U9520 (N_9520,N_8537,N_8752);
nor U9521 (N_9521,N_8667,N_8736);
xor U9522 (N_9522,N_8459,N_8605);
nand U9523 (N_9523,N_8571,N_8967);
or U9524 (N_9524,N_8292,N_8268);
or U9525 (N_9525,N_8880,N_8996);
and U9526 (N_9526,N_8544,N_8510);
nor U9527 (N_9527,N_8806,N_8795);
and U9528 (N_9528,N_8279,N_8335);
and U9529 (N_9529,N_8655,N_8893);
nor U9530 (N_9530,N_8929,N_8952);
and U9531 (N_9531,N_8532,N_8904);
nor U9532 (N_9532,N_8957,N_8550);
nand U9533 (N_9533,N_8535,N_8767);
nand U9534 (N_9534,N_8772,N_8370);
nand U9535 (N_9535,N_8939,N_8868);
and U9536 (N_9536,N_8638,N_8636);
nand U9537 (N_9537,N_8325,N_8838);
nor U9538 (N_9538,N_8281,N_8683);
or U9539 (N_9539,N_8702,N_8999);
or U9540 (N_9540,N_8380,N_8924);
nor U9541 (N_9541,N_8255,N_8679);
nor U9542 (N_9542,N_8597,N_8994);
nand U9543 (N_9543,N_8561,N_8417);
and U9544 (N_9544,N_8709,N_8955);
xnor U9545 (N_9545,N_8885,N_8890);
and U9546 (N_9546,N_8607,N_8888);
or U9547 (N_9547,N_8459,N_8830);
nand U9548 (N_9548,N_8600,N_8347);
or U9549 (N_9549,N_8608,N_8279);
or U9550 (N_9550,N_8702,N_8368);
nand U9551 (N_9551,N_8981,N_8717);
nor U9552 (N_9552,N_8443,N_8283);
or U9553 (N_9553,N_8712,N_8831);
or U9554 (N_9554,N_8692,N_8304);
nor U9555 (N_9555,N_8757,N_8312);
or U9556 (N_9556,N_8702,N_8704);
or U9557 (N_9557,N_8973,N_8942);
nand U9558 (N_9558,N_8625,N_8929);
nand U9559 (N_9559,N_8448,N_8809);
or U9560 (N_9560,N_8777,N_8935);
nand U9561 (N_9561,N_8891,N_8374);
and U9562 (N_9562,N_8702,N_8580);
and U9563 (N_9563,N_8717,N_8677);
nand U9564 (N_9564,N_8330,N_8672);
nand U9565 (N_9565,N_8874,N_8263);
and U9566 (N_9566,N_8774,N_8895);
or U9567 (N_9567,N_8932,N_8496);
and U9568 (N_9568,N_8401,N_8672);
nand U9569 (N_9569,N_8800,N_8539);
nand U9570 (N_9570,N_8500,N_8354);
nand U9571 (N_9571,N_8950,N_8785);
and U9572 (N_9572,N_8679,N_8266);
and U9573 (N_9573,N_8254,N_8957);
or U9574 (N_9574,N_8859,N_8668);
and U9575 (N_9575,N_8499,N_8322);
nand U9576 (N_9576,N_8438,N_8563);
or U9577 (N_9577,N_8735,N_8856);
and U9578 (N_9578,N_8845,N_8277);
and U9579 (N_9579,N_8682,N_8294);
or U9580 (N_9580,N_8816,N_8790);
nand U9581 (N_9581,N_8719,N_8741);
and U9582 (N_9582,N_8967,N_8662);
or U9583 (N_9583,N_8931,N_8766);
or U9584 (N_9584,N_8657,N_8534);
or U9585 (N_9585,N_8737,N_8748);
and U9586 (N_9586,N_8478,N_8740);
and U9587 (N_9587,N_8427,N_8587);
or U9588 (N_9588,N_8847,N_8673);
nor U9589 (N_9589,N_8911,N_8681);
and U9590 (N_9590,N_8798,N_8718);
or U9591 (N_9591,N_8960,N_8658);
or U9592 (N_9592,N_8405,N_8980);
and U9593 (N_9593,N_8947,N_8580);
nand U9594 (N_9594,N_8492,N_8713);
nor U9595 (N_9595,N_8520,N_8451);
or U9596 (N_9596,N_8890,N_8561);
nand U9597 (N_9597,N_8977,N_8955);
or U9598 (N_9598,N_8299,N_8476);
or U9599 (N_9599,N_8677,N_8387);
and U9600 (N_9600,N_8787,N_8755);
nor U9601 (N_9601,N_8889,N_8954);
or U9602 (N_9602,N_8264,N_8402);
or U9603 (N_9603,N_8912,N_8755);
nand U9604 (N_9604,N_8991,N_8455);
and U9605 (N_9605,N_8918,N_8765);
or U9606 (N_9606,N_8705,N_8937);
or U9607 (N_9607,N_8811,N_8910);
nor U9608 (N_9608,N_8323,N_8494);
nor U9609 (N_9609,N_8667,N_8962);
nand U9610 (N_9610,N_8879,N_8815);
nand U9611 (N_9611,N_8921,N_8406);
and U9612 (N_9612,N_8850,N_8290);
or U9613 (N_9613,N_8605,N_8404);
or U9614 (N_9614,N_8546,N_8328);
nor U9615 (N_9615,N_8393,N_8874);
and U9616 (N_9616,N_8595,N_8268);
or U9617 (N_9617,N_8828,N_8680);
or U9618 (N_9618,N_8377,N_8804);
and U9619 (N_9619,N_8304,N_8609);
xor U9620 (N_9620,N_8725,N_8494);
nand U9621 (N_9621,N_8784,N_8816);
or U9622 (N_9622,N_8619,N_8940);
nor U9623 (N_9623,N_8266,N_8567);
or U9624 (N_9624,N_8436,N_8888);
and U9625 (N_9625,N_8514,N_8824);
or U9626 (N_9626,N_8585,N_8810);
and U9627 (N_9627,N_8905,N_8368);
nor U9628 (N_9628,N_8283,N_8415);
nor U9629 (N_9629,N_8335,N_8871);
nand U9630 (N_9630,N_8987,N_8933);
nand U9631 (N_9631,N_8674,N_8334);
and U9632 (N_9632,N_8966,N_8728);
nand U9633 (N_9633,N_8590,N_8372);
or U9634 (N_9634,N_8308,N_8988);
and U9635 (N_9635,N_8609,N_8319);
or U9636 (N_9636,N_8665,N_8548);
nor U9637 (N_9637,N_8740,N_8940);
nand U9638 (N_9638,N_8712,N_8914);
and U9639 (N_9639,N_8826,N_8792);
nand U9640 (N_9640,N_8494,N_8270);
and U9641 (N_9641,N_8802,N_8690);
nor U9642 (N_9642,N_8974,N_8986);
and U9643 (N_9643,N_8262,N_8758);
and U9644 (N_9644,N_8392,N_8603);
nand U9645 (N_9645,N_8355,N_8805);
and U9646 (N_9646,N_8395,N_8984);
or U9647 (N_9647,N_8491,N_8274);
or U9648 (N_9648,N_8390,N_8577);
or U9649 (N_9649,N_8934,N_8300);
nand U9650 (N_9650,N_8608,N_8957);
and U9651 (N_9651,N_8393,N_8345);
nor U9652 (N_9652,N_8258,N_8284);
and U9653 (N_9653,N_8645,N_8835);
nand U9654 (N_9654,N_8269,N_8492);
nor U9655 (N_9655,N_8813,N_8737);
nor U9656 (N_9656,N_8633,N_8621);
nand U9657 (N_9657,N_8766,N_8397);
nand U9658 (N_9658,N_8293,N_8935);
and U9659 (N_9659,N_8726,N_8697);
and U9660 (N_9660,N_8656,N_8273);
or U9661 (N_9661,N_8626,N_8424);
nor U9662 (N_9662,N_8586,N_8522);
and U9663 (N_9663,N_8547,N_8902);
nor U9664 (N_9664,N_8433,N_8364);
nand U9665 (N_9665,N_8672,N_8699);
nand U9666 (N_9666,N_8891,N_8627);
nand U9667 (N_9667,N_8500,N_8804);
nor U9668 (N_9668,N_8321,N_8978);
or U9669 (N_9669,N_8612,N_8295);
and U9670 (N_9670,N_8776,N_8317);
nand U9671 (N_9671,N_8857,N_8841);
or U9672 (N_9672,N_8334,N_8385);
nand U9673 (N_9673,N_8984,N_8553);
or U9674 (N_9674,N_8315,N_8938);
nor U9675 (N_9675,N_8476,N_8753);
nand U9676 (N_9676,N_8264,N_8693);
or U9677 (N_9677,N_8404,N_8319);
nand U9678 (N_9678,N_8562,N_8677);
nor U9679 (N_9679,N_8308,N_8388);
nor U9680 (N_9680,N_8601,N_8551);
and U9681 (N_9681,N_8476,N_8527);
nand U9682 (N_9682,N_8905,N_8404);
nand U9683 (N_9683,N_8907,N_8815);
nand U9684 (N_9684,N_8395,N_8501);
and U9685 (N_9685,N_8724,N_8883);
and U9686 (N_9686,N_8323,N_8968);
and U9687 (N_9687,N_8938,N_8681);
nand U9688 (N_9688,N_8352,N_8415);
nand U9689 (N_9689,N_8583,N_8850);
or U9690 (N_9690,N_8473,N_8461);
or U9691 (N_9691,N_8493,N_8833);
nand U9692 (N_9692,N_8437,N_8523);
and U9693 (N_9693,N_8303,N_8936);
nor U9694 (N_9694,N_8927,N_8747);
nand U9695 (N_9695,N_8918,N_8383);
and U9696 (N_9696,N_8687,N_8707);
or U9697 (N_9697,N_8924,N_8618);
nand U9698 (N_9698,N_8464,N_8358);
nor U9699 (N_9699,N_8697,N_8292);
nor U9700 (N_9700,N_8726,N_8260);
or U9701 (N_9701,N_8326,N_8280);
xor U9702 (N_9702,N_8578,N_8965);
nor U9703 (N_9703,N_8861,N_8478);
nor U9704 (N_9704,N_8557,N_8392);
nand U9705 (N_9705,N_8991,N_8783);
and U9706 (N_9706,N_8276,N_8881);
or U9707 (N_9707,N_8779,N_8864);
nand U9708 (N_9708,N_8826,N_8837);
nand U9709 (N_9709,N_8411,N_8720);
nand U9710 (N_9710,N_8995,N_8461);
and U9711 (N_9711,N_8330,N_8366);
or U9712 (N_9712,N_8998,N_8683);
and U9713 (N_9713,N_8451,N_8638);
and U9714 (N_9714,N_8342,N_8830);
nand U9715 (N_9715,N_8808,N_8694);
nand U9716 (N_9716,N_8251,N_8634);
nand U9717 (N_9717,N_8713,N_8594);
nor U9718 (N_9718,N_8814,N_8937);
or U9719 (N_9719,N_8295,N_8888);
nor U9720 (N_9720,N_8479,N_8598);
and U9721 (N_9721,N_8939,N_8903);
nor U9722 (N_9722,N_8600,N_8579);
and U9723 (N_9723,N_8458,N_8381);
nor U9724 (N_9724,N_8789,N_8909);
nor U9725 (N_9725,N_8599,N_8357);
nand U9726 (N_9726,N_8952,N_8702);
nand U9727 (N_9727,N_8397,N_8396);
nor U9728 (N_9728,N_8515,N_8555);
nand U9729 (N_9729,N_8345,N_8284);
and U9730 (N_9730,N_8718,N_8902);
or U9731 (N_9731,N_8955,N_8975);
and U9732 (N_9732,N_8701,N_8837);
nor U9733 (N_9733,N_8430,N_8340);
or U9734 (N_9734,N_8776,N_8990);
nand U9735 (N_9735,N_8355,N_8296);
nor U9736 (N_9736,N_8600,N_8639);
nor U9737 (N_9737,N_8299,N_8365);
and U9738 (N_9738,N_8815,N_8392);
or U9739 (N_9739,N_8489,N_8266);
and U9740 (N_9740,N_8637,N_8864);
or U9741 (N_9741,N_8320,N_8875);
or U9742 (N_9742,N_8653,N_8934);
nor U9743 (N_9743,N_8932,N_8253);
nor U9744 (N_9744,N_8347,N_8719);
nor U9745 (N_9745,N_8659,N_8988);
nand U9746 (N_9746,N_8916,N_8461);
nand U9747 (N_9747,N_8826,N_8724);
nand U9748 (N_9748,N_8989,N_8277);
and U9749 (N_9749,N_8577,N_8335);
or U9750 (N_9750,N_9062,N_9679);
or U9751 (N_9751,N_9100,N_9708);
or U9752 (N_9752,N_9613,N_9334);
nor U9753 (N_9753,N_9279,N_9236);
nor U9754 (N_9754,N_9030,N_9588);
and U9755 (N_9755,N_9352,N_9194);
nor U9756 (N_9756,N_9168,N_9022);
nand U9757 (N_9757,N_9654,N_9589);
nor U9758 (N_9758,N_9649,N_9535);
and U9759 (N_9759,N_9544,N_9372);
or U9760 (N_9760,N_9726,N_9046);
or U9761 (N_9761,N_9149,N_9554);
nand U9762 (N_9762,N_9434,N_9411);
and U9763 (N_9763,N_9531,N_9447);
or U9764 (N_9764,N_9154,N_9604);
and U9765 (N_9765,N_9347,N_9387);
nand U9766 (N_9766,N_9078,N_9650);
or U9767 (N_9767,N_9182,N_9438);
and U9768 (N_9768,N_9227,N_9312);
or U9769 (N_9769,N_9349,N_9647);
nor U9770 (N_9770,N_9048,N_9306);
or U9771 (N_9771,N_9222,N_9590);
nor U9772 (N_9772,N_9692,N_9664);
or U9773 (N_9773,N_9052,N_9500);
nand U9774 (N_9774,N_9158,N_9415);
nor U9775 (N_9775,N_9666,N_9711);
nand U9776 (N_9776,N_9580,N_9719);
nand U9777 (N_9777,N_9739,N_9059);
nand U9778 (N_9778,N_9697,N_9574);
or U9779 (N_9779,N_9422,N_9437);
or U9780 (N_9780,N_9656,N_9319);
nand U9781 (N_9781,N_9218,N_9350);
nand U9782 (N_9782,N_9360,N_9569);
or U9783 (N_9783,N_9346,N_9088);
or U9784 (N_9784,N_9110,N_9672);
and U9785 (N_9785,N_9459,N_9506);
nand U9786 (N_9786,N_9691,N_9491);
nor U9787 (N_9787,N_9611,N_9746);
nor U9788 (N_9788,N_9577,N_9733);
nand U9789 (N_9789,N_9004,N_9181);
or U9790 (N_9790,N_9307,N_9639);
or U9791 (N_9791,N_9548,N_9384);
and U9792 (N_9792,N_9712,N_9495);
nor U9793 (N_9793,N_9038,N_9083);
and U9794 (N_9794,N_9351,N_9745);
and U9795 (N_9795,N_9573,N_9282);
or U9796 (N_9796,N_9278,N_9359);
nor U9797 (N_9797,N_9061,N_9419);
and U9798 (N_9798,N_9435,N_9338);
and U9799 (N_9799,N_9426,N_9680);
nor U9800 (N_9800,N_9157,N_9348);
and U9801 (N_9801,N_9003,N_9525);
and U9802 (N_9802,N_9231,N_9208);
nor U9803 (N_9803,N_9190,N_9578);
nand U9804 (N_9804,N_9114,N_9657);
nor U9805 (N_9805,N_9295,N_9374);
nor U9806 (N_9806,N_9311,N_9095);
nand U9807 (N_9807,N_9209,N_9166);
or U9808 (N_9808,N_9509,N_9188);
nor U9809 (N_9809,N_9695,N_9183);
and U9810 (N_9810,N_9392,N_9555);
and U9811 (N_9811,N_9394,N_9628);
nor U9812 (N_9812,N_9738,N_9047);
nor U9813 (N_9813,N_9579,N_9210);
or U9814 (N_9814,N_9482,N_9385);
or U9815 (N_9815,N_9550,N_9517);
nor U9816 (N_9816,N_9538,N_9226);
and U9817 (N_9817,N_9057,N_9451);
nor U9818 (N_9818,N_9725,N_9174);
nor U9819 (N_9819,N_9536,N_9532);
nor U9820 (N_9820,N_9335,N_9373);
or U9821 (N_9821,N_9136,N_9693);
nand U9822 (N_9822,N_9082,N_9406);
or U9823 (N_9823,N_9009,N_9309);
and U9824 (N_9824,N_9741,N_9408);
or U9825 (N_9825,N_9169,N_9262);
and U9826 (N_9826,N_9595,N_9642);
nand U9827 (N_9827,N_9742,N_9717);
nor U9828 (N_9828,N_9050,N_9248);
and U9829 (N_9829,N_9185,N_9571);
and U9830 (N_9830,N_9337,N_9594);
nor U9831 (N_9831,N_9698,N_9005);
and U9832 (N_9832,N_9681,N_9553);
nand U9833 (N_9833,N_9133,N_9081);
nand U9834 (N_9834,N_9146,N_9107);
or U9835 (N_9835,N_9453,N_9101);
nand U9836 (N_9836,N_9494,N_9161);
and U9837 (N_9837,N_9559,N_9006);
nand U9838 (N_9838,N_9035,N_9125);
and U9839 (N_9839,N_9292,N_9540);
nand U9840 (N_9840,N_9720,N_9123);
nand U9841 (N_9841,N_9497,N_9683);
nor U9842 (N_9842,N_9477,N_9106);
or U9843 (N_9843,N_9630,N_9070);
and U9844 (N_9844,N_9034,N_9000);
nor U9845 (N_9845,N_9322,N_9448);
or U9846 (N_9846,N_9180,N_9514);
or U9847 (N_9847,N_9736,N_9016);
and U9848 (N_9848,N_9220,N_9029);
and U9849 (N_9849,N_9598,N_9714);
nor U9850 (N_9850,N_9466,N_9685);
nor U9851 (N_9851,N_9033,N_9670);
nand U9852 (N_9852,N_9010,N_9245);
and U9853 (N_9853,N_9018,N_9480);
nand U9854 (N_9854,N_9336,N_9584);
and U9855 (N_9855,N_9327,N_9195);
or U9856 (N_9856,N_9472,N_9205);
or U9857 (N_9857,N_9104,N_9283);
or U9858 (N_9858,N_9244,N_9249);
nor U9859 (N_9859,N_9199,N_9476);
nand U9860 (N_9860,N_9475,N_9660);
or U9861 (N_9861,N_9743,N_9333);
or U9862 (N_9862,N_9483,N_9706);
nand U9863 (N_9863,N_9663,N_9017);
nand U9864 (N_9864,N_9400,N_9313);
and U9865 (N_9865,N_9456,N_9446);
nand U9866 (N_9866,N_9528,N_9069);
nand U9867 (N_9867,N_9324,N_9031);
and U9868 (N_9868,N_9441,N_9102);
xnor U9869 (N_9869,N_9063,N_9671);
nand U9870 (N_9870,N_9653,N_9658);
nor U9871 (N_9871,N_9417,N_9357);
nand U9872 (N_9872,N_9390,N_9533);
and U9873 (N_9873,N_9583,N_9235);
and U9874 (N_9874,N_9457,N_9523);
or U9875 (N_9875,N_9071,N_9191);
and U9876 (N_9876,N_9399,N_9382);
nand U9877 (N_9877,N_9619,N_9354);
nand U9878 (N_9878,N_9330,N_9305);
nand U9879 (N_9879,N_9566,N_9055);
nand U9880 (N_9880,N_9585,N_9316);
nor U9881 (N_9881,N_9513,N_9014);
and U9882 (N_9882,N_9694,N_9187);
or U9883 (N_9883,N_9460,N_9037);
and U9884 (N_9884,N_9612,N_9287);
and U9885 (N_9885,N_9511,N_9730);
nor U9886 (N_9886,N_9703,N_9586);
and U9887 (N_9887,N_9290,N_9223);
and U9888 (N_9888,N_9304,N_9512);
nor U9889 (N_9889,N_9458,N_9370);
or U9890 (N_9890,N_9433,N_9469);
nor U9891 (N_9891,N_9369,N_9464);
nand U9892 (N_9892,N_9302,N_9315);
and U9893 (N_9893,N_9635,N_9073);
or U9894 (N_9894,N_9049,N_9124);
and U9895 (N_9895,N_9644,N_9353);
and U9896 (N_9896,N_9380,N_9054);
nor U9897 (N_9897,N_9428,N_9496);
or U9898 (N_9898,N_9643,N_9277);
nor U9899 (N_9899,N_9443,N_9655);
and U9900 (N_9900,N_9255,N_9170);
and U9901 (N_9901,N_9117,N_9682);
or U9902 (N_9902,N_9620,N_9572);
or U9903 (N_9903,N_9651,N_9213);
and U9904 (N_9904,N_9724,N_9257);
nor U9905 (N_9905,N_9558,N_9616);
nand U9906 (N_9906,N_9293,N_9045);
and U9907 (N_9907,N_9246,N_9138);
nand U9908 (N_9908,N_9631,N_9383);
and U9909 (N_9909,N_9131,N_9515);
and U9910 (N_9910,N_9109,N_9240);
or U9911 (N_9911,N_9317,N_9020);
nor U9912 (N_9912,N_9075,N_9575);
and U9913 (N_9913,N_9111,N_9086);
or U9914 (N_9914,N_9707,N_9701);
and U9915 (N_9915,N_9108,N_9596);
and U9916 (N_9916,N_9524,N_9427);
nand U9917 (N_9917,N_9486,N_9715);
nand U9918 (N_9918,N_9404,N_9299);
nand U9919 (N_9919,N_9710,N_9044);
nand U9920 (N_9920,N_9025,N_9260);
nor U9921 (N_9921,N_9012,N_9144);
or U9922 (N_9922,N_9264,N_9310);
nand U9923 (N_9923,N_9709,N_9247);
nor U9924 (N_9924,N_9160,N_9243);
nor U9925 (N_9925,N_9275,N_9557);
or U9926 (N_9926,N_9068,N_9207);
and U9927 (N_9927,N_9675,N_9627);
nand U9928 (N_9928,N_9423,N_9470);
and U9929 (N_9929,N_9058,N_9405);
and U9930 (N_9930,N_9242,N_9652);
nand U9931 (N_9931,N_9605,N_9623);
and U9932 (N_9932,N_9172,N_9677);
nand U9933 (N_9933,N_9186,N_9219);
or U9934 (N_9934,N_9269,N_9542);
and U9935 (N_9935,N_9228,N_9455);
and U9936 (N_9936,N_9371,N_9375);
or U9937 (N_9937,N_9066,N_9547);
and U9938 (N_9938,N_9601,N_9060);
and U9939 (N_9939,N_9122,N_9481);
nand U9940 (N_9940,N_9197,N_9378);
nand U9941 (N_9941,N_9291,N_9702);
xnor U9942 (N_9942,N_9274,N_9252);
and U9943 (N_9943,N_9501,N_9502);
or U9944 (N_9944,N_9318,N_9521);
nor U9945 (N_9945,N_9718,N_9173);
nand U9946 (N_9946,N_9668,N_9254);
or U9947 (N_9947,N_9148,N_9238);
or U9948 (N_9948,N_9155,N_9356);
nor U9949 (N_9949,N_9080,N_9622);
nor U9950 (N_9950,N_9728,N_9265);
nor U9951 (N_9951,N_9273,N_9416);
nand U9952 (N_9952,N_9332,N_9401);
nor U9953 (N_9953,N_9699,N_9688);
nand U9954 (N_9954,N_9606,N_9549);
nor U9955 (N_9955,N_9039,N_9567);
nand U9956 (N_9956,N_9637,N_9722);
and U9957 (N_9957,N_9576,N_9256);
nor U9958 (N_9958,N_9429,N_9281);
nand U9959 (N_9959,N_9216,N_9345);
or U9960 (N_9960,N_9323,N_9505);
nand U9961 (N_9961,N_9503,N_9740);
nor U9962 (N_9962,N_9115,N_9541);
nor U9963 (N_9963,N_9492,N_9266);
nand U9964 (N_9964,N_9676,N_9632);
or U9965 (N_9965,N_9700,N_9539);
nand U9966 (N_9966,N_9355,N_9167);
nor U9967 (N_9967,N_9599,N_9179);
nand U9968 (N_9968,N_9690,N_9648);
nor U9969 (N_9969,N_9217,N_9203);
or U9970 (N_9970,N_9189,N_9530);
and U9971 (N_9971,N_9036,N_9563);
and U9972 (N_9972,N_9396,N_9079);
or U9973 (N_9973,N_9461,N_9546);
nor U9974 (N_9974,N_9625,N_9381);
and U9975 (N_9975,N_9468,N_9289);
nor U9976 (N_9976,N_9450,N_9723);
nor U9977 (N_9977,N_9271,N_9420);
and U9978 (N_9978,N_9713,N_9128);
nor U9979 (N_9979,N_9177,N_9561);
or U9980 (N_9980,N_9621,N_9072);
or U9981 (N_9981,N_9151,N_9617);
nand U9982 (N_9982,N_9032,N_9667);
nand U9983 (N_9983,N_9471,N_9522);
nand U9984 (N_9984,N_9041,N_9259);
and U9985 (N_9985,N_9484,N_9178);
or U9986 (N_9986,N_9552,N_9640);
and U9987 (N_9987,N_9234,N_9403);
nand U9988 (N_9988,N_9118,N_9184);
and U9989 (N_9989,N_9564,N_9444);
nand U9990 (N_9990,N_9294,N_9200);
or U9991 (N_9991,N_9325,N_9737);
nand U9992 (N_9992,N_9593,N_9092);
nor U9993 (N_9993,N_9363,N_9286);
or U9994 (N_9994,N_9196,N_9142);
or U9995 (N_9995,N_9303,N_9343);
nand U9996 (N_9996,N_9376,N_9734);
nand U9997 (N_9997,N_9721,N_9232);
nand U9998 (N_9998,N_9641,N_9626);
nand U9999 (N_9999,N_9421,N_9253);
and U10000 (N_10000,N_9087,N_9534);
nor U10001 (N_10001,N_9581,N_9013);
nand U10002 (N_10002,N_9366,N_9418);
nor U10003 (N_10003,N_9090,N_9089);
nor U10004 (N_10004,N_9145,N_9143);
or U10005 (N_10005,N_9120,N_9076);
or U10006 (N_10006,N_9085,N_9397);
nand U10007 (N_10007,N_9665,N_9452);
or U10008 (N_10008,N_9462,N_9021);
and U10009 (N_10009,N_9565,N_9056);
nand U10010 (N_10010,N_9233,N_9225);
and U10011 (N_10011,N_9206,N_9467);
nand U10012 (N_10012,N_9103,N_9308);
nand U10013 (N_10013,N_9127,N_9440);
or U10014 (N_10014,N_9430,N_9051);
or U10015 (N_10015,N_9026,N_9395);
and U10016 (N_10016,N_9749,N_9105);
nand U10017 (N_10017,N_9093,N_9704);
nor U10018 (N_10018,N_9171,N_9673);
nand U10019 (N_10019,N_9687,N_9053);
nand U10020 (N_10020,N_9272,N_9431);
and U10021 (N_10021,N_9602,N_9696);
nor U10022 (N_10022,N_9529,N_9727);
and U10023 (N_10023,N_9153,N_9600);
and U10024 (N_10024,N_9362,N_9748);
nor U10025 (N_10025,N_9498,N_9597);
nand U10026 (N_10026,N_9019,N_9340);
or U10027 (N_10027,N_9001,N_9258);
nand U10028 (N_10028,N_9008,N_9084);
and U10029 (N_10029,N_9570,N_9393);
nand U10030 (N_10030,N_9493,N_9636);
and U10031 (N_10031,N_9152,N_9659);
and U10032 (N_10032,N_9744,N_9121);
or U10033 (N_10033,N_9402,N_9268);
or U10034 (N_10034,N_9465,N_9474);
and U10035 (N_10035,N_9424,N_9662);
and U10036 (N_10036,N_9377,N_9119);
nor U10037 (N_10037,N_9747,N_9686);
nor U10038 (N_10038,N_9365,N_9661);
nor U10039 (N_10039,N_9328,N_9388);
and U10040 (N_10040,N_9398,N_9147);
and U10041 (N_10041,N_9214,N_9568);
and U10042 (N_10042,N_9634,N_9389);
nor U10043 (N_10043,N_9545,N_9267);
xor U10044 (N_10044,N_9684,N_9094);
or U10045 (N_10045,N_9301,N_9096);
and U10046 (N_10046,N_9716,N_9674);
nor U10047 (N_10047,N_9331,N_9410);
xor U10048 (N_10048,N_9358,N_9270);
nand U10049 (N_10049,N_9150,N_9134);
nand U10050 (N_10050,N_9463,N_9591);
nand U10051 (N_10051,N_9510,N_9519);
or U10052 (N_10052,N_9043,N_9202);
nor U10053 (N_10053,N_9141,N_9229);
or U10054 (N_10054,N_9162,N_9449);
nor U10055 (N_10055,N_9067,N_9615);
nand U10056 (N_10056,N_9250,N_9263);
xor U10057 (N_10057,N_9156,N_9064);
nand U10058 (N_10058,N_9163,N_9646);
nand U10059 (N_10059,N_9645,N_9298);
nor U10060 (N_10060,N_9139,N_9024);
and U10061 (N_10061,N_9488,N_9413);
or U10062 (N_10062,N_9490,N_9140);
and U10063 (N_10063,N_9516,N_9543);
and U10064 (N_10064,N_9074,N_9425);
nor U10065 (N_10065,N_9002,N_9116);
nor U10066 (N_10066,N_9176,N_9241);
or U10067 (N_10067,N_9237,N_9551);
nand U10068 (N_10068,N_9499,N_9409);
nand U10069 (N_10069,N_9669,N_9113);
or U10070 (N_10070,N_9386,N_9098);
nand U10071 (N_10071,N_9638,N_9344);
nand U10072 (N_10072,N_9454,N_9284);
nor U10073 (N_10073,N_9379,N_9520);
nand U10074 (N_10074,N_9230,N_9099);
or U10075 (N_10075,N_9341,N_9339);
or U10076 (N_10076,N_9091,N_9097);
and U10077 (N_10077,N_9473,N_9368);
nor U10078 (N_10078,N_9436,N_9624);
nor U10079 (N_10079,N_9023,N_9129);
and U10080 (N_10080,N_9508,N_9285);
nor U10081 (N_10081,N_9175,N_9633);
and U10082 (N_10082,N_9112,N_9261);
or U10083 (N_10083,N_9560,N_9582);
nor U10084 (N_10084,N_9007,N_9489);
or U10085 (N_10085,N_9592,N_9159);
or U10086 (N_10086,N_9537,N_9485);
and U10087 (N_10087,N_9126,N_9300);
nor U10088 (N_10088,N_9526,N_9280);
nand U10089 (N_10089,N_9608,N_9439);
and U10090 (N_10090,N_9732,N_9132);
nand U10091 (N_10091,N_9367,N_9297);
nor U10092 (N_10092,N_9296,N_9027);
nand U10093 (N_10093,N_9678,N_9705);
or U10094 (N_10094,N_9204,N_9556);
and U10095 (N_10095,N_9239,N_9212);
and U10096 (N_10096,N_9042,N_9314);
nand U10097 (N_10097,N_9445,N_9442);
nand U10098 (N_10098,N_9407,N_9527);
nand U10099 (N_10099,N_9040,N_9361);
nand U10100 (N_10100,N_9609,N_9211);
and U10101 (N_10101,N_9731,N_9165);
or U10102 (N_10102,N_9193,N_9478);
and U10103 (N_10103,N_9614,N_9130);
nor U10104 (N_10104,N_9135,N_9562);
and U10105 (N_10105,N_9320,N_9507);
nor U10106 (N_10106,N_9432,N_9629);
nor U10107 (N_10107,N_9224,N_9164);
and U10108 (N_10108,N_9618,N_9412);
nor U10109 (N_10109,N_9011,N_9326);
nand U10110 (N_10110,N_9215,N_9689);
nand U10111 (N_10111,N_9065,N_9607);
nor U10112 (N_10112,N_9414,N_9251);
nor U10113 (N_10113,N_9518,N_9735);
or U10114 (N_10114,N_9504,N_9603);
nand U10115 (N_10115,N_9198,N_9487);
and U10116 (N_10116,N_9479,N_9364);
nor U10117 (N_10117,N_9329,N_9288);
nand U10118 (N_10118,N_9587,N_9729);
and U10119 (N_10119,N_9391,N_9610);
nand U10120 (N_10120,N_9276,N_9221);
nand U10121 (N_10121,N_9077,N_9137);
nand U10122 (N_10122,N_9015,N_9192);
or U10123 (N_10123,N_9342,N_9028);
or U10124 (N_10124,N_9201,N_9321);
nor U10125 (N_10125,N_9442,N_9652);
nand U10126 (N_10126,N_9628,N_9244);
nand U10127 (N_10127,N_9294,N_9378);
nor U10128 (N_10128,N_9483,N_9192);
or U10129 (N_10129,N_9262,N_9526);
nor U10130 (N_10130,N_9273,N_9682);
nand U10131 (N_10131,N_9285,N_9490);
nand U10132 (N_10132,N_9147,N_9081);
xnor U10133 (N_10133,N_9498,N_9611);
or U10134 (N_10134,N_9516,N_9694);
nand U10135 (N_10135,N_9040,N_9550);
or U10136 (N_10136,N_9035,N_9241);
nand U10137 (N_10137,N_9291,N_9444);
or U10138 (N_10138,N_9446,N_9090);
nand U10139 (N_10139,N_9192,N_9273);
nor U10140 (N_10140,N_9700,N_9098);
nand U10141 (N_10141,N_9716,N_9722);
nand U10142 (N_10142,N_9223,N_9685);
nand U10143 (N_10143,N_9290,N_9476);
nor U10144 (N_10144,N_9121,N_9478);
and U10145 (N_10145,N_9740,N_9278);
or U10146 (N_10146,N_9059,N_9394);
or U10147 (N_10147,N_9654,N_9597);
nand U10148 (N_10148,N_9606,N_9161);
nand U10149 (N_10149,N_9164,N_9381);
and U10150 (N_10150,N_9732,N_9415);
and U10151 (N_10151,N_9197,N_9478);
nand U10152 (N_10152,N_9358,N_9242);
nand U10153 (N_10153,N_9741,N_9286);
or U10154 (N_10154,N_9232,N_9741);
or U10155 (N_10155,N_9046,N_9195);
and U10156 (N_10156,N_9015,N_9560);
nand U10157 (N_10157,N_9564,N_9256);
nand U10158 (N_10158,N_9128,N_9745);
or U10159 (N_10159,N_9083,N_9289);
or U10160 (N_10160,N_9333,N_9149);
and U10161 (N_10161,N_9236,N_9159);
nor U10162 (N_10162,N_9749,N_9468);
and U10163 (N_10163,N_9683,N_9240);
nor U10164 (N_10164,N_9274,N_9492);
or U10165 (N_10165,N_9543,N_9421);
and U10166 (N_10166,N_9233,N_9123);
and U10167 (N_10167,N_9195,N_9248);
nor U10168 (N_10168,N_9150,N_9177);
and U10169 (N_10169,N_9706,N_9197);
nand U10170 (N_10170,N_9304,N_9646);
nand U10171 (N_10171,N_9084,N_9718);
and U10172 (N_10172,N_9179,N_9722);
and U10173 (N_10173,N_9384,N_9213);
nor U10174 (N_10174,N_9210,N_9469);
nand U10175 (N_10175,N_9094,N_9300);
or U10176 (N_10176,N_9124,N_9354);
and U10177 (N_10177,N_9630,N_9568);
nor U10178 (N_10178,N_9243,N_9700);
nand U10179 (N_10179,N_9432,N_9607);
nand U10180 (N_10180,N_9315,N_9512);
nor U10181 (N_10181,N_9704,N_9163);
nand U10182 (N_10182,N_9490,N_9559);
nor U10183 (N_10183,N_9375,N_9259);
nand U10184 (N_10184,N_9264,N_9271);
nand U10185 (N_10185,N_9482,N_9136);
nand U10186 (N_10186,N_9649,N_9015);
nand U10187 (N_10187,N_9228,N_9011);
nand U10188 (N_10188,N_9058,N_9317);
nor U10189 (N_10189,N_9262,N_9712);
nand U10190 (N_10190,N_9015,N_9587);
and U10191 (N_10191,N_9246,N_9150);
nor U10192 (N_10192,N_9013,N_9224);
xnor U10193 (N_10193,N_9567,N_9673);
and U10194 (N_10194,N_9651,N_9401);
nand U10195 (N_10195,N_9484,N_9068);
and U10196 (N_10196,N_9570,N_9382);
nor U10197 (N_10197,N_9741,N_9466);
or U10198 (N_10198,N_9494,N_9152);
and U10199 (N_10199,N_9127,N_9709);
and U10200 (N_10200,N_9662,N_9459);
nand U10201 (N_10201,N_9097,N_9711);
nand U10202 (N_10202,N_9575,N_9535);
or U10203 (N_10203,N_9269,N_9112);
and U10204 (N_10204,N_9002,N_9406);
and U10205 (N_10205,N_9456,N_9469);
nand U10206 (N_10206,N_9372,N_9706);
and U10207 (N_10207,N_9484,N_9188);
nor U10208 (N_10208,N_9291,N_9717);
or U10209 (N_10209,N_9649,N_9078);
or U10210 (N_10210,N_9038,N_9402);
nor U10211 (N_10211,N_9032,N_9074);
nor U10212 (N_10212,N_9214,N_9224);
nor U10213 (N_10213,N_9077,N_9138);
or U10214 (N_10214,N_9108,N_9231);
and U10215 (N_10215,N_9438,N_9449);
and U10216 (N_10216,N_9402,N_9384);
and U10217 (N_10217,N_9734,N_9005);
nor U10218 (N_10218,N_9356,N_9400);
nand U10219 (N_10219,N_9104,N_9747);
nand U10220 (N_10220,N_9304,N_9699);
nor U10221 (N_10221,N_9460,N_9224);
nand U10222 (N_10222,N_9457,N_9662);
or U10223 (N_10223,N_9721,N_9319);
or U10224 (N_10224,N_9746,N_9546);
or U10225 (N_10225,N_9064,N_9648);
and U10226 (N_10226,N_9102,N_9603);
nand U10227 (N_10227,N_9443,N_9383);
and U10228 (N_10228,N_9692,N_9640);
or U10229 (N_10229,N_9069,N_9067);
nand U10230 (N_10230,N_9364,N_9170);
nor U10231 (N_10231,N_9289,N_9563);
nand U10232 (N_10232,N_9043,N_9719);
nor U10233 (N_10233,N_9265,N_9219);
xnor U10234 (N_10234,N_9505,N_9369);
or U10235 (N_10235,N_9000,N_9373);
nor U10236 (N_10236,N_9726,N_9453);
and U10237 (N_10237,N_9687,N_9417);
and U10238 (N_10238,N_9253,N_9337);
or U10239 (N_10239,N_9241,N_9140);
xor U10240 (N_10240,N_9272,N_9733);
or U10241 (N_10241,N_9717,N_9257);
and U10242 (N_10242,N_9285,N_9272);
and U10243 (N_10243,N_9220,N_9017);
and U10244 (N_10244,N_9713,N_9155);
nor U10245 (N_10245,N_9690,N_9006);
nor U10246 (N_10246,N_9582,N_9715);
nor U10247 (N_10247,N_9011,N_9053);
or U10248 (N_10248,N_9255,N_9717);
nand U10249 (N_10249,N_9014,N_9617);
or U10250 (N_10250,N_9657,N_9214);
and U10251 (N_10251,N_9618,N_9299);
xnor U10252 (N_10252,N_9025,N_9633);
or U10253 (N_10253,N_9721,N_9553);
and U10254 (N_10254,N_9692,N_9625);
nand U10255 (N_10255,N_9076,N_9262);
nand U10256 (N_10256,N_9569,N_9463);
or U10257 (N_10257,N_9444,N_9040);
nor U10258 (N_10258,N_9207,N_9566);
and U10259 (N_10259,N_9733,N_9444);
nor U10260 (N_10260,N_9482,N_9543);
nand U10261 (N_10261,N_9571,N_9630);
nor U10262 (N_10262,N_9086,N_9704);
or U10263 (N_10263,N_9129,N_9304);
nor U10264 (N_10264,N_9351,N_9337);
nor U10265 (N_10265,N_9008,N_9004);
nor U10266 (N_10266,N_9622,N_9594);
and U10267 (N_10267,N_9746,N_9605);
or U10268 (N_10268,N_9215,N_9077);
nand U10269 (N_10269,N_9328,N_9130);
nor U10270 (N_10270,N_9579,N_9125);
nand U10271 (N_10271,N_9423,N_9703);
or U10272 (N_10272,N_9744,N_9556);
nor U10273 (N_10273,N_9504,N_9289);
and U10274 (N_10274,N_9685,N_9252);
or U10275 (N_10275,N_9567,N_9650);
nand U10276 (N_10276,N_9540,N_9535);
and U10277 (N_10277,N_9546,N_9152);
nor U10278 (N_10278,N_9092,N_9726);
xnor U10279 (N_10279,N_9342,N_9142);
nand U10280 (N_10280,N_9035,N_9135);
and U10281 (N_10281,N_9082,N_9333);
or U10282 (N_10282,N_9003,N_9688);
nand U10283 (N_10283,N_9404,N_9702);
nand U10284 (N_10284,N_9492,N_9324);
nor U10285 (N_10285,N_9739,N_9297);
nand U10286 (N_10286,N_9643,N_9411);
and U10287 (N_10287,N_9404,N_9140);
and U10288 (N_10288,N_9707,N_9526);
and U10289 (N_10289,N_9084,N_9644);
or U10290 (N_10290,N_9518,N_9131);
nand U10291 (N_10291,N_9704,N_9306);
or U10292 (N_10292,N_9736,N_9719);
and U10293 (N_10293,N_9348,N_9706);
and U10294 (N_10294,N_9337,N_9504);
nand U10295 (N_10295,N_9164,N_9538);
or U10296 (N_10296,N_9019,N_9623);
nand U10297 (N_10297,N_9135,N_9519);
xnor U10298 (N_10298,N_9616,N_9245);
nand U10299 (N_10299,N_9261,N_9033);
and U10300 (N_10300,N_9395,N_9405);
and U10301 (N_10301,N_9308,N_9460);
and U10302 (N_10302,N_9386,N_9003);
nor U10303 (N_10303,N_9730,N_9652);
nor U10304 (N_10304,N_9434,N_9388);
or U10305 (N_10305,N_9742,N_9375);
nand U10306 (N_10306,N_9324,N_9098);
nand U10307 (N_10307,N_9352,N_9683);
or U10308 (N_10308,N_9429,N_9670);
nand U10309 (N_10309,N_9071,N_9527);
nor U10310 (N_10310,N_9444,N_9081);
xor U10311 (N_10311,N_9425,N_9746);
nor U10312 (N_10312,N_9368,N_9302);
or U10313 (N_10313,N_9045,N_9503);
or U10314 (N_10314,N_9113,N_9137);
nor U10315 (N_10315,N_9064,N_9673);
nand U10316 (N_10316,N_9373,N_9296);
nand U10317 (N_10317,N_9123,N_9261);
and U10318 (N_10318,N_9034,N_9746);
nor U10319 (N_10319,N_9363,N_9533);
or U10320 (N_10320,N_9472,N_9578);
nand U10321 (N_10321,N_9451,N_9526);
or U10322 (N_10322,N_9108,N_9651);
nand U10323 (N_10323,N_9583,N_9681);
nor U10324 (N_10324,N_9123,N_9167);
nand U10325 (N_10325,N_9291,N_9349);
nor U10326 (N_10326,N_9221,N_9498);
or U10327 (N_10327,N_9171,N_9690);
nor U10328 (N_10328,N_9062,N_9596);
xnor U10329 (N_10329,N_9551,N_9464);
nor U10330 (N_10330,N_9433,N_9737);
or U10331 (N_10331,N_9638,N_9382);
or U10332 (N_10332,N_9503,N_9301);
or U10333 (N_10333,N_9012,N_9289);
nor U10334 (N_10334,N_9429,N_9671);
nor U10335 (N_10335,N_9245,N_9612);
nor U10336 (N_10336,N_9695,N_9441);
nor U10337 (N_10337,N_9515,N_9489);
and U10338 (N_10338,N_9732,N_9041);
nor U10339 (N_10339,N_9513,N_9303);
nand U10340 (N_10340,N_9274,N_9159);
or U10341 (N_10341,N_9627,N_9667);
nand U10342 (N_10342,N_9315,N_9066);
nor U10343 (N_10343,N_9276,N_9130);
nor U10344 (N_10344,N_9557,N_9716);
or U10345 (N_10345,N_9728,N_9250);
nand U10346 (N_10346,N_9132,N_9459);
and U10347 (N_10347,N_9384,N_9102);
nor U10348 (N_10348,N_9078,N_9472);
nor U10349 (N_10349,N_9392,N_9487);
nor U10350 (N_10350,N_9147,N_9369);
nor U10351 (N_10351,N_9046,N_9377);
nand U10352 (N_10352,N_9041,N_9316);
nor U10353 (N_10353,N_9161,N_9619);
or U10354 (N_10354,N_9653,N_9584);
or U10355 (N_10355,N_9205,N_9261);
or U10356 (N_10356,N_9142,N_9061);
or U10357 (N_10357,N_9709,N_9488);
nor U10358 (N_10358,N_9571,N_9439);
or U10359 (N_10359,N_9583,N_9581);
or U10360 (N_10360,N_9112,N_9499);
nor U10361 (N_10361,N_9124,N_9710);
nand U10362 (N_10362,N_9315,N_9744);
nand U10363 (N_10363,N_9360,N_9668);
nor U10364 (N_10364,N_9535,N_9516);
nand U10365 (N_10365,N_9328,N_9168);
and U10366 (N_10366,N_9209,N_9268);
nor U10367 (N_10367,N_9027,N_9178);
nor U10368 (N_10368,N_9088,N_9094);
nor U10369 (N_10369,N_9388,N_9221);
nor U10370 (N_10370,N_9437,N_9081);
nor U10371 (N_10371,N_9130,N_9653);
or U10372 (N_10372,N_9565,N_9742);
or U10373 (N_10373,N_9720,N_9026);
nand U10374 (N_10374,N_9001,N_9689);
nor U10375 (N_10375,N_9569,N_9540);
and U10376 (N_10376,N_9282,N_9287);
and U10377 (N_10377,N_9084,N_9391);
nand U10378 (N_10378,N_9031,N_9103);
or U10379 (N_10379,N_9626,N_9698);
nor U10380 (N_10380,N_9642,N_9348);
or U10381 (N_10381,N_9671,N_9407);
or U10382 (N_10382,N_9668,N_9235);
and U10383 (N_10383,N_9298,N_9242);
nand U10384 (N_10384,N_9694,N_9508);
and U10385 (N_10385,N_9435,N_9269);
or U10386 (N_10386,N_9368,N_9420);
and U10387 (N_10387,N_9286,N_9678);
nand U10388 (N_10388,N_9383,N_9630);
nand U10389 (N_10389,N_9314,N_9587);
nand U10390 (N_10390,N_9088,N_9102);
and U10391 (N_10391,N_9628,N_9064);
or U10392 (N_10392,N_9139,N_9180);
nand U10393 (N_10393,N_9560,N_9366);
nand U10394 (N_10394,N_9138,N_9349);
nand U10395 (N_10395,N_9302,N_9406);
or U10396 (N_10396,N_9399,N_9042);
and U10397 (N_10397,N_9348,N_9478);
or U10398 (N_10398,N_9470,N_9280);
nor U10399 (N_10399,N_9102,N_9130);
or U10400 (N_10400,N_9250,N_9546);
nand U10401 (N_10401,N_9056,N_9713);
and U10402 (N_10402,N_9607,N_9057);
and U10403 (N_10403,N_9371,N_9589);
nor U10404 (N_10404,N_9657,N_9251);
or U10405 (N_10405,N_9277,N_9059);
and U10406 (N_10406,N_9310,N_9073);
or U10407 (N_10407,N_9504,N_9086);
nor U10408 (N_10408,N_9319,N_9275);
nand U10409 (N_10409,N_9635,N_9629);
nand U10410 (N_10410,N_9067,N_9454);
nand U10411 (N_10411,N_9684,N_9600);
nand U10412 (N_10412,N_9141,N_9595);
nor U10413 (N_10413,N_9526,N_9154);
nor U10414 (N_10414,N_9511,N_9010);
or U10415 (N_10415,N_9038,N_9608);
and U10416 (N_10416,N_9691,N_9463);
nor U10417 (N_10417,N_9000,N_9366);
or U10418 (N_10418,N_9084,N_9437);
nor U10419 (N_10419,N_9055,N_9102);
nor U10420 (N_10420,N_9029,N_9219);
nor U10421 (N_10421,N_9430,N_9529);
xor U10422 (N_10422,N_9503,N_9437);
or U10423 (N_10423,N_9664,N_9080);
and U10424 (N_10424,N_9156,N_9446);
and U10425 (N_10425,N_9740,N_9078);
nand U10426 (N_10426,N_9039,N_9695);
nand U10427 (N_10427,N_9606,N_9209);
and U10428 (N_10428,N_9434,N_9547);
and U10429 (N_10429,N_9671,N_9427);
nor U10430 (N_10430,N_9008,N_9641);
or U10431 (N_10431,N_9039,N_9145);
or U10432 (N_10432,N_9712,N_9248);
and U10433 (N_10433,N_9691,N_9198);
nand U10434 (N_10434,N_9041,N_9119);
nand U10435 (N_10435,N_9165,N_9730);
or U10436 (N_10436,N_9656,N_9563);
nor U10437 (N_10437,N_9225,N_9081);
nand U10438 (N_10438,N_9733,N_9417);
nand U10439 (N_10439,N_9565,N_9283);
or U10440 (N_10440,N_9514,N_9303);
nor U10441 (N_10441,N_9019,N_9397);
and U10442 (N_10442,N_9550,N_9667);
and U10443 (N_10443,N_9108,N_9647);
nand U10444 (N_10444,N_9206,N_9282);
nor U10445 (N_10445,N_9521,N_9354);
nor U10446 (N_10446,N_9575,N_9065);
nor U10447 (N_10447,N_9212,N_9332);
nor U10448 (N_10448,N_9194,N_9192);
and U10449 (N_10449,N_9539,N_9587);
nor U10450 (N_10450,N_9492,N_9157);
nor U10451 (N_10451,N_9006,N_9046);
or U10452 (N_10452,N_9326,N_9631);
nand U10453 (N_10453,N_9382,N_9733);
and U10454 (N_10454,N_9507,N_9497);
and U10455 (N_10455,N_9057,N_9179);
and U10456 (N_10456,N_9210,N_9652);
and U10457 (N_10457,N_9067,N_9572);
and U10458 (N_10458,N_9620,N_9340);
and U10459 (N_10459,N_9011,N_9482);
or U10460 (N_10460,N_9534,N_9092);
and U10461 (N_10461,N_9260,N_9251);
and U10462 (N_10462,N_9141,N_9146);
nand U10463 (N_10463,N_9726,N_9370);
or U10464 (N_10464,N_9564,N_9057);
and U10465 (N_10465,N_9721,N_9406);
nand U10466 (N_10466,N_9391,N_9069);
and U10467 (N_10467,N_9582,N_9074);
and U10468 (N_10468,N_9221,N_9081);
nor U10469 (N_10469,N_9648,N_9460);
or U10470 (N_10470,N_9263,N_9518);
and U10471 (N_10471,N_9271,N_9049);
nand U10472 (N_10472,N_9285,N_9701);
and U10473 (N_10473,N_9294,N_9145);
or U10474 (N_10474,N_9605,N_9551);
nand U10475 (N_10475,N_9196,N_9354);
and U10476 (N_10476,N_9547,N_9032);
or U10477 (N_10477,N_9179,N_9195);
and U10478 (N_10478,N_9193,N_9458);
and U10479 (N_10479,N_9358,N_9298);
or U10480 (N_10480,N_9044,N_9569);
and U10481 (N_10481,N_9003,N_9344);
nor U10482 (N_10482,N_9501,N_9019);
or U10483 (N_10483,N_9134,N_9007);
or U10484 (N_10484,N_9148,N_9633);
nand U10485 (N_10485,N_9365,N_9510);
or U10486 (N_10486,N_9253,N_9702);
nor U10487 (N_10487,N_9149,N_9581);
nor U10488 (N_10488,N_9211,N_9700);
nor U10489 (N_10489,N_9092,N_9469);
nor U10490 (N_10490,N_9607,N_9388);
nand U10491 (N_10491,N_9043,N_9097);
nand U10492 (N_10492,N_9337,N_9415);
nor U10493 (N_10493,N_9023,N_9381);
or U10494 (N_10494,N_9314,N_9503);
nor U10495 (N_10495,N_9603,N_9473);
or U10496 (N_10496,N_9073,N_9223);
nand U10497 (N_10497,N_9092,N_9462);
and U10498 (N_10498,N_9730,N_9384);
nand U10499 (N_10499,N_9518,N_9233);
nand U10500 (N_10500,N_10067,N_9947);
and U10501 (N_10501,N_9953,N_9849);
nand U10502 (N_10502,N_10153,N_10293);
nor U10503 (N_10503,N_9843,N_10047);
nand U10504 (N_10504,N_10408,N_10444);
and U10505 (N_10505,N_9973,N_10468);
nand U10506 (N_10506,N_10278,N_10482);
nand U10507 (N_10507,N_10222,N_9908);
nand U10508 (N_10508,N_10152,N_10435);
nand U10509 (N_10509,N_10422,N_10169);
and U10510 (N_10510,N_10127,N_10023);
nand U10511 (N_10511,N_10082,N_9889);
and U10512 (N_10512,N_10395,N_9836);
or U10513 (N_10513,N_10325,N_10328);
nand U10514 (N_10514,N_10072,N_10119);
nor U10515 (N_10515,N_10176,N_10296);
and U10516 (N_10516,N_10024,N_10002);
and U10517 (N_10517,N_10004,N_10077);
and U10518 (N_10518,N_10020,N_9971);
nand U10519 (N_10519,N_10146,N_10184);
or U10520 (N_10520,N_10148,N_10285);
nand U10521 (N_10521,N_10231,N_10490);
nand U10522 (N_10522,N_10027,N_10359);
nor U10523 (N_10523,N_10149,N_10173);
nand U10524 (N_10524,N_10415,N_10229);
nor U10525 (N_10525,N_10466,N_10262);
nand U10526 (N_10526,N_10459,N_10301);
nand U10527 (N_10527,N_10043,N_10015);
nor U10528 (N_10528,N_9978,N_10066);
or U10529 (N_10529,N_10268,N_9764);
nor U10530 (N_10530,N_10460,N_10236);
nand U10531 (N_10531,N_10085,N_9929);
or U10532 (N_10532,N_10202,N_9757);
xnor U10533 (N_10533,N_9844,N_10138);
nor U10534 (N_10534,N_9852,N_10336);
nor U10535 (N_10535,N_10496,N_10075);
and U10536 (N_10536,N_10356,N_9962);
and U10537 (N_10537,N_10239,N_9858);
nor U10538 (N_10538,N_9808,N_9893);
nand U10539 (N_10539,N_9802,N_9963);
or U10540 (N_10540,N_10070,N_9950);
nand U10541 (N_10541,N_10255,N_9898);
nand U10542 (N_10542,N_10011,N_10494);
nand U10543 (N_10543,N_10279,N_9816);
and U10544 (N_10544,N_9930,N_10489);
and U10545 (N_10545,N_9803,N_9912);
nand U10546 (N_10546,N_10495,N_10358);
xor U10547 (N_10547,N_10209,N_10025);
and U10548 (N_10548,N_9928,N_10432);
nor U10549 (N_10549,N_10197,N_10175);
or U10550 (N_10550,N_9940,N_10165);
nand U10551 (N_10551,N_9957,N_10150);
nor U10552 (N_10552,N_9961,N_9883);
and U10553 (N_10553,N_10414,N_9887);
nor U10554 (N_10554,N_10218,N_9993);
xnor U10555 (N_10555,N_10054,N_10396);
and U10556 (N_10556,N_9906,N_9872);
or U10557 (N_10557,N_9968,N_10102);
nor U10558 (N_10558,N_10322,N_10041);
and U10559 (N_10559,N_10330,N_10294);
xnor U10560 (N_10560,N_10284,N_10032);
and U10561 (N_10561,N_9865,N_9966);
and U10562 (N_10562,N_10309,N_9825);
nor U10563 (N_10563,N_9787,N_9987);
and U10564 (N_10564,N_10497,N_9926);
nand U10565 (N_10565,N_10340,N_9919);
nand U10566 (N_10566,N_9853,N_10472);
or U10567 (N_10567,N_10005,N_10090);
and U10568 (N_10568,N_10483,N_10334);
or U10569 (N_10569,N_9954,N_10323);
nand U10570 (N_10570,N_10196,N_10003);
or U10571 (N_10571,N_10326,N_10155);
and U10572 (N_10572,N_10170,N_10052);
xor U10573 (N_10573,N_9800,N_9925);
and U10574 (N_10574,N_9864,N_9877);
nor U10575 (N_10575,N_10192,N_10178);
and U10576 (N_10576,N_10462,N_9988);
and U10577 (N_10577,N_9900,N_9779);
nand U10578 (N_10578,N_10068,N_10303);
or U10579 (N_10579,N_9996,N_9861);
nor U10580 (N_10580,N_9923,N_9845);
nor U10581 (N_10581,N_9886,N_9760);
and U10582 (N_10582,N_9841,N_10225);
nand U10583 (N_10583,N_9897,N_10058);
and U10584 (N_10584,N_10089,N_10012);
nor U10585 (N_10585,N_10136,N_10131);
nand U10586 (N_10586,N_9927,N_10088);
and U10587 (N_10587,N_10282,N_10476);
nor U10588 (N_10588,N_9932,N_9851);
and U10589 (N_10589,N_10252,N_9944);
nor U10590 (N_10590,N_10306,N_10167);
and U10591 (N_10591,N_10064,N_10083);
nand U10592 (N_10592,N_10106,N_10122);
or U10593 (N_10593,N_10286,N_9870);
and U10594 (N_10594,N_10246,N_10061);
nor U10595 (N_10595,N_10276,N_9773);
and U10596 (N_10596,N_10139,N_9949);
nor U10597 (N_10597,N_9796,N_9982);
nor U10598 (N_10598,N_10186,N_10449);
and U10599 (N_10599,N_9890,N_10310);
nor U10600 (N_10600,N_10256,N_9960);
nand U10601 (N_10601,N_10393,N_9847);
nor U10602 (N_10602,N_10158,N_10187);
and U10603 (N_10603,N_10223,N_10345);
or U10604 (N_10604,N_10308,N_10248);
nor U10605 (N_10605,N_10200,N_10346);
nand U10606 (N_10606,N_10379,N_9995);
nor U10607 (N_10607,N_10313,N_9892);
and U10608 (N_10608,N_9876,N_9821);
or U10609 (N_10609,N_10441,N_10368);
or U10610 (N_10610,N_10295,N_10029);
or U10611 (N_10611,N_9917,N_10475);
nand U10612 (N_10612,N_10046,N_10215);
and U10613 (N_10613,N_9933,N_10166);
and U10614 (N_10614,N_9899,N_9922);
nor U10615 (N_10615,N_10055,N_10266);
or U10616 (N_10616,N_10172,N_10087);
nand U10617 (N_10617,N_9904,N_10477);
or U10618 (N_10618,N_9873,N_10144);
nor U10619 (N_10619,N_9989,N_10201);
and U10620 (N_10620,N_10493,N_10264);
or U10621 (N_10621,N_10314,N_10260);
nand U10622 (N_10622,N_10230,N_10190);
nor U10623 (N_10623,N_9780,N_10458);
or U10624 (N_10624,N_10171,N_9905);
nor U10625 (N_10625,N_10243,N_9918);
nand U10626 (N_10626,N_10084,N_10352);
nand U10627 (N_10627,N_9850,N_10374);
xnor U10628 (N_10628,N_10026,N_10143);
and U10629 (N_10629,N_9983,N_10307);
or U10630 (N_10630,N_9826,N_10220);
nor U10631 (N_10631,N_10219,N_10018);
nor U10632 (N_10632,N_9942,N_10344);
nor U10633 (N_10633,N_9814,N_10125);
nor U10634 (N_10634,N_9750,N_10233);
nor U10635 (N_10635,N_9763,N_9767);
or U10636 (N_10636,N_9920,N_10241);
and U10637 (N_10637,N_10244,N_10337);
or U10638 (N_10638,N_9797,N_9976);
nand U10639 (N_10639,N_10382,N_10259);
nand U10640 (N_10640,N_10179,N_9785);
nor U10641 (N_10641,N_10198,N_10288);
nand U10642 (N_10642,N_10351,N_9924);
nor U10643 (N_10643,N_10271,N_10329);
or U10644 (N_10644,N_10390,N_10370);
nand U10645 (N_10645,N_9761,N_10429);
and U10646 (N_10646,N_9972,N_10433);
and U10647 (N_10647,N_9879,N_10478);
and U10648 (N_10648,N_9986,N_9846);
nand U10649 (N_10649,N_10133,N_10380);
nor U10650 (N_10650,N_9751,N_10141);
nand U10651 (N_10651,N_9772,N_9762);
nor U10652 (N_10652,N_10180,N_9938);
and U10653 (N_10653,N_9948,N_9842);
or U10654 (N_10654,N_9874,N_10383);
nand U10655 (N_10655,N_10445,N_10321);
nor U10656 (N_10656,N_10080,N_9866);
nand U10657 (N_10657,N_9801,N_10471);
nand U10658 (N_10658,N_9791,N_10404);
nor U10659 (N_10659,N_10430,N_10487);
or U10660 (N_10660,N_10385,N_10203);
or U10661 (N_10661,N_9964,N_9774);
and U10662 (N_10662,N_10355,N_9820);
nor U10663 (N_10663,N_9969,N_10413);
nand U10664 (N_10664,N_10327,N_9768);
or U10665 (N_10665,N_10137,N_10436);
or U10666 (N_10666,N_9979,N_9792);
nand U10667 (N_10667,N_10121,N_10056);
nand U10668 (N_10668,N_10287,N_9867);
and U10669 (N_10669,N_10300,N_10074);
nor U10670 (N_10670,N_10378,N_9981);
or U10671 (N_10671,N_10134,N_10335);
and U10672 (N_10672,N_10315,N_10044);
and U10673 (N_10673,N_10124,N_10107);
nand U10674 (N_10674,N_9939,N_10120);
or U10675 (N_10675,N_10464,N_10417);
nor U10676 (N_10676,N_10037,N_10114);
xnor U10677 (N_10677,N_9848,N_10022);
nor U10678 (N_10678,N_10371,N_10272);
nor U10679 (N_10679,N_10484,N_10384);
or U10680 (N_10680,N_10049,N_10113);
nand U10681 (N_10681,N_10177,N_10492);
nor U10682 (N_10682,N_10110,N_9885);
nor U10683 (N_10683,N_10332,N_9752);
nand U10684 (N_10684,N_10410,N_10226);
nand U10685 (N_10685,N_10305,N_10250);
nand U10686 (N_10686,N_9936,N_10428);
nand U10687 (N_10687,N_10238,N_9856);
nand U10688 (N_10688,N_9888,N_10258);
or U10689 (N_10689,N_10103,N_9952);
or U10690 (N_10690,N_10001,N_10208);
or U10691 (N_10691,N_10304,N_9935);
and U10692 (N_10692,N_10425,N_9882);
nand U10693 (N_10693,N_9789,N_10245);
and U10694 (N_10694,N_9910,N_10028);
nor U10695 (N_10695,N_9788,N_10443);
nor U10696 (N_10696,N_9804,N_10420);
or U10697 (N_10697,N_10275,N_10031);
and U10698 (N_10698,N_10214,N_10096);
or U10699 (N_10699,N_10079,N_10183);
and U10700 (N_10700,N_10405,N_10160);
nand U10701 (N_10701,N_9869,N_10455);
nor U10702 (N_10702,N_9794,N_9891);
nand U10703 (N_10703,N_9937,N_10470);
xnor U10704 (N_10704,N_9753,N_9831);
nor U10705 (N_10705,N_9975,N_9799);
nor U10706 (N_10706,N_10481,N_10185);
or U10707 (N_10707,N_10213,N_10343);
nor U10708 (N_10708,N_10423,N_10499);
nor U10709 (N_10709,N_10257,N_9758);
nand U10710 (N_10710,N_10035,N_10129);
or U10711 (N_10711,N_10440,N_10453);
or U10712 (N_10712,N_10191,N_10253);
and U10713 (N_10713,N_10227,N_10485);
or U10714 (N_10714,N_10232,N_9991);
nand U10715 (N_10715,N_9777,N_10357);
nand U10716 (N_10716,N_10045,N_10463);
nor U10717 (N_10717,N_10115,N_10099);
nand U10718 (N_10718,N_9756,N_9863);
or U10719 (N_10719,N_10274,N_10094);
and U10720 (N_10720,N_10265,N_9999);
nor U10721 (N_10721,N_10142,N_10394);
or U10722 (N_10722,N_10311,N_10164);
nor U10723 (N_10723,N_9830,N_9965);
nand U10724 (N_10724,N_9824,N_10474);
and U10725 (N_10725,N_9818,N_10235);
or U10726 (N_10726,N_10254,N_10036);
nor U10727 (N_10727,N_9881,N_10350);
nor U10728 (N_10728,N_10159,N_10416);
nand U10729 (N_10729,N_10181,N_10210);
or U10730 (N_10730,N_10498,N_9829);
nor U10731 (N_10731,N_10442,N_9806);
and U10732 (N_10732,N_10317,N_10132);
and U10733 (N_10733,N_10418,N_10448);
nand U10734 (N_10734,N_9984,N_9857);
and U10735 (N_10735,N_10281,N_10062);
and U10736 (N_10736,N_9992,N_9833);
and U10737 (N_10737,N_9838,N_10362);
nand U10738 (N_10738,N_9781,N_9980);
nor U10739 (N_10739,N_9967,N_9997);
nor U10740 (N_10740,N_10277,N_9809);
nor U10741 (N_10741,N_10363,N_9812);
or U10742 (N_10742,N_10400,N_10205);
nand U10743 (N_10743,N_10348,N_10000);
and U10744 (N_10744,N_9878,N_10071);
nand U10745 (N_10745,N_10316,N_10069);
and U10746 (N_10746,N_10389,N_10040);
and U10747 (N_10747,N_10108,N_10078);
nand U10748 (N_10748,N_9786,N_9955);
nand U10749 (N_10749,N_10488,N_9793);
nand U10750 (N_10750,N_10193,N_10302);
and U10751 (N_10751,N_10421,N_9921);
or U10752 (N_10752,N_10365,N_10211);
and U10753 (N_10753,N_10109,N_10147);
nand U10754 (N_10754,N_10369,N_10216);
nor U10755 (N_10755,N_10439,N_10341);
nor U10756 (N_10756,N_10373,N_9934);
and U10757 (N_10757,N_9817,N_10398);
or U10758 (N_10758,N_10360,N_10375);
and U10759 (N_10759,N_9859,N_9784);
or U10760 (N_10760,N_10057,N_10409);
nor U10761 (N_10761,N_9909,N_10342);
and U10762 (N_10762,N_10269,N_9884);
or U10763 (N_10763,N_9970,N_10263);
or U10764 (N_10764,N_10364,N_10039);
and U10765 (N_10765,N_10467,N_10034);
nand U10766 (N_10766,N_10399,N_9766);
or U10767 (N_10767,N_9837,N_9823);
nor U10768 (N_10768,N_10480,N_10053);
and U10769 (N_10769,N_9770,N_10116);
or U10770 (N_10770,N_10093,N_10479);
nand U10771 (N_10771,N_10101,N_10412);
nor U10772 (N_10772,N_10299,N_9895);
nor U10773 (N_10773,N_10033,N_10098);
and U10774 (N_10774,N_10388,N_10411);
or U10775 (N_10775,N_9868,N_10240);
and U10776 (N_10776,N_9828,N_10491);
nor U10777 (N_10777,N_9896,N_9945);
and U10778 (N_10778,N_10457,N_10081);
or U10779 (N_10779,N_10189,N_10157);
and U10780 (N_10780,N_10473,N_10419);
nand U10781 (N_10781,N_10426,N_10204);
nor U10782 (N_10782,N_10059,N_9977);
and U10783 (N_10783,N_10130,N_10063);
and U10784 (N_10784,N_9822,N_10437);
and U10785 (N_10785,N_9985,N_10267);
nand U10786 (N_10786,N_9805,N_10249);
or U10787 (N_10787,N_9875,N_10104);
and U10788 (N_10788,N_9835,N_10283);
or U10789 (N_10789,N_10391,N_10401);
or U10790 (N_10790,N_9769,N_9807);
or U10791 (N_10791,N_9998,N_9931);
and U10792 (N_10792,N_10312,N_10469);
nand U10793 (N_10793,N_10261,N_10387);
nand U10794 (N_10794,N_10100,N_9855);
nor U10795 (N_10795,N_9903,N_10318);
nor U10796 (N_10796,N_9941,N_10403);
or U10797 (N_10797,N_10347,N_10438);
nor U10798 (N_10798,N_9783,N_10361);
nor U10799 (N_10799,N_10280,N_10456);
and U10800 (N_10800,N_9946,N_9871);
nand U10801 (N_10801,N_10486,N_10195);
nand U10802 (N_10802,N_9994,N_10427);
or U10803 (N_10803,N_10434,N_10123);
or U10804 (N_10804,N_10320,N_9754);
nand U10805 (N_10805,N_10095,N_10135);
or U10806 (N_10806,N_9880,N_9790);
or U10807 (N_10807,N_10016,N_10174);
or U10808 (N_10808,N_10048,N_10406);
nand U10809 (N_10809,N_10247,N_10006);
nor U10810 (N_10810,N_9862,N_10212);
or U10811 (N_10811,N_9759,N_10010);
nand U10812 (N_10812,N_10188,N_10156);
and U10813 (N_10813,N_9815,N_9755);
nor U10814 (N_10814,N_10465,N_10402);
or U10815 (N_10815,N_9798,N_10050);
and U10816 (N_10816,N_9907,N_10377);
and U10817 (N_10817,N_10161,N_9913);
nand U10818 (N_10818,N_9990,N_10182);
and U10819 (N_10819,N_9914,N_10091);
nor U10820 (N_10820,N_10117,N_9765);
nand U10821 (N_10821,N_10228,N_10030);
nor U10822 (N_10822,N_10446,N_10289);
and U10823 (N_10823,N_10424,N_9775);
nand U10824 (N_10824,N_10447,N_10038);
or U10825 (N_10825,N_10454,N_9771);
and U10826 (N_10826,N_10354,N_10128);
and U10827 (N_10827,N_10298,N_10111);
nand U10828 (N_10828,N_10060,N_10092);
nor U10829 (N_10829,N_10042,N_9839);
nand U10830 (N_10830,N_10331,N_10163);
nor U10831 (N_10831,N_9911,N_10145);
nor U10832 (N_10832,N_10234,N_9795);
nand U10833 (N_10833,N_10199,N_9854);
nor U10834 (N_10834,N_9782,N_10386);
nor U10835 (N_10835,N_10431,N_10251);
nor U10836 (N_10836,N_10297,N_10008);
nand U10837 (N_10837,N_10112,N_10339);
nand U10838 (N_10838,N_10461,N_10353);
and U10839 (N_10839,N_10017,N_9840);
nor U10840 (N_10840,N_9956,N_10207);
nor U10841 (N_10841,N_10162,N_10086);
nand U10842 (N_10842,N_10206,N_9894);
nor U10843 (N_10843,N_9832,N_10349);
and U10844 (N_10844,N_9915,N_9974);
nand U10845 (N_10845,N_10319,N_9959);
nand U10846 (N_10846,N_10290,N_10367);
or U10847 (N_10847,N_10452,N_10065);
nand U10848 (N_10848,N_10073,N_10126);
and U10849 (N_10849,N_10151,N_9813);
nand U10850 (N_10850,N_10097,N_9810);
or U10851 (N_10851,N_10407,N_9778);
nor U10852 (N_10852,N_10366,N_10013);
nand U10853 (N_10853,N_10194,N_10051);
or U10854 (N_10854,N_10237,N_10076);
or U10855 (N_10855,N_10270,N_9860);
nor U10856 (N_10856,N_10014,N_10372);
nor U10857 (N_10857,N_10009,N_9827);
nand U10858 (N_10858,N_10242,N_10451);
or U10859 (N_10859,N_9958,N_10291);
nand U10860 (N_10860,N_10392,N_10333);
or U10861 (N_10861,N_9811,N_10397);
nand U10862 (N_10862,N_10450,N_10292);
and U10863 (N_10863,N_9776,N_9901);
or U10864 (N_10864,N_9834,N_10273);
nand U10865 (N_10865,N_10021,N_10221);
and U10866 (N_10866,N_10140,N_10019);
nand U10867 (N_10867,N_9943,N_10105);
and U10868 (N_10868,N_9902,N_10324);
and U10869 (N_10869,N_10217,N_10154);
and U10870 (N_10870,N_9819,N_10007);
and U10871 (N_10871,N_10118,N_10224);
or U10872 (N_10872,N_10168,N_10376);
and U10873 (N_10873,N_10338,N_10381);
nor U10874 (N_10874,N_9916,N_9951);
or U10875 (N_10875,N_9832,N_9886);
xor U10876 (N_10876,N_10050,N_9920);
nor U10877 (N_10877,N_10404,N_10065);
nor U10878 (N_10878,N_9885,N_9933);
nor U10879 (N_10879,N_10342,N_10020);
or U10880 (N_10880,N_10290,N_10380);
and U10881 (N_10881,N_10134,N_10475);
and U10882 (N_10882,N_10381,N_9885);
nor U10883 (N_10883,N_10352,N_10117);
and U10884 (N_10884,N_10115,N_9841);
or U10885 (N_10885,N_9857,N_10030);
and U10886 (N_10886,N_9867,N_10483);
nor U10887 (N_10887,N_9804,N_10338);
nor U10888 (N_10888,N_10161,N_10368);
nand U10889 (N_10889,N_9926,N_10031);
nor U10890 (N_10890,N_10410,N_10268);
nand U10891 (N_10891,N_10245,N_9946);
or U10892 (N_10892,N_10220,N_10482);
nand U10893 (N_10893,N_10018,N_10240);
nand U10894 (N_10894,N_10420,N_10365);
nand U10895 (N_10895,N_10380,N_10145);
nand U10896 (N_10896,N_10465,N_9987);
and U10897 (N_10897,N_10467,N_10346);
and U10898 (N_10898,N_10004,N_10192);
or U10899 (N_10899,N_10245,N_10007);
and U10900 (N_10900,N_10225,N_9793);
or U10901 (N_10901,N_10060,N_9805);
nor U10902 (N_10902,N_9916,N_9959);
or U10903 (N_10903,N_10436,N_9756);
xor U10904 (N_10904,N_10106,N_10345);
or U10905 (N_10905,N_10455,N_10164);
or U10906 (N_10906,N_10371,N_10125);
nand U10907 (N_10907,N_10019,N_10408);
and U10908 (N_10908,N_9928,N_9851);
nor U10909 (N_10909,N_10285,N_10327);
nor U10910 (N_10910,N_10217,N_10233);
nand U10911 (N_10911,N_10298,N_10029);
nand U10912 (N_10912,N_10374,N_10289);
or U10913 (N_10913,N_10413,N_9755);
or U10914 (N_10914,N_9960,N_9837);
nand U10915 (N_10915,N_10488,N_10399);
nor U10916 (N_10916,N_9944,N_10293);
nor U10917 (N_10917,N_10193,N_10327);
and U10918 (N_10918,N_10064,N_9939);
and U10919 (N_10919,N_10124,N_9982);
nand U10920 (N_10920,N_10368,N_10082);
nand U10921 (N_10921,N_10335,N_9887);
nor U10922 (N_10922,N_10177,N_10040);
or U10923 (N_10923,N_9752,N_10357);
and U10924 (N_10924,N_10461,N_9987);
nand U10925 (N_10925,N_10045,N_9884);
or U10926 (N_10926,N_9860,N_9922);
nor U10927 (N_10927,N_10192,N_10207);
nand U10928 (N_10928,N_10016,N_10179);
and U10929 (N_10929,N_10150,N_10327);
nand U10930 (N_10930,N_10022,N_10118);
nor U10931 (N_10931,N_9897,N_10453);
nand U10932 (N_10932,N_10474,N_10254);
xnor U10933 (N_10933,N_9906,N_10051);
nor U10934 (N_10934,N_10351,N_10341);
nor U10935 (N_10935,N_10087,N_9873);
nand U10936 (N_10936,N_10186,N_9830);
or U10937 (N_10937,N_10187,N_10249);
nor U10938 (N_10938,N_9912,N_10372);
and U10939 (N_10939,N_9858,N_10068);
nor U10940 (N_10940,N_9950,N_9838);
and U10941 (N_10941,N_10214,N_9914);
and U10942 (N_10942,N_10071,N_10095);
or U10943 (N_10943,N_10371,N_9782);
and U10944 (N_10944,N_9846,N_10139);
nand U10945 (N_10945,N_10472,N_9775);
and U10946 (N_10946,N_9982,N_10489);
nor U10947 (N_10947,N_10048,N_10085);
nand U10948 (N_10948,N_10002,N_9943);
nand U10949 (N_10949,N_9913,N_9764);
and U10950 (N_10950,N_10196,N_10466);
and U10951 (N_10951,N_10349,N_9822);
and U10952 (N_10952,N_10172,N_9808);
or U10953 (N_10953,N_9763,N_10448);
nor U10954 (N_10954,N_10336,N_9931);
or U10955 (N_10955,N_9923,N_10211);
nand U10956 (N_10956,N_9811,N_10330);
or U10957 (N_10957,N_10140,N_9799);
or U10958 (N_10958,N_9999,N_9853);
or U10959 (N_10959,N_9941,N_10443);
nand U10960 (N_10960,N_10241,N_9991);
and U10961 (N_10961,N_9930,N_9890);
nand U10962 (N_10962,N_10490,N_9879);
nand U10963 (N_10963,N_10058,N_9798);
nor U10964 (N_10964,N_10144,N_10086);
nor U10965 (N_10965,N_9996,N_9791);
nand U10966 (N_10966,N_9804,N_9956);
nor U10967 (N_10967,N_10353,N_9931);
or U10968 (N_10968,N_10287,N_9770);
and U10969 (N_10969,N_10031,N_10250);
and U10970 (N_10970,N_10366,N_10069);
nor U10971 (N_10971,N_10409,N_9994);
and U10972 (N_10972,N_10263,N_10004);
nor U10973 (N_10973,N_9866,N_10022);
nand U10974 (N_10974,N_10140,N_10052);
and U10975 (N_10975,N_10180,N_10394);
nor U10976 (N_10976,N_9963,N_10458);
or U10977 (N_10977,N_10277,N_9804);
nand U10978 (N_10978,N_9837,N_10134);
or U10979 (N_10979,N_9754,N_10202);
and U10980 (N_10980,N_10333,N_10176);
nand U10981 (N_10981,N_10310,N_10093);
nand U10982 (N_10982,N_9888,N_10359);
or U10983 (N_10983,N_10384,N_9848);
nor U10984 (N_10984,N_10371,N_10325);
nor U10985 (N_10985,N_10017,N_10206);
nand U10986 (N_10986,N_9802,N_10461);
and U10987 (N_10987,N_9857,N_10328);
and U10988 (N_10988,N_10237,N_10281);
nor U10989 (N_10989,N_9938,N_9908);
or U10990 (N_10990,N_10091,N_10158);
and U10991 (N_10991,N_10326,N_10362);
nand U10992 (N_10992,N_10130,N_10013);
and U10993 (N_10993,N_9919,N_10401);
and U10994 (N_10994,N_10426,N_10419);
or U10995 (N_10995,N_10069,N_10056);
nand U10996 (N_10996,N_9772,N_9831);
or U10997 (N_10997,N_10004,N_9994);
or U10998 (N_10998,N_9995,N_9958);
nor U10999 (N_10999,N_9807,N_10170);
or U11000 (N_11000,N_10413,N_10411);
or U11001 (N_11001,N_10238,N_10283);
nor U11002 (N_11002,N_10041,N_10090);
and U11003 (N_11003,N_9875,N_10017);
nand U11004 (N_11004,N_10083,N_9926);
nor U11005 (N_11005,N_10419,N_9823);
and U11006 (N_11006,N_10063,N_10104);
nor U11007 (N_11007,N_9873,N_9891);
and U11008 (N_11008,N_10257,N_10285);
nor U11009 (N_11009,N_10065,N_9858);
nand U11010 (N_11010,N_9975,N_10325);
xnor U11011 (N_11011,N_10117,N_9768);
nand U11012 (N_11012,N_9760,N_10386);
or U11013 (N_11013,N_9991,N_9968);
nor U11014 (N_11014,N_10171,N_10013);
or U11015 (N_11015,N_10049,N_9908);
nand U11016 (N_11016,N_10261,N_10486);
nor U11017 (N_11017,N_9833,N_9958);
and U11018 (N_11018,N_9968,N_9871);
nor U11019 (N_11019,N_9885,N_10435);
nor U11020 (N_11020,N_10285,N_10365);
nand U11021 (N_11021,N_9758,N_9797);
nand U11022 (N_11022,N_9787,N_10018);
or U11023 (N_11023,N_10171,N_9976);
and U11024 (N_11024,N_9778,N_10200);
or U11025 (N_11025,N_9998,N_10376);
nor U11026 (N_11026,N_10412,N_9777);
nand U11027 (N_11027,N_9867,N_10445);
and U11028 (N_11028,N_10096,N_10411);
nand U11029 (N_11029,N_9959,N_9825);
and U11030 (N_11030,N_9841,N_10426);
nand U11031 (N_11031,N_10090,N_10448);
nand U11032 (N_11032,N_10228,N_9845);
or U11033 (N_11033,N_10403,N_10170);
nor U11034 (N_11034,N_9952,N_10403);
or U11035 (N_11035,N_9820,N_10043);
or U11036 (N_11036,N_10440,N_10139);
nor U11037 (N_11037,N_10377,N_10302);
and U11038 (N_11038,N_10494,N_10322);
nor U11039 (N_11039,N_10321,N_9836);
and U11040 (N_11040,N_9960,N_9935);
nand U11041 (N_11041,N_10008,N_9750);
and U11042 (N_11042,N_9840,N_10217);
nor U11043 (N_11043,N_10119,N_9952);
nand U11044 (N_11044,N_10086,N_10308);
nor U11045 (N_11045,N_9967,N_10445);
nand U11046 (N_11046,N_10071,N_10182);
nor U11047 (N_11047,N_9786,N_10450);
nand U11048 (N_11048,N_9909,N_10061);
nand U11049 (N_11049,N_9934,N_9898);
and U11050 (N_11050,N_9875,N_10463);
or U11051 (N_11051,N_10309,N_10001);
and U11052 (N_11052,N_9781,N_10413);
or U11053 (N_11053,N_10362,N_10240);
nor U11054 (N_11054,N_9964,N_9983);
and U11055 (N_11055,N_10282,N_10273);
or U11056 (N_11056,N_10225,N_9895);
and U11057 (N_11057,N_10310,N_10181);
or U11058 (N_11058,N_9866,N_10247);
and U11059 (N_11059,N_10365,N_10250);
nand U11060 (N_11060,N_10240,N_10227);
or U11061 (N_11061,N_10034,N_9911);
nand U11062 (N_11062,N_9915,N_10033);
and U11063 (N_11063,N_10334,N_10008);
nand U11064 (N_11064,N_10338,N_9903);
nor U11065 (N_11065,N_10406,N_9862);
or U11066 (N_11066,N_9758,N_10025);
or U11067 (N_11067,N_10184,N_10078);
and U11068 (N_11068,N_10499,N_9912);
or U11069 (N_11069,N_10474,N_10438);
or U11070 (N_11070,N_9812,N_9988);
nand U11071 (N_11071,N_9866,N_10191);
nor U11072 (N_11072,N_9762,N_10462);
and U11073 (N_11073,N_10010,N_10183);
nand U11074 (N_11074,N_10223,N_10469);
nor U11075 (N_11075,N_10048,N_10116);
and U11076 (N_11076,N_10338,N_9762);
or U11077 (N_11077,N_10489,N_10240);
and U11078 (N_11078,N_9776,N_10121);
nand U11079 (N_11079,N_9936,N_10208);
or U11080 (N_11080,N_10308,N_10224);
nand U11081 (N_11081,N_10401,N_10206);
nor U11082 (N_11082,N_9899,N_10163);
nand U11083 (N_11083,N_10073,N_9804);
nor U11084 (N_11084,N_9932,N_9884);
nand U11085 (N_11085,N_9760,N_9780);
and U11086 (N_11086,N_10301,N_9909);
or U11087 (N_11087,N_9870,N_9967);
and U11088 (N_11088,N_9994,N_10166);
nor U11089 (N_11089,N_10421,N_9773);
or U11090 (N_11090,N_10061,N_10160);
nand U11091 (N_11091,N_10175,N_9840);
nor U11092 (N_11092,N_9869,N_9987);
nand U11093 (N_11093,N_9915,N_10047);
nor U11094 (N_11094,N_10044,N_10287);
or U11095 (N_11095,N_10019,N_9934);
nor U11096 (N_11096,N_9947,N_10475);
nand U11097 (N_11097,N_9929,N_9885);
nand U11098 (N_11098,N_10341,N_10218);
nor U11099 (N_11099,N_10045,N_10227);
or U11100 (N_11100,N_10161,N_9875);
nand U11101 (N_11101,N_9906,N_9931);
nand U11102 (N_11102,N_10480,N_9973);
and U11103 (N_11103,N_9873,N_10331);
or U11104 (N_11104,N_9889,N_10474);
and U11105 (N_11105,N_10025,N_10434);
and U11106 (N_11106,N_10071,N_10412);
or U11107 (N_11107,N_10122,N_9916);
and U11108 (N_11108,N_10127,N_10319);
nand U11109 (N_11109,N_9963,N_9940);
nor U11110 (N_11110,N_10150,N_10197);
xnor U11111 (N_11111,N_10116,N_9893);
and U11112 (N_11112,N_10373,N_10038);
and U11113 (N_11113,N_9945,N_9814);
or U11114 (N_11114,N_9952,N_9987);
or U11115 (N_11115,N_9966,N_10284);
nor U11116 (N_11116,N_9856,N_10434);
nand U11117 (N_11117,N_10304,N_10480);
or U11118 (N_11118,N_9859,N_10035);
or U11119 (N_11119,N_9833,N_10077);
or U11120 (N_11120,N_9950,N_10440);
or U11121 (N_11121,N_10238,N_9797);
nand U11122 (N_11122,N_9805,N_10116);
or U11123 (N_11123,N_10059,N_10231);
or U11124 (N_11124,N_10383,N_10093);
and U11125 (N_11125,N_10270,N_10404);
or U11126 (N_11126,N_10365,N_10093);
xor U11127 (N_11127,N_9843,N_10373);
or U11128 (N_11128,N_10479,N_9962);
or U11129 (N_11129,N_9908,N_9812);
nor U11130 (N_11130,N_10377,N_10234);
or U11131 (N_11131,N_9762,N_10006);
nor U11132 (N_11132,N_9797,N_10092);
or U11133 (N_11133,N_9880,N_9995);
and U11134 (N_11134,N_9788,N_10182);
or U11135 (N_11135,N_10403,N_10128);
nor U11136 (N_11136,N_10471,N_10229);
nor U11137 (N_11137,N_10160,N_10134);
nand U11138 (N_11138,N_10238,N_10104);
nand U11139 (N_11139,N_10010,N_10225);
or U11140 (N_11140,N_10283,N_9767);
or U11141 (N_11141,N_10422,N_10061);
nor U11142 (N_11142,N_9935,N_10335);
or U11143 (N_11143,N_10263,N_10498);
and U11144 (N_11144,N_10470,N_10327);
nand U11145 (N_11145,N_10328,N_9757);
nand U11146 (N_11146,N_10371,N_10486);
nor U11147 (N_11147,N_9794,N_10417);
nand U11148 (N_11148,N_10455,N_9929);
nor U11149 (N_11149,N_9843,N_10360);
xor U11150 (N_11150,N_9890,N_9936);
nor U11151 (N_11151,N_10078,N_10334);
nand U11152 (N_11152,N_10356,N_10180);
nand U11153 (N_11153,N_10083,N_9860);
nand U11154 (N_11154,N_10034,N_9775);
or U11155 (N_11155,N_9922,N_9965);
nand U11156 (N_11156,N_10062,N_10362);
nor U11157 (N_11157,N_10121,N_10091);
and U11158 (N_11158,N_10369,N_9824);
nand U11159 (N_11159,N_9856,N_10400);
or U11160 (N_11160,N_10328,N_10442);
nand U11161 (N_11161,N_10278,N_10230);
nor U11162 (N_11162,N_9761,N_10294);
nor U11163 (N_11163,N_10361,N_10487);
and U11164 (N_11164,N_10253,N_10027);
and U11165 (N_11165,N_9980,N_10003);
or U11166 (N_11166,N_10215,N_10159);
nor U11167 (N_11167,N_9827,N_10177);
or U11168 (N_11168,N_10463,N_9950);
nand U11169 (N_11169,N_9985,N_10415);
nor U11170 (N_11170,N_10333,N_9867);
nor U11171 (N_11171,N_9956,N_9765);
and U11172 (N_11172,N_10285,N_10270);
nand U11173 (N_11173,N_10301,N_9807);
or U11174 (N_11174,N_10174,N_10062);
or U11175 (N_11175,N_9830,N_10417);
or U11176 (N_11176,N_10068,N_9904);
or U11177 (N_11177,N_9846,N_10215);
nand U11178 (N_11178,N_10236,N_10497);
and U11179 (N_11179,N_10021,N_10291);
nor U11180 (N_11180,N_9997,N_10440);
nand U11181 (N_11181,N_9869,N_10160);
xnor U11182 (N_11182,N_10442,N_10107);
or U11183 (N_11183,N_10255,N_10176);
and U11184 (N_11184,N_10383,N_10033);
and U11185 (N_11185,N_10021,N_10049);
or U11186 (N_11186,N_10350,N_10141);
nor U11187 (N_11187,N_9896,N_10312);
and U11188 (N_11188,N_10093,N_10067);
nand U11189 (N_11189,N_9807,N_9902);
nand U11190 (N_11190,N_9769,N_9970);
and U11191 (N_11191,N_9905,N_9995);
and U11192 (N_11192,N_10409,N_9768);
and U11193 (N_11193,N_10238,N_10404);
or U11194 (N_11194,N_10445,N_10158);
nand U11195 (N_11195,N_9774,N_9901);
or U11196 (N_11196,N_10164,N_9854);
nand U11197 (N_11197,N_9943,N_10079);
nor U11198 (N_11198,N_10467,N_9801);
or U11199 (N_11199,N_10070,N_9961);
nor U11200 (N_11200,N_9966,N_9830);
or U11201 (N_11201,N_10110,N_9818);
nor U11202 (N_11202,N_9890,N_10180);
nor U11203 (N_11203,N_9767,N_9861);
and U11204 (N_11204,N_9993,N_10295);
nor U11205 (N_11205,N_9927,N_10466);
xor U11206 (N_11206,N_9862,N_9763);
or U11207 (N_11207,N_10261,N_10408);
or U11208 (N_11208,N_9938,N_9874);
nor U11209 (N_11209,N_10444,N_9803);
or U11210 (N_11210,N_10162,N_10267);
nand U11211 (N_11211,N_10269,N_9967);
nor U11212 (N_11212,N_10409,N_10431);
nand U11213 (N_11213,N_10024,N_10401);
or U11214 (N_11214,N_10456,N_9878);
nand U11215 (N_11215,N_10191,N_10088);
xnor U11216 (N_11216,N_10094,N_10236);
nor U11217 (N_11217,N_9766,N_9762);
nand U11218 (N_11218,N_10141,N_9896);
or U11219 (N_11219,N_10192,N_10280);
and U11220 (N_11220,N_10313,N_10027);
nand U11221 (N_11221,N_10204,N_10447);
and U11222 (N_11222,N_10258,N_9771);
nand U11223 (N_11223,N_10060,N_9769);
and U11224 (N_11224,N_10316,N_10380);
or U11225 (N_11225,N_9811,N_10254);
or U11226 (N_11226,N_9992,N_10486);
nor U11227 (N_11227,N_10418,N_10051);
or U11228 (N_11228,N_10445,N_10223);
nand U11229 (N_11229,N_10330,N_9887);
and U11230 (N_11230,N_10118,N_9898);
nor U11231 (N_11231,N_10245,N_10064);
and U11232 (N_11232,N_9762,N_10387);
nor U11233 (N_11233,N_10439,N_10363);
nand U11234 (N_11234,N_9937,N_10427);
or U11235 (N_11235,N_10058,N_9813);
and U11236 (N_11236,N_10470,N_10386);
nor U11237 (N_11237,N_9835,N_10209);
nand U11238 (N_11238,N_10362,N_9754);
or U11239 (N_11239,N_10477,N_10334);
nor U11240 (N_11240,N_9791,N_9985);
nand U11241 (N_11241,N_9995,N_9977);
nand U11242 (N_11242,N_9922,N_10293);
nor U11243 (N_11243,N_10190,N_10290);
nand U11244 (N_11244,N_10279,N_9977);
and U11245 (N_11245,N_9831,N_10350);
and U11246 (N_11246,N_10319,N_9960);
nor U11247 (N_11247,N_9826,N_10124);
and U11248 (N_11248,N_10193,N_10081);
or U11249 (N_11249,N_9968,N_10469);
nand U11250 (N_11250,N_10827,N_10761);
or U11251 (N_11251,N_10590,N_10943);
nor U11252 (N_11252,N_10693,N_11082);
nand U11253 (N_11253,N_11119,N_10542);
or U11254 (N_11254,N_10909,N_11008);
and U11255 (N_11255,N_10661,N_11124);
or U11256 (N_11256,N_11074,N_10650);
and U11257 (N_11257,N_11175,N_11030);
and U11258 (N_11258,N_11021,N_10596);
or U11259 (N_11259,N_10981,N_10955);
nor U11260 (N_11260,N_10683,N_10531);
nand U11261 (N_11261,N_10830,N_11073);
nand U11262 (N_11262,N_10989,N_10824);
or U11263 (N_11263,N_11239,N_10715);
or U11264 (N_11264,N_10705,N_11229);
nand U11265 (N_11265,N_11240,N_11140);
and U11266 (N_11266,N_10828,N_11145);
nor U11267 (N_11267,N_10941,N_10740);
nor U11268 (N_11268,N_11069,N_11186);
nor U11269 (N_11269,N_11120,N_10626);
nor U11270 (N_11270,N_10518,N_10868);
or U11271 (N_11271,N_10887,N_10572);
xnor U11272 (N_11272,N_10832,N_10584);
nand U11273 (N_11273,N_10623,N_10805);
or U11274 (N_11274,N_10831,N_10569);
nor U11275 (N_11275,N_11224,N_10736);
nand U11276 (N_11276,N_10769,N_10587);
nor U11277 (N_11277,N_10894,N_11085);
nand U11278 (N_11278,N_11081,N_10781);
nor U11279 (N_11279,N_10651,N_10985);
or U11280 (N_11280,N_10525,N_11088);
nand U11281 (N_11281,N_10556,N_10956);
and U11282 (N_11282,N_10982,N_10822);
nor U11283 (N_11283,N_11153,N_10673);
or U11284 (N_11284,N_10557,N_10821);
nand U11285 (N_11285,N_10919,N_10706);
nor U11286 (N_11286,N_11003,N_10674);
nor U11287 (N_11287,N_10906,N_11206);
nor U11288 (N_11288,N_10599,N_10903);
and U11289 (N_11289,N_10561,N_10635);
or U11290 (N_11290,N_10534,N_10593);
and U11291 (N_11291,N_10809,N_10965);
nor U11292 (N_11292,N_11238,N_10928);
or U11293 (N_11293,N_11162,N_11109);
and U11294 (N_11294,N_11110,N_10806);
nand U11295 (N_11295,N_10767,N_10645);
nor U11296 (N_11296,N_10972,N_10775);
and U11297 (N_11297,N_10770,N_10864);
nor U11298 (N_11298,N_11084,N_10515);
or U11299 (N_11299,N_10627,N_10927);
or U11300 (N_11300,N_10966,N_10811);
and U11301 (N_11301,N_11004,N_10738);
nand U11302 (N_11302,N_10813,N_10753);
nor U11303 (N_11303,N_10984,N_10735);
nand U11304 (N_11304,N_10846,N_10664);
nand U11305 (N_11305,N_10792,N_11174);
nor U11306 (N_11306,N_11129,N_11149);
nand U11307 (N_11307,N_10737,N_11076);
nor U11308 (N_11308,N_10502,N_10964);
and U11309 (N_11309,N_10778,N_10672);
nor U11310 (N_11310,N_10883,N_10957);
nand U11311 (N_11311,N_10567,N_10568);
or U11312 (N_11312,N_11098,N_11080);
or U11313 (N_11313,N_10725,N_11198);
and U11314 (N_11314,N_10999,N_10891);
and U11315 (N_11315,N_11045,N_10639);
or U11316 (N_11316,N_10875,N_10657);
or U11317 (N_11317,N_11190,N_10527);
or U11318 (N_11318,N_10823,N_10577);
nor U11319 (N_11319,N_10871,N_11201);
xnor U11320 (N_11320,N_11007,N_11054);
or U11321 (N_11321,N_10698,N_11249);
or U11322 (N_11322,N_10837,N_10942);
and U11323 (N_11323,N_11043,N_10566);
nor U11324 (N_11324,N_10893,N_11099);
nor U11325 (N_11325,N_10520,N_10609);
or U11326 (N_11326,N_11115,N_10579);
or U11327 (N_11327,N_10659,N_10780);
nor U11328 (N_11328,N_10529,N_10930);
nor U11329 (N_11329,N_10773,N_10933);
and U11330 (N_11330,N_11134,N_10746);
and U11331 (N_11331,N_10717,N_10848);
nor U11332 (N_11332,N_11011,N_11068);
and U11333 (N_11333,N_11137,N_10558);
nand U11334 (N_11334,N_10851,N_10642);
and U11335 (N_11335,N_11049,N_11041);
and U11336 (N_11336,N_10797,N_11173);
nand U11337 (N_11337,N_11038,N_10656);
nor U11338 (N_11338,N_10631,N_10794);
or U11339 (N_11339,N_10583,N_10544);
or U11340 (N_11340,N_10829,N_10791);
nor U11341 (N_11341,N_11005,N_10712);
nand U11342 (N_11342,N_11237,N_10784);
nor U11343 (N_11343,N_11210,N_10582);
nor U11344 (N_11344,N_11023,N_10553);
nand U11345 (N_11345,N_11168,N_10872);
and U11346 (N_11346,N_11142,N_11188);
and U11347 (N_11347,N_10621,N_11169);
or U11348 (N_11348,N_11230,N_10905);
or U11349 (N_11349,N_11053,N_11170);
or U11350 (N_11350,N_10886,N_11086);
nand U11351 (N_11351,N_10597,N_10697);
nor U11352 (N_11352,N_10595,N_11079);
and U11353 (N_11353,N_11207,N_11136);
nand U11354 (N_11354,N_11101,N_10702);
and U11355 (N_11355,N_11058,N_11203);
and U11356 (N_11356,N_11245,N_10504);
or U11357 (N_11357,N_10853,N_10701);
nor U11358 (N_11358,N_11070,N_11111);
or U11359 (N_11359,N_10889,N_10611);
nand U11360 (N_11360,N_10793,N_10847);
nor U11361 (N_11361,N_11094,N_11220);
or U11362 (N_11362,N_10953,N_10812);
or U11363 (N_11363,N_10978,N_10990);
nor U11364 (N_11364,N_11143,N_10757);
and U11365 (N_11365,N_11225,N_10555);
nor U11366 (N_11366,N_11144,N_11231);
or U11367 (N_11367,N_10547,N_10779);
and U11368 (N_11368,N_10726,N_10947);
or U11369 (N_11369,N_10762,N_10676);
and U11370 (N_11370,N_11065,N_10714);
xnor U11371 (N_11371,N_10980,N_10900);
nor U11372 (N_11372,N_10898,N_10765);
nand U11373 (N_11373,N_10666,N_11218);
or U11374 (N_11374,N_10667,N_10517);
and U11375 (N_11375,N_11031,N_11107);
nor U11376 (N_11376,N_10692,N_10551);
and U11377 (N_11377,N_11091,N_11015);
and U11378 (N_11378,N_10731,N_11104);
or U11379 (N_11379,N_11171,N_10917);
or U11380 (N_11380,N_11095,N_10625);
nand U11381 (N_11381,N_10748,N_10968);
and U11382 (N_11382,N_11112,N_10749);
and U11383 (N_11383,N_11227,N_10854);
nor U11384 (N_11384,N_10739,N_11006);
and U11385 (N_11385,N_11184,N_11222);
and U11386 (N_11386,N_10546,N_10574);
xnor U11387 (N_11387,N_10804,N_10879);
and U11388 (N_11388,N_11044,N_10920);
and U11389 (N_11389,N_10637,N_10988);
nor U11390 (N_11390,N_10638,N_10818);
and U11391 (N_11391,N_11035,N_10888);
or U11392 (N_11392,N_10974,N_10573);
nand U11393 (N_11393,N_10810,N_10679);
and U11394 (N_11394,N_10799,N_11234);
nor U11395 (N_11395,N_10815,N_10663);
and U11396 (N_11396,N_10622,N_10633);
and U11397 (N_11397,N_11114,N_10973);
nor U11398 (N_11398,N_11146,N_10967);
nor U11399 (N_11399,N_10563,N_10899);
and U11400 (N_11400,N_10709,N_10616);
or U11401 (N_11401,N_11117,N_10533);
and U11402 (N_11402,N_11148,N_10653);
nor U11403 (N_11403,N_10742,N_10530);
nor U11404 (N_11404,N_11156,N_10850);
and U11405 (N_11405,N_10689,N_10992);
or U11406 (N_11406,N_10826,N_10862);
or U11407 (N_11407,N_10503,N_10509);
nand U11408 (N_11408,N_11017,N_10895);
nand U11409 (N_11409,N_10807,N_10764);
or U11410 (N_11410,N_10708,N_10758);
or U11411 (N_11411,N_10727,N_10925);
and U11412 (N_11412,N_11116,N_10877);
or U11413 (N_11413,N_11067,N_10858);
and U11414 (N_11414,N_10744,N_10628);
or U11415 (N_11415,N_11024,N_10840);
nand U11416 (N_11416,N_11236,N_10790);
nor U11417 (N_11417,N_11192,N_10641);
nand U11418 (N_11418,N_11241,N_10512);
or U11419 (N_11419,N_10922,N_11001);
nand U11420 (N_11420,N_10931,N_10820);
and U11421 (N_11421,N_11248,N_10685);
nand U11422 (N_11422,N_10844,N_10860);
and U11423 (N_11423,N_10695,N_11025);
nor U11424 (N_11424,N_10524,N_10729);
and U11425 (N_11425,N_10774,N_10662);
nand U11426 (N_11426,N_10669,N_10745);
or U11427 (N_11427,N_11193,N_10723);
and U11428 (N_11428,N_11150,N_11166);
or U11429 (N_11429,N_11215,N_10950);
and U11430 (N_11430,N_11185,N_10655);
nand U11431 (N_11431,N_10755,N_11177);
or U11432 (N_11432,N_10839,N_10677);
and U11433 (N_11433,N_10969,N_10940);
and U11434 (N_11434,N_10560,N_10733);
or U11435 (N_11435,N_10816,N_10924);
nor U11436 (N_11436,N_10934,N_11056);
nand U11437 (N_11437,N_10857,N_10722);
nor U11438 (N_11438,N_10977,N_10926);
and U11439 (N_11439,N_10771,N_11138);
nand U11440 (N_11440,N_10658,N_11200);
and U11441 (N_11441,N_10576,N_11059);
or U11442 (N_11442,N_11087,N_11046);
or U11443 (N_11443,N_10540,N_11057);
and U11444 (N_11444,N_11033,N_10814);
or U11445 (N_11445,N_11214,N_11176);
and U11446 (N_11446,N_10665,N_11100);
and U11447 (N_11447,N_10629,N_10766);
or U11448 (N_11448,N_10668,N_11194);
or U11449 (N_11449,N_10975,N_11232);
and U11450 (N_11450,N_11130,N_11055);
and U11451 (N_11451,N_10945,N_11147);
nand U11452 (N_11452,N_11092,N_11127);
or U11453 (N_11453,N_11040,N_10604);
xor U11454 (N_11454,N_11075,N_10852);
nor U11455 (N_11455,N_11118,N_11233);
and U11456 (N_11456,N_10798,N_10505);
nor U11457 (N_11457,N_10994,N_11014);
nand U11458 (N_11458,N_10976,N_10796);
nand U11459 (N_11459,N_11223,N_10939);
nor U11460 (N_11460,N_10588,N_10855);
nand U11461 (N_11461,N_10789,N_10719);
and U11462 (N_11462,N_10522,N_10591);
or U11463 (N_11463,N_10835,N_10526);
or U11464 (N_11464,N_10575,N_11189);
and U11465 (N_11465,N_10937,N_10983);
and U11466 (N_11466,N_11022,N_10537);
nor U11467 (N_11467,N_10949,N_11002);
nand U11468 (N_11468,N_10838,N_10648);
or U11469 (N_11469,N_10741,N_11018);
nor U11470 (N_11470,N_11126,N_10841);
or U11471 (N_11471,N_10506,N_10585);
nor U11472 (N_11472,N_10660,N_10720);
nor U11473 (N_11473,N_11243,N_10986);
and U11474 (N_11474,N_10690,N_10904);
or U11475 (N_11475,N_11205,N_11131);
and U11476 (N_11476,N_11122,N_10511);
nor U11477 (N_11477,N_11060,N_11202);
nand U11478 (N_11478,N_10795,N_11034);
or U11479 (N_11479,N_10682,N_10586);
nor U11480 (N_11480,N_10929,N_11219);
nand U11481 (N_11481,N_10699,N_10936);
and U11482 (N_11482,N_10721,N_11151);
and U11483 (N_11483,N_10594,N_11013);
or U11484 (N_11484,N_11152,N_10801);
and U11485 (N_11485,N_10911,N_10836);
nand U11486 (N_11486,N_10901,N_11213);
nand U11487 (N_11487,N_11113,N_10649);
or U11488 (N_11488,N_10550,N_11181);
and U11489 (N_11489,N_10600,N_10592);
nand U11490 (N_11490,N_11209,N_11036);
nand U11491 (N_11491,N_10747,N_10634);
nand U11492 (N_11492,N_11027,N_10787);
and U11493 (N_11493,N_10856,N_11009);
nor U11494 (N_11494,N_10866,N_10808);
or U11495 (N_11495,N_11196,N_10688);
nor U11496 (N_11496,N_11102,N_10777);
and U11497 (N_11497,N_10849,N_10549);
nor U11498 (N_11498,N_10918,N_11042);
nand U11499 (N_11499,N_10961,N_10863);
or U11500 (N_11500,N_10548,N_11204);
nand U11501 (N_11501,N_10958,N_10878);
or U11502 (N_11502,N_10552,N_10785);
nor U11503 (N_11503,N_10834,N_10508);
or U11504 (N_11504,N_10963,N_10754);
nor U11505 (N_11505,N_10786,N_10997);
nand U11506 (N_11506,N_10935,N_10885);
nor U11507 (N_11507,N_10681,N_10654);
nand U11508 (N_11508,N_11180,N_10865);
nor U11509 (N_11509,N_10896,N_10970);
nor U11510 (N_11510,N_10559,N_11244);
nor U11511 (N_11511,N_10734,N_10951);
or U11512 (N_11512,N_10914,N_11051);
and U11513 (N_11513,N_10962,N_10907);
nand U11514 (N_11514,N_10763,N_11048);
xnor U11515 (N_11515,N_11242,N_11216);
nor U11516 (N_11516,N_10516,N_11078);
nand U11517 (N_11517,N_10724,N_10716);
nand U11518 (N_11518,N_10678,N_11178);
and U11519 (N_11519,N_11106,N_10632);
or U11520 (N_11520,N_11155,N_10718);
and U11521 (N_11521,N_10691,N_10643);
nor U11522 (N_11522,N_10882,N_10539);
and U11523 (N_11523,N_10610,N_11063);
nor U11524 (N_11524,N_11064,N_11097);
and U11525 (N_11525,N_11029,N_11179);
or U11526 (N_11526,N_10687,N_10675);
nor U11527 (N_11527,N_10993,N_10845);
nor U11528 (N_11528,N_10536,N_10944);
nand U11529 (N_11529,N_10630,N_10908);
nor U11530 (N_11530,N_11195,N_10652);
and U11531 (N_11531,N_10759,N_10501);
or U11532 (N_11532,N_10680,N_10833);
nor U11533 (N_11533,N_10802,N_10783);
nor U11534 (N_11534,N_11172,N_11071);
and U11535 (N_11535,N_10694,N_10751);
or U11536 (N_11536,N_10636,N_11159);
and U11537 (N_11537,N_11226,N_11208);
nor U11538 (N_11538,N_10979,N_10843);
or U11539 (N_11539,N_11139,N_10601);
nor U11540 (N_11540,N_10580,N_10703);
or U11541 (N_11541,N_10768,N_10578);
nand U11542 (N_11542,N_10730,N_10646);
and U11543 (N_11543,N_10620,N_11183);
nand U11544 (N_11544,N_10910,N_11016);
nor U11545 (N_11545,N_10565,N_10644);
and U11546 (N_11546,N_11167,N_10874);
and U11547 (N_11547,N_11132,N_10605);
nor U11548 (N_11548,N_10897,N_10870);
or U11549 (N_11549,N_10528,N_10562);
or U11550 (N_11550,N_10523,N_10971);
nor U11551 (N_11551,N_10613,N_10817);
and U11552 (N_11552,N_10998,N_11246);
and U11553 (N_11553,N_10800,N_10684);
and U11554 (N_11554,N_11077,N_11191);
and U11555 (N_11555,N_10606,N_11211);
nand U11556 (N_11556,N_10615,N_10873);
nor U11557 (N_11557,N_10954,N_10869);
nand U11558 (N_11558,N_10500,N_10995);
nand U11559 (N_11559,N_10959,N_11039);
nor U11560 (N_11560,N_10880,N_10541);
nor U11561 (N_11561,N_11000,N_10987);
nor U11562 (N_11562,N_10603,N_10619);
nand U11563 (N_11563,N_10519,N_11066);
nand U11564 (N_11564,N_10624,N_10570);
and U11565 (N_11565,N_10960,N_10532);
nand U11566 (N_11566,N_10670,N_10612);
nor U11567 (N_11567,N_11133,N_10842);
nand U11568 (N_11568,N_11052,N_10617);
nand U11569 (N_11569,N_11221,N_10788);
nor U11570 (N_11570,N_11108,N_11154);
nand U11571 (N_11571,N_11128,N_11123);
or U11572 (N_11572,N_10732,N_10614);
nor U11573 (N_11573,N_10543,N_11093);
or U11574 (N_11574,N_11047,N_10756);
nor U11575 (N_11575,N_10598,N_10507);
and U11576 (N_11576,N_10890,N_10713);
and U11577 (N_11577,N_10696,N_10710);
nand U11578 (N_11578,N_11160,N_10607);
or U11579 (N_11579,N_10510,N_11182);
nor U11580 (N_11580,N_11103,N_11235);
nand U11581 (N_11581,N_10912,N_10819);
nand U11582 (N_11582,N_11187,N_11026);
or U11583 (N_11583,N_10946,N_10743);
nor U11584 (N_11584,N_10892,N_10513);
nand U11585 (N_11585,N_10825,N_11012);
or U11586 (N_11586,N_10752,N_11019);
nor U11587 (N_11587,N_10581,N_11163);
or U11588 (N_11588,N_11096,N_10952);
xor U11589 (N_11589,N_11199,N_10921);
nor U11590 (N_11590,N_10948,N_11164);
or U11591 (N_11591,N_11062,N_10521);
or U11592 (N_11592,N_10803,N_10867);
or U11593 (N_11593,N_10884,N_11089);
or U11594 (N_11594,N_11228,N_10571);
nand U11595 (N_11595,N_11061,N_10589);
and U11596 (N_11596,N_11217,N_10932);
nand U11597 (N_11597,N_10991,N_10538);
and U11598 (N_11598,N_10915,N_10772);
nor U11599 (N_11599,N_10640,N_11083);
nand U11600 (N_11600,N_11135,N_10618);
xnor U11601 (N_11601,N_11010,N_10996);
and U11602 (N_11602,N_10707,N_11247);
nand U11603 (N_11603,N_10728,N_11028);
nand U11604 (N_11604,N_11161,N_10902);
and U11605 (N_11605,N_11105,N_10750);
or U11606 (N_11606,N_11197,N_10881);
nor U11607 (N_11607,N_10923,N_11141);
and U11608 (N_11608,N_10647,N_10704);
xor U11609 (N_11609,N_11020,N_10776);
nor U11610 (N_11610,N_11125,N_10760);
nor U11611 (N_11611,N_10545,N_11090);
nand U11612 (N_11612,N_11158,N_11165);
and U11613 (N_11613,N_11050,N_10700);
nor U11614 (N_11614,N_10608,N_10876);
or U11615 (N_11615,N_10535,N_10859);
nand U11616 (N_11616,N_10686,N_10782);
or U11617 (N_11617,N_10602,N_11157);
or U11618 (N_11618,N_10671,N_11032);
nand U11619 (N_11619,N_10861,N_11212);
nand U11620 (N_11620,N_11072,N_11121);
and U11621 (N_11621,N_10554,N_10938);
nand U11622 (N_11622,N_11037,N_10916);
nor U11623 (N_11623,N_10514,N_10913);
and U11624 (N_11624,N_10711,N_10564);
or U11625 (N_11625,N_10517,N_10554);
or U11626 (N_11626,N_10571,N_10767);
and U11627 (N_11627,N_11063,N_11110);
nand U11628 (N_11628,N_10535,N_10655);
and U11629 (N_11629,N_10689,N_10554);
or U11630 (N_11630,N_11243,N_10981);
nand U11631 (N_11631,N_11151,N_10967);
or U11632 (N_11632,N_10807,N_11153);
nor U11633 (N_11633,N_10945,N_10806);
and U11634 (N_11634,N_10559,N_10940);
or U11635 (N_11635,N_11060,N_10949);
or U11636 (N_11636,N_10608,N_10524);
or U11637 (N_11637,N_10899,N_11114);
nor U11638 (N_11638,N_10775,N_11206);
nor U11639 (N_11639,N_10685,N_11223);
nand U11640 (N_11640,N_11093,N_10698);
and U11641 (N_11641,N_10999,N_10555);
or U11642 (N_11642,N_10527,N_10662);
and U11643 (N_11643,N_10603,N_11213);
or U11644 (N_11644,N_11130,N_10637);
nor U11645 (N_11645,N_10863,N_11113);
or U11646 (N_11646,N_11066,N_10613);
nand U11647 (N_11647,N_10844,N_11151);
or U11648 (N_11648,N_10876,N_10829);
nor U11649 (N_11649,N_10699,N_10955);
nor U11650 (N_11650,N_10538,N_10816);
nand U11651 (N_11651,N_11168,N_10547);
or U11652 (N_11652,N_11139,N_10610);
or U11653 (N_11653,N_10563,N_11223);
nand U11654 (N_11654,N_10643,N_10969);
nand U11655 (N_11655,N_10606,N_11208);
and U11656 (N_11656,N_11239,N_10801);
or U11657 (N_11657,N_10984,N_11245);
nor U11658 (N_11658,N_11132,N_11072);
and U11659 (N_11659,N_11144,N_10860);
or U11660 (N_11660,N_10581,N_10921);
or U11661 (N_11661,N_11177,N_10559);
and U11662 (N_11662,N_10783,N_11043);
and U11663 (N_11663,N_10857,N_10613);
or U11664 (N_11664,N_10734,N_10688);
and U11665 (N_11665,N_11104,N_11083);
and U11666 (N_11666,N_11226,N_11017);
nor U11667 (N_11667,N_10646,N_11157);
nor U11668 (N_11668,N_11156,N_10903);
nand U11669 (N_11669,N_10602,N_11209);
or U11670 (N_11670,N_10584,N_10687);
nand U11671 (N_11671,N_10744,N_10559);
or U11672 (N_11672,N_10631,N_11041);
and U11673 (N_11673,N_10615,N_10574);
nor U11674 (N_11674,N_11012,N_10902);
or U11675 (N_11675,N_10792,N_11166);
and U11676 (N_11676,N_10729,N_10544);
and U11677 (N_11677,N_10639,N_10780);
or U11678 (N_11678,N_10931,N_10923);
and U11679 (N_11679,N_11009,N_10825);
nor U11680 (N_11680,N_10840,N_10896);
nor U11681 (N_11681,N_10919,N_11154);
or U11682 (N_11682,N_11017,N_10553);
and U11683 (N_11683,N_10826,N_11247);
and U11684 (N_11684,N_10658,N_10785);
and U11685 (N_11685,N_10630,N_10769);
and U11686 (N_11686,N_10754,N_11091);
and U11687 (N_11687,N_11009,N_10982);
and U11688 (N_11688,N_10993,N_10968);
nand U11689 (N_11689,N_10993,N_10567);
nor U11690 (N_11690,N_11105,N_10681);
or U11691 (N_11691,N_10891,N_11141);
and U11692 (N_11692,N_10841,N_11248);
or U11693 (N_11693,N_11119,N_10514);
and U11694 (N_11694,N_10759,N_10728);
or U11695 (N_11695,N_10883,N_10512);
xnor U11696 (N_11696,N_10713,N_10711);
nor U11697 (N_11697,N_11205,N_11035);
or U11698 (N_11698,N_10985,N_11039);
or U11699 (N_11699,N_11083,N_10763);
nor U11700 (N_11700,N_10759,N_11236);
nand U11701 (N_11701,N_10557,N_10753);
nor U11702 (N_11702,N_11059,N_11151);
and U11703 (N_11703,N_10574,N_10658);
or U11704 (N_11704,N_10561,N_10865);
or U11705 (N_11705,N_11208,N_11014);
or U11706 (N_11706,N_11017,N_11139);
and U11707 (N_11707,N_11169,N_10819);
or U11708 (N_11708,N_10500,N_10742);
or U11709 (N_11709,N_11017,N_10619);
and U11710 (N_11710,N_11159,N_10527);
and U11711 (N_11711,N_10609,N_11197);
or U11712 (N_11712,N_10893,N_10515);
nor U11713 (N_11713,N_10910,N_10599);
and U11714 (N_11714,N_10574,N_10700);
nand U11715 (N_11715,N_10876,N_10639);
and U11716 (N_11716,N_10995,N_11139);
and U11717 (N_11717,N_10950,N_10884);
or U11718 (N_11718,N_10891,N_10808);
or U11719 (N_11719,N_10563,N_11084);
nor U11720 (N_11720,N_10684,N_11041);
nand U11721 (N_11721,N_10922,N_11024);
and U11722 (N_11722,N_10875,N_11166);
nor U11723 (N_11723,N_11098,N_10995);
nor U11724 (N_11724,N_11221,N_10545);
nand U11725 (N_11725,N_10734,N_10531);
and U11726 (N_11726,N_11126,N_11110);
or U11727 (N_11727,N_11037,N_11239);
nand U11728 (N_11728,N_10719,N_11149);
or U11729 (N_11729,N_10936,N_10988);
nor U11730 (N_11730,N_10745,N_10521);
nor U11731 (N_11731,N_10611,N_11057);
or U11732 (N_11732,N_11104,N_10720);
or U11733 (N_11733,N_10595,N_11163);
or U11734 (N_11734,N_11168,N_10514);
or U11735 (N_11735,N_10649,N_10991);
nand U11736 (N_11736,N_10634,N_10581);
nor U11737 (N_11737,N_10826,N_10692);
or U11738 (N_11738,N_10635,N_11117);
nand U11739 (N_11739,N_10931,N_10605);
nand U11740 (N_11740,N_11228,N_10553);
and U11741 (N_11741,N_10976,N_10613);
and U11742 (N_11742,N_10882,N_10860);
or U11743 (N_11743,N_10850,N_10679);
nand U11744 (N_11744,N_10571,N_11225);
and U11745 (N_11745,N_10500,N_10700);
nor U11746 (N_11746,N_10801,N_11180);
or U11747 (N_11747,N_10839,N_10648);
and U11748 (N_11748,N_10530,N_11084);
nor U11749 (N_11749,N_11072,N_10956);
nand U11750 (N_11750,N_10815,N_11205);
nand U11751 (N_11751,N_11092,N_10859);
nand U11752 (N_11752,N_11117,N_10545);
nor U11753 (N_11753,N_10666,N_10782);
or U11754 (N_11754,N_11015,N_10587);
nand U11755 (N_11755,N_10631,N_11093);
or U11756 (N_11756,N_10668,N_11202);
nand U11757 (N_11757,N_11197,N_11028);
nand U11758 (N_11758,N_10615,N_10863);
or U11759 (N_11759,N_10651,N_10862);
nand U11760 (N_11760,N_11063,N_11179);
nand U11761 (N_11761,N_11248,N_10613);
and U11762 (N_11762,N_10763,N_10909);
and U11763 (N_11763,N_10544,N_10684);
nor U11764 (N_11764,N_10621,N_10678);
nor U11765 (N_11765,N_10541,N_10572);
nand U11766 (N_11766,N_10849,N_10672);
nor U11767 (N_11767,N_10538,N_10762);
or U11768 (N_11768,N_11041,N_10648);
xor U11769 (N_11769,N_10871,N_10700);
or U11770 (N_11770,N_10873,N_11168);
nand U11771 (N_11771,N_11062,N_11067);
nand U11772 (N_11772,N_11010,N_11039);
nand U11773 (N_11773,N_10538,N_10550);
or U11774 (N_11774,N_10725,N_10778);
or U11775 (N_11775,N_10758,N_10631);
and U11776 (N_11776,N_10644,N_10617);
or U11777 (N_11777,N_10581,N_10550);
nor U11778 (N_11778,N_10876,N_11078);
or U11779 (N_11779,N_11236,N_11061);
and U11780 (N_11780,N_11160,N_10630);
nand U11781 (N_11781,N_11201,N_10543);
nand U11782 (N_11782,N_10920,N_10581);
and U11783 (N_11783,N_11169,N_10575);
or U11784 (N_11784,N_11230,N_11085);
or U11785 (N_11785,N_11116,N_10830);
nor U11786 (N_11786,N_10670,N_11181);
or U11787 (N_11787,N_10794,N_10948);
nand U11788 (N_11788,N_10835,N_11080);
nand U11789 (N_11789,N_10866,N_10897);
nand U11790 (N_11790,N_10709,N_11111);
and U11791 (N_11791,N_10629,N_10701);
nor U11792 (N_11792,N_10759,N_10826);
nand U11793 (N_11793,N_11126,N_10753);
or U11794 (N_11794,N_10633,N_10585);
nor U11795 (N_11795,N_11075,N_11123);
nor U11796 (N_11796,N_11112,N_10521);
or U11797 (N_11797,N_11035,N_10566);
nor U11798 (N_11798,N_11063,N_10673);
nand U11799 (N_11799,N_11094,N_10746);
and U11800 (N_11800,N_10677,N_10737);
or U11801 (N_11801,N_10681,N_10514);
nand U11802 (N_11802,N_10865,N_10510);
nand U11803 (N_11803,N_10985,N_10779);
or U11804 (N_11804,N_11119,N_10594);
or U11805 (N_11805,N_10579,N_11051);
or U11806 (N_11806,N_10976,N_11088);
and U11807 (N_11807,N_10522,N_10590);
and U11808 (N_11808,N_11141,N_10611);
nor U11809 (N_11809,N_10625,N_11212);
nand U11810 (N_11810,N_10777,N_10932);
or U11811 (N_11811,N_11043,N_10794);
nand U11812 (N_11812,N_11026,N_10650);
and U11813 (N_11813,N_10769,N_11143);
nand U11814 (N_11814,N_10645,N_10504);
and U11815 (N_11815,N_10895,N_10710);
and U11816 (N_11816,N_10978,N_10937);
or U11817 (N_11817,N_11081,N_10597);
and U11818 (N_11818,N_10882,N_11013);
or U11819 (N_11819,N_11146,N_10960);
nand U11820 (N_11820,N_10889,N_10615);
nand U11821 (N_11821,N_10794,N_10532);
and U11822 (N_11822,N_10987,N_10533);
nand U11823 (N_11823,N_10517,N_10811);
nor U11824 (N_11824,N_10725,N_10830);
nor U11825 (N_11825,N_10818,N_10836);
nand U11826 (N_11826,N_10809,N_10848);
nand U11827 (N_11827,N_10792,N_11014);
and U11828 (N_11828,N_10782,N_10949);
and U11829 (N_11829,N_10848,N_10571);
nand U11830 (N_11830,N_10884,N_10934);
nor U11831 (N_11831,N_10908,N_10550);
or U11832 (N_11832,N_11134,N_10612);
nor U11833 (N_11833,N_10919,N_11070);
or U11834 (N_11834,N_10530,N_10978);
nand U11835 (N_11835,N_11037,N_10869);
and U11836 (N_11836,N_10714,N_11027);
or U11837 (N_11837,N_10825,N_11023);
nor U11838 (N_11838,N_10829,N_11151);
nand U11839 (N_11839,N_10926,N_10576);
nand U11840 (N_11840,N_10661,N_10729);
and U11841 (N_11841,N_10734,N_10892);
and U11842 (N_11842,N_11033,N_10971);
nor U11843 (N_11843,N_11112,N_10740);
or U11844 (N_11844,N_10705,N_10911);
nand U11845 (N_11845,N_10511,N_10696);
and U11846 (N_11846,N_10629,N_10985);
nor U11847 (N_11847,N_10815,N_11039);
and U11848 (N_11848,N_11149,N_10550);
nor U11849 (N_11849,N_10920,N_11215);
and U11850 (N_11850,N_11005,N_10733);
or U11851 (N_11851,N_10647,N_11193);
nand U11852 (N_11852,N_10811,N_10604);
and U11853 (N_11853,N_11202,N_10511);
or U11854 (N_11854,N_11150,N_10645);
and U11855 (N_11855,N_10581,N_10654);
xor U11856 (N_11856,N_10692,N_10533);
or U11857 (N_11857,N_11163,N_11043);
or U11858 (N_11858,N_11078,N_10517);
nand U11859 (N_11859,N_11244,N_10802);
nand U11860 (N_11860,N_11216,N_11178);
nand U11861 (N_11861,N_10631,N_11187);
nor U11862 (N_11862,N_10686,N_10581);
and U11863 (N_11863,N_10955,N_10637);
and U11864 (N_11864,N_10630,N_10512);
and U11865 (N_11865,N_10697,N_10755);
and U11866 (N_11866,N_10795,N_11176);
nand U11867 (N_11867,N_10950,N_10647);
nor U11868 (N_11868,N_10980,N_10881);
nand U11869 (N_11869,N_10729,N_10533);
or U11870 (N_11870,N_11227,N_10781);
and U11871 (N_11871,N_10852,N_11018);
nand U11872 (N_11872,N_11160,N_11187);
and U11873 (N_11873,N_10941,N_11010);
nor U11874 (N_11874,N_11081,N_10553);
nor U11875 (N_11875,N_10998,N_11050);
and U11876 (N_11876,N_11235,N_10804);
nor U11877 (N_11877,N_10728,N_10914);
nor U11878 (N_11878,N_10797,N_11107);
nand U11879 (N_11879,N_10821,N_10742);
nor U11880 (N_11880,N_10500,N_10901);
or U11881 (N_11881,N_11171,N_10677);
and U11882 (N_11882,N_10657,N_11207);
and U11883 (N_11883,N_10858,N_10671);
and U11884 (N_11884,N_10661,N_10683);
nand U11885 (N_11885,N_10872,N_10621);
nor U11886 (N_11886,N_10985,N_11181);
nand U11887 (N_11887,N_10721,N_10769);
nor U11888 (N_11888,N_10592,N_10567);
and U11889 (N_11889,N_10641,N_10568);
xnor U11890 (N_11890,N_10586,N_10936);
nand U11891 (N_11891,N_11087,N_10895);
nor U11892 (N_11892,N_10797,N_10672);
xnor U11893 (N_11893,N_11081,N_10605);
or U11894 (N_11894,N_11211,N_10815);
nor U11895 (N_11895,N_10965,N_10691);
nor U11896 (N_11896,N_11104,N_10968);
nor U11897 (N_11897,N_10652,N_10706);
nor U11898 (N_11898,N_11123,N_10872);
xnor U11899 (N_11899,N_11106,N_11061);
nand U11900 (N_11900,N_10609,N_10906);
nor U11901 (N_11901,N_10546,N_10977);
nand U11902 (N_11902,N_10963,N_10870);
nor U11903 (N_11903,N_11007,N_10755);
or U11904 (N_11904,N_10649,N_10773);
or U11905 (N_11905,N_11014,N_10860);
nor U11906 (N_11906,N_11199,N_10720);
or U11907 (N_11907,N_11160,N_11072);
nor U11908 (N_11908,N_10945,N_10599);
nor U11909 (N_11909,N_11039,N_10998);
nand U11910 (N_11910,N_10943,N_10635);
and U11911 (N_11911,N_10684,N_10803);
xor U11912 (N_11912,N_10538,N_11202);
and U11913 (N_11913,N_10536,N_10505);
or U11914 (N_11914,N_10885,N_11028);
or U11915 (N_11915,N_10951,N_10557);
xor U11916 (N_11916,N_10859,N_10736);
nand U11917 (N_11917,N_10804,N_10851);
and U11918 (N_11918,N_10977,N_11139);
nand U11919 (N_11919,N_10686,N_10636);
nor U11920 (N_11920,N_10920,N_11153);
nor U11921 (N_11921,N_10549,N_10704);
nor U11922 (N_11922,N_10626,N_10910);
nor U11923 (N_11923,N_10729,N_10689);
or U11924 (N_11924,N_10952,N_10778);
and U11925 (N_11925,N_10753,N_10703);
nand U11926 (N_11926,N_10590,N_10939);
or U11927 (N_11927,N_11241,N_11047);
and U11928 (N_11928,N_10746,N_10966);
nand U11929 (N_11929,N_10907,N_11077);
nand U11930 (N_11930,N_10888,N_10672);
or U11931 (N_11931,N_11042,N_10527);
nor U11932 (N_11932,N_10820,N_10662);
nor U11933 (N_11933,N_11186,N_10530);
nand U11934 (N_11934,N_10903,N_11000);
nand U11935 (N_11935,N_11102,N_10751);
nand U11936 (N_11936,N_10791,N_10808);
and U11937 (N_11937,N_10910,N_10522);
nor U11938 (N_11938,N_10527,N_10798);
and U11939 (N_11939,N_11223,N_10816);
nor U11940 (N_11940,N_11016,N_11199);
or U11941 (N_11941,N_10698,N_10521);
nor U11942 (N_11942,N_10885,N_11222);
nand U11943 (N_11943,N_11064,N_10850);
nand U11944 (N_11944,N_10614,N_10962);
nand U11945 (N_11945,N_10927,N_11088);
nor U11946 (N_11946,N_11006,N_10946);
nand U11947 (N_11947,N_11137,N_11167);
and U11948 (N_11948,N_10764,N_11074);
and U11949 (N_11949,N_11195,N_10722);
nand U11950 (N_11950,N_10998,N_11240);
and U11951 (N_11951,N_11101,N_10532);
and U11952 (N_11952,N_10599,N_10789);
and U11953 (N_11953,N_11010,N_10959);
and U11954 (N_11954,N_11061,N_11091);
nand U11955 (N_11955,N_10987,N_10677);
or U11956 (N_11956,N_10740,N_10612);
and U11957 (N_11957,N_10699,N_10921);
and U11958 (N_11958,N_11228,N_11133);
and U11959 (N_11959,N_11027,N_10679);
nand U11960 (N_11960,N_11064,N_11157);
or U11961 (N_11961,N_10754,N_10875);
nor U11962 (N_11962,N_11041,N_10784);
and U11963 (N_11963,N_10984,N_11188);
or U11964 (N_11964,N_11135,N_11049);
and U11965 (N_11965,N_11232,N_11091);
nand U11966 (N_11966,N_11171,N_10564);
nand U11967 (N_11967,N_10683,N_11198);
and U11968 (N_11968,N_10778,N_10947);
nand U11969 (N_11969,N_11129,N_10595);
and U11970 (N_11970,N_10826,N_10964);
nand U11971 (N_11971,N_10646,N_11007);
and U11972 (N_11972,N_10972,N_10759);
nor U11973 (N_11973,N_11197,N_11070);
or U11974 (N_11974,N_10659,N_11094);
and U11975 (N_11975,N_11003,N_10747);
nor U11976 (N_11976,N_10856,N_11205);
or U11977 (N_11977,N_10524,N_10868);
and U11978 (N_11978,N_10800,N_10565);
nand U11979 (N_11979,N_11139,N_10602);
and U11980 (N_11980,N_11233,N_10891);
or U11981 (N_11981,N_11162,N_10645);
nor U11982 (N_11982,N_10557,N_10906);
nor U11983 (N_11983,N_11173,N_10556);
and U11984 (N_11984,N_10510,N_11008);
nand U11985 (N_11985,N_10911,N_10650);
nor U11986 (N_11986,N_10565,N_11015);
or U11987 (N_11987,N_11246,N_11170);
or U11988 (N_11988,N_10851,N_10697);
and U11989 (N_11989,N_10716,N_11083);
and U11990 (N_11990,N_10595,N_10709);
nor U11991 (N_11991,N_11001,N_10789);
or U11992 (N_11992,N_11174,N_10889);
nor U11993 (N_11993,N_11011,N_10958);
or U11994 (N_11994,N_11070,N_10733);
or U11995 (N_11995,N_10719,N_10794);
and U11996 (N_11996,N_10715,N_11189);
nor U11997 (N_11997,N_10769,N_10991);
nor U11998 (N_11998,N_10958,N_10716);
and U11999 (N_11999,N_10777,N_10566);
nand U12000 (N_12000,N_11772,N_11811);
or U12001 (N_12001,N_11611,N_11318);
nor U12002 (N_12002,N_11264,N_11769);
and U12003 (N_12003,N_11797,N_11253);
nand U12004 (N_12004,N_11274,N_11537);
or U12005 (N_12005,N_11900,N_11935);
or U12006 (N_12006,N_11677,N_11407);
and U12007 (N_12007,N_11712,N_11429);
nand U12008 (N_12008,N_11363,N_11637);
and U12009 (N_12009,N_11905,N_11566);
or U12010 (N_12010,N_11721,N_11853);
nand U12011 (N_12011,N_11970,N_11685);
or U12012 (N_12012,N_11804,N_11449);
nand U12013 (N_12013,N_11918,N_11865);
or U12014 (N_12014,N_11728,N_11377);
and U12015 (N_12015,N_11827,N_11436);
nor U12016 (N_12016,N_11636,N_11679);
and U12017 (N_12017,N_11846,N_11767);
nand U12018 (N_12018,N_11939,N_11945);
nand U12019 (N_12019,N_11604,N_11349);
nand U12020 (N_12020,N_11932,N_11366);
nand U12021 (N_12021,N_11940,N_11831);
nor U12022 (N_12022,N_11575,N_11285);
nor U12023 (N_12023,N_11718,N_11780);
and U12024 (N_12024,N_11740,N_11508);
and U12025 (N_12025,N_11507,N_11825);
nand U12026 (N_12026,N_11373,N_11713);
nor U12027 (N_12027,N_11787,N_11936);
nor U12028 (N_12028,N_11464,N_11505);
nor U12029 (N_12029,N_11334,N_11454);
nand U12030 (N_12030,N_11589,N_11708);
nand U12031 (N_12031,N_11823,N_11541);
and U12032 (N_12032,N_11852,N_11977);
and U12033 (N_12033,N_11903,N_11896);
and U12034 (N_12034,N_11697,N_11837);
or U12035 (N_12035,N_11961,N_11327);
nand U12036 (N_12036,N_11869,N_11529);
nand U12037 (N_12037,N_11564,N_11822);
nand U12038 (N_12038,N_11473,N_11562);
and U12039 (N_12039,N_11714,N_11886);
nand U12040 (N_12040,N_11283,N_11319);
nor U12041 (N_12041,N_11821,N_11969);
or U12042 (N_12042,N_11314,N_11751);
or U12043 (N_12043,N_11578,N_11286);
nand U12044 (N_12044,N_11581,N_11979);
nand U12045 (N_12045,N_11549,N_11983);
and U12046 (N_12046,N_11661,N_11615);
and U12047 (N_12047,N_11587,N_11756);
nor U12048 (N_12048,N_11870,N_11676);
and U12049 (N_12049,N_11986,N_11862);
or U12050 (N_12050,N_11388,N_11576);
or U12051 (N_12051,N_11660,N_11843);
and U12052 (N_12052,N_11262,N_11616);
nor U12053 (N_12053,N_11948,N_11813);
and U12054 (N_12054,N_11364,N_11659);
nor U12055 (N_12055,N_11799,N_11462);
and U12056 (N_12056,N_11622,N_11665);
or U12057 (N_12057,N_11923,N_11795);
nand U12058 (N_12058,N_11739,N_11331);
nand U12059 (N_12059,N_11968,N_11880);
and U12060 (N_12060,N_11536,N_11384);
or U12061 (N_12061,N_11858,N_11893);
nand U12062 (N_12062,N_11744,N_11819);
nor U12063 (N_12063,N_11810,N_11764);
or U12064 (N_12064,N_11488,N_11450);
nand U12065 (N_12065,N_11544,N_11674);
nor U12066 (N_12066,N_11621,N_11614);
or U12067 (N_12067,N_11806,N_11350);
or U12068 (N_12068,N_11733,N_11394);
and U12069 (N_12069,N_11548,N_11269);
and U12070 (N_12070,N_11402,N_11758);
nand U12071 (N_12071,N_11890,N_11609);
nor U12072 (N_12072,N_11586,N_11872);
nor U12073 (N_12073,N_11493,N_11704);
nand U12074 (N_12074,N_11761,N_11856);
and U12075 (N_12075,N_11812,N_11592);
nand U12076 (N_12076,N_11671,N_11854);
xnor U12077 (N_12077,N_11626,N_11376);
nand U12078 (N_12078,N_11382,N_11291);
and U12079 (N_12079,N_11563,N_11469);
nand U12080 (N_12080,N_11747,N_11398);
xor U12081 (N_12081,N_11686,N_11330);
nor U12082 (N_12082,N_11421,N_11642);
nor U12083 (N_12083,N_11259,N_11496);
and U12084 (N_12084,N_11460,N_11399);
nor U12085 (N_12085,N_11666,N_11989);
nor U12086 (N_12086,N_11768,N_11315);
and U12087 (N_12087,N_11420,N_11284);
and U12088 (N_12088,N_11328,N_11754);
or U12089 (N_12089,N_11683,N_11908);
and U12090 (N_12090,N_11500,N_11297);
or U12091 (N_12091,N_11667,N_11675);
nand U12092 (N_12092,N_11783,N_11838);
or U12093 (N_12093,N_11332,N_11424);
or U12094 (N_12094,N_11922,N_11802);
or U12095 (N_12095,N_11290,N_11835);
nand U12096 (N_12096,N_11702,N_11414);
or U12097 (N_12097,N_11289,N_11648);
or U12098 (N_12098,N_11278,N_11931);
nor U12099 (N_12099,N_11913,N_11478);
nor U12100 (N_12100,N_11817,N_11727);
nor U12101 (N_12101,N_11580,N_11486);
nor U12102 (N_12102,N_11796,N_11498);
nor U12103 (N_12103,N_11694,N_11574);
or U12104 (N_12104,N_11624,N_11958);
nand U12105 (N_12105,N_11742,N_11689);
and U12106 (N_12106,N_11816,N_11395);
nor U12107 (N_12107,N_11426,N_11620);
nand U12108 (N_12108,N_11401,N_11670);
or U12109 (N_12109,N_11474,N_11818);
and U12110 (N_12110,N_11326,N_11656);
and U12111 (N_12111,N_11565,N_11506);
or U12112 (N_12112,N_11465,N_11554);
and U12113 (N_12113,N_11730,N_11387);
nand U12114 (N_12114,N_11551,N_11260);
nand U12115 (N_12115,N_11413,N_11947);
and U12116 (N_12116,N_11658,N_11513);
and U12117 (N_12117,N_11834,N_11725);
nor U12118 (N_12118,N_11381,N_11801);
and U12119 (N_12119,N_11270,N_11515);
nor U12120 (N_12120,N_11815,N_11898);
or U12121 (N_12121,N_11791,N_11484);
nor U12122 (N_12122,N_11568,N_11706);
nand U12123 (N_12123,N_11993,N_11746);
or U12124 (N_12124,N_11850,N_11271);
nor U12125 (N_12125,N_11800,N_11311);
nand U12126 (N_12126,N_11552,N_11926);
and U12127 (N_12127,N_11964,N_11809);
nor U12128 (N_12128,N_11427,N_11999);
or U12129 (N_12129,N_11527,N_11481);
or U12130 (N_12130,N_11955,N_11298);
nand U12131 (N_12131,N_11530,N_11982);
or U12132 (N_12132,N_11444,N_11276);
and U12133 (N_12133,N_11409,N_11577);
and U12134 (N_12134,N_11655,N_11316);
nand U12135 (N_12135,N_11836,N_11902);
or U12136 (N_12136,N_11994,N_11597);
nand U12137 (N_12137,N_11663,N_11494);
nand U12138 (N_12138,N_11601,N_11695);
and U12139 (N_12139,N_11645,N_11353);
and U12140 (N_12140,N_11638,N_11531);
or U12141 (N_12141,N_11995,N_11790);
nand U12142 (N_12142,N_11960,N_11690);
or U12143 (N_12143,N_11786,N_11651);
nand U12144 (N_12144,N_11630,N_11881);
nor U12145 (N_12145,N_11520,N_11774);
and U12146 (N_12146,N_11504,N_11406);
and U12147 (N_12147,N_11653,N_11512);
nor U12148 (N_12148,N_11534,N_11482);
and U12149 (N_12149,N_11847,N_11897);
nor U12150 (N_12150,N_11591,N_11419);
nand U12151 (N_12151,N_11699,N_11347);
and U12152 (N_12152,N_11914,N_11701);
nor U12153 (N_12153,N_11405,N_11859);
nor U12154 (N_12154,N_11613,N_11803);
nand U12155 (N_12155,N_11480,N_11990);
nand U12156 (N_12156,N_11963,N_11627);
nor U12157 (N_12157,N_11573,N_11770);
and U12158 (N_12158,N_11499,N_11781);
nor U12159 (N_12159,N_11720,N_11807);
and U12160 (N_12160,N_11357,N_11719);
and U12161 (N_12161,N_11383,N_11703);
or U12162 (N_12162,N_11523,N_11631);
nand U12163 (N_12163,N_11680,N_11288);
nand U12164 (N_12164,N_11313,N_11771);
and U12165 (N_12165,N_11943,N_11974);
nand U12166 (N_12166,N_11841,N_11299);
nand U12167 (N_12167,N_11370,N_11673);
nand U12168 (N_12168,N_11477,N_11555);
nor U12169 (N_12169,N_11403,N_11973);
or U12170 (N_12170,N_11662,N_11681);
nor U12171 (N_12171,N_11441,N_11833);
nand U12172 (N_12172,N_11985,N_11877);
nand U12173 (N_12173,N_11337,N_11501);
or U12174 (N_12174,N_11250,N_11678);
nand U12175 (N_12175,N_11844,N_11321);
nor U12176 (N_12176,N_11468,N_11367);
nand U12177 (N_12177,N_11851,N_11691);
or U12178 (N_12178,N_11682,N_11792);
nand U12179 (N_12179,N_11304,N_11752);
and U12180 (N_12180,N_11561,N_11418);
or U12181 (N_12181,N_11503,N_11491);
nor U12182 (N_12182,N_11700,N_11348);
nand U12183 (N_12183,N_11981,N_11607);
or U12184 (N_12184,N_11976,N_11687);
xnor U12185 (N_12185,N_11866,N_11972);
or U12186 (N_12186,N_11322,N_11365);
or U12187 (N_12187,N_11845,N_11798);
nor U12188 (N_12188,N_11924,N_11617);
nor U12189 (N_12189,N_11602,N_11535);
or U12190 (N_12190,N_11839,N_11710);
and U12191 (N_12191,N_11997,N_11878);
nor U12192 (N_12192,N_11475,N_11448);
nor U12193 (N_12193,N_11855,N_11391);
and U12194 (N_12194,N_11916,N_11526);
and U12195 (N_12195,N_11594,N_11723);
or U12196 (N_12196,N_11988,N_11649);
nand U12197 (N_12197,N_11891,N_11868);
nand U12198 (N_12198,N_11268,N_11765);
nor U12199 (N_12199,N_11778,N_11921);
nand U12200 (N_12200,N_11492,N_11510);
and U12201 (N_12201,N_11652,N_11542);
nor U12202 (N_12202,N_11273,N_11389);
nand U12203 (N_12203,N_11688,N_11455);
or U12204 (N_12204,N_11832,N_11863);
and U12205 (N_12205,N_11867,N_11635);
nand U12206 (N_12206,N_11608,N_11292);
or U12207 (N_12207,N_11571,N_11282);
nor U12208 (N_12208,N_11934,N_11550);
xor U12209 (N_12209,N_11775,N_11920);
nand U12210 (N_12210,N_11452,N_11632);
nand U12211 (N_12211,N_11830,N_11814);
nand U12212 (N_12212,N_11709,N_11476);
or U12213 (N_12213,N_11466,N_11805);
and U12214 (N_12214,N_11749,N_11623);
nor U12215 (N_12215,N_11397,N_11303);
or U12216 (N_12216,N_11459,N_11996);
nor U12217 (N_12217,N_11335,N_11415);
and U12218 (N_12218,N_11748,N_11495);
nand U12219 (N_12219,N_11912,N_11762);
nor U12220 (N_12220,N_11559,N_11485);
nor U12221 (N_12221,N_11371,N_11640);
nand U12222 (N_12222,N_11490,N_11483);
nand U12223 (N_12223,N_11416,N_11600);
and U12224 (N_12224,N_11957,N_11669);
or U12225 (N_12225,N_11471,N_11430);
or U12226 (N_12226,N_11603,N_11309);
nand U12227 (N_12227,N_11808,N_11431);
xnor U12228 (N_12228,N_11650,N_11967);
nor U12229 (N_12229,N_11951,N_11522);
nand U12230 (N_12230,N_11287,N_11840);
nor U12231 (N_12231,N_11295,N_11511);
nand U12232 (N_12232,N_11518,N_11343);
nand U12233 (N_12233,N_11338,N_11412);
nor U12234 (N_12234,N_11975,N_11378);
or U12235 (N_12235,N_11323,N_11784);
nor U12236 (N_12236,N_11447,N_11528);
and U12237 (N_12237,N_11252,N_11938);
nand U12238 (N_12238,N_11711,N_11301);
nand U12239 (N_12239,N_11556,N_11788);
and U12240 (N_12240,N_11785,N_11737);
and U12241 (N_12241,N_11582,N_11255);
or U12242 (N_12242,N_11567,N_11992);
nor U12243 (N_12243,N_11824,N_11472);
and U12244 (N_12244,N_11928,N_11876);
or U12245 (N_12245,N_11759,N_11705);
or U12246 (N_12246,N_11917,N_11950);
or U12247 (N_12247,N_11857,N_11991);
nor U12248 (N_12248,N_11716,N_11606);
or U12249 (N_12249,N_11915,N_11425);
nor U12250 (N_12250,N_11306,N_11610);
nand U12251 (N_12251,N_11984,N_11553);
nand U12252 (N_12252,N_11386,N_11339);
or U12253 (N_12253,N_11467,N_11646);
nand U12254 (N_12254,N_11829,N_11417);
or U12255 (N_12255,N_11352,N_11341);
nor U12256 (N_12256,N_11453,N_11354);
or U12257 (N_12257,N_11965,N_11693);
nand U12258 (N_12258,N_11849,N_11410);
or U12259 (N_12259,N_11433,N_11873);
or U12260 (N_12260,N_11598,N_11432);
and U12261 (N_12261,N_11722,N_11296);
or U12262 (N_12262,N_11875,N_11572);
and U12263 (N_12263,N_11533,N_11910);
nor U12264 (N_12264,N_11539,N_11618);
and U12265 (N_12265,N_11351,N_11692);
and U12266 (N_12266,N_11628,N_11281);
or U12267 (N_12267,N_11525,N_11595);
nor U12268 (N_12268,N_11547,N_11509);
and U12269 (N_12269,N_11929,N_11585);
and U12270 (N_12270,N_11599,N_11736);
or U12271 (N_12271,N_11445,N_11446);
or U12272 (N_12272,N_11435,N_11633);
and U12273 (N_12273,N_11941,N_11317);
and U12274 (N_12274,N_11346,N_11753);
nor U12275 (N_12275,N_11664,N_11442);
nor U12276 (N_12276,N_11361,N_11324);
or U12277 (N_12277,N_11773,N_11743);
and U12278 (N_12278,N_11794,N_11369);
and U12279 (N_12279,N_11971,N_11715);
or U12280 (N_12280,N_11634,N_11385);
nor U12281 (N_12281,N_11254,N_11750);
and U12282 (N_12282,N_11895,N_11428);
or U12283 (N_12283,N_11596,N_11942);
nand U12284 (N_12284,N_11540,N_11732);
nor U12285 (N_12285,N_11300,N_11280);
nor U12286 (N_12286,N_11888,N_11279);
nand U12287 (N_12287,N_11521,N_11390);
or U12288 (N_12288,N_11777,N_11735);
nor U12289 (N_12289,N_11310,N_11724);
nand U12290 (N_12290,N_11776,N_11393);
or U12291 (N_12291,N_11543,N_11590);
nand U12292 (N_12292,N_11266,N_11358);
nor U12293 (N_12293,N_11456,N_11698);
xnor U12294 (N_12294,N_11355,N_11930);
or U12295 (N_12295,N_11707,N_11763);
and U12296 (N_12296,N_11502,N_11643);
or U12297 (N_12297,N_11396,N_11277);
or U12298 (N_12298,N_11294,N_11345);
nand U12299 (N_12299,N_11901,N_11871);
and U12300 (N_12300,N_11340,N_11404);
and U12301 (N_12301,N_11411,N_11438);
nand U12302 (N_12302,N_11359,N_11570);
or U12303 (N_12303,N_11258,N_11487);
nor U12304 (N_12304,N_11911,N_11557);
or U12305 (N_12305,N_11879,N_11760);
and U12306 (N_12306,N_11738,N_11944);
and U12307 (N_12307,N_11644,N_11434);
nand U12308 (N_12308,N_11612,N_11887);
nor U12309 (N_12309,N_11293,N_11439);
nor U12310 (N_12310,N_11883,N_11463);
or U12311 (N_12311,N_11729,N_11789);
and U12312 (N_12312,N_11305,N_11379);
or U12313 (N_12313,N_11842,N_11619);
and U12314 (N_12314,N_11479,N_11257);
nor U12315 (N_12315,N_11362,N_11755);
or U12316 (N_12316,N_11583,N_11959);
and U12317 (N_12317,N_11909,N_11745);
or U12318 (N_12318,N_11422,N_11892);
and U12319 (N_12319,N_11907,N_11717);
and U12320 (N_12320,N_11588,N_11333);
xor U12321 (N_12321,N_11437,N_11927);
and U12322 (N_12322,N_11368,N_11949);
and U12323 (N_12323,N_11489,N_11956);
nand U12324 (N_12324,N_11325,N_11933);
and U12325 (N_12325,N_11726,N_11461);
or U12326 (N_12326,N_11925,N_11356);
or U12327 (N_12327,N_11848,N_11312);
nor U12328 (N_12328,N_11864,N_11906);
nor U12329 (N_12329,N_11684,N_11641);
or U12330 (N_12330,N_11558,N_11904);
nor U12331 (N_12331,N_11593,N_11560);
nand U12332 (N_12332,N_11440,N_11374);
and U12333 (N_12333,N_11629,N_11605);
nor U12334 (N_12334,N_11263,N_11826);
or U12335 (N_12335,N_11946,N_11400);
or U12336 (N_12336,N_11443,N_11579);
nor U12337 (N_12337,N_11757,N_11952);
nor U12338 (N_12338,N_11980,N_11256);
or U12339 (N_12339,N_11874,N_11546);
nand U12340 (N_12340,N_11451,N_11307);
nor U12341 (N_12341,N_11919,N_11820);
or U12342 (N_12342,N_11657,N_11654);
nor U12343 (N_12343,N_11423,N_11828);
or U12344 (N_12344,N_11514,N_11894);
nor U12345 (N_12345,N_11308,N_11261);
nor U12346 (N_12346,N_11779,N_11734);
nor U12347 (N_12347,N_11524,N_11978);
nor U12348 (N_12348,N_11731,N_11889);
nand U12349 (N_12349,N_11344,N_11265);
or U12350 (N_12350,N_11408,N_11998);
nand U12351 (N_12351,N_11267,N_11336);
and U12352 (N_12352,N_11885,N_11782);
nand U12353 (N_12353,N_11625,N_11457);
and U12354 (N_12354,N_11320,N_11360);
nor U12355 (N_12355,N_11899,N_11639);
nor U12356 (N_12356,N_11584,N_11251);
nor U12357 (N_12357,N_11380,N_11860);
nor U12358 (N_12358,N_11741,N_11329);
nor U12359 (N_12359,N_11647,N_11954);
nor U12360 (N_12360,N_11516,N_11375);
or U12361 (N_12361,N_11302,N_11884);
or U12362 (N_12362,N_11766,N_11882);
nand U12363 (N_12363,N_11966,N_11987);
nand U12364 (N_12364,N_11861,N_11672);
or U12365 (N_12365,N_11668,N_11342);
nand U12366 (N_12366,N_11470,N_11545);
nand U12367 (N_12367,N_11793,N_11696);
or U12368 (N_12368,N_11962,N_11458);
nor U12369 (N_12369,N_11937,N_11497);
nand U12370 (N_12370,N_11392,N_11372);
nor U12371 (N_12371,N_11532,N_11569);
nand U12372 (N_12372,N_11538,N_11272);
nor U12373 (N_12373,N_11275,N_11953);
nand U12374 (N_12374,N_11517,N_11519);
nor U12375 (N_12375,N_11860,N_11532);
and U12376 (N_12376,N_11252,N_11509);
and U12377 (N_12377,N_11683,N_11922);
and U12378 (N_12378,N_11454,N_11998);
or U12379 (N_12379,N_11962,N_11688);
and U12380 (N_12380,N_11955,N_11491);
or U12381 (N_12381,N_11314,N_11767);
nor U12382 (N_12382,N_11376,N_11390);
nand U12383 (N_12383,N_11339,N_11692);
or U12384 (N_12384,N_11789,N_11619);
nand U12385 (N_12385,N_11388,N_11574);
or U12386 (N_12386,N_11846,N_11716);
and U12387 (N_12387,N_11576,N_11643);
or U12388 (N_12388,N_11481,N_11279);
nor U12389 (N_12389,N_11938,N_11524);
or U12390 (N_12390,N_11712,N_11695);
nand U12391 (N_12391,N_11737,N_11535);
nand U12392 (N_12392,N_11673,N_11822);
nor U12393 (N_12393,N_11810,N_11620);
nand U12394 (N_12394,N_11486,N_11637);
nor U12395 (N_12395,N_11822,N_11549);
nor U12396 (N_12396,N_11771,N_11956);
nor U12397 (N_12397,N_11497,N_11768);
or U12398 (N_12398,N_11995,N_11936);
nor U12399 (N_12399,N_11733,N_11534);
nor U12400 (N_12400,N_11540,N_11762);
or U12401 (N_12401,N_11932,N_11519);
nand U12402 (N_12402,N_11994,N_11977);
and U12403 (N_12403,N_11366,N_11494);
or U12404 (N_12404,N_11685,N_11308);
nand U12405 (N_12405,N_11426,N_11690);
nor U12406 (N_12406,N_11412,N_11774);
nor U12407 (N_12407,N_11428,N_11292);
nand U12408 (N_12408,N_11891,N_11324);
or U12409 (N_12409,N_11575,N_11454);
nand U12410 (N_12410,N_11848,N_11774);
or U12411 (N_12411,N_11353,N_11960);
nor U12412 (N_12412,N_11609,N_11597);
nor U12413 (N_12413,N_11795,N_11842);
nand U12414 (N_12414,N_11780,N_11753);
and U12415 (N_12415,N_11501,N_11389);
and U12416 (N_12416,N_11541,N_11456);
nor U12417 (N_12417,N_11325,N_11832);
nand U12418 (N_12418,N_11598,N_11296);
or U12419 (N_12419,N_11769,N_11960);
and U12420 (N_12420,N_11349,N_11448);
or U12421 (N_12421,N_11668,N_11705);
nor U12422 (N_12422,N_11562,N_11994);
nor U12423 (N_12423,N_11307,N_11281);
nand U12424 (N_12424,N_11959,N_11988);
nand U12425 (N_12425,N_11306,N_11689);
nor U12426 (N_12426,N_11910,N_11657);
nor U12427 (N_12427,N_11674,N_11596);
nor U12428 (N_12428,N_11257,N_11557);
nor U12429 (N_12429,N_11597,N_11447);
or U12430 (N_12430,N_11256,N_11309);
nand U12431 (N_12431,N_11412,N_11512);
or U12432 (N_12432,N_11902,N_11868);
nand U12433 (N_12433,N_11517,N_11281);
and U12434 (N_12434,N_11335,N_11475);
or U12435 (N_12435,N_11961,N_11399);
nor U12436 (N_12436,N_11622,N_11957);
nor U12437 (N_12437,N_11447,N_11719);
and U12438 (N_12438,N_11650,N_11446);
and U12439 (N_12439,N_11494,N_11891);
nand U12440 (N_12440,N_11785,N_11891);
nor U12441 (N_12441,N_11819,N_11413);
and U12442 (N_12442,N_11261,N_11924);
nand U12443 (N_12443,N_11404,N_11438);
and U12444 (N_12444,N_11897,N_11601);
and U12445 (N_12445,N_11750,N_11618);
or U12446 (N_12446,N_11968,N_11712);
or U12447 (N_12447,N_11425,N_11836);
and U12448 (N_12448,N_11519,N_11344);
or U12449 (N_12449,N_11338,N_11890);
or U12450 (N_12450,N_11458,N_11341);
nor U12451 (N_12451,N_11469,N_11479);
or U12452 (N_12452,N_11276,N_11420);
or U12453 (N_12453,N_11690,N_11381);
and U12454 (N_12454,N_11865,N_11794);
nand U12455 (N_12455,N_11661,N_11934);
nor U12456 (N_12456,N_11836,N_11612);
nor U12457 (N_12457,N_11643,N_11681);
xor U12458 (N_12458,N_11614,N_11429);
or U12459 (N_12459,N_11833,N_11836);
or U12460 (N_12460,N_11952,N_11726);
or U12461 (N_12461,N_11930,N_11933);
and U12462 (N_12462,N_11634,N_11844);
or U12463 (N_12463,N_11513,N_11854);
and U12464 (N_12464,N_11359,N_11716);
or U12465 (N_12465,N_11659,N_11571);
nand U12466 (N_12466,N_11931,N_11302);
or U12467 (N_12467,N_11507,N_11471);
or U12468 (N_12468,N_11352,N_11489);
nand U12469 (N_12469,N_11652,N_11464);
nor U12470 (N_12470,N_11455,N_11451);
and U12471 (N_12471,N_11857,N_11281);
or U12472 (N_12472,N_11625,N_11979);
nand U12473 (N_12473,N_11934,N_11902);
nor U12474 (N_12474,N_11826,N_11918);
and U12475 (N_12475,N_11812,N_11985);
nand U12476 (N_12476,N_11791,N_11382);
nor U12477 (N_12477,N_11731,N_11840);
nor U12478 (N_12478,N_11988,N_11722);
nand U12479 (N_12479,N_11600,N_11534);
nand U12480 (N_12480,N_11386,N_11741);
nand U12481 (N_12481,N_11351,N_11516);
nor U12482 (N_12482,N_11815,N_11953);
and U12483 (N_12483,N_11842,N_11920);
or U12484 (N_12484,N_11471,N_11728);
nor U12485 (N_12485,N_11623,N_11306);
and U12486 (N_12486,N_11519,N_11356);
or U12487 (N_12487,N_11507,N_11384);
nand U12488 (N_12488,N_11861,N_11961);
or U12489 (N_12489,N_11835,N_11541);
or U12490 (N_12490,N_11389,N_11921);
nand U12491 (N_12491,N_11495,N_11937);
nand U12492 (N_12492,N_11327,N_11258);
nor U12493 (N_12493,N_11296,N_11566);
or U12494 (N_12494,N_11731,N_11375);
nor U12495 (N_12495,N_11505,N_11768);
or U12496 (N_12496,N_11931,N_11843);
or U12497 (N_12497,N_11792,N_11755);
or U12498 (N_12498,N_11757,N_11550);
or U12499 (N_12499,N_11697,N_11900);
or U12500 (N_12500,N_11764,N_11436);
nor U12501 (N_12501,N_11716,N_11722);
nor U12502 (N_12502,N_11532,N_11515);
and U12503 (N_12503,N_11320,N_11750);
nand U12504 (N_12504,N_11987,N_11795);
or U12505 (N_12505,N_11514,N_11538);
nand U12506 (N_12506,N_11396,N_11356);
and U12507 (N_12507,N_11374,N_11416);
and U12508 (N_12508,N_11472,N_11717);
or U12509 (N_12509,N_11889,N_11906);
nand U12510 (N_12510,N_11567,N_11399);
or U12511 (N_12511,N_11802,N_11437);
nor U12512 (N_12512,N_11973,N_11829);
nor U12513 (N_12513,N_11760,N_11969);
nor U12514 (N_12514,N_11776,N_11440);
and U12515 (N_12515,N_11338,N_11551);
and U12516 (N_12516,N_11585,N_11877);
nor U12517 (N_12517,N_11649,N_11864);
nand U12518 (N_12518,N_11336,N_11415);
and U12519 (N_12519,N_11826,N_11665);
and U12520 (N_12520,N_11322,N_11755);
or U12521 (N_12521,N_11307,N_11508);
and U12522 (N_12522,N_11329,N_11848);
nand U12523 (N_12523,N_11373,N_11944);
and U12524 (N_12524,N_11762,N_11980);
nand U12525 (N_12525,N_11690,N_11639);
nand U12526 (N_12526,N_11713,N_11584);
nor U12527 (N_12527,N_11549,N_11984);
xnor U12528 (N_12528,N_11583,N_11321);
or U12529 (N_12529,N_11574,N_11506);
nand U12530 (N_12530,N_11858,N_11528);
nand U12531 (N_12531,N_11558,N_11261);
or U12532 (N_12532,N_11993,N_11331);
and U12533 (N_12533,N_11621,N_11635);
or U12534 (N_12534,N_11638,N_11823);
or U12535 (N_12535,N_11591,N_11620);
and U12536 (N_12536,N_11550,N_11795);
nand U12537 (N_12537,N_11451,N_11967);
and U12538 (N_12538,N_11298,N_11601);
or U12539 (N_12539,N_11348,N_11735);
and U12540 (N_12540,N_11372,N_11874);
or U12541 (N_12541,N_11384,N_11582);
nor U12542 (N_12542,N_11286,N_11697);
and U12543 (N_12543,N_11441,N_11512);
nor U12544 (N_12544,N_11768,N_11700);
nor U12545 (N_12545,N_11771,N_11520);
or U12546 (N_12546,N_11448,N_11614);
and U12547 (N_12547,N_11546,N_11317);
nor U12548 (N_12548,N_11362,N_11531);
nand U12549 (N_12549,N_11772,N_11813);
and U12550 (N_12550,N_11947,N_11981);
nand U12551 (N_12551,N_11855,N_11496);
or U12552 (N_12552,N_11846,N_11581);
or U12553 (N_12553,N_11467,N_11980);
nand U12554 (N_12554,N_11596,N_11286);
or U12555 (N_12555,N_11625,N_11255);
and U12556 (N_12556,N_11852,N_11473);
and U12557 (N_12557,N_11516,N_11532);
or U12558 (N_12558,N_11571,N_11497);
nor U12559 (N_12559,N_11559,N_11869);
and U12560 (N_12560,N_11971,N_11381);
or U12561 (N_12561,N_11463,N_11529);
and U12562 (N_12562,N_11294,N_11259);
or U12563 (N_12563,N_11935,N_11668);
nor U12564 (N_12564,N_11736,N_11530);
nand U12565 (N_12565,N_11363,N_11632);
nand U12566 (N_12566,N_11400,N_11598);
and U12567 (N_12567,N_11414,N_11618);
nor U12568 (N_12568,N_11435,N_11886);
or U12569 (N_12569,N_11362,N_11691);
nor U12570 (N_12570,N_11415,N_11723);
nand U12571 (N_12571,N_11918,N_11888);
nor U12572 (N_12572,N_11563,N_11356);
or U12573 (N_12573,N_11527,N_11342);
or U12574 (N_12574,N_11961,N_11688);
nand U12575 (N_12575,N_11312,N_11951);
nor U12576 (N_12576,N_11705,N_11616);
nand U12577 (N_12577,N_11435,N_11698);
and U12578 (N_12578,N_11537,N_11502);
and U12579 (N_12579,N_11990,N_11978);
nand U12580 (N_12580,N_11935,N_11953);
and U12581 (N_12581,N_11961,N_11550);
or U12582 (N_12582,N_11696,N_11352);
nor U12583 (N_12583,N_11490,N_11789);
or U12584 (N_12584,N_11984,N_11560);
or U12585 (N_12585,N_11686,N_11982);
nand U12586 (N_12586,N_11475,N_11316);
nand U12587 (N_12587,N_11699,N_11954);
xnor U12588 (N_12588,N_11423,N_11482);
nor U12589 (N_12589,N_11955,N_11704);
nor U12590 (N_12590,N_11996,N_11630);
or U12591 (N_12591,N_11866,N_11690);
nand U12592 (N_12592,N_11482,N_11644);
nand U12593 (N_12593,N_11991,N_11880);
nor U12594 (N_12594,N_11821,N_11841);
or U12595 (N_12595,N_11408,N_11551);
nor U12596 (N_12596,N_11437,N_11941);
and U12597 (N_12597,N_11536,N_11893);
nor U12598 (N_12598,N_11762,N_11903);
or U12599 (N_12599,N_11718,N_11426);
or U12600 (N_12600,N_11479,N_11737);
or U12601 (N_12601,N_11752,N_11284);
and U12602 (N_12602,N_11880,N_11945);
or U12603 (N_12603,N_11352,N_11276);
and U12604 (N_12604,N_11488,N_11900);
or U12605 (N_12605,N_11511,N_11853);
nand U12606 (N_12606,N_11350,N_11276);
or U12607 (N_12607,N_11907,N_11459);
nand U12608 (N_12608,N_11414,N_11997);
and U12609 (N_12609,N_11992,N_11488);
nor U12610 (N_12610,N_11450,N_11545);
and U12611 (N_12611,N_11932,N_11272);
and U12612 (N_12612,N_11803,N_11360);
or U12613 (N_12613,N_11689,N_11519);
and U12614 (N_12614,N_11480,N_11510);
or U12615 (N_12615,N_11391,N_11895);
and U12616 (N_12616,N_11764,N_11331);
nor U12617 (N_12617,N_11368,N_11749);
nor U12618 (N_12618,N_11751,N_11313);
nand U12619 (N_12619,N_11427,N_11713);
nor U12620 (N_12620,N_11390,N_11974);
or U12621 (N_12621,N_11956,N_11661);
or U12622 (N_12622,N_11480,N_11495);
or U12623 (N_12623,N_11870,N_11851);
or U12624 (N_12624,N_11479,N_11795);
xnor U12625 (N_12625,N_11983,N_11528);
nand U12626 (N_12626,N_11936,N_11356);
nand U12627 (N_12627,N_11600,N_11709);
and U12628 (N_12628,N_11290,N_11556);
nand U12629 (N_12629,N_11842,N_11475);
nor U12630 (N_12630,N_11640,N_11387);
nand U12631 (N_12631,N_11908,N_11917);
or U12632 (N_12632,N_11365,N_11339);
and U12633 (N_12633,N_11855,N_11407);
nand U12634 (N_12634,N_11808,N_11506);
nor U12635 (N_12635,N_11631,N_11698);
nand U12636 (N_12636,N_11471,N_11523);
nand U12637 (N_12637,N_11635,N_11594);
nor U12638 (N_12638,N_11887,N_11663);
nor U12639 (N_12639,N_11818,N_11648);
nor U12640 (N_12640,N_11571,N_11251);
and U12641 (N_12641,N_11709,N_11469);
or U12642 (N_12642,N_11954,N_11425);
nand U12643 (N_12643,N_11887,N_11549);
and U12644 (N_12644,N_11770,N_11609);
nor U12645 (N_12645,N_11796,N_11303);
nand U12646 (N_12646,N_11546,N_11736);
or U12647 (N_12647,N_11838,N_11516);
nor U12648 (N_12648,N_11271,N_11867);
nand U12649 (N_12649,N_11428,N_11443);
nand U12650 (N_12650,N_11986,N_11305);
and U12651 (N_12651,N_11946,N_11862);
nor U12652 (N_12652,N_11797,N_11620);
nand U12653 (N_12653,N_11638,N_11439);
xor U12654 (N_12654,N_11579,N_11629);
nor U12655 (N_12655,N_11488,N_11494);
nor U12656 (N_12656,N_11435,N_11733);
nor U12657 (N_12657,N_11806,N_11759);
nand U12658 (N_12658,N_11298,N_11342);
and U12659 (N_12659,N_11494,N_11676);
nor U12660 (N_12660,N_11853,N_11947);
or U12661 (N_12661,N_11396,N_11599);
nand U12662 (N_12662,N_11541,N_11716);
nand U12663 (N_12663,N_11552,N_11923);
and U12664 (N_12664,N_11392,N_11557);
nand U12665 (N_12665,N_11417,N_11866);
nand U12666 (N_12666,N_11569,N_11993);
and U12667 (N_12667,N_11895,N_11858);
and U12668 (N_12668,N_11649,N_11415);
and U12669 (N_12669,N_11948,N_11505);
and U12670 (N_12670,N_11440,N_11903);
xor U12671 (N_12671,N_11288,N_11410);
nor U12672 (N_12672,N_11509,N_11314);
and U12673 (N_12673,N_11850,N_11595);
nand U12674 (N_12674,N_11324,N_11796);
nor U12675 (N_12675,N_11399,N_11305);
or U12676 (N_12676,N_11374,N_11896);
or U12677 (N_12677,N_11741,N_11697);
nor U12678 (N_12678,N_11349,N_11830);
and U12679 (N_12679,N_11300,N_11284);
or U12680 (N_12680,N_11630,N_11334);
or U12681 (N_12681,N_11308,N_11970);
nor U12682 (N_12682,N_11622,N_11627);
or U12683 (N_12683,N_11671,N_11812);
and U12684 (N_12684,N_11394,N_11610);
nor U12685 (N_12685,N_11391,N_11746);
nand U12686 (N_12686,N_11822,N_11814);
or U12687 (N_12687,N_11558,N_11889);
nor U12688 (N_12688,N_11274,N_11766);
nor U12689 (N_12689,N_11648,N_11251);
or U12690 (N_12690,N_11395,N_11792);
or U12691 (N_12691,N_11673,N_11317);
or U12692 (N_12692,N_11730,N_11969);
or U12693 (N_12693,N_11297,N_11550);
nand U12694 (N_12694,N_11497,N_11801);
and U12695 (N_12695,N_11261,N_11483);
nand U12696 (N_12696,N_11660,N_11930);
nand U12697 (N_12697,N_11655,N_11307);
nor U12698 (N_12698,N_11838,N_11471);
or U12699 (N_12699,N_11913,N_11699);
nor U12700 (N_12700,N_11353,N_11405);
nand U12701 (N_12701,N_11750,N_11864);
nor U12702 (N_12702,N_11993,N_11728);
nor U12703 (N_12703,N_11995,N_11683);
nand U12704 (N_12704,N_11819,N_11855);
nand U12705 (N_12705,N_11936,N_11709);
nor U12706 (N_12706,N_11272,N_11747);
nand U12707 (N_12707,N_11357,N_11744);
nand U12708 (N_12708,N_11816,N_11458);
or U12709 (N_12709,N_11298,N_11933);
or U12710 (N_12710,N_11359,N_11870);
nand U12711 (N_12711,N_11856,N_11489);
or U12712 (N_12712,N_11960,N_11392);
nand U12713 (N_12713,N_11710,N_11432);
nand U12714 (N_12714,N_11937,N_11617);
nand U12715 (N_12715,N_11734,N_11765);
nor U12716 (N_12716,N_11578,N_11654);
nand U12717 (N_12717,N_11508,N_11548);
and U12718 (N_12718,N_11590,N_11940);
and U12719 (N_12719,N_11473,N_11349);
or U12720 (N_12720,N_11587,N_11419);
nand U12721 (N_12721,N_11776,N_11340);
nor U12722 (N_12722,N_11683,N_11462);
nand U12723 (N_12723,N_11428,N_11564);
nand U12724 (N_12724,N_11898,N_11308);
or U12725 (N_12725,N_11889,N_11849);
nor U12726 (N_12726,N_11909,N_11471);
or U12727 (N_12727,N_11407,N_11682);
nand U12728 (N_12728,N_11456,N_11500);
and U12729 (N_12729,N_11827,N_11698);
and U12730 (N_12730,N_11634,N_11474);
and U12731 (N_12731,N_11468,N_11854);
and U12732 (N_12732,N_11811,N_11927);
and U12733 (N_12733,N_11844,N_11340);
or U12734 (N_12734,N_11684,N_11925);
and U12735 (N_12735,N_11252,N_11575);
nand U12736 (N_12736,N_11742,N_11706);
and U12737 (N_12737,N_11506,N_11322);
nor U12738 (N_12738,N_11952,N_11813);
nor U12739 (N_12739,N_11382,N_11704);
and U12740 (N_12740,N_11884,N_11904);
and U12741 (N_12741,N_11325,N_11825);
or U12742 (N_12742,N_11388,N_11553);
and U12743 (N_12743,N_11947,N_11698);
or U12744 (N_12744,N_11460,N_11255);
or U12745 (N_12745,N_11780,N_11757);
and U12746 (N_12746,N_11496,N_11666);
nand U12747 (N_12747,N_11898,N_11679);
or U12748 (N_12748,N_11537,N_11404);
or U12749 (N_12749,N_11973,N_11600);
and U12750 (N_12750,N_12057,N_12056);
nor U12751 (N_12751,N_12353,N_12654);
nand U12752 (N_12752,N_12539,N_12704);
or U12753 (N_12753,N_12435,N_12323);
nor U12754 (N_12754,N_12581,N_12660);
or U12755 (N_12755,N_12598,N_12216);
and U12756 (N_12756,N_12518,N_12081);
nor U12757 (N_12757,N_12426,N_12271);
or U12758 (N_12758,N_12662,N_12441);
nand U12759 (N_12759,N_12264,N_12146);
or U12760 (N_12760,N_12329,N_12445);
nor U12761 (N_12761,N_12507,N_12675);
nand U12762 (N_12762,N_12156,N_12100);
nand U12763 (N_12763,N_12212,N_12269);
nor U12764 (N_12764,N_12711,N_12177);
or U12765 (N_12765,N_12709,N_12721);
nand U12766 (N_12766,N_12682,N_12548);
or U12767 (N_12767,N_12279,N_12288);
nand U12768 (N_12768,N_12553,N_12127);
nand U12769 (N_12769,N_12311,N_12701);
nand U12770 (N_12770,N_12023,N_12229);
and U12771 (N_12771,N_12604,N_12684);
or U12772 (N_12772,N_12064,N_12738);
nor U12773 (N_12773,N_12298,N_12187);
nor U12774 (N_12774,N_12728,N_12535);
or U12775 (N_12775,N_12195,N_12729);
nor U12776 (N_12776,N_12228,N_12392);
and U12777 (N_12777,N_12226,N_12166);
or U12778 (N_12778,N_12063,N_12199);
or U12779 (N_12779,N_12310,N_12230);
or U12780 (N_12780,N_12054,N_12115);
nand U12781 (N_12781,N_12494,N_12748);
nor U12782 (N_12782,N_12651,N_12039);
or U12783 (N_12783,N_12284,N_12712);
and U12784 (N_12784,N_12138,N_12066);
nand U12785 (N_12785,N_12597,N_12048);
and U12786 (N_12786,N_12674,N_12415);
or U12787 (N_12787,N_12324,N_12136);
nor U12788 (N_12788,N_12050,N_12382);
and U12789 (N_12789,N_12217,N_12591);
or U12790 (N_12790,N_12019,N_12293);
and U12791 (N_12791,N_12302,N_12013);
or U12792 (N_12792,N_12473,N_12128);
and U12793 (N_12793,N_12008,N_12648);
or U12794 (N_12794,N_12133,N_12386);
and U12795 (N_12795,N_12582,N_12289);
and U12796 (N_12796,N_12710,N_12594);
nand U12797 (N_12797,N_12234,N_12544);
or U12798 (N_12798,N_12266,N_12458);
and U12799 (N_12799,N_12678,N_12257);
and U12800 (N_12800,N_12732,N_12120);
or U12801 (N_12801,N_12315,N_12419);
nand U12802 (N_12802,N_12049,N_12639);
and U12803 (N_12803,N_12222,N_12479);
nor U12804 (N_12804,N_12537,N_12683);
or U12805 (N_12805,N_12698,N_12555);
nor U12806 (N_12806,N_12188,N_12287);
and U12807 (N_12807,N_12189,N_12538);
or U12808 (N_12808,N_12291,N_12554);
nor U12809 (N_12809,N_12181,N_12546);
nand U12810 (N_12810,N_12277,N_12655);
nand U12811 (N_12811,N_12616,N_12540);
and U12812 (N_12812,N_12275,N_12454);
and U12813 (N_12813,N_12080,N_12154);
nand U12814 (N_12814,N_12645,N_12169);
or U12815 (N_12815,N_12613,N_12573);
nand U12816 (N_12816,N_12493,N_12103);
and U12817 (N_12817,N_12032,N_12240);
and U12818 (N_12818,N_12101,N_12305);
nand U12819 (N_12819,N_12432,N_12263);
nor U12820 (N_12820,N_12631,N_12237);
nor U12821 (N_12821,N_12326,N_12153);
xor U12822 (N_12822,N_12061,N_12468);
nor U12823 (N_12823,N_12492,N_12213);
nor U12824 (N_12824,N_12708,N_12089);
and U12825 (N_12825,N_12145,N_12715);
nor U12826 (N_12826,N_12515,N_12241);
and U12827 (N_12827,N_12502,N_12418);
and U12828 (N_12828,N_12440,N_12235);
nor U12829 (N_12829,N_12409,N_12065);
and U12830 (N_12830,N_12472,N_12427);
and U12831 (N_12831,N_12131,N_12641);
nor U12832 (N_12832,N_12163,N_12112);
nor U12833 (N_12833,N_12547,N_12095);
nand U12834 (N_12834,N_12281,N_12086);
and U12835 (N_12835,N_12031,N_12692);
or U12836 (N_12836,N_12190,N_12303);
xnor U12837 (N_12837,N_12077,N_12193);
or U12838 (N_12838,N_12149,N_12429);
or U12839 (N_12839,N_12612,N_12344);
or U12840 (N_12840,N_12376,N_12511);
and U12841 (N_12841,N_12044,N_12088);
or U12842 (N_12842,N_12076,N_12703);
nor U12843 (N_12843,N_12624,N_12245);
and U12844 (N_12844,N_12723,N_12041);
and U12845 (N_12845,N_12521,N_12233);
nor U12846 (N_12846,N_12564,N_12680);
or U12847 (N_12847,N_12135,N_12716);
nand U12848 (N_12848,N_12151,N_12215);
nand U12849 (N_12849,N_12238,N_12173);
and U12850 (N_12850,N_12697,N_12105);
or U12851 (N_12851,N_12366,N_12236);
and U12852 (N_12852,N_12431,N_12200);
and U12853 (N_12853,N_12357,N_12733);
and U12854 (N_12854,N_12300,N_12693);
and U12855 (N_12855,N_12242,N_12513);
nor U12856 (N_12856,N_12390,N_12260);
or U12857 (N_12857,N_12621,N_12691);
and U12858 (N_12858,N_12576,N_12068);
nand U12859 (N_12859,N_12037,N_12003);
or U12860 (N_12860,N_12070,N_12223);
and U12861 (N_12861,N_12626,N_12208);
and U12862 (N_12862,N_12335,N_12198);
nand U12863 (N_12863,N_12667,N_12273);
nor U12864 (N_12864,N_12542,N_12417);
and U12865 (N_12865,N_12219,N_12380);
and U12866 (N_12866,N_12336,N_12423);
or U12867 (N_12867,N_12010,N_12410);
or U12868 (N_12868,N_12157,N_12451);
nor U12869 (N_12869,N_12206,N_12178);
and U12870 (N_12870,N_12456,N_12465);
nor U12871 (N_12871,N_12455,N_12497);
nor U12872 (N_12872,N_12561,N_12253);
nor U12873 (N_12873,N_12268,N_12498);
and U12874 (N_12874,N_12543,N_12259);
or U12875 (N_12875,N_12171,N_12139);
nand U12876 (N_12876,N_12608,N_12227);
nor U12877 (N_12877,N_12001,N_12144);
and U12878 (N_12878,N_12038,N_12285);
nor U12879 (N_12879,N_12255,N_12421);
and U12880 (N_12880,N_12349,N_12098);
nor U12881 (N_12881,N_12736,N_12580);
and U12882 (N_12882,N_12730,N_12352);
and U12883 (N_12883,N_12307,N_12125);
nand U12884 (N_12884,N_12114,N_12487);
and U12885 (N_12885,N_12405,N_12205);
nand U12886 (N_12886,N_12747,N_12588);
or U12887 (N_12887,N_12265,N_12474);
xor U12888 (N_12888,N_12749,N_12517);
xor U12889 (N_12889,N_12152,N_12119);
and U12890 (N_12890,N_12278,N_12345);
and U12891 (N_12891,N_12183,N_12677);
nand U12892 (N_12892,N_12516,N_12143);
nor U12893 (N_12893,N_12276,N_12447);
nor U12894 (N_12894,N_12433,N_12182);
and U12895 (N_12895,N_12396,N_12571);
nor U12896 (N_12896,N_12179,N_12665);
nand U12897 (N_12897,N_12055,N_12280);
nand U12898 (N_12898,N_12681,N_12658);
nand U12899 (N_12899,N_12282,N_12015);
nand U12900 (N_12900,N_12043,N_12130);
nor U12901 (N_12901,N_12122,N_12123);
nand U12902 (N_12902,N_12734,N_12485);
and U12903 (N_12903,N_12406,N_12342);
and U12904 (N_12904,N_12559,N_12186);
nor U12905 (N_12905,N_12514,N_12332);
or U12906 (N_12906,N_12155,N_12393);
or U12907 (N_12907,N_12168,N_12231);
or U12908 (N_12908,N_12113,N_12262);
or U12909 (N_12909,N_12073,N_12094);
or U12910 (N_12910,N_12358,N_12207);
nand U12911 (N_12911,N_12110,N_12254);
nand U12912 (N_12912,N_12522,N_12132);
nor U12913 (N_12913,N_12078,N_12642);
and U12914 (N_12914,N_12140,N_12197);
or U12915 (N_12915,N_12337,N_12046);
and U12916 (N_12916,N_12014,N_12314);
and U12917 (N_12917,N_12165,N_12368);
nor U12918 (N_12918,N_12702,N_12209);
nand U12919 (N_12919,N_12283,N_12439);
and U12920 (N_12920,N_12534,N_12121);
nor U12921 (N_12921,N_12673,N_12731);
nor U12922 (N_12922,N_12270,N_12087);
nor U12923 (N_12923,N_12569,N_12586);
and U12924 (N_12924,N_12656,N_12695);
and U12925 (N_12925,N_12220,N_12661);
nand U12926 (N_12926,N_12011,N_12536);
nor U12927 (N_12927,N_12478,N_12629);
nand U12928 (N_12928,N_12218,N_12028);
nor U12929 (N_12929,N_12638,N_12587);
or U12930 (N_12930,N_12148,N_12483);
and U12931 (N_12931,N_12664,N_12556);
nand U12932 (N_12932,N_12117,N_12420);
nor U12933 (N_12933,N_12202,N_12462);
nand U12934 (N_12934,N_12615,N_12707);
and U12935 (N_12935,N_12690,N_12243);
or U12936 (N_12936,N_12557,N_12640);
nor U12937 (N_12937,N_12051,N_12742);
or U12938 (N_12938,N_12083,N_12005);
and U12939 (N_12939,N_12290,N_12109);
nand U12940 (N_12940,N_12325,N_12356);
and U12941 (N_12941,N_12167,N_12312);
and U12942 (N_12942,N_12689,N_12413);
or U12943 (N_12943,N_12510,N_12176);
nand U12944 (N_12944,N_12676,N_12652);
and U12945 (N_12945,N_12446,N_12365);
nor U12946 (N_12946,N_12496,N_12568);
or U12947 (N_12947,N_12036,N_12566);
and U12948 (N_12948,N_12308,N_12351);
nor U12949 (N_12949,N_12603,N_12339);
nand U12950 (N_12950,N_12040,N_12004);
nand U12951 (N_12951,N_12450,N_12074);
and U12952 (N_12952,N_12428,N_12668);
or U12953 (N_12953,N_12622,N_12142);
and U12954 (N_12954,N_12469,N_12482);
or U12955 (N_12955,N_12726,N_12071);
nand U12956 (N_12956,N_12304,N_12623);
xnor U12957 (N_12957,N_12346,N_12718);
and U12958 (N_12958,N_12210,N_12360);
xor U12959 (N_12959,N_12286,N_12574);
and U12960 (N_12960,N_12274,N_12299);
nor U12961 (N_12961,N_12481,N_12745);
nand U12962 (N_12962,N_12505,N_12267);
and U12963 (N_12963,N_12625,N_12714);
nand U12964 (N_12964,N_12449,N_12118);
nand U12965 (N_12965,N_12079,N_12509);
or U12966 (N_12966,N_12434,N_12694);
and U12967 (N_12967,N_12328,N_12545);
and U12968 (N_12968,N_12388,N_12414);
and U12969 (N_12969,N_12012,N_12592);
and U12970 (N_12970,N_12599,N_12221);
nor U12971 (N_12971,N_12137,N_12725);
and U12972 (N_12972,N_12425,N_12609);
nor U12973 (N_12973,N_12422,N_12744);
nor U12974 (N_12974,N_12175,N_12649);
nor U12975 (N_12975,N_12343,N_12045);
nand U12976 (N_12976,N_12700,N_12593);
and U12977 (N_12977,N_12464,N_12102);
nor U12978 (N_12978,N_12348,N_12585);
nor U12979 (N_12979,N_12141,N_12035);
nor U12980 (N_12980,N_12552,N_12696);
or U12981 (N_12981,N_12111,N_12192);
nor U12982 (N_12982,N_12589,N_12448);
nand U12983 (N_12983,N_12584,N_12203);
nand U12984 (N_12984,N_12490,N_12488);
nand U12985 (N_12985,N_12318,N_12363);
or U12986 (N_12986,N_12252,N_12532);
nand U12987 (N_12987,N_12605,N_12634);
nor U12988 (N_12988,N_12172,N_12508);
or U12989 (N_12989,N_12397,N_12575);
and U12990 (N_12990,N_12258,N_12006);
or U12991 (N_12991,N_12579,N_12412);
nor U12992 (N_12992,N_12249,N_12021);
nor U12993 (N_12993,N_12350,N_12411);
nand U12994 (N_12994,N_12741,N_12630);
nor U12995 (N_12995,N_12387,N_12327);
nand U12996 (N_12996,N_12129,N_12367);
and U12997 (N_12997,N_12672,N_12407);
or U12998 (N_12998,N_12436,N_12457);
nor U12999 (N_12999,N_12317,N_12164);
or U13000 (N_13000,N_12191,N_12256);
nor U13001 (N_13001,N_12408,N_12637);
nor U13002 (N_13002,N_12194,N_12463);
nand U13003 (N_13003,N_12669,N_12644);
or U13004 (N_13004,N_12529,N_12364);
or U13005 (N_13005,N_12523,N_12400);
nor U13006 (N_13006,N_12602,N_12359);
and U13007 (N_13007,N_12085,N_12403);
nor U13008 (N_13008,N_12058,N_12116);
or U13009 (N_13009,N_12467,N_12685);
and U13010 (N_13010,N_12550,N_12016);
nor U13011 (N_13011,N_12477,N_12453);
nor U13012 (N_13012,N_12309,N_12562);
or U13013 (N_13013,N_12106,N_12746);
and U13014 (N_13014,N_12371,N_12577);
and U13015 (N_13015,N_12666,N_12082);
or U13016 (N_13016,N_12059,N_12520);
nand U13017 (N_13017,N_12124,N_12062);
nor U13018 (N_13018,N_12180,N_12601);
or U13019 (N_13019,N_12161,N_12444);
nor U13020 (N_13020,N_12531,N_12296);
and U13021 (N_13021,N_12635,N_12533);
nand U13022 (N_13022,N_12373,N_12354);
nand U13023 (N_13023,N_12201,N_12247);
nand U13024 (N_13024,N_12033,N_12204);
or U13025 (N_13025,N_12657,N_12370);
and U13026 (N_13026,N_12459,N_12026);
nand U13027 (N_13027,N_12381,N_12294);
nor U13028 (N_13028,N_12007,N_12024);
and U13029 (N_13029,N_12160,N_12184);
nor U13030 (N_13030,N_12740,N_12093);
xor U13031 (N_13031,N_12670,N_12743);
and U13032 (N_13032,N_12042,N_12334);
nor U13033 (N_13033,N_12355,N_12052);
nand U13034 (N_13034,N_12362,N_12452);
nor U13035 (N_13035,N_12025,N_12313);
and U13036 (N_13036,N_12404,N_12600);
nor U13037 (N_13037,N_12570,N_12541);
or U13038 (N_13038,N_12687,N_12075);
nand U13039 (N_13039,N_12484,N_12567);
nand U13040 (N_13040,N_12688,N_12306);
and U13041 (N_13041,N_12107,N_12643);
nand U13042 (N_13042,N_12398,N_12633);
and U13043 (N_13043,N_12379,N_12526);
or U13044 (N_13044,N_12647,N_12663);
nor U13045 (N_13045,N_12369,N_12385);
nor U13046 (N_13046,N_12147,N_12196);
and U13047 (N_13047,N_12470,N_12372);
nor U13048 (N_13048,N_12512,N_12471);
and U13049 (N_13049,N_12491,N_12319);
or U13050 (N_13050,N_12506,N_12091);
or U13051 (N_13051,N_12020,N_12430);
nor U13052 (N_13052,N_12560,N_12316);
nor U13053 (N_13053,N_12292,N_12174);
and U13054 (N_13054,N_12606,N_12719);
and U13055 (N_13055,N_12248,N_12578);
or U13056 (N_13056,N_12027,N_12361);
and U13057 (N_13057,N_12524,N_12424);
or U13058 (N_13058,N_12558,N_12530);
nand U13059 (N_13059,N_12653,N_12659);
nor U13060 (N_13060,N_12500,N_12097);
nor U13061 (N_13061,N_12295,N_12565);
nand U13062 (N_13062,N_12320,N_12232);
nand U13063 (N_13063,N_12029,N_12126);
nand U13064 (N_13064,N_12519,N_12739);
xnor U13065 (N_13065,N_12727,N_12159);
or U13066 (N_13066,N_12583,N_12475);
and U13067 (N_13067,N_12214,N_12009);
nand U13068 (N_13068,N_12170,N_12341);
or U13069 (N_13069,N_12374,N_12347);
and U13070 (N_13070,N_12053,N_12394);
or U13071 (N_13071,N_12443,N_12720);
nor U13072 (N_13072,N_12620,N_12646);
or U13073 (N_13073,N_12628,N_12722);
or U13074 (N_13074,N_12461,N_12486);
nand U13075 (N_13075,N_12618,N_12416);
nor U13076 (N_13076,N_12504,N_12717);
nand U13077 (N_13077,N_12384,N_12002);
or U13078 (N_13078,N_12096,N_12377);
nor U13079 (N_13079,N_12466,N_12162);
nor U13080 (N_13080,N_12735,N_12596);
or U13081 (N_13081,N_12699,N_12724);
or U13082 (N_13082,N_12383,N_12017);
and U13083 (N_13083,N_12636,N_12158);
nand U13084 (N_13084,N_12251,N_12084);
nor U13085 (N_13085,N_12501,N_12099);
or U13086 (N_13086,N_12000,N_12617);
or U13087 (N_13087,N_12244,N_12090);
nand U13088 (N_13088,N_12590,N_12060);
nor U13089 (N_13089,N_12437,N_12671);
or U13090 (N_13090,N_12442,N_12503);
or U13091 (N_13091,N_12528,N_12402);
nor U13092 (N_13092,N_12340,N_12614);
nand U13093 (N_13093,N_12034,N_12679);
nor U13094 (N_13094,N_12018,N_12104);
nand U13095 (N_13095,N_12333,N_12331);
nand U13096 (N_13096,N_12391,N_12338);
nor U13097 (N_13097,N_12632,N_12389);
nand U13098 (N_13098,N_12401,N_12272);
nand U13099 (N_13099,N_12072,N_12321);
and U13100 (N_13100,N_12525,N_12395);
nor U13101 (N_13101,N_12611,N_12460);
and U13102 (N_13102,N_12022,N_12047);
and U13103 (N_13103,N_12527,N_12480);
and U13104 (N_13104,N_12134,N_12250);
nor U13105 (N_13105,N_12261,N_12499);
nor U13106 (N_13106,N_12030,N_12150);
and U13107 (N_13107,N_12619,N_12322);
nor U13108 (N_13108,N_12476,N_12595);
nand U13109 (N_13109,N_12737,N_12092);
and U13110 (N_13110,N_12495,N_12607);
and U13111 (N_13111,N_12551,N_12297);
nand U13112 (N_13112,N_12185,N_12610);
or U13113 (N_13113,N_12650,N_12489);
or U13114 (N_13114,N_12069,N_12239);
or U13115 (N_13115,N_12627,N_12686);
or U13116 (N_13116,N_12399,N_12301);
and U13117 (N_13117,N_12067,N_12713);
or U13118 (N_13118,N_12330,N_12705);
nand U13119 (N_13119,N_12563,N_12108);
nand U13120 (N_13120,N_12224,N_12211);
nand U13121 (N_13121,N_12246,N_12572);
nand U13122 (N_13122,N_12438,N_12375);
nand U13123 (N_13123,N_12706,N_12225);
nand U13124 (N_13124,N_12549,N_12378);
nand U13125 (N_13125,N_12290,N_12281);
or U13126 (N_13126,N_12161,N_12036);
or U13127 (N_13127,N_12429,N_12079);
or U13128 (N_13128,N_12227,N_12365);
nand U13129 (N_13129,N_12232,N_12686);
or U13130 (N_13130,N_12427,N_12652);
and U13131 (N_13131,N_12707,N_12264);
nor U13132 (N_13132,N_12688,N_12354);
or U13133 (N_13133,N_12209,N_12366);
and U13134 (N_13134,N_12675,N_12352);
and U13135 (N_13135,N_12063,N_12099);
nor U13136 (N_13136,N_12023,N_12389);
and U13137 (N_13137,N_12331,N_12608);
and U13138 (N_13138,N_12718,N_12466);
nor U13139 (N_13139,N_12310,N_12652);
or U13140 (N_13140,N_12690,N_12122);
nor U13141 (N_13141,N_12168,N_12592);
and U13142 (N_13142,N_12317,N_12351);
and U13143 (N_13143,N_12526,N_12142);
or U13144 (N_13144,N_12329,N_12384);
or U13145 (N_13145,N_12435,N_12680);
nand U13146 (N_13146,N_12267,N_12180);
and U13147 (N_13147,N_12629,N_12242);
and U13148 (N_13148,N_12642,N_12726);
and U13149 (N_13149,N_12210,N_12239);
and U13150 (N_13150,N_12346,N_12603);
and U13151 (N_13151,N_12400,N_12297);
nor U13152 (N_13152,N_12175,N_12530);
nor U13153 (N_13153,N_12397,N_12466);
and U13154 (N_13154,N_12049,N_12215);
nand U13155 (N_13155,N_12715,N_12160);
and U13156 (N_13156,N_12625,N_12285);
nor U13157 (N_13157,N_12428,N_12654);
nand U13158 (N_13158,N_12541,N_12274);
nand U13159 (N_13159,N_12410,N_12398);
and U13160 (N_13160,N_12367,N_12141);
and U13161 (N_13161,N_12606,N_12523);
or U13162 (N_13162,N_12478,N_12571);
nand U13163 (N_13163,N_12117,N_12671);
and U13164 (N_13164,N_12294,N_12604);
or U13165 (N_13165,N_12047,N_12610);
nor U13166 (N_13166,N_12619,N_12479);
nor U13167 (N_13167,N_12307,N_12140);
and U13168 (N_13168,N_12601,N_12572);
and U13169 (N_13169,N_12607,N_12564);
and U13170 (N_13170,N_12749,N_12717);
and U13171 (N_13171,N_12234,N_12648);
nor U13172 (N_13172,N_12262,N_12257);
and U13173 (N_13173,N_12370,N_12406);
or U13174 (N_13174,N_12230,N_12514);
nand U13175 (N_13175,N_12243,N_12565);
or U13176 (N_13176,N_12524,N_12080);
and U13177 (N_13177,N_12117,N_12547);
or U13178 (N_13178,N_12087,N_12228);
and U13179 (N_13179,N_12035,N_12175);
nand U13180 (N_13180,N_12455,N_12029);
or U13181 (N_13181,N_12239,N_12223);
and U13182 (N_13182,N_12143,N_12230);
or U13183 (N_13183,N_12244,N_12474);
nand U13184 (N_13184,N_12675,N_12367);
or U13185 (N_13185,N_12356,N_12433);
nor U13186 (N_13186,N_12623,N_12068);
or U13187 (N_13187,N_12709,N_12614);
xor U13188 (N_13188,N_12071,N_12460);
and U13189 (N_13189,N_12053,N_12205);
nor U13190 (N_13190,N_12080,N_12542);
nand U13191 (N_13191,N_12503,N_12440);
or U13192 (N_13192,N_12533,N_12435);
or U13193 (N_13193,N_12286,N_12285);
or U13194 (N_13194,N_12670,N_12032);
nand U13195 (N_13195,N_12207,N_12556);
nor U13196 (N_13196,N_12097,N_12162);
nor U13197 (N_13197,N_12647,N_12110);
and U13198 (N_13198,N_12586,N_12236);
nand U13199 (N_13199,N_12087,N_12597);
or U13200 (N_13200,N_12076,N_12320);
nor U13201 (N_13201,N_12337,N_12048);
nor U13202 (N_13202,N_12577,N_12532);
or U13203 (N_13203,N_12489,N_12030);
nand U13204 (N_13204,N_12403,N_12134);
or U13205 (N_13205,N_12544,N_12365);
nand U13206 (N_13206,N_12191,N_12351);
or U13207 (N_13207,N_12029,N_12050);
and U13208 (N_13208,N_12024,N_12126);
nor U13209 (N_13209,N_12726,N_12180);
nor U13210 (N_13210,N_12223,N_12090);
nand U13211 (N_13211,N_12318,N_12707);
and U13212 (N_13212,N_12319,N_12525);
and U13213 (N_13213,N_12262,N_12226);
nor U13214 (N_13214,N_12086,N_12100);
nand U13215 (N_13215,N_12264,N_12312);
nand U13216 (N_13216,N_12469,N_12260);
nand U13217 (N_13217,N_12084,N_12638);
or U13218 (N_13218,N_12041,N_12101);
and U13219 (N_13219,N_12408,N_12467);
nor U13220 (N_13220,N_12274,N_12509);
nand U13221 (N_13221,N_12261,N_12731);
and U13222 (N_13222,N_12642,N_12748);
nand U13223 (N_13223,N_12545,N_12735);
nor U13224 (N_13224,N_12277,N_12335);
and U13225 (N_13225,N_12703,N_12725);
xnor U13226 (N_13226,N_12351,N_12687);
or U13227 (N_13227,N_12056,N_12046);
nor U13228 (N_13228,N_12269,N_12493);
and U13229 (N_13229,N_12360,N_12329);
or U13230 (N_13230,N_12385,N_12439);
nand U13231 (N_13231,N_12368,N_12178);
nor U13232 (N_13232,N_12578,N_12080);
nand U13233 (N_13233,N_12426,N_12232);
nor U13234 (N_13234,N_12748,N_12460);
or U13235 (N_13235,N_12544,N_12492);
and U13236 (N_13236,N_12314,N_12472);
and U13237 (N_13237,N_12078,N_12537);
nand U13238 (N_13238,N_12038,N_12059);
nand U13239 (N_13239,N_12203,N_12108);
and U13240 (N_13240,N_12125,N_12654);
nand U13241 (N_13241,N_12355,N_12478);
nand U13242 (N_13242,N_12115,N_12629);
and U13243 (N_13243,N_12041,N_12281);
nor U13244 (N_13244,N_12731,N_12387);
nor U13245 (N_13245,N_12368,N_12667);
or U13246 (N_13246,N_12581,N_12631);
and U13247 (N_13247,N_12441,N_12091);
nor U13248 (N_13248,N_12003,N_12508);
nor U13249 (N_13249,N_12116,N_12163);
and U13250 (N_13250,N_12420,N_12326);
nor U13251 (N_13251,N_12159,N_12164);
and U13252 (N_13252,N_12593,N_12646);
nand U13253 (N_13253,N_12211,N_12086);
nor U13254 (N_13254,N_12561,N_12377);
or U13255 (N_13255,N_12638,N_12602);
nand U13256 (N_13256,N_12358,N_12131);
nand U13257 (N_13257,N_12548,N_12710);
and U13258 (N_13258,N_12112,N_12185);
and U13259 (N_13259,N_12626,N_12679);
and U13260 (N_13260,N_12205,N_12401);
or U13261 (N_13261,N_12383,N_12121);
nand U13262 (N_13262,N_12463,N_12666);
nor U13263 (N_13263,N_12416,N_12005);
and U13264 (N_13264,N_12737,N_12146);
nor U13265 (N_13265,N_12577,N_12736);
nand U13266 (N_13266,N_12143,N_12087);
and U13267 (N_13267,N_12606,N_12536);
or U13268 (N_13268,N_12664,N_12037);
nand U13269 (N_13269,N_12748,N_12104);
or U13270 (N_13270,N_12666,N_12248);
or U13271 (N_13271,N_12331,N_12248);
and U13272 (N_13272,N_12327,N_12383);
and U13273 (N_13273,N_12577,N_12476);
nand U13274 (N_13274,N_12235,N_12641);
nand U13275 (N_13275,N_12212,N_12386);
nand U13276 (N_13276,N_12259,N_12030);
nand U13277 (N_13277,N_12317,N_12139);
nand U13278 (N_13278,N_12172,N_12236);
and U13279 (N_13279,N_12046,N_12457);
nor U13280 (N_13280,N_12274,N_12642);
or U13281 (N_13281,N_12233,N_12330);
xor U13282 (N_13282,N_12445,N_12050);
nor U13283 (N_13283,N_12290,N_12490);
xor U13284 (N_13284,N_12476,N_12126);
nor U13285 (N_13285,N_12090,N_12384);
nand U13286 (N_13286,N_12684,N_12351);
or U13287 (N_13287,N_12048,N_12290);
nor U13288 (N_13288,N_12532,N_12561);
nor U13289 (N_13289,N_12226,N_12676);
and U13290 (N_13290,N_12061,N_12623);
or U13291 (N_13291,N_12076,N_12604);
nand U13292 (N_13292,N_12592,N_12202);
or U13293 (N_13293,N_12371,N_12116);
nor U13294 (N_13294,N_12057,N_12487);
nor U13295 (N_13295,N_12737,N_12461);
and U13296 (N_13296,N_12527,N_12531);
nand U13297 (N_13297,N_12179,N_12536);
and U13298 (N_13298,N_12520,N_12132);
nor U13299 (N_13299,N_12393,N_12222);
nand U13300 (N_13300,N_12635,N_12009);
nor U13301 (N_13301,N_12582,N_12067);
or U13302 (N_13302,N_12635,N_12390);
and U13303 (N_13303,N_12429,N_12354);
and U13304 (N_13304,N_12565,N_12061);
nand U13305 (N_13305,N_12040,N_12403);
or U13306 (N_13306,N_12620,N_12729);
nor U13307 (N_13307,N_12349,N_12484);
nand U13308 (N_13308,N_12336,N_12046);
or U13309 (N_13309,N_12648,N_12605);
and U13310 (N_13310,N_12045,N_12061);
and U13311 (N_13311,N_12185,N_12654);
nand U13312 (N_13312,N_12255,N_12407);
or U13313 (N_13313,N_12185,N_12317);
or U13314 (N_13314,N_12028,N_12488);
nand U13315 (N_13315,N_12021,N_12033);
and U13316 (N_13316,N_12052,N_12746);
nor U13317 (N_13317,N_12592,N_12258);
nor U13318 (N_13318,N_12563,N_12617);
and U13319 (N_13319,N_12470,N_12233);
or U13320 (N_13320,N_12183,N_12106);
nor U13321 (N_13321,N_12412,N_12086);
nor U13322 (N_13322,N_12627,N_12611);
nand U13323 (N_13323,N_12245,N_12203);
xnor U13324 (N_13324,N_12162,N_12614);
nand U13325 (N_13325,N_12501,N_12156);
or U13326 (N_13326,N_12355,N_12085);
nand U13327 (N_13327,N_12478,N_12667);
nor U13328 (N_13328,N_12720,N_12693);
or U13329 (N_13329,N_12659,N_12446);
and U13330 (N_13330,N_12419,N_12638);
nor U13331 (N_13331,N_12704,N_12741);
and U13332 (N_13332,N_12438,N_12488);
or U13333 (N_13333,N_12266,N_12029);
and U13334 (N_13334,N_12539,N_12094);
or U13335 (N_13335,N_12323,N_12458);
or U13336 (N_13336,N_12149,N_12534);
nand U13337 (N_13337,N_12278,N_12569);
nand U13338 (N_13338,N_12133,N_12328);
and U13339 (N_13339,N_12411,N_12391);
nand U13340 (N_13340,N_12674,N_12715);
nand U13341 (N_13341,N_12380,N_12300);
and U13342 (N_13342,N_12352,N_12069);
nand U13343 (N_13343,N_12517,N_12271);
and U13344 (N_13344,N_12100,N_12302);
xnor U13345 (N_13345,N_12368,N_12674);
or U13346 (N_13346,N_12681,N_12619);
nand U13347 (N_13347,N_12494,N_12347);
or U13348 (N_13348,N_12618,N_12700);
and U13349 (N_13349,N_12193,N_12410);
or U13350 (N_13350,N_12687,N_12611);
nor U13351 (N_13351,N_12389,N_12233);
and U13352 (N_13352,N_12513,N_12478);
or U13353 (N_13353,N_12377,N_12453);
or U13354 (N_13354,N_12085,N_12574);
nor U13355 (N_13355,N_12440,N_12287);
nand U13356 (N_13356,N_12311,N_12322);
nand U13357 (N_13357,N_12497,N_12739);
nor U13358 (N_13358,N_12021,N_12388);
nor U13359 (N_13359,N_12521,N_12730);
nor U13360 (N_13360,N_12548,N_12300);
nand U13361 (N_13361,N_12309,N_12638);
or U13362 (N_13362,N_12063,N_12461);
and U13363 (N_13363,N_12631,N_12655);
xor U13364 (N_13364,N_12566,N_12225);
nand U13365 (N_13365,N_12441,N_12697);
nand U13366 (N_13366,N_12058,N_12173);
nor U13367 (N_13367,N_12050,N_12242);
and U13368 (N_13368,N_12220,N_12294);
nand U13369 (N_13369,N_12670,N_12699);
nand U13370 (N_13370,N_12438,N_12344);
or U13371 (N_13371,N_12089,N_12227);
or U13372 (N_13372,N_12205,N_12443);
nand U13373 (N_13373,N_12544,N_12079);
and U13374 (N_13374,N_12531,N_12055);
or U13375 (N_13375,N_12640,N_12357);
nor U13376 (N_13376,N_12068,N_12371);
nand U13377 (N_13377,N_12332,N_12386);
or U13378 (N_13378,N_12242,N_12530);
nor U13379 (N_13379,N_12140,N_12654);
or U13380 (N_13380,N_12272,N_12347);
or U13381 (N_13381,N_12478,N_12651);
and U13382 (N_13382,N_12383,N_12448);
nor U13383 (N_13383,N_12629,N_12380);
and U13384 (N_13384,N_12353,N_12365);
nand U13385 (N_13385,N_12013,N_12419);
or U13386 (N_13386,N_12083,N_12160);
or U13387 (N_13387,N_12494,N_12681);
or U13388 (N_13388,N_12678,N_12508);
nand U13389 (N_13389,N_12086,N_12355);
and U13390 (N_13390,N_12133,N_12742);
and U13391 (N_13391,N_12639,N_12347);
and U13392 (N_13392,N_12435,N_12116);
or U13393 (N_13393,N_12321,N_12659);
nor U13394 (N_13394,N_12481,N_12476);
nor U13395 (N_13395,N_12538,N_12312);
and U13396 (N_13396,N_12482,N_12548);
and U13397 (N_13397,N_12096,N_12259);
nor U13398 (N_13398,N_12395,N_12166);
and U13399 (N_13399,N_12684,N_12309);
nor U13400 (N_13400,N_12022,N_12374);
or U13401 (N_13401,N_12595,N_12291);
nand U13402 (N_13402,N_12112,N_12194);
nand U13403 (N_13403,N_12497,N_12501);
or U13404 (N_13404,N_12622,N_12439);
and U13405 (N_13405,N_12503,N_12654);
and U13406 (N_13406,N_12603,N_12391);
nand U13407 (N_13407,N_12687,N_12585);
nor U13408 (N_13408,N_12356,N_12075);
and U13409 (N_13409,N_12131,N_12559);
nand U13410 (N_13410,N_12710,N_12361);
nand U13411 (N_13411,N_12599,N_12310);
nor U13412 (N_13412,N_12247,N_12327);
and U13413 (N_13413,N_12637,N_12040);
and U13414 (N_13414,N_12303,N_12528);
nand U13415 (N_13415,N_12169,N_12273);
nor U13416 (N_13416,N_12542,N_12372);
or U13417 (N_13417,N_12604,N_12650);
and U13418 (N_13418,N_12067,N_12396);
or U13419 (N_13419,N_12391,N_12239);
and U13420 (N_13420,N_12307,N_12540);
or U13421 (N_13421,N_12732,N_12311);
and U13422 (N_13422,N_12141,N_12669);
nor U13423 (N_13423,N_12100,N_12639);
or U13424 (N_13424,N_12032,N_12210);
nand U13425 (N_13425,N_12748,N_12302);
nand U13426 (N_13426,N_12176,N_12337);
and U13427 (N_13427,N_12667,N_12636);
or U13428 (N_13428,N_12396,N_12361);
or U13429 (N_13429,N_12436,N_12408);
nor U13430 (N_13430,N_12462,N_12540);
nand U13431 (N_13431,N_12563,N_12169);
and U13432 (N_13432,N_12452,N_12088);
nor U13433 (N_13433,N_12343,N_12426);
nor U13434 (N_13434,N_12631,N_12342);
xnor U13435 (N_13435,N_12537,N_12562);
and U13436 (N_13436,N_12353,N_12529);
nor U13437 (N_13437,N_12318,N_12560);
or U13438 (N_13438,N_12168,N_12538);
nor U13439 (N_13439,N_12447,N_12317);
or U13440 (N_13440,N_12241,N_12521);
nor U13441 (N_13441,N_12210,N_12684);
nor U13442 (N_13442,N_12221,N_12546);
and U13443 (N_13443,N_12234,N_12330);
nand U13444 (N_13444,N_12571,N_12363);
nand U13445 (N_13445,N_12494,N_12245);
or U13446 (N_13446,N_12587,N_12501);
nor U13447 (N_13447,N_12385,N_12296);
nand U13448 (N_13448,N_12506,N_12742);
nor U13449 (N_13449,N_12115,N_12036);
nor U13450 (N_13450,N_12047,N_12703);
nor U13451 (N_13451,N_12413,N_12618);
or U13452 (N_13452,N_12509,N_12653);
or U13453 (N_13453,N_12746,N_12154);
and U13454 (N_13454,N_12376,N_12600);
nor U13455 (N_13455,N_12409,N_12016);
or U13456 (N_13456,N_12083,N_12001);
nand U13457 (N_13457,N_12114,N_12670);
nand U13458 (N_13458,N_12290,N_12646);
nor U13459 (N_13459,N_12100,N_12290);
and U13460 (N_13460,N_12602,N_12655);
nor U13461 (N_13461,N_12615,N_12484);
nor U13462 (N_13462,N_12024,N_12230);
or U13463 (N_13463,N_12108,N_12533);
nor U13464 (N_13464,N_12358,N_12476);
and U13465 (N_13465,N_12549,N_12309);
nand U13466 (N_13466,N_12062,N_12608);
or U13467 (N_13467,N_12312,N_12078);
or U13468 (N_13468,N_12031,N_12300);
and U13469 (N_13469,N_12694,N_12733);
and U13470 (N_13470,N_12712,N_12269);
nor U13471 (N_13471,N_12185,N_12673);
and U13472 (N_13472,N_12712,N_12307);
nand U13473 (N_13473,N_12578,N_12079);
nor U13474 (N_13474,N_12001,N_12487);
and U13475 (N_13475,N_12061,N_12580);
nor U13476 (N_13476,N_12193,N_12578);
or U13477 (N_13477,N_12656,N_12049);
or U13478 (N_13478,N_12524,N_12327);
nor U13479 (N_13479,N_12156,N_12210);
and U13480 (N_13480,N_12645,N_12117);
and U13481 (N_13481,N_12409,N_12607);
and U13482 (N_13482,N_12620,N_12456);
nand U13483 (N_13483,N_12045,N_12435);
and U13484 (N_13484,N_12627,N_12413);
nor U13485 (N_13485,N_12660,N_12721);
and U13486 (N_13486,N_12090,N_12395);
nand U13487 (N_13487,N_12731,N_12591);
nand U13488 (N_13488,N_12604,N_12451);
and U13489 (N_13489,N_12202,N_12626);
or U13490 (N_13490,N_12070,N_12504);
nand U13491 (N_13491,N_12515,N_12473);
or U13492 (N_13492,N_12214,N_12206);
nand U13493 (N_13493,N_12111,N_12506);
xnor U13494 (N_13494,N_12455,N_12692);
and U13495 (N_13495,N_12440,N_12283);
or U13496 (N_13496,N_12497,N_12240);
or U13497 (N_13497,N_12225,N_12580);
and U13498 (N_13498,N_12287,N_12138);
nor U13499 (N_13499,N_12082,N_12462);
or U13500 (N_13500,N_12985,N_12976);
nand U13501 (N_13501,N_12758,N_13428);
or U13502 (N_13502,N_12920,N_13269);
nor U13503 (N_13503,N_13413,N_13482);
or U13504 (N_13504,N_12944,N_12861);
and U13505 (N_13505,N_13388,N_13405);
nand U13506 (N_13506,N_13013,N_12785);
or U13507 (N_13507,N_12755,N_12889);
nor U13508 (N_13508,N_13445,N_13422);
or U13509 (N_13509,N_12827,N_13462);
nor U13510 (N_13510,N_13147,N_13120);
or U13511 (N_13511,N_13232,N_12899);
or U13512 (N_13512,N_13281,N_13054);
nor U13513 (N_13513,N_12965,N_13478);
and U13514 (N_13514,N_12845,N_13392);
nand U13515 (N_13515,N_13200,N_13471);
or U13516 (N_13516,N_13035,N_13167);
nand U13517 (N_13517,N_12967,N_13144);
or U13518 (N_13518,N_12959,N_13334);
and U13519 (N_13519,N_12906,N_13240);
nand U13520 (N_13520,N_13172,N_13412);
or U13521 (N_13521,N_13248,N_13131);
or U13522 (N_13522,N_13489,N_12879);
nand U13523 (N_13523,N_12805,N_13457);
nand U13524 (N_13524,N_13123,N_12975);
or U13525 (N_13525,N_13355,N_12886);
nand U13526 (N_13526,N_13448,N_13215);
nand U13527 (N_13527,N_12860,N_13365);
xnor U13528 (N_13528,N_12999,N_13488);
nand U13529 (N_13529,N_13330,N_12995);
and U13530 (N_13530,N_13094,N_13235);
and U13531 (N_13531,N_13310,N_13254);
or U13532 (N_13532,N_13197,N_12790);
and U13533 (N_13533,N_12918,N_13111);
nor U13534 (N_13534,N_13370,N_13433);
and U13535 (N_13535,N_13188,N_12838);
nand U13536 (N_13536,N_13325,N_13135);
nand U13537 (N_13537,N_13132,N_12907);
or U13538 (N_13538,N_12777,N_13446);
nand U13539 (N_13539,N_13491,N_13026);
or U13540 (N_13540,N_13395,N_12974);
and U13541 (N_13541,N_12816,N_12983);
nand U13542 (N_13542,N_13309,N_12941);
and U13543 (N_13543,N_13307,N_12798);
nand U13544 (N_13544,N_13487,N_12882);
nand U13545 (N_13545,N_12839,N_13225);
nor U13546 (N_13546,N_13202,N_12997);
and U13547 (N_13547,N_12817,N_13377);
and U13548 (N_13548,N_13440,N_12964);
nand U13549 (N_13549,N_13192,N_12802);
nor U13550 (N_13550,N_12856,N_13461);
or U13551 (N_13551,N_13436,N_13088);
nor U13552 (N_13552,N_13438,N_13027);
nand U13553 (N_13553,N_12836,N_12949);
and U13554 (N_13554,N_12915,N_13483);
or U13555 (N_13555,N_12822,N_13110);
nand U13556 (N_13556,N_13250,N_12771);
nor U13557 (N_13557,N_13329,N_12801);
or U13558 (N_13558,N_13317,N_12939);
nor U13559 (N_13559,N_13300,N_13162);
nand U13560 (N_13560,N_13205,N_13425);
and U13561 (N_13561,N_13157,N_12951);
or U13562 (N_13562,N_13391,N_13453);
nand U13563 (N_13563,N_13118,N_12929);
and U13564 (N_13564,N_13015,N_12911);
nor U13565 (N_13565,N_12862,N_13020);
and U13566 (N_13566,N_13130,N_13077);
and U13567 (N_13567,N_13382,N_12966);
nor U13568 (N_13568,N_13140,N_13262);
nand U13569 (N_13569,N_13459,N_13229);
or U13570 (N_13570,N_13348,N_13354);
nand U13571 (N_13571,N_13010,N_13369);
and U13572 (N_13572,N_13091,N_12853);
and U13573 (N_13573,N_12787,N_13170);
nor U13574 (N_13574,N_13148,N_13237);
and U13575 (N_13575,N_13275,N_12783);
or U13576 (N_13576,N_13164,N_13253);
nand U13577 (N_13577,N_13326,N_13302);
nand U13578 (N_13578,N_13117,N_13180);
and U13579 (N_13579,N_12992,N_12952);
nand U13580 (N_13580,N_13420,N_13342);
nor U13581 (N_13581,N_13485,N_13469);
or U13582 (N_13582,N_13203,N_12973);
or U13583 (N_13583,N_13086,N_13336);
and U13584 (N_13584,N_12767,N_13360);
and U13585 (N_13585,N_12796,N_13021);
nor U13586 (N_13586,N_12931,N_13181);
nor U13587 (N_13587,N_13076,N_13107);
nor U13588 (N_13588,N_13353,N_13373);
or U13589 (N_13589,N_13198,N_12979);
or U13590 (N_13590,N_12812,N_12971);
or U13591 (N_13591,N_13340,N_13109);
nor U13592 (N_13592,N_13152,N_12900);
and U13593 (N_13593,N_12769,N_13403);
or U13594 (N_13594,N_12823,N_13318);
nand U13595 (N_13595,N_12909,N_13447);
and U13596 (N_13596,N_13492,N_12884);
nor U13597 (N_13597,N_13092,N_13289);
or U13598 (N_13598,N_13243,N_13264);
and U13599 (N_13599,N_13137,N_13190);
and U13600 (N_13600,N_13146,N_13093);
nor U13601 (N_13601,N_13233,N_13335);
or U13602 (N_13602,N_12828,N_13345);
and U13603 (N_13603,N_13291,N_12814);
nor U13604 (N_13604,N_13087,N_13106);
or U13605 (N_13605,N_12818,N_13038);
xor U13606 (N_13606,N_13383,N_13134);
nor U13607 (N_13607,N_13333,N_13443);
and U13608 (N_13608,N_13299,N_12766);
and U13609 (N_13609,N_12922,N_12854);
and U13610 (N_13610,N_12926,N_12978);
and U13611 (N_13611,N_13372,N_13430);
xor U13612 (N_13612,N_13227,N_12935);
and U13613 (N_13613,N_13398,N_13286);
and U13614 (N_13614,N_13356,N_13418);
and U13615 (N_13615,N_12924,N_13173);
and U13616 (N_13616,N_13400,N_13136);
nor U13617 (N_13617,N_13217,N_13401);
nand U13618 (N_13618,N_13272,N_13016);
nor U13619 (N_13619,N_12994,N_12969);
nand U13620 (N_13620,N_12940,N_13151);
and U13621 (N_13621,N_13359,N_12848);
and U13622 (N_13622,N_13085,N_13404);
nor U13623 (N_13623,N_13429,N_12768);
and U13624 (N_13624,N_13175,N_13458);
and U13625 (N_13625,N_12987,N_13384);
nor U13626 (N_13626,N_12989,N_12923);
or U13627 (N_13627,N_13411,N_13319);
and U13628 (N_13628,N_12855,N_13211);
and U13629 (N_13629,N_13075,N_13285);
or U13630 (N_13630,N_12968,N_12874);
and U13631 (N_13631,N_12819,N_13268);
or U13632 (N_13632,N_13025,N_12869);
or U13633 (N_13633,N_13399,N_13174);
nor U13634 (N_13634,N_13207,N_13049);
nor U13635 (N_13635,N_13150,N_13274);
nand U13636 (N_13636,N_13468,N_13176);
and U13637 (N_13637,N_13257,N_13009);
nand U13638 (N_13638,N_12916,N_13368);
nand U13639 (N_13639,N_12793,N_13361);
and U13640 (N_13640,N_12808,N_13431);
nand U13641 (N_13641,N_12942,N_12998);
nand U13642 (N_13642,N_12880,N_13260);
xor U13643 (N_13643,N_12866,N_13407);
nand U13644 (N_13644,N_13273,N_13244);
nand U13645 (N_13645,N_12847,N_13432);
nor U13646 (N_13646,N_13100,N_13113);
nor U13647 (N_13647,N_13182,N_13321);
nand U13648 (N_13648,N_13474,N_13078);
nand U13649 (N_13649,N_13320,N_13350);
nor U13650 (N_13650,N_13141,N_12763);
nand U13651 (N_13651,N_13246,N_13393);
and U13652 (N_13652,N_12779,N_13160);
nor U13653 (N_13653,N_13270,N_13464);
nor U13654 (N_13654,N_13331,N_12774);
nand U13655 (N_13655,N_13218,N_13213);
nor U13656 (N_13656,N_12864,N_13105);
nand U13657 (N_13657,N_13071,N_13435);
and U13658 (N_13658,N_13024,N_13366);
or U13659 (N_13659,N_13470,N_13357);
xnor U13660 (N_13660,N_13138,N_13067);
or U13661 (N_13661,N_13278,N_12938);
nand U13662 (N_13662,N_13389,N_12833);
nand U13663 (N_13663,N_12908,N_13011);
nor U13664 (N_13664,N_12858,N_13259);
and U13665 (N_13665,N_13362,N_13060);
nand U13666 (N_13666,N_13158,N_13014);
or U13667 (N_13667,N_13466,N_13378);
or U13668 (N_13668,N_13165,N_12986);
nor U13669 (N_13669,N_13096,N_12895);
or U13670 (N_13670,N_13312,N_13284);
nor U13671 (N_13671,N_13454,N_12753);
nor U13672 (N_13672,N_13417,N_12868);
nand U13673 (N_13673,N_13031,N_13245);
nand U13674 (N_13674,N_13338,N_12803);
or U13675 (N_13675,N_13301,N_13044);
or U13676 (N_13676,N_13292,N_13328);
and U13677 (N_13677,N_13481,N_13099);
and U13678 (N_13678,N_12914,N_12844);
or U13679 (N_13679,N_12825,N_13479);
or U13680 (N_13680,N_12961,N_13496);
and U13681 (N_13681,N_12843,N_13406);
or U13682 (N_13682,N_12821,N_13293);
and U13683 (N_13683,N_12933,N_12917);
and U13684 (N_13684,N_12757,N_13064);
or U13685 (N_13685,N_12878,N_13012);
nor U13686 (N_13686,N_13102,N_13287);
nor U13687 (N_13687,N_12958,N_13062);
nand U13688 (N_13688,N_13121,N_12988);
and U13689 (N_13689,N_13374,N_12863);
nand U13690 (N_13690,N_13222,N_13452);
nand U13691 (N_13691,N_13179,N_13019);
nor U13692 (N_13692,N_13005,N_13006);
and U13693 (N_13693,N_13041,N_13081);
and U13694 (N_13694,N_13122,N_13212);
and U13695 (N_13695,N_13097,N_13280);
or U13696 (N_13696,N_12934,N_13421);
nand U13697 (N_13697,N_12780,N_13056);
or U13698 (N_13698,N_13294,N_12993);
nand U13699 (N_13699,N_13456,N_13112);
nor U13700 (N_13700,N_13143,N_12772);
nor U13701 (N_13701,N_13022,N_13476);
nand U13702 (N_13702,N_13344,N_13234);
or U13703 (N_13703,N_13467,N_12813);
nand U13704 (N_13704,N_13042,N_13313);
or U13705 (N_13705,N_12789,N_13206);
and U13706 (N_13706,N_13163,N_12782);
xnor U13707 (N_13707,N_12751,N_13032);
nor U13708 (N_13708,N_13339,N_12857);
or U13709 (N_13709,N_12752,N_12897);
and U13710 (N_13710,N_13437,N_12764);
and U13711 (N_13711,N_13367,N_13178);
or U13712 (N_13712,N_12794,N_12811);
or U13713 (N_13713,N_13073,N_12829);
or U13714 (N_13714,N_12877,N_13463);
and U13715 (N_13715,N_13104,N_13166);
nand U13716 (N_13716,N_13415,N_12791);
or U13717 (N_13717,N_13002,N_12797);
nor U13718 (N_13718,N_13186,N_13480);
nor U13719 (N_13719,N_13477,N_12842);
or U13720 (N_13720,N_13171,N_12936);
nand U13721 (N_13721,N_12902,N_13155);
or U13722 (N_13722,N_13195,N_13231);
or U13723 (N_13723,N_13139,N_13189);
and U13724 (N_13724,N_13039,N_12851);
or U13725 (N_13725,N_12883,N_13379);
nor U13726 (N_13726,N_12826,N_12996);
and U13727 (N_13727,N_13057,N_13265);
nand U13728 (N_13728,N_13089,N_13177);
nand U13729 (N_13729,N_13442,N_13380);
and U13730 (N_13730,N_13126,N_13169);
and U13731 (N_13731,N_13376,N_13423);
and U13732 (N_13732,N_13266,N_12800);
nor U13733 (N_13733,N_13305,N_13303);
and U13734 (N_13734,N_12792,N_12765);
or U13735 (N_13735,N_12913,N_13204);
nor U13736 (N_13736,N_12840,N_13059);
nand U13737 (N_13737,N_12865,N_13224);
or U13738 (N_13738,N_13018,N_13416);
or U13739 (N_13739,N_13043,N_13494);
nor U13740 (N_13740,N_12948,N_13133);
or U13741 (N_13741,N_13346,N_13271);
or U13742 (N_13742,N_12946,N_12891);
nand U13743 (N_13743,N_13115,N_12852);
or U13744 (N_13744,N_13238,N_13068);
nor U13745 (N_13745,N_13475,N_13324);
or U13746 (N_13746,N_12770,N_13154);
or U13747 (N_13747,N_12873,N_12898);
and U13748 (N_13748,N_12972,N_13079);
and U13749 (N_13749,N_12953,N_12799);
or U13750 (N_13750,N_13114,N_13397);
nand U13751 (N_13751,N_12990,N_12809);
and U13752 (N_13752,N_13125,N_13072);
nand U13753 (N_13753,N_13220,N_13315);
or U13754 (N_13754,N_12982,N_13101);
and U13755 (N_13755,N_12778,N_13290);
nor U13756 (N_13756,N_13036,N_13352);
xor U13757 (N_13757,N_13095,N_12831);
nor U13758 (N_13758,N_12956,N_13277);
nand U13759 (N_13759,N_13082,N_12788);
or U13760 (N_13760,N_13098,N_13451);
or U13761 (N_13761,N_13124,N_12919);
and U13762 (N_13762,N_13047,N_12815);
and U13763 (N_13763,N_13033,N_13194);
nor U13764 (N_13764,N_12773,N_12921);
nand U13765 (N_13765,N_13298,N_12810);
or U13766 (N_13766,N_13490,N_12804);
nor U13767 (N_13767,N_12981,N_12962);
and U13768 (N_13768,N_12903,N_13048);
nor U13769 (N_13769,N_13046,N_13424);
nor U13770 (N_13770,N_13156,N_13055);
and U13771 (N_13771,N_13444,N_12837);
nand U13772 (N_13772,N_12781,N_13050);
and U13773 (N_13773,N_13001,N_13053);
nor U13774 (N_13774,N_13028,N_13385);
or U13775 (N_13775,N_12859,N_12945);
nand U13776 (N_13776,N_13267,N_13441);
nor U13777 (N_13777,N_13185,N_13003);
or U13778 (N_13778,N_12888,N_13375);
or U13779 (N_13779,N_13247,N_12784);
and U13780 (N_13780,N_12832,N_13484);
nand U13781 (N_13781,N_12887,N_13037);
and U13782 (N_13782,N_12977,N_13108);
or U13783 (N_13783,N_13023,N_13201);
or U13784 (N_13784,N_13450,N_13261);
and U13785 (N_13785,N_13351,N_12960);
nor U13786 (N_13786,N_12830,N_13127);
and U13787 (N_13787,N_12943,N_13061);
nor U13788 (N_13788,N_13343,N_13030);
and U13789 (N_13789,N_13323,N_13396);
nand U13790 (N_13790,N_12876,N_12954);
and U13791 (N_13791,N_12756,N_13486);
nand U13792 (N_13792,N_13223,N_12991);
nand U13793 (N_13793,N_12925,N_12905);
and U13794 (N_13794,N_13145,N_13034);
or U13795 (N_13795,N_13080,N_13239);
nand U13796 (N_13796,N_12937,N_12947);
and U13797 (N_13797,N_13439,N_13304);
nor U13798 (N_13798,N_12754,N_13210);
nand U13799 (N_13799,N_13337,N_13187);
nor U13800 (N_13800,N_13465,N_12872);
or U13801 (N_13801,N_13308,N_12850);
xor U13802 (N_13802,N_12759,N_13381);
and U13803 (N_13803,N_12807,N_12875);
and U13804 (N_13804,N_13000,N_13084);
and U13805 (N_13805,N_13371,N_13449);
nor U13806 (N_13806,N_13394,N_12760);
and U13807 (N_13807,N_12834,N_12896);
or U13808 (N_13808,N_13161,N_13322);
nand U13809 (N_13809,N_12871,N_12932);
or U13810 (N_13810,N_13159,N_13347);
nor U13811 (N_13811,N_13341,N_13142);
nand U13812 (N_13812,N_13316,N_13363);
nand U13813 (N_13813,N_13258,N_12984);
nor U13814 (N_13814,N_12904,N_13065);
nand U13815 (N_13815,N_13069,N_13103);
nand U13816 (N_13816,N_13473,N_12955);
nor U13817 (N_13817,N_13007,N_13153);
nand U13818 (N_13818,N_13332,N_12980);
and U13819 (N_13819,N_13029,N_13252);
or U13820 (N_13820,N_13358,N_13236);
or U13821 (N_13821,N_13004,N_13311);
nor U13822 (N_13822,N_13184,N_12841);
and U13823 (N_13823,N_13455,N_13349);
nor U13824 (N_13824,N_13434,N_13149);
nand U13825 (N_13825,N_12867,N_12750);
nand U13826 (N_13826,N_13066,N_12890);
or U13827 (N_13827,N_13414,N_13498);
or U13828 (N_13828,N_13279,N_12910);
nor U13829 (N_13829,N_13472,N_13051);
and U13830 (N_13830,N_13387,N_13297);
or U13831 (N_13831,N_13497,N_13256);
xor U13832 (N_13832,N_12927,N_13410);
and U13833 (N_13833,N_13242,N_13074);
or U13834 (N_13834,N_12824,N_12806);
nor U13835 (N_13835,N_12761,N_13045);
nand U13836 (N_13836,N_13196,N_12892);
and U13837 (N_13837,N_13386,N_13209);
and U13838 (N_13838,N_12901,N_12776);
nand U13839 (N_13839,N_12963,N_13128);
or U13840 (N_13840,N_13306,N_13419);
xnor U13841 (N_13841,N_12893,N_13495);
xor U13842 (N_13842,N_13219,N_13426);
and U13843 (N_13843,N_13402,N_13070);
or U13844 (N_13844,N_13221,N_13255);
nor U13845 (N_13845,N_12795,N_13228);
and U13846 (N_13846,N_13327,N_12970);
or U13847 (N_13847,N_13364,N_13408);
and U13848 (N_13848,N_13119,N_13314);
or U13849 (N_13849,N_12762,N_13193);
and U13850 (N_13850,N_13040,N_13409);
or U13851 (N_13851,N_13199,N_13282);
or U13852 (N_13852,N_13283,N_13251);
or U13853 (N_13853,N_13083,N_12930);
nand U13854 (N_13854,N_13017,N_12846);
or U13855 (N_13855,N_13129,N_12786);
or U13856 (N_13856,N_13052,N_13295);
nand U13857 (N_13857,N_12928,N_13390);
nor U13858 (N_13858,N_13427,N_13230);
nor U13859 (N_13859,N_12849,N_12957);
or U13860 (N_13860,N_13216,N_13208);
and U13861 (N_13861,N_13168,N_13183);
or U13862 (N_13862,N_13296,N_12881);
nand U13863 (N_13863,N_13263,N_13288);
and U13864 (N_13864,N_13116,N_13008);
or U13865 (N_13865,N_13090,N_13058);
or U13866 (N_13866,N_13460,N_12775);
nand U13867 (N_13867,N_13063,N_12885);
nor U13868 (N_13868,N_12870,N_13499);
and U13869 (N_13869,N_13214,N_13191);
nor U13870 (N_13870,N_13249,N_12894);
nor U13871 (N_13871,N_12835,N_13276);
or U13872 (N_13872,N_12820,N_13241);
or U13873 (N_13873,N_13493,N_12912);
nor U13874 (N_13874,N_13226,N_12950);
and U13875 (N_13875,N_12904,N_13341);
nor U13876 (N_13876,N_12803,N_13231);
nor U13877 (N_13877,N_13074,N_12958);
and U13878 (N_13878,N_13048,N_12982);
and U13879 (N_13879,N_13402,N_13104);
nand U13880 (N_13880,N_13483,N_13033);
nor U13881 (N_13881,N_13408,N_12826);
nor U13882 (N_13882,N_13097,N_13116);
nor U13883 (N_13883,N_13141,N_12834);
or U13884 (N_13884,N_13271,N_13063);
nor U13885 (N_13885,N_13494,N_13004);
nand U13886 (N_13886,N_13022,N_13264);
or U13887 (N_13887,N_13155,N_12988);
and U13888 (N_13888,N_13023,N_13005);
and U13889 (N_13889,N_12842,N_13121);
nand U13890 (N_13890,N_13495,N_13029);
or U13891 (N_13891,N_13363,N_12831);
and U13892 (N_13892,N_13157,N_12921);
nand U13893 (N_13893,N_13229,N_13005);
or U13894 (N_13894,N_13380,N_13245);
or U13895 (N_13895,N_13461,N_13411);
nor U13896 (N_13896,N_13260,N_13417);
or U13897 (N_13897,N_13309,N_12871);
xnor U13898 (N_13898,N_13396,N_13339);
nor U13899 (N_13899,N_13087,N_12807);
nor U13900 (N_13900,N_13034,N_12779);
or U13901 (N_13901,N_12766,N_13237);
or U13902 (N_13902,N_13210,N_13259);
xor U13903 (N_13903,N_13099,N_13233);
nor U13904 (N_13904,N_13408,N_12803);
nand U13905 (N_13905,N_13394,N_13472);
nor U13906 (N_13906,N_13214,N_13066);
nand U13907 (N_13907,N_13291,N_13260);
or U13908 (N_13908,N_13364,N_13342);
nor U13909 (N_13909,N_13227,N_13097);
and U13910 (N_13910,N_12796,N_13019);
nor U13911 (N_13911,N_12840,N_13139);
and U13912 (N_13912,N_13376,N_13056);
nor U13913 (N_13913,N_12955,N_13069);
or U13914 (N_13914,N_13174,N_12958);
nand U13915 (N_13915,N_12982,N_13381);
and U13916 (N_13916,N_12966,N_13158);
nor U13917 (N_13917,N_13201,N_13496);
and U13918 (N_13918,N_12985,N_12897);
xor U13919 (N_13919,N_13450,N_12967);
and U13920 (N_13920,N_13233,N_13044);
nand U13921 (N_13921,N_13165,N_12945);
and U13922 (N_13922,N_12976,N_13161);
nand U13923 (N_13923,N_13004,N_12976);
and U13924 (N_13924,N_13491,N_13102);
and U13925 (N_13925,N_13156,N_13107);
or U13926 (N_13926,N_13117,N_13289);
and U13927 (N_13927,N_13270,N_13114);
nor U13928 (N_13928,N_13194,N_12903);
nand U13929 (N_13929,N_13128,N_12784);
nor U13930 (N_13930,N_13468,N_13297);
nor U13931 (N_13931,N_12986,N_13383);
nand U13932 (N_13932,N_13475,N_12793);
or U13933 (N_13933,N_13239,N_13307);
and U13934 (N_13934,N_13075,N_13363);
or U13935 (N_13935,N_12769,N_12863);
and U13936 (N_13936,N_13163,N_13111);
nand U13937 (N_13937,N_13297,N_13278);
and U13938 (N_13938,N_13483,N_13073);
nor U13939 (N_13939,N_13174,N_12849);
nand U13940 (N_13940,N_12801,N_12981);
nand U13941 (N_13941,N_13251,N_13389);
or U13942 (N_13942,N_12778,N_12827);
or U13943 (N_13943,N_13316,N_13345);
nor U13944 (N_13944,N_12954,N_13453);
or U13945 (N_13945,N_12750,N_13317);
nor U13946 (N_13946,N_13426,N_13337);
nor U13947 (N_13947,N_13286,N_13071);
nand U13948 (N_13948,N_12957,N_12911);
and U13949 (N_13949,N_13184,N_12866);
or U13950 (N_13950,N_12842,N_12785);
or U13951 (N_13951,N_13248,N_13068);
or U13952 (N_13952,N_13346,N_13304);
nand U13953 (N_13953,N_13027,N_12967);
or U13954 (N_13954,N_12836,N_13030);
nand U13955 (N_13955,N_13457,N_12762);
nor U13956 (N_13956,N_12967,N_12936);
nand U13957 (N_13957,N_13454,N_12870);
or U13958 (N_13958,N_12924,N_13269);
and U13959 (N_13959,N_12756,N_12923);
nand U13960 (N_13960,N_13229,N_13278);
nor U13961 (N_13961,N_13486,N_13101);
and U13962 (N_13962,N_13151,N_13041);
nand U13963 (N_13963,N_13169,N_13449);
and U13964 (N_13964,N_13407,N_13205);
nand U13965 (N_13965,N_13417,N_13269);
nand U13966 (N_13966,N_13248,N_12902);
nand U13967 (N_13967,N_12786,N_12994);
nor U13968 (N_13968,N_12878,N_13454);
xor U13969 (N_13969,N_12920,N_12946);
and U13970 (N_13970,N_13255,N_12766);
nand U13971 (N_13971,N_13026,N_13140);
and U13972 (N_13972,N_13360,N_12919);
or U13973 (N_13973,N_13375,N_12912);
or U13974 (N_13974,N_13069,N_13493);
and U13975 (N_13975,N_13120,N_13111);
and U13976 (N_13976,N_12919,N_12796);
and U13977 (N_13977,N_13164,N_13336);
nand U13978 (N_13978,N_12927,N_13247);
nor U13979 (N_13979,N_12975,N_13007);
xor U13980 (N_13980,N_13089,N_12994);
nand U13981 (N_13981,N_13171,N_12842);
and U13982 (N_13982,N_13319,N_13168);
nor U13983 (N_13983,N_12800,N_12875);
and U13984 (N_13984,N_13200,N_13169);
or U13985 (N_13985,N_13377,N_13289);
nor U13986 (N_13986,N_12765,N_13482);
nor U13987 (N_13987,N_13389,N_13218);
and U13988 (N_13988,N_13188,N_13031);
xnor U13989 (N_13989,N_13255,N_13130);
nor U13990 (N_13990,N_13340,N_12797);
nor U13991 (N_13991,N_13214,N_13185);
nor U13992 (N_13992,N_13235,N_13002);
or U13993 (N_13993,N_12828,N_13306);
nand U13994 (N_13994,N_13257,N_13164);
nor U13995 (N_13995,N_13229,N_12979);
nand U13996 (N_13996,N_13342,N_13438);
xnor U13997 (N_13997,N_12831,N_12811);
nand U13998 (N_13998,N_13207,N_13201);
and U13999 (N_13999,N_13367,N_13498);
nor U14000 (N_14000,N_13302,N_13487);
nor U14001 (N_14001,N_13279,N_13167);
or U14002 (N_14002,N_13104,N_13335);
nor U14003 (N_14003,N_13130,N_13327);
xor U14004 (N_14004,N_12915,N_13179);
nor U14005 (N_14005,N_13221,N_13000);
and U14006 (N_14006,N_13228,N_13319);
nand U14007 (N_14007,N_12769,N_13120);
and U14008 (N_14008,N_13086,N_12777);
or U14009 (N_14009,N_13141,N_12914);
and U14010 (N_14010,N_13263,N_13428);
and U14011 (N_14011,N_12881,N_13399);
nor U14012 (N_14012,N_13043,N_13473);
nor U14013 (N_14013,N_12762,N_13352);
or U14014 (N_14014,N_13386,N_13170);
nand U14015 (N_14015,N_13171,N_12878);
nand U14016 (N_14016,N_13209,N_13434);
or U14017 (N_14017,N_13264,N_13262);
nor U14018 (N_14018,N_13170,N_13190);
nand U14019 (N_14019,N_13343,N_13392);
and U14020 (N_14020,N_13298,N_13134);
or U14021 (N_14021,N_13099,N_13052);
nand U14022 (N_14022,N_12939,N_13207);
nand U14023 (N_14023,N_12757,N_13314);
nand U14024 (N_14024,N_12791,N_13218);
nand U14025 (N_14025,N_13132,N_13056);
or U14026 (N_14026,N_13076,N_13342);
nand U14027 (N_14027,N_12892,N_13384);
nor U14028 (N_14028,N_13174,N_12810);
xnor U14029 (N_14029,N_13404,N_13298);
or U14030 (N_14030,N_13228,N_13045);
and U14031 (N_14031,N_12993,N_13097);
nand U14032 (N_14032,N_12876,N_13235);
nor U14033 (N_14033,N_13332,N_12990);
nor U14034 (N_14034,N_12838,N_12985);
nor U14035 (N_14035,N_12901,N_12978);
nand U14036 (N_14036,N_13384,N_13459);
nor U14037 (N_14037,N_12984,N_13380);
or U14038 (N_14038,N_13210,N_13113);
and U14039 (N_14039,N_13251,N_13255);
or U14040 (N_14040,N_13389,N_12938);
nand U14041 (N_14041,N_13092,N_13245);
or U14042 (N_14042,N_13044,N_12794);
nor U14043 (N_14043,N_12908,N_12833);
or U14044 (N_14044,N_12857,N_12832);
or U14045 (N_14045,N_13179,N_12912);
nor U14046 (N_14046,N_12827,N_12905);
nand U14047 (N_14047,N_13380,N_13287);
and U14048 (N_14048,N_12826,N_13411);
and U14049 (N_14049,N_13220,N_12873);
or U14050 (N_14050,N_12782,N_12828);
xnor U14051 (N_14051,N_13139,N_13143);
and U14052 (N_14052,N_13334,N_12821);
or U14053 (N_14053,N_12934,N_13415);
or U14054 (N_14054,N_13204,N_12917);
or U14055 (N_14055,N_13400,N_13352);
nand U14056 (N_14056,N_12770,N_12990);
and U14057 (N_14057,N_13316,N_12832);
xor U14058 (N_14058,N_13020,N_13127);
or U14059 (N_14059,N_12878,N_13075);
nand U14060 (N_14060,N_13127,N_12758);
nor U14061 (N_14061,N_13311,N_13247);
nand U14062 (N_14062,N_13465,N_13317);
nor U14063 (N_14063,N_12854,N_13228);
nand U14064 (N_14064,N_12802,N_13383);
nor U14065 (N_14065,N_12813,N_13283);
xor U14066 (N_14066,N_13176,N_13144);
nand U14067 (N_14067,N_13204,N_13176);
or U14068 (N_14068,N_13251,N_12806);
nor U14069 (N_14069,N_12955,N_12751);
or U14070 (N_14070,N_12781,N_13271);
or U14071 (N_14071,N_12900,N_13443);
nand U14072 (N_14072,N_13465,N_13475);
nor U14073 (N_14073,N_12970,N_12776);
or U14074 (N_14074,N_13099,N_13265);
nor U14075 (N_14075,N_13092,N_13201);
nor U14076 (N_14076,N_13006,N_12790);
or U14077 (N_14077,N_13360,N_12782);
nand U14078 (N_14078,N_13293,N_13125);
nor U14079 (N_14079,N_12969,N_13286);
nand U14080 (N_14080,N_13344,N_13484);
or U14081 (N_14081,N_12919,N_12781);
and U14082 (N_14082,N_13078,N_13310);
or U14083 (N_14083,N_12870,N_13099);
nand U14084 (N_14084,N_13369,N_12952);
or U14085 (N_14085,N_13186,N_13283);
nor U14086 (N_14086,N_13367,N_12755);
nor U14087 (N_14087,N_13380,N_12875);
nand U14088 (N_14088,N_12887,N_13430);
nand U14089 (N_14089,N_13350,N_13448);
or U14090 (N_14090,N_13429,N_12767);
and U14091 (N_14091,N_13392,N_13212);
nor U14092 (N_14092,N_13242,N_13196);
or U14093 (N_14093,N_13167,N_13129);
xor U14094 (N_14094,N_12995,N_13213);
nor U14095 (N_14095,N_12858,N_12970);
or U14096 (N_14096,N_13209,N_13039);
nor U14097 (N_14097,N_13383,N_13246);
nor U14098 (N_14098,N_13281,N_13148);
or U14099 (N_14099,N_13182,N_12885);
nor U14100 (N_14100,N_13442,N_13418);
and U14101 (N_14101,N_13318,N_13411);
nor U14102 (N_14102,N_13331,N_12753);
nor U14103 (N_14103,N_12766,N_13095);
xnor U14104 (N_14104,N_13241,N_13342);
and U14105 (N_14105,N_12813,N_13448);
and U14106 (N_14106,N_12949,N_13406);
and U14107 (N_14107,N_13179,N_13397);
or U14108 (N_14108,N_12915,N_13494);
nand U14109 (N_14109,N_13378,N_13387);
nor U14110 (N_14110,N_13333,N_12819);
nand U14111 (N_14111,N_12801,N_12754);
nor U14112 (N_14112,N_12941,N_13349);
or U14113 (N_14113,N_13358,N_13093);
nor U14114 (N_14114,N_13361,N_12898);
or U14115 (N_14115,N_12835,N_13055);
and U14116 (N_14116,N_13363,N_13048);
nand U14117 (N_14117,N_12768,N_13227);
and U14118 (N_14118,N_13025,N_13419);
or U14119 (N_14119,N_13293,N_12967);
and U14120 (N_14120,N_12931,N_13178);
and U14121 (N_14121,N_12904,N_12767);
nand U14122 (N_14122,N_13230,N_12792);
or U14123 (N_14123,N_13060,N_13167);
nand U14124 (N_14124,N_13286,N_13195);
nand U14125 (N_14125,N_13181,N_13047);
or U14126 (N_14126,N_13156,N_13270);
xnor U14127 (N_14127,N_13071,N_12809);
nand U14128 (N_14128,N_13401,N_13325);
nand U14129 (N_14129,N_13428,N_13350);
nand U14130 (N_14130,N_12764,N_13195);
nor U14131 (N_14131,N_13234,N_13384);
and U14132 (N_14132,N_13343,N_12913);
and U14133 (N_14133,N_13490,N_13019);
or U14134 (N_14134,N_13070,N_13381);
nand U14135 (N_14135,N_13013,N_13192);
xor U14136 (N_14136,N_13217,N_12770);
or U14137 (N_14137,N_13426,N_13431);
nand U14138 (N_14138,N_13161,N_12754);
or U14139 (N_14139,N_12864,N_13035);
nor U14140 (N_14140,N_13221,N_12798);
or U14141 (N_14141,N_13207,N_13474);
and U14142 (N_14142,N_12895,N_12897);
or U14143 (N_14143,N_13261,N_12893);
nor U14144 (N_14144,N_12779,N_12900);
and U14145 (N_14145,N_12899,N_12959);
nand U14146 (N_14146,N_12983,N_12931);
and U14147 (N_14147,N_13063,N_12993);
nor U14148 (N_14148,N_12991,N_13221);
or U14149 (N_14149,N_13462,N_13082);
and U14150 (N_14150,N_13351,N_12852);
or U14151 (N_14151,N_13054,N_13178);
nor U14152 (N_14152,N_13038,N_13419);
nor U14153 (N_14153,N_13065,N_13482);
or U14154 (N_14154,N_13450,N_13374);
nor U14155 (N_14155,N_13323,N_12986);
or U14156 (N_14156,N_13083,N_13470);
nor U14157 (N_14157,N_13050,N_13370);
nand U14158 (N_14158,N_12788,N_12932);
or U14159 (N_14159,N_13435,N_13144);
and U14160 (N_14160,N_13132,N_13229);
and U14161 (N_14161,N_12755,N_13463);
nand U14162 (N_14162,N_13456,N_13432);
nor U14163 (N_14163,N_12784,N_13327);
or U14164 (N_14164,N_13020,N_13287);
or U14165 (N_14165,N_13212,N_13286);
nand U14166 (N_14166,N_12847,N_13024);
nand U14167 (N_14167,N_13297,N_12913);
nand U14168 (N_14168,N_13419,N_13006);
nand U14169 (N_14169,N_13340,N_13293);
and U14170 (N_14170,N_13051,N_12848);
or U14171 (N_14171,N_12882,N_12972);
nor U14172 (N_14172,N_13397,N_13400);
and U14173 (N_14173,N_12976,N_13294);
or U14174 (N_14174,N_13282,N_12821);
nor U14175 (N_14175,N_13241,N_13220);
or U14176 (N_14176,N_13412,N_13403);
and U14177 (N_14177,N_13364,N_13313);
or U14178 (N_14178,N_13196,N_13051);
and U14179 (N_14179,N_13465,N_12791);
and U14180 (N_14180,N_13371,N_13328);
nand U14181 (N_14181,N_13180,N_13485);
nand U14182 (N_14182,N_13485,N_13408);
and U14183 (N_14183,N_13350,N_13177);
or U14184 (N_14184,N_13367,N_12814);
or U14185 (N_14185,N_13006,N_13299);
nor U14186 (N_14186,N_12803,N_13094);
nand U14187 (N_14187,N_12773,N_12909);
nor U14188 (N_14188,N_12780,N_12794);
and U14189 (N_14189,N_13022,N_13487);
nand U14190 (N_14190,N_13245,N_12776);
and U14191 (N_14191,N_13370,N_13453);
or U14192 (N_14192,N_13196,N_13142);
or U14193 (N_14193,N_13497,N_13433);
nor U14194 (N_14194,N_13004,N_13147);
and U14195 (N_14195,N_13424,N_13284);
nand U14196 (N_14196,N_12920,N_12913);
nor U14197 (N_14197,N_13369,N_13323);
nand U14198 (N_14198,N_12956,N_13100);
or U14199 (N_14199,N_12881,N_12842);
nor U14200 (N_14200,N_13324,N_12866);
and U14201 (N_14201,N_12774,N_12897);
nor U14202 (N_14202,N_13021,N_13176);
nand U14203 (N_14203,N_13291,N_13109);
or U14204 (N_14204,N_13209,N_12905);
and U14205 (N_14205,N_12774,N_13219);
and U14206 (N_14206,N_13251,N_13232);
nand U14207 (N_14207,N_13077,N_13084);
and U14208 (N_14208,N_12818,N_13301);
nor U14209 (N_14209,N_12835,N_13296);
nor U14210 (N_14210,N_12810,N_12807);
or U14211 (N_14211,N_13226,N_13479);
or U14212 (N_14212,N_13186,N_13479);
and U14213 (N_14213,N_12940,N_12962);
nand U14214 (N_14214,N_13443,N_12930);
nand U14215 (N_14215,N_13140,N_12865);
nand U14216 (N_14216,N_13323,N_13378);
and U14217 (N_14217,N_13133,N_12944);
or U14218 (N_14218,N_13277,N_13180);
or U14219 (N_14219,N_13420,N_13004);
and U14220 (N_14220,N_13353,N_12863);
nand U14221 (N_14221,N_13240,N_13262);
and U14222 (N_14222,N_12914,N_13093);
or U14223 (N_14223,N_12839,N_13307);
nand U14224 (N_14224,N_13230,N_13241);
or U14225 (N_14225,N_13402,N_12831);
or U14226 (N_14226,N_13176,N_13052);
or U14227 (N_14227,N_13322,N_12766);
nand U14228 (N_14228,N_13321,N_13430);
nor U14229 (N_14229,N_13258,N_13194);
nand U14230 (N_14230,N_13189,N_13120);
or U14231 (N_14231,N_13143,N_12940);
or U14232 (N_14232,N_13118,N_13376);
nor U14233 (N_14233,N_13181,N_13197);
and U14234 (N_14234,N_13061,N_13429);
or U14235 (N_14235,N_13108,N_13060);
nand U14236 (N_14236,N_13039,N_13196);
or U14237 (N_14237,N_13379,N_13458);
nand U14238 (N_14238,N_13292,N_13461);
nor U14239 (N_14239,N_13439,N_12882);
or U14240 (N_14240,N_13046,N_13020);
nor U14241 (N_14241,N_13466,N_13374);
xor U14242 (N_14242,N_12995,N_13243);
nor U14243 (N_14243,N_13380,N_13045);
nor U14244 (N_14244,N_13280,N_13141);
or U14245 (N_14245,N_13308,N_13370);
and U14246 (N_14246,N_13419,N_12925);
or U14247 (N_14247,N_12821,N_12931);
nor U14248 (N_14248,N_13194,N_13164);
nor U14249 (N_14249,N_13140,N_13008);
and U14250 (N_14250,N_13865,N_13904);
and U14251 (N_14251,N_14145,N_13656);
nand U14252 (N_14252,N_13868,N_13636);
and U14253 (N_14253,N_13559,N_13926);
nor U14254 (N_14254,N_14097,N_13852);
or U14255 (N_14255,N_13693,N_13823);
nor U14256 (N_14256,N_13661,N_13505);
nand U14257 (N_14257,N_13531,N_13522);
nand U14258 (N_14258,N_14189,N_13795);
or U14259 (N_14259,N_14058,N_14209);
or U14260 (N_14260,N_13980,N_13681);
and U14261 (N_14261,N_13844,N_14013);
or U14262 (N_14262,N_13793,N_14221);
nor U14263 (N_14263,N_14152,N_13939);
or U14264 (N_14264,N_14077,N_13897);
and U14265 (N_14265,N_14089,N_13553);
nand U14266 (N_14266,N_13851,N_13564);
nand U14267 (N_14267,N_14102,N_13557);
nand U14268 (N_14268,N_13975,N_13994);
nor U14269 (N_14269,N_13736,N_13790);
nand U14270 (N_14270,N_13612,N_14178);
or U14271 (N_14271,N_13896,N_14092);
nand U14272 (N_14272,N_14166,N_14136);
and U14273 (N_14273,N_13739,N_13958);
nand U14274 (N_14274,N_14001,N_14017);
nand U14275 (N_14275,N_13758,N_13573);
and U14276 (N_14276,N_14227,N_14184);
nand U14277 (N_14277,N_13668,N_14248);
nor U14278 (N_14278,N_14067,N_13762);
nor U14279 (N_14279,N_13831,N_14146);
and U14280 (N_14280,N_13746,N_13922);
or U14281 (N_14281,N_13783,N_14037);
nand U14282 (N_14282,N_13871,N_13696);
nand U14283 (N_14283,N_13627,N_14132);
nand U14284 (N_14284,N_13749,N_13691);
nor U14285 (N_14285,N_13658,N_13609);
or U14286 (N_14286,N_13745,N_14150);
and U14287 (N_14287,N_14085,N_13524);
and U14288 (N_14288,N_14055,N_14099);
nand U14289 (N_14289,N_14235,N_14086);
nand U14290 (N_14290,N_14045,N_13504);
and U14291 (N_14291,N_13638,N_13796);
or U14292 (N_14292,N_14105,N_13833);
nor U14293 (N_14293,N_13990,N_13672);
and U14294 (N_14294,N_13754,N_13590);
or U14295 (N_14295,N_14149,N_14009);
nor U14296 (N_14296,N_14021,N_13792);
and U14297 (N_14297,N_13677,N_13953);
nor U14298 (N_14298,N_13785,N_13845);
and U14299 (N_14299,N_13921,N_13918);
or U14300 (N_14300,N_13512,N_14175);
and U14301 (N_14301,N_13560,N_13680);
or U14302 (N_14302,N_14199,N_14204);
and U14303 (N_14303,N_13563,N_13521);
or U14304 (N_14304,N_13752,N_14128);
nand U14305 (N_14305,N_14056,N_13731);
nor U14306 (N_14306,N_13525,N_13848);
nand U14307 (N_14307,N_13878,N_13641);
nand U14308 (N_14308,N_13809,N_13963);
nand U14309 (N_14309,N_13961,N_14074);
and U14310 (N_14310,N_14238,N_13695);
nand U14311 (N_14311,N_14114,N_13606);
nor U14312 (N_14312,N_13789,N_13890);
and U14313 (N_14313,N_13702,N_13633);
nor U14314 (N_14314,N_14063,N_13917);
and U14315 (N_14315,N_13712,N_13782);
xor U14316 (N_14316,N_13721,N_13663);
or U14317 (N_14317,N_13876,N_14088);
and U14318 (N_14318,N_13838,N_13503);
and U14319 (N_14319,N_14211,N_13931);
nand U14320 (N_14320,N_13808,N_13608);
nand U14321 (N_14321,N_14030,N_13613);
nor U14322 (N_14322,N_14006,N_13935);
and U14323 (N_14323,N_14070,N_13583);
and U14324 (N_14324,N_13856,N_14080);
nand U14325 (N_14325,N_13965,N_13631);
nand U14326 (N_14326,N_14069,N_13892);
nor U14327 (N_14327,N_13624,N_13690);
nand U14328 (N_14328,N_13944,N_13863);
nor U14329 (N_14329,N_14143,N_13618);
xor U14330 (N_14330,N_14072,N_14222);
nand U14331 (N_14331,N_13832,N_13692);
and U14332 (N_14332,N_13725,N_14148);
or U14333 (N_14333,N_14142,N_13942);
and U14334 (N_14334,N_13924,N_14025);
or U14335 (N_14335,N_13686,N_14188);
or U14336 (N_14336,N_13854,N_13555);
nand U14337 (N_14337,N_14062,N_13665);
nor U14338 (N_14338,N_14109,N_13666);
or U14339 (N_14339,N_14126,N_14223);
and U14340 (N_14340,N_14071,N_14024);
or U14341 (N_14341,N_13886,N_13533);
nor U14342 (N_14342,N_13649,N_13518);
or U14343 (N_14343,N_13750,N_13600);
or U14344 (N_14344,N_13577,N_13585);
nor U14345 (N_14345,N_13799,N_13826);
and U14346 (N_14346,N_13623,N_13891);
or U14347 (N_14347,N_13900,N_14120);
and U14348 (N_14348,N_13718,N_13753);
nand U14349 (N_14349,N_14231,N_13914);
nand U14350 (N_14350,N_13913,N_13956);
nand U14351 (N_14351,N_14113,N_14028);
nand U14352 (N_14352,N_13962,N_13574);
and U14353 (N_14353,N_13598,N_13902);
nand U14354 (N_14354,N_13787,N_13594);
or U14355 (N_14355,N_13768,N_13540);
or U14356 (N_14356,N_13757,N_13737);
nor U14357 (N_14357,N_13673,N_13669);
or U14358 (N_14358,N_13628,N_13544);
or U14359 (N_14359,N_13558,N_13930);
nor U14360 (N_14360,N_13614,N_13858);
nor U14361 (N_14361,N_13776,N_13949);
xnor U14362 (N_14362,N_13951,N_14242);
and U14363 (N_14363,N_14049,N_13571);
nand U14364 (N_14364,N_14234,N_13836);
and U14365 (N_14365,N_13777,N_14139);
nor U14366 (N_14366,N_13507,N_14073);
nor U14367 (N_14367,N_14215,N_14208);
or U14368 (N_14368,N_13542,N_14106);
or U14369 (N_14369,N_14031,N_13659);
nand U14370 (N_14370,N_14236,N_14064);
nor U14371 (N_14371,N_14046,N_14047);
and U14372 (N_14372,N_13637,N_13760);
nand U14373 (N_14373,N_13539,N_14134);
or U14374 (N_14374,N_13643,N_13778);
nand U14375 (N_14375,N_13955,N_13864);
or U14376 (N_14376,N_13806,N_14110);
nand U14377 (N_14377,N_13981,N_14008);
or U14378 (N_14378,N_13671,N_13640);
nor U14379 (N_14379,N_14138,N_13717);
nor U14380 (N_14380,N_13932,N_14082);
nor U14381 (N_14381,N_13967,N_13706);
and U14382 (N_14382,N_13991,N_13543);
nor U14383 (N_14383,N_13622,N_13748);
and U14384 (N_14384,N_13804,N_13572);
xnor U14385 (N_14385,N_13945,N_13866);
or U14386 (N_14386,N_13709,N_13732);
nand U14387 (N_14387,N_13687,N_14052);
xor U14388 (N_14388,N_13916,N_14048);
nor U14389 (N_14389,N_14107,N_13625);
and U14390 (N_14390,N_14026,N_14194);
xnor U14391 (N_14391,N_14198,N_13895);
or U14392 (N_14392,N_14193,N_14016);
and U14393 (N_14393,N_14053,N_13581);
nor U14394 (N_14394,N_13678,N_13905);
nor U14395 (N_14395,N_14172,N_13846);
or U14396 (N_14396,N_13984,N_13860);
or U14397 (N_14397,N_14054,N_13950);
and U14398 (N_14398,N_13873,N_13646);
nand U14399 (N_14399,N_14224,N_13840);
or U14400 (N_14400,N_14141,N_13697);
and U14401 (N_14401,N_13551,N_13626);
nand U14402 (N_14402,N_13893,N_13791);
or U14403 (N_14403,N_14029,N_13982);
nor U14404 (N_14404,N_14144,N_14101);
nor U14405 (N_14405,N_14212,N_13816);
nor U14406 (N_14406,N_14133,N_13647);
nand U14407 (N_14407,N_13645,N_13676);
nor U14408 (N_14408,N_13713,N_13546);
nand U14409 (N_14409,N_13933,N_13969);
nand U14410 (N_14410,N_13894,N_13923);
and U14411 (N_14411,N_13710,N_13517);
nor U14412 (N_14412,N_13767,N_13780);
and U14413 (N_14413,N_14081,N_13513);
and U14414 (N_14414,N_13977,N_14004);
or U14415 (N_14415,N_13857,N_14038);
nand U14416 (N_14416,N_13867,N_13747);
or U14417 (N_14417,N_13814,N_13934);
nor U14418 (N_14418,N_13520,N_14066);
and U14419 (N_14419,N_13537,N_14083);
nand U14420 (N_14420,N_14197,N_14168);
nand U14421 (N_14421,N_14057,N_13774);
nand U14422 (N_14422,N_14103,N_13759);
and U14423 (N_14423,N_13781,N_14127);
nor U14424 (N_14424,N_13674,N_14018);
or U14425 (N_14425,N_14007,N_14160);
xnor U14426 (N_14426,N_13586,N_13909);
nand U14427 (N_14427,N_13527,N_13535);
nand U14428 (N_14428,N_14156,N_13908);
nor U14429 (N_14429,N_14201,N_13604);
nor U14430 (N_14430,N_14164,N_14230);
or U14431 (N_14431,N_14161,N_13515);
nor U14432 (N_14432,N_13595,N_13810);
nor U14433 (N_14433,N_14091,N_13570);
or U14434 (N_14434,N_13502,N_13738);
nor U14435 (N_14435,N_14068,N_13599);
or U14436 (N_14436,N_13529,N_14122);
or U14437 (N_14437,N_13642,N_14035);
and U14438 (N_14438,N_13538,N_14015);
nor U14439 (N_14439,N_14182,N_13834);
and U14440 (N_14440,N_13591,N_13730);
nor U14441 (N_14441,N_14163,N_13763);
and U14442 (N_14442,N_14170,N_13993);
nor U14443 (N_14443,N_14185,N_13741);
and U14444 (N_14444,N_13519,N_13728);
and U14445 (N_14445,N_13651,N_13801);
nor U14446 (N_14446,N_13516,N_14214);
nor U14447 (N_14447,N_14196,N_13510);
or U14448 (N_14448,N_14243,N_14210);
or U14449 (N_14449,N_13828,N_13850);
nand U14450 (N_14450,N_13662,N_13584);
nand U14451 (N_14451,N_13534,N_14003);
or U14452 (N_14452,N_13569,N_14032);
nand U14453 (N_14453,N_13648,N_13634);
nand U14454 (N_14454,N_13987,N_13880);
nand U14455 (N_14455,N_14247,N_13530);
nor U14456 (N_14456,N_13632,N_14219);
or U14457 (N_14457,N_13772,N_13972);
and U14458 (N_14458,N_13797,N_13575);
and U14459 (N_14459,N_13862,N_13509);
or U14460 (N_14460,N_13941,N_14041);
nor U14461 (N_14461,N_13506,N_14249);
nor U14462 (N_14462,N_13970,N_13639);
nand U14463 (N_14463,N_13996,N_14162);
and U14464 (N_14464,N_14179,N_13592);
and U14465 (N_14465,N_13605,N_13587);
xor U14466 (N_14466,N_13619,N_13755);
or U14467 (N_14467,N_13715,N_13705);
and U14468 (N_14468,N_13620,N_13700);
or U14469 (N_14469,N_14002,N_13957);
nand U14470 (N_14470,N_13500,N_13784);
or U14471 (N_14471,N_13742,N_14093);
nor U14472 (N_14472,N_13839,N_13903);
and U14473 (N_14473,N_14129,N_13578);
nand U14474 (N_14474,N_13820,N_14061);
nand U14475 (N_14475,N_13769,N_13607);
and U14476 (N_14476,N_13565,N_13885);
nor U14477 (N_14477,N_13847,N_14096);
nand U14478 (N_14478,N_13803,N_14218);
or U14479 (N_14479,N_13819,N_13960);
and U14480 (N_14480,N_14180,N_14241);
nand U14481 (N_14481,N_14213,N_13910);
and U14482 (N_14482,N_13554,N_13964);
nor U14483 (N_14483,N_13729,N_13925);
or U14484 (N_14484,N_13998,N_13561);
nand U14485 (N_14485,N_14033,N_14153);
nand U14486 (N_14486,N_13567,N_13859);
nand U14487 (N_14487,N_14155,N_13603);
or U14488 (N_14488,N_13978,N_14183);
or U14489 (N_14489,N_13765,N_13694);
or U14490 (N_14490,N_13911,N_13654);
nand U14491 (N_14491,N_14005,N_13966);
and U14492 (N_14492,N_13853,N_13727);
or U14493 (N_14493,N_14011,N_14169);
nor U14494 (N_14494,N_14022,N_13899);
nor U14495 (N_14495,N_13670,N_13568);
or U14496 (N_14496,N_13744,N_13869);
nand U14497 (N_14497,N_14078,N_13508);
nor U14498 (N_14498,N_14147,N_14117);
nor U14499 (N_14499,N_14216,N_14228);
or U14500 (N_14500,N_14076,N_13734);
or U14501 (N_14501,N_13827,N_13875);
or U14502 (N_14502,N_14019,N_13794);
or U14503 (N_14503,N_13779,N_14090);
nor U14504 (N_14504,N_13582,N_14118);
nor U14505 (N_14505,N_13788,N_13733);
nand U14506 (N_14506,N_13621,N_13989);
or U14507 (N_14507,N_14246,N_14023);
and U14508 (N_14508,N_13817,N_13974);
nand U14509 (N_14509,N_13901,N_13675);
and U14510 (N_14510,N_13997,N_13689);
nor U14511 (N_14511,N_13714,N_14165);
nor U14512 (N_14512,N_13927,N_13881);
and U14513 (N_14513,N_13655,N_13948);
nand U14514 (N_14514,N_14154,N_13684);
nor U14515 (N_14515,N_14119,N_14191);
or U14516 (N_14516,N_14237,N_13889);
nand U14517 (N_14517,N_13855,N_13940);
or U14518 (N_14518,N_13716,N_14220);
or U14519 (N_14519,N_13830,N_13835);
xnor U14520 (N_14520,N_13682,N_13635);
and U14521 (N_14521,N_14167,N_14229);
or U14522 (N_14522,N_13579,N_13685);
nor U14523 (N_14523,N_13986,N_14012);
and U14524 (N_14524,N_13528,N_14060);
and U14525 (N_14525,N_13679,N_13811);
nor U14526 (N_14526,N_13861,N_13617);
or U14527 (N_14527,N_14158,N_13707);
and U14528 (N_14528,N_13650,N_13616);
nor U14529 (N_14529,N_14159,N_14217);
or U14530 (N_14530,N_14206,N_13735);
and U14531 (N_14531,N_13514,N_13536);
nand U14532 (N_14532,N_14115,N_13701);
nand U14533 (N_14533,N_14137,N_14202);
or U14534 (N_14534,N_13629,N_13601);
and U14535 (N_14535,N_13704,N_14173);
nand U14536 (N_14536,N_13644,N_14014);
nand U14537 (N_14537,N_14094,N_13708);
nor U14538 (N_14538,N_14044,N_14157);
nor U14539 (N_14539,N_14121,N_13597);
nor U14540 (N_14540,N_13630,N_13983);
and U14541 (N_14541,N_14020,N_14050);
or U14542 (N_14542,N_13818,N_14177);
and U14543 (N_14543,N_13929,N_13973);
and U14544 (N_14544,N_14084,N_13841);
and U14545 (N_14545,N_14190,N_13883);
nor U14546 (N_14546,N_13959,N_14098);
or U14547 (N_14547,N_13683,N_13766);
nor U14548 (N_14548,N_13872,N_13660);
nor U14549 (N_14549,N_14027,N_13593);
nand U14550 (N_14550,N_13771,N_13798);
nand U14551 (N_14551,N_14059,N_14225);
and U14552 (N_14552,N_13813,N_13764);
nor U14553 (N_14553,N_13611,N_13775);
and U14554 (N_14554,N_14116,N_13541);
nor U14555 (N_14555,N_13724,N_13824);
or U14556 (N_14556,N_13532,N_13610);
or U14557 (N_14557,N_14125,N_13887);
nand U14558 (N_14558,N_14040,N_13898);
and U14559 (N_14559,N_14075,N_13552);
nor U14560 (N_14560,N_13698,N_13843);
nor U14561 (N_14561,N_13526,N_14111);
nand U14562 (N_14562,N_14036,N_13907);
nand U14563 (N_14563,N_14171,N_13812);
and U14564 (N_14564,N_14151,N_13968);
and U14565 (N_14565,N_14043,N_13985);
nor U14566 (N_14566,N_14192,N_14010);
or U14567 (N_14567,N_13877,N_13703);
nor U14568 (N_14568,N_14200,N_13615);
and U14569 (N_14569,N_14112,N_14042);
nor U14570 (N_14570,N_14186,N_13545);
or U14571 (N_14571,N_13979,N_13912);
nand U14572 (N_14572,N_13936,N_13770);
nor U14573 (N_14573,N_13773,N_13588);
or U14574 (N_14574,N_14135,N_14000);
and U14575 (N_14575,N_13802,N_13751);
nand U14576 (N_14576,N_13882,N_14124);
or U14577 (N_14577,N_13501,N_14205);
nor U14578 (N_14578,N_13726,N_14130);
nor U14579 (N_14579,N_13723,N_14087);
nand U14580 (N_14580,N_13566,N_13849);
or U14581 (N_14581,N_14174,N_14240);
and U14582 (N_14582,N_13743,N_13919);
nand U14583 (N_14583,N_14226,N_13825);
and U14584 (N_14584,N_13722,N_14176);
or U14585 (N_14585,N_13870,N_13562);
or U14586 (N_14586,N_13837,N_13988);
or U14587 (N_14587,N_13999,N_13884);
and U14588 (N_14588,N_14131,N_13576);
nor U14589 (N_14589,N_13711,N_13937);
nor U14590 (N_14590,N_13952,N_13954);
nand U14591 (N_14591,N_14140,N_13920);
and U14592 (N_14592,N_14108,N_13667);
nand U14593 (N_14593,N_13971,N_13596);
and U14594 (N_14594,N_13547,N_13879);
and U14595 (N_14595,N_13740,N_13549);
nand U14596 (N_14596,N_13602,N_14065);
nand U14597 (N_14597,N_13906,N_13652);
nor U14598 (N_14598,N_14239,N_14207);
and U14599 (N_14599,N_14195,N_13976);
nand U14600 (N_14600,N_14233,N_13928);
or U14601 (N_14601,N_14079,N_14100);
nor U14602 (N_14602,N_13805,N_14244);
nor U14603 (N_14603,N_14039,N_13807);
and U14604 (N_14604,N_13992,N_13786);
and U14605 (N_14605,N_14203,N_13523);
nand U14606 (N_14606,N_14034,N_13756);
or U14607 (N_14607,N_13550,N_14095);
or U14608 (N_14608,N_13938,N_13548);
nor U14609 (N_14609,N_13580,N_13995);
or U14610 (N_14610,N_13888,N_13815);
and U14611 (N_14611,N_14123,N_13822);
nand U14612 (N_14612,N_13915,N_13761);
nand U14613 (N_14613,N_14181,N_13720);
nor U14614 (N_14614,N_13842,N_13821);
nand U14615 (N_14615,N_13657,N_14245);
nor U14616 (N_14616,N_13664,N_13589);
and U14617 (N_14617,N_14187,N_14104);
nor U14618 (N_14618,N_13829,N_14232);
and U14619 (N_14619,N_13653,N_13800);
or U14620 (N_14620,N_13688,N_13719);
or U14621 (N_14621,N_13511,N_14051);
or U14622 (N_14622,N_13946,N_13947);
and U14623 (N_14623,N_13556,N_13943);
and U14624 (N_14624,N_13699,N_13874);
and U14625 (N_14625,N_13940,N_13794);
or U14626 (N_14626,N_14055,N_13663);
nand U14627 (N_14627,N_13721,N_13785);
and U14628 (N_14628,N_13620,N_13893);
nor U14629 (N_14629,N_14123,N_14170);
or U14630 (N_14630,N_14199,N_13509);
or U14631 (N_14631,N_13842,N_13869);
nand U14632 (N_14632,N_14163,N_13575);
nor U14633 (N_14633,N_14089,N_14152);
nand U14634 (N_14634,N_13948,N_13723);
nor U14635 (N_14635,N_14224,N_14014);
nand U14636 (N_14636,N_14173,N_13607);
nand U14637 (N_14637,N_13887,N_14030);
nor U14638 (N_14638,N_14162,N_14098);
nand U14639 (N_14639,N_14012,N_13514);
or U14640 (N_14640,N_13550,N_14038);
and U14641 (N_14641,N_14209,N_14179);
nor U14642 (N_14642,N_14209,N_14022);
nor U14643 (N_14643,N_14067,N_13520);
nor U14644 (N_14644,N_13978,N_14126);
nand U14645 (N_14645,N_13670,N_14137);
nor U14646 (N_14646,N_13652,N_14110);
nand U14647 (N_14647,N_13903,N_13702);
nor U14648 (N_14648,N_13816,N_13813);
or U14649 (N_14649,N_13588,N_13561);
or U14650 (N_14650,N_13809,N_13516);
or U14651 (N_14651,N_13655,N_13536);
nor U14652 (N_14652,N_14115,N_14112);
nor U14653 (N_14653,N_14155,N_14223);
nor U14654 (N_14654,N_13902,N_13762);
or U14655 (N_14655,N_13586,N_13977);
or U14656 (N_14656,N_13527,N_14225);
nand U14657 (N_14657,N_13820,N_13875);
nand U14658 (N_14658,N_13953,N_13631);
nor U14659 (N_14659,N_13705,N_13538);
nor U14660 (N_14660,N_13745,N_13872);
or U14661 (N_14661,N_13794,N_13950);
nor U14662 (N_14662,N_14215,N_13732);
nand U14663 (N_14663,N_13927,N_14031);
or U14664 (N_14664,N_13797,N_13588);
and U14665 (N_14665,N_14087,N_14118);
nor U14666 (N_14666,N_13634,N_13876);
nor U14667 (N_14667,N_13901,N_13811);
and U14668 (N_14668,N_14143,N_14183);
nand U14669 (N_14669,N_14214,N_14195);
or U14670 (N_14670,N_13717,N_14037);
and U14671 (N_14671,N_13716,N_13622);
and U14672 (N_14672,N_14116,N_13547);
or U14673 (N_14673,N_13654,N_13961);
and U14674 (N_14674,N_13875,N_13688);
nand U14675 (N_14675,N_13513,N_13545);
nand U14676 (N_14676,N_13865,N_13957);
and U14677 (N_14677,N_13568,N_14051);
nor U14678 (N_14678,N_14051,N_13925);
or U14679 (N_14679,N_14224,N_13954);
nand U14680 (N_14680,N_14107,N_14171);
nand U14681 (N_14681,N_13928,N_13560);
and U14682 (N_14682,N_13631,N_13883);
nand U14683 (N_14683,N_13839,N_14192);
nand U14684 (N_14684,N_13726,N_14117);
nand U14685 (N_14685,N_13759,N_13515);
nand U14686 (N_14686,N_14085,N_13622);
nor U14687 (N_14687,N_13815,N_13507);
nand U14688 (N_14688,N_13540,N_13573);
and U14689 (N_14689,N_13638,N_14120);
nor U14690 (N_14690,N_13993,N_13855);
nand U14691 (N_14691,N_13950,N_13865);
nor U14692 (N_14692,N_14123,N_14060);
nor U14693 (N_14693,N_13764,N_14019);
nor U14694 (N_14694,N_13706,N_14123);
or U14695 (N_14695,N_13943,N_14188);
nor U14696 (N_14696,N_14094,N_13771);
and U14697 (N_14697,N_13566,N_13721);
nor U14698 (N_14698,N_13878,N_13923);
nor U14699 (N_14699,N_13939,N_14143);
and U14700 (N_14700,N_13711,N_14006);
and U14701 (N_14701,N_13649,N_14081);
or U14702 (N_14702,N_14175,N_13851);
nand U14703 (N_14703,N_13893,N_14240);
or U14704 (N_14704,N_13548,N_14112);
nor U14705 (N_14705,N_13507,N_13724);
and U14706 (N_14706,N_13557,N_13861);
nand U14707 (N_14707,N_14177,N_13694);
nand U14708 (N_14708,N_13996,N_13991);
or U14709 (N_14709,N_14209,N_14110);
and U14710 (N_14710,N_14024,N_13929);
and U14711 (N_14711,N_14050,N_13902);
xnor U14712 (N_14712,N_14144,N_14021);
and U14713 (N_14713,N_13958,N_13505);
or U14714 (N_14714,N_13961,N_14114);
nand U14715 (N_14715,N_13980,N_13814);
nand U14716 (N_14716,N_14247,N_13962);
nor U14717 (N_14717,N_13934,N_13563);
nand U14718 (N_14718,N_13747,N_13713);
or U14719 (N_14719,N_13947,N_13973);
or U14720 (N_14720,N_13985,N_13697);
xor U14721 (N_14721,N_13634,N_14059);
nor U14722 (N_14722,N_13705,N_14065);
or U14723 (N_14723,N_14130,N_14206);
xnor U14724 (N_14724,N_14193,N_14126);
and U14725 (N_14725,N_13710,N_13620);
and U14726 (N_14726,N_13796,N_14139);
nor U14727 (N_14727,N_13909,N_13792);
nor U14728 (N_14728,N_13683,N_13609);
nand U14729 (N_14729,N_13635,N_13960);
nor U14730 (N_14730,N_13870,N_13753);
or U14731 (N_14731,N_13957,N_13525);
and U14732 (N_14732,N_13691,N_13877);
nand U14733 (N_14733,N_13992,N_13868);
and U14734 (N_14734,N_14078,N_14011);
nor U14735 (N_14735,N_14150,N_13749);
nor U14736 (N_14736,N_14135,N_14085);
or U14737 (N_14737,N_13663,N_13828);
nand U14738 (N_14738,N_13691,N_14009);
and U14739 (N_14739,N_13576,N_13824);
and U14740 (N_14740,N_13779,N_13959);
nor U14741 (N_14741,N_13639,N_14212);
and U14742 (N_14742,N_13597,N_14211);
nor U14743 (N_14743,N_14105,N_13791);
or U14744 (N_14744,N_14157,N_14245);
nor U14745 (N_14745,N_14110,N_13923);
or U14746 (N_14746,N_14016,N_13972);
nand U14747 (N_14747,N_14234,N_14218);
or U14748 (N_14748,N_13609,N_13617);
and U14749 (N_14749,N_13684,N_13882);
and U14750 (N_14750,N_14196,N_13766);
or U14751 (N_14751,N_13906,N_14030);
or U14752 (N_14752,N_14043,N_14068);
and U14753 (N_14753,N_13613,N_13782);
nand U14754 (N_14754,N_13889,N_13657);
or U14755 (N_14755,N_14198,N_13619);
and U14756 (N_14756,N_13513,N_13717);
and U14757 (N_14757,N_14184,N_13886);
nor U14758 (N_14758,N_13894,N_14137);
nor U14759 (N_14759,N_13999,N_13777);
and U14760 (N_14760,N_13848,N_14198);
nor U14761 (N_14761,N_14037,N_13747);
nand U14762 (N_14762,N_13640,N_14171);
nand U14763 (N_14763,N_13876,N_13894);
or U14764 (N_14764,N_13953,N_14047);
or U14765 (N_14765,N_14135,N_14032);
nor U14766 (N_14766,N_13611,N_14130);
nand U14767 (N_14767,N_13846,N_13709);
or U14768 (N_14768,N_13516,N_13595);
and U14769 (N_14769,N_14234,N_13676);
and U14770 (N_14770,N_14057,N_13765);
and U14771 (N_14771,N_13634,N_13595);
or U14772 (N_14772,N_13755,N_14176);
or U14773 (N_14773,N_13557,N_13791);
nand U14774 (N_14774,N_13989,N_13988);
and U14775 (N_14775,N_13506,N_13736);
nor U14776 (N_14776,N_14138,N_13798);
nand U14777 (N_14777,N_13504,N_14151);
nor U14778 (N_14778,N_14144,N_13785);
and U14779 (N_14779,N_13504,N_14088);
nor U14780 (N_14780,N_13967,N_13732);
and U14781 (N_14781,N_13878,N_13693);
or U14782 (N_14782,N_13858,N_14111);
nand U14783 (N_14783,N_13923,N_13505);
nand U14784 (N_14784,N_13914,N_14190);
and U14785 (N_14785,N_13647,N_13510);
and U14786 (N_14786,N_13843,N_14100);
nor U14787 (N_14787,N_13994,N_13738);
nor U14788 (N_14788,N_13932,N_13729);
nor U14789 (N_14789,N_14137,N_14175);
nand U14790 (N_14790,N_14100,N_13571);
or U14791 (N_14791,N_14173,N_13527);
or U14792 (N_14792,N_14241,N_13736);
and U14793 (N_14793,N_13948,N_13695);
nor U14794 (N_14794,N_13909,N_13847);
nor U14795 (N_14795,N_14135,N_13613);
nand U14796 (N_14796,N_13932,N_13686);
nand U14797 (N_14797,N_14184,N_14230);
and U14798 (N_14798,N_13899,N_13932);
nor U14799 (N_14799,N_13937,N_13586);
or U14800 (N_14800,N_13533,N_13513);
nand U14801 (N_14801,N_13958,N_14166);
or U14802 (N_14802,N_13944,N_13914);
or U14803 (N_14803,N_14121,N_13525);
and U14804 (N_14804,N_13881,N_13905);
or U14805 (N_14805,N_13998,N_14164);
and U14806 (N_14806,N_14217,N_13933);
nand U14807 (N_14807,N_13936,N_14105);
and U14808 (N_14808,N_14243,N_13930);
or U14809 (N_14809,N_14202,N_13501);
nor U14810 (N_14810,N_13598,N_13737);
and U14811 (N_14811,N_13513,N_14227);
or U14812 (N_14812,N_14191,N_14220);
nor U14813 (N_14813,N_13567,N_14123);
and U14814 (N_14814,N_14054,N_13887);
nand U14815 (N_14815,N_13974,N_13602);
and U14816 (N_14816,N_13724,N_14043);
or U14817 (N_14817,N_14162,N_13603);
nand U14818 (N_14818,N_13815,N_13513);
and U14819 (N_14819,N_14188,N_13815);
nand U14820 (N_14820,N_14092,N_13956);
nand U14821 (N_14821,N_14120,N_13632);
and U14822 (N_14822,N_14189,N_13590);
and U14823 (N_14823,N_14072,N_14235);
and U14824 (N_14824,N_14020,N_13507);
nand U14825 (N_14825,N_14062,N_13596);
or U14826 (N_14826,N_13542,N_13976);
or U14827 (N_14827,N_14134,N_13589);
or U14828 (N_14828,N_14192,N_14070);
or U14829 (N_14829,N_13608,N_13651);
nand U14830 (N_14830,N_13953,N_13573);
nor U14831 (N_14831,N_13711,N_14204);
nor U14832 (N_14832,N_13731,N_13799);
nand U14833 (N_14833,N_13675,N_14013);
nor U14834 (N_14834,N_14246,N_14071);
or U14835 (N_14835,N_13669,N_13915);
nand U14836 (N_14836,N_13917,N_14002);
nand U14837 (N_14837,N_13946,N_13612);
nand U14838 (N_14838,N_13530,N_13525);
or U14839 (N_14839,N_14095,N_13735);
nor U14840 (N_14840,N_13680,N_13919);
nand U14841 (N_14841,N_13799,N_14135);
and U14842 (N_14842,N_14030,N_13650);
or U14843 (N_14843,N_13678,N_13651);
or U14844 (N_14844,N_13522,N_13672);
nor U14845 (N_14845,N_13613,N_13691);
nand U14846 (N_14846,N_13557,N_13945);
and U14847 (N_14847,N_13981,N_13757);
or U14848 (N_14848,N_13790,N_13682);
or U14849 (N_14849,N_14117,N_14013);
or U14850 (N_14850,N_13500,N_13869);
nand U14851 (N_14851,N_14124,N_13956);
or U14852 (N_14852,N_13762,N_14083);
or U14853 (N_14853,N_13577,N_14134);
nand U14854 (N_14854,N_13565,N_13666);
and U14855 (N_14855,N_14137,N_13905);
and U14856 (N_14856,N_14057,N_13860);
and U14857 (N_14857,N_13680,N_13803);
nor U14858 (N_14858,N_13619,N_14078);
nor U14859 (N_14859,N_14006,N_14012);
and U14860 (N_14860,N_13795,N_13887);
and U14861 (N_14861,N_13950,N_13540);
or U14862 (N_14862,N_13517,N_14059);
or U14863 (N_14863,N_14214,N_13629);
or U14864 (N_14864,N_13547,N_13962);
nand U14865 (N_14865,N_13728,N_13975);
nand U14866 (N_14866,N_13582,N_13574);
or U14867 (N_14867,N_13713,N_13719);
or U14868 (N_14868,N_13798,N_14220);
or U14869 (N_14869,N_13521,N_14185);
or U14870 (N_14870,N_13679,N_14104);
nand U14871 (N_14871,N_13892,N_14133);
or U14872 (N_14872,N_13790,N_13611);
nor U14873 (N_14873,N_14234,N_14080);
and U14874 (N_14874,N_13807,N_14129);
or U14875 (N_14875,N_14017,N_13851);
nor U14876 (N_14876,N_13789,N_13928);
or U14877 (N_14877,N_13785,N_13812);
nor U14878 (N_14878,N_13976,N_14185);
or U14879 (N_14879,N_13817,N_14098);
nor U14880 (N_14880,N_13853,N_13947);
nand U14881 (N_14881,N_13524,N_14236);
and U14882 (N_14882,N_13569,N_14212);
xnor U14883 (N_14883,N_13670,N_13697);
or U14884 (N_14884,N_13748,N_13758);
or U14885 (N_14885,N_13716,N_13571);
nand U14886 (N_14886,N_14095,N_14033);
or U14887 (N_14887,N_13854,N_13892);
nand U14888 (N_14888,N_13810,N_14028);
and U14889 (N_14889,N_14123,N_13613);
and U14890 (N_14890,N_13962,N_14006);
nor U14891 (N_14891,N_13870,N_14020);
and U14892 (N_14892,N_13614,N_14068);
nor U14893 (N_14893,N_13531,N_13724);
nand U14894 (N_14894,N_13665,N_13934);
and U14895 (N_14895,N_13927,N_13838);
or U14896 (N_14896,N_13689,N_13595);
or U14897 (N_14897,N_14205,N_13500);
and U14898 (N_14898,N_13731,N_13738);
and U14899 (N_14899,N_13575,N_13800);
nand U14900 (N_14900,N_14225,N_13832);
nor U14901 (N_14901,N_13655,N_14019);
or U14902 (N_14902,N_13968,N_13628);
nor U14903 (N_14903,N_14136,N_13837);
nand U14904 (N_14904,N_13582,N_14007);
or U14905 (N_14905,N_13982,N_14089);
and U14906 (N_14906,N_13929,N_13945);
or U14907 (N_14907,N_13578,N_13506);
and U14908 (N_14908,N_14040,N_14058);
and U14909 (N_14909,N_13744,N_13509);
and U14910 (N_14910,N_13577,N_14170);
or U14911 (N_14911,N_13524,N_13720);
or U14912 (N_14912,N_13838,N_13846);
nand U14913 (N_14913,N_14039,N_13826);
or U14914 (N_14914,N_13577,N_13582);
nand U14915 (N_14915,N_13929,N_13665);
and U14916 (N_14916,N_13946,N_13941);
nor U14917 (N_14917,N_14221,N_13844);
or U14918 (N_14918,N_13977,N_13974);
or U14919 (N_14919,N_14001,N_13865);
or U14920 (N_14920,N_14184,N_13538);
and U14921 (N_14921,N_14136,N_13877);
and U14922 (N_14922,N_14114,N_14021);
and U14923 (N_14923,N_13846,N_14012);
nand U14924 (N_14924,N_13656,N_14054);
nor U14925 (N_14925,N_14106,N_14035);
or U14926 (N_14926,N_13729,N_13515);
nor U14927 (N_14927,N_13773,N_14026);
nor U14928 (N_14928,N_14174,N_13850);
nor U14929 (N_14929,N_13972,N_13544);
or U14930 (N_14930,N_13638,N_13504);
nand U14931 (N_14931,N_14035,N_13794);
or U14932 (N_14932,N_14115,N_13636);
nor U14933 (N_14933,N_13839,N_13694);
and U14934 (N_14934,N_14194,N_13882);
or U14935 (N_14935,N_14232,N_13879);
nand U14936 (N_14936,N_13623,N_14094);
nand U14937 (N_14937,N_13942,N_13571);
or U14938 (N_14938,N_14218,N_14150);
nand U14939 (N_14939,N_13536,N_13904);
and U14940 (N_14940,N_13903,N_13619);
nor U14941 (N_14941,N_14121,N_14207);
or U14942 (N_14942,N_13736,N_13694);
nor U14943 (N_14943,N_13890,N_14067);
or U14944 (N_14944,N_13684,N_14150);
and U14945 (N_14945,N_13718,N_13507);
nor U14946 (N_14946,N_14028,N_14135);
nand U14947 (N_14947,N_13838,N_13533);
xnor U14948 (N_14948,N_14188,N_14175);
and U14949 (N_14949,N_14175,N_13543);
and U14950 (N_14950,N_13776,N_14144);
or U14951 (N_14951,N_14079,N_13890);
xnor U14952 (N_14952,N_13802,N_13651);
or U14953 (N_14953,N_14018,N_14102);
nand U14954 (N_14954,N_13594,N_14208);
nor U14955 (N_14955,N_14048,N_14233);
xor U14956 (N_14956,N_13654,N_14191);
or U14957 (N_14957,N_14155,N_13703);
nor U14958 (N_14958,N_13907,N_14205);
or U14959 (N_14959,N_14237,N_13707);
nor U14960 (N_14960,N_14089,N_14181);
nor U14961 (N_14961,N_14239,N_13747);
nor U14962 (N_14962,N_13573,N_14188);
or U14963 (N_14963,N_13543,N_13856);
nand U14964 (N_14964,N_13740,N_14076);
or U14965 (N_14965,N_13831,N_13549);
nand U14966 (N_14966,N_13594,N_13855);
or U14967 (N_14967,N_13776,N_13920);
or U14968 (N_14968,N_13521,N_13827);
nor U14969 (N_14969,N_13705,N_14077);
and U14970 (N_14970,N_13726,N_14119);
and U14971 (N_14971,N_13906,N_13677);
or U14972 (N_14972,N_14249,N_13775);
nor U14973 (N_14973,N_13516,N_14194);
or U14974 (N_14974,N_13748,N_14128);
nor U14975 (N_14975,N_13526,N_13659);
nand U14976 (N_14976,N_13712,N_13789);
or U14977 (N_14977,N_13603,N_13975);
nor U14978 (N_14978,N_13987,N_13528);
nand U14979 (N_14979,N_14138,N_13805);
nand U14980 (N_14980,N_13625,N_13984);
or U14981 (N_14981,N_13736,N_13992);
or U14982 (N_14982,N_13653,N_13923);
nand U14983 (N_14983,N_13659,N_13709);
and U14984 (N_14984,N_13988,N_13907);
or U14985 (N_14985,N_13813,N_13918);
nor U14986 (N_14986,N_13882,N_13678);
and U14987 (N_14987,N_14004,N_13801);
and U14988 (N_14988,N_13844,N_13605);
nor U14989 (N_14989,N_14026,N_13864);
and U14990 (N_14990,N_13739,N_13651);
nand U14991 (N_14991,N_13541,N_14132);
nand U14992 (N_14992,N_13720,N_13814);
nand U14993 (N_14993,N_13785,N_14030);
nor U14994 (N_14994,N_13659,N_13865);
or U14995 (N_14995,N_14049,N_13923);
and U14996 (N_14996,N_14086,N_14077);
nor U14997 (N_14997,N_14017,N_13570);
and U14998 (N_14998,N_14068,N_14086);
nor U14999 (N_14999,N_14145,N_14009);
nor UO_0 (O_0,N_14679,N_14335);
and UO_1 (O_1,N_14776,N_14361);
nor UO_2 (O_2,N_14357,N_14408);
nand UO_3 (O_3,N_14797,N_14689);
nor UO_4 (O_4,N_14559,N_14629);
or UO_5 (O_5,N_14294,N_14342);
or UO_6 (O_6,N_14626,N_14803);
or UO_7 (O_7,N_14817,N_14707);
nor UO_8 (O_8,N_14321,N_14724);
nor UO_9 (O_9,N_14719,N_14251);
and UO_10 (O_10,N_14762,N_14270);
or UO_11 (O_11,N_14372,N_14483);
nor UO_12 (O_12,N_14538,N_14594);
nor UO_13 (O_13,N_14250,N_14819);
nand UO_14 (O_14,N_14501,N_14863);
and UO_15 (O_15,N_14539,N_14926);
or UO_16 (O_16,N_14288,N_14944);
and UO_17 (O_17,N_14692,N_14468);
nor UO_18 (O_18,N_14605,N_14971);
nand UO_19 (O_19,N_14578,N_14826);
nor UO_20 (O_20,N_14535,N_14607);
nand UO_21 (O_21,N_14814,N_14945);
or UO_22 (O_22,N_14507,N_14347);
or UO_23 (O_23,N_14889,N_14955);
nor UO_24 (O_24,N_14767,N_14477);
or UO_25 (O_25,N_14406,N_14654);
or UO_26 (O_26,N_14359,N_14916);
and UO_27 (O_27,N_14484,N_14741);
nand UO_28 (O_28,N_14424,N_14365);
or UO_29 (O_29,N_14515,N_14287);
and UO_30 (O_30,N_14274,N_14792);
or UO_31 (O_31,N_14779,N_14986);
nor UO_32 (O_32,N_14476,N_14950);
or UO_33 (O_33,N_14447,N_14960);
nand UO_34 (O_34,N_14352,N_14329);
or UO_35 (O_35,N_14835,N_14290);
and UO_36 (O_36,N_14513,N_14465);
or UO_37 (O_37,N_14269,N_14573);
nand UO_38 (O_38,N_14624,N_14920);
and UO_39 (O_39,N_14580,N_14587);
nand UO_40 (O_40,N_14557,N_14475);
or UO_41 (O_41,N_14646,N_14543);
and UO_42 (O_42,N_14678,N_14600);
and UO_43 (O_43,N_14804,N_14421);
nor UO_44 (O_44,N_14256,N_14518);
and UO_45 (O_45,N_14997,N_14768);
and UO_46 (O_46,N_14610,N_14387);
or UO_47 (O_47,N_14621,N_14892);
and UO_48 (O_48,N_14490,N_14497);
nor UO_49 (O_49,N_14729,N_14571);
or UO_50 (O_50,N_14656,N_14973);
nor UO_51 (O_51,N_14591,N_14749);
or UO_52 (O_52,N_14635,N_14579);
nand UO_53 (O_53,N_14902,N_14806);
and UO_54 (O_54,N_14853,N_14907);
nand UO_55 (O_55,N_14681,N_14422);
xnor UO_56 (O_56,N_14284,N_14851);
nor UO_57 (O_57,N_14978,N_14439);
nand UO_58 (O_58,N_14252,N_14348);
nor UO_59 (O_59,N_14417,N_14377);
or UO_60 (O_60,N_14500,N_14487);
and UO_61 (O_61,N_14264,N_14954);
nor UO_62 (O_62,N_14878,N_14316);
nand UO_63 (O_63,N_14838,N_14530);
or UO_64 (O_64,N_14991,N_14868);
xor UO_65 (O_65,N_14470,N_14981);
nand UO_66 (O_66,N_14650,N_14875);
or UO_67 (O_67,N_14737,N_14313);
and UO_68 (O_68,N_14567,N_14930);
nand UO_69 (O_69,N_14998,N_14904);
nand UO_70 (O_70,N_14888,N_14731);
nand UO_71 (O_71,N_14636,N_14935);
and UO_72 (O_72,N_14818,N_14478);
and UO_73 (O_73,N_14325,N_14672);
nand UO_74 (O_74,N_14680,N_14469);
or UO_75 (O_75,N_14574,N_14642);
nand UO_76 (O_76,N_14534,N_14428);
nand UO_77 (O_77,N_14298,N_14932);
nand UO_78 (O_78,N_14569,N_14871);
nor UO_79 (O_79,N_14315,N_14379);
nor UO_80 (O_80,N_14402,N_14657);
and UO_81 (O_81,N_14625,N_14403);
or UO_82 (O_82,N_14346,N_14975);
or UO_83 (O_83,N_14989,N_14604);
nor UO_84 (O_84,N_14616,N_14738);
and UO_85 (O_85,N_14718,N_14485);
nor UO_86 (O_86,N_14582,N_14671);
nor UO_87 (O_87,N_14267,N_14339);
or UO_88 (O_88,N_14698,N_14524);
or UO_89 (O_89,N_14392,N_14992);
or UO_90 (O_90,N_14683,N_14963);
nor UO_91 (O_91,N_14669,N_14766);
and UO_92 (O_92,N_14383,N_14536);
nand UO_93 (O_93,N_14412,N_14602);
nor UO_94 (O_94,N_14714,N_14828);
or UO_95 (O_95,N_14541,N_14556);
nand UO_96 (O_96,N_14301,N_14299);
nand UO_97 (O_97,N_14854,N_14885);
or UO_98 (O_98,N_14957,N_14702);
nor UO_99 (O_99,N_14910,N_14293);
and UO_100 (O_100,N_14418,N_14364);
nor UO_101 (O_101,N_14940,N_14425);
or UO_102 (O_102,N_14805,N_14987);
and UO_103 (O_103,N_14744,N_14946);
or UO_104 (O_104,N_14612,N_14486);
nand UO_105 (O_105,N_14684,N_14967);
or UO_106 (O_106,N_14464,N_14782);
or UO_107 (O_107,N_14943,N_14503);
or UO_108 (O_108,N_14560,N_14708);
and UO_109 (O_109,N_14880,N_14929);
and UO_110 (O_110,N_14481,N_14864);
nand UO_111 (O_111,N_14493,N_14323);
and UO_112 (O_112,N_14699,N_14462);
nand UO_113 (O_113,N_14273,N_14385);
or UO_114 (O_114,N_14344,N_14925);
nand UO_115 (O_115,N_14908,N_14627);
or UO_116 (O_116,N_14791,N_14399);
and UO_117 (O_117,N_14471,N_14753);
or UO_118 (O_118,N_14407,N_14821);
or UO_119 (O_119,N_14865,N_14923);
or UO_120 (O_120,N_14965,N_14676);
nand UO_121 (O_121,N_14832,N_14409);
or UO_122 (O_122,N_14816,N_14453);
or UO_123 (O_123,N_14599,N_14354);
nand UO_124 (O_124,N_14834,N_14461);
and UO_125 (O_125,N_14746,N_14951);
nor UO_126 (O_126,N_14652,N_14972);
and UO_127 (O_127,N_14961,N_14688);
or UO_128 (O_128,N_14917,N_14317);
nand UO_129 (O_129,N_14262,N_14488);
nor UO_130 (O_130,N_14271,N_14905);
nand UO_131 (O_131,N_14445,N_14393);
or UO_132 (O_132,N_14673,N_14691);
and UO_133 (O_133,N_14455,N_14793);
nand UO_134 (O_134,N_14644,N_14886);
nand UO_135 (O_135,N_14995,N_14716);
and UO_136 (O_136,N_14894,N_14632);
and UO_137 (O_137,N_14494,N_14386);
and UO_138 (O_138,N_14953,N_14523);
nor UO_139 (O_139,N_14775,N_14537);
or UO_140 (O_140,N_14528,N_14341);
or UO_141 (O_141,N_14451,N_14748);
nor UO_142 (O_142,N_14585,N_14436);
nand UO_143 (O_143,N_14983,N_14275);
nor UO_144 (O_144,N_14979,N_14442);
or UO_145 (O_145,N_14457,N_14295);
nand UO_146 (O_146,N_14400,N_14913);
or UO_147 (O_147,N_14977,N_14253);
nor UO_148 (O_148,N_14686,N_14933);
and UO_149 (O_149,N_14473,N_14340);
or UO_150 (O_150,N_14328,N_14550);
nand UO_151 (O_151,N_14939,N_14314);
and UO_152 (O_152,N_14677,N_14291);
nor UO_153 (O_153,N_14405,N_14670);
nand UO_154 (O_154,N_14728,N_14467);
nand UO_155 (O_155,N_14261,N_14282);
nor UO_156 (O_156,N_14320,N_14414);
and UO_157 (O_157,N_14934,N_14896);
or UO_158 (O_158,N_14815,N_14463);
or UO_159 (O_159,N_14770,N_14480);
nor UO_160 (O_160,N_14773,N_14496);
nand UO_161 (O_161,N_14968,N_14527);
nor UO_162 (O_162,N_14549,N_14394);
nor UO_163 (O_163,N_14956,N_14586);
and UO_164 (O_164,N_14959,N_14350);
and UO_165 (O_165,N_14846,N_14659);
or UO_166 (O_166,N_14890,N_14787);
nor UO_167 (O_167,N_14371,N_14278);
nand UO_168 (O_168,N_14837,N_14564);
nor UO_169 (O_169,N_14649,N_14730);
nand UO_170 (O_170,N_14502,N_14300);
nand UO_171 (O_171,N_14643,N_14709);
nand UO_172 (O_172,N_14936,N_14623);
or UO_173 (O_173,N_14568,N_14958);
nor UO_174 (O_174,N_14362,N_14544);
nand UO_175 (O_175,N_14307,N_14745);
and UO_176 (O_176,N_14446,N_14382);
and UO_177 (O_177,N_14389,N_14812);
and UO_178 (O_178,N_14272,N_14640);
and UO_179 (O_179,N_14847,N_14430);
nand UO_180 (O_180,N_14444,N_14735);
nor UO_181 (O_181,N_14268,N_14774);
and UO_182 (O_182,N_14474,N_14498);
and UO_183 (O_183,N_14631,N_14994);
xor UO_184 (O_184,N_14566,N_14696);
or UO_185 (O_185,N_14750,N_14843);
xnor UO_186 (O_186,N_14825,N_14663);
xnor UO_187 (O_187,N_14322,N_14859);
nand UO_188 (O_188,N_14778,N_14460);
nand UO_189 (O_189,N_14976,N_14807);
or UO_190 (O_190,N_14796,N_14398);
nor UO_191 (O_191,N_14615,N_14491);
nand UO_192 (O_192,N_14742,N_14420);
and UO_193 (O_193,N_14260,N_14531);
nand UO_194 (O_194,N_14682,N_14302);
nor UO_195 (O_195,N_14280,N_14358);
nor UO_196 (O_196,N_14630,N_14822);
nand UO_197 (O_197,N_14751,N_14784);
nand UO_198 (O_198,N_14740,N_14440);
or UO_199 (O_199,N_14540,N_14380);
or UO_200 (O_200,N_14924,N_14369);
nor UO_201 (O_201,N_14769,N_14254);
and UO_202 (O_202,N_14721,N_14589);
nand UO_203 (O_203,N_14982,N_14370);
and UO_204 (O_204,N_14700,N_14829);
nor UO_205 (O_205,N_14918,N_14355);
and UO_206 (O_206,N_14561,N_14609);
nor UO_207 (O_207,N_14618,N_14633);
xor UO_208 (O_208,N_14510,N_14433);
or UO_209 (O_209,N_14532,N_14772);
and UO_210 (O_210,N_14548,N_14529);
or UO_211 (O_211,N_14704,N_14525);
nand UO_212 (O_212,N_14984,N_14620);
and UO_213 (O_213,N_14900,N_14508);
nor UO_214 (O_214,N_14519,N_14373);
and UO_215 (O_215,N_14426,N_14701);
nand UO_216 (O_216,N_14596,N_14309);
nor UO_217 (O_217,N_14712,N_14520);
and UO_218 (O_218,N_14551,N_14877);
nor UO_219 (O_219,N_14622,N_14927);
nand UO_220 (O_220,N_14660,N_14651);
nor UO_221 (O_221,N_14823,N_14754);
nand UO_222 (O_222,N_14397,N_14411);
and UO_223 (O_223,N_14697,N_14283);
nand UO_224 (O_224,N_14788,N_14914);
or UO_225 (O_225,N_14458,N_14506);
nand UO_226 (O_226,N_14427,N_14584);
and UO_227 (O_227,N_14281,N_14820);
nor UO_228 (O_228,N_14969,N_14466);
or UO_229 (O_229,N_14619,N_14855);
or UO_230 (O_230,N_14833,N_14306);
nor UO_231 (O_231,N_14448,N_14653);
nor UO_232 (O_232,N_14570,N_14555);
or UO_233 (O_233,N_14576,N_14909);
nand UO_234 (O_234,N_14598,N_14592);
or UO_235 (O_235,N_14512,N_14789);
nor UO_236 (O_236,N_14658,N_14723);
nor UO_237 (O_237,N_14343,N_14808);
or UO_238 (O_238,N_14297,N_14831);
and UO_239 (O_239,N_14454,N_14732);
and UO_240 (O_240,N_14876,N_14588);
or UO_241 (O_241,N_14947,N_14824);
and UO_242 (O_242,N_14813,N_14840);
and UO_243 (O_243,N_14608,N_14665);
xor UO_244 (O_244,N_14511,N_14265);
or UO_245 (O_245,N_14552,N_14949);
nor UO_246 (O_246,N_14988,N_14590);
xor UO_247 (O_247,N_14879,N_14416);
or UO_248 (O_248,N_14257,N_14715);
or UO_249 (O_249,N_14891,N_14441);
and UO_250 (O_250,N_14710,N_14330);
nand UO_251 (O_251,N_14499,N_14783);
nand UO_252 (O_252,N_14811,N_14459);
or UO_253 (O_253,N_14861,N_14495);
nor UO_254 (O_254,N_14810,N_14964);
or UO_255 (O_255,N_14872,N_14993);
nor UO_256 (O_256,N_14733,N_14996);
and UO_257 (O_257,N_14351,N_14554);
nor UO_258 (O_258,N_14279,N_14856);
or UO_259 (O_259,N_14395,N_14419);
and UO_260 (O_260,N_14318,N_14517);
nand UO_261 (O_261,N_14366,N_14761);
nand UO_262 (O_262,N_14952,N_14606);
and UO_263 (O_263,N_14258,N_14572);
and UO_264 (O_264,N_14693,N_14324);
or UO_265 (O_265,N_14867,N_14563);
nor UO_266 (O_266,N_14869,N_14575);
nor UO_267 (O_267,N_14514,N_14547);
and UO_268 (O_268,N_14664,N_14848);
nand UO_269 (O_269,N_14786,N_14897);
or UO_270 (O_270,N_14388,N_14899);
or UO_271 (O_271,N_14690,N_14938);
or UO_272 (O_272,N_14452,N_14637);
nand UO_273 (O_273,N_14844,N_14648);
nand UO_274 (O_274,N_14887,N_14668);
nand UO_275 (O_275,N_14970,N_14780);
nor UO_276 (O_276,N_14345,N_14752);
nand UO_277 (O_277,N_14628,N_14747);
nand UO_278 (O_278,N_14734,N_14311);
nor UO_279 (O_279,N_14333,N_14915);
nand UO_280 (O_280,N_14331,N_14800);
and UO_281 (O_281,N_14327,N_14390);
or UO_282 (O_282,N_14546,N_14381);
or UO_283 (O_283,N_14276,N_14882);
nor UO_284 (O_284,N_14836,N_14966);
or UO_285 (O_285,N_14312,N_14305);
nand UO_286 (O_286,N_14263,N_14901);
or UO_287 (O_287,N_14694,N_14553);
nand UO_288 (O_288,N_14368,N_14726);
nand UO_289 (O_289,N_14758,N_14911);
nand UO_290 (O_290,N_14756,N_14349);
nand UO_291 (O_291,N_14285,N_14286);
or UO_292 (O_292,N_14980,N_14713);
or UO_293 (O_293,N_14472,N_14505);
or UO_294 (O_294,N_14809,N_14990);
nand UO_295 (O_295,N_14893,N_14337);
or UO_296 (O_296,N_14912,N_14795);
and UO_297 (O_297,N_14647,N_14743);
xor UO_298 (O_298,N_14941,N_14948);
or UO_299 (O_299,N_14777,N_14326);
nor UO_300 (O_300,N_14296,N_14802);
nor UO_301 (O_301,N_14883,N_14655);
and UO_302 (O_302,N_14931,N_14542);
nand UO_303 (O_303,N_14903,N_14391);
nand UO_304 (O_304,N_14866,N_14259);
and UO_305 (O_305,N_14906,N_14850);
and UO_306 (O_306,N_14667,N_14581);
and UO_307 (O_307,N_14852,N_14401);
nor UO_308 (O_308,N_14661,N_14675);
nand UO_309 (O_309,N_14641,N_14597);
nand UO_310 (O_310,N_14858,N_14614);
and UO_311 (O_311,N_14739,N_14849);
or UO_312 (O_312,N_14759,N_14839);
nand UO_313 (O_313,N_14277,N_14611);
or UO_314 (O_314,N_14356,N_14404);
nor UO_315 (O_315,N_14479,N_14727);
nor UO_316 (O_316,N_14895,N_14492);
or UO_317 (O_317,N_14725,N_14617);
or UO_318 (O_318,N_14798,N_14558);
nand UO_319 (O_319,N_14429,N_14292);
or UO_320 (O_320,N_14974,N_14999);
nand UO_321 (O_321,N_14937,N_14862);
nor UO_322 (O_322,N_14881,N_14378);
nor UO_323 (O_323,N_14645,N_14593);
and UO_324 (O_324,N_14545,N_14841);
nor UO_325 (O_325,N_14830,N_14674);
nand UO_326 (O_326,N_14985,N_14794);
and UO_327 (O_327,N_14565,N_14771);
and UO_328 (O_328,N_14873,N_14685);
nor UO_329 (O_329,N_14711,N_14334);
nand UO_330 (O_330,N_14583,N_14310);
or UO_331 (O_331,N_14703,N_14336);
or UO_332 (O_332,N_14415,N_14942);
nand UO_333 (O_333,N_14360,N_14706);
or UO_334 (O_334,N_14308,N_14332);
or UO_335 (O_335,N_14375,N_14736);
nor UO_336 (O_336,N_14919,N_14504);
nand UO_337 (O_337,N_14603,N_14962);
or UO_338 (O_338,N_14764,N_14720);
or UO_339 (O_339,N_14423,N_14434);
nor UO_340 (O_340,N_14521,N_14781);
or UO_341 (O_341,N_14533,N_14790);
and UO_342 (O_342,N_14613,N_14662);
or UO_343 (O_343,N_14874,N_14456);
or UO_344 (O_344,N_14634,N_14438);
nand UO_345 (O_345,N_14705,N_14928);
nor UO_346 (O_346,N_14842,N_14717);
and UO_347 (O_347,N_14255,N_14367);
nand UO_348 (O_348,N_14431,N_14363);
nor UO_349 (O_349,N_14595,N_14450);
nor UO_350 (O_350,N_14639,N_14289);
nand UO_351 (O_351,N_14449,N_14577);
nand UO_352 (O_352,N_14763,N_14845);
and UO_353 (O_353,N_14922,N_14516);
and UO_354 (O_354,N_14687,N_14437);
and UO_355 (O_355,N_14522,N_14857);
nand UO_356 (O_356,N_14443,N_14338);
nand UO_357 (O_357,N_14860,N_14353);
or UO_358 (O_358,N_14638,N_14601);
or UO_359 (O_359,N_14410,N_14760);
nor UO_360 (O_360,N_14799,N_14304);
and UO_361 (O_361,N_14785,N_14526);
or UO_362 (O_362,N_14435,N_14722);
nand UO_363 (O_363,N_14695,N_14884);
and UO_364 (O_364,N_14482,N_14562);
and UO_365 (O_365,N_14757,N_14765);
nor UO_366 (O_366,N_14396,N_14384);
and UO_367 (O_367,N_14898,N_14266);
and UO_368 (O_368,N_14413,N_14801);
nand UO_369 (O_369,N_14870,N_14489);
or UO_370 (O_370,N_14827,N_14755);
nor UO_371 (O_371,N_14509,N_14921);
nor UO_372 (O_372,N_14319,N_14303);
nor UO_373 (O_373,N_14666,N_14376);
or UO_374 (O_374,N_14432,N_14374);
or UO_375 (O_375,N_14622,N_14860);
nor UO_376 (O_376,N_14700,N_14532);
or UO_377 (O_377,N_14692,N_14729);
nor UO_378 (O_378,N_14855,N_14904);
and UO_379 (O_379,N_14738,N_14544);
and UO_380 (O_380,N_14992,N_14455);
or UO_381 (O_381,N_14676,N_14804);
nand UO_382 (O_382,N_14681,N_14814);
or UO_383 (O_383,N_14749,N_14599);
and UO_384 (O_384,N_14937,N_14789);
nand UO_385 (O_385,N_14349,N_14285);
and UO_386 (O_386,N_14961,N_14983);
and UO_387 (O_387,N_14564,N_14551);
and UO_388 (O_388,N_14731,N_14458);
nand UO_389 (O_389,N_14564,N_14548);
xnor UO_390 (O_390,N_14277,N_14434);
and UO_391 (O_391,N_14586,N_14533);
or UO_392 (O_392,N_14677,N_14768);
nand UO_393 (O_393,N_14667,N_14349);
nor UO_394 (O_394,N_14888,N_14837);
and UO_395 (O_395,N_14699,N_14488);
nor UO_396 (O_396,N_14335,N_14971);
and UO_397 (O_397,N_14270,N_14959);
nand UO_398 (O_398,N_14424,N_14649);
and UO_399 (O_399,N_14606,N_14320);
or UO_400 (O_400,N_14833,N_14879);
nand UO_401 (O_401,N_14669,N_14620);
and UO_402 (O_402,N_14578,N_14990);
nor UO_403 (O_403,N_14568,N_14858);
and UO_404 (O_404,N_14498,N_14605);
xor UO_405 (O_405,N_14702,N_14534);
or UO_406 (O_406,N_14835,N_14514);
nand UO_407 (O_407,N_14555,N_14414);
nand UO_408 (O_408,N_14315,N_14422);
and UO_409 (O_409,N_14637,N_14455);
or UO_410 (O_410,N_14612,N_14557);
and UO_411 (O_411,N_14551,N_14372);
nand UO_412 (O_412,N_14923,N_14307);
nand UO_413 (O_413,N_14398,N_14502);
nor UO_414 (O_414,N_14328,N_14646);
nand UO_415 (O_415,N_14904,N_14931);
and UO_416 (O_416,N_14857,N_14439);
and UO_417 (O_417,N_14904,N_14445);
and UO_418 (O_418,N_14354,N_14857);
nand UO_419 (O_419,N_14933,N_14285);
nor UO_420 (O_420,N_14915,N_14416);
or UO_421 (O_421,N_14551,N_14785);
nor UO_422 (O_422,N_14552,N_14959);
and UO_423 (O_423,N_14735,N_14652);
nand UO_424 (O_424,N_14552,N_14862);
nand UO_425 (O_425,N_14492,N_14725);
or UO_426 (O_426,N_14861,N_14300);
nor UO_427 (O_427,N_14818,N_14707);
nor UO_428 (O_428,N_14717,N_14350);
and UO_429 (O_429,N_14961,N_14349);
nand UO_430 (O_430,N_14319,N_14994);
and UO_431 (O_431,N_14365,N_14307);
nor UO_432 (O_432,N_14666,N_14388);
and UO_433 (O_433,N_14459,N_14498);
nand UO_434 (O_434,N_14273,N_14320);
nor UO_435 (O_435,N_14395,N_14830);
nor UO_436 (O_436,N_14709,N_14613);
nor UO_437 (O_437,N_14375,N_14755);
and UO_438 (O_438,N_14828,N_14630);
and UO_439 (O_439,N_14373,N_14514);
nor UO_440 (O_440,N_14901,N_14643);
nor UO_441 (O_441,N_14684,N_14617);
and UO_442 (O_442,N_14948,N_14265);
nor UO_443 (O_443,N_14926,N_14282);
nor UO_444 (O_444,N_14434,N_14714);
nor UO_445 (O_445,N_14766,N_14755);
nor UO_446 (O_446,N_14917,N_14810);
or UO_447 (O_447,N_14630,N_14288);
and UO_448 (O_448,N_14399,N_14967);
and UO_449 (O_449,N_14957,N_14643);
and UO_450 (O_450,N_14593,N_14755);
nand UO_451 (O_451,N_14945,N_14279);
or UO_452 (O_452,N_14327,N_14662);
nand UO_453 (O_453,N_14555,N_14911);
or UO_454 (O_454,N_14984,N_14751);
or UO_455 (O_455,N_14983,N_14379);
or UO_456 (O_456,N_14434,N_14781);
nor UO_457 (O_457,N_14549,N_14603);
or UO_458 (O_458,N_14893,N_14388);
and UO_459 (O_459,N_14574,N_14887);
nand UO_460 (O_460,N_14582,N_14921);
or UO_461 (O_461,N_14289,N_14446);
and UO_462 (O_462,N_14300,N_14958);
nor UO_463 (O_463,N_14745,N_14489);
nand UO_464 (O_464,N_14388,N_14697);
nand UO_465 (O_465,N_14996,N_14958);
nor UO_466 (O_466,N_14953,N_14380);
or UO_467 (O_467,N_14562,N_14481);
and UO_468 (O_468,N_14526,N_14310);
nand UO_469 (O_469,N_14630,N_14420);
and UO_470 (O_470,N_14474,N_14966);
or UO_471 (O_471,N_14898,N_14922);
and UO_472 (O_472,N_14483,N_14817);
and UO_473 (O_473,N_14632,N_14278);
nor UO_474 (O_474,N_14629,N_14478);
nor UO_475 (O_475,N_14736,N_14498);
and UO_476 (O_476,N_14609,N_14782);
or UO_477 (O_477,N_14447,N_14738);
or UO_478 (O_478,N_14729,N_14420);
nor UO_479 (O_479,N_14987,N_14875);
nor UO_480 (O_480,N_14633,N_14915);
and UO_481 (O_481,N_14346,N_14573);
or UO_482 (O_482,N_14853,N_14641);
or UO_483 (O_483,N_14407,N_14602);
nand UO_484 (O_484,N_14820,N_14651);
nor UO_485 (O_485,N_14558,N_14499);
or UO_486 (O_486,N_14879,N_14595);
and UO_487 (O_487,N_14916,N_14674);
nor UO_488 (O_488,N_14569,N_14848);
nor UO_489 (O_489,N_14945,N_14631);
nand UO_490 (O_490,N_14819,N_14731);
or UO_491 (O_491,N_14689,N_14690);
or UO_492 (O_492,N_14395,N_14439);
nor UO_493 (O_493,N_14951,N_14279);
or UO_494 (O_494,N_14286,N_14621);
nor UO_495 (O_495,N_14959,N_14836);
nand UO_496 (O_496,N_14280,N_14835);
and UO_497 (O_497,N_14292,N_14418);
nor UO_498 (O_498,N_14869,N_14652);
and UO_499 (O_499,N_14496,N_14668);
nand UO_500 (O_500,N_14792,N_14512);
nand UO_501 (O_501,N_14968,N_14615);
nand UO_502 (O_502,N_14860,N_14771);
nor UO_503 (O_503,N_14916,N_14797);
nor UO_504 (O_504,N_14733,N_14782);
or UO_505 (O_505,N_14849,N_14864);
and UO_506 (O_506,N_14754,N_14584);
and UO_507 (O_507,N_14811,N_14552);
nand UO_508 (O_508,N_14774,N_14607);
or UO_509 (O_509,N_14782,N_14310);
and UO_510 (O_510,N_14438,N_14269);
nand UO_511 (O_511,N_14633,N_14968);
and UO_512 (O_512,N_14272,N_14752);
nand UO_513 (O_513,N_14908,N_14839);
or UO_514 (O_514,N_14385,N_14915);
and UO_515 (O_515,N_14633,N_14756);
nor UO_516 (O_516,N_14590,N_14547);
or UO_517 (O_517,N_14692,N_14705);
nor UO_518 (O_518,N_14765,N_14595);
or UO_519 (O_519,N_14665,N_14821);
nor UO_520 (O_520,N_14488,N_14672);
and UO_521 (O_521,N_14675,N_14715);
or UO_522 (O_522,N_14382,N_14726);
nand UO_523 (O_523,N_14829,N_14592);
and UO_524 (O_524,N_14554,N_14953);
or UO_525 (O_525,N_14300,N_14266);
nor UO_526 (O_526,N_14673,N_14781);
nand UO_527 (O_527,N_14303,N_14383);
nand UO_528 (O_528,N_14252,N_14721);
and UO_529 (O_529,N_14704,N_14622);
nor UO_530 (O_530,N_14853,N_14335);
nand UO_531 (O_531,N_14440,N_14668);
and UO_532 (O_532,N_14745,N_14934);
or UO_533 (O_533,N_14485,N_14324);
and UO_534 (O_534,N_14304,N_14612);
nand UO_535 (O_535,N_14814,N_14686);
or UO_536 (O_536,N_14855,N_14443);
and UO_537 (O_537,N_14634,N_14268);
and UO_538 (O_538,N_14942,N_14959);
nor UO_539 (O_539,N_14737,N_14454);
nor UO_540 (O_540,N_14410,N_14815);
nor UO_541 (O_541,N_14500,N_14708);
nand UO_542 (O_542,N_14786,N_14919);
nand UO_543 (O_543,N_14255,N_14892);
nor UO_544 (O_544,N_14254,N_14409);
nand UO_545 (O_545,N_14769,N_14761);
and UO_546 (O_546,N_14888,N_14287);
nand UO_547 (O_547,N_14359,N_14883);
and UO_548 (O_548,N_14642,N_14594);
nand UO_549 (O_549,N_14365,N_14380);
or UO_550 (O_550,N_14788,N_14261);
nor UO_551 (O_551,N_14686,N_14919);
and UO_552 (O_552,N_14678,N_14442);
or UO_553 (O_553,N_14392,N_14989);
and UO_554 (O_554,N_14766,N_14891);
or UO_555 (O_555,N_14877,N_14478);
nor UO_556 (O_556,N_14538,N_14748);
and UO_557 (O_557,N_14572,N_14575);
or UO_558 (O_558,N_14415,N_14448);
nand UO_559 (O_559,N_14657,N_14618);
nor UO_560 (O_560,N_14502,N_14977);
and UO_561 (O_561,N_14773,N_14694);
or UO_562 (O_562,N_14920,N_14825);
nand UO_563 (O_563,N_14931,N_14373);
nand UO_564 (O_564,N_14867,N_14912);
nand UO_565 (O_565,N_14894,N_14965);
nand UO_566 (O_566,N_14378,N_14928);
or UO_567 (O_567,N_14981,N_14490);
nand UO_568 (O_568,N_14458,N_14778);
nor UO_569 (O_569,N_14640,N_14404);
and UO_570 (O_570,N_14635,N_14552);
and UO_571 (O_571,N_14491,N_14543);
or UO_572 (O_572,N_14779,N_14321);
or UO_573 (O_573,N_14736,N_14944);
nor UO_574 (O_574,N_14722,N_14935);
and UO_575 (O_575,N_14861,N_14829);
and UO_576 (O_576,N_14866,N_14815);
nand UO_577 (O_577,N_14698,N_14433);
nand UO_578 (O_578,N_14719,N_14859);
nor UO_579 (O_579,N_14609,N_14862);
nand UO_580 (O_580,N_14589,N_14317);
and UO_581 (O_581,N_14870,N_14480);
and UO_582 (O_582,N_14983,N_14571);
or UO_583 (O_583,N_14254,N_14443);
nor UO_584 (O_584,N_14864,N_14761);
nor UO_585 (O_585,N_14763,N_14593);
or UO_586 (O_586,N_14899,N_14851);
or UO_587 (O_587,N_14804,N_14514);
nor UO_588 (O_588,N_14812,N_14617);
and UO_589 (O_589,N_14977,N_14606);
and UO_590 (O_590,N_14775,N_14503);
or UO_591 (O_591,N_14694,N_14460);
and UO_592 (O_592,N_14977,N_14552);
nand UO_593 (O_593,N_14569,N_14811);
nand UO_594 (O_594,N_14779,N_14587);
nor UO_595 (O_595,N_14757,N_14394);
or UO_596 (O_596,N_14653,N_14472);
or UO_597 (O_597,N_14369,N_14624);
and UO_598 (O_598,N_14738,N_14393);
and UO_599 (O_599,N_14716,N_14501);
or UO_600 (O_600,N_14592,N_14732);
and UO_601 (O_601,N_14496,N_14924);
nand UO_602 (O_602,N_14402,N_14413);
nand UO_603 (O_603,N_14670,N_14734);
nand UO_604 (O_604,N_14948,N_14789);
and UO_605 (O_605,N_14454,N_14959);
and UO_606 (O_606,N_14735,N_14323);
nand UO_607 (O_607,N_14801,N_14841);
or UO_608 (O_608,N_14447,N_14277);
nand UO_609 (O_609,N_14648,N_14561);
nand UO_610 (O_610,N_14480,N_14961);
and UO_611 (O_611,N_14588,N_14644);
nor UO_612 (O_612,N_14253,N_14630);
nor UO_613 (O_613,N_14320,N_14741);
nor UO_614 (O_614,N_14622,N_14489);
and UO_615 (O_615,N_14855,N_14617);
and UO_616 (O_616,N_14333,N_14929);
and UO_617 (O_617,N_14980,N_14736);
and UO_618 (O_618,N_14900,N_14503);
nand UO_619 (O_619,N_14545,N_14809);
or UO_620 (O_620,N_14873,N_14609);
and UO_621 (O_621,N_14821,N_14968);
nand UO_622 (O_622,N_14669,N_14820);
and UO_623 (O_623,N_14285,N_14653);
nand UO_624 (O_624,N_14481,N_14311);
or UO_625 (O_625,N_14650,N_14938);
and UO_626 (O_626,N_14487,N_14666);
nor UO_627 (O_627,N_14438,N_14667);
or UO_628 (O_628,N_14816,N_14503);
nor UO_629 (O_629,N_14549,N_14361);
or UO_630 (O_630,N_14321,N_14452);
or UO_631 (O_631,N_14805,N_14250);
and UO_632 (O_632,N_14875,N_14905);
and UO_633 (O_633,N_14961,N_14911);
nand UO_634 (O_634,N_14499,N_14550);
or UO_635 (O_635,N_14663,N_14960);
and UO_636 (O_636,N_14660,N_14945);
nand UO_637 (O_637,N_14875,N_14698);
and UO_638 (O_638,N_14947,N_14827);
nor UO_639 (O_639,N_14583,N_14724);
nand UO_640 (O_640,N_14991,N_14827);
nand UO_641 (O_641,N_14991,N_14736);
or UO_642 (O_642,N_14877,N_14427);
or UO_643 (O_643,N_14579,N_14974);
nand UO_644 (O_644,N_14555,N_14827);
or UO_645 (O_645,N_14883,N_14619);
nand UO_646 (O_646,N_14956,N_14424);
nand UO_647 (O_647,N_14407,N_14463);
nand UO_648 (O_648,N_14355,N_14633);
nand UO_649 (O_649,N_14577,N_14745);
nor UO_650 (O_650,N_14509,N_14989);
nand UO_651 (O_651,N_14289,N_14997);
nor UO_652 (O_652,N_14510,N_14828);
nor UO_653 (O_653,N_14878,N_14769);
and UO_654 (O_654,N_14837,N_14727);
nand UO_655 (O_655,N_14536,N_14984);
or UO_656 (O_656,N_14661,N_14573);
or UO_657 (O_657,N_14672,N_14589);
nand UO_658 (O_658,N_14383,N_14851);
nand UO_659 (O_659,N_14684,N_14287);
nand UO_660 (O_660,N_14778,N_14862);
or UO_661 (O_661,N_14953,N_14376);
nor UO_662 (O_662,N_14667,N_14369);
nor UO_663 (O_663,N_14703,N_14805);
nor UO_664 (O_664,N_14535,N_14368);
nand UO_665 (O_665,N_14356,N_14716);
and UO_666 (O_666,N_14406,N_14426);
and UO_667 (O_667,N_14611,N_14386);
and UO_668 (O_668,N_14576,N_14859);
and UO_669 (O_669,N_14877,N_14405);
nor UO_670 (O_670,N_14447,N_14254);
or UO_671 (O_671,N_14866,N_14944);
nand UO_672 (O_672,N_14429,N_14695);
or UO_673 (O_673,N_14503,N_14863);
nand UO_674 (O_674,N_14616,N_14599);
nor UO_675 (O_675,N_14279,N_14446);
or UO_676 (O_676,N_14723,N_14352);
and UO_677 (O_677,N_14598,N_14850);
or UO_678 (O_678,N_14499,N_14941);
and UO_679 (O_679,N_14820,N_14809);
and UO_680 (O_680,N_14944,N_14890);
nand UO_681 (O_681,N_14289,N_14582);
nor UO_682 (O_682,N_14420,N_14994);
or UO_683 (O_683,N_14677,N_14755);
and UO_684 (O_684,N_14757,N_14724);
nand UO_685 (O_685,N_14265,N_14852);
nand UO_686 (O_686,N_14448,N_14496);
and UO_687 (O_687,N_14329,N_14859);
and UO_688 (O_688,N_14837,N_14856);
nand UO_689 (O_689,N_14537,N_14316);
nor UO_690 (O_690,N_14273,N_14659);
or UO_691 (O_691,N_14605,N_14348);
nand UO_692 (O_692,N_14879,N_14329);
and UO_693 (O_693,N_14715,N_14373);
nor UO_694 (O_694,N_14334,N_14394);
nor UO_695 (O_695,N_14411,N_14738);
nand UO_696 (O_696,N_14293,N_14806);
nand UO_697 (O_697,N_14691,N_14964);
nor UO_698 (O_698,N_14376,N_14371);
or UO_699 (O_699,N_14279,N_14954);
nand UO_700 (O_700,N_14481,N_14898);
and UO_701 (O_701,N_14962,N_14565);
nand UO_702 (O_702,N_14745,N_14381);
nor UO_703 (O_703,N_14596,N_14766);
or UO_704 (O_704,N_14380,N_14288);
nand UO_705 (O_705,N_14457,N_14529);
nand UO_706 (O_706,N_14290,N_14774);
nor UO_707 (O_707,N_14679,N_14587);
or UO_708 (O_708,N_14799,N_14623);
and UO_709 (O_709,N_14539,N_14840);
nor UO_710 (O_710,N_14338,N_14638);
nor UO_711 (O_711,N_14990,N_14644);
nand UO_712 (O_712,N_14981,N_14363);
nand UO_713 (O_713,N_14867,N_14459);
and UO_714 (O_714,N_14710,N_14281);
nand UO_715 (O_715,N_14915,N_14295);
nand UO_716 (O_716,N_14742,N_14263);
nor UO_717 (O_717,N_14893,N_14364);
nor UO_718 (O_718,N_14758,N_14545);
and UO_719 (O_719,N_14498,N_14347);
or UO_720 (O_720,N_14758,N_14742);
or UO_721 (O_721,N_14268,N_14390);
nor UO_722 (O_722,N_14306,N_14724);
and UO_723 (O_723,N_14256,N_14505);
and UO_724 (O_724,N_14808,N_14259);
or UO_725 (O_725,N_14345,N_14372);
nor UO_726 (O_726,N_14442,N_14796);
nand UO_727 (O_727,N_14477,N_14647);
and UO_728 (O_728,N_14963,N_14826);
nor UO_729 (O_729,N_14337,N_14914);
or UO_730 (O_730,N_14674,N_14874);
or UO_731 (O_731,N_14681,N_14516);
nor UO_732 (O_732,N_14716,N_14407);
and UO_733 (O_733,N_14632,N_14687);
nor UO_734 (O_734,N_14297,N_14815);
nor UO_735 (O_735,N_14301,N_14554);
nand UO_736 (O_736,N_14582,N_14264);
and UO_737 (O_737,N_14495,N_14572);
nand UO_738 (O_738,N_14799,N_14880);
or UO_739 (O_739,N_14442,N_14396);
nor UO_740 (O_740,N_14267,N_14331);
nand UO_741 (O_741,N_14409,N_14897);
or UO_742 (O_742,N_14417,N_14917);
or UO_743 (O_743,N_14437,N_14260);
nand UO_744 (O_744,N_14401,N_14526);
and UO_745 (O_745,N_14802,N_14306);
and UO_746 (O_746,N_14283,N_14263);
nand UO_747 (O_747,N_14880,N_14677);
or UO_748 (O_748,N_14434,N_14550);
and UO_749 (O_749,N_14764,N_14387);
xnor UO_750 (O_750,N_14562,N_14690);
and UO_751 (O_751,N_14476,N_14513);
nor UO_752 (O_752,N_14371,N_14883);
and UO_753 (O_753,N_14932,N_14850);
or UO_754 (O_754,N_14531,N_14692);
and UO_755 (O_755,N_14412,N_14385);
nand UO_756 (O_756,N_14774,N_14967);
nor UO_757 (O_757,N_14743,N_14856);
nor UO_758 (O_758,N_14850,N_14459);
or UO_759 (O_759,N_14528,N_14971);
and UO_760 (O_760,N_14292,N_14491);
or UO_761 (O_761,N_14791,N_14621);
nand UO_762 (O_762,N_14715,N_14252);
or UO_763 (O_763,N_14807,N_14718);
nand UO_764 (O_764,N_14413,N_14567);
and UO_765 (O_765,N_14788,N_14562);
nor UO_766 (O_766,N_14389,N_14846);
nor UO_767 (O_767,N_14396,N_14267);
and UO_768 (O_768,N_14510,N_14551);
nor UO_769 (O_769,N_14397,N_14843);
nand UO_770 (O_770,N_14553,N_14745);
nor UO_771 (O_771,N_14389,N_14581);
nand UO_772 (O_772,N_14270,N_14709);
nand UO_773 (O_773,N_14805,N_14458);
or UO_774 (O_774,N_14993,N_14767);
nor UO_775 (O_775,N_14280,N_14977);
and UO_776 (O_776,N_14256,N_14885);
nand UO_777 (O_777,N_14847,N_14669);
and UO_778 (O_778,N_14596,N_14752);
and UO_779 (O_779,N_14598,N_14322);
nand UO_780 (O_780,N_14562,N_14763);
or UO_781 (O_781,N_14543,N_14384);
nand UO_782 (O_782,N_14654,N_14958);
nor UO_783 (O_783,N_14635,N_14855);
or UO_784 (O_784,N_14290,N_14947);
nand UO_785 (O_785,N_14919,N_14903);
nand UO_786 (O_786,N_14370,N_14443);
nand UO_787 (O_787,N_14948,N_14262);
nand UO_788 (O_788,N_14778,N_14429);
and UO_789 (O_789,N_14793,N_14891);
and UO_790 (O_790,N_14873,N_14646);
nor UO_791 (O_791,N_14907,N_14330);
nor UO_792 (O_792,N_14803,N_14435);
and UO_793 (O_793,N_14767,N_14700);
nor UO_794 (O_794,N_14619,N_14950);
and UO_795 (O_795,N_14930,N_14892);
nand UO_796 (O_796,N_14280,N_14711);
nand UO_797 (O_797,N_14726,N_14862);
or UO_798 (O_798,N_14656,N_14759);
or UO_799 (O_799,N_14994,N_14512);
nand UO_800 (O_800,N_14434,N_14790);
or UO_801 (O_801,N_14537,N_14301);
nor UO_802 (O_802,N_14931,N_14315);
or UO_803 (O_803,N_14634,N_14967);
nand UO_804 (O_804,N_14914,N_14324);
or UO_805 (O_805,N_14746,N_14521);
nand UO_806 (O_806,N_14574,N_14545);
nand UO_807 (O_807,N_14645,N_14388);
and UO_808 (O_808,N_14990,N_14312);
and UO_809 (O_809,N_14830,N_14273);
nand UO_810 (O_810,N_14500,N_14604);
nor UO_811 (O_811,N_14828,N_14722);
nor UO_812 (O_812,N_14627,N_14527);
or UO_813 (O_813,N_14813,N_14689);
nand UO_814 (O_814,N_14907,N_14304);
and UO_815 (O_815,N_14447,N_14334);
nor UO_816 (O_816,N_14625,N_14735);
nand UO_817 (O_817,N_14833,N_14512);
or UO_818 (O_818,N_14386,N_14603);
nand UO_819 (O_819,N_14321,N_14327);
or UO_820 (O_820,N_14969,N_14840);
nand UO_821 (O_821,N_14258,N_14414);
or UO_822 (O_822,N_14479,N_14495);
nand UO_823 (O_823,N_14710,N_14516);
nor UO_824 (O_824,N_14671,N_14666);
and UO_825 (O_825,N_14952,N_14967);
nand UO_826 (O_826,N_14513,N_14481);
or UO_827 (O_827,N_14284,N_14321);
nor UO_828 (O_828,N_14665,N_14997);
nand UO_829 (O_829,N_14768,N_14771);
and UO_830 (O_830,N_14884,N_14849);
nor UO_831 (O_831,N_14970,N_14867);
and UO_832 (O_832,N_14898,N_14926);
or UO_833 (O_833,N_14485,N_14481);
nand UO_834 (O_834,N_14437,N_14580);
and UO_835 (O_835,N_14631,N_14325);
and UO_836 (O_836,N_14586,N_14397);
nand UO_837 (O_837,N_14690,N_14353);
and UO_838 (O_838,N_14325,N_14500);
nor UO_839 (O_839,N_14545,N_14333);
nand UO_840 (O_840,N_14620,N_14297);
and UO_841 (O_841,N_14817,N_14851);
xor UO_842 (O_842,N_14385,N_14853);
nand UO_843 (O_843,N_14983,N_14292);
and UO_844 (O_844,N_14803,N_14284);
nand UO_845 (O_845,N_14380,N_14301);
or UO_846 (O_846,N_14996,N_14256);
or UO_847 (O_847,N_14365,N_14668);
or UO_848 (O_848,N_14406,N_14764);
or UO_849 (O_849,N_14642,N_14958);
nand UO_850 (O_850,N_14904,N_14599);
or UO_851 (O_851,N_14483,N_14386);
and UO_852 (O_852,N_14674,N_14375);
nand UO_853 (O_853,N_14838,N_14689);
and UO_854 (O_854,N_14868,N_14347);
nand UO_855 (O_855,N_14528,N_14939);
nor UO_856 (O_856,N_14903,N_14567);
or UO_857 (O_857,N_14760,N_14608);
nand UO_858 (O_858,N_14713,N_14727);
or UO_859 (O_859,N_14533,N_14990);
xor UO_860 (O_860,N_14417,N_14662);
nor UO_861 (O_861,N_14746,N_14827);
and UO_862 (O_862,N_14596,N_14963);
and UO_863 (O_863,N_14885,N_14411);
or UO_864 (O_864,N_14397,N_14949);
nor UO_865 (O_865,N_14692,N_14932);
nor UO_866 (O_866,N_14714,N_14341);
and UO_867 (O_867,N_14431,N_14468);
or UO_868 (O_868,N_14719,N_14736);
nand UO_869 (O_869,N_14446,N_14420);
and UO_870 (O_870,N_14779,N_14311);
or UO_871 (O_871,N_14605,N_14440);
nand UO_872 (O_872,N_14891,N_14444);
nand UO_873 (O_873,N_14673,N_14315);
or UO_874 (O_874,N_14616,N_14487);
nor UO_875 (O_875,N_14799,N_14308);
nand UO_876 (O_876,N_14544,N_14974);
and UO_877 (O_877,N_14602,N_14366);
nand UO_878 (O_878,N_14402,N_14547);
or UO_879 (O_879,N_14865,N_14263);
or UO_880 (O_880,N_14293,N_14826);
or UO_881 (O_881,N_14417,N_14621);
or UO_882 (O_882,N_14740,N_14386);
nand UO_883 (O_883,N_14368,N_14746);
nand UO_884 (O_884,N_14628,N_14334);
and UO_885 (O_885,N_14749,N_14565);
nand UO_886 (O_886,N_14786,N_14477);
and UO_887 (O_887,N_14399,N_14592);
nor UO_888 (O_888,N_14770,N_14632);
nor UO_889 (O_889,N_14615,N_14725);
and UO_890 (O_890,N_14653,N_14322);
nand UO_891 (O_891,N_14957,N_14655);
nand UO_892 (O_892,N_14514,N_14838);
or UO_893 (O_893,N_14387,N_14879);
nand UO_894 (O_894,N_14545,N_14342);
and UO_895 (O_895,N_14482,N_14631);
or UO_896 (O_896,N_14904,N_14463);
or UO_897 (O_897,N_14459,N_14906);
nand UO_898 (O_898,N_14414,N_14859);
and UO_899 (O_899,N_14775,N_14603);
nor UO_900 (O_900,N_14565,N_14344);
and UO_901 (O_901,N_14272,N_14996);
nor UO_902 (O_902,N_14690,N_14525);
nor UO_903 (O_903,N_14586,N_14284);
or UO_904 (O_904,N_14332,N_14869);
nand UO_905 (O_905,N_14328,N_14926);
nand UO_906 (O_906,N_14729,N_14615);
or UO_907 (O_907,N_14997,N_14971);
and UO_908 (O_908,N_14880,N_14265);
and UO_909 (O_909,N_14710,N_14547);
nand UO_910 (O_910,N_14441,N_14912);
xor UO_911 (O_911,N_14918,N_14598);
and UO_912 (O_912,N_14574,N_14656);
nand UO_913 (O_913,N_14512,N_14813);
and UO_914 (O_914,N_14602,N_14658);
or UO_915 (O_915,N_14905,N_14843);
nor UO_916 (O_916,N_14630,N_14318);
nor UO_917 (O_917,N_14829,N_14905);
nand UO_918 (O_918,N_14322,N_14403);
or UO_919 (O_919,N_14471,N_14780);
and UO_920 (O_920,N_14398,N_14811);
nor UO_921 (O_921,N_14555,N_14710);
nand UO_922 (O_922,N_14791,N_14764);
nand UO_923 (O_923,N_14662,N_14687);
nand UO_924 (O_924,N_14465,N_14879);
nand UO_925 (O_925,N_14317,N_14490);
nand UO_926 (O_926,N_14354,N_14861);
nor UO_927 (O_927,N_14518,N_14767);
and UO_928 (O_928,N_14701,N_14577);
nand UO_929 (O_929,N_14407,N_14572);
and UO_930 (O_930,N_14558,N_14995);
and UO_931 (O_931,N_14470,N_14543);
and UO_932 (O_932,N_14586,N_14578);
or UO_933 (O_933,N_14559,N_14797);
and UO_934 (O_934,N_14747,N_14253);
or UO_935 (O_935,N_14788,N_14637);
nand UO_936 (O_936,N_14497,N_14804);
nor UO_937 (O_937,N_14396,N_14511);
xnor UO_938 (O_938,N_14810,N_14271);
or UO_939 (O_939,N_14366,N_14378);
nor UO_940 (O_940,N_14252,N_14826);
or UO_941 (O_941,N_14409,N_14358);
xnor UO_942 (O_942,N_14431,N_14721);
nand UO_943 (O_943,N_14528,N_14967);
nand UO_944 (O_944,N_14438,N_14947);
nand UO_945 (O_945,N_14681,N_14793);
or UO_946 (O_946,N_14972,N_14632);
nand UO_947 (O_947,N_14762,N_14561);
nand UO_948 (O_948,N_14606,N_14967);
nand UO_949 (O_949,N_14782,N_14709);
or UO_950 (O_950,N_14540,N_14405);
nor UO_951 (O_951,N_14391,N_14999);
and UO_952 (O_952,N_14943,N_14843);
and UO_953 (O_953,N_14685,N_14976);
nor UO_954 (O_954,N_14605,N_14494);
and UO_955 (O_955,N_14561,N_14746);
nor UO_956 (O_956,N_14833,N_14417);
nand UO_957 (O_957,N_14325,N_14743);
nor UO_958 (O_958,N_14744,N_14313);
or UO_959 (O_959,N_14805,N_14732);
and UO_960 (O_960,N_14405,N_14862);
and UO_961 (O_961,N_14645,N_14810);
nand UO_962 (O_962,N_14555,N_14772);
nor UO_963 (O_963,N_14788,N_14845);
and UO_964 (O_964,N_14970,N_14428);
nand UO_965 (O_965,N_14617,N_14770);
and UO_966 (O_966,N_14536,N_14712);
or UO_967 (O_967,N_14984,N_14991);
or UO_968 (O_968,N_14794,N_14616);
and UO_969 (O_969,N_14520,N_14347);
xnor UO_970 (O_970,N_14427,N_14539);
nor UO_971 (O_971,N_14905,N_14783);
or UO_972 (O_972,N_14383,N_14562);
nor UO_973 (O_973,N_14297,N_14851);
or UO_974 (O_974,N_14883,N_14767);
nand UO_975 (O_975,N_14336,N_14675);
and UO_976 (O_976,N_14645,N_14656);
and UO_977 (O_977,N_14911,N_14360);
nand UO_978 (O_978,N_14845,N_14935);
nand UO_979 (O_979,N_14358,N_14407);
nand UO_980 (O_980,N_14629,N_14503);
and UO_981 (O_981,N_14966,N_14573);
nor UO_982 (O_982,N_14716,N_14857);
nor UO_983 (O_983,N_14783,N_14889);
or UO_984 (O_984,N_14354,N_14813);
nand UO_985 (O_985,N_14966,N_14493);
nor UO_986 (O_986,N_14680,N_14707);
nand UO_987 (O_987,N_14914,N_14947);
nand UO_988 (O_988,N_14562,N_14475);
and UO_989 (O_989,N_14587,N_14743);
or UO_990 (O_990,N_14472,N_14384);
nor UO_991 (O_991,N_14907,N_14449);
and UO_992 (O_992,N_14918,N_14334);
nor UO_993 (O_993,N_14638,N_14509);
and UO_994 (O_994,N_14485,N_14338);
or UO_995 (O_995,N_14284,N_14349);
or UO_996 (O_996,N_14954,N_14309);
nand UO_997 (O_997,N_14774,N_14809);
or UO_998 (O_998,N_14722,N_14926);
nand UO_999 (O_999,N_14545,N_14648);
nor UO_1000 (O_1000,N_14602,N_14547);
nand UO_1001 (O_1001,N_14370,N_14451);
or UO_1002 (O_1002,N_14397,N_14960);
or UO_1003 (O_1003,N_14332,N_14346);
nor UO_1004 (O_1004,N_14444,N_14284);
and UO_1005 (O_1005,N_14461,N_14427);
nand UO_1006 (O_1006,N_14674,N_14467);
nand UO_1007 (O_1007,N_14598,N_14962);
and UO_1008 (O_1008,N_14877,N_14677);
or UO_1009 (O_1009,N_14833,N_14414);
nand UO_1010 (O_1010,N_14765,N_14827);
or UO_1011 (O_1011,N_14745,N_14944);
nor UO_1012 (O_1012,N_14670,N_14351);
nand UO_1013 (O_1013,N_14728,N_14546);
nand UO_1014 (O_1014,N_14883,N_14449);
or UO_1015 (O_1015,N_14458,N_14296);
nand UO_1016 (O_1016,N_14331,N_14920);
and UO_1017 (O_1017,N_14881,N_14289);
nand UO_1018 (O_1018,N_14573,N_14668);
or UO_1019 (O_1019,N_14773,N_14304);
and UO_1020 (O_1020,N_14427,N_14879);
or UO_1021 (O_1021,N_14323,N_14633);
nor UO_1022 (O_1022,N_14414,N_14742);
or UO_1023 (O_1023,N_14885,N_14707);
nor UO_1024 (O_1024,N_14251,N_14482);
nor UO_1025 (O_1025,N_14692,N_14826);
nand UO_1026 (O_1026,N_14945,N_14502);
and UO_1027 (O_1027,N_14949,N_14859);
nand UO_1028 (O_1028,N_14579,N_14421);
or UO_1029 (O_1029,N_14577,N_14669);
nor UO_1030 (O_1030,N_14310,N_14704);
nand UO_1031 (O_1031,N_14714,N_14336);
nor UO_1032 (O_1032,N_14271,N_14948);
nand UO_1033 (O_1033,N_14251,N_14474);
nor UO_1034 (O_1034,N_14646,N_14624);
or UO_1035 (O_1035,N_14472,N_14739);
nand UO_1036 (O_1036,N_14565,N_14790);
nor UO_1037 (O_1037,N_14927,N_14262);
nand UO_1038 (O_1038,N_14669,N_14434);
and UO_1039 (O_1039,N_14312,N_14815);
and UO_1040 (O_1040,N_14606,N_14276);
or UO_1041 (O_1041,N_14918,N_14761);
nand UO_1042 (O_1042,N_14702,N_14256);
and UO_1043 (O_1043,N_14833,N_14569);
nor UO_1044 (O_1044,N_14725,N_14474);
nor UO_1045 (O_1045,N_14389,N_14351);
nor UO_1046 (O_1046,N_14772,N_14339);
and UO_1047 (O_1047,N_14653,N_14598);
nand UO_1048 (O_1048,N_14894,N_14827);
and UO_1049 (O_1049,N_14478,N_14361);
nand UO_1050 (O_1050,N_14463,N_14930);
nor UO_1051 (O_1051,N_14813,N_14724);
or UO_1052 (O_1052,N_14753,N_14827);
or UO_1053 (O_1053,N_14401,N_14689);
or UO_1054 (O_1054,N_14435,N_14854);
and UO_1055 (O_1055,N_14579,N_14395);
and UO_1056 (O_1056,N_14963,N_14580);
nand UO_1057 (O_1057,N_14650,N_14282);
nand UO_1058 (O_1058,N_14677,N_14744);
nand UO_1059 (O_1059,N_14477,N_14958);
nor UO_1060 (O_1060,N_14387,N_14929);
nor UO_1061 (O_1061,N_14806,N_14758);
and UO_1062 (O_1062,N_14816,N_14622);
and UO_1063 (O_1063,N_14626,N_14722);
and UO_1064 (O_1064,N_14568,N_14582);
nand UO_1065 (O_1065,N_14596,N_14901);
and UO_1066 (O_1066,N_14931,N_14505);
and UO_1067 (O_1067,N_14577,N_14860);
nor UO_1068 (O_1068,N_14660,N_14671);
nand UO_1069 (O_1069,N_14863,N_14989);
nand UO_1070 (O_1070,N_14345,N_14582);
nor UO_1071 (O_1071,N_14500,N_14669);
or UO_1072 (O_1072,N_14446,N_14757);
xor UO_1073 (O_1073,N_14691,N_14325);
xor UO_1074 (O_1074,N_14903,N_14673);
and UO_1075 (O_1075,N_14676,N_14811);
nand UO_1076 (O_1076,N_14426,N_14813);
nor UO_1077 (O_1077,N_14290,N_14851);
nand UO_1078 (O_1078,N_14603,N_14915);
nor UO_1079 (O_1079,N_14924,N_14542);
and UO_1080 (O_1080,N_14988,N_14335);
nor UO_1081 (O_1081,N_14752,N_14747);
nor UO_1082 (O_1082,N_14285,N_14956);
nand UO_1083 (O_1083,N_14489,N_14356);
nand UO_1084 (O_1084,N_14398,N_14476);
and UO_1085 (O_1085,N_14964,N_14714);
nand UO_1086 (O_1086,N_14644,N_14362);
nand UO_1087 (O_1087,N_14930,N_14912);
or UO_1088 (O_1088,N_14953,N_14970);
and UO_1089 (O_1089,N_14989,N_14682);
nor UO_1090 (O_1090,N_14617,N_14595);
or UO_1091 (O_1091,N_14871,N_14661);
or UO_1092 (O_1092,N_14342,N_14762);
and UO_1093 (O_1093,N_14490,N_14815);
xor UO_1094 (O_1094,N_14766,N_14307);
nor UO_1095 (O_1095,N_14967,N_14672);
nand UO_1096 (O_1096,N_14362,N_14818);
nor UO_1097 (O_1097,N_14498,N_14849);
nor UO_1098 (O_1098,N_14470,N_14947);
nand UO_1099 (O_1099,N_14864,N_14897);
nor UO_1100 (O_1100,N_14497,N_14402);
nor UO_1101 (O_1101,N_14885,N_14364);
or UO_1102 (O_1102,N_14780,N_14290);
nand UO_1103 (O_1103,N_14645,N_14862);
and UO_1104 (O_1104,N_14751,N_14996);
or UO_1105 (O_1105,N_14649,N_14508);
and UO_1106 (O_1106,N_14411,N_14365);
nand UO_1107 (O_1107,N_14544,N_14856);
and UO_1108 (O_1108,N_14457,N_14357);
or UO_1109 (O_1109,N_14407,N_14890);
nor UO_1110 (O_1110,N_14892,N_14572);
nor UO_1111 (O_1111,N_14282,N_14855);
nor UO_1112 (O_1112,N_14583,N_14403);
and UO_1113 (O_1113,N_14846,N_14285);
and UO_1114 (O_1114,N_14641,N_14780);
nor UO_1115 (O_1115,N_14299,N_14965);
and UO_1116 (O_1116,N_14500,N_14803);
and UO_1117 (O_1117,N_14685,N_14844);
nor UO_1118 (O_1118,N_14319,N_14571);
nor UO_1119 (O_1119,N_14518,N_14565);
and UO_1120 (O_1120,N_14435,N_14471);
or UO_1121 (O_1121,N_14861,N_14347);
and UO_1122 (O_1122,N_14667,N_14522);
nor UO_1123 (O_1123,N_14663,N_14461);
nor UO_1124 (O_1124,N_14369,N_14441);
and UO_1125 (O_1125,N_14520,N_14250);
or UO_1126 (O_1126,N_14594,N_14727);
or UO_1127 (O_1127,N_14523,N_14297);
nor UO_1128 (O_1128,N_14928,N_14463);
or UO_1129 (O_1129,N_14790,N_14960);
nor UO_1130 (O_1130,N_14694,N_14865);
or UO_1131 (O_1131,N_14896,N_14816);
nor UO_1132 (O_1132,N_14984,N_14270);
and UO_1133 (O_1133,N_14330,N_14995);
nand UO_1134 (O_1134,N_14926,N_14478);
or UO_1135 (O_1135,N_14693,N_14576);
and UO_1136 (O_1136,N_14846,N_14917);
and UO_1137 (O_1137,N_14513,N_14993);
nand UO_1138 (O_1138,N_14695,N_14503);
or UO_1139 (O_1139,N_14932,N_14601);
or UO_1140 (O_1140,N_14345,N_14738);
and UO_1141 (O_1141,N_14276,N_14623);
nor UO_1142 (O_1142,N_14407,N_14949);
nand UO_1143 (O_1143,N_14978,N_14876);
nor UO_1144 (O_1144,N_14495,N_14830);
nand UO_1145 (O_1145,N_14607,N_14280);
nand UO_1146 (O_1146,N_14887,N_14706);
nor UO_1147 (O_1147,N_14603,N_14439);
nor UO_1148 (O_1148,N_14822,N_14281);
and UO_1149 (O_1149,N_14552,N_14279);
and UO_1150 (O_1150,N_14742,N_14550);
and UO_1151 (O_1151,N_14474,N_14543);
or UO_1152 (O_1152,N_14312,N_14978);
nor UO_1153 (O_1153,N_14512,N_14530);
nand UO_1154 (O_1154,N_14263,N_14828);
nand UO_1155 (O_1155,N_14876,N_14991);
or UO_1156 (O_1156,N_14581,N_14710);
and UO_1157 (O_1157,N_14953,N_14589);
nor UO_1158 (O_1158,N_14923,N_14849);
or UO_1159 (O_1159,N_14523,N_14867);
or UO_1160 (O_1160,N_14535,N_14846);
or UO_1161 (O_1161,N_14748,N_14853);
nand UO_1162 (O_1162,N_14634,N_14285);
or UO_1163 (O_1163,N_14551,N_14270);
or UO_1164 (O_1164,N_14677,N_14978);
or UO_1165 (O_1165,N_14669,N_14517);
and UO_1166 (O_1166,N_14478,N_14252);
and UO_1167 (O_1167,N_14391,N_14528);
and UO_1168 (O_1168,N_14994,N_14818);
or UO_1169 (O_1169,N_14575,N_14879);
nand UO_1170 (O_1170,N_14700,N_14506);
and UO_1171 (O_1171,N_14463,N_14794);
nand UO_1172 (O_1172,N_14925,N_14992);
nand UO_1173 (O_1173,N_14282,N_14506);
nand UO_1174 (O_1174,N_14656,N_14848);
nand UO_1175 (O_1175,N_14505,N_14346);
and UO_1176 (O_1176,N_14953,N_14762);
and UO_1177 (O_1177,N_14504,N_14759);
nand UO_1178 (O_1178,N_14836,N_14429);
nor UO_1179 (O_1179,N_14367,N_14599);
nor UO_1180 (O_1180,N_14704,N_14488);
and UO_1181 (O_1181,N_14733,N_14953);
nand UO_1182 (O_1182,N_14602,N_14436);
nand UO_1183 (O_1183,N_14255,N_14292);
and UO_1184 (O_1184,N_14821,N_14270);
nand UO_1185 (O_1185,N_14254,N_14932);
nand UO_1186 (O_1186,N_14752,N_14390);
or UO_1187 (O_1187,N_14413,N_14327);
nor UO_1188 (O_1188,N_14990,N_14670);
nor UO_1189 (O_1189,N_14613,N_14399);
nor UO_1190 (O_1190,N_14511,N_14583);
and UO_1191 (O_1191,N_14435,N_14254);
nor UO_1192 (O_1192,N_14434,N_14605);
or UO_1193 (O_1193,N_14368,N_14665);
or UO_1194 (O_1194,N_14583,N_14882);
nand UO_1195 (O_1195,N_14923,N_14317);
and UO_1196 (O_1196,N_14423,N_14604);
or UO_1197 (O_1197,N_14881,N_14496);
and UO_1198 (O_1198,N_14908,N_14647);
nand UO_1199 (O_1199,N_14490,N_14907);
and UO_1200 (O_1200,N_14329,N_14812);
and UO_1201 (O_1201,N_14366,N_14804);
and UO_1202 (O_1202,N_14811,N_14783);
nand UO_1203 (O_1203,N_14596,N_14362);
nor UO_1204 (O_1204,N_14834,N_14927);
nor UO_1205 (O_1205,N_14397,N_14350);
or UO_1206 (O_1206,N_14985,N_14421);
nor UO_1207 (O_1207,N_14304,N_14893);
nor UO_1208 (O_1208,N_14393,N_14804);
nand UO_1209 (O_1209,N_14398,N_14644);
nand UO_1210 (O_1210,N_14464,N_14596);
or UO_1211 (O_1211,N_14977,N_14383);
nor UO_1212 (O_1212,N_14885,N_14610);
or UO_1213 (O_1213,N_14776,N_14913);
and UO_1214 (O_1214,N_14675,N_14627);
and UO_1215 (O_1215,N_14615,N_14365);
nand UO_1216 (O_1216,N_14539,N_14497);
nand UO_1217 (O_1217,N_14802,N_14768);
nand UO_1218 (O_1218,N_14327,N_14550);
nor UO_1219 (O_1219,N_14682,N_14755);
and UO_1220 (O_1220,N_14936,N_14824);
or UO_1221 (O_1221,N_14987,N_14301);
nand UO_1222 (O_1222,N_14477,N_14432);
nand UO_1223 (O_1223,N_14413,N_14853);
nand UO_1224 (O_1224,N_14621,N_14495);
nand UO_1225 (O_1225,N_14544,N_14294);
and UO_1226 (O_1226,N_14496,N_14318);
nor UO_1227 (O_1227,N_14695,N_14391);
nand UO_1228 (O_1228,N_14501,N_14504);
and UO_1229 (O_1229,N_14839,N_14535);
nand UO_1230 (O_1230,N_14494,N_14465);
or UO_1231 (O_1231,N_14899,N_14667);
and UO_1232 (O_1232,N_14409,N_14426);
or UO_1233 (O_1233,N_14384,N_14819);
or UO_1234 (O_1234,N_14893,N_14840);
nor UO_1235 (O_1235,N_14942,N_14826);
and UO_1236 (O_1236,N_14607,N_14440);
nand UO_1237 (O_1237,N_14823,N_14346);
nor UO_1238 (O_1238,N_14853,N_14785);
and UO_1239 (O_1239,N_14901,N_14260);
or UO_1240 (O_1240,N_14534,N_14404);
nand UO_1241 (O_1241,N_14564,N_14395);
and UO_1242 (O_1242,N_14371,N_14913);
nor UO_1243 (O_1243,N_14721,N_14383);
nand UO_1244 (O_1244,N_14260,N_14711);
or UO_1245 (O_1245,N_14261,N_14826);
nor UO_1246 (O_1246,N_14651,N_14602);
nand UO_1247 (O_1247,N_14689,N_14724);
or UO_1248 (O_1248,N_14704,N_14853);
or UO_1249 (O_1249,N_14633,N_14867);
nor UO_1250 (O_1250,N_14786,N_14916);
and UO_1251 (O_1251,N_14612,N_14633);
nor UO_1252 (O_1252,N_14447,N_14266);
and UO_1253 (O_1253,N_14722,N_14973);
or UO_1254 (O_1254,N_14733,N_14277);
nor UO_1255 (O_1255,N_14645,N_14340);
or UO_1256 (O_1256,N_14297,N_14444);
nor UO_1257 (O_1257,N_14578,N_14605);
nand UO_1258 (O_1258,N_14591,N_14677);
or UO_1259 (O_1259,N_14910,N_14335);
nor UO_1260 (O_1260,N_14493,N_14716);
nor UO_1261 (O_1261,N_14916,N_14276);
and UO_1262 (O_1262,N_14628,N_14928);
nand UO_1263 (O_1263,N_14664,N_14635);
nor UO_1264 (O_1264,N_14779,N_14954);
nand UO_1265 (O_1265,N_14509,N_14828);
or UO_1266 (O_1266,N_14896,N_14367);
nor UO_1267 (O_1267,N_14925,N_14454);
and UO_1268 (O_1268,N_14794,N_14380);
or UO_1269 (O_1269,N_14293,N_14616);
or UO_1270 (O_1270,N_14736,N_14669);
nand UO_1271 (O_1271,N_14436,N_14657);
nor UO_1272 (O_1272,N_14694,N_14295);
nand UO_1273 (O_1273,N_14480,N_14310);
nand UO_1274 (O_1274,N_14872,N_14674);
nor UO_1275 (O_1275,N_14944,N_14462);
and UO_1276 (O_1276,N_14358,N_14638);
and UO_1277 (O_1277,N_14339,N_14985);
nand UO_1278 (O_1278,N_14611,N_14925);
or UO_1279 (O_1279,N_14599,N_14832);
and UO_1280 (O_1280,N_14702,N_14678);
and UO_1281 (O_1281,N_14837,N_14531);
nor UO_1282 (O_1282,N_14558,N_14346);
or UO_1283 (O_1283,N_14710,N_14453);
nand UO_1284 (O_1284,N_14798,N_14359);
nor UO_1285 (O_1285,N_14662,N_14269);
and UO_1286 (O_1286,N_14485,N_14719);
nand UO_1287 (O_1287,N_14302,N_14956);
and UO_1288 (O_1288,N_14685,N_14506);
nand UO_1289 (O_1289,N_14266,N_14692);
nor UO_1290 (O_1290,N_14428,N_14741);
and UO_1291 (O_1291,N_14750,N_14669);
nand UO_1292 (O_1292,N_14956,N_14492);
nor UO_1293 (O_1293,N_14318,N_14972);
nand UO_1294 (O_1294,N_14332,N_14502);
or UO_1295 (O_1295,N_14860,N_14321);
or UO_1296 (O_1296,N_14947,N_14526);
or UO_1297 (O_1297,N_14691,N_14592);
nand UO_1298 (O_1298,N_14615,N_14777);
and UO_1299 (O_1299,N_14777,N_14372);
nor UO_1300 (O_1300,N_14474,N_14648);
nand UO_1301 (O_1301,N_14577,N_14951);
nand UO_1302 (O_1302,N_14691,N_14852);
nor UO_1303 (O_1303,N_14932,N_14461);
nor UO_1304 (O_1304,N_14617,N_14720);
or UO_1305 (O_1305,N_14483,N_14485);
nand UO_1306 (O_1306,N_14620,N_14863);
or UO_1307 (O_1307,N_14586,N_14674);
and UO_1308 (O_1308,N_14267,N_14473);
nor UO_1309 (O_1309,N_14950,N_14842);
and UO_1310 (O_1310,N_14478,N_14721);
or UO_1311 (O_1311,N_14498,N_14352);
or UO_1312 (O_1312,N_14443,N_14880);
nand UO_1313 (O_1313,N_14423,N_14803);
nor UO_1314 (O_1314,N_14626,N_14706);
or UO_1315 (O_1315,N_14773,N_14946);
nor UO_1316 (O_1316,N_14886,N_14750);
nand UO_1317 (O_1317,N_14261,N_14877);
nor UO_1318 (O_1318,N_14826,N_14858);
and UO_1319 (O_1319,N_14546,N_14600);
nand UO_1320 (O_1320,N_14309,N_14658);
or UO_1321 (O_1321,N_14492,N_14886);
nor UO_1322 (O_1322,N_14842,N_14525);
nand UO_1323 (O_1323,N_14686,N_14705);
nor UO_1324 (O_1324,N_14920,N_14918);
or UO_1325 (O_1325,N_14378,N_14698);
or UO_1326 (O_1326,N_14595,N_14728);
nand UO_1327 (O_1327,N_14840,N_14980);
or UO_1328 (O_1328,N_14579,N_14348);
or UO_1329 (O_1329,N_14343,N_14792);
nand UO_1330 (O_1330,N_14419,N_14436);
and UO_1331 (O_1331,N_14286,N_14422);
or UO_1332 (O_1332,N_14380,N_14277);
and UO_1333 (O_1333,N_14662,N_14307);
nand UO_1334 (O_1334,N_14926,N_14501);
and UO_1335 (O_1335,N_14965,N_14653);
nor UO_1336 (O_1336,N_14655,N_14506);
xnor UO_1337 (O_1337,N_14409,N_14456);
or UO_1338 (O_1338,N_14277,N_14788);
and UO_1339 (O_1339,N_14714,N_14543);
or UO_1340 (O_1340,N_14897,N_14487);
nand UO_1341 (O_1341,N_14635,N_14261);
and UO_1342 (O_1342,N_14733,N_14298);
or UO_1343 (O_1343,N_14260,N_14795);
or UO_1344 (O_1344,N_14294,N_14470);
nand UO_1345 (O_1345,N_14726,N_14570);
nand UO_1346 (O_1346,N_14558,N_14983);
nand UO_1347 (O_1347,N_14268,N_14266);
nor UO_1348 (O_1348,N_14678,N_14750);
nand UO_1349 (O_1349,N_14445,N_14370);
nand UO_1350 (O_1350,N_14255,N_14979);
nand UO_1351 (O_1351,N_14508,N_14790);
and UO_1352 (O_1352,N_14312,N_14660);
and UO_1353 (O_1353,N_14271,N_14523);
or UO_1354 (O_1354,N_14534,N_14287);
nand UO_1355 (O_1355,N_14733,N_14790);
nor UO_1356 (O_1356,N_14320,N_14467);
and UO_1357 (O_1357,N_14624,N_14904);
nor UO_1358 (O_1358,N_14780,N_14473);
or UO_1359 (O_1359,N_14257,N_14411);
and UO_1360 (O_1360,N_14282,N_14821);
or UO_1361 (O_1361,N_14783,N_14557);
nand UO_1362 (O_1362,N_14916,N_14316);
and UO_1363 (O_1363,N_14898,N_14510);
nand UO_1364 (O_1364,N_14781,N_14800);
or UO_1365 (O_1365,N_14616,N_14925);
or UO_1366 (O_1366,N_14344,N_14520);
nand UO_1367 (O_1367,N_14455,N_14878);
xor UO_1368 (O_1368,N_14956,N_14605);
nor UO_1369 (O_1369,N_14570,N_14264);
nand UO_1370 (O_1370,N_14377,N_14881);
nand UO_1371 (O_1371,N_14488,N_14343);
nand UO_1372 (O_1372,N_14396,N_14919);
nor UO_1373 (O_1373,N_14784,N_14668);
nand UO_1374 (O_1374,N_14751,N_14830);
or UO_1375 (O_1375,N_14850,N_14475);
or UO_1376 (O_1376,N_14673,N_14908);
nand UO_1377 (O_1377,N_14832,N_14702);
nand UO_1378 (O_1378,N_14338,N_14384);
or UO_1379 (O_1379,N_14492,N_14793);
or UO_1380 (O_1380,N_14527,N_14534);
and UO_1381 (O_1381,N_14612,N_14666);
nand UO_1382 (O_1382,N_14571,N_14759);
nor UO_1383 (O_1383,N_14428,N_14298);
nand UO_1384 (O_1384,N_14343,N_14530);
nand UO_1385 (O_1385,N_14667,N_14911);
and UO_1386 (O_1386,N_14820,N_14940);
nand UO_1387 (O_1387,N_14952,N_14332);
and UO_1388 (O_1388,N_14920,N_14941);
or UO_1389 (O_1389,N_14658,N_14325);
and UO_1390 (O_1390,N_14847,N_14998);
nand UO_1391 (O_1391,N_14925,N_14631);
nand UO_1392 (O_1392,N_14863,N_14594);
nand UO_1393 (O_1393,N_14766,N_14638);
or UO_1394 (O_1394,N_14580,N_14946);
nand UO_1395 (O_1395,N_14376,N_14789);
or UO_1396 (O_1396,N_14909,N_14632);
nor UO_1397 (O_1397,N_14302,N_14769);
nor UO_1398 (O_1398,N_14286,N_14701);
or UO_1399 (O_1399,N_14547,N_14465);
and UO_1400 (O_1400,N_14307,N_14879);
and UO_1401 (O_1401,N_14281,N_14917);
or UO_1402 (O_1402,N_14828,N_14705);
or UO_1403 (O_1403,N_14684,N_14923);
nand UO_1404 (O_1404,N_14761,N_14399);
nor UO_1405 (O_1405,N_14582,N_14359);
or UO_1406 (O_1406,N_14675,N_14742);
nand UO_1407 (O_1407,N_14936,N_14966);
or UO_1408 (O_1408,N_14855,N_14876);
xor UO_1409 (O_1409,N_14830,N_14422);
and UO_1410 (O_1410,N_14914,N_14253);
nand UO_1411 (O_1411,N_14254,N_14560);
nor UO_1412 (O_1412,N_14824,N_14918);
and UO_1413 (O_1413,N_14414,N_14441);
and UO_1414 (O_1414,N_14755,N_14479);
or UO_1415 (O_1415,N_14556,N_14307);
nand UO_1416 (O_1416,N_14706,N_14250);
and UO_1417 (O_1417,N_14573,N_14320);
nor UO_1418 (O_1418,N_14525,N_14288);
or UO_1419 (O_1419,N_14602,N_14421);
and UO_1420 (O_1420,N_14730,N_14272);
nor UO_1421 (O_1421,N_14701,N_14827);
nand UO_1422 (O_1422,N_14995,N_14968);
nand UO_1423 (O_1423,N_14639,N_14621);
and UO_1424 (O_1424,N_14853,N_14400);
nand UO_1425 (O_1425,N_14311,N_14298);
nor UO_1426 (O_1426,N_14732,N_14636);
and UO_1427 (O_1427,N_14678,N_14397);
nor UO_1428 (O_1428,N_14827,N_14587);
or UO_1429 (O_1429,N_14323,N_14683);
nand UO_1430 (O_1430,N_14818,N_14625);
nand UO_1431 (O_1431,N_14609,N_14892);
nor UO_1432 (O_1432,N_14786,N_14572);
or UO_1433 (O_1433,N_14718,N_14892);
and UO_1434 (O_1434,N_14356,N_14672);
and UO_1435 (O_1435,N_14892,N_14915);
or UO_1436 (O_1436,N_14275,N_14887);
or UO_1437 (O_1437,N_14731,N_14638);
nor UO_1438 (O_1438,N_14429,N_14953);
nor UO_1439 (O_1439,N_14290,N_14775);
nor UO_1440 (O_1440,N_14828,N_14536);
nor UO_1441 (O_1441,N_14478,N_14632);
nand UO_1442 (O_1442,N_14678,N_14800);
nor UO_1443 (O_1443,N_14486,N_14265);
nor UO_1444 (O_1444,N_14937,N_14764);
and UO_1445 (O_1445,N_14535,N_14899);
or UO_1446 (O_1446,N_14702,N_14712);
and UO_1447 (O_1447,N_14946,N_14706);
or UO_1448 (O_1448,N_14278,N_14971);
and UO_1449 (O_1449,N_14512,N_14364);
and UO_1450 (O_1450,N_14910,N_14785);
or UO_1451 (O_1451,N_14466,N_14664);
or UO_1452 (O_1452,N_14978,N_14355);
or UO_1453 (O_1453,N_14568,N_14927);
or UO_1454 (O_1454,N_14500,N_14819);
and UO_1455 (O_1455,N_14287,N_14513);
nor UO_1456 (O_1456,N_14871,N_14750);
nor UO_1457 (O_1457,N_14336,N_14486);
nor UO_1458 (O_1458,N_14502,N_14795);
or UO_1459 (O_1459,N_14949,N_14339);
nor UO_1460 (O_1460,N_14413,N_14896);
nand UO_1461 (O_1461,N_14661,N_14345);
and UO_1462 (O_1462,N_14398,N_14444);
nor UO_1463 (O_1463,N_14836,N_14480);
nor UO_1464 (O_1464,N_14526,N_14445);
nand UO_1465 (O_1465,N_14939,N_14447);
and UO_1466 (O_1466,N_14531,N_14439);
and UO_1467 (O_1467,N_14490,N_14814);
nand UO_1468 (O_1468,N_14936,N_14958);
xor UO_1469 (O_1469,N_14849,N_14980);
nor UO_1470 (O_1470,N_14259,N_14702);
or UO_1471 (O_1471,N_14449,N_14495);
nor UO_1472 (O_1472,N_14695,N_14549);
or UO_1473 (O_1473,N_14619,N_14736);
and UO_1474 (O_1474,N_14565,N_14774);
and UO_1475 (O_1475,N_14525,N_14951);
and UO_1476 (O_1476,N_14623,N_14319);
nor UO_1477 (O_1477,N_14431,N_14485);
nand UO_1478 (O_1478,N_14343,N_14863);
and UO_1479 (O_1479,N_14269,N_14840);
nor UO_1480 (O_1480,N_14282,N_14446);
or UO_1481 (O_1481,N_14659,N_14402);
nor UO_1482 (O_1482,N_14933,N_14662);
or UO_1483 (O_1483,N_14775,N_14543);
or UO_1484 (O_1484,N_14274,N_14544);
nand UO_1485 (O_1485,N_14275,N_14905);
nor UO_1486 (O_1486,N_14972,N_14889);
nor UO_1487 (O_1487,N_14637,N_14723);
nor UO_1488 (O_1488,N_14876,N_14689);
or UO_1489 (O_1489,N_14803,N_14982);
nor UO_1490 (O_1490,N_14674,N_14784);
nand UO_1491 (O_1491,N_14568,N_14776);
or UO_1492 (O_1492,N_14445,N_14328);
nand UO_1493 (O_1493,N_14284,N_14612);
or UO_1494 (O_1494,N_14286,N_14550);
or UO_1495 (O_1495,N_14558,N_14329);
and UO_1496 (O_1496,N_14510,N_14654);
xnor UO_1497 (O_1497,N_14881,N_14643);
nor UO_1498 (O_1498,N_14999,N_14835);
and UO_1499 (O_1499,N_14846,N_14449);
nand UO_1500 (O_1500,N_14885,N_14670);
nand UO_1501 (O_1501,N_14860,N_14997);
nand UO_1502 (O_1502,N_14781,N_14850);
or UO_1503 (O_1503,N_14594,N_14788);
nand UO_1504 (O_1504,N_14841,N_14298);
and UO_1505 (O_1505,N_14441,N_14538);
nand UO_1506 (O_1506,N_14816,N_14812);
nor UO_1507 (O_1507,N_14931,N_14280);
or UO_1508 (O_1508,N_14810,N_14438);
nand UO_1509 (O_1509,N_14586,N_14386);
nand UO_1510 (O_1510,N_14428,N_14345);
or UO_1511 (O_1511,N_14442,N_14807);
nand UO_1512 (O_1512,N_14763,N_14987);
nor UO_1513 (O_1513,N_14842,N_14794);
nand UO_1514 (O_1514,N_14364,N_14435);
and UO_1515 (O_1515,N_14852,N_14948);
and UO_1516 (O_1516,N_14720,N_14907);
nand UO_1517 (O_1517,N_14453,N_14263);
or UO_1518 (O_1518,N_14523,N_14689);
or UO_1519 (O_1519,N_14819,N_14759);
nor UO_1520 (O_1520,N_14439,N_14915);
nor UO_1521 (O_1521,N_14865,N_14618);
and UO_1522 (O_1522,N_14711,N_14442);
or UO_1523 (O_1523,N_14250,N_14917);
nand UO_1524 (O_1524,N_14433,N_14643);
nand UO_1525 (O_1525,N_14277,N_14759);
nor UO_1526 (O_1526,N_14410,N_14941);
and UO_1527 (O_1527,N_14927,N_14584);
nand UO_1528 (O_1528,N_14966,N_14260);
or UO_1529 (O_1529,N_14253,N_14488);
and UO_1530 (O_1530,N_14720,N_14643);
or UO_1531 (O_1531,N_14586,N_14877);
or UO_1532 (O_1532,N_14279,N_14626);
nor UO_1533 (O_1533,N_14784,N_14673);
or UO_1534 (O_1534,N_14373,N_14549);
and UO_1535 (O_1535,N_14920,N_14656);
or UO_1536 (O_1536,N_14841,N_14504);
and UO_1537 (O_1537,N_14444,N_14458);
or UO_1538 (O_1538,N_14736,N_14531);
nand UO_1539 (O_1539,N_14962,N_14819);
nor UO_1540 (O_1540,N_14661,N_14406);
or UO_1541 (O_1541,N_14318,N_14390);
or UO_1542 (O_1542,N_14737,N_14281);
nand UO_1543 (O_1543,N_14559,N_14701);
and UO_1544 (O_1544,N_14987,N_14837);
and UO_1545 (O_1545,N_14415,N_14746);
nor UO_1546 (O_1546,N_14556,N_14388);
or UO_1547 (O_1547,N_14819,N_14868);
or UO_1548 (O_1548,N_14640,N_14742);
nor UO_1549 (O_1549,N_14612,N_14366);
nor UO_1550 (O_1550,N_14908,N_14857);
nor UO_1551 (O_1551,N_14454,N_14355);
nand UO_1552 (O_1552,N_14523,N_14376);
nand UO_1553 (O_1553,N_14992,N_14743);
nand UO_1554 (O_1554,N_14777,N_14359);
nor UO_1555 (O_1555,N_14544,N_14345);
or UO_1556 (O_1556,N_14628,N_14753);
or UO_1557 (O_1557,N_14889,N_14904);
nor UO_1558 (O_1558,N_14305,N_14401);
and UO_1559 (O_1559,N_14269,N_14349);
or UO_1560 (O_1560,N_14667,N_14627);
and UO_1561 (O_1561,N_14599,N_14666);
or UO_1562 (O_1562,N_14990,N_14387);
nor UO_1563 (O_1563,N_14308,N_14276);
or UO_1564 (O_1564,N_14256,N_14898);
nand UO_1565 (O_1565,N_14846,N_14789);
nand UO_1566 (O_1566,N_14374,N_14694);
nand UO_1567 (O_1567,N_14353,N_14668);
or UO_1568 (O_1568,N_14648,N_14918);
nor UO_1569 (O_1569,N_14570,N_14290);
and UO_1570 (O_1570,N_14471,N_14340);
nor UO_1571 (O_1571,N_14500,N_14609);
or UO_1572 (O_1572,N_14458,N_14396);
nor UO_1573 (O_1573,N_14965,N_14649);
nor UO_1574 (O_1574,N_14963,N_14719);
nand UO_1575 (O_1575,N_14663,N_14431);
nor UO_1576 (O_1576,N_14612,N_14569);
and UO_1577 (O_1577,N_14985,N_14966);
nand UO_1578 (O_1578,N_14681,N_14597);
and UO_1579 (O_1579,N_14787,N_14349);
nor UO_1580 (O_1580,N_14528,N_14892);
nor UO_1581 (O_1581,N_14556,N_14722);
or UO_1582 (O_1582,N_14435,N_14896);
nor UO_1583 (O_1583,N_14346,N_14289);
or UO_1584 (O_1584,N_14961,N_14501);
or UO_1585 (O_1585,N_14921,N_14618);
nand UO_1586 (O_1586,N_14686,N_14683);
or UO_1587 (O_1587,N_14446,N_14899);
and UO_1588 (O_1588,N_14609,N_14931);
and UO_1589 (O_1589,N_14511,N_14619);
and UO_1590 (O_1590,N_14254,N_14706);
and UO_1591 (O_1591,N_14999,N_14596);
nor UO_1592 (O_1592,N_14675,N_14917);
nand UO_1593 (O_1593,N_14794,N_14636);
or UO_1594 (O_1594,N_14698,N_14682);
and UO_1595 (O_1595,N_14815,N_14798);
or UO_1596 (O_1596,N_14941,N_14994);
nand UO_1597 (O_1597,N_14453,N_14851);
nand UO_1598 (O_1598,N_14691,N_14521);
nand UO_1599 (O_1599,N_14829,N_14642);
and UO_1600 (O_1600,N_14593,N_14739);
nand UO_1601 (O_1601,N_14805,N_14615);
nor UO_1602 (O_1602,N_14733,N_14793);
nor UO_1603 (O_1603,N_14925,N_14558);
nand UO_1604 (O_1604,N_14395,N_14603);
nor UO_1605 (O_1605,N_14270,N_14942);
or UO_1606 (O_1606,N_14257,N_14945);
nand UO_1607 (O_1607,N_14692,N_14739);
or UO_1608 (O_1608,N_14269,N_14813);
and UO_1609 (O_1609,N_14644,N_14837);
or UO_1610 (O_1610,N_14824,N_14949);
and UO_1611 (O_1611,N_14425,N_14373);
nor UO_1612 (O_1612,N_14618,N_14412);
and UO_1613 (O_1613,N_14881,N_14658);
and UO_1614 (O_1614,N_14491,N_14482);
nand UO_1615 (O_1615,N_14327,N_14909);
and UO_1616 (O_1616,N_14423,N_14562);
and UO_1617 (O_1617,N_14536,N_14723);
and UO_1618 (O_1618,N_14739,N_14780);
and UO_1619 (O_1619,N_14472,N_14255);
xnor UO_1620 (O_1620,N_14622,N_14311);
and UO_1621 (O_1621,N_14968,N_14686);
nor UO_1622 (O_1622,N_14866,N_14382);
or UO_1623 (O_1623,N_14748,N_14383);
nand UO_1624 (O_1624,N_14752,N_14614);
and UO_1625 (O_1625,N_14763,N_14594);
or UO_1626 (O_1626,N_14677,N_14339);
or UO_1627 (O_1627,N_14879,N_14689);
and UO_1628 (O_1628,N_14765,N_14794);
nor UO_1629 (O_1629,N_14327,N_14549);
nor UO_1630 (O_1630,N_14528,N_14990);
or UO_1631 (O_1631,N_14919,N_14305);
nor UO_1632 (O_1632,N_14877,N_14252);
or UO_1633 (O_1633,N_14796,N_14440);
nand UO_1634 (O_1634,N_14661,N_14564);
nand UO_1635 (O_1635,N_14873,N_14573);
or UO_1636 (O_1636,N_14548,N_14693);
and UO_1637 (O_1637,N_14292,N_14442);
and UO_1638 (O_1638,N_14810,N_14497);
nand UO_1639 (O_1639,N_14545,N_14384);
and UO_1640 (O_1640,N_14862,N_14331);
and UO_1641 (O_1641,N_14490,N_14740);
and UO_1642 (O_1642,N_14341,N_14819);
nor UO_1643 (O_1643,N_14262,N_14578);
and UO_1644 (O_1644,N_14343,N_14909);
or UO_1645 (O_1645,N_14529,N_14600);
xor UO_1646 (O_1646,N_14967,N_14605);
nand UO_1647 (O_1647,N_14250,N_14705);
nor UO_1648 (O_1648,N_14417,N_14820);
and UO_1649 (O_1649,N_14518,N_14834);
or UO_1650 (O_1650,N_14641,N_14600);
nor UO_1651 (O_1651,N_14943,N_14959);
nand UO_1652 (O_1652,N_14765,N_14777);
and UO_1653 (O_1653,N_14701,N_14774);
and UO_1654 (O_1654,N_14733,N_14456);
nor UO_1655 (O_1655,N_14262,N_14309);
nand UO_1656 (O_1656,N_14684,N_14564);
nand UO_1657 (O_1657,N_14525,N_14336);
nand UO_1658 (O_1658,N_14521,N_14416);
or UO_1659 (O_1659,N_14470,N_14539);
nor UO_1660 (O_1660,N_14618,N_14946);
nand UO_1661 (O_1661,N_14724,N_14308);
xor UO_1662 (O_1662,N_14930,N_14867);
nand UO_1663 (O_1663,N_14580,N_14673);
nand UO_1664 (O_1664,N_14703,N_14496);
or UO_1665 (O_1665,N_14495,N_14262);
nor UO_1666 (O_1666,N_14377,N_14962);
nor UO_1667 (O_1667,N_14919,N_14861);
nor UO_1668 (O_1668,N_14862,N_14751);
and UO_1669 (O_1669,N_14758,N_14741);
nand UO_1670 (O_1670,N_14866,N_14476);
nor UO_1671 (O_1671,N_14256,N_14422);
or UO_1672 (O_1672,N_14905,N_14273);
and UO_1673 (O_1673,N_14273,N_14864);
nor UO_1674 (O_1674,N_14487,N_14796);
or UO_1675 (O_1675,N_14489,N_14410);
and UO_1676 (O_1676,N_14457,N_14786);
nand UO_1677 (O_1677,N_14853,N_14649);
and UO_1678 (O_1678,N_14828,N_14318);
or UO_1679 (O_1679,N_14619,N_14829);
and UO_1680 (O_1680,N_14988,N_14257);
nor UO_1681 (O_1681,N_14938,N_14998);
or UO_1682 (O_1682,N_14999,N_14438);
xnor UO_1683 (O_1683,N_14697,N_14420);
and UO_1684 (O_1684,N_14539,N_14853);
nor UO_1685 (O_1685,N_14711,N_14624);
and UO_1686 (O_1686,N_14933,N_14994);
or UO_1687 (O_1687,N_14883,N_14648);
and UO_1688 (O_1688,N_14335,N_14565);
and UO_1689 (O_1689,N_14275,N_14563);
nand UO_1690 (O_1690,N_14365,N_14341);
and UO_1691 (O_1691,N_14515,N_14947);
nand UO_1692 (O_1692,N_14516,N_14577);
nand UO_1693 (O_1693,N_14352,N_14262);
and UO_1694 (O_1694,N_14268,N_14618);
or UO_1695 (O_1695,N_14294,N_14425);
or UO_1696 (O_1696,N_14578,N_14461);
or UO_1697 (O_1697,N_14666,N_14476);
nor UO_1698 (O_1698,N_14377,N_14842);
nand UO_1699 (O_1699,N_14495,N_14966);
and UO_1700 (O_1700,N_14274,N_14537);
and UO_1701 (O_1701,N_14355,N_14974);
and UO_1702 (O_1702,N_14290,N_14299);
nand UO_1703 (O_1703,N_14413,N_14606);
nand UO_1704 (O_1704,N_14537,N_14699);
or UO_1705 (O_1705,N_14425,N_14839);
nor UO_1706 (O_1706,N_14991,N_14426);
and UO_1707 (O_1707,N_14397,N_14579);
nor UO_1708 (O_1708,N_14829,N_14751);
nor UO_1709 (O_1709,N_14297,N_14979);
nor UO_1710 (O_1710,N_14266,N_14857);
xor UO_1711 (O_1711,N_14296,N_14688);
nor UO_1712 (O_1712,N_14737,N_14706);
nand UO_1713 (O_1713,N_14671,N_14805);
or UO_1714 (O_1714,N_14302,N_14679);
and UO_1715 (O_1715,N_14308,N_14425);
and UO_1716 (O_1716,N_14374,N_14985);
nor UO_1717 (O_1717,N_14713,N_14278);
nor UO_1718 (O_1718,N_14368,N_14632);
nor UO_1719 (O_1719,N_14830,N_14521);
or UO_1720 (O_1720,N_14513,N_14809);
and UO_1721 (O_1721,N_14564,N_14794);
or UO_1722 (O_1722,N_14409,N_14778);
nand UO_1723 (O_1723,N_14394,N_14812);
or UO_1724 (O_1724,N_14753,N_14294);
nor UO_1725 (O_1725,N_14949,N_14479);
or UO_1726 (O_1726,N_14961,N_14293);
or UO_1727 (O_1727,N_14829,N_14986);
nor UO_1728 (O_1728,N_14980,N_14752);
and UO_1729 (O_1729,N_14454,N_14718);
nor UO_1730 (O_1730,N_14728,N_14257);
or UO_1731 (O_1731,N_14459,N_14601);
nand UO_1732 (O_1732,N_14431,N_14936);
and UO_1733 (O_1733,N_14507,N_14881);
nand UO_1734 (O_1734,N_14330,N_14685);
nor UO_1735 (O_1735,N_14475,N_14682);
nor UO_1736 (O_1736,N_14649,N_14348);
and UO_1737 (O_1737,N_14354,N_14427);
nand UO_1738 (O_1738,N_14747,N_14480);
nand UO_1739 (O_1739,N_14926,N_14824);
nor UO_1740 (O_1740,N_14838,N_14466);
or UO_1741 (O_1741,N_14260,N_14973);
nand UO_1742 (O_1742,N_14254,N_14262);
and UO_1743 (O_1743,N_14332,N_14670);
or UO_1744 (O_1744,N_14458,N_14291);
nor UO_1745 (O_1745,N_14390,N_14429);
or UO_1746 (O_1746,N_14338,N_14420);
and UO_1747 (O_1747,N_14636,N_14489);
and UO_1748 (O_1748,N_14796,N_14651);
nand UO_1749 (O_1749,N_14624,N_14471);
nor UO_1750 (O_1750,N_14337,N_14906);
and UO_1751 (O_1751,N_14329,N_14663);
and UO_1752 (O_1752,N_14540,N_14372);
and UO_1753 (O_1753,N_14358,N_14895);
nor UO_1754 (O_1754,N_14613,N_14459);
nand UO_1755 (O_1755,N_14252,N_14662);
and UO_1756 (O_1756,N_14827,N_14274);
nor UO_1757 (O_1757,N_14439,N_14677);
nand UO_1758 (O_1758,N_14556,N_14360);
and UO_1759 (O_1759,N_14378,N_14264);
nand UO_1760 (O_1760,N_14915,N_14944);
and UO_1761 (O_1761,N_14987,N_14372);
nand UO_1762 (O_1762,N_14963,N_14574);
or UO_1763 (O_1763,N_14944,N_14359);
nand UO_1764 (O_1764,N_14437,N_14592);
nor UO_1765 (O_1765,N_14933,N_14433);
and UO_1766 (O_1766,N_14706,N_14671);
and UO_1767 (O_1767,N_14479,N_14825);
and UO_1768 (O_1768,N_14456,N_14280);
nand UO_1769 (O_1769,N_14689,N_14280);
or UO_1770 (O_1770,N_14756,N_14842);
or UO_1771 (O_1771,N_14419,N_14590);
or UO_1772 (O_1772,N_14306,N_14689);
nand UO_1773 (O_1773,N_14306,N_14919);
or UO_1774 (O_1774,N_14702,N_14279);
or UO_1775 (O_1775,N_14532,N_14805);
nor UO_1776 (O_1776,N_14390,N_14812);
or UO_1777 (O_1777,N_14498,N_14889);
nor UO_1778 (O_1778,N_14551,N_14817);
nand UO_1779 (O_1779,N_14938,N_14918);
or UO_1780 (O_1780,N_14499,N_14444);
nand UO_1781 (O_1781,N_14710,N_14421);
and UO_1782 (O_1782,N_14592,N_14974);
nor UO_1783 (O_1783,N_14919,N_14725);
or UO_1784 (O_1784,N_14890,N_14911);
nand UO_1785 (O_1785,N_14526,N_14905);
nor UO_1786 (O_1786,N_14881,N_14555);
nor UO_1787 (O_1787,N_14653,N_14647);
nor UO_1788 (O_1788,N_14608,N_14873);
and UO_1789 (O_1789,N_14424,N_14824);
or UO_1790 (O_1790,N_14535,N_14628);
nor UO_1791 (O_1791,N_14533,N_14636);
nand UO_1792 (O_1792,N_14613,N_14993);
nor UO_1793 (O_1793,N_14501,N_14627);
nand UO_1794 (O_1794,N_14924,N_14996);
nor UO_1795 (O_1795,N_14789,N_14666);
and UO_1796 (O_1796,N_14297,N_14647);
and UO_1797 (O_1797,N_14482,N_14769);
and UO_1798 (O_1798,N_14608,N_14320);
nand UO_1799 (O_1799,N_14847,N_14333);
or UO_1800 (O_1800,N_14269,N_14867);
and UO_1801 (O_1801,N_14347,N_14300);
and UO_1802 (O_1802,N_14727,N_14638);
or UO_1803 (O_1803,N_14879,N_14577);
nand UO_1804 (O_1804,N_14460,N_14602);
or UO_1805 (O_1805,N_14452,N_14621);
nor UO_1806 (O_1806,N_14602,N_14857);
or UO_1807 (O_1807,N_14949,N_14563);
or UO_1808 (O_1808,N_14475,N_14502);
and UO_1809 (O_1809,N_14801,N_14772);
and UO_1810 (O_1810,N_14697,N_14691);
nor UO_1811 (O_1811,N_14440,N_14392);
nand UO_1812 (O_1812,N_14910,N_14405);
or UO_1813 (O_1813,N_14421,N_14899);
nor UO_1814 (O_1814,N_14683,N_14590);
or UO_1815 (O_1815,N_14738,N_14271);
or UO_1816 (O_1816,N_14469,N_14719);
nor UO_1817 (O_1817,N_14733,N_14690);
nor UO_1818 (O_1818,N_14310,N_14270);
and UO_1819 (O_1819,N_14275,N_14527);
nor UO_1820 (O_1820,N_14555,N_14531);
nand UO_1821 (O_1821,N_14267,N_14947);
and UO_1822 (O_1822,N_14930,N_14589);
nor UO_1823 (O_1823,N_14699,N_14771);
nor UO_1824 (O_1824,N_14727,N_14893);
nand UO_1825 (O_1825,N_14780,N_14849);
nor UO_1826 (O_1826,N_14675,N_14343);
nor UO_1827 (O_1827,N_14734,N_14961);
and UO_1828 (O_1828,N_14819,N_14751);
nor UO_1829 (O_1829,N_14320,N_14950);
or UO_1830 (O_1830,N_14801,N_14993);
or UO_1831 (O_1831,N_14755,N_14481);
or UO_1832 (O_1832,N_14783,N_14858);
nand UO_1833 (O_1833,N_14836,N_14860);
nor UO_1834 (O_1834,N_14519,N_14317);
and UO_1835 (O_1835,N_14742,N_14875);
nand UO_1836 (O_1836,N_14343,N_14507);
nor UO_1837 (O_1837,N_14596,N_14744);
nand UO_1838 (O_1838,N_14598,N_14638);
or UO_1839 (O_1839,N_14991,N_14851);
nand UO_1840 (O_1840,N_14376,N_14386);
nand UO_1841 (O_1841,N_14665,N_14958);
and UO_1842 (O_1842,N_14744,N_14466);
or UO_1843 (O_1843,N_14873,N_14761);
nand UO_1844 (O_1844,N_14524,N_14660);
and UO_1845 (O_1845,N_14856,N_14251);
nand UO_1846 (O_1846,N_14466,N_14768);
or UO_1847 (O_1847,N_14972,N_14282);
or UO_1848 (O_1848,N_14910,N_14351);
nand UO_1849 (O_1849,N_14319,N_14876);
and UO_1850 (O_1850,N_14649,N_14866);
nand UO_1851 (O_1851,N_14872,N_14369);
or UO_1852 (O_1852,N_14639,N_14958);
and UO_1853 (O_1853,N_14461,N_14528);
nor UO_1854 (O_1854,N_14800,N_14842);
nand UO_1855 (O_1855,N_14534,N_14728);
nand UO_1856 (O_1856,N_14755,N_14304);
nand UO_1857 (O_1857,N_14885,N_14298);
nor UO_1858 (O_1858,N_14697,N_14532);
nand UO_1859 (O_1859,N_14608,N_14569);
nand UO_1860 (O_1860,N_14300,N_14955);
or UO_1861 (O_1861,N_14926,N_14728);
or UO_1862 (O_1862,N_14895,N_14994);
nor UO_1863 (O_1863,N_14862,N_14451);
nand UO_1864 (O_1864,N_14258,N_14289);
or UO_1865 (O_1865,N_14524,N_14446);
nor UO_1866 (O_1866,N_14390,N_14987);
or UO_1867 (O_1867,N_14978,N_14461);
and UO_1868 (O_1868,N_14650,N_14720);
nor UO_1869 (O_1869,N_14267,N_14989);
or UO_1870 (O_1870,N_14575,N_14983);
nor UO_1871 (O_1871,N_14410,N_14467);
or UO_1872 (O_1872,N_14504,N_14283);
nor UO_1873 (O_1873,N_14727,N_14359);
nand UO_1874 (O_1874,N_14900,N_14720);
or UO_1875 (O_1875,N_14915,N_14355);
nor UO_1876 (O_1876,N_14261,N_14720);
nor UO_1877 (O_1877,N_14560,N_14982);
nand UO_1878 (O_1878,N_14866,N_14363);
nor UO_1879 (O_1879,N_14890,N_14539);
nor UO_1880 (O_1880,N_14357,N_14789);
and UO_1881 (O_1881,N_14469,N_14437);
or UO_1882 (O_1882,N_14284,N_14844);
nor UO_1883 (O_1883,N_14394,N_14797);
and UO_1884 (O_1884,N_14873,N_14717);
and UO_1885 (O_1885,N_14482,N_14384);
and UO_1886 (O_1886,N_14575,N_14724);
or UO_1887 (O_1887,N_14605,N_14450);
nor UO_1888 (O_1888,N_14756,N_14918);
and UO_1889 (O_1889,N_14258,N_14692);
nand UO_1890 (O_1890,N_14999,N_14367);
or UO_1891 (O_1891,N_14891,N_14288);
nand UO_1892 (O_1892,N_14819,N_14985);
nor UO_1893 (O_1893,N_14574,N_14636);
nor UO_1894 (O_1894,N_14845,N_14453);
xor UO_1895 (O_1895,N_14913,N_14270);
nor UO_1896 (O_1896,N_14707,N_14527);
nand UO_1897 (O_1897,N_14664,N_14437);
and UO_1898 (O_1898,N_14613,N_14702);
nand UO_1899 (O_1899,N_14904,N_14688);
or UO_1900 (O_1900,N_14469,N_14807);
or UO_1901 (O_1901,N_14308,N_14292);
nand UO_1902 (O_1902,N_14619,N_14252);
nor UO_1903 (O_1903,N_14552,N_14950);
or UO_1904 (O_1904,N_14781,N_14671);
nand UO_1905 (O_1905,N_14718,N_14348);
and UO_1906 (O_1906,N_14266,N_14814);
nand UO_1907 (O_1907,N_14882,N_14348);
nor UO_1908 (O_1908,N_14253,N_14588);
and UO_1909 (O_1909,N_14338,N_14503);
and UO_1910 (O_1910,N_14604,N_14845);
and UO_1911 (O_1911,N_14823,N_14415);
nor UO_1912 (O_1912,N_14443,N_14807);
nor UO_1913 (O_1913,N_14993,N_14343);
or UO_1914 (O_1914,N_14495,N_14349);
nor UO_1915 (O_1915,N_14330,N_14523);
nand UO_1916 (O_1916,N_14630,N_14929);
nand UO_1917 (O_1917,N_14272,N_14406);
nor UO_1918 (O_1918,N_14490,N_14319);
and UO_1919 (O_1919,N_14407,N_14934);
and UO_1920 (O_1920,N_14977,N_14749);
or UO_1921 (O_1921,N_14277,N_14648);
nand UO_1922 (O_1922,N_14779,N_14352);
nor UO_1923 (O_1923,N_14503,N_14406);
nand UO_1924 (O_1924,N_14726,N_14587);
nand UO_1925 (O_1925,N_14351,N_14427);
nor UO_1926 (O_1926,N_14417,N_14671);
and UO_1927 (O_1927,N_14506,N_14417);
or UO_1928 (O_1928,N_14720,N_14822);
nand UO_1929 (O_1929,N_14557,N_14477);
and UO_1930 (O_1930,N_14773,N_14675);
nand UO_1931 (O_1931,N_14342,N_14979);
nand UO_1932 (O_1932,N_14981,N_14300);
nor UO_1933 (O_1933,N_14618,N_14347);
nor UO_1934 (O_1934,N_14447,N_14882);
or UO_1935 (O_1935,N_14997,N_14825);
or UO_1936 (O_1936,N_14555,N_14680);
nor UO_1937 (O_1937,N_14593,N_14906);
nor UO_1938 (O_1938,N_14275,N_14769);
or UO_1939 (O_1939,N_14272,N_14427);
or UO_1940 (O_1940,N_14483,N_14944);
or UO_1941 (O_1941,N_14601,N_14586);
nor UO_1942 (O_1942,N_14620,N_14404);
nor UO_1943 (O_1943,N_14262,N_14699);
nor UO_1944 (O_1944,N_14528,N_14529);
nand UO_1945 (O_1945,N_14880,N_14673);
or UO_1946 (O_1946,N_14856,N_14694);
nand UO_1947 (O_1947,N_14501,N_14522);
or UO_1948 (O_1948,N_14401,N_14472);
nor UO_1949 (O_1949,N_14783,N_14330);
and UO_1950 (O_1950,N_14462,N_14398);
and UO_1951 (O_1951,N_14984,N_14465);
or UO_1952 (O_1952,N_14860,N_14259);
or UO_1953 (O_1953,N_14652,N_14477);
and UO_1954 (O_1954,N_14840,N_14718);
nand UO_1955 (O_1955,N_14630,N_14295);
nor UO_1956 (O_1956,N_14717,N_14854);
and UO_1957 (O_1957,N_14529,N_14959);
nand UO_1958 (O_1958,N_14753,N_14359);
nand UO_1959 (O_1959,N_14848,N_14739);
or UO_1960 (O_1960,N_14447,N_14412);
nor UO_1961 (O_1961,N_14482,N_14380);
or UO_1962 (O_1962,N_14495,N_14471);
nor UO_1963 (O_1963,N_14683,N_14252);
or UO_1964 (O_1964,N_14586,N_14276);
nor UO_1965 (O_1965,N_14567,N_14471);
or UO_1966 (O_1966,N_14377,N_14464);
nor UO_1967 (O_1967,N_14695,N_14307);
nand UO_1968 (O_1968,N_14685,N_14548);
and UO_1969 (O_1969,N_14747,N_14913);
and UO_1970 (O_1970,N_14978,N_14840);
and UO_1971 (O_1971,N_14624,N_14285);
or UO_1972 (O_1972,N_14566,N_14785);
and UO_1973 (O_1973,N_14282,N_14879);
and UO_1974 (O_1974,N_14960,N_14673);
and UO_1975 (O_1975,N_14861,N_14895);
or UO_1976 (O_1976,N_14751,N_14879);
or UO_1977 (O_1977,N_14762,N_14800);
nand UO_1978 (O_1978,N_14543,N_14954);
or UO_1979 (O_1979,N_14507,N_14367);
and UO_1980 (O_1980,N_14268,N_14943);
nor UO_1981 (O_1981,N_14395,N_14521);
and UO_1982 (O_1982,N_14881,N_14509);
nor UO_1983 (O_1983,N_14453,N_14837);
and UO_1984 (O_1984,N_14908,N_14508);
nand UO_1985 (O_1985,N_14900,N_14610);
and UO_1986 (O_1986,N_14835,N_14760);
nor UO_1987 (O_1987,N_14462,N_14422);
nand UO_1988 (O_1988,N_14839,N_14553);
nor UO_1989 (O_1989,N_14408,N_14625);
nand UO_1990 (O_1990,N_14329,N_14448);
or UO_1991 (O_1991,N_14881,N_14941);
nor UO_1992 (O_1992,N_14919,N_14969);
nand UO_1993 (O_1993,N_14621,N_14333);
and UO_1994 (O_1994,N_14466,N_14482);
nand UO_1995 (O_1995,N_14771,N_14451);
nor UO_1996 (O_1996,N_14902,N_14767);
nand UO_1997 (O_1997,N_14758,N_14533);
nand UO_1998 (O_1998,N_14740,N_14388);
or UO_1999 (O_1999,N_14608,N_14947);
endmodule